magic
tech sky130A
magscale 1 2
timestamp 1628437904
<< nwell >>
rect -512 1248 2 1760
<< pwell >>
rect -490 670 -12 1094
<< nmos >>
rect -216 678 -186 1078
rect -122 678 -92 1078
<< pmos >>
rect -216 1298 -186 1698
rect -122 1298 -92 1698
<< ndiff >>
rect -274 1066 -216 1078
rect -274 690 -262 1066
rect -228 690 -216 1066
rect -274 678 -216 690
rect -186 1066 -122 1078
rect -186 690 -168 1066
rect -134 690 -122 1066
rect -186 678 -122 690
rect -92 1066 -34 1078
rect -92 690 -80 1066
rect -46 690 -34 1066
rect -92 678 -34 690
<< pdiff >>
rect -274 1686 -216 1698
rect -274 1310 -262 1686
rect -228 1310 -216 1686
rect -274 1298 -216 1310
rect -186 1686 -122 1698
rect -186 1310 -168 1686
rect -134 1310 -122 1686
rect -186 1298 -122 1310
rect -92 1686 -34 1698
rect -92 1310 -80 1686
rect -46 1310 -34 1686
rect -92 1298 -34 1310
<< ndiffc >>
rect -262 690 -228 1066
rect -168 690 -134 1066
rect -80 690 -46 1066
<< pdiffc >>
rect -262 1310 -228 1686
rect -168 1310 -134 1686
rect -80 1310 -46 1686
<< psubdiffcont >>
rect -454 766 -360 980
<< nsubdiffcont >>
rect -436 1392 -360 1598
<< poly >>
rect -216 1698 -186 1724
rect -122 1698 -92 1724
rect -216 1264 -186 1298
rect -302 1250 -186 1264
rect -302 1218 -284 1250
rect -226 1218 -186 1250
rect -302 1206 -186 1218
rect -216 1078 -186 1206
rect -122 1178 -92 1298
rect -144 1164 -50 1178
rect -144 1132 -126 1164
rect -68 1132 -50 1164
rect -144 1120 -50 1132
rect -122 1078 -92 1120
rect -216 652 -186 678
rect -122 652 -92 678
<< polycont >>
rect -284 1218 -226 1250
rect -126 1132 -68 1164
<< locali >>
rect -262 1686 -228 1702
rect -454 1598 -340 1620
rect -454 1392 -436 1598
rect -360 1392 -340 1598
rect -454 1374 -340 1392
rect -262 1294 -228 1310
rect -174 1686 -134 1702
rect -174 1310 -168 1686
rect -174 1294 -134 1310
rect -80 1686 -46 1702
rect -80 1294 -46 1310
rect -300 1218 -294 1252
rect -220 1218 -210 1252
rect -142 1132 -132 1166
rect -58 1132 -52 1166
rect -262 1066 -228 1082
rect -472 980 -344 1002
rect -472 766 -454 980
rect -360 766 -344 980
rect -472 750 -344 766
rect -262 674 -228 690
rect -174 1066 -134 1082
rect -174 690 -168 1066
rect -174 674 -134 690
rect -80 1066 -46 1082
rect -80 674 -46 690
<< viali >>
rect -436 1392 -360 1598
rect -262 1310 -228 1686
rect -168 1310 -134 1686
rect -80 1310 -46 1686
rect -294 1250 -220 1258
rect -294 1218 -284 1250
rect -284 1218 -226 1250
rect -226 1218 -220 1250
rect -294 1212 -220 1218
rect -132 1164 -58 1172
rect -132 1132 -126 1164
rect -126 1132 -68 1164
rect -68 1132 -58 1164
rect -132 1126 -58 1132
rect -454 766 -360 980
rect -262 690 -228 1066
rect -168 690 -134 1066
rect -80 690 -46 1066
<< metal1 >>
rect -284 1842 -274 1866
rect -414 1792 -274 1842
rect -204 1792 -194 1866
rect -102 1792 -92 1866
rect -22 1792 -12 1866
rect -414 1790 -222 1792
rect -102 1790 -40 1792
rect -414 1610 -374 1790
rect -268 1686 -222 1790
rect -442 1598 -354 1610
rect -442 1392 -436 1598
rect -360 1392 -354 1598
rect -442 1380 -354 1392
rect -268 1310 -262 1686
rect -228 1310 -222 1686
rect -268 1298 -222 1310
rect -180 1686 -128 1698
rect -180 1310 -168 1686
rect -134 1310 -128 1686
rect -306 1258 -208 1264
rect -306 1212 -294 1258
rect -220 1212 -208 1258
rect -180 1258 -128 1310
rect -86 1686 -40 1790
rect -86 1310 -80 1686
rect -46 1310 -40 1686
rect -86 1298 -40 1310
rect -180 1218 18 1258
rect -306 1206 -208 1212
rect -144 1172 -46 1178
rect -144 1126 -132 1172
rect -58 1126 -46 1172
rect -144 1120 -46 1126
rect -18 1078 18 1218
rect -268 1066 -222 1078
rect -460 980 -354 992
rect -460 766 -454 980
rect -360 766 -354 980
rect -460 754 -354 766
rect -432 634 -372 754
rect -268 690 -262 1066
rect -228 690 -222 1066
rect -268 638 -222 690
rect -180 1066 -128 1078
rect -180 690 -168 1066
rect -134 690 -128 1066
rect -180 678 -128 690
rect -86 1066 18 1078
rect -86 690 -80 1066
rect -46 1038 18 1066
rect -46 690 -40 1038
rect -86 678 -40 690
rect -288 634 -278 638
rect -432 570 -278 634
rect -288 552 -278 570
rect -194 552 -184 638
<< via1 >>
rect -274 1792 -204 1866
rect -92 1792 -22 1866
rect -278 552 -194 638
<< metal2 >>
rect -280 1872 -196 1882
rect -280 1776 -196 1786
rect -98 1872 -14 1882
rect -98 1776 -14 1786
rect -278 638 -194 648
rect -278 542 -194 552
<< via2 >>
rect -280 1866 -196 1872
rect -280 1792 -274 1866
rect -274 1792 -204 1866
rect -204 1792 -196 1866
rect -280 1786 -196 1792
rect -98 1866 -14 1872
rect -98 1792 -92 1866
rect -92 1792 -22 1866
rect -22 1792 -14 1866
rect -98 1786 -14 1792
rect -278 552 -194 638
<< metal3 >>
rect -290 1872 -186 1877
rect -290 1786 -280 1872
rect -196 1786 -186 1872
rect -290 1781 -186 1786
rect -108 1872 -4 1877
rect -108 1786 -98 1872
rect -14 1786 -4 1872
rect -108 1781 -4 1786
rect -288 638 -184 643
rect -288 552 -278 638
rect -194 552 -184 638
rect -288 547 -184 552
<< via3 >>
rect -280 1786 -196 1872
rect -98 1786 -14 1872
rect -278 552 -194 638
<< metal4 >>
rect -286 1872 -4 1882
rect -286 1786 -280 1872
rect -196 1786 -98 1872
rect -14 1786 -4 1872
rect -286 1778 -4 1786
rect -288 638 -18 648
rect -288 552 -278 638
rect -194 552 -18 638
rect -288 544 -18 552
<< labels >>
flabel metal4 -166 1838 -166 1838 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal4 -88 570 -88 570 0 FreeSans 1600 0 0 0 vss
port 4 nsew
flabel metal1 4 1174 4 1174 0 FreeSans 1600 0 0 0 out
port 3 nsew
flabel viali -112 1146 -112 1146 0 FreeSans 1600 0 0 0 A
port 2 nsew
flabel viali -270 1226 -270 1226 0 FreeSans 1600 0 0 0 B
port 1 nsew
<< end >>
