* NGSPICE file created from floor_plan.ext - technology: sky130A


* Top level circuit floor_plan

X0 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2 a_677477_25371# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4 a_677477_25371# a_673159_24981# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X11 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X12 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X15 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X16 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X17 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X20 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X21 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X22 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X23 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X24 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X25 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X26 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X27 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X28 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X29 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X30 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X31 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X32 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X33 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X34 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X35 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X36 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X37 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X38 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X39 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X40 w_692190_39881# a_664155_35747# a_692386_37781# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X41 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X42 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X43 a_677477_25371# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X44 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X45 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X46 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X47 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X48 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X49 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X50 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X51 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X52 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X53 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X54 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X55 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X56 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X57 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X58 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X59 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X60 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X61 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X62 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X63 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X64 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X65 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X66 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X67 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X68 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X69 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X70 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X71 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X72 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X73 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X74 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X75 w_719104_5922# a_719858_6024# a_722600_2050# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X76 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X77 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X78 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X79 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X80 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X81 a_725512_82134# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X82 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X83 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X84 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X85 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X86 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X87 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X88 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X89 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X90 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X91 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X92 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X93 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X94 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X95 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X96 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X97 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X98 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X99 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X100 w_693353_20554# a_682038_37869# a_693549_25370# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X101 w_649931_37947# a_693549_25370# a_694493_20773# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X102 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X103 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X104 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X105 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X106 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X107 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X108 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X109 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X110 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X111 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X112 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X113 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X114 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X115 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X116 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X117 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X118 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X119 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X120 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X121 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X122 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X123 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X124 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X125 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X126 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X127 a_719858_78562# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X128 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X129 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X130 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X131 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X132 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X133 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X134 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X135 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X136 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X137 a_725512_8976# a_719900_5846# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X138 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X139 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X140 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X141 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X142 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X143 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X144 w_649931_37947# a_693549_25370# a_694493_20773# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X145 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X146 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X147 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X148 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X149 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X150 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X151 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X152 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X153 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X154 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X155 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X156 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X157 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X158 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X159 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X160 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X161 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X162 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X163 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X164 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X165 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X166 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X167 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X168 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X169 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X170 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X171 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X172 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X173 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X174 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X175 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X176 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X177 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X178 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X179 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X180 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X181 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X182 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X183 a_679806_37869# a_682459_41330# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=1.4e+06u
X184 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X185 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X186 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X187 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X188 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X189 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X190 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X191 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X192 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X193 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X194 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X195 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X196 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X197 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X198 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X199 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X200 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X201 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X202 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X203 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X204 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X205 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X206 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X207 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X208 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X209 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X210 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X211 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X212 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X213 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X214 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X215 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X216 w_693353_61507# a_682038_37869# a_693549_59407# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X217 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X218 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X219 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X220 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X221 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X222 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X223 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X224 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X225 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X226 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X227 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X228 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X229 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X230 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X231 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X232 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X233 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X234 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X235 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X236 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X237 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X238 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X239 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X240 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X241 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X242 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X243 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X244 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X245 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X246 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X247 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X248 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X249 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X250 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X251 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X252 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X253 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X254 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X255 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X256 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X257 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X258 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X259 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X260 a_664355_46657# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X261 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X262 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X263 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X264 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X265 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X266 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X267 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X268 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X269 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X270 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X271 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X272 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X273 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X274 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X275 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X276 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X277 w_677281_61507# a_664155_35747# a_678421_59495# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X278 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X279 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X280 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X281 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X282 w_649931_37947# a_677477_59407# a_677477_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X283 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X284 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X285 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X286 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X287 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X288 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X289 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X290 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X291 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X292 a_677477_59407# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X293 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X294 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X295 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X296 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X297 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X298 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X299 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X300 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X301 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X302 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X303 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X304 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X305 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X306 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X307 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X308 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X309 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X310 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X311 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X312 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X313 a_693549_59407# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X314 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X315 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X316 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X317 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X318 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X319 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X320 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X321 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X322 w_649931_37947# a_663411_33525# a_664355_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X323 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X324 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X325 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X326 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X327 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X328 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X329 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X330 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X331 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X332 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X333 a_675258_42633# a_676490_42315# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X334 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X335 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X336 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X337 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X338 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X339 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X340 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X341 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X342 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X343 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X344 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X345 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X346 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X347 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X348 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X349 w_649931_37947# a_663411_33525# a_664355_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X350 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X351 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X352 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X353 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X354 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X355 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X356 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X357 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X358 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X359 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X360 a_650141_38543# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X361 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X362 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X363 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X364 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X365 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X366 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X367 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X368 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X369 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X370 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X371 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X372 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X373 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X374 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X375 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X376 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X377 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X378 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X379 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X380 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X381 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X382 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X383 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X384 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X385 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X386 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X387 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X388 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X389 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X390 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X391 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X392 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X393 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X394 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X395 w_678666_39881# a_676490_44223# a_678862_37781# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X396 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X397 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X398 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X399 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X400 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X401 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X402 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X403 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X404 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X405 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X406 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X407 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X408 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X409 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X410 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X411 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X412 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X413 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X414 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X415 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X416 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X417 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X418 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X419 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X420 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X421 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X422 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X423 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X424 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X425 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X426 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X427 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X428 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X429 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X430 a_678421_20774# a_664155_35747# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X431 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X432 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X433 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X434 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X435 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X436 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X437 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X438 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X439 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X440 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X441 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X442 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X443 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X444 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X445 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X446 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X447 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X448 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X449 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X450 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X451 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X452 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X453 a_692386_37781# a_664155_35747# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X454 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X455 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X456 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X457 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X458 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X459 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X460 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X461 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X462 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X463 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X464 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X465 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X466 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X467 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X468 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X469 a_677477_59407# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X470 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X471 w_649931_37947# a_677477_59407# a_678421_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X472 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X473 a_719858_80608# a_719332_79990# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X474 w_649931_37947# a_650053_38143# a_650141_46551# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X475 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X476 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X477 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X478 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X479 w_649931_37947# a_677477_25371# a_678421_20774# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X480 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X481 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X482 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X483 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X484 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X485 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X486 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X487 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X488 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X489 w_649931_37947# a_693549_59407# a_694493_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X490 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X491 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X492 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X493 a_650141_44263# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X494 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X495 a_694493_59495# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X496 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X497 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X498 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X499 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X500 a_719742_79090# a_722600_82134# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X501 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X502 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X503 a_693549_59407# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X504 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X505 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X506 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X507 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X508 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X509 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X510 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X511 a_663411_33525# a_662413_39580# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X512 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X513 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X514 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X515 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X516 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X517 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X518 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X519 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X520 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X521 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X522 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X523 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X524 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X525 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X526 a_725512_8976# a_719900_5846# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X527 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X528 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X529 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X530 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X531 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X532 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X533 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X534 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X535 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X536 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X537 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X538 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X539 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X540 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X541 a_650053_38143# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X542 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X543 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X544 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X545 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X546 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X547 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X548 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X549 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X550 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X551 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X552 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X553 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X554 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X555 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X556 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X557 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X558 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X559 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X560 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X561 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X562 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X563 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X564 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X565 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X566 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X567 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X568 a_664355_46657# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X569 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X570 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X571 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X572 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X573 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X574 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X575 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X576 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X577 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X578 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X579 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X580 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X581 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X582 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X583 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X584 w_663215_35625# a_664155_35747# a_664355_33613# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X585 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X586 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X587 a_678421_20774# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X588 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X589 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X590 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X591 w_649931_37947# a_719742_79090# a_725512_82134# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X592 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X593 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X594 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X595 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X596 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X597 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X598 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X599 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X600 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X601 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X602 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X603 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X604 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X605 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X606 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X607 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X608 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X609 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X610 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X611 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X612 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X613 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X614 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X615 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X616 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X617 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X618 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X619 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X620 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X621 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X622 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X623 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X624 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X625 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X626 w_692190_39881# a_693130_40003# a_693330_37869# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X627 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X628 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X629 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X630 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X631 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X632 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X633 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X634 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X635 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X636 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X637 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X638 a_675315_85767# a_674997_87199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X639 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X640 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X641 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X642 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X643 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X644 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X645 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X646 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X647 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X648 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X649 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X650 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X651 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X652 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X653 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X654 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X655 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X656 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X657 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X658 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X659 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X660 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X661 w_677281_20555# a_673159_24981# a_677477_25371# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X662 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X663 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X664 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X665 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X666 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X667 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X668 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X669 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X670 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X671 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X672 a_725512_8976# a_719900_5846# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X673 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X674 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X675 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X676 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X677 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X678 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X679 w_649931_37947# a_719900_80508# a_725512_73584# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X680 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X681 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X682 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X683 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X684 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X685 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X686 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X687 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X688 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X689 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X690 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X691 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X692 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X693 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X694 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X695 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X696 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X697 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X698 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X699 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X700 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X701 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X702 a_693549_25370# a_682038_37869# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X703 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X704 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X705 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X706 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X707 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X708 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X709 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X710 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X711 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X712 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X713 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X714 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X715 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X716 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X717 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X718 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X719 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X720 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X721 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X722 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X723 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X724 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X725 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X726 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X727 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X728 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X729 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X730 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X731 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X732 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X733 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X734 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X735 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X736 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X737 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X738 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X739 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X740 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X741 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X742 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X743 w_649931_37947# a_678862_37781# a_678862_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X744 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X745 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X746 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X747 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X748 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X749 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X750 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X751 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X752 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X753 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X754 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X755 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X756 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X757 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X758 w_649931_37947# a_663411_51254# a_663411_51254# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X759 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X760 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X761 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X762 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X763 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X764 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X765 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X766 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X767 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X768 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X769 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X770 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X771 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X772 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X773 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X774 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X775 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X776 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X777 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X778 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X779 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X780 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X781 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X782 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X783 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X784 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X785 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X786 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X787 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X788 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X789 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X790 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X791 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X792 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X793 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X794 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X795 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X796 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X797 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X798 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X799 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X800 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X801 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X802 a_677477_25371# a_673159_24981# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X803 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X804 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X805 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X806 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X807 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X808 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X809 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X810 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X811 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X812 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X813 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X814 a_693549_59407# a_682038_37869# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X815 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X816 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X817 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X818 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X819 w_649931_37947# a_693549_59407# a_693549_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X820 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X821 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X822 a_682038_37869# a_693130_40003# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X823 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X824 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X825 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X826 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X827 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X828 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X829 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X830 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X831 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X832 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X833 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X834 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X835 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X836 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X837 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X838 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X839 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X840 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X841 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X842 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X843 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X844 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X845 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X846 w_678666_39881# a_676490_44223# a_678862_37781# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X847 a_677477_25371# a_673159_24981# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X848 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X849 a_679806_37869# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X850 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X851 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X852 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X853 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X854 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X855 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X856 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X857 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X858 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X859 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X860 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X861 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X862 w_649931_37947# a_677477_59407# a_677477_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X863 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X864 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X865 a_650141_47695# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X866 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X867 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X868 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X869 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X870 a_693549_25370# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X871 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X872 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X873 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X874 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X875 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X876 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X877 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X878 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X879 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X880 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X881 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X882 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X883 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X884 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X885 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X886 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X887 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X888 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X889 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X890 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X891 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X892 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X893 a_719742_79090# a_722600_82134# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X894 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X895 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X896 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X897 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X898 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X899 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X900 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X901 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X902 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X903 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X904 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X905 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X906 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X907 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X908 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X909 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X910 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X911 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X912 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X913 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X914 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X915 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X916 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X917 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X918 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X919 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X920 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X921 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X922 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X923 w_649931_37947# a_650053_38143# a_650141_39687# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X924 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X925 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X926 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X927 w_649931_37947# a_677477_59407# a_678421_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X928 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X929 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X930 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X931 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X932 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X933 a_675633_n1233# a_675951_199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X934 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X935 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X936 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X937 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X938 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X939 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X940 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X941 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X942 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X943 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X944 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X945 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X946 w_693353_20554# a_680653_25459# a_694493_20773# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X947 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X948 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X949 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X950 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X951 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X952 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X953 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X954 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X955 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X956 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X957 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X958 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X959 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X960 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X961 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X962 w_719104_5922# a_722600_75208# a_719900_80508# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X963 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X964 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X965 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X966 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X967 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X968 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X969 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X970 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X971 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X972 a_693330_37869# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X973 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X974 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X975 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X976 w_677281_20555# a_664155_35747# a_678421_20774# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X977 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X978 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X979 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X980 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X981 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X982 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X983 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X984 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X985 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X986 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X987 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X988 a_679806_37869# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X989 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X990 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X991 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X992 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X993 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X994 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X995 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X996 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X997 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X998 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X999 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1000 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1001 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1002 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1003 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1004 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X1005 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1006 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1007 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1008 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1009 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1010 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1011 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1012 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1013 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1014 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1015 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1016 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1017 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1018 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1019 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1020 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1021 w_649931_37947# a_719900_5846# a_725512_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1022 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1023 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1024 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1025 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1026 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1027 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1028 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1029 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1030 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1031 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1032 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1033 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1034 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1035 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1036 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1037 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1038 w_649931_37947# a_722600_8976# a_719900_5846# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1039 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1040 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1041 a_677477_59407# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1042 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1043 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1044 w_693353_61507# a_680653_59495# a_694493_59495# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1045 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1046 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1047 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1048 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1049 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1050 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1051 w_649931_37947# a_722600_2050# a_719742_7264# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1052 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1053 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1054 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1055 a_693549_59407# a_682038_37869# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1056 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1057 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1058 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1059 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1060 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1061 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1062 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1063 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1064 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1065 a_694493_59495# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1066 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1067 a_694493_20773# a_680653_25459# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1068 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1069 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1070 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1071 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1072 a_664355_33613# a_664155_35747# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1073 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1074 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1075 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1076 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1077 a_693330_37869# a_693130_40003# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1078 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1079 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1080 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1081 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1082 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1083 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1084 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1085 a_725512_82134# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1086 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1087 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1088 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1089 w_663215_35625# a_664155_35747# a_664355_33613# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1090 a_679806_37869# a_664155_35747# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1091 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1092 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1093 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1094 w_649931_37947# a_678862_37781# a_679806_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1095 w_719104_5922# a_696725_59495# a_719858_79182# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1096 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1097 w_663215_46438# a_663411_46560# a_663411_51254# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1098 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1099 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1100 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1101 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1102 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1103 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1104 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1105 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1106 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1107 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1108 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1109 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1110 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1111 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1112 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1113 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1114 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1115 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1116 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1117 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1118 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X1119 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1120 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1121 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1122 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1123 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1124 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1125 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1126 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1127 w_719104_5922# a_722600_8976# a_719900_5846# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1128 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1129 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1130 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1131 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1132 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1133 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1134 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1135 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1136 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1137 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1138 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1139 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1140 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1141 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1142 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1143 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1144 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1145 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1146 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1147 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1148 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1149 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1150 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1151 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1152 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1153 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1154 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1155 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1156 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1157 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1158 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1159 a_725512_73584# a_719900_80508# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1160 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1161 w_677281_61507# a_673159_61357# a_677477_59407# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1162 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1163 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1164 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1165 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1166 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1167 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1168 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1169 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1170 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1171 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1172 a_693549_25370# a_682038_37869# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1173 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1174 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1175 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1176 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1177 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1178 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1179 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1180 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1181 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1182 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1183 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1184 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1185 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1186 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1187 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1188 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1189 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1190 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1191 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1192 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1193 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1194 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1195 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1196 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1197 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1198 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1199 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1200 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1201 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1202 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1203 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1204 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1205 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1206 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1207 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1208 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1209 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1210 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1211 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1212 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1213 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1214 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1215 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1216 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1217 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1218 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1219 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1220 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1221 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1222 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1223 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1224 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1225 a_676490_44223# a_682038_37869# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X1226 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1227 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1228 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1229 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1230 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1231 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1232 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1233 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1234 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1235 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1236 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1237 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1238 w_693353_61507# a_680653_59495# a_694493_59495# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1239 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1240 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1241 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1242 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1243 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1244 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1245 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1246 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1247 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1248 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1249 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1250 w_649931_37947# a_650053_38143# a_650141_38543# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1251 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1252 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1253 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1254 w_693353_20554# a_682038_37869# a_693549_25370# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1255 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1256 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1257 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1258 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1259 w_649931_37947# a_663411_51254# a_664355_46657# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1260 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1261 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1262 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1263 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1264 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1265 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1266 a_694493_20773# a_680653_25459# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1267 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1268 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1269 w_649931_37947# a_650053_38143# a_650141_41975# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1270 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1271 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1272 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1273 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1274 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1275 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1276 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1277 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1278 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1279 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1280 w_649931_37947# a_663411_51254# a_664355_46657# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1281 a_663411_51254# a_663411_46560# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1282 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1283 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1284 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1285 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1286 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1287 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1288 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1289 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1290 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1291 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1292 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1293 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1294 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1295 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1296 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1297 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1298 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1299 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1300 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1301 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1302 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1303 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1304 a_719900_5846# a_722600_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1305 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1306 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1307 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1308 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1309 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1310 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1311 w_719104_5922# a_722600_2050# a_719742_7264# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1312 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1313 a_675258_43269# a_676490_43587# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X1314 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1315 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1316 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1317 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1318 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1319 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1320 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1321 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1322 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1323 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1324 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1325 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1326 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1327 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1328 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1329 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1330 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1331 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1332 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1333 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1334 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1335 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1336 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1337 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1338 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1339 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1340 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1341 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1342 a_664355_33613# a_664155_35747# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1343 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1344 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1345 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1346 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1347 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1348 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1349 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1350 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1351 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1352 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1353 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1354 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1355 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1356 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1357 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1358 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1359 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1360 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1361 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1362 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1363 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1364 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1365 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1366 a_677477_59407# a_673159_61357# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1367 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1368 w_649931_37947# a_663411_33525# a_663411_33525# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1369 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1370 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1371 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1372 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1373 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1374 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1375 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1376 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1377 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1378 w_693353_20554# a_680653_25459# a_694493_20773# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1379 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1380 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1381 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1382 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1383 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1384 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1385 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1386 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1387 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1388 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1389 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1390 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1391 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1392 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1393 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1394 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1395 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1396 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1397 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1398 a_694493_59495# a_680653_59495# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1399 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1400 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1401 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1402 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1403 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1404 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1405 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1406 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1407 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1408 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1409 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1410 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1411 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1412 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1413 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1414 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1415 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1416 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1417 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1418 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1419 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1420 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1421 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1422 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1423 a_650141_44263# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1424 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1425 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1426 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1427 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1428 a_681073_63341# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=3e+07u
X1429 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1430 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1431 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1432 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1433 w_692190_39881# a_693130_40003# a_693330_37869# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1434 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1435 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1436 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1437 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1438 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1439 a_678421_59495# a_664155_35747# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1440 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1441 a_678862_37781# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1442 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1443 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1444 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X1445 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X1446 w_649931_37947# a_722600_8976# a_719900_5846# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1447 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1448 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1449 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1450 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1451 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1452 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1453 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1454 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1455 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1456 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1457 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1458 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1459 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1460 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1461 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1462 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1463 a_694493_20773# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1464 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1465 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1466 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1467 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1468 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1469 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1470 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1471 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1472 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1473 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1474 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1475 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1476 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1477 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1478 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1479 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1480 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1481 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1482 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1483 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1484 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1485 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1486 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1487 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1488 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1489 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1490 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1491 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1492 a_725512_n974# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1493 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1494 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1495 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1496 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1497 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1498 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1499 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1500 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1501 a_673159_59449# a_663411_46560# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X1502 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1503 a_725512_82134# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1504 a_719742_7264# a_722600_2050# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1505 w_649931_37947# a_692386_37781# a_693330_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1506 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1507 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1508 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1509 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1510 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1511 a_693330_37869# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1512 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1513 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1514 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1515 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1516 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1517 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1518 a_719858_6830# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1519 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1520 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1521 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1522 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1523 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1524 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1525 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1526 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1527 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1528 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1529 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1530 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1531 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1532 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1533 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1534 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1535 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1536 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1537 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1538 a_725512_n974# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1539 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1540 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1541 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1542 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1543 a_673159_60721# a_674591_61039# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X1544 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1545 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1546 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1547 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1548 w_663215_35625# a_662413_39580# a_663411_33525# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1549 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1550 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1551 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1552 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1553 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1554 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1555 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1556 w_663215_46438# a_662095_39580# a_664355_46657# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1557 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1558 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1559 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1560 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1561 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1562 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1563 a_679806_37869# a_664155_35747# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1564 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1565 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1566 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1567 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1568 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1569 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1570 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1571 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1572 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1573 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1574 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1575 a_663411_33525# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1576 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1577 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1578 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1579 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1580 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1581 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1582 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1583 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1584 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1585 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1586 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1587 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1588 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1589 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1590 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1591 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1592 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1593 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1594 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1595 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1596 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1597 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1598 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1599 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1600 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1601 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1602 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1603 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1604 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1605 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1606 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1607 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1608 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1609 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1610 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1611 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1612 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1613 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1614 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1615 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1616 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X1617 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1618 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1619 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1620 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1621 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1622 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1623 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1624 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1625 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1626 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1627 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1628 a_664355_33613# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1629 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1630 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1631 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1632 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1633 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1634 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1635 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1636 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1637 a_673159_25935# a_674591_25617# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X1638 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1639 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1640 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1641 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1642 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1643 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1644 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1645 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1646 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1647 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1648 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1649 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1650 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1651 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1652 a_725512_82134# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1653 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1654 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1655 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1656 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1657 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1658 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1659 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1660 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1661 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1662 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1663 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1664 a_693549_59407# a_682038_37869# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1665 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1666 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1667 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1668 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1669 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1670 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1671 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1672 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1673 w_649931_37947# a_693549_59407# a_694493_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1674 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1675 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1676 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1677 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1678 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1679 w_649931_37947# a_693549_25370# a_693549_25370# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1680 a_650141_39687# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1681 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1682 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1683 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1684 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1685 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1686 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1687 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1688 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1689 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1690 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1691 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1692 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1693 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1694 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1695 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1696 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1697 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1698 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1699 w_678666_39881# a_676490_44223# a_678862_37781# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1700 w_692190_39881# a_664155_35747# a_692386_37781# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1701 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1702 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1703 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1704 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1705 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1706 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1707 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1708 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1709 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1710 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1711 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1712 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1713 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1714 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1715 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1716 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1717 w_677281_61507# a_664155_35747# a_678421_59495# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1718 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1719 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1720 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1721 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1722 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1723 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1724 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1725 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1726 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1727 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1728 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1729 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1730 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1731 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1732 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1733 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1734 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1735 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1736 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1737 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1738 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1739 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1740 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1741 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1742 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1743 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1744 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1745 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1746 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1747 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X1748 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1749 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1750 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1751 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1752 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1753 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1754 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1755 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1756 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1757 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1758 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1759 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1760 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1761 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1762 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1763 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1764 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1765 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1766 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1767 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1768 w_649931_37947# a_692386_37781# a_692386_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1769 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1770 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1771 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1772 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1773 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1774 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1775 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1776 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1777 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1778 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1779 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1780 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1781 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1782 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1783 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1784 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1785 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1786 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1787 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1788 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1789 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1790 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1791 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1792 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1793 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1794 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1795 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1796 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1797 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1798 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1799 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1800 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1801 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1802 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1803 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1804 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1805 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1806 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1807 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1808 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1809 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1810 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1811 w_649931_37947# a_650053_38143# a_650141_47695# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X1812 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1813 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1814 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1815 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1816 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1817 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1818 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1819 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1820 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1821 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X1822 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1823 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1824 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1825 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1826 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1827 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1828 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1829 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1830 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1831 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1832 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1833 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1834 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1835 w_678666_39881# a_664155_35747# a_679806_37869# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1836 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1837 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1838 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1839 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1840 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1841 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1842 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1843 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1844 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1845 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1846 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1847 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1848 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1849 a_664355_46657# a_662095_39580# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1850 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1851 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1852 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1853 w_649931_37947# a_663411_51254# a_663411_51254# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1854 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1855 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1856 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1857 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1858 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1859 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1860 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1861 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1862 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1863 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1864 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1865 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1866 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1867 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1868 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1869 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1870 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1871 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1872 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1873 a_678862_37781# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1874 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1875 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1876 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1877 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1878 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1879 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1880 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1881 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1882 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1883 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1884 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1885 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1886 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1887 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1888 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1889 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1890 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1891 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1892 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1893 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1894 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1895 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1896 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1897 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1898 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1899 a_719858_6024# a_719900_5846# a_719858_5404# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1900 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1901 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1902 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1903 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1904 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1905 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1906 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1907 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1908 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1909 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1910 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1911 a_663411_33525# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1912 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1913 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1914 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1915 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1916 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1917 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1918 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1919 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1920 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1921 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1922 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1923 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1924 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1925 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1926 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1927 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1928 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1929 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1930 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1931 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1932 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1933 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1934 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1935 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1936 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1937 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1938 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1939 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1940 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1941 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1942 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1943 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1944 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1945 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1946 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1947 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1948 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1949 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1950 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1951 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1952 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1953 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1954 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1955 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1956 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1957 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1958 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1959 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1960 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1961 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1962 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1963 a_693330_37869# a_693130_40003# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1964 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1965 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1966 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1967 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1968 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1969 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1970 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1971 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1972 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1973 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1974 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1975 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1976 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1977 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1978 a_679806_37869# a_664155_35747# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1979 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1980 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1981 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1982 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1983 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1984 a_676490_44223# a_682038_37869# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X1985 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1986 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1987 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1988 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1989 a_678862_37781# a_676490_44223# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1990 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1991 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1992 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1993 w_649931_37947# a_678862_37781# a_678862_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1994 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1995 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1996 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X1997 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X1998 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1999 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2000 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2001 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2002 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X2003 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2004 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2005 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2006 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2007 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2008 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2009 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2010 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2011 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2012 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2013 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2014 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2015 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2016 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2017 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2018 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2019 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2020 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2021 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2022 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2023 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2024 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2025 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2026 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2027 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2028 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2029 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2030 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2031 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2032 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2033 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2034 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2035 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2036 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2037 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2038 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2039 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2040 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2041 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2042 w_649931_37947# a_719742_79090# a_725512_82134# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2043 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2044 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2045 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2046 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2047 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2048 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2049 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2050 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2051 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2052 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2053 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2054 a_663411_51254# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2055 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2056 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2057 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2058 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2059 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2060 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2061 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2062 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2063 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2064 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2065 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2066 w_677281_61507# a_673159_61357# a_677477_59407# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2067 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2068 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2069 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2070 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2071 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2072 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2073 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2074 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2075 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2076 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2077 a_725512_n974# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2078 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2079 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2080 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2081 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2082 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2083 a_678421_59495# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2084 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2085 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2086 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2087 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2088 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2089 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2090 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2091 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2092 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2093 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2094 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2095 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2096 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2097 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2098 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2099 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2100 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2101 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2102 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2103 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2104 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2105 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2106 a_650141_40831# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2107 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2108 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2109 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2110 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2111 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2112 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2113 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2114 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2115 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2116 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2117 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2118 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2119 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2120 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2121 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2122 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2123 w_663215_46438# a_662095_39580# a_664355_46657# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2124 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2125 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2126 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2127 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2128 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2129 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2130 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2131 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2132 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2133 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2134 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2135 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2136 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2137 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2138 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2139 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2140 a_725512_8976# a_719900_5846# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2141 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2142 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2143 w_649931_37947# a_650053_38143# a_650141_45407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2144 w_649931_37947# a_663411_33525# a_664355_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2145 w_649931_37947# a_719900_80508# a_725512_73584# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2146 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2147 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2148 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2149 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2150 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2151 a_692386_37781# a_664155_35747# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2152 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2153 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2154 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2155 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2156 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2157 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2158 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2159 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2160 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2161 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2162 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2163 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2164 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2165 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2166 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2167 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2168 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2169 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2170 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2171 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2172 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2173 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2174 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2175 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2176 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2177 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2178 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2179 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2180 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2181 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2182 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2183 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2184 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2185 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2186 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2187 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2188 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2189 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2190 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2191 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2192 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2193 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2194 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2195 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2196 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2197 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2198 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2199 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2200 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2201 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2202 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2203 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2204 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2205 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2206 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2207 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2208 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2209 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2210 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2211 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2212 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2213 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2214 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2215 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2216 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2217 a_692386_37781# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2218 a_663411_33525# a_662413_39580# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2219 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2220 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2221 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2222 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2223 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2224 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2225 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2226 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2227 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2228 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2229 w_649931_37947# a_650053_38143# a_650053_38143# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2230 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2231 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2232 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2233 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2234 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2235 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2236 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2237 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2238 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2239 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2240 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2241 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2242 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2243 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2244 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2245 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2246 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2247 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2248 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2249 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2250 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2251 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2252 a_667251_37508# a_662413_39580# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X2253 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2254 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2255 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2256 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2257 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2258 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2259 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2260 a_693330_37869# a_693130_40003# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2261 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2262 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2263 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2264 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2265 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2266 w_719104_5922# a_719858_79988# a_722600_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2267 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2268 a_650141_45407# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2269 w_649931_37947# a_650053_38143# a_650141_38543# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2270 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2271 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2272 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2273 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2274 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2275 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2276 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2277 a_677477_59407# a_673159_61357# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2278 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2279 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2280 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2281 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2282 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2283 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2284 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2285 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2286 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2287 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2288 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2289 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2290 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2291 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2292 w_649931_37947# a_650053_38143# a_650141_41975# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2293 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2294 w_649931_37947# a_677477_25371# a_677477_25371# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2295 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2296 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2297 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2298 a_677477_25371# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2299 w_649931_37947# a_719900_80508# a_725512_73584# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2300 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2301 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2302 a_677477_25371# a_673159_24981# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2303 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2304 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2305 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2306 a_694493_59495# a_680653_59495# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2307 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2308 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2309 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2310 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2311 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2312 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2313 a_719858_6830# a_696725_25458# a_719858_7450# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2314 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2315 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2316 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2317 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2318 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2319 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2320 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2321 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2322 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2323 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2324 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2325 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2326 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2327 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2328 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2329 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2330 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2331 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2332 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2333 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2334 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2335 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2336 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2337 w_649931_37947# a_692386_37781# a_692386_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2338 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2339 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2340 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2341 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2342 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2343 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2344 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2345 a_677477_25371# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2346 w_692190_39881# a_693130_40003# a_693330_37869# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2347 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2348 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2349 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2350 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2351 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2352 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2353 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2354 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2355 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2356 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2357 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2358 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2359 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2360 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2361 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2362 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2363 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2364 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2365 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2366 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2367 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2368 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2369 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2370 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2371 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2372 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2373 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2374 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2375 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2376 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2377 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2378 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2379 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2380 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2381 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2382 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2383 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2384 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2385 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2386 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2387 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2388 a_693549_59407# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2389 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2390 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2391 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2392 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2393 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2394 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2395 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2396 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2397 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2398 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2399 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2400 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2401 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2402 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2403 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2404 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2405 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2406 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2407 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2408 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2409 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2410 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2411 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2412 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2413 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2414 w_649931_37947# a_692386_37781# a_693330_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2415 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2416 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2417 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2418 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2419 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2420 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2421 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2422 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2423 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2424 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2425 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2426 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2427 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2428 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2429 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2430 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2431 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2432 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2433 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2434 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2435 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2436 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2437 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2438 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2439 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2440 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2441 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2442 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2443 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2444 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2445 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2446 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2447 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2448 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2449 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2450 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2451 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2452 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2453 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2454 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2455 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2456 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2457 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2458 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2459 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2460 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2461 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2462 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2463 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2464 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2465 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2466 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2467 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2468 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2469 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2470 a_722600_2050# a_719858_6024# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2471 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2472 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2473 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2474 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2475 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2476 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2477 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2478 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2479 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2480 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2481 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2482 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2483 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2484 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2485 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2486 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2487 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2488 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2489 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2490 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2491 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2492 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2493 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2494 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2495 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X2496 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2497 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2498 a_677477_25371# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2499 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2500 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2501 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2502 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2503 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2504 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2505 w_649931_37947# a_677477_25371# a_678421_20774# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2506 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2507 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2508 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2509 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2510 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2511 w_677281_20555# a_664155_35747# a_678421_20774# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2512 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2513 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2514 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2515 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2516 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2517 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2518 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2519 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2520 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2521 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2522 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2523 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2524 a_719742_79090# a_722600_82134# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2525 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2526 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2527 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2528 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2529 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2530 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2531 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2532 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2533 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2534 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2535 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2536 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2537 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2538 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2539 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2540 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2541 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2542 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2543 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2544 a_692386_37781# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2545 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2546 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2547 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2548 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2549 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2550 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2551 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2552 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2553 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2554 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2555 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2556 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2557 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2558 w_649931_37947# a_677477_25371# a_678421_20774# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2559 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2560 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2561 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2562 a_725512_8976# a_719900_5846# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2563 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2564 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2565 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2566 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2567 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2568 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2569 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2570 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2571 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2572 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2573 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2574 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2575 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2576 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2577 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2578 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2579 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2580 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2581 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2582 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2583 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2584 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2585 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2586 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2587 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2588 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2589 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2590 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2591 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2592 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2593 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2594 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2595 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2596 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2597 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2598 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2599 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2600 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2601 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2602 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2603 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2604 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2605 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2606 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2607 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2608 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2609 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2610 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2611 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2612 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2613 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2614 w_649931_37947# a_693549_25370# a_694493_20773# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2615 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2616 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2617 a_694493_20773# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2618 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2619 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2620 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2621 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2622 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2623 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2624 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2625 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2626 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2627 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2628 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2629 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2630 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2631 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2632 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2633 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2634 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2635 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2636 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2637 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2638 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2639 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2640 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2641 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2642 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2643 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2644 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2645 w_677281_61507# a_673159_61357# a_677477_59407# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2646 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2647 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2648 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2649 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2650 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2651 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2652 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2653 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2654 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2655 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2656 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2657 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2658 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2659 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2660 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2661 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2662 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2663 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2664 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2665 a_678421_20774# a_664155_35747# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2666 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2667 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2668 a_694493_20773# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2669 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2670 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2671 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2672 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2673 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2674 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2675 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2676 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2677 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2678 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2679 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2680 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2681 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2682 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2683 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2684 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2685 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2686 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2687 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2688 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2689 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2690 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2691 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2692 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2693 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2694 a_675258_41997# a_676490_42315# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X2695 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2696 a_664355_46657# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2697 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2698 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2699 a_725512_73584# a_719900_80508# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2700 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2701 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2702 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2703 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2704 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2705 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2706 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2707 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2708 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2709 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2710 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2711 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2712 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2713 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2714 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2715 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2716 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2717 a_650141_39687# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2718 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2719 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2720 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2721 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2722 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2723 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2724 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2725 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2726 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2727 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2728 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2729 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2730 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2731 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2732 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2733 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2734 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2735 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2736 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2737 w_649931_37947# a_719900_80508# a_725512_73584# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2738 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2739 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2740 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2741 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2742 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2743 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2744 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2745 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2746 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2747 a_673159_26571# a_666587_33613# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X2748 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2749 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2750 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2751 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2752 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2753 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X2754 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2755 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2756 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2757 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2758 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2759 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2760 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2761 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2762 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2763 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2764 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2765 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2766 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2767 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2768 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2769 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2770 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2771 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2772 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2773 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2774 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2775 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2776 w_678666_39881# a_676490_44223# a_678862_37781# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2777 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2778 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2779 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2780 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2781 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2782 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2783 w_663215_35625# a_662413_39580# a_663411_33525# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2784 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2785 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2786 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2787 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2788 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2789 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2790 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2791 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2792 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2793 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2794 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2795 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2796 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2797 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2798 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2799 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2800 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2801 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2802 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2803 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2804 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2805 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2806 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2807 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2808 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2809 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2810 w_649931_37947# a_677477_59407# a_677477_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2811 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2812 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2813 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2814 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2815 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2816 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2817 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2818 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2819 a_677477_59407# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2820 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2821 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2822 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2823 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2824 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2825 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2826 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2827 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2828 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2829 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2830 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2831 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2832 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2833 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2834 w_649931_37947# a_693549_25370# a_693549_25370# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2835 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2836 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2837 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2838 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2839 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2840 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2841 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2842 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2843 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2844 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2845 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2846 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2847 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2848 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2849 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2850 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2851 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2852 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2853 w_649931_37947# a_650053_38143# a_650141_47695# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2854 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2855 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2856 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2857 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2858 a_664355_33613# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2859 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2860 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2861 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2862 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2863 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2864 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2865 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2866 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2867 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2868 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2869 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2870 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2871 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2872 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2873 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2874 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2875 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2876 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2877 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2878 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2879 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2880 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2881 w_649931_37947# a_693549_25370# a_693549_25370# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2882 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2883 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2884 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2885 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2886 w_649931_37947# a_678862_37781# a_679806_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2887 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2888 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2889 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2890 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2891 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2892 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2893 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2894 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2895 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2896 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2897 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2898 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2899 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2900 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2901 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2902 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2903 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2904 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2905 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X2906 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2907 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2908 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2909 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2910 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2911 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2912 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2913 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2914 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2915 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2916 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2917 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2918 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2919 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2920 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2921 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2922 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2923 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2924 a_678862_37781# a_676490_44223# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2925 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2926 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2927 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2928 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2929 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2930 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2931 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2932 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2933 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2934 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2935 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2936 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2937 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2938 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2939 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2940 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2941 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2942 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2943 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2944 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2945 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2946 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2947 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2948 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2949 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2950 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2951 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2952 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2953 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2954 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2955 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2956 w_677281_20555# a_664155_35747# a_678421_20774# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2957 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2958 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2959 a_693549_25370# a_682038_37869# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2960 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2961 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2962 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2963 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2964 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2965 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2966 a_663411_33525# a_662413_39580# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2967 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2968 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2969 a_663411_51254# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2970 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2971 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2972 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2973 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2974 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2975 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2976 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2977 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2978 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2979 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2980 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2981 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2982 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2983 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2984 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X2985 w_663215_35625# a_664155_35747# a_664355_33613# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2986 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2987 w_678666_39881# a_664155_35747# a_679806_37869# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2988 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2989 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2990 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2991 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2992 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2993 a_677477_59407# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2994 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2995 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2996 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2997 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2998 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2999 w_649931_37947# a_677477_59407# a_678421_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3000 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3001 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3002 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3003 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3004 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3005 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3006 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3007 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3008 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3009 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3010 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3011 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3012 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3013 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3014 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3015 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3016 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3017 a_719858_6024# a_719332_5566# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3018 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3019 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3020 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3021 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3022 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3023 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3024 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3025 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3026 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3027 a_694493_59495# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3028 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3029 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3030 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3031 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3032 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3033 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3034 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3035 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3036 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3037 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3038 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3039 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3040 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3041 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3042 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3043 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3044 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3045 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3046 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3047 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3048 w_649931_37947# a_663411_33525# a_663411_33525# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3049 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3050 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3051 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3052 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3053 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3054 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3055 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3056 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3057 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3058 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3059 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3060 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3061 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3062 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3063 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3064 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3065 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3066 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3067 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3068 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3069 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3070 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3071 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3072 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3073 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3074 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3075 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3076 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3077 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3078 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3079 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3080 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3081 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3082 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3083 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3084 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3085 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3086 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3087 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3088 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3089 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3090 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3091 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3092 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3093 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3094 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3095 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3096 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3097 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3098 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3099 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3100 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3101 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3102 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3103 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3104 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3105 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3106 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3107 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3108 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3109 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3110 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3111 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3112 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3113 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3114 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3115 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3116 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3117 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3118 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3119 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3120 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3121 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3122 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3123 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3124 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3125 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3126 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3127 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3128 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3129 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3130 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3131 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3132 a_722600_75208# a_719858_79182# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3133 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3134 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3135 a_725512_n974# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3136 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3137 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3138 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3139 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3140 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3141 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3142 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3143 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3144 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3145 a_664355_33613# a_664155_35747# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3146 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3147 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3148 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3149 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X3150 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3151 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3152 w_649931_37947# a_677477_25371# a_678421_20774# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3153 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3154 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3155 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3156 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3157 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3158 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3159 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3160 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3161 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3162 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3163 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3164 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3165 a_673159_60085# a_674591_59767# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X3166 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3167 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3168 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3169 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3170 w_693353_20554# a_680653_25459# a_694493_20773# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3171 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3172 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3173 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3174 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3175 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3176 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3177 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3178 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3179 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3180 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3181 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3182 a_678421_59495# a_681073_63341# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=2.8e+06u
X3183 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3184 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3185 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3186 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3187 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3188 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3189 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3190 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3191 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3192 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3193 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3194 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3195 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3196 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3197 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3198 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3199 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3200 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3201 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3202 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3203 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3204 a_725512_82134# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3205 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3206 w_649931_37947# a_663411_51254# a_664355_46657# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3207 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3208 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3209 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3210 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3211 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3212 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3213 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3214 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3215 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3216 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3217 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3218 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3219 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3220 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3221 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3222 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3223 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3224 a_650141_46551# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3225 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3226 a_677477_25371# a_673159_24981# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3227 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3228 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3229 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3230 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3231 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3232 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3233 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3234 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3235 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3236 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3237 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3238 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3239 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3240 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3241 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3242 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3243 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3244 a_693549_59407# a_682038_37869# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3245 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3246 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3247 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3248 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3249 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3250 w_649931_37947# a_650053_38143# a_650053_38143# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3251 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3252 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3253 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3254 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3255 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3256 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3257 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3258 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3259 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3260 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3261 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3262 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3263 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3264 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3265 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3266 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3267 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3268 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3269 a_673159_24981# a_674591_24981# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X3270 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3271 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3272 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3273 a_663411_51254# a_663411_46560# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3274 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3275 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3276 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3277 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3278 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3279 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3280 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3281 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3282 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3283 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3284 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3285 a_667251_37508# a_666587_33613# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X3286 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3287 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3288 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3289 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3290 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3291 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3292 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3293 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3294 w_649931_37947# a_650053_38143# a_650141_38543# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3295 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3296 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3297 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3298 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3299 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3300 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3301 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3302 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3303 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3304 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3305 w_649931_37947# a_677477_59407# a_677477_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3306 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3307 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3308 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3309 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3310 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3311 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3312 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3313 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3314 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3315 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3316 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3317 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3318 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3319 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3320 w_649931_37947# a_650053_38143# a_650141_41975# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3321 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3322 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3323 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3324 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3325 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3326 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3327 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3328 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3329 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3330 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3331 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3332 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3333 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3334 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3335 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3336 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3337 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3338 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3339 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3340 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3341 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3342 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3343 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3344 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3345 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3346 w_649931_37947# a_663411_33525# a_663411_33525# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3347 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3348 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3349 w_663215_35625# a_662413_39580# a_663411_33525# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3350 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3351 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3352 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3353 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3354 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3355 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3356 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3357 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3358 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3359 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3360 a_662095_38148# a_662095_39580# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X3361 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3362 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3363 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3364 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3365 a_679806_37869# a_664155_35747# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3366 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3367 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3368 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3369 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3370 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3371 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3372 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3373 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3374 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3375 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3376 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3377 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3378 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3379 a_693549_25370# a_682038_37869# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3380 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3381 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3382 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3383 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3384 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3385 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3386 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3387 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3388 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3389 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3390 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3391 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3392 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3393 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3394 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3395 w_649931_37947# a_693549_59407# a_693549_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3396 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3397 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3398 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3399 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3400 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3401 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3402 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3403 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3404 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3405 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3406 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3407 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3408 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3409 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3410 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3411 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3412 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3413 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3414 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3415 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3416 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3417 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3418 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3419 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3420 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3421 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3422 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3423 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3424 a_679806_37869# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3425 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3426 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3427 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3428 w_677281_20555# a_664155_35747# a_678421_20774# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3429 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3430 w_649931_37947# a_678862_37781# a_678862_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3431 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3432 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3433 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3434 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3435 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3436 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3437 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3438 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3439 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3440 a_677477_59407# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3441 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3442 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3443 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3444 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3445 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3446 a_719742_7264# a_722600_2050# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3447 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3448 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3449 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3450 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3451 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3452 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3453 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3454 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3455 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3456 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3457 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3458 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3459 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3460 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3461 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3462 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3463 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3464 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3465 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3466 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3467 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3468 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3469 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3470 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3471 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3472 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3473 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3474 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3475 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3476 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3477 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3478 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3479 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3480 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3481 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3482 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3483 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3484 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3485 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3486 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3487 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3488 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3489 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3490 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3491 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3492 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3493 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3494 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3495 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3496 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3497 w_719104_5922# a_722600_82134# a_719742_79090# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3498 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3499 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3500 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3501 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3502 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3503 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3504 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3505 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3506 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3507 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3508 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3509 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3510 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3511 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3512 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3513 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3514 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3515 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3516 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3517 a_694493_20773# a_680653_25459# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3518 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3519 a_664355_33613# a_664155_35747# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3520 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3521 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3522 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3523 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3524 a_719900_5846# a_722600_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3525 a_663411_33525# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3526 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3527 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3528 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3529 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3530 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3531 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3532 a_650141_41975# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3533 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3534 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3535 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3536 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3537 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3538 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3539 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3540 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3541 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3542 w_663215_46438# a_663411_46560# a_663411_51254# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3543 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3544 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3545 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3546 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3547 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3548 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3549 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3550 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3551 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3552 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3553 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3554 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3555 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3556 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3557 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3558 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3559 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3560 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3561 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3562 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3563 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3564 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3565 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3566 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3567 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3568 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3569 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3570 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3571 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3572 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3573 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3574 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3575 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3576 a_719900_80508# a_722600_75208# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3577 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3578 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3579 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3580 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3581 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3582 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3583 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3584 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3585 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3586 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3587 a_725512_82134# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3588 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3589 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3590 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3591 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3592 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3593 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3594 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3595 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3596 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3597 a_678421_59495# a_664155_35747# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3598 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3599 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3600 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3601 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3602 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3603 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3604 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3605 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3606 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3607 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3608 w_678666_39881# a_664155_35747# a_679806_37869# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3609 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3610 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3611 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3612 w_677281_61507# a_673159_61357# a_677477_59407# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3613 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3614 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3615 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3616 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3617 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3618 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3619 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3620 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3621 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3622 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3623 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3624 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3625 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3626 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3627 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3628 w_649931_37947# a_677477_59407# a_678421_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3629 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3630 a_694493_59495# a_680653_59495# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3631 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3632 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3633 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3634 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3635 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3636 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3637 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3638 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3639 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3640 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3641 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3642 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3643 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3644 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3645 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3646 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3647 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3648 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3649 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3650 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3651 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3652 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3653 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3654 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3655 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3656 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3657 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3658 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3659 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3660 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3661 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3662 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3663 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3664 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3665 w_649931_37947# a_650053_38143# a_650141_40831# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3666 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3667 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3668 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3669 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3670 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3671 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3672 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3673 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3674 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3675 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3676 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3677 a_693330_37869# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3678 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3679 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3680 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3681 w_649931_37947# a_719900_5846# a_725512_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3682 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3683 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3684 w_649931_37947# a_678862_37781# a_679806_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3685 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3686 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3687 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X3688 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3689 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3690 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3691 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3692 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3693 a_679806_37869# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3694 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3695 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3696 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3697 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3698 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3699 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3700 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3701 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3702 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3703 a_650141_39687# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3704 a_725512_n974# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3705 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3706 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3707 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3708 w_719104_5922# a_722600_8976# a_719900_5846# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3709 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3710 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3711 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3712 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3713 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3714 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3715 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3716 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3717 a_719742_7264# a_722600_2050# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3718 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3719 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3720 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3721 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3722 w_693353_20554# a_682038_37869# a_693549_25370# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3723 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3724 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3725 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3726 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3727 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3728 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3729 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3730 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3731 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3732 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3733 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3734 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3735 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3736 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3737 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3738 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3739 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3740 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3741 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3742 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3743 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3744 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3745 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3746 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3747 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3748 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3749 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3750 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3751 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3752 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3753 a_663411_51254# a_663411_46560# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3754 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3755 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3756 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3757 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3758 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3759 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3760 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3761 a_675258_43269# a_676490_42951# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X3762 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3763 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3764 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3765 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3766 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3767 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3768 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3769 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3770 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3771 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3772 a_677477_59407# a_673159_61357# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3773 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3774 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3775 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3776 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3777 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3778 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3779 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3780 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3781 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3782 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3783 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3784 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3785 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3786 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3787 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3788 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3789 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3790 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3791 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3792 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3793 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3794 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3795 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3796 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3797 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3798 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3799 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3800 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3801 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3802 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3803 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3804 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3805 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3806 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3807 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3808 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3809 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3810 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3811 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3812 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3813 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3814 w_649931_37947# a_719900_80508# a_725512_73584# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3815 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3816 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3817 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3818 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3819 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3820 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3821 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3822 w_649931_37947# a_722600_75208# a_719900_80508# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3823 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3824 a_677477_59407# a_673159_61357# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3825 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3826 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3827 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3828 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3829 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3830 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3831 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3832 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3833 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3834 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3835 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3836 a_663411_33525# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3837 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3838 w_649931_37947# a_650053_38143# a_650141_47695# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3839 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3840 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3841 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3842 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3843 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3844 w_693353_61507# a_682038_37869# a_693549_59407# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3845 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3846 w_677281_20555# a_673159_24981# a_677477_25371# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3847 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X3848 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3849 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3850 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3851 a_676269_n1233# a_675951_199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X3852 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3853 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3854 a_681073_22635# a_678421_20774# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=2.8e+06u
X3855 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3856 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3857 a_694493_59495# a_680653_59495# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3858 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3859 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3860 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3861 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3862 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3863 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3864 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3865 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3866 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3867 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3868 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3869 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3870 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3871 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3872 a_664355_46657# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3873 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3874 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3875 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3876 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3877 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3878 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3879 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3880 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3881 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3882 w_678666_39881# a_664155_35747# a_679806_37869# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3883 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3884 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3885 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3886 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3887 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3888 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3889 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3890 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3891 w_649931_37947# a_719742_7264# a_725512_n974# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3892 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3893 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3894 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3895 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3896 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3897 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3898 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3899 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3900 w_663215_46438# a_662095_39580# a_664355_46657# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3901 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3902 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3903 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3904 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3905 w_719104_5922# a_722600_2050# a_719742_7264# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3906 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3907 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3908 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3909 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3910 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3911 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3912 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3913 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3914 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3915 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3916 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3917 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3918 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3919 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3920 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3921 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3922 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3923 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3924 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3925 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3926 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3927 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3928 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3929 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3930 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3931 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3932 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3933 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3934 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3935 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3936 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3937 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3938 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3939 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3940 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3941 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3942 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3943 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3944 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3945 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3946 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3947 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3948 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3949 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3950 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3951 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3952 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3953 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3954 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3955 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3956 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3957 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3958 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3959 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3960 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3961 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3962 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3963 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3964 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3965 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3966 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3967 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3968 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3969 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3970 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3971 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3972 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3973 w_677281_61507# a_664155_35747# a_678421_59495# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3974 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3975 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3976 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3977 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X3978 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3979 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3980 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3981 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3982 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3983 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3984 a_694493_20773# a_680653_25459# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3985 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3986 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3987 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3988 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3989 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3990 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3991 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3992 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3993 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3994 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3995 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3996 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X3997 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3998 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3999 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4000 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4001 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4002 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4003 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4004 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4005 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4006 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4007 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4008 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4009 w_663215_46438# a_662095_39580# a_664355_46657# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4010 w_649931_37947# a_693549_59407# a_693549_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4011 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4012 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4013 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4014 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4015 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4016 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4017 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4018 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4019 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4020 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4021 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4022 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4023 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X4024 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4025 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4026 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4027 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4028 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4029 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4030 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4031 a_693330_37869# a_693130_40003# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4032 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4033 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4034 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4035 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4036 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4037 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4038 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4039 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4040 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4041 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4042 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4043 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4044 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4045 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4046 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4047 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4048 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4049 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4050 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4051 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4052 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4053 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4054 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4055 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4056 a_650141_38543# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4057 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4058 a_725512_n974# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4059 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4060 w_649931_37947# a_663411_51254# a_663411_51254# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4061 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4062 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4063 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4064 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4065 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4066 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4067 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4068 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4069 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4070 a_673159_25299# a_674591_25617# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X4071 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4072 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4073 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4074 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4075 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4076 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4077 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4078 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4079 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4080 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4081 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4082 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4083 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4084 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4085 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X4086 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4087 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4088 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4089 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4090 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4091 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4092 a_693330_37869# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4093 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4094 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4095 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4096 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4097 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4098 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4099 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4100 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4101 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4102 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4103 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4104 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4105 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4106 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4107 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4108 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4109 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4110 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4111 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4112 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4113 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4114 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4115 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4116 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4117 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4118 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4119 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4120 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4121 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4122 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4123 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4124 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4125 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4126 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4127 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4128 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4129 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4130 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4131 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4132 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4133 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4134 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4135 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4136 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4137 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4138 a_664355_46657# a_662095_39580# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4139 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4140 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4141 w_678666_39881# a_676490_44223# a_678862_37781# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4142 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4143 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4144 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4145 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4146 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4147 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4148 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4149 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4150 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4151 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4152 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4153 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4154 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4155 w_649931_37947# a_663411_33525# a_664355_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4156 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4157 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4158 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4159 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4160 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4161 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4162 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4163 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4164 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X4165 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4166 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4167 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4168 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4169 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4170 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4171 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4172 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4173 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4174 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4175 a_678421_20774# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4176 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4177 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4178 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4179 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4180 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4181 a_678421_20774# a_664155_35747# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4182 a_676490_44223# a_682038_37869# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X4183 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4184 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4185 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4186 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4187 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4188 w_649931_37947# a_650053_38143# a_650141_46551# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4189 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4190 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4191 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4192 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4193 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4194 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4195 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4196 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4197 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4198 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4199 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4200 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4201 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4202 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4203 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4204 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4205 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4206 a_725512_8976# a_719900_5846# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4207 w_649931_37947# a_692386_37781# a_693330_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4208 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4209 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4210 w_693353_20554# a_682038_37869# a_693549_25370# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4211 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4212 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4213 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4214 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4215 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4216 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4217 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4218 w_649931_37947# a_650053_38143# a_650053_38143# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4219 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4220 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4221 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4222 a_678421_20774# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4223 w_649931_37947# a_722600_75208# a_719900_80508# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4224 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4225 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4226 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4227 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4228 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4229 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4230 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4231 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4232 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4233 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4234 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4235 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4236 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4237 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4238 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4239 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4240 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4241 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4242 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4243 a_678421_59495# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4244 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4245 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4246 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4247 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4248 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4249 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4250 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4251 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4252 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4253 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4254 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4255 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4256 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4257 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4258 w_649931_37947# a_693549_59407# a_694493_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4259 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4260 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4261 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4262 a_694493_59495# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4263 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4264 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4265 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4266 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4267 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4268 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4269 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4270 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4271 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4272 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4273 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4274 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4275 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4276 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4277 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4278 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4279 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4280 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4281 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4282 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4283 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4284 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4285 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4286 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4287 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4288 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4289 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4290 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4291 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4292 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4293 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4294 a_676490_44223# a_682038_37869# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X4295 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4296 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4297 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4298 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4299 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4300 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4301 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4302 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4303 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4304 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4305 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4306 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4307 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4308 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4309 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4310 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4311 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4312 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4313 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4314 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4315 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4316 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4317 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4318 w_693353_61507# a_682038_37869# a_693549_59407# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4319 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4320 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4321 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4322 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4323 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4324 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4325 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4326 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4327 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4328 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4329 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4330 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4331 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4332 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4333 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4334 w_663215_46438# a_663411_46560# a_663411_51254# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4335 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4336 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4337 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4338 w_649931_37947# a_663411_51254# a_663411_51254# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4339 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4340 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4341 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4342 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4343 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4344 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4345 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4346 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4347 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4348 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4349 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4350 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4351 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4352 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4353 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4354 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4355 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4356 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4357 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4358 a_719858_79182# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4359 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4360 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4361 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4362 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4363 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4364 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4365 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4366 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4367 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4368 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4369 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4370 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4371 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4372 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4373 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4374 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4375 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4376 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4377 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4378 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4379 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4380 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4381 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4382 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4383 w_649931_37947# a_693549_25370# a_693549_25370# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4384 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4385 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4386 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4387 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4388 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4389 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4390 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4391 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4392 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4393 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4394 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4395 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4396 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4397 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4398 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4399 a_693330_37869# a_693130_40003# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4400 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4401 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4402 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4403 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4404 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4405 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4406 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4407 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4408 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4409 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4410 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4411 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4412 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4413 a_679806_37869# a_664155_35747# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4414 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4415 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4416 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4417 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4418 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4419 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4420 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4421 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4422 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4423 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4424 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4425 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4426 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4427 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4428 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4429 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4430 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4431 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4432 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4433 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4434 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4435 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4436 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4437 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4438 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4439 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4440 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4441 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4442 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4443 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4444 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4445 w_649931_37947# a_719742_7264# a_725512_n974# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4446 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4447 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4448 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4449 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4450 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4451 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4452 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4453 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4454 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4455 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4456 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4457 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4458 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4459 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4460 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4461 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4462 w_649931_37947# a_693549_59407# a_693549_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4463 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4464 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4465 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4466 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4467 a_693549_25370# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4468 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4469 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4470 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4471 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4472 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4473 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4474 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4475 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4476 w_649931_37947# a_692386_37781# a_692386_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4477 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4478 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4479 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4480 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4481 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4482 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4483 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4484 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4485 w_649931_37947# a_650053_38143# a_650141_44263# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4486 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4487 w_649931_37947# a_722600_82134# a_719742_79090# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4488 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4489 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4490 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4491 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4492 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4493 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4494 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4495 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4496 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4497 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4498 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4499 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4500 w_678666_39881# a_676490_44223# a_678862_37781# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4501 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4502 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4503 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4504 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4505 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4506 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4507 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4508 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4509 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4510 a_650141_41975# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4511 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4512 a_693549_25370# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4513 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4514 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4515 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4516 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4517 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4518 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4519 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4520 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4521 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4522 a_678862_37781# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4523 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4524 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4525 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4526 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4527 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4528 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4529 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4530 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4531 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4532 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4533 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4534 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4535 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4536 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4537 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4538 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4539 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4540 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4541 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4542 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4543 a_663411_51254# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4544 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4545 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4546 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4547 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4548 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4549 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4550 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4551 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4552 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4553 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4554 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4555 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4556 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4557 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4558 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4559 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4560 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4561 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4562 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4563 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4564 w_649931_37947# a_678862_37781# a_678862_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4565 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4566 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4567 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4568 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4569 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4570 a_678862_37781# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4571 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4572 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4573 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4574 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4575 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4576 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4577 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4578 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4579 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4580 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4581 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4582 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4583 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4584 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4585 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4586 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4587 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4588 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4589 a_650141_47695# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4590 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4591 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4592 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4593 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4594 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4595 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4596 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4597 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4598 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4599 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4600 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4601 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4602 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4603 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4604 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4605 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4606 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4607 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4608 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4609 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4610 w_649931_37947# a_663411_51254# a_664355_46657# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4611 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4612 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4613 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4614 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4615 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4616 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4617 a_663411_33525# a_662413_39580# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4618 a_678862_37781# a_676490_44223# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4619 w_649931_37947# a_650053_38143# a_650141_40831# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4620 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4621 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4622 a_677477_59407# a_673159_61357# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4623 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4624 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4625 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4626 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4627 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4628 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4629 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4630 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4631 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4632 a_678421_59495# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4633 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4634 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4635 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4636 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4637 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4638 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4639 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4640 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4641 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4642 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4643 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4644 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4645 w_649931_37947# a_693549_25370# a_694493_20773# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4646 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4647 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4648 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4649 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4650 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4651 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4652 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4653 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4654 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4655 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4656 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4657 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4658 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4659 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4660 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4661 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4662 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4663 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4664 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4665 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4666 w_649931_37947# a_719742_79090# a_725512_82134# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4667 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4668 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4669 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4670 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4671 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4672 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4673 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4674 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4675 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4676 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4677 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4678 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4679 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4680 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4681 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4682 w_649931_37947# a_693549_25370# a_694493_20773# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4683 a_664355_33613# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4684 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4685 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4686 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4687 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4688 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4689 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4690 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4691 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4692 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4693 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4694 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4695 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4696 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4697 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4698 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4699 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4700 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4701 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4702 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4703 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4704 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4705 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4706 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4707 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4708 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4709 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4710 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4711 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4712 w_719104_5922# a_696725_25458# a_719858_6830# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4713 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4714 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4715 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4716 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4717 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4718 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4719 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4720 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4721 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4722 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4723 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4724 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4725 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4726 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4727 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4728 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4729 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4730 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4731 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4732 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4733 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4734 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4735 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4736 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4737 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4738 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4739 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4740 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4741 a_678421_20774# a_664155_35747# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4742 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4743 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4744 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4745 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4746 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4747 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4748 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4749 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4750 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4751 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4752 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4753 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4754 w_677281_20555# a_673159_24981# a_677477_25371# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4755 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4756 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4757 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4758 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4759 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4760 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4761 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4762 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4763 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4764 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4765 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4766 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4767 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4768 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4769 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4770 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4771 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4772 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4773 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4774 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4775 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4776 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4777 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4778 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4779 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4780 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4781 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4782 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4783 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4784 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4785 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4786 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4787 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4788 a_663411_51254# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4789 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4790 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4791 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4792 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4793 w_677281_61507# a_664155_35747# a_678421_59495# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4794 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4795 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4796 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4797 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4798 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4799 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4800 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4801 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4802 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4803 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4804 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4805 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4806 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4807 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4808 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4809 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4810 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4811 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4812 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4813 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X4814 a_677477_25371# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4815 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4816 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4817 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4818 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4819 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4820 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4821 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4822 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4823 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4824 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4825 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4826 a_674997_n1233# a_673159_24981# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X4827 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4828 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4829 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4830 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4831 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4832 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4833 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4834 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4835 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4836 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4837 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4838 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4839 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4840 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4841 w_649931_37947# a_693549_59407# a_694493_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4842 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4843 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4844 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4845 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4846 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4847 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4848 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4849 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4850 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4851 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4852 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4853 a_692386_37781# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4854 w_649931_37947# a_722600_82134# a_719742_79090# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4855 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4856 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4857 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4858 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4859 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4860 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4861 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4862 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4863 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4864 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4865 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4866 w_649931_37947# a_663411_33525# a_663411_33525# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4867 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4868 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4869 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4870 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4871 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4872 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4873 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4874 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4875 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4876 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4877 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4878 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4879 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4880 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4881 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4882 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4883 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4884 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4885 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4886 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4887 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4888 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4889 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4890 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4891 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4892 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4893 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4894 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4895 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4896 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4897 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4898 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4899 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4900 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4901 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4902 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4903 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4904 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4905 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4906 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4907 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4908 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4909 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4910 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4911 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4912 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4913 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4914 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4915 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4916 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4917 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4918 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4919 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4920 a_664355_33613# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4921 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4922 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4923 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4924 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4925 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4926 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4927 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4928 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4929 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4930 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4931 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4932 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4933 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4934 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4935 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4936 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4937 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4938 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4939 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4940 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4941 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4942 w_649931_37947# a_677477_25371# a_677477_25371# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4943 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4944 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4945 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4946 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4947 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4948 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4949 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4950 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4951 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4952 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4953 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4954 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4955 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4956 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4957 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4958 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4959 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4960 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X4961 a_677477_25371# a_673159_24981# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4962 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4963 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X4964 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4965 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4966 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4967 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4968 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4969 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4970 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X4971 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4972 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4973 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4974 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4975 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4976 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4977 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4978 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4979 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4980 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4981 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4982 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4983 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4984 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4985 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4986 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4987 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4988 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4989 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4990 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4991 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4992 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4993 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4994 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4995 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4996 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4997 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4998 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4999 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5000 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5001 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5002 a_650141_38543# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5003 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5004 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5005 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X5006 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5007 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5008 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5009 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5010 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5011 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5012 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5013 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5014 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5015 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5016 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5017 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5018 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5019 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5020 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5021 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5022 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5023 w_649931_37947# a_677477_25371# a_678421_20774# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5024 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5025 a_678421_20774# a_664155_35747# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5026 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5027 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5028 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5029 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5030 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5031 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5032 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5033 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5034 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X5035 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5036 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5037 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5038 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5039 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5040 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5041 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5042 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5043 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5044 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5045 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5046 a_693549_25370# a_682038_37869# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5047 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5048 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5049 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5050 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5051 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5052 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5053 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5054 a_722600_8976# a_719858_6830# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5055 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5056 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5057 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5058 w_649931_37947# a_692386_37781# a_693330_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5059 w_693353_20554# a_680653_25459# a_694493_20773# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5060 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5061 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5062 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5063 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5064 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5065 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5066 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5067 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5068 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5069 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5070 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5071 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5072 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5073 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5074 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5075 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5076 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5077 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5078 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5079 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5080 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X5081 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5082 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5083 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5084 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5085 a_676905_n1233# a_676587_199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X5086 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5087 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5088 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5089 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5090 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5091 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5092 w_719104_5922# a_722600_82134# a_719742_79090# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5093 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5094 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5095 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5096 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5097 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5098 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5099 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5100 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5101 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5102 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5103 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5104 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5105 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5106 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5107 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5108 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5109 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5110 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5111 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5112 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5113 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5114 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5115 w_649931_37947# a_719900_5846# a_725512_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5116 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5117 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5118 a_694493_20773# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5119 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5120 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5121 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5122 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5123 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5124 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5125 w_649931_37947# a_650053_38143# a_650141_46551# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5126 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5127 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5128 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5129 w_663215_35625# a_662413_39580# a_663411_33525# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5130 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5131 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5132 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5133 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5134 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5135 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5136 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5137 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5138 a_677477_25371# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5139 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5140 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5141 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5142 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5143 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5144 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5145 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5146 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5147 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5148 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5149 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5150 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5151 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5152 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5153 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5154 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5155 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5156 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5157 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5158 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5159 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5160 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5161 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5162 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5163 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5164 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5165 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5166 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5167 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5168 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5169 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5170 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5171 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5172 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5173 a_719900_80508# a_722600_75208# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5174 w_693353_61507# a_682038_37869# a_693549_59407# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5175 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5176 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5177 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5178 w_693353_61507# a_680653_59495# a_694493_59495# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5179 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5180 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5181 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5182 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5183 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5184 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5185 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5186 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5187 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5188 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5189 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5190 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5191 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5192 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5193 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5194 a_725512_82134# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5195 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5196 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5197 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5198 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5199 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5200 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5201 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5202 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5203 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5204 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5205 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5206 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5207 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5208 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5209 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5210 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5211 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5212 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5213 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5214 a_664355_33613# a_664155_35747# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5215 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5216 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5217 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5218 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5219 a_722600_8976# a_719858_6830# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5220 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5221 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5222 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5223 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5224 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5225 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5226 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5227 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5228 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5229 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5230 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5231 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5232 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5233 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5234 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5235 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5236 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5237 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5238 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5239 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5240 a_662095_38148# a_662413_39580# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X5241 a_678421_59495# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5242 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5243 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5244 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5245 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5246 a_722600_2050# a_719858_6024# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5247 w_649931_37947# a_693549_25370# a_694493_20773# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5248 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5249 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5250 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5251 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5252 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5253 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5254 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5255 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5256 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5257 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5258 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5259 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5260 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5261 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5262 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5263 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5264 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5265 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5266 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5267 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5268 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5269 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5270 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5271 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5272 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5273 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5274 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5275 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5276 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5277 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5278 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5279 a_678862_37781# a_676490_44223# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5280 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5281 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5282 w_649931_37947# a_719900_5846# a_725512_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5283 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5284 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5285 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5286 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5287 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5288 a_725512_73584# a_719900_80508# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5289 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5290 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5291 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X5292 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5293 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5294 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5295 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5296 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5297 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5298 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5299 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5300 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5301 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5302 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5303 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5304 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5305 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5306 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5307 w_649931_37947# a_677477_25371# a_677477_25371# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5308 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5309 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5310 a_677477_59407# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5311 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5312 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5313 w_677281_20555# a_673159_24981# a_677477_25371# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5314 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5315 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5316 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5317 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5318 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5319 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5320 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5321 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5322 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5323 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5324 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5325 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5326 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5327 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5328 a_693549_25370# a_682038_37869# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5329 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5330 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5331 w_649931_37947# a_693549_25370# a_693549_25370# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5332 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5333 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5334 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5335 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5336 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5337 a_663411_33525# a_662413_39580# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5338 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5339 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5340 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5341 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5342 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5343 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5344 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5345 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5346 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5347 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5348 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5349 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5350 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5351 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5352 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5353 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5354 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5355 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5356 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5357 w_649931_37947# a_677477_25371# a_677477_25371# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5358 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5359 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5360 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5361 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5362 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5363 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5364 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5365 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5366 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5367 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5368 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5369 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5370 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5371 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5372 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5373 w_649931_37947# a_692386_37781# a_692386_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5374 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5375 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5376 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5377 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5378 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5379 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5380 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5381 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5382 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5383 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5384 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5385 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5386 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5387 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5388 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5389 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5390 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5391 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5392 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5393 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5394 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5395 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5396 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5397 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5398 a_675258_43905# a_676490_44223# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X5399 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5400 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5401 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5402 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5403 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5404 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5405 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5406 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5407 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5408 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5409 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5410 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5411 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5412 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5413 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5414 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5415 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5416 w_649931_37947# a_719900_80508# a_725512_73584# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5417 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5418 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5419 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5420 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5421 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5422 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5423 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5424 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5425 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5426 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5427 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5428 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5429 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5430 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5431 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5432 w_649931_37947# a_719742_7264# a_725512_n974# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5433 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5434 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5435 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5436 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5437 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5438 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5439 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5440 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5441 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5442 a_693549_59407# a_682038_37869# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5443 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5444 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5445 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5446 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5447 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5448 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5449 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5450 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5451 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5452 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5453 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5454 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5455 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5456 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5457 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5458 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5459 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5460 a_650141_41975# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5461 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5462 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5463 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5464 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5465 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5466 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5467 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5468 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5469 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5470 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5471 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5472 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5473 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5474 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5475 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5476 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5477 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5478 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5479 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5480 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5481 w_663215_35625# a_664155_35747# a_664355_33613# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5482 w_692190_39881# a_664155_35747# a_692386_37781# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5483 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5484 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5485 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5486 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5487 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5488 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5489 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5490 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5491 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5492 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5493 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5494 a_678862_37781# a_676490_44223# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5495 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5496 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5497 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5498 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5499 a_664355_33613# a_664155_35747# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5500 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5501 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5502 w_649931_37947# a_678862_37781# a_679806_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5503 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5504 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5505 w_719104_5922# a_722600_82134# a_719742_79090# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5506 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5507 w_649931_37947# a_677477_59407# a_678421_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5508 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5509 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5510 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5511 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5512 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5513 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5514 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5515 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5516 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5517 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5518 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5519 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5520 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5521 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5522 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5523 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5524 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5525 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5526 w_693353_20554# a_680653_25459# a_694493_20773# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5527 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5528 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5529 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5530 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5531 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5532 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5533 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5534 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5535 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5536 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5537 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5538 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5539 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5540 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5541 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5542 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5543 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5544 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5545 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5546 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5547 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5548 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5549 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5550 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5551 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5552 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5553 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5554 a_650141_47695# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5555 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5556 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5557 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5558 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5559 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5560 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5561 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5562 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5563 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5564 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5565 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5566 a_692386_37781# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5567 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5568 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5569 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5570 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5571 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5572 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5573 a_676490_44223# a_682038_37869# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X5574 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5575 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5576 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5577 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5578 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5579 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5580 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5581 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5582 a_678421_59495# a_664155_35747# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5583 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5584 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5585 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5586 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5587 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5588 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5589 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5590 w_649931_37947# a_650053_38143# a_650141_40831# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5591 a_719900_80508# a_722600_75208# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5592 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5593 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5594 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5595 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5596 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5597 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5598 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5599 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5600 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5601 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5602 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5603 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5604 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5605 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5606 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5607 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5608 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5609 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5610 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5611 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5612 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5613 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5614 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5615 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5616 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5617 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5618 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5619 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5620 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5621 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5622 a_663411_51254# a_663411_46560# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5623 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5624 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5625 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5626 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5627 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5628 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5629 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5630 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5631 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5632 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5633 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5634 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5635 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5636 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5637 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X5638 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5639 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5640 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5641 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5642 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5643 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5644 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5645 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5646 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5647 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5648 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5649 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5650 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5651 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5652 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5653 w_693353_61507# a_680653_59495# a_694493_59495# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5654 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5655 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5656 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5657 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5658 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5659 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5660 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5661 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5662 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5663 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5664 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5665 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X5666 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5667 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5668 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5669 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5670 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5671 a_725512_8976# a_719900_5846# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5672 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5673 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5674 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5675 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5676 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5677 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5678 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5679 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5680 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5681 a_694493_20773# a_680653_25459# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5682 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5683 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5684 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5685 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5686 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5687 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5688 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5689 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5690 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5691 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5692 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5693 a_692386_37781# a_664155_35747# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5694 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5695 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5696 a_719900_5846# a_722600_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5697 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5698 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5699 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5700 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5701 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5702 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5703 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5704 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5705 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5706 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5707 w_649931_37947# a_719900_5846# a_725512_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5708 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5709 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5710 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5711 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5712 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5713 w_663215_35625# a_662413_39580# a_663411_33525# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5714 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5715 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5716 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5717 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5718 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5719 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5720 a_664355_46657# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5721 w_663215_46438# a_662095_39580# a_664355_46657# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5722 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5723 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5724 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5725 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5726 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5727 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5728 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5729 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5730 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5731 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5732 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5733 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5734 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5735 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5736 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5737 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5738 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5739 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5740 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5741 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5742 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5743 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5744 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5745 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5746 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5747 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5748 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5749 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X5750 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5751 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5752 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5753 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5754 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5755 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5756 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5757 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5758 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5759 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5760 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5761 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5762 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5763 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5764 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5765 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5766 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5767 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5768 a_650053_38143# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5769 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5770 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5771 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5772 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5773 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5774 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5775 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5776 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5777 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5778 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5779 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5780 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5781 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5782 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5783 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5784 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5785 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5786 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5787 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5788 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5789 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5790 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5791 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5792 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5793 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5794 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5795 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5796 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X5797 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5798 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5799 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5800 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5801 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5802 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5803 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5804 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5805 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5806 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5807 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5808 w_649931_37947# a_677477_59407# a_677477_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5809 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5810 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5811 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5812 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5813 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5814 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5815 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5816 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5817 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5818 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5819 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5820 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5821 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5822 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5823 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5824 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5825 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5826 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5827 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5828 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5829 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5830 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5831 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5832 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5833 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5834 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5835 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5836 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5837 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5838 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5839 a_676269_n1233# a_676587_199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X5840 w_649931_37947# a_719900_80508# a_725512_73584# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5841 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5842 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5843 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5844 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5845 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5846 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5847 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5848 a_650141_40831# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5849 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5850 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5851 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5852 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5853 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5854 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5855 w_719104_5922# a_722600_8976# a_719900_5846# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5856 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5857 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5858 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5859 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5860 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5861 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5862 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5863 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5864 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5865 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5866 w_678666_39881# a_676490_44223# a_678862_37781# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5867 w_649931_37947# a_650053_38143# a_650141_45407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5868 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5869 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5870 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5871 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5872 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5873 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5874 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5875 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5876 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5877 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5878 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5879 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5880 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5881 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5882 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5883 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5884 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5885 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5886 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5887 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5888 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5889 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5890 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5891 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5892 w_649931_37947# a_693549_59407# a_693549_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5893 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5894 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5895 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5896 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5897 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5898 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5899 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5900 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5901 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5902 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5903 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5904 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X5905 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5906 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5907 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5908 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5909 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5910 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5911 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5912 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5913 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5914 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5915 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5916 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5917 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5918 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5919 w_649931_37947# a_663411_51254# a_663411_51254# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5920 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5921 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5922 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5923 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5924 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5925 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5926 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5927 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5928 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5929 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5930 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5931 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5932 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5933 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5934 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5935 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5936 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5937 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5938 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5939 w_649931_37947# a_678862_37781# a_678862_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5940 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5941 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5942 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5943 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5944 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5945 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5946 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X5947 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5948 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5949 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5950 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5951 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5952 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5953 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5954 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5955 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5956 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5957 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5958 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5959 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5960 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5961 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5962 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5963 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5964 a_664355_46657# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5965 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5966 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5967 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5968 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5969 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5970 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5971 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5972 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5973 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5974 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5975 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5976 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5977 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5978 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X5979 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5980 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5981 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5982 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5983 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5984 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5985 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5986 w_649931_37947# a_663411_33525# a_664355_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5987 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5988 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5989 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5990 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5991 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5992 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5993 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5994 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5995 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5996 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5997 a_650141_45407# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5998 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5999 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6000 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6001 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6002 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6003 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6004 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6005 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6006 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6007 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6008 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6009 a_650141_38543# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6010 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6011 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6012 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6013 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6014 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6015 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6016 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6017 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6018 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6019 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6020 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6021 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6022 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6023 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6024 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6025 w_649931_37947# a_719742_7264# a_725512_n974# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6026 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6027 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6028 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6029 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6030 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6031 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6032 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6033 a_719900_5846# a_722600_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6034 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6035 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6036 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6037 w_719104_5922# a_722600_2050# a_719742_7264# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6038 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6039 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6040 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6041 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6042 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6043 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6044 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6045 a_676587_85767# a_676269_87199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X6046 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6047 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6048 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6049 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6050 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6051 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6052 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6053 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6054 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6055 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6056 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6057 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6058 w_649931_37947# a_663411_33525# a_664355_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6059 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6060 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6061 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6062 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6063 a_679806_37869# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6064 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6065 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6066 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6067 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6068 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6069 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6070 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6071 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6072 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6073 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6074 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6075 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6076 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6077 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6078 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6079 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6080 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6081 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6082 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6083 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6084 a_676490_44223# a_682038_37869# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X6085 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6086 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6087 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6088 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6089 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6090 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6091 w_693353_61507# a_680653_59495# a_694493_59495# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6092 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6093 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6094 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6095 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6096 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6097 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6098 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6099 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6100 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6101 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6102 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6103 a_693549_59407# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6104 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6105 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6106 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6107 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6108 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6109 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6110 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6111 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6112 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6113 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6114 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6115 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6116 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6117 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6118 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6119 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6120 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6121 a_682459_41330# a_682038_37869# sky130_fd_pr__cap_mim_m3_1 l=1.8e+07u w=2.7e+07u
X6122 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6123 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6124 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6125 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6126 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6127 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6128 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6129 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6130 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6131 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6132 a_693330_37869# a_693130_40003# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6133 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6134 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6135 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6136 w_677281_61507# a_664155_35747# a_678421_59495# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6137 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6138 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6139 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6140 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6141 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6142 w_649931_37947# a_650053_38143# a_650141_46551# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6143 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6144 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6145 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6146 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6147 a_679806_37869# a_664155_35747# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6148 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6149 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6150 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6151 a_677477_59407# a_673159_61357# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6152 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6153 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6154 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6155 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6156 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6157 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6158 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6159 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6160 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6161 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6162 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6163 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6164 w_649931_37947# a_650053_38143# a_650141_39687# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6165 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6166 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6167 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6168 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6169 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6170 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6171 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6172 w_649931_37947# a_719742_79090# a_725512_82134# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6173 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6174 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6175 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6176 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6177 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X6178 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6179 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6180 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6181 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6182 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6183 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6184 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6185 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6186 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6187 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6188 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6189 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6190 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6191 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6192 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6193 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6194 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6195 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6196 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6197 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6198 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6199 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6200 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6201 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6202 w_719104_5922# a_719900_5846# a_719858_6024# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6203 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6204 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6205 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6206 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6207 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6208 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6209 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6210 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6211 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6212 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6213 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6214 a_693330_37869# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6215 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6216 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6217 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6218 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6219 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6220 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6221 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6222 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6223 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6224 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6225 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6226 a_725512_n974# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6227 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6228 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6229 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6230 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6231 a_679806_37869# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6232 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6233 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6234 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6235 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6236 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6237 w_677281_20555# a_673159_24981# a_677477_25371# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6238 a_719742_7264# a_722600_2050# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6239 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6240 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6241 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6242 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6243 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6244 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6245 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6246 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6247 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6248 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6249 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6250 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6251 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6252 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6253 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6254 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6255 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6256 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6257 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6258 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6259 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6260 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6261 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6262 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6263 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6264 a_664355_46657# a_662095_39580# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6265 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6266 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6267 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6268 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6269 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6270 w_678666_39881# a_664155_35747# a_679806_37869# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6271 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6272 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6273 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6274 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6275 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6276 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6277 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6278 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6279 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6280 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6281 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6282 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6283 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6284 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6285 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6286 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6287 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6288 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6289 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6290 w_663215_46438# a_662095_39580# a_664355_46657# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6291 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6292 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6293 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6294 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6295 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6296 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6297 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6298 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6299 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6300 a_668545_37217# a_666587_33613# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=1.4e+07u
X6301 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6302 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6303 a_678421_20774# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6304 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6305 a_678421_20774# a_664155_35747# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6306 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6307 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6308 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6309 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6310 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6311 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6312 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6313 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6314 w_649931_37947# a_693549_59407# a_694493_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6315 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6316 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6317 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6318 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6319 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6320 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6321 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6322 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6323 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6324 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6325 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6326 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6327 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6328 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6329 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6330 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6331 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6332 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6333 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6334 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6335 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6336 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6337 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6338 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6339 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6340 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6341 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6342 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6343 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6344 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6345 w_649931_37947# a_719742_79090# a_725512_82134# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6346 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6347 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6348 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6349 a_678421_20774# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6350 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6351 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6352 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6353 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6354 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6355 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6356 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6357 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6358 w_649931_37947# a_678862_37781# a_679806_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6359 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6360 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6361 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6362 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6363 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6364 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6365 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6366 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6367 w_677281_61507# a_664155_35747# a_678421_59495# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6368 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6369 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6370 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6371 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6372 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6373 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X6374 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6375 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6376 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6377 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6378 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6379 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6380 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6381 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6382 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6383 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6384 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6385 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6386 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6387 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6388 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6389 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6390 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6391 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6392 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6393 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6394 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6395 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6396 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6397 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6398 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6399 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6400 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6401 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6402 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6403 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6404 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6405 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6406 w_692190_39881# a_664155_35747# a_692386_37781# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6407 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6408 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6409 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6410 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6411 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6412 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6413 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6414 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6415 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6416 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6417 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6418 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6419 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6420 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6421 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6422 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6423 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6424 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6425 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6426 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6427 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6428 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6429 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6430 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6431 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6432 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6433 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6434 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6435 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6436 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6437 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6438 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6439 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X6440 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6441 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6442 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6443 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6444 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6445 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6446 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6447 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6448 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6449 w_649931_37947# a_677477_59407# a_677477_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6450 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6451 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6452 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6453 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6454 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6455 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6456 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6457 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6458 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6459 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6460 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6461 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6462 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6463 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6464 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6465 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6466 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6467 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6468 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6469 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6470 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6471 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6472 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6473 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6474 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6475 w_649931_37947# a_663411_51254# a_664355_46657# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6476 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6477 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6478 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6479 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6480 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6481 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6482 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6483 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6484 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6485 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6486 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6487 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6488 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6489 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6490 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6491 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6492 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6493 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6494 a_678421_59495# a_664155_35747# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6495 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6496 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6497 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6498 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6499 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6500 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6501 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6502 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6503 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6504 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6505 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6506 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6507 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6508 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6509 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6510 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6511 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6512 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6513 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6514 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6515 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6516 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6517 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6518 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6519 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6520 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6521 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6522 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6523 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6524 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6525 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6526 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6527 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6528 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6529 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6530 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6531 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6532 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6533 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6534 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6535 a_664355_46657# a_662095_39580# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6536 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6537 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6538 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6539 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6540 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6541 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6542 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6543 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6544 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6545 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6546 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6547 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6548 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6549 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6550 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6551 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6552 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6553 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6554 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6555 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6556 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6557 a_650141_47695# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6558 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6559 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6560 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6561 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6562 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6563 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6564 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6565 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6566 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6567 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6568 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6569 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6570 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6571 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6572 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6573 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6574 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6575 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6576 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6577 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6578 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6579 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6580 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6581 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6582 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6583 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6584 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6585 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6586 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6587 a_693549_25370# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6588 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6589 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6590 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6591 a_692386_37781# a_664155_35747# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6592 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6593 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6594 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6595 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6596 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6597 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6598 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6599 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6600 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6601 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6602 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6603 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6604 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6605 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6606 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6607 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6608 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6609 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6610 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6611 w_649931_37947# a_663411_33525# a_663411_33525# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6612 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6613 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6614 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6615 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6616 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6617 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6618 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6619 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6620 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6621 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6622 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6623 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6624 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6625 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6626 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6627 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6628 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6629 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6630 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6631 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6632 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6633 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6634 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6635 a_693549_25370# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6636 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6637 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6638 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6639 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6640 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6641 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6642 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6643 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6644 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6645 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6646 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6647 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6648 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6649 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6650 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6651 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6652 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6653 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6654 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6655 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6656 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6657 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6658 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6659 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6660 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6661 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6662 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6663 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6664 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6665 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6666 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6667 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6668 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6669 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6670 a_673159_60721# a_674591_60403# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X6671 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6672 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6673 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6674 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6675 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6676 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6677 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6678 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6679 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6680 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6681 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6682 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6683 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6684 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6685 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6686 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6687 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6688 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6689 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6690 a_650141_44263# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6691 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6692 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6693 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6694 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6695 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6696 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6697 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6698 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6699 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6700 a_725512_82134# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6701 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6702 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6703 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6704 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6705 a_678421_20774# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6706 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6707 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6708 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6709 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6710 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6711 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6712 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6713 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6714 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6715 w_693353_61507# a_682038_37869# a_693549_59407# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6716 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6717 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6718 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6719 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6720 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6721 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6722 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6723 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6724 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6725 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6726 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6727 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6728 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6729 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6730 w_663215_46438# a_663411_46560# a_663411_51254# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6731 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6732 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6733 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6734 w_649931_37947# a_719742_79090# a_725512_82134# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6735 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6736 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6737 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6738 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6739 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6740 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6741 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6742 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6743 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6744 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6745 a_693330_37869# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6746 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6747 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6748 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6749 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6750 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6751 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6752 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6753 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6754 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6755 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6756 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6757 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6758 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6759 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6760 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6761 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6762 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6763 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6764 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6765 a_678421_59495# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6766 w_677281_61507# a_673159_61357# a_677477_59407# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6767 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6768 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6769 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6770 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6771 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6772 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6773 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6774 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6775 w_649931_37947# a_677477_59407# a_678421_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6776 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6777 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6778 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X6779 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6780 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6781 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6782 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6783 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6784 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6785 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6786 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6787 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6788 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6789 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6790 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6791 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6792 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6793 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6794 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6795 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6796 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6797 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6798 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6799 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6800 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6801 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6802 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6803 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6804 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6805 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6806 w_649931_37947# a_719900_5846# a_725512_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6807 w_649931_37947# a_693549_59407# a_694493_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6808 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6809 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6810 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6811 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6812 a_694493_59495# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6813 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6814 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6815 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6816 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6817 a_663411_33525# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6818 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6819 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6820 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6821 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6822 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6823 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6824 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6825 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6826 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6827 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6828 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6829 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6830 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6831 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6832 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6833 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6834 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6835 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6836 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6837 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6838 a_664355_33613# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6839 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6840 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6841 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6842 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6843 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6844 a_650141_40831# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6845 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6846 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6847 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6848 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6849 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6850 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6851 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6852 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6853 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6854 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6855 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6856 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6857 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6858 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6859 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6860 w_693353_20554# a_682038_37869# a_693549_25370# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6861 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6862 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6863 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6864 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6865 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6866 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6867 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6868 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6869 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6870 w_649931_37947# a_650053_38143# a_650141_45407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6871 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6872 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6873 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6874 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6875 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6876 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6877 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6878 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6879 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6880 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6881 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6882 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6883 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6884 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6885 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6886 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6887 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6888 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6889 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6890 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6891 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6892 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6893 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6894 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6895 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6896 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6897 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6898 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6899 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6900 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6901 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X6902 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6903 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6904 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6905 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6906 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6907 w_663215_35625# a_662413_39580# a_663411_33525# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6908 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6909 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6910 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6911 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6912 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6913 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6914 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6915 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6916 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6917 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6918 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6919 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6920 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6921 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6922 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6923 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6924 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6925 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6926 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6927 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6928 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6929 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6930 a_650141_46551# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6931 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6932 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6933 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6934 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6935 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6936 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6937 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6938 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6939 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6940 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6941 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6942 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6943 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X6944 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6945 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6946 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6947 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6948 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6949 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6950 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6951 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6952 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6953 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6954 a_725512_73584# a_719900_80508# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6955 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6956 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6957 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6958 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6959 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6960 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6961 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6962 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6963 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6964 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6965 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6966 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6967 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6968 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6969 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6970 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6971 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6972 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6973 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6974 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6975 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6976 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6977 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6978 a_650141_45407# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6979 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6980 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6981 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6982 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X6983 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6984 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6985 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X6986 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6987 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6988 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6989 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6990 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X6991 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6992 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6993 w_649931_37947# a_693549_59407# a_693549_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6994 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6995 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6996 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6997 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6998 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6999 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7000 a_693549_25370# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7001 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7002 w_719104_5922# a_719858_79182# a_722600_75208# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7003 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7004 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7005 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7006 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7007 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7008 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7009 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7010 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7011 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7012 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7013 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7014 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7015 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7016 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7017 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7018 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7019 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7020 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7021 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7022 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7023 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7024 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7025 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7026 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7027 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7028 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7029 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7030 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7031 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7032 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7033 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7034 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7035 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7036 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7037 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7038 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7039 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7040 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7041 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7042 a_678862_37781# a_676490_44223# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7043 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7044 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7045 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7046 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7047 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7048 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7049 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7050 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7051 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7052 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7053 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7054 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7055 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7056 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7057 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7058 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7059 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7060 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7061 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7062 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7063 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7064 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7065 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7066 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7067 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7068 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7069 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7070 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7071 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7072 w_649931_37947# a_663411_51254# a_664355_46657# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7073 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7074 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7075 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7076 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7077 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7078 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7079 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7080 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7081 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7082 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7083 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7084 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7085 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7086 a_663411_33525# a_662413_39580# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7087 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7088 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7089 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7090 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7091 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7092 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7093 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7094 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7095 a_678862_37781# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7096 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7097 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7098 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7099 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7100 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7101 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7102 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7103 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7104 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7105 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7106 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7107 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7108 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7109 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7110 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7111 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7112 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7113 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7114 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7115 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7116 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7117 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7118 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7119 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7120 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7121 a_675258_41997# a_676490_41997# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X7122 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7123 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7124 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7125 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7126 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7127 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7128 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7129 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7130 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7131 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7132 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7133 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7134 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7135 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7136 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7137 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7138 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7139 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7140 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7141 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7142 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7143 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7144 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7145 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7146 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7147 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7148 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7149 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7150 w_719104_5922# a_722600_82134# a_719742_79090# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7151 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7152 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7153 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7154 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7155 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7156 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7157 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7158 a_678421_20774# a_664155_35747# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7159 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7160 a_678862_37781# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7161 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7162 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7163 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7164 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7165 a_678421_59495# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7166 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7167 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7168 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7169 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7170 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7171 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7172 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7173 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7174 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7175 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7176 w_649931_37947# a_693549_25370# a_694493_20773# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7177 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7178 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X7179 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7180 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7181 a_694493_20773# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7182 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7183 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7184 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7185 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7186 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7187 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7188 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7189 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7190 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7191 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7192 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7193 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7194 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7195 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7196 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7197 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7198 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7199 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7200 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7201 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7202 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7203 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7204 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7205 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7206 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7207 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7208 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7209 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7210 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7211 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7212 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7213 w_649931_37947# a_678862_37781# a_678862_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7214 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7215 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7216 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7217 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7218 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7219 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7220 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7221 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7222 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7223 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7224 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7225 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7226 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7227 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7228 w_649931_37947# a_692386_37781# a_693330_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7229 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7230 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7231 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7232 a_694493_20773# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7233 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7234 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7235 a_719900_80508# a_722600_75208# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7236 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7237 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7238 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7239 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7240 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7241 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7242 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7243 a_675258_43905# a_676490_43587# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X7244 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7245 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7246 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7247 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7248 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7249 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7250 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7251 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7252 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7253 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7254 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7255 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7256 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7257 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7258 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7259 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7260 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7261 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7262 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7263 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7264 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7265 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7266 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7267 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7268 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7269 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7270 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7271 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7272 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7273 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7274 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7275 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7276 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7277 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7278 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7279 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7280 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7281 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7282 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7283 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7284 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7285 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7286 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7287 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7288 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7289 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7290 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7291 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7292 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7293 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7294 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7295 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7296 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7297 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7298 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7299 w_677281_20555# a_664155_35747# a_678421_20774# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7300 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7301 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7302 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7303 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7304 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7305 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7306 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7307 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7308 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7309 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7310 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7311 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7312 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7313 a_677477_25371# a_673159_24981# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7314 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7315 w_719104_5922# a_719900_80508# a_719858_79988# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7316 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7317 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7318 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7319 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7320 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7321 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7322 a_719900_5846# a_722600_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7323 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7324 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7325 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7326 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7327 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7328 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7329 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7330 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7331 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7332 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7333 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7334 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7335 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7336 w_663215_35625# a_664155_35747# a_664355_33613# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7337 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7338 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7339 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7340 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7341 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7342 w_692190_39881# a_693130_40003# a_693330_37869# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7343 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7344 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7345 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7346 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7347 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7348 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7349 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7350 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7351 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7352 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7353 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7354 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7355 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7356 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7357 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7358 a_663411_51254# a_663411_46560# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7359 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7360 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7361 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7362 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7363 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7364 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7365 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7366 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7367 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7368 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7369 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7370 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7371 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7372 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7373 a_678421_59495# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7374 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7375 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7376 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7377 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7378 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7379 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7380 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7381 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7382 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7383 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7384 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7385 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7386 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7387 a_668545_48760# a_663411_46560# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=1.4e+07u
X7388 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7389 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7390 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7391 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7392 a_668545_48760# a_664355_46657# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=500000u
X7393 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7394 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7395 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7396 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7397 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7398 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7399 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7400 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7401 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7402 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7403 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7404 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7405 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7406 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7407 a_694493_59495# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7408 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7409 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7410 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7411 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7412 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7413 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7414 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7415 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7416 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7417 a_719332_79990# a_696725_59495# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7418 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7419 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7420 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7421 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7422 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7423 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7424 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7425 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7426 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7427 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7428 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7429 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7430 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7431 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7432 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7433 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7434 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7435 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7436 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7437 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7438 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7439 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7440 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7441 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7442 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7443 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7444 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7445 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7446 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7447 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X7448 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7449 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7450 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7451 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7452 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7453 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7454 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7455 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7456 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7457 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7458 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7459 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7460 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7461 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7462 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7463 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7464 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7465 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7466 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7467 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7468 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7469 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7470 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7471 a_693549_25370# a_682038_37869# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7472 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7473 w_649931_37947# a_719900_80508# a_725512_73584# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7474 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7475 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7476 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7477 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7478 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7479 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7480 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7481 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7482 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7483 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7484 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7485 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7486 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7487 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7488 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7489 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7490 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7491 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7492 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7493 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7494 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7495 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7496 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7497 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7498 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7499 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7500 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7501 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7502 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7503 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7504 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7505 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7506 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7507 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7508 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7509 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7510 w_649931_37947# a_692386_37781# a_692386_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7511 a_677477_25371# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7512 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7513 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7514 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7515 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7516 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7517 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7518 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7519 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7520 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7521 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7522 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7523 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7524 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7525 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7526 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7527 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7528 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7529 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7530 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7531 w_677281_20555# a_664155_35747# a_678421_20774# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7532 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7533 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7534 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7535 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7536 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7537 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7538 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7539 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7540 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7541 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7542 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7543 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7544 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7545 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7546 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7547 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7548 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7549 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7550 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7551 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7552 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7553 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7554 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7555 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7556 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7557 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7558 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7559 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7560 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7561 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7562 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7563 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7564 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7565 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7566 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7567 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7568 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7569 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7570 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7571 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7572 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7573 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7574 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7575 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7576 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7577 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7578 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7579 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7580 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7581 a_693549_59407# a_682038_37869# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7582 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7583 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7584 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7585 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7586 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7587 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7588 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7589 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7590 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7591 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7592 w_693353_61507# a_680653_59495# a_694493_59495# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7593 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7594 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7595 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7596 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7597 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7598 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7599 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7600 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7601 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7602 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7603 w_649931_37947# a_719742_7264# a_725512_n974# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7604 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7605 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7606 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7607 w_649931_37947# a_693549_59407# a_693549_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7608 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7609 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7610 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7611 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7612 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7613 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7614 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7615 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7616 w_649931_37947# a_663411_51254# a_663411_51254# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7617 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7618 w_692190_39881# a_664155_35747# a_692386_37781# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7619 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7620 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7621 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7622 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7623 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7624 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7625 a_694493_20773# a_680653_25459# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7626 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7627 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7628 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7629 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7630 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7631 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7632 a_664355_33613# a_664155_35747# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7633 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7634 a_663411_33525# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7635 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7636 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7637 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7638 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7639 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7640 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7641 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7642 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7643 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7644 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7645 w_677281_61507# a_673159_61357# a_677477_59407# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7646 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7647 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7648 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7649 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7650 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7651 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7652 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7653 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7654 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7655 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7656 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7657 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7658 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7659 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7660 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7661 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7662 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7663 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7664 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7665 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7666 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7667 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7668 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7669 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7670 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7671 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7672 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7673 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7674 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7675 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7676 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7677 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7678 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7679 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7680 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7681 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7682 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7683 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7684 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7685 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7686 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7687 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7688 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7689 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7690 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7691 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7692 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7693 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7694 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7695 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7696 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7697 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7698 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7699 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7700 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7701 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7702 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7703 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7704 w_649931_37947# a_677477_25371# a_678421_20774# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7705 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7706 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7707 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7708 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7709 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7710 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7711 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7712 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7713 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7714 a_678421_59495# a_664155_35747# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7715 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7716 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7717 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7718 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7719 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7720 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7721 w_693353_20554# a_680653_25459# a_694493_20773# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7722 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7723 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7724 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7725 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7726 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7727 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7728 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7729 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7730 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7731 a_694493_59495# a_680653_59495# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7732 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7733 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7734 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7735 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7736 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7737 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7738 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7739 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7740 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7741 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7742 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7743 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7744 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7745 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7746 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7747 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7748 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7749 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7750 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7751 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7752 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7753 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7754 a_719858_79182# a_696725_59495# a_719858_78562# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7755 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7756 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7757 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7758 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7759 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7760 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7761 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7762 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7763 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7764 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7765 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7766 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7767 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7768 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7769 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7770 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7771 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7772 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7773 a_725512_n974# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7774 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7775 a_675951_85767# a_676269_87199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X7776 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7777 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7778 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7779 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7780 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7781 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7782 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7783 w_649931_37947# a_719742_79090# a_725512_82134# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7784 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7785 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7786 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7787 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X7788 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7789 a_650141_40831# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7790 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7791 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7792 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7793 a_694493_20773# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7794 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7795 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7796 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7797 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7798 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7799 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7800 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7801 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7802 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7803 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7804 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7805 a_663411_51254# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7806 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7807 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7808 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7809 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7810 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7811 w_693353_20554# a_682038_37869# a_693549_25370# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7812 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7813 a_674997_n1233# a_675315_199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X7814 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7815 w_649931_37947# a_650053_38143# a_650141_45407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7816 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7817 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7818 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7819 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7820 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7821 a_664355_46657# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7822 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7823 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7824 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7825 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7826 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7827 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7828 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7829 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7830 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7831 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7832 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7833 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7834 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7835 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7836 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7837 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7838 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7839 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7840 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7841 w_649931_37947# a_677477_25371# a_677477_25371# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7842 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7843 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7844 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7845 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7846 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7847 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7848 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7849 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7850 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7851 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7852 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7853 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7854 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X7855 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7856 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7857 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7858 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7859 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7860 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7861 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7862 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7863 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7864 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7865 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7866 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7867 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7868 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7869 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7870 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7871 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7872 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7873 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7874 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7875 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7876 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7877 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7878 w_663215_35625# a_664155_35747# a_664355_33613# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7879 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7880 a_650141_46551# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7881 a_664355_33613# a_668545_37217# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=500000u
X7882 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7883 w_649931_37947# a_663411_33525# a_664355_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7884 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7885 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7886 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7887 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7888 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7889 w_663215_46438# a_663411_46560# a_663411_51254# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7890 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7891 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7892 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7893 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7894 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X7895 a_678862_37781# a_676490_44223# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7896 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7897 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7898 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7899 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7900 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7901 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7902 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7903 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7904 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7905 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7906 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7907 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7908 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7909 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7910 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7911 a_692386_37781# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7912 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7913 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7914 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7915 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7916 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7917 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7918 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7919 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7920 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7921 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7922 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X7923 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7924 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7925 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7926 w_693353_61507# a_682038_37869# a_693549_59407# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7927 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7928 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7929 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7930 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7931 a_650141_45407# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7932 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7933 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7934 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7935 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7936 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7937 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7938 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7939 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7940 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7941 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7942 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7943 a_722600_75208# a_719858_79182# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7944 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7945 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7946 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7947 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7948 w_677281_61507# a_673159_61357# a_677477_59407# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7949 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7950 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7951 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7952 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7953 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7954 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7955 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7956 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7957 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7958 a_693130_40003# a_676490_41997# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=9e+06u
X7959 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7960 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7961 w_678666_39881# a_664155_35747# a_679806_37869# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7962 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7963 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7964 a_676587_85767# a_676905_87199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X7965 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7966 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7967 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7968 a_678421_59495# a_664155_35747# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7969 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7970 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7971 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7972 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7973 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7974 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7975 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7976 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7977 w_649931_37947# a_693549_25370# a_693549_25370# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7978 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7979 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7980 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7981 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7982 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7983 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7984 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7985 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7986 a_725512_73584# a_719900_80508# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7987 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7988 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7989 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7990 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7991 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7992 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7993 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X7994 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7995 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7996 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7997 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7998 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7999 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8000 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8001 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8002 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8003 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8004 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8005 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8006 a_675951_85767# a_675633_87199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X8007 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8008 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8009 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8010 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8011 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8012 a_692386_37781# a_664155_35747# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8013 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8014 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8015 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8016 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8017 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8018 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8019 w_649931_37947# a_692386_37781# a_692386_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8020 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8021 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8022 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8023 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8024 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8025 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8026 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8027 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8028 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8029 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8030 w_649931_37947# a_678862_37781# a_679806_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8031 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8032 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8033 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8034 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8035 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8036 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8037 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8038 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8039 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8040 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8041 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8042 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8043 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8044 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8045 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8046 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8047 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8048 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8049 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8050 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8051 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8052 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8053 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8054 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8055 a_694493_20773# a_680653_25459# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8056 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8057 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8058 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8059 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8060 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8061 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8062 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8063 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8064 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8065 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8066 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8067 a_663411_51254# a_663411_46560# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8068 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8069 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8070 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8071 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8072 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8073 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8074 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8075 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8076 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8077 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8078 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8079 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8080 w_663215_46438# a_662095_39580# a_664355_46657# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8081 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8082 a_663411_51254# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8083 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8084 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8085 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8086 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8087 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8088 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8089 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8090 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8091 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8092 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8093 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8094 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8095 w_649931_37947# a_692386_37781# a_693330_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8096 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8097 a_719858_79988# a_719900_80508# a_719858_80608# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8098 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8099 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8100 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8101 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8102 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8103 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8104 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8105 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8106 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8107 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8108 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8109 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8110 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8111 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8112 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8113 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8114 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8115 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8116 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8117 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8118 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8119 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8120 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8121 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8122 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8123 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8124 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8125 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8126 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8127 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8128 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8129 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8130 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8131 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8132 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8133 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8134 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8135 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8136 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8137 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8138 a_677477_59407# a_673159_61357# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8139 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8140 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8141 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8142 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8143 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8144 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8145 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8146 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8147 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8148 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8149 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8150 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8151 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8152 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8153 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8154 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8155 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8156 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8157 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8158 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8159 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8160 a_719900_5846# a_722600_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8161 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8162 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8163 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8164 w_719104_5922# a_722600_75208# a_719900_80508# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8165 w_649931_37947# a_650053_38143# a_650141_44263# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8166 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8167 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8168 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8169 a_694493_59495# a_680653_59495# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8170 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8171 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8172 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8173 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8174 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8175 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8176 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8177 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8178 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8179 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8180 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8181 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8182 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8183 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8184 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8185 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8186 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8187 a_693549_59407# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8188 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8189 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8190 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8191 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8192 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8193 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8194 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8195 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8196 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8197 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8198 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8199 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8200 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8201 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8202 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8203 w_692190_39881# a_693130_40003# a_693330_37869# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8204 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8205 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8206 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8207 w_692190_39881# a_693130_40003# a_693330_37869# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8208 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8209 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8210 a_692386_37781# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8211 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8212 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8213 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8214 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8215 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8216 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8217 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8218 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8219 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8220 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8221 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8222 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8223 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8224 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8225 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8226 a_664355_46657# a_662095_39580# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8227 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8228 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8229 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8230 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8231 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8232 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8233 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8234 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8235 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8236 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8237 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8238 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8239 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8240 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8241 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8242 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8243 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8244 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8245 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8246 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8247 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8248 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8249 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8250 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8251 a_725512_8976# a_719900_5846# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8252 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8253 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8254 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8255 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8256 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8257 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8258 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8259 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8260 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8261 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8262 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8263 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8264 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8265 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8266 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8267 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8268 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8269 a_719332_5566# a_696725_25458# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8270 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8271 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8272 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8273 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8274 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8275 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8276 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8277 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8278 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8279 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8280 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8281 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8282 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8283 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8284 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8285 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8286 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8287 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8288 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8289 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8290 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8291 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8292 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8293 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8294 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8295 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8296 w_649931_37947# a_677477_59407# a_677477_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8297 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8298 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8299 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8300 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8301 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8302 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8303 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8304 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8305 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8306 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8307 a_673159_26571# a_674591_26253# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X8308 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8309 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8310 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8311 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8312 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8313 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8314 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8315 a_725512_n974# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8316 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8317 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8318 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8319 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8320 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8321 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8322 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8323 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8324 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8325 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8326 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8327 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8328 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8329 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8330 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8331 a_719742_7264# a_722600_2050# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8332 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8333 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8334 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8335 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8336 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8337 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8338 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8339 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8340 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8341 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8342 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8343 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8344 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8345 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8346 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8347 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8348 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8349 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8350 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8351 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8352 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8353 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8354 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8355 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8356 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8357 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8358 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8359 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8360 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8361 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8362 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8363 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8364 w_649931_37947# a_719900_5846# a_725512_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8365 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8366 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8367 a_725512_73584# a_719900_80508# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8368 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8369 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8370 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8371 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8372 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8373 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8374 a_719900_80508# a_722600_75208# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8375 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8376 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8377 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8378 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8379 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8380 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8381 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8382 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8383 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8384 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8385 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8386 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8387 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8388 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8389 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8390 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8391 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8392 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8393 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8394 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8395 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8396 w_663215_46438# a_663411_46560# a_663411_51254# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8397 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8398 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8399 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8400 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8401 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8402 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8403 w_649931_37947# a_663411_33525# a_663411_33525# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8404 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8405 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8406 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8407 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8408 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8409 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8410 w_649931_37947# a_650053_38143# a_650141_38543# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8411 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8412 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8413 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8414 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8415 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8416 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8417 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8418 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8419 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8420 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8421 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8422 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8423 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8424 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8425 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8426 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8427 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8428 w_649931_37947# a_650053_38143# a_650141_41975# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8429 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8430 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8431 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8432 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8433 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8434 w_692190_39881# a_664155_35747# a_692386_37781# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8435 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8436 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8437 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8438 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8439 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8440 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8441 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8442 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8443 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8444 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8445 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8446 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8447 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8448 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8449 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8450 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8451 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8452 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8453 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8454 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8455 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8456 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8457 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8458 a_664355_33613# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8459 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8460 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8461 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8462 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8463 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8464 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8465 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8466 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8467 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8468 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8469 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8470 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8471 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8472 w_649931_37947# a_719742_7264# a_725512_n974# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8473 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8474 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8475 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8476 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8477 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8478 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8479 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8480 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8481 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8482 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8483 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8484 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8485 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8486 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8487 w_693353_20554# a_682038_37869# a_693549_25370# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8488 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8489 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8490 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8491 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8492 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8493 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8494 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8495 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8496 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8497 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8498 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8499 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8500 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8501 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8502 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8503 a_725512_73584# a_719900_80508# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8504 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8505 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8506 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8507 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8508 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8509 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8510 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8511 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8512 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8513 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8514 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8515 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8516 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8517 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8518 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8519 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8520 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8521 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8522 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8523 w_649931_37947# a_678862_37781# a_678862_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8524 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8525 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8526 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8527 a_678421_59495# a_664155_35747# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8528 a_676490_44223# a_682038_37869# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X8529 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8530 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8531 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8532 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8533 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8534 w_649931_37947# a_677477_59407# a_677477_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8535 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8536 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8537 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8538 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8539 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8540 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8541 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8542 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8543 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8544 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8545 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8546 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8547 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8548 a_694493_59495# a_680653_59495# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8549 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8550 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8551 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8552 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8553 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8554 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8555 a_693549_59407# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8556 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8557 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8558 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8559 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8560 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8561 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8562 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8563 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8564 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8565 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8566 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8567 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8568 a_664355_46657# a_662095_39580# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8569 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8570 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8571 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8572 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8573 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8574 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8575 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8576 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8577 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8578 a_722600_82134# a_719858_79988# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8579 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8580 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8581 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8582 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8583 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8584 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8585 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8586 a_663411_33525# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8587 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8588 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8589 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8590 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8591 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8592 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8593 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8594 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8595 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8596 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8597 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8598 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8599 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8600 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8601 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8602 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8603 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8604 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8605 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8606 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8607 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8608 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8609 w_661727_40249# a_650141_38543# a_650141_38543# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8610 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8611 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8612 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8613 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8614 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8615 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8616 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8617 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8618 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8619 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8620 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8621 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8622 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8623 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8624 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8625 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8626 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8627 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8628 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8629 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8630 w_649931_37947# a_663411_33525# a_663411_33525# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8631 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8632 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8633 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8634 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8635 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8636 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8637 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8638 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8639 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8640 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8641 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8642 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8643 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8644 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8645 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8646 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8647 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8648 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8649 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8650 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8651 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8652 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8653 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8654 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8655 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8656 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8657 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8658 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8659 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8660 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8661 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8662 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8663 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8664 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8665 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8666 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8667 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8668 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8669 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8670 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X8671 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8672 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8673 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8674 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8675 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8676 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8677 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8678 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8679 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8680 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8681 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8682 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8683 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8684 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8685 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8686 w_692190_39881# a_664155_35747# a_692386_37781# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8687 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8688 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8689 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8690 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8691 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8692 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8693 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8694 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8695 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8696 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8697 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8698 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8699 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8700 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8701 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8702 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8703 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8704 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8705 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8706 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8707 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8708 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8709 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8710 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8711 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8712 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8713 a_677477_59407# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8714 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8715 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8716 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8717 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8718 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8719 a_675258_42633# a_676490_42951# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X8720 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8721 a_678421_20774# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8722 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8723 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8724 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8725 w_649931_37947# a_677477_25371# a_678421_20774# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8726 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8727 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8728 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8729 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8730 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8731 w_649931_37947# a_719900_5846# a_725512_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8732 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8733 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8734 w_677281_20555# a_664155_35747# a_678421_20774# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8735 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8736 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8737 w_693353_61507# a_682038_37869# a_693549_59407# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8738 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8739 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8740 w_649931_37947# a_693549_59407# a_694493_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8741 a_694493_59495# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8742 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8743 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8744 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8745 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8746 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8747 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8748 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8749 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8750 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8751 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8752 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8753 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8754 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8755 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8756 w_661727_40249# a_650141_46551# a_650141_46551# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8757 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8758 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8759 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8760 a_693330_37869# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8761 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8762 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8763 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8764 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8765 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8766 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8767 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8768 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8769 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8770 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8771 w_649931_37947# a_677477_25371# a_678421_20774# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8772 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8773 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8774 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8775 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8776 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8777 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8778 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8779 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8780 a_679806_37869# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8781 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8782 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8783 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8784 a_650141_46551# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8785 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8786 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8787 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8788 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8789 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8790 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8791 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8792 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8793 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8794 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8795 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8796 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8797 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8798 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8799 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8800 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8801 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8802 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8803 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8804 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8805 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X8806 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8807 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8808 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8809 a_650141_39687# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8810 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8811 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8812 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8813 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8814 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8815 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8816 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8817 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8818 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8819 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8820 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8821 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8822 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8823 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8824 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8825 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8826 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8827 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8828 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8829 w_649931_37947# a_663411_51254# a_664355_46657# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8830 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8831 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8832 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8833 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8834 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8835 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8836 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8837 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8838 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8839 a_692386_37781# a_664155_35747# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8840 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8841 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8842 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8843 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8844 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8845 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8846 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8847 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8848 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8849 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8850 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8851 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8852 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8853 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8854 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8855 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8856 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8857 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8858 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8859 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8860 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8861 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8862 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8863 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8864 a_725512_n974# a_719742_7264# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8865 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8866 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8867 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8868 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8869 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8870 w_649931_37947# a_719900_80508# a_725512_73584# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8871 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8872 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8873 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8874 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8875 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8876 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8877 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8878 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8879 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8880 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8881 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8882 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8883 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8884 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8885 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8886 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8887 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8888 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8889 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8890 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8891 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8892 a_650141_45407# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8893 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8894 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8895 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8896 a_692386_37781# a_664155_35747# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8897 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8898 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8899 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8900 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8901 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8902 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8903 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8904 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8905 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8906 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8907 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8908 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8909 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8910 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X8911 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8912 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8913 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8914 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8915 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8916 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8917 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8918 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8919 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8920 a_663411_33525# a_662413_39580# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8921 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8922 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8923 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8924 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8925 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8926 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8927 a_664355_46657# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8928 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8929 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8930 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8931 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8932 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8933 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8934 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8935 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8936 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8937 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8938 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8939 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8940 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8941 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8942 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8943 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8944 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8945 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8946 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8947 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8948 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8949 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8950 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8951 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8952 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8953 w_649931_37947# a_650053_38143# a_650141_47695# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8954 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8955 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8956 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8957 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8958 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8959 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8960 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8961 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8962 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8963 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8964 a_673159_60085# a_674591_60403# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X8965 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8966 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8967 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8968 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8969 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8970 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8971 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8972 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8973 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8974 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X8975 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8976 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8977 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8978 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8979 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8980 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8981 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8982 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8983 a_673159_25299# a_674591_24981# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X8984 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8985 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8986 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8987 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8988 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8989 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8990 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8991 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8992 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X8993 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8994 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8995 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X8996 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8997 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8998 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8999 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9000 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9001 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9002 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9003 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9004 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9005 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9006 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9007 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9008 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9009 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9010 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9011 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9012 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9013 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9014 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9015 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9016 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9017 a_681073_22635# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=1.4e+07u
X9018 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9019 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9020 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9021 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9022 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9023 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9024 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9025 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9026 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9027 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9028 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9029 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9030 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9031 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9032 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9033 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9034 a_679806_37869# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9035 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9036 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9037 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9038 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9039 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9040 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9041 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9042 a_650141_47695# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9043 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9044 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9045 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9046 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9047 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9048 a_719742_79090# a_722600_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9049 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9050 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9051 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9052 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9053 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9054 a_693549_25370# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9055 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9056 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9057 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9058 w_692190_39881# a_693130_40003# a_693330_37869# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9059 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9060 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9061 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9062 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9063 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9064 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9065 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9066 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9067 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9068 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9069 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9070 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9071 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9072 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9073 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9074 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9075 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9076 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9077 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9078 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9079 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9080 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9081 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9082 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9083 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9084 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9085 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9086 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9087 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9088 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9089 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9090 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9091 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9092 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9093 w_677281_61507# a_673159_61357# a_677477_59407# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9094 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9095 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9096 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9097 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9098 w_677281_20555# a_673159_24981# a_677477_25371# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9099 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9100 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9101 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9102 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9103 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9104 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9105 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9106 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9107 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9108 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9109 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9110 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9111 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9112 w_649931_37947# a_650053_38143# a_650141_44263# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9113 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9114 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9115 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9116 a_678421_20774# a_664155_35747# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9117 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9118 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9119 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9120 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9121 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9122 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9123 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9124 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9125 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9126 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9127 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9128 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9129 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9130 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9131 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9132 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9133 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9134 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9135 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9136 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9137 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9138 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9139 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9140 w_649931_37947# a_663411_51254# a_663411_51254# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9141 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9142 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9143 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9144 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9145 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9146 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9147 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9148 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9149 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9150 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9151 a_679806_37869# a_664155_35747# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9152 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9153 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9154 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9155 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9156 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9157 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9158 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9159 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9160 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9161 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9162 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9163 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9164 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9165 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9166 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9167 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9168 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9169 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9170 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9171 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9172 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9173 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9174 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9175 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9176 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9177 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9178 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9179 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9180 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9181 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9182 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9183 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9184 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9185 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9186 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9187 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9188 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9189 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9190 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9191 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9192 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9193 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9194 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9195 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9196 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9197 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9198 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9199 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9200 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9201 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9202 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9203 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9204 a_693549_59407# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9205 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9206 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9207 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9208 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9209 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9210 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9211 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9212 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9213 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9214 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9215 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9216 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9217 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9218 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9219 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9220 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9221 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9222 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9223 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9224 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9225 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9226 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X9227 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9228 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9229 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9230 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9231 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9232 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9233 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9234 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9235 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9236 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9237 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9238 w_663215_35625# a_662413_39580# a_663411_33525# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9239 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9240 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9241 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9242 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9243 a_722600_82134# a_719858_79988# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9244 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9245 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9246 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9247 a_678421_59495# a_677477_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9248 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9249 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9250 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9251 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9252 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9253 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9254 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9255 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9256 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9257 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9258 w_649931_37947# a_677477_59407# a_678421_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9259 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9260 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9261 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9262 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9263 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9264 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9265 w_661727_40249# a_650141_41975# a_650141_41975# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9266 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9267 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9268 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9269 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9270 a_725512_82134# a_719742_79090# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9271 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9272 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9273 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9274 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9275 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9276 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9277 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9278 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9279 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9280 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9281 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9282 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9283 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9284 a_694493_59495# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9285 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9286 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9287 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9288 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9289 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9290 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9291 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9292 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9293 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9294 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9295 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9296 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9297 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9298 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9299 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9300 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9301 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9302 w_649931_37947# a_663411_33525# a_664355_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9303 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9304 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9305 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9306 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9307 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9308 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9309 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9310 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9311 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9312 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9313 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9314 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9315 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9316 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9317 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9318 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9319 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9320 a_677477_25371# a_673159_24981# w_677281_20555# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9321 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9322 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9323 a_678421_20774# a_677477_25371# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9324 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9325 w_649931_37947# a_678862_37781# a_679806_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9326 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9327 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9328 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9329 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9330 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9331 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9332 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9333 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9334 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9335 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9336 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9337 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9338 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9339 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9340 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9341 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9342 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9343 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9344 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9345 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9346 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9347 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9348 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9349 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9350 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9351 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9352 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9353 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9354 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9355 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9356 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9357 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9358 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9359 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9360 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9361 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9362 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9363 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9364 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9365 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9366 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9367 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9368 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9369 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9370 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9371 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9372 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9373 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9374 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9375 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9376 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9377 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9378 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9379 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9380 w_649931_37947# a_650053_38143# a_650053_38143# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9381 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9382 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9383 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9384 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9385 a_719858_6830# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9386 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9387 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9388 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9389 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9390 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9391 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9392 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9393 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9394 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9395 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9396 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9397 w_649931_37947# a_719742_79090# a_725512_82134# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9398 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9399 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9400 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9401 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9402 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9403 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9404 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9405 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9406 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9407 a_650141_39687# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9408 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9409 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9410 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9411 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9412 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9413 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9414 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9415 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9416 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9417 w_649931_37947# a_693549_59407# a_694493_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9418 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9419 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9420 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9421 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9422 w_693353_20554# a_680653_25459# a_694493_20773# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9423 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9424 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9425 w_649931_37947# a_722600_2050# a_719742_7264# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9426 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9427 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9428 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9429 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9430 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9431 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9432 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9433 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9434 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9435 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9436 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9437 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9438 a_693549_25370# a_682038_37869# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9439 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9440 a_650053_38143# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9441 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9442 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9443 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9444 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9445 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9446 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9447 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9448 a_663411_33525# a_662413_39580# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9449 w_678666_39881# a_664155_35747# a_679806_37869# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9450 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9451 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9452 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9453 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9454 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9455 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9456 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9457 w_649931_37947# a_663411_51254# a_663411_51254# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9458 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9459 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9460 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9461 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9462 w_692190_39881# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9463 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9464 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9465 a_719332_79990# a_696725_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9466 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9467 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9468 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9469 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9470 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9471 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9472 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9473 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9474 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9475 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9476 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9477 w_678666_39881# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9478 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9479 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9480 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9481 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9482 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9483 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9484 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9485 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9486 w_677281_61507# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9487 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9488 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9489 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9490 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9491 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9492 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9493 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9494 w_649931_37947# a_693549_59407# a_693549_59407# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9495 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9496 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9497 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9498 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9499 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9500 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9501 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9502 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9503 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9504 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9505 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9506 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9507 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9508 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9509 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9510 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9511 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9512 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9513 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9514 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9515 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9516 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9517 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9518 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9519 a_663411_33525# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9520 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9521 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9522 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9523 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9524 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9525 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9526 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9527 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9528 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9529 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9530 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9531 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9532 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9533 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9534 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9535 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9536 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9537 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9538 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9539 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9540 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9541 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9542 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9543 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9544 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9545 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9546 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9547 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9548 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9549 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9550 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9551 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9552 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9553 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9554 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9555 a_693549_59407# a_682038_37869# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9556 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9557 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9558 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9559 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9560 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9561 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9562 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9563 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9564 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9565 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9566 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9567 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9568 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9569 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9570 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9571 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9572 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9573 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9574 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9575 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9576 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9577 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9578 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9579 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9580 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9581 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9582 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9583 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9584 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9585 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9586 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9587 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9588 w_663215_35625# a_664155_35747# a_664355_33613# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9589 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9590 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9591 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9592 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9593 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9594 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9595 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9596 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9597 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9598 a_678862_37781# a_676490_44223# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9599 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9600 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9601 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9602 a_719858_5404# a_719332_5566# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X9603 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9604 a_719742_7264# a_722600_2050# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9605 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9606 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9607 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9608 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9609 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9610 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9611 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9612 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9613 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9614 a_693549_25370# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9615 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9616 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9617 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9618 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9619 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9620 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9621 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9622 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9623 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9624 w_661727_40249# a_650141_44263# w_692190_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9625 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9626 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9627 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9628 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9629 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9630 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9631 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9632 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9633 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9634 w_693353_20554# a_680653_25459# a_694493_20773# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9635 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9636 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9637 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9638 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9639 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9640 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9641 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9642 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9643 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9644 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9645 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9646 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9647 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9648 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9649 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9650 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9651 a_663411_51254# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9652 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9653 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9654 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9655 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9656 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9657 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9658 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9659 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9660 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9661 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9662 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9663 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9664 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9665 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9666 a_678862_37781# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9667 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9668 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9669 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9670 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9671 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9672 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9673 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9674 w_677281_20555# a_664155_35747# a_678421_20774# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9675 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X9676 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9677 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9678 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9679 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9680 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9681 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9682 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9683 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9684 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9685 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9686 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9687 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9688 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9689 a_666587_33613# a_664355_33613# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9690 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9691 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9692 a_694493_20773# a_693549_25370# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9693 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9694 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9695 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9696 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9697 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9698 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9699 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9700 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9701 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9702 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9703 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9704 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9705 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9706 w_663215_35625# a_664155_35747# a_664355_33613# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9707 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9708 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9709 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9710 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9711 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9712 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9713 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9714 a_719742_79090# a_722600_82134# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9715 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9716 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9717 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9718 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9719 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9720 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9721 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9722 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9723 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9724 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9725 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9726 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9727 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9728 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9729 a_678862_37781# a_678862_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9730 a_663411_51254# a_663411_46560# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9731 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9732 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9733 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9734 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9735 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9736 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9737 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9738 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X9739 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9740 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9741 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9742 a_693330_37869# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9743 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9744 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9745 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9746 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9747 a_675315_85767# a_675633_87199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X9748 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9749 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9750 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9751 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9752 w_693353_61507# a_680653_59495# a_694493_59495# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9753 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9754 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9755 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9756 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9757 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9758 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9759 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9760 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9761 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9762 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9763 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9764 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9765 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X9766 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9767 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9768 a_725512_82134# a_719742_79090# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9769 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9770 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9771 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9772 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9773 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9774 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9775 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9776 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9777 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9778 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9779 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9780 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9781 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9782 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9783 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9784 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9785 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9786 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9787 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9788 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9789 a_650141_38543# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9790 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9791 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9792 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9793 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9794 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9795 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9796 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9797 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9798 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9799 w_719104_5922# a_722600_75208# a_719900_80508# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9800 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9801 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9802 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9803 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9804 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9805 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9806 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9807 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9808 a_675633_n1233# a_675315_199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X9809 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9810 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9811 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9812 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9813 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9814 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9815 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9816 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9817 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9818 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9819 w_649931_37947# a_719742_79090# a_725512_82134# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9820 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9821 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9822 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9823 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9824 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9825 w_649931_37947# a_693549_25370# a_694493_20773# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9826 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9827 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9828 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9829 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9830 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9831 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9832 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9833 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9834 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9835 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9836 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9837 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9838 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9839 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9840 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9841 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9842 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9843 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9844 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9845 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9846 w_649931_37947# a_650053_38143# a_650141_39687# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9847 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9848 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9849 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9850 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9851 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9852 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9853 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9854 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9855 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9856 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9857 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9858 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9859 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9860 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9861 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9862 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9863 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9864 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9865 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9866 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9867 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9868 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9869 a_664355_33613# a_664155_35747# w_663215_35625# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9870 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9871 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9872 a_693330_37869# a_693130_40003# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9873 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9874 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9875 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9876 w_649931_37947# a_692386_37781# a_693330_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9877 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9878 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9879 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9880 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9881 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9882 a_676490_44223# a_682038_37869# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X9883 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9884 w_693353_61507# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9885 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9886 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9887 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9888 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9889 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9890 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9891 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9892 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9893 w_719104_5922# a_722600_8976# a_719900_5846# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9894 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9895 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9896 w_661727_40249# a_650141_40831# a_650141_40831# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9897 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9898 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9899 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9900 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9901 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9902 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9903 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9904 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9905 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9906 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9907 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9908 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9909 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9910 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9911 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9912 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9913 w_649931_37947# a_677477_59407# a_678421_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9914 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9915 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9916 a_696725_59495# a_694493_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9917 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9918 a_725512_8976# a_719900_5846# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9919 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9920 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9921 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9922 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9923 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9924 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9925 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9926 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9927 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9928 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9929 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9930 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9931 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9932 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9933 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9934 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9935 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9936 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9937 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9938 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9939 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9940 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9941 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9942 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9943 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9944 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9945 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9946 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9947 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9948 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9949 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9950 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9951 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9952 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9953 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9954 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9955 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9956 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9957 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9958 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X9959 a_693330_37869# a_697520_41473# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=500000u
X9960 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9961 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9962 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9963 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9964 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9965 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9966 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X9967 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9968 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9969 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9970 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9971 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9972 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9973 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9974 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9975 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9976 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9977 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9978 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9979 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9980 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9981 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9982 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9983 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9984 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9985 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9986 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9987 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9988 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9989 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9990 w_661727_40249# a_650141_46551# a_680653_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9991 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9992 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9993 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9994 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9995 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9996 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9997 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9998 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9999 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10000 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10001 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10002 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10003 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10004 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10005 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10006 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10007 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10008 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10009 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10010 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10011 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10012 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10013 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10014 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10015 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10016 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10017 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10018 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10019 w_649931_37947# a_679806_37869# a_682038_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10020 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10021 a_719858_7450# a_719742_7264# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10022 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10023 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10024 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10025 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10026 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10027 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10028 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10029 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10030 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10031 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10032 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10033 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10034 a_673159_59449# a_674591_59767# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10035 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10036 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10037 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10038 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10039 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10040 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10041 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10042 a_725512_73584# a_719900_80508# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10043 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10044 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10045 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10046 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10047 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10048 a_719900_80508# a_722600_75208# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10049 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10050 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10051 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10052 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10053 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10054 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10055 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10056 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10057 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10058 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10059 w_649931_37947# a_693549_25370# a_693549_25370# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10060 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10061 w_649931_37947# a_719742_7264# a_725512_n974# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10062 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10063 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10064 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10065 w_663215_35625# a_662413_39580# a_663411_33525# w_663215_35625# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10066 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10067 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10068 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10069 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10070 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10071 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10072 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10073 w_719104_5922# a_722600_2050# a_719742_7264# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10074 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10075 a_679806_37869# a_664155_35747# w_678666_39881# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10076 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10077 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10078 a_673159_61357# a_674591_61039# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10079 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10080 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10081 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10082 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10083 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10084 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10085 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10086 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10087 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10088 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10089 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10090 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10091 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10092 a_678421_59495# a_664155_35747# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10093 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10094 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10095 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10096 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10097 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10098 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10099 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10100 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10101 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10102 w_649931_37947# a_693549_25370# a_693549_25370# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10103 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10104 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10105 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10106 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10107 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10108 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10109 w_649931_37947# a_719742_7264# a_725512_n974# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10110 a_697520_41473# a_676490_41997# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=1.4e+07u
X10111 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10112 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10113 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10114 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10115 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10116 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10117 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10118 a_694493_59495# a_680653_59495# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10119 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10120 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10121 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10122 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10123 a_673159_61357# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X10124 w_661727_40249# a_650141_41975# a_682038_37869# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10125 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10126 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10127 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10128 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10129 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10130 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10131 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10132 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10133 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10134 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10135 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10136 w_649931_37947# a_650053_38143# a_650141_44263# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X10137 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10138 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10139 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10140 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10141 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10142 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10143 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10144 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10145 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10146 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10147 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10148 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10149 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10150 w_649931_37947# a_692386_37781# a_692386_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10151 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10152 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10153 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10154 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10155 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10156 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10157 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10158 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10159 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10160 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10161 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10162 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10163 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10164 w_661727_40249# a_650141_47695# w_693353_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10165 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10166 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10167 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10168 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10169 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10170 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10171 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10172 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10173 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10174 w_661727_40249# a_650141_41975# w_678666_39881# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10175 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10176 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10177 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10178 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10179 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10180 a_681073_22635# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=3e+07u
X10181 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10182 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10183 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10184 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10185 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10186 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10187 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10188 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10189 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10190 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10191 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10192 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10193 a_696725_59495# a_650141_47695# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10194 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10195 w_693353_20554# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10196 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10197 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10198 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10199 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10200 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10201 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10202 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10203 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10204 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10205 w_719104_5922# a_722600_75208# a_719900_80508# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10206 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10207 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10208 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10209 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10210 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10211 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10212 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10213 a_681073_63341# a_680653_59495# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=1.4e+07u
X10214 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10215 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10216 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10217 w_649931_37947# a_678862_37781# a_678862_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10218 w_677281_61507# a_664155_35747# a_678421_59495# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10219 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10220 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10221 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10222 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10223 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10224 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10225 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10226 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10227 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10228 a_694493_20773# a_680653_25459# w_693353_20554# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10229 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10230 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10231 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10232 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10233 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10234 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10235 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10236 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10237 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10238 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10239 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10240 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10241 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10242 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10243 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10244 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10245 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10246 a_696725_25458# a_650141_38543# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10247 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10248 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10249 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10250 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10251 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10252 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10253 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10254 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10255 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10256 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10257 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10258 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10259 w_663215_46438# a_663411_46560# a_663411_51254# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10260 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10261 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10262 a_719332_5566# a_696725_25458# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10263 a_650141_40831# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10264 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10265 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10266 a_650141_41975# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10267 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10268 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10269 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10270 w_661727_40249# a_650141_45407# a_663411_46560# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10271 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10272 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10273 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10274 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10275 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10276 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10277 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10278 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10279 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10280 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10281 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10282 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10283 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10284 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10285 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10286 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10287 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10288 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10289 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10290 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10291 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10292 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10293 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10294 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10295 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10296 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10297 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10298 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10299 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10300 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10301 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10302 w_693353_61507# a_682038_37869# a_693549_59407# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10303 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10304 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10305 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10306 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10307 w_677281_20555# a_673159_24981# a_677477_25371# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10308 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10309 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10310 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10311 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10312 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10313 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10314 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10315 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10316 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10317 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10318 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10319 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10320 w_649931_37947# a_663411_51254# a_664355_46657# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10321 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10322 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10323 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10324 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10325 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10326 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10327 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10328 a_676490_41997# a_693330_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10329 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10330 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10331 w_678666_39881# a_664155_35747# a_679806_37869# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10332 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10333 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10334 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10335 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10336 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10337 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10338 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10339 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10340 w_678666_39881# a_676490_44223# a_678862_37781# w_678666_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10341 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10342 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10343 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10344 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10345 a_664355_46657# a_662095_39580# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10346 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10347 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10348 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10349 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10350 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10351 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10352 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10353 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10354 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10355 a_650141_44263# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10356 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10357 w_661727_40249# a_650141_40831# a_666587_33613# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10358 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10359 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10360 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10361 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10362 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10363 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10364 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10365 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10366 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10367 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10368 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10369 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10370 a_650141_44263# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X10371 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10372 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10373 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10374 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10375 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10376 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10377 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10378 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10379 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10380 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10381 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10382 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10383 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10384 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10385 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10386 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10387 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10388 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10389 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10390 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10391 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10392 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10393 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10394 w_661727_40249# a_650141_44263# a_676490_41997# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10395 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10396 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10397 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10398 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10399 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10400 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10401 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10402 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10403 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10404 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10405 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10406 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10407 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10408 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10409 w_649931_37947# a_725512_8976# a_730362_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10410 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10411 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10412 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10413 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10414 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10415 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10416 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10417 a_664355_33613# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10418 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10419 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10420 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10421 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10422 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10423 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10424 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10425 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10426 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10427 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10428 w_649931_37947# a_694493_59495# a_696725_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10429 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10430 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10431 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10432 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10433 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10434 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10435 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10436 a_650053_38143# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X10437 a_682038_37869# a_679806_37869# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10438 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10439 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10440 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10441 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10442 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10443 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10444 w_649931_37947# a_719900_5846# a_725512_8976# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10445 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10446 a_680653_25459# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10447 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10448 w_693353_20554# a_682038_37869# a_693549_25370# w_693353_20554# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10449 a_725512_73584# a_719900_80508# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10450 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10451 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10452 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10453 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10454 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10455 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10456 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10457 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10458 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10459 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10460 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10461 w_663215_35625# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10462 a_693549_59407# a_682038_37869# w_693353_61507# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10463 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10464 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10465 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10466 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10467 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10468 a_673159_24981# a_680653_25459# sky130_fd_pr__cap_mim_m3_1 l=1.75e+07u w=1.75e+07u
X10469 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10470 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10471 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10472 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10473 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10474 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10475 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10476 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10477 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10478 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10479 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10480 a_663411_51254# a_663411_46560# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10481 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10482 a_680653_25459# a_678421_20774# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10483 a_719858_6024# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10484 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10485 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10486 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10487 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10488 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10489 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10490 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10491 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10492 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10493 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10494 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10495 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10496 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10497 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10498 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10499 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10500 w_692190_39881# a_664155_35747# a_692386_37781# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10501 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10502 a_677477_59407# a_673159_61357# w_677281_61507# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10503 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10504 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10505 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10506 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10507 w_649931_37947# a_677477_25371# a_677477_25371# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10508 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10509 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10510 w_661727_40249# a_650141_39687# a_650141_39687# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10511 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10512 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10513 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10514 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10515 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10516 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10517 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10518 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10519 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10520 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10521 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10522 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10523 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10524 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10525 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10526 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10527 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10528 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10529 a_719858_79988# a_719332_79990# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10530 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10531 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10532 w_719104_5922# a_719742_7264# a_725512_n974# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10533 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10534 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10535 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10536 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10537 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10538 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10539 w_719104_5922# a_719900_80508# a_725512_73584# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10540 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10541 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10542 w_649931_37947# a_693330_37869# a_676490_41997# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10543 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10544 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10545 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10546 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10547 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10548 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10549 a_663411_51254# a_663411_51254# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10550 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10551 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10552 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10553 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10554 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10555 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10556 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10557 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10558 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10559 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10560 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10561 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10562 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10563 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10564 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10565 a_676490_41997# a_650141_44263# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10566 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10567 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10568 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10569 w_649931_37947# a_692386_37781# a_692386_37781# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10570 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10571 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10572 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10573 a_692386_37781# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10574 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10575 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10576 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10577 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10578 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10579 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10580 a_725512_8976# a_719900_5846# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10581 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10582 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10583 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10584 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10585 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10586 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10587 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10588 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10589 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10590 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10591 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10592 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10593 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10594 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10595 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10596 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10597 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10598 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10599 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10600 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10601 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10602 w_649931_37947# a_678421_20774# a_680653_25459# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10603 a_682038_37869# a_650141_41975# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10604 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10605 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10606 w_661727_40249# a_650141_45407# a_650141_45407# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10607 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10608 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10609 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10610 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10611 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10612 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10613 w_692190_39881# a_693130_40003# a_693330_37869# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10614 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10615 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10616 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10617 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10618 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10619 a_680653_59495# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10620 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10621 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10622 w_649931_37947# a_663411_33525# a_663411_33525# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10623 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10624 w_663215_46438# a_662095_39580# a_664355_46657# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10625 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10626 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10627 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10628 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10629 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10630 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10631 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10632 w_663215_46438# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10633 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10634 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10635 a_664355_33613# a_663411_33525# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10636 a_696725_25458# a_694493_20773# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10637 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10638 a_664355_46657# a_662095_39580# w_663215_46438# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10639 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10640 a_680653_59495# a_678421_59495# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10641 w_661727_40249# a_650141_39687# a_680653_25459# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10642 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10643 a_650141_46551# a_650141_46551# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10644 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10645 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10646 w_649931_37947# a_677477_25371# a_677477_25371# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10647 w_661727_40249# a_650141_47695# a_696725_59495# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10648 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10649 w_677281_20555# a_673159_24981# a_677477_25371# w_677281_20555# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10650 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10651 w_693353_61507# a_680653_59495# a_694493_59495# w_693353_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10652 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10653 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10654 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10655 w_719104_5922# a_725512_73584# a_730362_67500# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10656 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10657 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10658 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10659 w_661727_40249# a_650141_39687# w_677281_20555# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10660 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10661 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10662 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10663 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10664 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10665 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10666 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10667 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10668 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10669 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10670 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10671 w_661727_40249# a_650141_38543# w_693353_20554# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10672 w_661727_40249# a_650141_46551# w_677281_61507# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10673 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10674 a_650141_41975# a_650053_38143# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X10675 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10676 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10677 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10678 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10679 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10680 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10681 w_649931_37947# a_719742_7264# a_725512_n974# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10682 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10683 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10684 w_661727_40249# a_650141_44263# a_650141_44263# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10685 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10686 w_649931_37947# a_677477_25371# a_677477_25371# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10687 a_692386_37781# a_664155_35747# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10688 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10689 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10690 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10691 w_677281_61507# a_664155_35747# a_678421_59495# w_677281_61507# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10692 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10693 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10694 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10695 w_649931_37947# a_678862_37781# a_679806_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10696 a_730362_67500# a_725512_73584# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10697 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10698 w_677281_20555# a_650141_39687# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10699 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10700 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10701 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10702 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10703 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10704 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10705 w_649931_37947# a_725512_73584# a_730362_67500# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10706 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10707 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10708 w_661727_40249# a_650141_47695# a_650141_47695# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10709 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10710 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10711 a_673159_25935# a_674591_26253# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10712 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10713 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10714 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10715 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10716 w_661727_40249# a_650141_38543# a_696725_25458# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10717 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10718 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10719 w_719104_5922# a_719900_5846# a_725512_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10720 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10721 w_719104_5922# a_719742_79090# a_725512_82134# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10722 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10723 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10724 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10725 a_719742_79090# a_722600_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10726 a_719858_79988# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10727 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10728 a_663411_46560# a_664355_46657# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10729 w_719104_5922# a_725512_8976# a_730362_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10730 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10731 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10732 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10733 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10734 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10735 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10736 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10737 a_693549_59407# a_693549_59407# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10738 w_719104_5922# a_719858_6830# a_722600_8976# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10739 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10740 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10741 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10742 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10743 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10744 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10745 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10746 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10747 a_666587_33613# a_650141_40831# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10748 w_649931_37947# a_664355_46657# a_663411_46560# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10749 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10750 w_649931_37947# w_719104_5922# sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.6e+07u
X10751 a_693330_37869# a_693130_40003# w_692190_39881# w_692190_39881# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10752 a_692386_37781# a_692386_37781# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10753 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10754 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10755 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10756 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10757 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10758 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10759 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10760 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10761 w_649931_37947# a_692386_37781# a_693330_37869# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10762 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10763 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10764 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10765 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10766 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10767 a_650053_38143# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10768 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10769 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10770 a_676905_87199# a_725512_82134# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10771 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10772 w_661727_40249# a_650141_40831# w_663215_35625# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10773 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10774 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10775 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10776 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10777 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10778 a_730362_8976# a_725512_8976# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10779 a_663411_46560# a_650141_45407# w_661727_40249# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10780 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10781 w_661727_40249# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10782 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10783 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10784 a_673159_61357# a_674997_87199# w_649931_37947# sky130_fd_pr__res_xhigh_po w=350000u l=5e+06u
X10785 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10786 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10787 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10788 a_730362_67500# a_725512_73584# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10789 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10790 a_719858_79182# w_649931_37947# sky130_fd_pr__cap_mim_m3_1 l=1.775e+07u w=1.775e+07u
X10791 w_649931_37947# a_650053_38143# a_650141_40831# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X10792 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10793 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10794 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10795 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10796 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10797 a_725512_73584# a_719900_80508# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10798 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10799 a_676905_n1233# a_725512_n974# w_649931_37947# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10800 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10801 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10802 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10803 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10804 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10805 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10806 a_676905_n1233# a_730362_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10807 w_719104_5922# w_649931_37947# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
X10808 w_649931_37947# a_725512_82134# a_676905_87199# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10809 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10810 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10811 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10812 a_730362_8976# a_725512_8976# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10813 w_661727_40249# a_650141_45407# w_663215_46438# w_661727_40249# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10814 w_649931_37947# a_664355_33613# a_666587_33613# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10815 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10816 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10817 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10818 w_649931_37947# a_694493_20773# a_696725_25458# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10819 w_663215_46438# a_663411_46560# a_663411_51254# w_663215_46438# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10820 w_649931_37947# a_650053_38143# a_650141_39687# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X10821 w_649931_37947# a_725512_n974# a_676905_n1233# w_649931_37947# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10822 a_676905_87199# a_730362_67500# w_719104_5922# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10823 w_649931_37947# a_678421_59495# a_680653_59495# w_649931_37947# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10824 w_719104_5922# a_730362_8976# a_676905_n1233# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10825 w_719104_5922# a_730362_67500# a_676905_87199# w_719104_5922# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
.end

