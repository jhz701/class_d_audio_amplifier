magic
tech sky130A
magscale 1 2
timestamp 1627023368
<< nwell >>
rect -6920 -876 22100 2988
rect 6092 -5416 9088 -1386
<< pwell >>
rect 2384 4554 12798 7190
rect 13577 -5087 13979 -3331
rect 6704 -8194 8478 -5578
<< pmoslvt >>
rect -6428 1656 -6028 2456
rect -5840 1656 -5440 2456
rect -5252 1656 -4852 2456
rect -4664 1656 -4264 2456
rect -4076 1656 -3676 2456
rect -3488 1656 -3088 2456
rect -2900 1656 -2500 2456
rect -2312 1656 -1912 2456
rect -1724 1656 -1324 2456
rect -1136 1656 -736 2456
rect -548 1656 -148 2456
rect 40 1656 440 2456
rect 628 1656 1028 2456
rect 1216 1656 1616 2456
rect 1804 1656 2204 2456
rect 2392 1656 2792 2456
rect 2980 1656 3380 2456
rect 3568 1656 3968 2456
rect 4156 1656 4556 2456
rect 4744 1656 5144 2456
rect 5332 1656 5732 2456
rect 5920 1656 6320 2456
rect 6508 1656 6908 2456
rect 7096 1656 7496 2456
rect 7684 1656 8084 2456
rect 8272 1656 8672 2456
rect 8860 1656 9260 2456
rect 9448 1656 9848 2456
rect 10036 1656 10436 2456
rect 10624 1656 11024 2456
rect 11212 1656 11612 2456
rect 11800 1656 12200 2456
rect 12388 1656 12788 2456
rect 12976 1656 13376 2456
rect 13564 1656 13964 2456
rect 14152 1656 14552 2456
rect 14740 1656 15140 2456
rect 15328 1656 15728 2456
rect 15916 1656 16316 2456
rect 16504 1656 16904 2456
rect 17092 1656 17492 2456
rect 17680 1656 18080 2456
rect 18268 1656 18668 2456
rect 18856 1656 19256 2456
rect 19444 1656 19844 2456
rect 20032 1656 20432 2456
rect 20620 1656 21020 2456
rect 21208 1656 21608 2456
rect -6428 656 -6028 1456
rect -5840 656 -5440 1456
rect -5252 656 -4852 1456
rect -4664 656 -4264 1456
rect -4076 656 -3676 1456
rect -3488 656 -3088 1456
rect -2900 656 -2500 1456
rect -2312 656 -1912 1456
rect -1724 656 -1324 1456
rect -1136 656 -736 1456
rect -548 656 -148 1456
rect 40 656 440 1456
rect 628 656 1028 1456
rect 1216 656 1616 1456
rect 1804 656 2204 1456
rect 2392 656 2792 1456
rect 2980 656 3380 1456
rect 3568 656 3968 1456
rect 4156 656 4556 1456
rect 4744 656 5144 1456
rect 5332 656 5732 1456
rect 5920 656 6320 1456
rect 6508 656 6908 1456
rect 7096 656 7496 1456
rect 7684 656 8084 1456
rect 8272 656 8672 1456
rect 8860 656 9260 1456
rect 9448 656 9848 1456
rect 10036 656 10436 1456
rect 10624 656 11024 1456
rect 11212 656 11612 1456
rect 11800 656 12200 1456
rect 12388 656 12788 1456
rect 12976 656 13376 1456
rect 13564 656 13964 1456
rect 14152 656 14552 1456
rect 14740 656 15140 1456
rect 15328 656 15728 1456
rect 15916 656 16316 1456
rect 16504 656 16904 1456
rect 17092 656 17492 1456
rect 17680 656 18080 1456
rect 18268 656 18668 1456
rect 18856 656 19256 1456
rect 19444 656 19844 1456
rect 20032 656 20432 1456
rect 20620 656 21020 1456
rect 21208 656 21608 1456
rect -6428 -344 -6028 456
rect -5840 -344 -5440 456
rect -5252 -344 -4852 456
rect -4664 -344 -4264 456
rect -4076 -344 -3676 456
rect -3488 -344 -3088 456
rect -2900 -344 -2500 456
rect -2312 -344 -1912 456
rect -1724 -344 -1324 456
rect -1136 -344 -736 456
rect -548 -344 -148 456
rect 40 -344 440 456
rect 628 -344 1028 456
rect 1216 -344 1616 456
rect 1804 -344 2204 456
rect 2392 -344 2792 456
rect 2980 -344 3380 456
rect 3568 -344 3968 456
rect 4156 -344 4556 456
rect 4744 -344 5144 456
rect 5332 -344 5732 456
rect 5920 -344 6320 456
rect 6508 -344 6908 456
rect 7096 -344 7496 456
rect 7684 -344 8084 456
rect 8272 -344 8672 456
rect 8860 -344 9260 456
rect 9448 -344 9848 456
rect 10036 -344 10436 456
rect 10624 -344 11024 456
rect 11212 -344 11612 456
rect 11800 -344 12200 456
rect 12388 -344 12788 456
rect 12976 -344 13376 456
rect 13564 -344 13964 456
rect 14152 -344 14552 456
rect 14740 -344 15140 456
rect 15328 -344 15728 456
rect 15916 -344 16316 456
rect 16504 -344 16904 456
rect 17092 -344 17492 456
rect 17680 -344 18080 456
rect 18268 -344 18668 456
rect 18856 -344 19256 456
rect 19444 -344 19844 456
rect 20032 -344 20432 456
rect 20620 -344 21020 456
rect 21208 -344 21608 456
rect 6624 -2790 6694 -1990
rect 6890 -2790 6960 -1990
rect 7156 -2790 7226 -1990
rect 7422 -2790 7492 -1990
rect 7688 -2790 7758 -1990
rect 7954 -2790 8024 -1990
rect 8220 -2790 8290 -1990
rect 8486 -2790 8556 -1990
rect 6624 -3800 6694 -3000
rect 6890 -3800 6960 -3000
rect 7156 -3800 7226 -3000
rect 7422 -3800 7492 -3000
rect 7688 -3800 7758 -3000
rect 7954 -3800 8024 -3000
rect 8220 -3800 8290 -3000
rect 8486 -3800 8556 -3000
rect 6624 -4810 6694 -4010
rect 6890 -4810 6960 -4010
rect 7156 -4810 7226 -4010
rect 7422 -4810 7492 -4010
rect 7688 -4810 7758 -4010
rect 7954 -4810 8024 -4010
rect 8220 -4810 8290 -4010
rect 8486 -4810 8556 -4010
<< nmoslvt >>
rect 2876 5976 2946 6576
rect 3116 5976 3186 6576
rect 3356 5976 3426 6576
rect 3596 5976 3666 6576
rect 3836 5976 3906 6576
rect 4076 5976 4146 6576
rect 4316 5976 4386 6576
rect 4556 5976 4626 6576
rect 4796 5976 4866 6576
rect 5036 5976 5106 6576
rect 5276 5976 5346 6576
rect 5516 5976 5586 6576
rect 5756 5976 5826 6576
rect 5996 5976 6066 6576
rect 6236 5976 6306 6576
rect 6476 5976 6546 6576
rect 6716 5976 6786 6576
rect 6956 5976 7026 6576
rect 7196 5976 7266 6576
rect 7436 5976 7506 6576
rect 7676 5976 7746 6576
rect 7916 5976 7986 6576
rect 8156 5976 8226 6576
rect 8396 5976 8466 6576
rect 8636 5976 8706 6576
rect 8876 5976 8946 6576
rect 9116 5976 9186 6576
rect 9356 5976 9426 6576
rect 9596 5976 9666 6576
rect 9836 5976 9906 6576
rect 10076 5976 10146 6576
rect 10316 5976 10386 6576
rect 10556 5976 10626 6576
rect 10796 5976 10866 6576
rect 11036 5976 11106 6576
rect 11276 5976 11346 6576
rect 11516 5976 11586 6576
rect 11756 5976 11826 6576
rect 11996 5976 12066 6576
rect 12236 5976 12306 6576
rect 2876 5168 2946 5768
rect 3116 5168 3186 5768
rect 3356 5168 3426 5768
rect 3596 5168 3666 5768
rect 3836 5168 3906 5768
rect 4076 5168 4146 5768
rect 4316 5168 4386 5768
rect 4556 5168 4626 5768
rect 4796 5168 4866 5768
rect 5036 5168 5106 5768
rect 5276 5168 5346 5768
rect 5516 5168 5586 5768
rect 5756 5168 5826 5768
rect 5996 5168 6066 5768
rect 6236 5168 6306 5768
rect 6476 5168 6546 5768
rect 6716 5168 6786 5768
rect 6956 5168 7026 5768
rect 7196 5168 7266 5768
rect 7436 5168 7506 5768
rect 7676 5168 7746 5768
rect 7916 5168 7986 5768
rect 8156 5168 8226 5768
rect 8396 5168 8466 5768
rect 8636 5168 8706 5768
rect 8876 5168 8946 5768
rect 9116 5168 9186 5768
rect 9356 5168 9426 5768
rect 9596 5168 9666 5768
rect 9836 5168 9906 5768
rect 10076 5168 10146 5768
rect 10316 5168 10386 5768
rect 10556 5168 10626 5768
rect 10796 5168 10866 5768
rect 11036 5168 11106 5768
rect 11276 5168 11346 5768
rect 11516 5168 11586 5768
rect 11756 5168 11826 5768
rect 11996 5168 12066 5768
rect 12236 5168 12306 5768
rect 7196 -6782 7266 -6182
rect 7436 -6782 7506 -6182
rect 7676 -6782 7746 -6182
rect 7916 -6782 7986 -6182
rect 7196 -7590 7266 -6990
rect 7436 -7590 7506 -6990
rect 7676 -7590 7746 -6990
rect 7916 -7590 7986 -6990
<< ndiff >>
rect 2818 6564 2876 6576
rect 2818 5988 2830 6564
rect 2864 5988 2876 6564
rect 2818 5976 2876 5988
rect 2946 6564 3004 6576
rect 2946 5988 2958 6564
rect 2992 5988 3004 6564
rect 2946 5976 3004 5988
rect 3058 6564 3116 6576
rect 3058 5988 3070 6564
rect 3104 5988 3116 6564
rect 3058 5976 3116 5988
rect 3186 6564 3244 6576
rect 3186 5988 3198 6564
rect 3232 5988 3244 6564
rect 3186 5976 3244 5988
rect 3298 6564 3356 6576
rect 3298 5988 3310 6564
rect 3344 5988 3356 6564
rect 3298 5976 3356 5988
rect 3426 6564 3484 6576
rect 3426 5988 3438 6564
rect 3472 5988 3484 6564
rect 3426 5976 3484 5988
rect 3538 6564 3596 6576
rect 3538 5988 3550 6564
rect 3584 5988 3596 6564
rect 3538 5976 3596 5988
rect 3666 6564 3724 6576
rect 3666 5988 3678 6564
rect 3712 5988 3724 6564
rect 3666 5976 3724 5988
rect 3778 6564 3836 6576
rect 3778 5988 3790 6564
rect 3824 5988 3836 6564
rect 3778 5976 3836 5988
rect 3906 6564 3964 6576
rect 3906 5988 3918 6564
rect 3952 5988 3964 6564
rect 3906 5976 3964 5988
rect 4018 6564 4076 6576
rect 4018 5988 4030 6564
rect 4064 5988 4076 6564
rect 4018 5976 4076 5988
rect 4146 6564 4204 6576
rect 4146 5988 4158 6564
rect 4192 5988 4204 6564
rect 4146 5976 4204 5988
rect 4258 6564 4316 6576
rect 4258 5988 4270 6564
rect 4304 5988 4316 6564
rect 4258 5976 4316 5988
rect 4386 6564 4444 6576
rect 4386 5988 4398 6564
rect 4432 5988 4444 6564
rect 4386 5976 4444 5988
rect 4498 6564 4556 6576
rect 4498 5988 4510 6564
rect 4544 5988 4556 6564
rect 4498 5976 4556 5988
rect 4626 6564 4684 6576
rect 4626 5988 4638 6564
rect 4672 5988 4684 6564
rect 4626 5976 4684 5988
rect 4738 6564 4796 6576
rect 4738 5988 4750 6564
rect 4784 5988 4796 6564
rect 4738 5976 4796 5988
rect 4866 6564 4924 6576
rect 4866 5988 4878 6564
rect 4912 5988 4924 6564
rect 4866 5976 4924 5988
rect 4978 6564 5036 6576
rect 4978 5988 4990 6564
rect 5024 5988 5036 6564
rect 4978 5976 5036 5988
rect 5106 6564 5164 6576
rect 5106 5988 5118 6564
rect 5152 5988 5164 6564
rect 5106 5976 5164 5988
rect 5218 6564 5276 6576
rect 5218 5988 5230 6564
rect 5264 5988 5276 6564
rect 5218 5976 5276 5988
rect 5346 6564 5404 6576
rect 5346 5988 5358 6564
rect 5392 5988 5404 6564
rect 5346 5976 5404 5988
rect 5458 6564 5516 6576
rect 5458 5988 5470 6564
rect 5504 5988 5516 6564
rect 5458 5976 5516 5988
rect 5586 6564 5644 6576
rect 5586 5988 5598 6564
rect 5632 5988 5644 6564
rect 5586 5976 5644 5988
rect 5698 6564 5756 6576
rect 5698 5988 5710 6564
rect 5744 5988 5756 6564
rect 5698 5976 5756 5988
rect 5826 6564 5884 6576
rect 5826 5988 5838 6564
rect 5872 5988 5884 6564
rect 5826 5976 5884 5988
rect 5938 6564 5996 6576
rect 5938 5988 5950 6564
rect 5984 5988 5996 6564
rect 5938 5976 5996 5988
rect 6066 6564 6124 6576
rect 6066 5988 6078 6564
rect 6112 5988 6124 6564
rect 6066 5976 6124 5988
rect 6178 6564 6236 6576
rect 6178 5988 6190 6564
rect 6224 5988 6236 6564
rect 6178 5976 6236 5988
rect 6306 6564 6364 6576
rect 6306 5988 6318 6564
rect 6352 5988 6364 6564
rect 6306 5976 6364 5988
rect 6418 6564 6476 6576
rect 6418 5988 6430 6564
rect 6464 5988 6476 6564
rect 6418 5976 6476 5988
rect 6546 6564 6604 6576
rect 6546 5988 6558 6564
rect 6592 5988 6604 6564
rect 6546 5976 6604 5988
rect 6658 6564 6716 6576
rect 6658 5988 6670 6564
rect 6704 5988 6716 6564
rect 6658 5976 6716 5988
rect 6786 6564 6844 6576
rect 6786 5988 6798 6564
rect 6832 5988 6844 6564
rect 6786 5976 6844 5988
rect 6898 6564 6956 6576
rect 6898 5988 6910 6564
rect 6944 5988 6956 6564
rect 6898 5976 6956 5988
rect 7026 6564 7084 6576
rect 7026 5988 7038 6564
rect 7072 5988 7084 6564
rect 7026 5976 7084 5988
rect 7138 6564 7196 6576
rect 7138 5988 7150 6564
rect 7184 5988 7196 6564
rect 7138 5976 7196 5988
rect 7266 6564 7324 6576
rect 7266 5988 7278 6564
rect 7312 5988 7324 6564
rect 7266 5976 7324 5988
rect 7378 6564 7436 6576
rect 7378 5988 7390 6564
rect 7424 5988 7436 6564
rect 7378 5976 7436 5988
rect 7506 6564 7564 6576
rect 7506 5988 7518 6564
rect 7552 5988 7564 6564
rect 7506 5976 7564 5988
rect 7618 6564 7676 6576
rect 7618 5988 7630 6564
rect 7664 5988 7676 6564
rect 7618 5976 7676 5988
rect 7746 6564 7804 6576
rect 7746 5988 7758 6564
rect 7792 5988 7804 6564
rect 7746 5976 7804 5988
rect 7858 6564 7916 6576
rect 7858 5988 7870 6564
rect 7904 5988 7916 6564
rect 7858 5976 7916 5988
rect 7986 6564 8044 6576
rect 7986 5988 7998 6564
rect 8032 5988 8044 6564
rect 7986 5976 8044 5988
rect 8098 6564 8156 6576
rect 8098 5988 8110 6564
rect 8144 5988 8156 6564
rect 8098 5976 8156 5988
rect 8226 6564 8284 6576
rect 8226 5988 8238 6564
rect 8272 5988 8284 6564
rect 8226 5976 8284 5988
rect 8338 6564 8396 6576
rect 8338 5988 8350 6564
rect 8384 5988 8396 6564
rect 8338 5976 8396 5988
rect 8466 6564 8524 6576
rect 8466 5988 8478 6564
rect 8512 5988 8524 6564
rect 8466 5976 8524 5988
rect 8578 6564 8636 6576
rect 8578 5988 8590 6564
rect 8624 5988 8636 6564
rect 8578 5976 8636 5988
rect 8706 6564 8764 6576
rect 8706 5988 8718 6564
rect 8752 5988 8764 6564
rect 8706 5976 8764 5988
rect 8818 6564 8876 6576
rect 8818 5988 8830 6564
rect 8864 5988 8876 6564
rect 8818 5976 8876 5988
rect 8946 6564 9004 6576
rect 8946 5988 8958 6564
rect 8992 5988 9004 6564
rect 8946 5976 9004 5988
rect 9058 6564 9116 6576
rect 9058 5988 9070 6564
rect 9104 5988 9116 6564
rect 9058 5976 9116 5988
rect 9186 6564 9244 6576
rect 9186 5988 9198 6564
rect 9232 5988 9244 6564
rect 9186 5976 9244 5988
rect 9298 6564 9356 6576
rect 9298 5988 9310 6564
rect 9344 5988 9356 6564
rect 9298 5976 9356 5988
rect 9426 6564 9484 6576
rect 9426 5988 9438 6564
rect 9472 5988 9484 6564
rect 9426 5976 9484 5988
rect 9538 6564 9596 6576
rect 9538 5988 9550 6564
rect 9584 5988 9596 6564
rect 9538 5976 9596 5988
rect 9666 6564 9724 6576
rect 9666 5988 9678 6564
rect 9712 5988 9724 6564
rect 9666 5976 9724 5988
rect 9778 6564 9836 6576
rect 9778 5988 9790 6564
rect 9824 5988 9836 6564
rect 9778 5976 9836 5988
rect 9906 6564 9964 6576
rect 9906 5988 9918 6564
rect 9952 5988 9964 6564
rect 9906 5976 9964 5988
rect 10018 6564 10076 6576
rect 10018 5988 10030 6564
rect 10064 5988 10076 6564
rect 10018 5976 10076 5988
rect 10146 6564 10204 6576
rect 10146 5988 10158 6564
rect 10192 5988 10204 6564
rect 10146 5976 10204 5988
rect 10258 6564 10316 6576
rect 10258 5988 10270 6564
rect 10304 5988 10316 6564
rect 10258 5976 10316 5988
rect 10386 6564 10444 6576
rect 10386 5988 10398 6564
rect 10432 5988 10444 6564
rect 10386 5976 10444 5988
rect 10498 6564 10556 6576
rect 10498 5988 10510 6564
rect 10544 5988 10556 6564
rect 10498 5976 10556 5988
rect 10626 6564 10684 6576
rect 10626 5988 10638 6564
rect 10672 5988 10684 6564
rect 10626 5976 10684 5988
rect 10738 6564 10796 6576
rect 10738 5988 10750 6564
rect 10784 5988 10796 6564
rect 10738 5976 10796 5988
rect 10866 6564 10924 6576
rect 10866 5988 10878 6564
rect 10912 5988 10924 6564
rect 10866 5976 10924 5988
rect 10978 6564 11036 6576
rect 10978 5988 10990 6564
rect 11024 5988 11036 6564
rect 10978 5976 11036 5988
rect 11106 6564 11164 6576
rect 11106 5988 11118 6564
rect 11152 5988 11164 6564
rect 11106 5976 11164 5988
rect 11218 6564 11276 6576
rect 11218 5988 11230 6564
rect 11264 5988 11276 6564
rect 11218 5976 11276 5988
rect 11346 6564 11404 6576
rect 11346 5988 11358 6564
rect 11392 5988 11404 6564
rect 11346 5976 11404 5988
rect 11458 6564 11516 6576
rect 11458 5988 11470 6564
rect 11504 5988 11516 6564
rect 11458 5976 11516 5988
rect 11586 6564 11644 6576
rect 11586 5988 11598 6564
rect 11632 5988 11644 6564
rect 11586 5976 11644 5988
rect 11698 6564 11756 6576
rect 11698 5988 11710 6564
rect 11744 5988 11756 6564
rect 11698 5976 11756 5988
rect 11826 6564 11884 6576
rect 11826 5988 11838 6564
rect 11872 5988 11884 6564
rect 11826 5976 11884 5988
rect 11938 6564 11996 6576
rect 11938 5988 11950 6564
rect 11984 5988 11996 6564
rect 11938 5976 11996 5988
rect 12066 6564 12124 6576
rect 12066 5988 12078 6564
rect 12112 5988 12124 6564
rect 12066 5976 12124 5988
rect 12178 6564 12236 6576
rect 12178 5988 12190 6564
rect 12224 5988 12236 6564
rect 12178 5976 12236 5988
rect 12306 6564 12364 6576
rect 12306 5988 12318 6564
rect 12352 5988 12364 6564
rect 12306 5976 12364 5988
rect 2818 5756 2876 5768
rect 2818 5180 2830 5756
rect 2864 5180 2876 5756
rect 2818 5168 2876 5180
rect 2946 5756 3004 5768
rect 2946 5180 2958 5756
rect 2992 5180 3004 5756
rect 2946 5168 3004 5180
rect 3058 5756 3116 5768
rect 3058 5180 3070 5756
rect 3104 5180 3116 5756
rect 3058 5168 3116 5180
rect 3186 5756 3244 5768
rect 3186 5180 3198 5756
rect 3232 5180 3244 5756
rect 3186 5168 3244 5180
rect 3298 5756 3356 5768
rect 3298 5180 3310 5756
rect 3344 5180 3356 5756
rect 3298 5168 3356 5180
rect 3426 5756 3484 5768
rect 3426 5180 3438 5756
rect 3472 5180 3484 5756
rect 3426 5168 3484 5180
rect 3538 5756 3596 5768
rect 3538 5180 3550 5756
rect 3584 5180 3596 5756
rect 3538 5168 3596 5180
rect 3666 5756 3724 5768
rect 3666 5180 3678 5756
rect 3712 5180 3724 5756
rect 3666 5168 3724 5180
rect 3778 5756 3836 5768
rect 3778 5180 3790 5756
rect 3824 5180 3836 5756
rect 3778 5168 3836 5180
rect 3906 5756 3964 5768
rect 3906 5180 3918 5756
rect 3952 5180 3964 5756
rect 3906 5168 3964 5180
rect 4018 5756 4076 5768
rect 4018 5180 4030 5756
rect 4064 5180 4076 5756
rect 4018 5168 4076 5180
rect 4146 5756 4204 5768
rect 4146 5180 4158 5756
rect 4192 5180 4204 5756
rect 4146 5168 4204 5180
rect 4258 5756 4316 5768
rect 4258 5180 4270 5756
rect 4304 5180 4316 5756
rect 4258 5168 4316 5180
rect 4386 5756 4444 5768
rect 4386 5180 4398 5756
rect 4432 5180 4444 5756
rect 4386 5168 4444 5180
rect 4498 5756 4556 5768
rect 4498 5180 4510 5756
rect 4544 5180 4556 5756
rect 4498 5168 4556 5180
rect 4626 5756 4684 5768
rect 4626 5180 4638 5756
rect 4672 5180 4684 5756
rect 4626 5168 4684 5180
rect 4738 5756 4796 5768
rect 4738 5180 4750 5756
rect 4784 5180 4796 5756
rect 4738 5168 4796 5180
rect 4866 5756 4924 5768
rect 4866 5180 4878 5756
rect 4912 5180 4924 5756
rect 4866 5168 4924 5180
rect 4978 5756 5036 5768
rect 4978 5180 4990 5756
rect 5024 5180 5036 5756
rect 4978 5168 5036 5180
rect 5106 5756 5164 5768
rect 5106 5180 5118 5756
rect 5152 5180 5164 5756
rect 5106 5168 5164 5180
rect 5218 5756 5276 5768
rect 5218 5180 5230 5756
rect 5264 5180 5276 5756
rect 5218 5168 5276 5180
rect 5346 5756 5404 5768
rect 5346 5180 5358 5756
rect 5392 5180 5404 5756
rect 5346 5168 5404 5180
rect 5458 5756 5516 5768
rect 5458 5180 5470 5756
rect 5504 5180 5516 5756
rect 5458 5168 5516 5180
rect 5586 5756 5644 5768
rect 5586 5180 5598 5756
rect 5632 5180 5644 5756
rect 5586 5168 5644 5180
rect 5698 5756 5756 5768
rect 5698 5180 5710 5756
rect 5744 5180 5756 5756
rect 5698 5168 5756 5180
rect 5826 5756 5884 5768
rect 5826 5180 5838 5756
rect 5872 5180 5884 5756
rect 5826 5168 5884 5180
rect 5938 5756 5996 5768
rect 5938 5180 5950 5756
rect 5984 5180 5996 5756
rect 5938 5168 5996 5180
rect 6066 5756 6124 5768
rect 6066 5180 6078 5756
rect 6112 5180 6124 5756
rect 6066 5168 6124 5180
rect 6178 5756 6236 5768
rect 6178 5180 6190 5756
rect 6224 5180 6236 5756
rect 6178 5168 6236 5180
rect 6306 5756 6364 5768
rect 6306 5180 6318 5756
rect 6352 5180 6364 5756
rect 6306 5168 6364 5180
rect 6418 5756 6476 5768
rect 6418 5180 6430 5756
rect 6464 5180 6476 5756
rect 6418 5168 6476 5180
rect 6546 5756 6604 5768
rect 6546 5180 6558 5756
rect 6592 5180 6604 5756
rect 6546 5168 6604 5180
rect 6658 5756 6716 5768
rect 6658 5180 6670 5756
rect 6704 5180 6716 5756
rect 6658 5168 6716 5180
rect 6786 5756 6844 5768
rect 6786 5180 6798 5756
rect 6832 5180 6844 5756
rect 6786 5168 6844 5180
rect 6898 5756 6956 5768
rect 6898 5180 6910 5756
rect 6944 5180 6956 5756
rect 6898 5168 6956 5180
rect 7026 5756 7084 5768
rect 7026 5180 7038 5756
rect 7072 5180 7084 5756
rect 7026 5168 7084 5180
rect 7138 5756 7196 5768
rect 7138 5180 7150 5756
rect 7184 5180 7196 5756
rect 7138 5168 7196 5180
rect 7266 5756 7324 5768
rect 7266 5180 7278 5756
rect 7312 5180 7324 5756
rect 7266 5168 7324 5180
rect 7378 5756 7436 5768
rect 7378 5180 7390 5756
rect 7424 5180 7436 5756
rect 7378 5168 7436 5180
rect 7506 5756 7564 5768
rect 7506 5180 7518 5756
rect 7552 5180 7564 5756
rect 7506 5168 7564 5180
rect 7618 5756 7676 5768
rect 7618 5180 7630 5756
rect 7664 5180 7676 5756
rect 7618 5168 7676 5180
rect 7746 5756 7804 5768
rect 7746 5180 7758 5756
rect 7792 5180 7804 5756
rect 7746 5168 7804 5180
rect 7858 5756 7916 5768
rect 7858 5180 7870 5756
rect 7904 5180 7916 5756
rect 7858 5168 7916 5180
rect 7986 5756 8044 5768
rect 7986 5180 7998 5756
rect 8032 5180 8044 5756
rect 7986 5168 8044 5180
rect 8098 5756 8156 5768
rect 8098 5180 8110 5756
rect 8144 5180 8156 5756
rect 8098 5168 8156 5180
rect 8226 5756 8284 5768
rect 8226 5180 8238 5756
rect 8272 5180 8284 5756
rect 8226 5168 8284 5180
rect 8338 5756 8396 5768
rect 8338 5180 8350 5756
rect 8384 5180 8396 5756
rect 8338 5168 8396 5180
rect 8466 5756 8524 5768
rect 8466 5180 8478 5756
rect 8512 5180 8524 5756
rect 8466 5168 8524 5180
rect 8578 5756 8636 5768
rect 8578 5180 8590 5756
rect 8624 5180 8636 5756
rect 8578 5168 8636 5180
rect 8706 5756 8764 5768
rect 8706 5180 8718 5756
rect 8752 5180 8764 5756
rect 8706 5168 8764 5180
rect 8818 5756 8876 5768
rect 8818 5180 8830 5756
rect 8864 5180 8876 5756
rect 8818 5168 8876 5180
rect 8946 5756 9004 5768
rect 8946 5180 8958 5756
rect 8992 5180 9004 5756
rect 8946 5168 9004 5180
rect 9058 5756 9116 5768
rect 9058 5180 9070 5756
rect 9104 5180 9116 5756
rect 9058 5168 9116 5180
rect 9186 5756 9244 5768
rect 9186 5180 9198 5756
rect 9232 5180 9244 5756
rect 9186 5168 9244 5180
rect 9298 5756 9356 5768
rect 9298 5180 9310 5756
rect 9344 5180 9356 5756
rect 9298 5168 9356 5180
rect 9426 5756 9484 5768
rect 9426 5180 9438 5756
rect 9472 5180 9484 5756
rect 9426 5168 9484 5180
rect 9538 5756 9596 5768
rect 9538 5180 9550 5756
rect 9584 5180 9596 5756
rect 9538 5168 9596 5180
rect 9666 5756 9724 5768
rect 9666 5180 9678 5756
rect 9712 5180 9724 5756
rect 9666 5168 9724 5180
rect 9778 5756 9836 5768
rect 9778 5180 9790 5756
rect 9824 5180 9836 5756
rect 9778 5168 9836 5180
rect 9906 5756 9964 5768
rect 9906 5180 9918 5756
rect 9952 5180 9964 5756
rect 9906 5168 9964 5180
rect 10018 5756 10076 5768
rect 10018 5180 10030 5756
rect 10064 5180 10076 5756
rect 10018 5168 10076 5180
rect 10146 5756 10204 5768
rect 10146 5180 10158 5756
rect 10192 5180 10204 5756
rect 10146 5168 10204 5180
rect 10258 5756 10316 5768
rect 10258 5180 10270 5756
rect 10304 5180 10316 5756
rect 10258 5168 10316 5180
rect 10386 5756 10444 5768
rect 10386 5180 10398 5756
rect 10432 5180 10444 5756
rect 10386 5168 10444 5180
rect 10498 5756 10556 5768
rect 10498 5180 10510 5756
rect 10544 5180 10556 5756
rect 10498 5168 10556 5180
rect 10626 5756 10684 5768
rect 10626 5180 10638 5756
rect 10672 5180 10684 5756
rect 10626 5168 10684 5180
rect 10738 5756 10796 5768
rect 10738 5180 10750 5756
rect 10784 5180 10796 5756
rect 10738 5168 10796 5180
rect 10866 5756 10924 5768
rect 10866 5180 10878 5756
rect 10912 5180 10924 5756
rect 10866 5168 10924 5180
rect 10978 5756 11036 5768
rect 10978 5180 10990 5756
rect 11024 5180 11036 5756
rect 10978 5168 11036 5180
rect 11106 5756 11164 5768
rect 11106 5180 11118 5756
rect 11152 5180 11164 5756
rect 11106 5168 11164 5180
rect 11218 5756 11276 5768
rect 11218 5180 11230 5756
rect 11264 5180 11276 5756
rect 11218 5168 11276 5180
rect 11346 5756 11404 5768
rect 11346 5180 11358 5756
rect 11392 5180 11404 5756
rect 11346 5168 11404 5180
rect 11458 5756 11516 5768
rect 11458 5180 11470 5756
rect 11504 5180 11516 5756
rect 11458 5168 11516 5180
rect 11586 5756 11644 5768
rect 11586 5180 11598 5756
rect 11632 5180 11644 5756
rect 11586 5168 11644 5180
rect 11698 5756 11756 5768
rect 11698 5180 11710 5756
rect 11744 5180 11756 5756
rect 11698 5168 11756 5180
rect 11826 5756 11884 5768
rect 11826 5180 11838 5756
rect 11872 5180 11884 5756
rect 11826 5168 11884 5180
rect 11938 5756 11996 5768
rect 11938 5180 11950 5756
rect 11984 5180 11996 5756
rect 11938 5168 11996 5180
rect 12066 5756 12124 5768
rect 12066 5180 12078 5756
rect 12112 5180 12124 5756
rect 12066 5168 12124 5180
rect 12178 5756 12236 5768
rect 12178 5180 12190 5756
rect 12224 5180 12236 5756
rect 12178 5168 12236 5180
rect 12306 5756 12364 5768
rect 12306 5180 12318 5756
rect 12352 5180 12364 5756
rect 12306 5168 12364 5180
rect 7138 -6194 7196 -6182
rect 7138 -6770 7150 -6194
rect 7184 -6770 7196 -6194
rect 7138 -6782 7196 -6770
rect 7266 -6194 7324 -6182
rect 7266 -6770 7278 -6194
rect 7312 -6770 7324 -6194
rect 7266 -6782 7324 -6770
rect 7378 -6194 7436 -6182
rect 7378 -6770 7390 -6194
rect 7424 -6770 7436 -6194
rect 7378 -6782 7436 -6770
rect 7506 -6194 7564 -6182
rect 7506 -6770 7518 -6194
rect 7552 -6770 7564 -6194
rect 7506 -6782 7564 -6770
rect 7618 -6194 7676 -6182
rect 7618 -6770 7630 -6194
rect 7664 -6770 7676 -6194
rect 7618 -6782 7676 -6770
rect 7746 -6194 7804 -6182
rect 7746 -6770 7758 -6194
rect 7792 -6770 7804 -6194
rect 7746 -6782 7804 -6770
rect 7858 -6194 7916 -6182
rect 7858 -6770 7870 -6194
rect 7904 -6770 7916 -6194
rect 7858 -6782 7916 -6770
rect 7986 -6194 8044 -6182
rect 7986 -6770 7998 -6194
rect 8032 -6770 8044 -6194
rect 7986 -6782 8044 -6770
rect 7138 -7002 7196 -6990
rect 7138 -7578 7150 -7002
rect 7184 -7578 7196 -7002
rect 7138 -7590 7196 -7578
rect 7266 -7002 7324 -6990
rect 7266 -7578 7278 -7002
rect 7312 -7578 7324 -7002
rect 7266 -7590 7324 -7578
rect 7378 -7002 7436 -6990
rect 7378 -7578 7390 -7002
rect 7424 -7578 7436 -7002
rect 7378 -7590 7436 -7578
rect 7506 -7002 7564 -6990
rect 7506 -7578 7518 -7002
rect 7552 -7578 7564 -7002
rect 7506 -7590 7564 -7578
rect 7618 -7002 7676 -6990
rect 7618 -7578 7630 -7002
rect 7664 -7578 7676 -7002
rect 7618 -7590 7676 -7578
rect 7746 -7002 7804 -6990
rect 7746 -7578 7758 -7002
rect 7792 -7578 7804 -7002
rect 7746 -7590 7804 -7578
rect 7858 -7002 7916 -6990
rect 7858 -7578 7870 -7002
rect 7904 -7578 7916 -7002
rect 7858 -7590 7916 -7578
rect 7986 -7002 8044 -6990
rect 7986 -7578 7998 -7002
rect 8032 -7578 8044 -7002
rect 7986 -7590 8044 -7578
<< pdiff >>
rect -6486 2444 -6428 2456
rect -6486 1668 -6474 2444
rect -6440 1668 -6428 2444
rect -6486 1656 -6428 1668
rect -6028 2444 -5970 2456
rect -6028 1668 -6016 2444
rect -5982 1668 -5970 2444
rect -6028 1656 -5970 1668
rect -5898 2444 -5840 2456
rect -5898 1668 -5886 2444
rect -5852 1668 -5840 2444
rect -5898 1656 -5840 1668
rect -5440 2444 -5382 2456
rect -5440 1668 -5428 2444
rect -5394 1668 -5382 2444
rect -5440 1656 -5382 1668
rect -5310 2444 -5252 2456
rect -5310 1668 -5298 2444
rect -5264 1668 -5252 2444
rect -5310 1656 -5252 1668
rect -4852 2444 -4794 2456
rect -4852 1668 -4840 2444
rect -4806 1668 -4794 2444
rect -4852 1656 -4794 1668
rect -4722 2444 -4664 2456
rect -4722 1668 -4710 2444
rect -4676 1668 -4664 2444
rect -4722 1656 -4664 1668
rect -4264 2444 -4206 2456
rect -4264 1668 -4252 2444
rect -4218 1668 -4206 2444
rect -4264 1656 -4206 1668
rect -4134 2444 -4076 2456
rect -4134 1668 -4122 2444
rect -4088 1668 -4076 2444
rect -4134 1656 -4076 1668
rect -3676 2444 -3618 2456
rect -3676 1668 -3664 2444
rect -3630 1668 -3618 2444
rect -3676 1656 -3618 1668
rect -3546 2444 -3488 2456
rect -3546 1668 -3534 2444
rect -3500 1668 -3488 2444
rect -3546 1656 -3488 1668
rect -3088 2444 -3030 2456
rect -3088 1668 -3076 2444
rect -3042 1668 -3030 2444
rect -3088 1656 -3030 1668
rect -2958 2444 -2900 2456
rect -2958 1668 -2946 2444
rect -2912 1668 -2900 2444
rect -2958 1656 -2900 1668
rect -2500 2444 -2442 2456
rect -2500 1668 -2488 2444
rect -2454 1668 -2442 2444
rect -2500 1656 -2442 1668
rect -2370 2444 -2312 2456
rect -2370 1668 -2358 2444
rect -2324 1668 -2312 2444
rect -2370 1656 -2312 1668
rect -1912 2444 -1854 2456
rect -1912 1668 -1900 2444
rect -1866 1668 -1854 2444
rect -1912 1656 -1854 1668
rect -1782 2444 -1724 2456
rect -1782 1668 -1770 2444
rect -1736 1668 -1724 2444
rect -1782 1656 -1724 1668
rect -1324 2444 -1266 2456
rect -1324 1668 -1312 2444
rect -1278 1668 -1266 2444
rect -1324 1656 -1266 1668
rect -1194 2444 -1136 2456
rect -1194 1668 -1182 2444
rect -1148 1668 -1136 2444
rect -1194 1656 -1136 1668
rect -736 2444 -678 2456
rect -736 1668 -724 2444
rect -690 1668 -678 2444
rect -736 1656 -678 1668
rect -606 2444 -548 2456
rect -606 1668 -594 2444
rect -560 1668 -548 2444
rect -606 1656 -548 1668
rect -148 2444 -90 2456
rect -148 1668 -136 2444
rect -102 1668 -90 2444
rect -148 1656 -90 1668
rect -18 2444 40 2456
rect -18 1668 -6 2444
rect 28 1668 40 2444
rect -18 1656 40 1668
rect 440 2444 498 2456
rect 440 1668 452 2444
rect 486 1668 498 2444
rect 440 1656 498 1668
rect 570 2444 628 2456
rect 570 1668 582 2444
rect 616 1668 628 2444
rect 570 1656 628 1668
rect 1028 2444 1086 2456
rect 1028 1668 1040 2444
rect 1074 1668 1086 2444
rect 1028 1656 1086 1668
rect 1158 2444 1216 2456
rect 1158 1668 1170 2444
rect 1204 1668 1216 2444
rect 1158 1656 1216 1668
rect 1616 2444 1674 2456
rect 1616 1668 1628 2444
rect 1662 1668 1674 2444
rect 1616 1656 1674 1668
rect 1746 2444 1804 2456
rect 1746 1668 1758 2444
rect 1792 1668 1804 2444
rect 1746 1656 1804 1668
rect 2204 2444 2262 2456
rect 2204 1668 2216 2444
rect 2250 1668 2262 2444
rect 2204 1656 2262 1668
rect 2334 2444 2392 2456
rect 2334 1668 2346 2444
rect 2380 1668 2392 2444
rect 2334 1656 2392 1668
rect 2792 2444 2850 2456
rect 2792 1668 2804 2444
rect 2838 1668 2850 2444
rect 2792 1656 2850 1668
rect 2922 2444 2980 2456
rect 2922 1668 2934 2444
rect 2968 1668 2980 2444
rect 2922 1656 2980 1668
rect 3380 2444 3438 2456
rect 3380 1668 3392 2444
rect 3426 1668 3438 2444
rect 3380 1656 3438 1668
rect 3510 2444 3568 2456
rect 3510 1668 3522 2444
rect 3556 1668 3568 2444
rect 3510 1656 3568 1668
rect 3968 2444 4026 2456
rect 3968 1668 3980 2444
rect 4014 1668 4026 2444
rect 3968 1656 4026 1668
rect 4098 2444 4156 2456
rect 4098 1668 4110 2444
rect 4144 1668 4156 2444
rect 4098 1656 4156 1668
rect 4556 2444 4614 2456
rect 4556 1668 4568 2444
rect 4602 1668 4614 2444
rect 4556 1656 4614 1668
rect 4686 2444 4744 2456
rect 4686 1668 4698 2444
rect 4732 1668 4744 2444
rect 4686 1656 4744 1668
rect 5144 2444 5202 2456
rect 5144 1668 5156 2444
rect 5190 1668 5202 2444
rect 5144 1656 5202 1668
rect 5274 2444 5332 2456
rect 5274 1668 5286 2444
rect 5320 1668 5332 2444
rect 5274 1656 5332 1668
rect 5732 2444 5790 2456
rect 5732 1668 5744 2444
rect 5778 1668 5790 2444
rect 5732 1656 5790 1668
rect 5862 2444 5920 2456
rect 5862 1668 5874 2444
rect 5908 1668 5920 2444
rect 5862 1656 5920 1668
rect 6320 2444 6378 2456
rect 6320 1668 6332 2444
rect 6366 1668 6378 2444
rect 6320 1656 6378 1668
rect 6450 2444 6508 2456
rect 6450 1668 6462 2444
rect 6496 1668 6508 2444
rect 6450 1656 6508 1668
rect 6908 2444 6966 2456
rect 6908 1668 6920 2444
rect 6954 1668 6966 2444
rect 6908 1656 6966 1668
rect 7038 2444 7096 2456
rect 7038 1668 7050 2444
rect 7084 1668 7096 2444
rect 7038 1656 7096 1668
rect 7496 2444 7554 2456
rect 7496 1668 7508 2444
rect 7542 1668 7554 2444
rect 7496 1656 7554 1668
rect 7626 2444 7684 2456
rect 7626 1668 7638 2444
rect 7672 1668 7684 2444
rect 7626 1656 7684 1668
rect 8084 2444 8142 2456
rect 8084 1668 8096 2444
rect 8130 1668 8142 2444
rect 8084 1656 8142 1668
rect 8214 2444 8272 2456
rect 8214 1668 8226 2444
rect 8260 1668 8272 2444
rect 8214 1656 8272 1668
rect 8672 2444 8730 2456
rect 8672 1668 8684 2444
rect 8718 1668 8730 2444
rect 8672 1656 8730 1668
rect 8802 2444 8860 2456
rect 8802 1668 8814 2444
rect 8848 1668 8860 2444
rect 8802 1656 8860 1668
rect 9260 2444 9318 2456
rect 9260 1668 9272 2444
rect 9306 1668 9318 2444
rect 9260 1656 9318 1668
rect 9390 2444 9448 2456
rect 9390 1668 9402 2444
rect 9436 1668 9448 2444
rect 9390 1656 9448 1668
rect 9848 2444 9906 2456
rect 9848 1668 9860 2444
rect 9894 1668 9906 2444
rect 9848 1656 9906 1668
rect 9978 2444 10036 2456
rect 9978 1668 9990 2444
rect 10024 1668 10036 2444
rect 9978 1656 10036 1668
rect 10436 2444 10494 2456
rect 10436 1668 10448 2444
rect 10482 1668 10494 2444
rect 10436 1656 10494 1668
rect 10566 2444 10624 2456
rect 10566 1668 10578 2444
rect 10612 1668 10624 2444
rect 10566 1656 10624 1668
rect 11024 2444 11082 2456
rect 11024 1668 11036 2444
rect 11070 1668 11082 2444
rect 11024 1656 11082 1668
rect 11154 2444 11212 2456
rect 11154 1668 11166 2444
rect 11200 1668 11212 2444
rect 11154 1656 11212 1668
rect 11612 2444 11670 2456
rect 11612 1668 11624 2444
rect 11658 1668 11670 2444
rect 11612 1656 11670 1668
rect 11742 2444 11800 2456
rect 11742 1668 11754 2444
rect 11788 1668 11800 2444
rect 11742 1656 11800 1668
rect 12200 2444 12258 2456
rect 12200 1668 12212 2444
rect 12246 1668 12258 2444
rect 12200 1656 12258 1668
rect 12330 2444 12388 2456
rect 12330 1668 12342 2444
rect 12376 1668 12388 2444
rect 12330 1656 12388 1668
rect 12788 2444 12846 2456
rect 12788 1668 12800 2444
rect 12834 1668 12846 2444
rect 12788 1656 12846 1668
rect 12918 2444 12976 2456
rect 12918 1668 12930 2444
rect 12964 1668 12976 2444
rect 12918 1656 12976 1668
rect 13376 2444 13434 2456
rect 13376 1668 13388 2444
rect 13422 1668 13434 2444
rect 13376 1656 13434 1668
rect 13506 2444 13564 2456
rect 13506 1668 13518 2444
rect 13552 1668 13564 2444
rect 13506 1656 13564 1668
rect 13964 2444 14022 2456
rect 13964 1668 13976 2444
rect 14010 1668 14022 2444
rect 13964 1656 14022 1668
rect 14094 2444 14152 2456
rect 14094 1668 14106 2444
rect 14140 1668 14152 2444
rect 14094 1656 14152 1668
rect 14552 2444 14610 2456
rect 14552 1668 14564 2444
rect 14598 1668 14610 2444
rect 14552 1656 14610 1668
rect 14682 2444 14740 2456
rect 14682 1668 14694 2444
rect 14728 1668 14740 2444
rect 14682 1656 14740 1668
rect 15140 2444 15198 2456
rect 15140 1668 15152 2444
rect 15186 1668 15198 2444
rect 15140 1656 15198 1668
rect 15270 2444 15328 2456
rect 15270 1668 15282 2444
rect 15316 1668 15328 2444
rect 15270 1656 15328 1668
rect 15728 2444 15786 2456
rect 15728 1668 15740 2444
rect 15774 1668 15786 2444
rect 15728 1656 15786 1668
rect 15858 2444 15916 2456
rect 15858 1668 15870 2444
rect 15904 1668 15916 2444
rect 15858 1656 15916 1668
rect 16316 2444 16374 2456
rect 16316 1668 16328 2444
rect 16362 1668 16374 2444
rect 16316 1656 16374 1668
rect 16446 2444 16504 2456
rect 16446 1668 16458 2444
rect 16492 1668 16504 2444
rect 16446 1656 16504 1668
rect 16904 2444 16962 2456
rect 16904 1668 16916 2444
rect 16950 1668 16962 2444
rect 16904 1656 16962 1668
rect 17034 2444 17092 2456
rect 17034 1668 17046 2444
rect 17080 1668 17092 2444
rect 17034 1656 17092 1668
rect 17492 2444 17550 2456
rect 17492 1668 17504 2444
rect 17538 1668 17550 2444
rect 17492 1656 17550 1668
rect 17622 2444 17680 2456
rect 17622 1668 17634 2444
rect 17668 1668 17680 2444
rect 17622 1656 17680 1668
rect 18080 2444 18138 2456
rect 18080 1668 18092 2444
rect 18126 1668 18138 2444
rect 18080 1656 18138 1668
rect 18210 2444 18268 2456
rect 18210 1668 18222 2444
rect 18256 1668 18268 2444
rect 18210 1656 18268 1668
rect 18668 2444 18726 2456
rect 18668 1668 18680 2444
rect 18714 1668 18726 2444
rect 18668 1656 18726 1668
rect 18798 2444 18856 2456
rect 18798 1668 18810 2444
rect 18844 1668 18856 2444
rect 18798 1656 18856 1668
rect 19256 2444 19314 2456
rect 19256 1668 19268 2444
rect 19302 1668 19314 2444
rect 19256 1656 19314 1668
rect 19386 2444 19444 2456
rect 19386 1668 19398 2444
rect 19432 1668 19444 2444
rect 19386 1656 19444 1668
rect 19844 2444 19902 2456
rect 19844 1668 19856 2444
rect 19890 1668 19902 2444
rect 19844 1656 19902 1668
rect 19974 2444 20032 2456
rect 19974 1668 19986 2444
rect 20020 1668 20032 2444
rect 19974 1656 20032 1668
rect 20432 2444 20490 2456
rect 20432 1668 20444 2444
rect 20478 1668 20490 2444
rect 20432 1656 20490 1668
rect 20562 2444 20620 2456
rect 20562 1668 20574 2444
rect 20608 1668 20620 2444
rect 20562 1656 20620 1668
rect 21020 2444 21078 2456
rect 21020 1668 21032 2444
rect 21066 1668 21078 2444
rect 21020 1656 21078 1668
rect 21150 2444 21208 2456
rect 21150 1668 21162 2444
rect 21196 1668 21208 2444
rect 21150 1656 21208 1668
rect 21608 2444 21666 2456
rect 21608 1668 21620 2444
rect 21654 1668 21666 2444
rect 21608 1656 21666 1668
rect -6486 1444 -6428 1456
rect -6486 668 -6474 1444
rect -6440 668 -6428 1444
rect -6486 656 -6428 668
rect -6028 1444 -5970 1456
rect -6028 668 -6016 1444
rect -5982 668 -5970 1444
rect -6028 656 -5970 668
rect -5898 1444 -5840 1456
rect -5898 668 -5886 1444
rect -5852 668 -5840 1444
rect -5898 656 -5840 668
rect -5440 1444 -5382 1456
rect -5440 668 -5428 1444
rect -5394 668 -5382 1444
rect -5440 656 -5382 668
rect -5310 1444 -5252 1456
rect -5310 668 -5298 1444
rect -5264 668 -5252 1444
rect -5310 656 -5252 668
rect -4852 1444 -4794 1456
rect -4852 668 -4840 1444
rect -4806 668 -4794 1444
rect -4852 656 -4794 668
rect -4722 1444 -4664 1456
rect -4722 668 -4710 1444
rect -4676 668 -4664 1444
rect -4722 656 -4664 668
rect -4264 1444 -4206 1456
rect -4264 668 -4252 1444
rect -4218 668 -4206 1444
rect -4264 656 -4206 668
rect -4134 1444 -4076 1456
rect -4134 668 -4122 1444
rect -4088 668 -4076 1444
rect -4134 656 -4076 668
rect -3676 1444 -3618 1456
rect -3676 668 -3664 1444
rect -3630 668 -3618 1444
rect -3676 656 -3618 668
rect -3546 1444 -3488 1456
rect -3546 668 -3534 1444
rect -3500 668 -3488 1444
rect -3546 656 -3488 668
rect -3088 1444 -3030 1456
rect -3088 668 -3076 1444
rect -3042 668 -3030 1444
rect -3088 656 -3030 668
rect -2958 1444 -2900 1456
rect -2958 668 -2946 1444
rect -2912 668 -2900 1444
rect -2958 656 -2900 668
rect -2500 1444 -2442 1456
rect -2500 668 -2488 1444
rect -2454 668 -2442 1444
rect -2500 656 -2442 668
rect -2370 1444 -2312 1456
rect -2370 668 -2358 1444
rect -2324 668 -2312 1444
rect -2370 656 -2312 668
rect -1912 1444 -1854 1456
rect -1912 668 -1900 1444
rect -1866 668 -1854 1444
rect -1912 656 -1854 668
rect -1782 1444 -1724 1456
rect -1782 668 -1770 1444
rect -1736 668 -1724 1444
rect -1782 656 -1724 668
rect -1324 1444 -1266 1456
rect -1324 668 -1312 1444
rect -1278 668 -1266 1444
rect -1324 656 -1266 668
rect -1194 1444 -1136 1456
rect -1194 668 -1182 1444
rect -1148 668 -1136 1444
rect -1194 656 -1136 668
rect -736 1444 -678 1456
rect -736 668 -724 1444
rect -690 668 -678 1444
rect -736 656 -678 668
rect -606 1444 -548 1456
rect -606 668 -594 1444
rect -560 668 -548 1444
rect -606 656 -548 668
rect -148 1444 -90 1456
rect -148 668 -136 1444
rect -102 668 -90 1444
rect -148 656 -90 668
rect -18 1444 40 1456
rect -18 668 -6 1444
rect 28 668 40 1444
rect -18 656 40 668
rect 440 1444 498 1456
rect 440 668 452 1444
rect 486 668 498 1444
rect 440 656 498 668
rect 570 1444 628 1456
rect 570 668 582 1444
rect 616 668 628 1444
rect 570 656 628 668
rect 1028 1444 1086 1456
rect 1028 668 1040 1444
rect 1074 668 1086 1444
rect 1028 656 1086 668
rect 1158 1444 1216 1456
rect 1158 668 1170 1444
rect 1204 668 1216 1444
rect 1158 656 1216 668
rect 1616 1444 1674 1456
rect 1616 668 1628 1444
rect 1662 668 1674 1444
rect 1616 656 1674 668
rect 1746 1444 1804 1456
rect 1746 668 1758 1444
rect 1792 668 1804 1444
rect 1746 656 1804 668
rect 2204 1444 2262 1456
rect 2204 668 2216 1444
rect 2250 668 2262 1444
rect 2204 656 2262 668
rect 2334 1444 2392 1456
rect 2334 668 2346 1444
rect 2380 668 2392 1444
rect 2334 656 2392 668
rect 2792 1444 2850 1456
rect 2792 668 2804 1444
rect 2838 668 2850 1444
rect 2792 656 2850 668
rect 2922 1444 2980 1456
rect 2922 668 2934 1444
rect 2968 668 2980 1444
rect 2922 656 2980 668
rect 3380 1444 3438 1456
rect 3380 668 3392 1444
rect 3426 668 3438 1444
rect 3380 656 3438 668
rect 3510 1444 3568 1456
rect 3510 668 3522 1444
rect 3556 668 3568 1444
rect 3510 656 3568 668
rect 3968 1444 4026 1456
rect 3968 668 3980 1444
rect 4014 668 4026 1444
rect 3968 656 4026 668
rect 4098 1444 4156 1456
rect 4098 668 4110 1444
rect 4144 668 4156 1444
rect 4098 656 4156 668
rect 4556 1444 4614 1456
rect 4556 668 4568 1444
rect 4602 668 4614 1444
rect 4556 656 4614 668
rect 4686 1444 4744 1456
rect 4686 668 4698 1444
rect 4732 668 4744 1444
rect 4686 656 4744 668
rect 5144 1444 5202 1456
rect 5144 668 5156 1444
rect 5190 668 5202 1444
rect 5144 656 5202 668
rect 5274 1444 5332 1456
rect 5274 668 5286 1444
rect 5320 668 5332 1444
rect 5274 656 5332 668
rect 5732 1444 5790 1456
rect 5732 668 5744 1444
rect 5778 668 5790 1444
rect 5732 656 5790 668
rect 5862 1444 5920 1456
rect 5862 668 5874 1444
rect 5908 668 5920 1444
rect 5862 656 5920 668
rect 6320 1444 6378 1456
rect 6320 668 6332 1444
rect 6366 668 6378 1444
rect 6320 656 6378 668
rect 6450 1444 6508 1456
rect 6450 668 6462 1444
rect 6496 668 6508 1444
rect 6450 656 6508 668
rect 6908 1444 6966 1456
rect 6908 668 6920 1444
rect 6954 668 6966 1444
rect 6908 656 6966 668
rect 7038 1444 7096 1456
rect 7038 668 7050 1444
rect 7084 668 7096 1444
rect 7038 656 7096 668
rect 7496 1444 7554 1456
rect 7496 668 7508 1444
rect 7542 668 7554 1444
rect 7496 656 7554 668
rect 7626 1444 7684 1456
rect 7626 668 7638 1444
rect 7672 668 7684 1444
rect 7626 656 7684 668
rect 8084 1444 8142 1456
rect 8084 668 8096 1444
rect 8130 668 8142 1444
rect 8084 656 8142 668
rect 8214 1444 8272 1456
rect 8214 668 8226 1444
rect 8260 668 8272 1444
rect 8214 656 8272 668
rect 8672 1444 8730 1456
rect 8672 668 8684 1444
rect 8718 668 8730 1444
rect 8672 656 8730 668
rect 8802 1444 8860 1456
rect 8802 668 8814 1444
rect 8848 668 8860 1444
rect 8802 656 8860 668
rect 9260 1444 9318 1456
rect 9260 668 9272 1444
rect 9306 668 9318 1444
rect 9260 656 9318 668
rect 9390 1444 9448 1456
rect 9390 668 9402 1444
rect 9436 668 9448 1444
rect 9390 656 9448 668
rect 9848 1444 9906 1456
rect 9848 668 9860 1444
rect 9894 668 9906 1444
rect 9848 656 9906 668
rect 9978 1444 10036 1456
rect 9978 668 9990 1444
rect 10024 668 10036 1444
rect 9978 656 10036 668
rect 10436 1444 10494 1456
rect 10436 668 10448 1444
rect 10482 668 10494 1444
rect 10436 656 10494 668
rect 10566 1444 10624 1456
rect 10566 668 10578 1444
rect 10612 668 10624 1444
rect 10566 656 10624 668
rect 11024 1444 11082 1456
rect 11024 668 11036 1444
rect 11070 668 11082 1444
rect 11024 656 11082 668
rect 11154 1444 11212 1456
rect 11154 668 11166 1444
rect 11200 668 11212 1444
rect 11154 656 11212 668
rect 11612 1444 11670 1456
rect 11612 668 11624 1444
rect 11658 668 11670 1444
rect 11612 656 11670 668
rect 11742 1444 11800 1456
rect 11742 668 11754 1444
rect 11788 668 11800 1444
rect 11742 656 11800 668
rect 12200 1444 12258 1456
rect 12200 668 12212 1444
rect 12246 668 12258 1444
rect 12200 656 12258 668
rect 12330 1444 12388 1456
rect 12330 668 12342 1444
rect 12376 668 12388 1444
rect 12330 656 12388 668
rect 12788 1444 12846 1456
rect 12788 668 12800 1444
rect 12834 668 12846 1444
rect 12788 656 12846 668
rect 12918 1444 12976 1456
rect 12918 668 12930 1444
rect 12964 668 12976 1444
rect 12918 656 12976 668
rect 13376 1444 13434 1456
rect 13376 668 13388 1444
rect 13422 668 13434 1444
rect 13376 656 13434 668
rect 13506 1444 13564 1456
rect 13506 668 13518 1444
rect 13552 668 13564 1444
rect 13506 656 13564 668
rect 13964 1444 14022 1456
rect 13964 668 13976 1444
rect 14010 668 14022 1444
rect 13964 656 14022 668
rect 14094 1444 14152 1456
rect 14094 668 14106 1444
rect 14140 668 14152 1444
rect 14094 656 14152 668
rect 14552 1444 14610 1456
rect 14552 668 14564 1444
rect 14598 668 14610 1444
rect 14552 656 14610 668
rect 14682 1444 14740 1456
rect 14682 668 14694 1444
rect 14728 668 14740 1444
rect 14682 656 14740 668
rect 15140 1444 15198 1456
rect 15140 668 15152 1444
rect 15186 668 15198 1444
rect 15140 656 15198 668
rect 15270 1444 15328 1456
rect 15270 668 15282 1444
rect 15316 668 15328 1444
rect 15270 656 15328 668
rect 15728 1444 15786 1456
rect 15728 668 15740 1444
rect 15774 668 15786 1444
rect 15728 656 15786 668
rect 15858 1444 15916 1456
rect 15858 668 15870 1444
rect 15904 668 15916 1444
rect 15858 656 15916 668
rect 16316 1444 16374 1456
rect 16316 668 16328 1444
rect 16362 668 16374 1444
rect 16316 656 16374 668
rect 16446 1444 16504 1456
rect 16446 668 16458 1444
rect 16492 668 16504 1444
rect 16446 656 16504 668
rect 16904 1444 16962 1456
rect 16904 668 16916 1444
rect 16950 668 16962 1444
rect 16904 656 16962 668
rect 17034 1444 17092 1456
rect 17034 668 17046 1444
rect 17080 668 17092 1444
rect 17034 656 17092 668
rect 17492 1444 17550 1456
rect 17492 668 17504 1444
rect 17538 668 17550 1444
rect 17492 656 17550 668
rect 17622 1444 17680 1456
rect 17622 668 17634 1444
rect 17668 668 17680 1444
rect 17622 656 17680 668
rect 18080 1444 18138 1456
rect 18080 668 18092 1444
rect 18126 668 18138 1444
rect 18080 656 18138 668
rect 18210 1444 18268 1456
rect 18210 668 18222 1444
rect 18256 668 18268 1444
rect 18210 656 18268 668
rect 18668 1444 18726 1456
rect 18668 668 18680 1444
rect 18714 668 18726 1444
rect 18668 656 18726 668
rect 18798 1444 18856 1456
rect 18798 668 18810 1444
rect 18844 668 18856 1444
rect 18798 656 18856 668
rect 19256 1444 19314 1456
rect 19256 668 19268 1444
rect 19302 668 19314 1444
rect 19256 656 19314 668
rect 19386 1444 19444 1456
rect 19386 668 19398 1444
rect 19432 668 19444 1444
rect 19386 656 19444 668
rect 19844 1444 19902 1456
rect 19844 668 19856 1444
rect 19890 668 19902 1444
rect 19844 656 19902 668
rect 19974 1444 20032 1456
rect 19974 668 19986 1444
rect 20020 668 20032 1444
rect 19974 656 20032 668
rect 20432 1444 20490 1456
rect 20432 668 20444 1444
rect 20478 668 20490 1444
rect 20432 656 20490 668
rect 20562 1444 20620 1456
rect 20562 668 20574 1444
rect 20608 668 20620 1444
rect 20562 656 20620 668
rect 21020 1444 21078 1456
rect 21020 668 21032 1444
rect 21066 668 21078 1444
rect 21020 656 21078 668
rect 21150 1444 21208 1456
rect 21150 668 21162 1444
rect 21196 668 21208 1444
rect 21150 656 21208 668
rect 21608 1444 21666 1456
rect 21608 668 21620 1444
rect 21654 668 21666 1444
rect 21608 656 21666 668
rect -6486 444 -6428 456
rect -6486 -332 -6474 444
rect -6440 -332 -6428 444
rect -6486 -344 -6428 -332
rect -6028 444 -5970 456
rect -6028 -332 -6016 444
rect -5982 -332 -5970 444
rect -6028 -344 -5970 -332
rect -5898 444 -5840 456
rect -5898 -332 -5886 444
rect -5852 -332 -5840 444
rect -5898 -344 -5840 -332
rect -5440 444 -5382 456
rect -5440 -332 -5428 444
rect -5394 -332 -5382 444
rect -5440 -344 -5382 -332
rect -5310 444 -5252 456
rect -5310 -332 -5298 444
rect -5264 -332 -5252 444
rect -5310 -344 -5252 -332
rect -4852 444 -4794 456
rect -4852 -332 -4840 444
rect -4806 -332 -4794 444
rect -4852 -344 -4794 -332
rect -4722 444 -4664 456
rect -4722 -332 -4710 444
rect -4676 -332 -4664 444
rect -4722 -344 -4664 -332
rect -4264 444 -4206 456
rect -4264 -332 -4252 444
rect -4218 -332 -4206 444
rect -4264 -344 -4206 -332
rect -4134 444 -4076 456
rect -4134 -332 -4122 444
rect -4088 -332 -4076 444
rect -4134 -344 -4076 -332
rect -3676 444 -3618 456
rect -3676 -332 -3664 444
rect -3630 -332 -3618 444
rect -3676 -344 -3618 -332
rect -3546 444 -3488 456
rect -3546 -332 -3534 444
rect -3500 -332 -3488 444
rect -3546 -344 -3488 -332
rect -3088 444 -3030 456
rect -3088 -332 -3076 444
rect -3042 -332 -3030 444
rect -3088 -344 -3030 -332
rect -2958 444 -2900 456
rect -2958 -332 -2946 444
rect -2912 -332 -2900 444
rect -2958 -344 -2900 -332
rect -2500 444 -2442 456
rect -2500 -332 -2488 444
rect -2454 -332 -2442 444
rect -2500 -344 -2442 -332
rect -2370 444 -2312 456
rect -2370 -332 -2358 444
rect -2324 -332 -2312 444
rect -2370 -344 -2312 -332
rect -1912 444 -1854 456
rect -1912 -332 -1900 444
rect -1866 -332 -1854 444
rect -1912 -344 -1854 -332
rect -1782 444 -1724 456
rect -1782 -332 -1770 444
rect -1736 -332 -1724 444
rect -1782 -344 -1724 -332
rect -1324 444 -1266 456
rect -1324 -332 -1312 444
rect -1278 -332 -1266 444
rect -1324 -344 -1266 -332
rect -1194 444 -1136 456
rect -1194 -332 -1182 444
rect -1148 -332 -1136 444
rect -1194 -344 -1136 -332
rect -736 444 -678 456
rect -736 -332 -724 444
rect -690 -332 -678 444
rect -736 -344 -678 -332
rect -606 444 -548 456
rect -606 -332 -594 444
rect -560 -332 -548 444
rect -606 -344 -548 -332
rect -148 444 -90 456
rect -148 -332 -136 444
rect -102 -332 -90 444
rect -148 -344 -90 -332
rect -18 444 40 456
rect -18 -332 -6 444
rect 28 -332 40 444
rect -18 -344 40 -332
rect 440 444 498 456
rect 440 -332 452 444
rect 486 -332 498 444
rect 440 -344 498 -332
rect 570 444 628 456
rect 570 -332 582 444
rect 616 -332 628 444
rect 570 -344 628 -332
rect 1028 444 1086 456
rect 1028 -332 1040 444
rect 1074 -332 1086 444
rect 1028 -344 1086 -332
rect 1158 444 1216 456
rect 1158 -332 1170 444
rect 1204 -332 1216 444
rect 1158 -344 1216 -332
rect 1616 444 1674 456
rect 1616 -332 1628 444
rect 1662 -332 1674 444
rect 1616 -344 1674 -332
rect 1746 444 1804 456
rect 1746 -332 1758 444
rect 1792 -332 1804 444
rect 1746 -344 1804 -332
rect 2204 444 2262 456
rect 2204 -332 2216 444
rect 2250 -332 2262 444
rect 2204 -344 2262 -332
rect 2334 444 2392 456
rect 2334 -332 2346 444
rect 2380 -332 2392 444
rect 2334 -344 2392 -332
rect 2792 444 2850 456
rect 2792 -332 2804 444
rect 2838 -332 2850 444
rect 2792 -344 2850 -332
rect 2922 444 2980 456
rect 2922 -332 2934 444
rect 2968 -332 2980 444
rect 2922 -344 2980 -332
rect 3380 444 3438 456
rect 3380 -332 3392 444
rect 3426 -332 3438 444
rect 3380 -344 3438 -332
rect 3510 444 3568 456
rect 3510 -332 3522 444
rect 3556 -332 3568 444
rect 3510 -344 3568 -332
rect 3968 444 4026 456
rect 3968 -332 3980 444
rect 4014 -332 4026 444
rect 3968 -344 4026 -332
rect 4098 444 4156 456
rect 4098 -332 4110 444
rect 4144 -332 4156 444
rect 4098 -344 4156 -332
rect 4556 444 4614 456
rect 4556 -332 4568 444
rect 4602 -332 4614 444
rect 4556 -344 4614 -332
rect 4686 444 4744 456
rect 4686 -332 4698 444
rect 4732 -332 4744 444
rect 4686 -344 4744 -332
rect 5144 444 5202 456
rect 5144 -332 5156 444
rect 5190 -332 5202 444
rect 5144 -344 5202 -332
rect 5274 444 5332 456
rect 5274 -332 5286 444
rect 5320 -332 5332 444
rect 5274 -344 5332 -332
rect 5732 444 5790 456
rect 5732 -332 5744 444
rect 5778 -332 5790 444
rect 5732 -344 5790 -332
rect 5862 444 5920 456
rect 5862 -332 5874 444
rect 5908 -332 5920 444
rect 5862 -344 5920 -332
rect 6320 444 6378 456
rect 6320 -332 6332 444
rect 6366 -332 6378 444
rect 6320 -344 6378 -332
rect 6450 444 6508 456
rect 6450 -332 6462 444
rect 6496 -332 6508 444
rect 6450 -344 6508 -332
rect 6908 444 6966 456
rect 6908 -332 6920 444
rect 6954 -332 6966 444
rect 6908 -344 6966 -332
rect 7038 444 7096 456
rect 7038 -332 7050 444
rect 7084 -332 7096 444
rect 7038 -344 7096 -332
rect 7496 444 7554 456
rect 7496 -332 7508 444
rect 7542 -332 7554 444
rect 7496 -344 7554 -332
rect 7626 444 7684 456
rect 7626 -332 7638 444
rect 7672 -332 7684 444
rect 7626 -344 7684 -332
rect 8084 444 8142 456
rect 8084 -332 8096 444
rect 8130 -332 8142 444
rect 8084 -344 8142 -332
rect 8214 444 8272 456
rect 8214 -332 8226 444
rect 8260 -332 8272 444
rect 8214 -344 8272 -332
rect 8672 444 8730 456
rect 8672 -332 8684 444
rect 8718 -332 8730 444
rect 8672 -344 8730 -332
rect 8802 444 8860 456
rect 8802 -332 8814 444
rect 8848 -332 8860 444
rect 8802 -344 8860 -332
rect 9260 444 9318 456
rect 9260 -332 9272 444
rect 9306 -332 9318 444
rect 9260 -344 9318 -332
rect 9390 444 9448 456
rect 9390 -332 9402 444
rect 9436 -332 9448 444
rect 9390 -344 9448 -332
rect 9848 444 9906 456
rect 9848 -332 9860 444
rect 9894 -332 9906 444
rect 9848 -344 9906 -332
rect 9978 444 10036 456
rect 9978 -332 9990 444
rect 10024 -332 10036 444
rect 9978 -344 10036 -332
rect 10436 444 10494 456
rect 10436 -332 10448 444
rect 10482 -332 10494 444
rect 10436 -344 10494 -332
rect 10566 444 10624 456
rect 10566 -332 10578 444
rect 10612 -332 10624 444
rect 10566 -344 10624 -332
rect 11024 444 11082 456
rect 11024 -332 11036 444
rect 11070 -332 11082 444
rect 11024 -344 11082 -332
rect 11154 444 11212 456
rect 11154 -332 11166 444
rect 11200 -332 11212 444
rect 11154 -344 11212 -332
rect 11612 444 11670 456
rect 11612 -332 11624 444
rect 11658 -332 11670 444
rect 11612 -344 11670 -332
rect 11742 444 11800 456
rect 11742 -332 11754 444
rect 11788 -332 11800 444
rect 11742 -344 11800 -332
rect 12200 444 12258 456
rect 12200 -332 12212 444
rect 12246 -332 12258 444
rect 12200 -344 12258 -332
rect 12330 444 12388 456
rect 12330 -332 12342 444
rect 12376 -332 12388 444
rect 12330 -344 12388 -332
rect 12788 444 12846 456
rect 12788 -332 12800 444
rect 12834 -332 12846 444
rect 12788 -344 12846 -332
rect 12918 444 12976 456
rect 12918 -332 12930 444
rect 12964 -332 12976 444
rect 12918 -344 12976 -332
rect 13376 444 13434 456
rect 13376 -332 13388 444
rect 13422 -332 13434 444
rect 13376 -344 13434 -332
rect 13506 444 13564 456
rect 13506 -332 13518 444
rect 13552 -332 13564 444
rect 13506 -344 13564 -332
rect 13964 444 14022 456
rect 13964 -332 13976 444
rect 14010 -332 14022 444
rect 13964 -344 14022 -332
rect 14094 444 14152 456
rect 14094 -332 14106 444
rect 14140 -332 14152 444
rect 14094 -344 14152 -332
rect 14552 444 14610 456
rect 14552 -332 14564 444
rect 14598 -332 14610 444
rect 14552 -344 14610 -332
rect 14682 444 14740 456
rect 14682 -332 14694 444
rect 14728 -332 14740 444
rect 14682 -344 14740 -332
rect 15140 444 15198 456
rect 15140 -332 15152 444
rect 15186 -332 15198 444
rect 15140 -344 15198 -332
rect 15270 444 15328 456
rect 15270 -332 15282 444
rect 15316 -332 15328 444
rect 15270 -344 15328 -332
rect 15728 444 15786 456
rect 15728 -332 15740 444
rect 15774 -332 15786 444
rect 15728 -344 15786 -332
rect 15858 444 15916 456
rect 15858 -332 15870 444
rect 15904 -332 15916 444
rect 15858 -344 15916 -332
rect 16316 444 16374 456
rect 16316 -332 16328 444
rect 16362 -332 16374 444
rect 16316 -344 16374 -332
rect 16446 444 16504 456
rect 16446 -332 16458 444
rect 16492 -332 16504 444
rect 16446 -344 16504 -332
rect 16904 444 16962 456
rect 16904 -332 16916 444
rect 16950 -332 16962 444
rect 16904 -344 16962 -332
rect 17034 444 17092 456
rect 17034 -332 17046 444
rect 17080 -332 17092 444
rect 17034 -344 17092 -332
rect 17492 444 17550 456
rect 17492 -332 17504 444
rect 17538 -332 17550 444
rect 17492 -344 17550 -332
rect 17622 444 17680 456
rect 17622 -332 17634 444
rect 17668 -332 17680 444
rect 17622 -344 17680 -332
rect 18080 444 18138 456
rect 18080 -332 18092 444
rect 18126 -332 18138 444
rect 18080 -344 18138 -332
rect 18210 444 18268 456
rect 18210 -332 18222 444
rect 18256 -332 18268 444
rect 18210 -344 18268 -332
rect 18668 444 18726 456
rect 18668 -332 18680 444
rect 18714 -332 18726 444
rect 18668 -344 18726 -332
rect 18798 444 18856 456
rect 18798 -332 18810 444
rect 18844 -332 18856 444
rect 18798 -344 18856 -332
rect 19256 444 19314 456
rect 19256 -332 19268 444
rect 19302 -332 19314 444
rect 19256 -344 19314 -332
rect 19386 444 19444 456
rect 19386 -332 19398 444
rect 19432 -332 19444 444
rect 19386 -344 19444 -332
rect 19844 444 19902 456
rect 19844 -332 19856 444
rect 19890 -332 19902 444
rect 19844 -344 19902 -332
rect 19974 444 20032 456
rect 19974 -332 19986 444
rect 20020 -332 20032 444
rect 19974 -344 20032 -332
rect 20432 444 20490 456
rect 20432 -332 20444 444
rect 20478 -332 20490 444
rect 20432 -344 20490 -332
rect 20562 444 20620 456
rect 20562 -332 20574 444
rect 20608 -332 20620 444
rect 20562 -344 20620 -332
rect 21020 444 21078 456
rect 21020 -332 21032 444
rect 21066 -332 21078 444
rect 21020 -344 21078 -332
rect 21150 444 21208 456
rect 21150 -332 21162 444
rect 21196 -332 21208 444
rect 21150 -344 21208 -332
rect 21608 444 21666 456
rect 21608 -332 21620 444
rect 21654 -332 21666 444
rect 21608 -344 21666 -332
rect 6566 -2002 6624 -1990
rect 6566 -2778 6578 -2002
rect 6612 -2778 6624 -2002
rect 6566 -2790 6624 -2778
rect 6694 -2002 6752 -1990
rect 6694 -2778 6706 -2002
rect 6740 -2778 6752 -2002
rect 6694 -2790 6752 -2778
rect 6832 -2002 6890 -1990
rect 6832 -2778 6844 -2002
rect 6878 -2778 6890 -2002
rect 6832 -2790 6890 -2778
rect 6960 -2002 7018 -1990
rect 6960 -2778 6972 -2002
rect 7006 -2778 7018 -2002
rect 6960 -2790 7018 -2778
rect 7098 -2002 7156 -1990
rect 7098 -2778 7110 -2002
rect 7144 -2778 7156 -2002
rect 7098 -2790 7156 -2778
rect 7226 -2002 7284 -1990
rect 7226 -2778 7238 -2002
rect 7272 -2778 7284 -2002
rect 7226 -2790 7284 -2778
rect 7364 -2002 7422 -1990
rect 7364 -2778 7376 -2002
rect 7410 -2778 7422 -2002
rect 7364 -2790 7422 -2778
rect 7492 -2002 7550 -1990
rect 7492 -2778 7504 -2002
rect 7538 -2778 7550 -2002
rect 7492 -2790 7550 -2778
rect 7630 -2002 7688 -1990
rect 7630 -2778 7642 -2002
rect 7676 -2778 7688 -2002
rect 7630 -2790 7688 -2778
rect 7758 -2002 7816 -1990
rect 7758 -2778 7770 -2002
rect 7804 -2778 7816 -2002
rect 7758 -2790 7816 -2778
rect 7896 -2002 7954 -1990
rect 7896 -2778 7908 -2002
rect 7942 -2778 7954 -2002
rect 7896 -2790 7954 -2778
rect 8024 -2002 8082 -1990
rect 8024 -2778 8036 -2002
rect 8070 -2778 8082 -2002
rect 8024 -2790 8082 -2778
rect 8162 -2002 8220 -1990
rect 8162 -2778 8174 -2002
rect 8208 -2778 8220 -2002
rect 8162 -2790 8220 -2778
rect 8290 -2002 8348 -1990
rect 8290 -2778 8302 -2002
rect 8336 -2778 8348 -2002
rect 8290 -2790 8348 -2778
rect 8428 -2002 8486 -1990
rect 8428 -2778 8440 -2002
rect 8474 -2778 8486 -2002
rect 8428 -2790 8486 -2778
rect 8556 -2002 8614 -1990
rect 8556 -2778 8568 -2002
rect 8602 -2778 8614 -2002
rect 8556 -2790 8614 -2778
rect 6566 -3012 6624 -3000
rect 6566 -3788 6578 -3012
rect 6612 -3788 6624 -3012
rect 6566 -3800 6624 -3788
rect 6694 -3012 6752 -3000
rect 6694 -3788 6706 -3012
rect 6740 -3788 6752 -3012
rect 6694 -3800 6752 -3788
rect 6832 -3012 6890 -3000
rect 6832 -3788 6844 -3012
rect 6878 -3788 6890 -3012
rect 6832 -3800 6890 -3788
rect 6960 -3012 7018 -3000
rect 6960 -3788 6972 -3012
rect 7006 -3788 7018 -3012
rect 6960 -3800 7018 -3788
rect 7098 -3012 7156 -3000
rect 7098 -3788 7110 -3012
rect 7144 -3788 7156 -3012
rect 7098 -3800 7156 -3788
rect 7226 -3012 7284 -3000
rect 7226 -3788 7238 -3012
rect 7272 -3788 7284 -3012
rect 7226 -3800 7284 -3788
rect 7364 -3012 7422 -3000
rect 7364 -3788 7376 -3012
rect 7410 -3788 7422 -3012
rect 7364 -3800 7422 -3788
rect 7492 -3012 7550 -3000
rect 7492 -3788 7504 -3012
rect 7538 -3788 7550 -3012
rect 7492 -3800 7550 -3788
rect 7630 -3012 7688 -3000
rect 7630 -3788 7642 -3012
rect 7676 -3788 7688 -3012
rect 7630 -3800 7688 -3788
rect 7758 -3012 7816 -3000
rect 7758 -3788 7770 -3012
rect 7804 -3788 7816 -3012
rect 7758 -3800 7816 -3788
rect 7896 -3012 7954 -3000
rect 7896 -3788 7908 -3012
rect 7942 -3788 7954 -3012
rect 7896 -3800 7954 -3788
rect 8024 -3012 8082 -3000
rect 8024 -3788 8036 -3012
rect 8070 -3788 8082 -3012
rect 8024 -3800 8082 -3788
rect 8162 -3012 8220 -3000
rect 8162 -3788 8174 -3012
rect 8208 -3788 8220 -3012
rect 8162 -3800 8220 -3788
rect 8290 -3012 8348 -3000
rect 8290 -3788 8302 -3012
rect 8336 -3788 8348 -3012
rect 8290 -3800 8348 -3788
rect 8428 -3012 8486 -3000
rect 8428 -3788 8440 -3012
rect 8474 -3788 8486 -3012
rect 8428 -3800 8486 -3788
rect 8556 -3012 8614 -3000
rect 8556 -3788 8568 -3012
rect 8602 -3788 8614 -3012
rect 8556 -3800 8614 -3788
rect 6566 -4022 6624 -4010
rect 6566 -4798 6578 -4022
rect 6612 -4798 6624 -4022
rect 6566 -4810 6624 -4798
rect 6694 -4022 6752 -4010
rect 6694 -4798 6706 -4022
rect 6740 -4798 6752 -4022
rect 6694 -4810 6752 -4798
rect 6832 -4022 6890 -4010
rect 6832 -4798 6844 -4022
rect 6878 -4798 6890 -4022
rect 6832 -4810 6890 -4798
rect 6960 -4022 7018 -4010
rect 6960 -4798 6972 -4022
rect 7006 -4798 7018 -4022
rect 6960 -4810 7018 -4798
rect 7098 -4022 7156 -4010
rect 7098 -4798 7110 -4022
rect 7144 -4798 7156 -4022
rect 7098 -4810 7156 -4798
rect 7226 -4022 7284 -4010
rect 7226 -4798 7238 -4022
rect 7272 -4798 7284 -4022
rect 7226 -4810 7284 -4798
rect 7364 -4022 7422 -4010
rect 7364 -4798 7376 -4022
rect 7410 -4798 7422 -4022
rect 7364 -4810 7422 -4798
rect 7492 -4022 7550 -4010
rect 7492 -4798 7504 -4022
rect 7538 -4798 7550 -4022
rect 7492 -4810 7550 -4798
rect 7630 -4022 7688 -4010
rect 7630 -4798 7642 -4022
rect 7676 -4798 7688 -4022
rect 7630 -4810 7688 -4798
rect 7758 -4022 7816 -4010
rect 7758 -4798 7770 -4022
rect 7804 -4798 7816 -4022
rect 7758 -4810 7816 -4798
rect 7896 -4022 7954 -4010
rect 7896 -4798 7908 -4022
rect 7942 -4798 7954 -4022
rect 7896 -4810 7954 -4798
rect 8024 -4022 8082 -4010
rect 8024 -4798 8036 -4022
rect 8070 -4798 8082 -4022
rect 8024 -4810 8082 -4798
rect 8162 -4022 8220 -4010
rect 8162 -4798 8174 -4022
rect 8208 -4798 8220 -4022
rect 8162 -4810 8220 -4798
rect 8290 -4022 8348 -4010
rect 8290 -4798 8302 -4022
rect 8336 -4798 8348 -4022
rect 8290 -4810 8348 -4798
rect 8428 -4022 8486 -4010
rect 8428 -4798 8440 -4022
rect 8474 -4798 8486 -4022
rect 8428 -4810 8486 -4798
rect 8556 -4022 8614 -4010
rect 8556 -4798 8568 -4022
rect 8602 -4798 8614 -4022
rect 8556 -4810 8614 -4798
<< ndiffc >>
rect 2830 5988 2864 6564
rect 2958 5988 2992 6564
rect 3070 5988 3104 6564
rect 3198 5988 3232 6564
rect 3310 5988 3344 6564
rect 3438 5988 3472 6564
rect 3550 5988 3584 6564
rect 3678 5988 3712 6564
rect 3790 5988 3824 6564
rect 3918 5988 3952 6564
rect 4030 5988 4064 6564
rect 4158 5988 4192 6564
rect 4270 5988 4304 6564
rect 4398 5988 4432 6564
rect 4510 5988 4544 6564
rect 4638 5988 4672 6564
rect 4750 5988 4784 6564
rect 4878 5988 4912 6564
rect 4990 5988 5024 6564
rect 5118 5988 5152 6564
rect 5230 5988 5264 6564
rect 5358 5988 5392 6564
rect 5470 5988 5504 6564
rect 5598 5988 5632 6564
rect 5710 5988 5744 6564
rect 5838 5988 5872 6564
rect 5950 5988 5984 6564
rect 6078 5988 6112 6564
rect 6190 5988 6224 6564
rect 6318 5988 6352 6564
rect 6430 5988 6464 6564
rect 6558 5988 6592 6564
rect 6670 5988 6704 6564
rect 6798 5988 6832 6564
rect 6910 5988 6944 6564
rect 7038 5988 7072 6564
rect 7150 5988 7184 6564
rect 7278 5988 7312 6564
rect 7390 5988 7424 6564
rect 7518 5988 7552 6564
rect 7630 5988 7664 6564
rect 7758 5988 7792 6564
rect 7870 5988 7904 6564
rect 7998 5988 8032 6564
rect 8110 5988 8144 6564
rect 8238 5988 8272 6564
rect 8350 5988 8384 6564
rect 8478 5988 8512 6564
rect 8590 5988 8624 6564
rect 8718 5988 8752 6564
rect 8830 5988 8864 6564
rect 8958 5988 8992 6564
rect 9070 5988 9104 6564
rect 9198 5988 9232 6564
rect 9310 5988 9344 6564
rect 9438 5988 9472 6564
rect 9550 5988 9584 6564
rect 9678 5988 9712 6564
rect 9790 5988 9824 6564
rect 9918 5988 9952 6564
rect 10030 5988 10064 6564
rect 10158 5988 10192 6564
rect 10270 5988 10304 6564
rect 10398 5988 10432 6564
rect 10510 5988 10544 6564
rect 10638 5988 10672 6564
rect 10750 5988 10784 6564
rect 10878 5988 10912 6564
rect 10990 5988 11024 6564
rect 11118 5988 11152 6564
rect 11230 5988 11264 6564
rect 11358 5988 11392 6564
rect 11470 5988 11504 6564
rect 11598 5988 11632 6564
rect 11710 5988 11744 6564
rect 11838 5988 11872 6564
rect 11950 5988 11984 6564
rect 12078 5988 12112 6564
rect 12190 5988 12224 6564
rect 12318 5988 12352 6564
rect 2830 5180 2864 5756
rect 2958 5180 2992 5756
rect 3070 5180 3104 5756
rect 3198 5180 3232 5756
rect 3310 5180 3344 5756
rect 3438 5180 3472 5756
rect 3550 5180 3584 5756
rect 3678 5180 3712 5756
rect 3790 5180 3824 5756
rect 3918 5180 3952 5756
rect 4030 5180 4064 5756
rect 4158 5180 4192 5756
rect 4270 5180 4304 5756
rect 4398 5180 4432 5756
rect 4510 5180 4544 5756
rect 4638 5180 4672 5756
rect 4750 5180 4784 5756
rect 4878 5180 4912 5756
rect 4990 5180 5024 5756
rect 5118 5180 5152 5756
rect 5230 5180 5264 5756
rect 5358 5180 5392 5756
rect 5470 5180 5504 5756
rect 5598 5180 5632 5756
rect 5710 5180 5744 5756
rect 5838 5180 5872 5756
rect 5950 5180 5984 5756
rect 6078 5180 6112 5756
rect 6190 5180 6224 5756
rect 6318 5180 6352 5756
rect 6430 5180 6464 5756
rect 6558 5180 6592 5756
rect 6670 5180 6704 5756
rect 6798 5180 6832 5756
rect 6910 5180 6944 5756
rect 7038 5180 7072 5756
rect 7150 5180 7184 5756
rect 7278 5180 7312 5756
rect 7390 5180 7424 5756
rect 7518 5180 7552 5756
rect 7630 5180 7664 5756
rect 7758 5180 7792 5756
rect 7870 5180 7904 5756
rect 7998 5180 8032 5756
rect 8110 5180 8144 5756
rect 8238 5180 8272 5756
rect 8350 5180 8384 5756
rect 8478 5180 8512 5756
rect 8590 5180 8624 5756
rect 8718 5180 8752 5756
rect 8830 5180 8864 5756
rect 8958 5180 8992 5756
rect 9070 5180 9104 5756
rect 9198 5180 9232 5756
rect 9310 5180 9344 5756
rect 9438 5180 9472 5756
rect 9550 5180 9584 5756
rect 9678 5180 9712 5756
rect 9790 5180 9824 5756
rect 9918 5180 9952 5756
rect 10030 5180 10064 5756
rect 10158 5180 10192 5756
rect 10270 5180 10304 5756
rect 10398 5180 10432 5756
rect 10510 5180 10544 5756
rect 10638 5180 10672 5756
rect 10750 5180 10784 5756
rect 10878 5180 10912 5756
rect 10990 5180 11024 5756
rect 11118 5180 11152 5756
rect 11230 5180 11264 5756
rect 11358 5180 11392 5756
rect 11470 5180 11504 5756
rect 11598 5180 11632 5756
rect 11710 5180 11744 5756
rect 11838 5180 11872 5756
rect 11950 5180 11984 5756
rect 12078 5180 12112 5756
rect 12190 5180 12224 5756
rect 12318 5180 12352 5756
rect 7150 -6770 7184 -6194
rect 7278 -6770 7312 -6194
rect 7390 -6770 7424 -6194
rect 7518 -6770 7552 -6194
rect 7630 -6770 7664 -6194
rect 7758 -6770 7792 -6194
rect 7870 -6770 7904 -6194
rect 7998 -6770 8032 -6194
rect 7150 -7578 7184 -7002
rect 7278 -7578 7312 -7002
rect 7390 -7578 7424 -7002
rect 7518 -7578 7552 -7002
rect 7630 -7578 7664 -7002
rect 7758 -7578 7792 -7002
rect 7870 -7578 7904 -7002
rect 7998 -7578 8032 -7002
<< pdiffc >>
rect -6474 1668 -6440 2444
rect -6016 1668 -5982 2444
rect -5886 1668 -5852 2444
rect -5428 1668 -5394 2444
rect -5298 1668 -5264 2444
rect -4840 1668 -4806 2444
rect -4710 1668 -4676 2444
rect -4252 1668 -4218 2444
rect -4122 1668 -4088 2444
rect -3664 1668 -3630 2444
rect -3534 1668 -3500 2444
rect -3076 1668 -3042 2444
rect -2946 1668 -2912 2444
rect -2488 1668 -2454 2444
rect -2358 1668 -2324 2444
rect -1900 1668 -1866 2444
rect -1770 1668 -1736 2444
rect -1312 1668 -1278 2444
rect -1182 1668 -1148 2444
rect -724 1668 -690 2444
rect -594 1668 -560 2444
rect -136 1668 -102 2444
rect -6 1668 28 2444
rect 452 1668 486 2444
rect 582 1668 616 2444
rect 1040 1668 1074 2444
rect 1170 1668 1204 2444
rect 1628 1668 1662 2444
rect 1758 1668 1792 2444
rect 2216 1668 2250 2444
rect 2346 1668 2380 2444
rect 2804 1668 2838 2444
rect 2934 1668 2968 2444
rect 3392 1668 3426 2444
rect 3522 1668 3556 2444
rect 3980 1668 4014 2444
rect 4110 1668 4144 2444
rect 4568 1668 4602 2444
rect 4698 1668 4732 2444
rect 5156 1668 5190 2444
rect 5286 1668 5320 2444
rect 5744 1668 5778 2444
rect 5874 1668 5908 2444
rect 6332 1668 6366 2444
rect 6462 1668 6496 2444
rect 6920 1668 6954 2444
rect 7050 1668 7084 2444
rect 7508 1668 7542 2444
rect 7638 1668 7672 2444
rect 8096 1668 8130 2444
rect 8226 1668 8260 2444
rect 8684 1668 8718 2444
rect 8814 1668 8848 2444
rect 9272 1668 9306 2444
rect 9402 1668 9436 2444
rect 9860 1668 9894 2444
rect 9990 1668 10024 2444
rect 10448 1668 10482 2444
rect 10578 1668 10612 2444
rect 11036 1668 11070 2444
rect 11166 1668 11200 2444
rect 11624 1668 11658 2444
rect 11754 1668 11788 2444
rect 12212 1668 12246 2444
rect 12342 1668 12376 2444
rect 12800 1668 12834 2444
rect 12930 1668 12964 2444
rect 13388 1668 13422 2444
rect 13518 1668 13552 2444
rect 13976 1668 14010 2444
rect 14106 1668 14140 2444
rect 14564 1668 14598 2444
rect 14694 1668 14728 2444
rect 15152 1668 15186 2444
rect 15282 1668 15316 2444
rect 15740 1668 15774 2444
rect 15870 1668 15904 2444
rect 16328 1668 16362 2444
rect 16458 1668 16492 2444
rect 16916 1668 16950 2444
rect 17046 1668 17080 2444
rect 17504 1668 17538 2444
rect 17634 1668 17668 2444
rect 18092 1668 18126 2444
rect 18222 1668 18256 2444
rect 18680 1668 18714 2444
rect 18810 1668 18844 2444
rect 19268 1668 19302 2444
rect 19398 1668 19432 2444
rect 19856 1668 19890 2444
rect 19986 1668 20020 2444
rect 20444 1668 20478 2444
rect 20574 1668 20608 2444
rect 21032 1668 21066 2444
rect 21162 1668 21196 2444
rect 21620 1668 21654 2444
rect -6474 668 -6440 1444
rect -6016 668 -5982 1444
rect -5886 668 -5852 1444
rect -5428 668 -5394 1444
rect -5298 668 -5264 1444
rect -4840 668 -4806 1444
rect -4710 668 -4676 1444
rect -4252 668 -4218 1444
rect -4122 668 -4088 1444
rect -3664 668 -3630 1444
rect -3534 668 -3500 1444
rect -3076 668 -3042 1444
rect -2946 668 -2912 1444
rect -2488 668 -2454 1444
rect -2358 668 -2324 1444
rect -1900 668 -1866 1444
rect -1770 668 -1736 1444
rect -1312 668 -1278 1444
rect -1182 668 -1148 1444
rect -724 668 -690 1444
rect -594 668 -560 1444
rect -136 668 -102 1444
rect -6 668 28 1444
rect 452 668 486 1444
rect 582 668 616 1444
rect 1040 668 1074 1444
rect 1170 668 1204 1444
rect 1628 668 1662 1444
rect 1758 668 1792 1444
rect 2216 668 2250 1444
rect 2346 668 2380 1444
rect 2804 668 2838 1444
rect 2934 668 2968 1444
rect 3392 668 3426 1444
rect 3522 668 3556 1444
rect 3980 668 4014 1444
rect 4110 668 4144 1444
rect 4568 668 4602 1444
rect 4698 668 4732 1444
rect 5156 668 5190 1444
rect 5286 668 5320 1444
rect 5744 668 5778 1444
rect 5874 668 5908 1444
rect 6332 668 6366 1444
rect 6462 668 6496 1444
rect 6920 668 6954 1444
rect 7050 668 7084 1444
rect 7508 668 7542 1444
rect 7638 668 7672 1444
rect 8096 668 8130 1444
rect 8226 668 8260 1444
rect 8684 668 8718 1444
rect 8814 668 8848 1444
rect 9272 668 9306 1444
rect 9402 668 9436 1444
rect 9860 668 9894 1444
rect 9990 668 10024 1444
rect 10448 668 10482 1444
rect 10578 668 10612 1444
rect 11036 668 11070 1444
rect 11166 668 11200 1444
rect 11624 668 11658 1444
rect 11754 668 11788 1444
rect 12212 668 12246 1444
rect 12342 668 12376 1444
rect 12800 668 12834 1444
rect 12930 668 12964 1444
rect 13388 668 13422 1444
rect 13518 668 13552 1444
rect 13976 668 14010 1444
rect 14106 668 14140 1444
rect 14564 668 14598 1444
rect 14694 668 14728 1444
rect 15152 668 15186 1444
rect 15282 668 15316 1444
rect 15740 668 15774 1444
rect 15870 668 15904 1444
rect 16328 668 16362 1444
rect 16458 668 16492 1444
rect 16916 668 16950 1444
rect 17046 668 17080 1444
rect 17504 668 17538 1444
rect 17634 668 17668 1444
rect 18092 668 18126 1444
rect 18222 668 18256 1444
rect 18680 668 18714 1444
rect 18810 668 18844 1444
rect 19268 668 19302 1444
rect 19398 668 19432 1444
rect 19856 668 19890 1444
rect 19986 668 20020 1444
rect 20444 668 20478 1444
rect 20574 668 20608 1444
rect 21032 668 21066 1444
rect 21162 668 21196 1444
rect 21620 668 21654 1444
rect -6474 -332 -6440 444
rect -6016 -332 -5982 444
rect -5886 -332 -5852 444
rect -5428 -332 -5394 444
rect -5298 -332 -5264 444
rect -4840 -332 -4806 444
rect -4710 -332 -4676 444
rect -4252 -332 -4218 444
rect -4122 -332 -4088 444
rect -3664 -332 -3630 444
rect -3534 -332 -3500 444
rect -3076 -332 -3042 444
rect -2946 -332 -2912 444
rect -2488 -332 -2454 444
rect -2358 -332 -2324 444
rect -1900 -332 -1866 444
rect -1770 -332 -1736 444
rect -1312 -332 -1278 444
rect -1182 -332 -1148 444
rect -724 -332 -690 444
rect -594 -332 -560 444
rect -136 -332 -102 444
rect -6 -332 28 444
rect 452 -332 486 444
rect 582 -332 616 444
rect 1040 -332 1074 444
rect 1170 -332 1204 444
rect 1628 -332 1662 444
rect 1758 -332 1792 444
rect 2216 -332 2250 444
rect 2346 -332 2380 444
rect 2804 -332 2838 444
rect 2934 -332 2968 444
rect 3392 -332 3426 444
rect 3522 -332 3556 444
rect 3980 -332 4014 444
rect 4110 -332 4144 444
rect 4568 -332 4602 444
rect 4698 -332 4732 444
rect 5156 -332 5190 444
rect 5286 -332 5320 444
rect 5744 -332 5778 444
rect 5874 -332 5908 444
rect 6332 -332 6366 444
rect 6462 -332 6496 444
rect 6920 -332 6954 444
rect 7050 -332 7084 444
rect 7508 -332 7542 444
rect 7638 -332 7672 444
rect 8096 -332 8130 444
rect 8226 -332 8260 444
rect 8684 -332 8718 444
rect 8814 -332 8848 444
rect 9272 -332 9306 444
rect 9402 -332 9436 444
rect 9860 -332 9894 444
rect 9990 -332 10024 444
rect 10448 -332 10482 444
rect 10578 -332 10612 444
rect 11036 -332 11070 444
rect 11166 -332 11200 444
rect 11624 -332 11658 444
rect 11754 -332 11788 444
rect 12212 -332 12246 444
rect 12342 -332 12376 444
rect 12800 -332 12834 444
rect 12930 -332 12964 444
rect 13388 -332 13422 444
rect 13518 -332 13552 444
rect 13976 -332 14010 444
rect 14106 -332 14140 444
rect 14564 -332 14598 444
rect 14694 -332 14728 444
rect 15152 -332 15186 444
rect 15282 -332 15316 444
rect 15740 -332 15774 444
rect 15870 -332 15904 444
rect 16328 -332 16362 444
rect 16458 -332 16492 444
rect 16916 -332 16950 444
rect 17046 -332 17080 444
rect 17504 -332 17538 444
rect 17634 -332 17668 444
rect 18092 -332 18126 444
rect 18222 -332 18256 444
rect 18680 -332 18714 444
rect 18810 -332 18844 444
rect 19268 -332 19302 444
rect 19398 -332 19432 444
rect 19856 -332 19890 444
rect 19986 -332 20020 444
rect 20444 -332 20478 444
rect 20574 -332 20608 444
rect 21032 -332 21066 444
rect 21162 -332 21196 444
rect 21620 -332 21654 444
rect 6578 -2778 6612 -2002
rect 6706 -2778 6740 -2002
rect 6844 -2778 6878 -2002
rect 6972 -2778 7006 -2002
rect 7110 -2778 7144 -2002
rect 7238 -2778 7272 -2002
rect 7376 -2778 7410 -2002
rect 7504 -2778 7538 -2002
rect 7642 -2778 7676 -2002
rect 7770 -2778 7804 -2002
rect 7908 -2778 7942 -2002
rect 8036 -2778 8070 -2002
rect 8174 -2778 8208 -2002
rect 8302 -2778 8336 -2002
rect 8440 -2778 8474 -2002
rect 8568 -2778 8602 -2002
rect 6578 -3788 6612 -3012
rect 6706 -3788 6740 -3012
rect 6844 -3788 6878 -3012
rect 6972 -3788 7006 -3012
rect 7110 -3788 7144 -3012
rect 7238 -3788 7272 -3012
rect 7376 -3788 7410 -3012
rect 7504 -3788 7538 -3012
rect 7642 -3788 7676 -3012
rect 7770 -3788 7804 -3012
rect 7908 -3788 7942 -3012
rect 8036 -3788 8070 -3012
rect 8174 -3788 8208 -3012
rect 8302 -3788 8336 -3012
rect 8440 -3788 8474 -3012
rect 8568 -3788 8602 -3012
rect 6578 -4798 6612 -4022
rect 6706 -4798 6740 -4022
rect 6844 -4798 6878 -4022
rect 6972 -4798 7006 -4022
rect 7110 -4798 7144 -4022
rect 7238 -4798 7272 -4022
rect 7376 -4798 7410 -4022
rect 7504 -4798 7538 -4022
rect 7642 -4798 7676 -4022
rect 7770 -4798 7804 -4022
rect 7908 -4798 7942 -4022
rect 8036 -4798 8070 -4022
rect 8174 -4798 8208 -4022
rect 8302 -4798 8336 -4022
rect 8440 -4798 8474 -4022
rect 8568 -4798 8602 -4022
<< psubdiff >>
rect 13613 -3401 13709 -3367
rect 13847 -3401 13943 -3367
rect 13613 -3463 13647 -3401
rect 13909 -3463 13943 -3401
rect 13613 -5017 13647 -4955
rect 13909 -5017 13943 -4955
rect 13613 -5051 13709 -5017
rect 13847 -5051 13943 -5017
<< nsubdiff >>
rect 6192 -1520 6226 -1486
rect 8954 -1520 8988 -1486
rect 6192 -5316 6226 -5282
rect 8954 -5316 8988 -5282
<< psubdiffcont >>
rect 2572 7056 12610 7090
rect 2484 4742 2518 7022
rect 12664 4742 12698 7024
rect 2518 4654 12664 4688
rect 13709 -3401 13847 -3367
rect 13613 -4955 13647 -3463
rect 13909 -4955 13943 -3463
rect 13709 -5051 13847 -5017
rect 6950 -5712 8160 -5678
rect 6804 -8060 6838 -5712
rect 8344 -8060 8378 -5712
rect 6962 -8094 8172 -8060
<< nsubdiffcont >>
rect -6660 2854 21862 2888
rect -6820 -722 -6786 2826
rect 21966 -688 22000 2860
rect -6702 -776 21912 -742
rect 6226 -1520 8954 -1486
rect 6192 -5282 6226 -1520
rect 8954 -5282 8988 -1520
rect 6226 -5316 8954 -5282
<< poly >>
rect 2876 6746 2946 6756
rect 2876 6614 2892 6746
rect 2930 6614 2946 6746
rect 2876 6576 2946 6614
rect 3116 6746 3186 6756
rect 3116 6614 3132 6746
rect 3170 6614 3186 6746
rect 3116 6576 3186 6614
rect 3356 6746 3426 6756
rect 3356 6614 3372 6746
rect 3410 6614 3426 6746
rect 3356 6576 3426 6614
rect 3596 6746 3666 6756
rect 3596 6614 3612 6746
rect 3650 6614 3666 6746
rect 3596 6576 3666 6614
rect 3836 6746 3906 6756
rect 3836 6614 3852 6746
rect 3890 6614 3906 6746
rect 3836 6576 3906 6614
rect 4076 6746 4146 6756
rect 4076 6614 4092 6746
rect 4130 6614 4146 6746
rect 4076 6576 4146 6614
rect 4316 6746 4386 6756
rect 4316 6614 4332 6746
rect 4370 6614 4386 6746
rect 4316 6576 4386 6614
rect 4556 6746 4626 6756
rect 4556 6614 4572 6746
rect 4610 6614 4626 6746
rect 4556 6576 4626 6614
rect 4796 6746 4866 6756
rect 4796 6614 4812 6746
rect 4850 6614 4866 6746
rect 4796 6576 4866 6614
rect 5036 6746 5106 6756
rect 5036 6614 5052 6746
rect 5090 6614 5106 6746
rect 5036 6576 5106 6614
rect 5276 6746 5346 6756
rect 5276 6614 5292 6746
rect 5330 6614 5346 6746
rect 5276 6576 5346 6614
rect 5516 6746 5586 6756
rect 5516 6614 5532 6746
rect 5570 6614 5586 6746
rect 5516 6576 5586 6614
rect 5756 6746 5826 6756
rect 5756 6614 5772 6746
rect 5810 6614 5826 6746
rect 5756 6576 5826 6614
rect 5996 6746 6066 6756
rect 5996 6614 6012 6746
rect 6050 6614 6066 6746
rect 5996 6576 6066 6614
rect 6236 6746 6306 6756
rect 6236 6614 6252 6746
rect 6290 6614 6306 6746
rect 6236 6576 6306 6614
rect 6476 6746 6546 6756
rect 6476 6614 6492 6746
rect 6530 6614 6546 6746
rect 6476 6576 6546 6614
rect 6716 6746 6786 6756
rect 6716 6614 6732 6746
rect 6770 6614 6786 6746
rect 6716 6576 6786 6614
rect 6956 6746 7026 6756
rect 6956 6614 6972 6746
rect 7010 6614 7026 6746
rect 6956 6576 7026 6614
rect 7196 6746 7266 6756
rect 7196 6614 7212 6746
rect 7250 6614 7266 6746
rect 7196 6576 7266 6614
rect 7436 6746 7506 6756
rect 7436 6614 7452 6746
rect 7490 6614 7506 6746
rect 7436 6576 7506 6614
rect 7676 6746 7746 6756
rect 7676 6614 7692 6746
rect 7730 6614 7746 6746
rect 7676 6576 7746 6614
rect 7916 6746 7986 6756
rect 7916 6614 7932 6746
rect 7970 6614 7986 6746
rect 7916 6576 7986 6614
rect 8156 6746 8226 6756
rect 8156 6614 8172 6746
rect 8210 6614 8226 6746
rect 8156 6576 8226 6614
rect 8396 6746 8466 6756
rect 8396 6614 8412 6746
rect 8450 6614 8466 6746
rect 8396 6576 8466 6614
rect 8636 6746 8706 6756
rect 8636 6614 8652 6746
rect 8690 6614 8706 6746
rect 8636 6576 8706 6614
rect 8876 6746 8946 6756
rect 8876 6614 8892 6746
rect 8930 6614 8946 6746
rect 8876 6576 8946 6614
rect 9116 6746 9186 6756
rect 9116 6614 9132 6746
rect 9170 6614 9186 6746
rect 9116 6576 9186 6614
rect 9356 6746 9426 6756
rect 9356 6614 9372 6746
rect 9410 6614 9426 6746
rect 9356 6576 9426 6614
rect 9596 6746 9666 6756
rect 9596 6614 9612 6746
rect 9650 6614 9666 6746
rect 9596 6576 9666 6614
rect 9836 6746 9906 6756
rect 9836 6614 9852 6746
rect 9890 6614 9906 6746
rect 9836 6576 9906 6614
rect 10076 6746 10146 6756
rect 10076 6614 10092 6746
rect 10130 6614 10146 6746
rect 10076 6576 10146 6614
rect 10316 6746 10386 6756
rect 10316 6614 10332 6746
rect 10370 6614 10386 6746
rect 10316 6576 10386 6614
rect 10556 6746 10626 6756
rect 10556 6614 10572 6746
rect 10610 6614 10626 6746
rect 10556 6576 10626 6614
rect 10796 6746 10866 6756
rect 10796 6614 10812 6746
rect 10850 6614 10866 6746
rect 10796 6576 10866 6614
rect 11036 6746 11106 6756
rect 11036 6614 11052 6746
rect 11090 6614 11106 6746
rect 11036 6576 11106 6614
rect 11276 6746 11346 6756
rect 11276 6614 11292 6746
rect 11330 6614 11346 6746
rect 11276 6576 11346 6614
rect 11516 6746 11586 6756
rect 11516 6614 11532 6746
rect 11570 6614 11586 6746
rect 11516 6576 11586 6614
rect 11756 6746 11826 6756
rect 11756 6614 11772 6746
rect 11810 6614 11826 6746
rect 11756 6576 11826 6614
rect 11996 6746 12066 6756
rect 11996 6614 12012 6746
rect 12050 6614 12066 6746
rect 11996 6576 12066 6614
rect 12236 6746 12306 6756
rect 12236 6614 12252 6746
rect 12290 6614 12306 6746
rect 12236 6576 12306 6614
rect 2876 5938 2946 5976
rect 2876 5806 2892 5938
rect 2930 5806 2946 5938
rect 2876 5768 2946 5806
rect 3116 5938 3186 5976
rect 3116 5806 3132 5938
rect 3170 5806 3186 5938
rect 3116 5768 3186 5806
rect 3356 5938 3426 5976
rect 3356 5806 3372 5938
rect 3410 5806 3426 5938
rect 3356 5768 3426 5806
rect 3596 5938 3666 5976
rect 3596 5806 3612 5938
rect 3650 5806 3666 5938
rect 3596 5768 3666 5806
rect 3836 5938 3906 5976
rect 3836 5806 3852 5938
rect 3890 5806 3906 5938
rect 3836 5768 3906 5806
rect 4076 5938 4146 5976
rect 4076 5806 4092 5938
rect 4130 5806 4146 5938
rect 4076 5768 4146 5806
rect 4316 5938 4386 5976
rect 4316 5806 4332 5938
rect 4370 5806 4386 5938
rect 4316 5768 4386 5806
rect 4556 5938 4626 5976
rect 4556 5806 4572 5938
rect 4610 5806 4626 5938
rect 4556 5768 4626 5806
rect 4796 5938 4866 5976
rect 4796 5806 4812 5938
rect 4850 5806 4866 5938
rect 4796 5768 4866 5806
rect 5036 5938 5106 5976
rect 5036 5806 5052 5938
rect 5090 5806 5106 5938
rect 5036 5768 5106 5806
rect 5276 5938 5346 5976
rect 5276 5806 5292 5938
rect 5330 5806 5346 5938
rect 5276 5768 5346 5806
rect 5516 5938 5586 5976
rect 5516 5806 5532 5938
rect 5570 5806 5586 5938
rect 5516 5768 5586 5806
rect 5756 5938 5826 5976
rect 5756 5806 5772 5938
rect 5810 5806 5826 5938
rect 5756 5768 5826 5806
rect 5996 5938 6066 5976
rect 5996 5806 6012 5938
rect 6050 5806 6066 5938
rect 5996 5768 6066 5806
rect 6236 5938 6306 5976
rect 6236 5806 6252 5938
rect 6290 5806 6306 5938
rect 6236 5768 6306 5806
rect 6476 5938 6546 5976
rect 6476 5806 6492 5938
rect 6530 5806 6546 5938
rect 6476 5768 6546 5806
rect 6716 5938 6786 5976
rect 6716 5806 6732 5938
rect 6770 5806 6786 5938
rect 6716 5768 6786 5806
rect 6956 5938 7026 5976
rect 6956 5806 6972 5938
rect 7010 5806 7026 5938
rect 6956 5768 7026 5806
rect 7196 5938 7266 5976
rect 7196 5806 7212 5938
rect 7250 5806 7266 5938
rect 7196 5768 7266 5806
rect 7436 5938 7506 5976
rect 7436 5806 7452 5938
rect 7490 5806 7506 5938
rect 7436 5768 7506 5806
rect 7676 5938 7746 5976
rect 7676 5806 7692 5938
rect 7730 5806 7746 5938
rect 7676 5768 7746 5806
rect 7916 5938 7986 5976
rect 7916 5806 7932 5938
rect 7970 5806 7986 5938
rect 7916 5768 7986 5806
rect 8156 5938 8226 5976
rect 8156 5806 8172 5938
rect 8210 5806 8226 5938
rect 8156 5768 8226 5806
rect 8396 5938 8466 5976
rect 8396 5806 8412 5938
rect 8450 5806 8466 5938
rect 8396 5768 8466 5806
rect 8636 5938 8706 5976
rect 8636 5806 8652 5938
rect 8690 5806 8706 5938
rect 8636 5768 8706 5806
rect 8876 5938 8946 5976
rect 8876 5806 8892 5938
rect 8930 5806 8946 5938
rect 8876 5768 8946 5806
rect 9116 5938 9186 5976
rect 9116 5806 9132 5938
rect 9170 5806 9186 5938
rect 9116 5768 9186 5806
rect 9356 5938 9426 5976
rect 9356 5806 9372 5938
rect 9410 5806 9426 5938
rect 9356 5768 9426 5806
rect 9596 5938 9666 5976
rect 9596 5806 9612 5938
rect 9650 5806 9666 5938
rect 9596 5768 9666 5806
rect 9836 5938 9906 5976
rect 9836 5806 9852 5938
rect 9890 5806 9906 5938
rect 9836 5768 9906 5806
rect 10076 5938 10146 5976
rect 10076 5806 10092 5938
rect 10130 5806 10146 5938
rect 10076 5768 10146 5806
rect 10316 5938 10386 5976
rect 10316 5806 10332 5938
rect 10370 5806 10386 5938
rect 10316 5768 10386 5806
rect 10556 5938 10626 5976
rect 10556 5806 10572 5938
rect 10610 5806 10626 5938
rect 10556 5768 10626 5806
rect 10796 5938 10866 5976
rect 10796 5806 10812 5938
rect 10850 5806 10866 5938
rect 10796 5768 10866 5806
rect 11036 5938 11106 5976
rect 11036 5806 11052 5938
rect 11090 5806 11106 5938
rect 11036 5768 11106 5806
rect 11276 5938 11346 5976
rect 11276 5806 11292 5938
rect 11330 5806 11346 5938
rect 11276 5768 11346 5806
rect 11516 5938 11586 5976
rect 11516 5806 11532 5938
rect 11570 5806 11586 5938
rect 11516 5768 11586 5806
rect 11756 5938 11826 5976
rect 11756 5806 11772 5938
rect 11810 5806 11826 5938
rect 11756 5768 11826 5806
rect 11996 5938 12066 5976
rect 11996 5806 12012 5938
rect 12050 5806 12066 5938
rect 11996 5768 12066 5806
rect 12236 5938 12306 5976
rect 12236 5806 12252 5938
rect 12290 5806 12306 5938
rect 12236 5768 12306 5806
rect 2876 5130 2946 5168
rect 2876 4998 2892 5130
rect 2930 4998 2946 5130
rect 2876 4988 2946 4998
rect 3116 5130 3186 5168
rect 3116 4998 3132 5130
rect 3170 4998 3186 5130
rect 3116 4988 3186 4998
rect 3356 5130 3426 5168
rect 3356 4998 3372 5130
rect 3410 4998 3426 5130
rect 3356 4988 3426 4998
rect 3596 5130 3666 5168
rect 3596 4998 3612 5130
rect 3650 4998 3666 5130
rect 3596 4988 3666 4998
rect 3836 5130 3906 5168
rect 3836 4998 3852 5130
rect 3890 4998 3906 5130
rect 3836 4988 3906 4998
rect 4076 5130 4146 5168
rect 4076 4998 4092 5130
rect 4130 4998 4146 5130
rect 4076 4988 4146 4998
rect 4316 5130 4386 5168
rect 4316 4998 4332 5130
rect 4370 4998 4386 5130
rect 4316 4988 4386 4998
rect 4556 5130 4626 5168
rect 4556 4998 4572 5130
rect 4610 4998 4626 5130
rect 4556 4988 4626 4998
rect 4796 5130 4866 5168
rect 4796 4998 4812 5130
rect 4850 4998 4866 5130
rect 4796 4988 4866 4998
rect 5036 5130 5106 5168
rect 5036 4998 5052 5130
rect 5090 4998 5106 5130
rect 5036 4988 5106 4998
rect 5276 5130 5346 5168
rect 5276 4998 5292 5130
rect 5330 4998 5346 5130
rect 5276 4988 5346 4998
rect 5516 5130 5586 5168
rect 5516 4998 5532 5130
rect 5570 4998 5586 5130
rect 5516 4988 5586 4998
rect 5756 5130 5826 5168
rect 5756 4998 5772 5130
rect 5810 4998 5826 5130
rect 5756 4988 5826 4998
rect 5996 5130 6066 5168
rect 5996 4998 6012 5130
rect 6050 4998 6066 5130
rect 5996 4988 6066 4998
rect 6236 5130 6306 5168
rect 6236 4998 6252 5130
rect 6290 4998 6306 5130
rect 6236 4988 6306 4998
rect 6476 5130 6546 5168
rect 6476 4998 6492 5130
rect 6530 4998 6546 5130
rect 6476 4988 6546 4998
rect 6716 5130 6786 5168
rect 6716 4998 6732 5130
rect 6770 4998 6786 5130
rect 6716 4988 6786 4998
rect 6956 5130 7026 5168
rect 6956 4998 6972 5130
rect 7010 4998 7026 5130
rect 6956 4988 7026 4998
rect 7196 5130 7266 5168
rect 7196 4998 7212 5130
rect 7250 4998 7266 5130
rect 7196 4988 7266 4998
rect 7436 5130 7506 5168
rect 7436 4998 7452 5130
rect 7490 4998 7506 5130
rect 7436 4988 7506 4998
rect 7676 5130 7746 5168
rect 7676 4998 7692 5130
rect 7730 4998 7746 5130
rect 7676 4988 7746 4998
rect 7916 5130 7986 5168
rect 7916 4998 7932 5130
rect 7970 4998 7986 5130
rect 7916 4988 7986 4998
rect 8156 5130 8226 5168
rect 8156 4998 8172 5130
rect 8210 4998 8226 5130
rect 8156 4988 8226 4998
rect 8396 5130 8466 5168
rect 8396 4998 8412 5130
rect 8450 4998 8466 5130
rect 8396 4988 8466 4998
rect 8636 5130 8706 5168
rect 8636 4998 8652 5130
rect 8690 4998 8706 5130
rect 8636 4988 8706 4998
rect 8876 5130 8946 5168
rect 8876 4998 8892 5130
rect 8930 4998 8946 5130
rect 8876 4988 8946 4998
rect 9116 5130 9186 5168
rect 9116 4998 9132 5130
rect 9170 4998 9186 5130
rect 9116 4988 9186 4998
rect 9356 5130 9426 5168
rect 9356 4998 9372 5130
rect 9410 4998 9426 5130
rect 9356 4988 9426 4998
rect 9596 5130 9666 5168
rect 9596 4998 9612 5130
rect 9650 4998 9666 5130
rect 9596 4988 9666 4998
rect 9836 5130 9906 5168
rect 9836 4998 9852 5130
rect 9890 4998 9906 5130
rect 9836 4988 9906 4998
rect 10076 5130 10146 5168
rect 10076 4998 10092 5130
rect 10130 4998 10146 5130
rect 10076 4988 10146 4998
rect 10316 5130 10386 5168
rect 10316 4998 10332 5130
rect 10370 4998 10386 5130
rect 10316 4988 10386 4998
rect 10556 5130 10626 5168
rect 10556 4998 10572 5130
rect 10610 4998 10626 5130
rect 10556 4988 10626 4998
rect 10796 5130 10866 5168
rect 10796 4998 10812 5130
rect 10850 4998 10866 5130
rect 10796 4988 10866 4998
rect 11036 5130 11106 5168
rect 11036 4998 11052 5130
rect 11090 4998 11106 5130
rect 11036 4988 11106 4998
rect 11276 5130 11346 5168
rect 11276 4998 11292 5130
rect 11330 4998 11346 5130
rect 11276 4988 11346 4998
rect 11516 5130 11586 5168
rect 11516 4998 11532 5130
rect 11570 4998 11586 5130
rect 11516 4988 11586 4998
rect 11756 5130 11826 5168
rect 11756 4998 11772 5130
rect 11810 4998 11826 5130
rect 11756 4988 11826 4998
rect 11996 5130 12066 5168
rect 11996 4998 12012 5130
rect 12050 4998 12066 5130
rect 11996 4988 12066 4998
rect 12236 5130 12306 5168
rect 12236 4998 12252 5130
rect 12290 4998 12306 5130
rect 12236 4988 12306 4998
rect -6428 2537 -6028 2553
rect -6428 2503 -6412 2537
rect -6044 2503 -6028 2537
rect -6428 2456 -6028 2503
rect -5840 2537 -5440 2553
rect -5840 2503 -5824 2537
rect -5456 2503 -5440 2537
rect -5840 2456 -5440 2503
rect -5252 2537 -4852 2553
rect -5252 2503 -5236 2537
rect -4868 2503 -4852 2537
rect -5252 2456 -4852 2503
rect -4664 2537 -4264 2553
rect -4664 2503 -4648 2537
rect -4280 2503 -4264 2537
rect -4664 2456 -4264 2503
rect -4076 2537 -3676 2553
rect -4076 2503 -4060 2537
rect -3692 2503 -3676 2537
rect -4076 2456 -3676 2503
rect -3488 2537 -3088 2553
rect -3488 2503 -3472 2537
rect -3104 2503 -3088 2537
rect -3488 2456 -3088 2503
rect -2900 2537 -2500 2553
rect -2900 2503 -2884 2537
rect -2516 2503 -2500 2537
rect -2900 2456 -2500 2503
rect -2312 2537 -1912 2553
rect -2312 2503 -2296 2537
rect -1928 2503 -1912 2537
rect -2312 2456 -1912 2503
rect -1724 2537 -1324 2553
rect -1724 2503 -1708 2537
rect -1340 2503 -1324 2537
rect -1724 2456 -1324 2503
rect -1136 2537 -736 2553
rect -1136 2503 -1120 2537
rect -752 2503 -736 2537
rect -1136 2456 -736 2503
rect -548 2537 -148 2553
rect -548 2503 -532 2537
rect -164 2503 -148 2537
rect -548 2456 -148 2503
rect 40 2537 440 2553
rect 40 2503 56 2537
rect 424 2503 440 2537
rect 40 2456 440 2503
rect 628 2537 1028 2553
rect 628 2503 644 2537
rect 1012 2503 1028 2537
rect 628 2456 1028 2503
rect 1216 2537 1616 2553
rect 1216 2503 1232 2537
rect 1600 2503 1616 2537
rect 1216 2456 1616 2503
rect 1804 2537 2204 2553
rect 1804 2503 1820 2537
rect 2188 2503 2204 2537
rect 1804 2456 2204 2503
rect 2392 2537 2792 2553
rect 2392 2503 2408 2537
rect 2776 2503 2792 2537
rect 2392 2456 2792 2503
rect 2980 2537 3380 2553
rect 2980 2503 2996 2537
rect 3364 2503 3380 2537
rect 2980 2456 3380 2503
rect 3568 2537 3968 2553
rect 3568 2503 3584 2537
rect 3952 2503 3968 2537
rect 3568 2456 3968 2503
rect 4156 2537 4556 2553
rect 4156 2503 4172 2537
rect 4540 2503 4556 2537
rect 4156 2456 4556 2503
rect 4744 2537 5144 2553
rect 4744 2503 4760 2537
rect 5128 2503 5144 2537
rect 4744 2456 5144 2503
rect 5332 2537 5732 2553
rect 5332 2503 5348 2537
rect 5716 2503 5732 2537
rect 5332 2456 5732 2503
rect 5920 2537 6320 2553
rect 5920 2503 5936 2537
rect 6304 2503 6320 2537
rect 5920 2456 6320 2503
rect 6508 2537 6908 2553
rect 6508 2503 6524 2537
rect 6892 2503 6908 2537
rect 6508 2456 6908 2503
rect 7096 2537 7496 2553
rect 7096 2503 7112 2537
rect 7480 2503 7496 2537
rect 7096 2456 7496 2503
rect 7684 2537 8084 2553
rect 7684 2503 7700 2537
rect 8068 2503 8084 2537
rect 7684 2456 8084 2503
rect 8272 2537 8672 2553
rect 8272 2503 8288 2537
rect 8656 2503 8672 2537
rect 8272 2456 8672 2503
rect 8860 2537 9260 2553
rect 8860 2503 8876 2537
rect 9244 2503 9260 2537
rect 8860 2456 9260 2503
rect 9448 2537 9848 2553
rect 9448 2503 9464 2537
rect 9832 2503 9848 2537
rect 9448 2456 9848 2503
rect 10036 2537 10436 2553
rect 10036 2503 10052 2537
rect 10420 2503 10436 2537
rect 10036 2456 10436 2503
rect 10624 2537 11024 2553
rect 10624 2503 10640 2537
rect 11008 2503 11024 2537
rect 10624 2456 11024 2503
rect 11212 2537 11612 2553
rect 11212 2503 11228 2537
rect 11596 2503 11612 2537
rect 11212 2456 11612 2503
rect 11800 2537 12200 2553
rect 11800 2503 11816 2537
rect 12184 2503 12200 2537
rect 11800 2456 12200 2503
rect 12388 2537 12788 2553
rect 12388 2503 12404 2537
rect 12772 2503 12788 2537
rect 12388 2456 12788 2503
rect 12976 2537 13376 2553
rect 12976 2503 12992 2537
rect 13360 2503 13376 2537
rect 12976 2456 13376 2503
rect 13564 2537 13964 2553
rect 13564 2503 13580 2537
rect 13948 2503 13964 2537
rect 13564 2456 13964 2503
rect 14152 2537 14552 2553
rect 14152 2503 14168 2537
rect 14536 2503 14552 2537
rect 14152 2456 14552 2503
rect 14740 2537 15140 2553
rect 14740 2503 14756 2537
rect 15124 2503 15140 2537
rect 14740 2456 15140 2503
rect 15328 2537 15728 2553
rect 15328 2503 15344 2537
rect 15712 2503 15728 2537
rect 15328 2456 15728 2503
rect 15916 2537 16316 2553
rect 15916 2503 15932 2537
rect 16300 2503 16316 2537
rect 15916 2456 16316 2503
rect 16504 2537 16904 2553
rect 16504 2503 16520 2537
rect 16888 2503 16904 2537
rect 16504 2456 16904 2503
rect 17092 2537 17492 2553
rect 17092 2503 17108 2537
rect 17476 2503 17492 2537
rect 17092 2456 17492 2503
rect 17680 2537 18080 2553
rect 17680 2503 17696 2537
rect 18064 2503 18080 2537
rect 17680 2456 18080 2503
rect 18268 2537 18668 2553
rect 18268 2503 18284 2537
rect 18652 2503 18668 2537
rect 18268 2456 18668 2503
rect 18856 2537 19256 2553
rect 18856 2503 18872 2537
rect 19240 2503 19256 2537
rect 18856 2456 19256 2503
rect 19444 2537 19844 2553
rect 19444 2503 19460 2537
rect 19828 2503 19844 2537
rect 19444 2456 19844 2503
rect 20032 2537 20432 2553
rect 20032 2503 20048 2537
rect 20416 2503 20432 2537
rect 20032 2456 20432 2503
rect 20620 2537 21020 2553
rect 20620 2503 20636 2537
rect 21004 2503 21020 2537
rect 20620 2456 21020 2503
rect 21208 2537 21608 2553
rect 21208 2503 21224 2537
rect 21592 2503 21608 2537
rect 21208 2456 21608 2503
rect -6428 1609 -6028 1656
rect -6428 1575 -6412 1609
rect -6044 1575 -6028 1609
rect -6428 1537 -6028 1575
rect -6428 1503 -6412 1537
rect -6044 1503 -6028 1537
rect -6428 1456 -6028 1503
rect -5840 1609 -5440 1656
rect -5840 1575 -5824 1609
rect -5456 1575 -5440 1609
rect -5840 1537 -5440 1575
rect -5840 1503 -5824 1537
rect -5456 1503 -5440 1537
rect -5840 1456 -5440 1503
rect -5252 1609 -4852 1656
rect -5252 1575 -5236 1609
rect -4868 1575 -4852 1609
rect -5252 1537 -4852 1575
rect -5252 1503 -5236 1537
rect -4868 1503 -4852 1537
rect -5252 1456 -4852 1503
rect -4664 1609 -4264 1656
rect -4664 1575 -4648 1609
rect -4280 1575 -4264 1609
rect -4664 1537 -4264 1575
rect -4664 1503 -4648 1537
rect -4280 1503 -4264 1537
rect -4664 1456 -4264 1503
rect -4076 1609 -3676 1656
rect -4076 1575 -4060 1609
rect -3692 1575 -3676 1609
rect -4076 1537 -3676 1575
rect -4076 1503 -4060 1537
rect -3692 1503 -3676 1537
rect -4076 1456 -3676 1503
rect -3488 1609 -3088 1656
rect -3488 1575 -3472 1609
rect -3104 1575 -3088 1609
rect -3488 1537 -3088 1575
rect -3488 1503 -3472 1537
rect -3104 1503 -3088 1537
rect -3488 1456 -3088 1503
rect -2900 1609 -2500 1656
rect -2900 1575 -2884 1609
rect -2516 1575 -2500 1609
rect -2900 1537 -2500 1575
rect -2900 1503 -2884 1537
rect -2516 1503 -2500 1537
rect -2900 1456 -2500 1503
rect -2312 1609 -1912 1656
rect -2312 1575 -2296 1609
rect -1928 1575 -1912 1609
rect -2312 1537 -1912 1575
rect -2312 1503 -2296 1537
rect -1928 1503 -1912 1537
rect -2312 1456 -1912 1503
rect -1724 1609 -1324 1656
rect -1724 1575 -1708 1609
rect -1340 1575 -1324 1609
rect -1724 1537 -1324 1575
rect -1724 1503 -1708 1537
rect -1340 1503 -1324 1537
rect -1724 1456 -1324 1503
rect -1136 1609 -736 1656
rect -1136 1575 -1120 1609
rect -752 1575 -736 1609
rect -1136 1537 -736 1575
rect -1136 1503 -1120 1537
rect -752 1503 -736 1537
rect -1136 1456 -736 1503
rect -548 1609 -148 1656
rect -548 1575 -532 1609
rect -164 1575 -148 1609
rect -548 1537 -148 1575
rect -548 1503 -532 1537
rect -164 1503 -148 1537
rect -548 1456 -148 1503
rect 40 1609 440 1656
rect 40 1575 56 1609
rect 424 1575 440 1609
rect 40 1537 440 1575
rect 40 1503 56 1537
rect 424 1503 440 1537
rect 40 1456 440 1503
rect 628 1609 1028 1656
rect 628 1575 644 1609
rect 1012 1575 1028 1609
rect 628 1537 1028 1575
rect 628 1503 644 1537
rect 1012 1503 1028 1537
rect 628 1456 1028 1503
rect 1216 1609 1616 1656
rect 1216 1575 1232 1609
rect 1600 1575 1616 1609
rect 1216 1537 1616 1575
rect 1216 1503 1232 1537
rect 1600 1503 1616 1537
rect 1216 1456 1616 1503
rect 1804 1609 2204 1656
rect 1804 1575 1820 1609
rect 2188 1575 2204 1609
rect 1804 1537 2204 1575
rect 1804 1503 1820 1537
rect 2188 1503 2204 1537
rect 1804 1456 2204 1503
rect 2392 1609 2792 1656
rect 2392 1575 2408 1609
rect 2776 1575 2792 1609
rect 2392 1537 2792 1575
rect 2392 1503 2408 1537
rect 2776 1503 2792 1537
rect 2392 1456 2792 1503
rect 2980 1609 3380 1656
rect 2980 1575 2996 1609
rect 3364 1575 3380 1609
rect 2980 1537 3380 1575
rect 2980 1503 2996 1537
rect 3364 1503 3380 1537
rect 2980 1456 3380 1503
rect 3568 1609 3968 1656
rect 3568 1575 3584 1609
rect 3952 1575 3968 1609
rect 3568 1537 3968 1575
rect 3568 1503 3584 1537
rect 3952 1503 3968 1537
rect 3568 1456 3968 1503
rect 4156 1609 4556 1656
rect 4156 1575 4172 1609
rect 4540 1575 4556 1609
rect 4156 1537 4556 1575
rect 4156 1503 4172 1537
rect 4540 1503 4556 1537
rect 4156 1456 4556 1503
rect 4744 1609 5144 1656
rect 4744 1575 4760 1609
rect 5128 1575 5144 1609
rect 4744 1537 5144 1575
rect 4744 1503 4760 1537
rect 5128 1503 5144 1537
rect 4744 1456 5144 1503
rect 5332 1609 5732 1656
rect 5332 1575 5348 1609
rect 5716 1575 5732 1609
rect 5332 1537 5732 1575
rect 5332 1503 5348 1537
rect 5716 1503 5732 1537
rect 5332 1456 5732 1503
rect 5920 1609 6320 1656
rect 5920 1575 5936 1609
rect 6304 1575 6320 1609
rect 5920 1537 6320 1575
rect 5920 1503 5936 1537
rect 6304 1503 6320 1537
rect 5920 1456 6320 1503
rect 6508 1609 6908 1656
rect 6508 1575 6524 1609
rect 6892 1575 6908 1609
rect 6508 1537 6908 1575
rect 6508 1503 6524 1537
rect 6892 1503 6908 1537
rect 6508 1456 6908 1503
rect 7096 1609 7496 1656
rect 7096 1575 7112 1609
rect 7480 1575 7496 1609
rect 7096 1537 7496 1575
rect 7096 1503 7112 1537
rect 7480 1503 7496 1537
rect 7096 1456 7496 1503
rect 7684 1609 8084 1656
rect 7684 1575 7700 1609
rect 8068 1575 8084 1609
rect 7684 1537 8084 1575
rect 7684 1503 7700 1537
rect 8068 1503 8084 1537
rect 7684 1456 8084 1503
rect 8272 1609 8672 1656
rect 8272 1575 8288 1609
rect 8656 1575 8672 1609
rect 8272 1537 8672 1575
rect 8272 1503 8288 1537
rect 8656 1503 8672 1537
rect 8272 1456 8672 1503
rect 8860 1609 9260 1656
rect 8860 1575 8876 1609
rect 9244 1575 9260 1609
rect 8860 1537 9260 1575
rect 8860 1503 8876 1537
rect 9244 1503 9260 1537
rect 8860 1456 9260 1503
rect 9448 1609 9848 1656
rect 9448 1575 9464 1609
rect 9832 1575 9848 1609
rect 9448 1537 9848 1575
rect 9448 1503 9464 1537
rect 9832 1503 9848 1537
rect 9448 1456 9848 1503
rect 10036 1609 10436 1656
rect 10036 1575 10052 1609
rect 10420 1575 10436 1609
rect 10036 1537 10436 1575
rect 10036 1503 10052 1537
rect 10420 1503 10436 1537
rect 10036 1456 10436 1503
rect 10624 1609 11024 1656
rect 10624 1575 10640 1609
rect 11008 1575 11024 1609
rect 10624 1537 11024 1575
rect 10624 1503 10640 1537
rect 11008 1503 11024 1537
rect 10624 1456 11024 1503
rect 11212 1609 11612 1656
rect 11212 1575 11228 1609
rect 11596 1575 11612 1609
rect 11212 1537 11612 1575
rect 11212 1503 11228 1537
rect 11596 1503 11612 1537
rect 11212 1456 11612 1503
rect 11800 1609 12200 1656
rect 11800 1575 11816 1609
rect 12184 1575 12200 1609
rect 11800 1537 12200 1575
rect 11800 1503 11816 1537
rect 12184 1503 12200 1537
rect 11800 1456 12200 1503
rect 12388 1609 12788 1656
rect 12388 1575 12404 1609
rect 12772 1575 12788 1609
rect 12388 1537 12788 1575
rect 12388 1503 12404 1537
rect 12772 1503 12788 1537
rect 12388 1456 12788 1503
rect 12976 1609 13376 1656
rect 12976 1575 12992 1609
rect 13360 1575 13376 1609
rect 12976 1537 13376 1575
rect 12976 1503 12992 1537
rect 13360 1503 13376 1537
rect 12976 1456 13376 1503
rect 13564 1609 13964 1656
rect 13564 1575 13580 1609
rect 13948 1575 13964 1609
rect 13564 1537 13964 1575
rect 13564 1503 13580 1537
rect 13948 1503 13964 1537
rect 13564 1456 13964 1503
rect 14152 1609 14552 1656
rect 14152 1575 14168 1609
rect 14536 1575 14552 1609
rect 14152 1537 14552 1575
rect 14152 1503 14168 1537
rect 14536 1503 14552 1537
rect 14152 1456 14552 1503
rect 14740 1609 15140 1656
rect 14740 1575 14756 1609
rect 15124 1575 15140 1609
rect 14740 1537 15140 1575
rect 14740 1503 14756 1537
rect 15124 1503 15140 1537
rect 14740 1456 15140 1503
rect 15328 1609 15728 1656
rect 15328 1575 15344 1609
rect 15712 1575 15728 1609
rect 15328 1537 15728 1575
rect 15328 1503 15344 1537
rect 15712 1503 15728 1537
rect 15328 1456 15728 1503
rect 15916 1609 16316 1656
rect 15916 1575 15932 1609
rect 16300 1575 16316 1609
rect 15916 1537 16316 1575
rect 15916 1503 15932 1537
rect 16300 1503 16316 1537
rect 15916 1456 16316 1503
rect 16504 1609 16904 1656
rect 16504 1575 16520 1609
rect 16888 1575 16904 1609
rect 16504 1537 16904 1575
rect 16504 1503 16520 1537
rect 16888 1503 16904 1537
rect 16504 1456 16904 1503
rect 17092 1609 17492 1656
rect 17092 1575 17108 1609
rect 17476 1575 17492 1609
rect 17092 1537 17492 1575
rect 17092 1503 17108 1537
rect 17476 1503 17492 1537
rect 17092 1456 17492 1503
rect 17680 1609 18080 1656
rect 17680 1575 17696 1609
rect 18064 1575 18080 1609
rect 17680 1537 18080 1575
rect 17680 1503 17696 1537
rect 18064 1503 18080 1537
rect 17680 1456 18080 1503
rect 18268 1609 18668 1656
rect 18268 1575 18284 1609
rect 18652 1575 18668 1609
rect 18268 1537 18668 1575
rect 18268 1503 18284 1537
rect 18652 1503 18668 1537
rect 18268 1456 18668 1503
rect 18856 1609 19256 1656
rect 18856 1575 18872 1609
rect 19240 1575 19256 1609
rect 18856 1537 19256 1575
rect 18856 1503 18872 1537
rect 19240 1503 19256 1537
rect 18856 1456 19256 1503
rect 19444 1609 19844 1656
rect 19444 1575 19460 1609
rect 19828 1575 19844 1609
rect 19444 1537 19844 1575
rect 19444 1503 19460 1537
rect 19828 1503 19844 1537
rect 19444 1456 19844 1503
rect 20032 1609 20432 1656
rect 20032 1575 20048 1609
rect 20416 1575 20432 1609
rect 20032 1537 20432 1575
rect 20032 1503 20048 1537
rect 20416 1503 20432 1537
rect 20032 1456 20432 1503
rect 20620 1609 21020 1656
rect 20620 1575 20636 1609
rect 21004 1575 21020 1609
rect 20620 1537 21020 1575
rect 20620 1503 20636 1537
rect 21004 1503 21020 1537
rect 20620 1456 21020 1503
rect 21208 1609 21608 1656
rect 21208 1575 21224 1609
rect 21592 1575 21608 1609
rect 21208 1537 21608 1575
rect 21208 1503 21224 1537
rect 21592 1503 21608 1537
rect 21208 1456 21608 1503
rect -6428 609 -6028 656
rect -6428 575 -6412 609
rect -6044 575 -6028 609
rect -6428 537 -6028 575
rect -6428 503 -6412 537
rect -6044 503 -6028 537
rect -6428 456 -6028 503
rect -5840 609 -5440 656
rect -5840 575 -5824 609
rect -5456 575 -5440 609
rect -5840 537 -5440 575
rect -5840 503 -5824 537
rect -5456 503 -5440 537
rect -5840 456 -5440 503
rect -5252 609 -4852 656
rect -5252 575 -5236 609
rect -4868 575 -4852 609
rect -5252 537 -4852 575
rect -5252 503 -5236 537
rect -4868 503 -4852 537
rect -5252 456 -4852 503
rect -4664 609 -4264 656
rect -4664 575 -4648 609
rect -4280 575 -4264 609
rect -4664 537 -4264 575
rect -4664 503 -4648 537
rect -4280 503 -4264 537
rect -4664 456 -4264 503
rect -4076 609 -3676 656
rect -4076 575 -4060 609
rect -3692 575 -3676 609
rect -4076 537 -3676 575
rect -4076 503 -4060 537
rect -3692 503 -3676 537
rect -4076 456 -3676 503
rect -3488 609 -3088 656
rect -3488 575 -3472 609
rect -3104 575 -3088 609
rect -3488 537 -3088 575
rect -3488 503 -3472 537
rect -3104 503 -3088 537
rect -3488 456 -3088 503
rect -2900 609 -2500 656
rect -2900 575 -2884 609
rect -2516 575 -2500 609
rect -2900 537 -2500 575
rect -2900 503 -2884 537
rect -2516 503 -2500 537
rect -2900 456 -2500 503
rect -2312 609 -1912 656
rect -2312 575 -2296 609
rect -1928 575 -1912 609
rect -2312 537 -1912 575
rect -2312 503 -2296 537
rect -1928 503 -1912 537
rect -2312 456 -1912 503
rect -1724 609 -1324 656
rect -1724 575 -1708 609
rect -1340 575 -1324 609
rect -1724 537 -1324 575
rect -1724 503 -1708 537
rect -1340 503 -1324 537
rect -1724 456 -1324 503
rect -1136 609 -736 656
rect -1136 575 -1120 609
rect -752 575 -736 609
rect -1136 537 -736 575
rect -1136 503 -1120 537
rect -752 503 -736 537
rect -1136 456 -736 503
rect -548 609 -148 656
rect -548 575 -532 609
rect -164 575 -148 609
rect -548 537 -148 575
rect -548 503 -532 537
rect -164 503 -148 537
rect -548 456 -148 503
rect 40 609 440 656
rect 40 575 56 609
rect 424 575 440 609
rect 40 537 440 575
rect 40 503 56 537
rect 424 503 440 537
rect 40 456 440 503
rect 628 609 1028 656
rect 628 575 644 609
rect 1012 575 1028 609
rect 628 537 1028 575
rect 628 503 644 537
rect 1012 503 1028 537
rect 628 456 1028 503
rect 1216 609 1616 656
rect 1216 575 1232 609
rect 1600 575 1616 609
rect 1216 537 1616 575
rect 1216 503 1232 537
rect 1600 503 1616 537
rect 1216 456 1616 503
rect 1804 609 2204 656
rect 1804 575 1820 609
rect 2188 575 2204 609
rect 1804 537 2204 575
rect 1804 503 1820 537
rect 2188 503 2204 537
rect 1804 456 2204 503
rect 2392 609 2792 656
rect 2392 575 2408 609
rect 2776 575 2792 609
rect 2392 537 2792 575
rect 2392 503 2408 537
rect 2776 503 2792 537
rect 2392 456 2792 503
rect 2980 609 3380 656
rect 2980 575 2996 609
rect 3364 575 3380 609
rect 2980 537 3380 575
rect 2980 503 2996 537
rect 3364 503 3380 537
rect 2980 456 3380 503
rect 3568 609 3968 656
rect 3568 575 3584 609
rect 3952 575 3968 609
rect 3568 537 3968 575
rect 3568 503 3584 537
rect 3952 503 3968 537
rect 3568 456 3968 503
rect 4156 609 4556 656
rect 4156 575 4172 609
rect 4540 575 4556 609
rect 4156 537 4556 575
rect 4156 503 4172 537
rect 4540 503 4556 537
rect 4156 456 4556 503
rect 4744 609 5144 656
rect 4744 575 4760 609
rect 5128 575 5144 609
rect 4744 537 5144 575
rect 4744 503 4760 537
rect 5128 503 5144 537
rect 4744 456 5144 503
rect 5332 609 5732 656
rect 5332 575 5348 609
rect 5716 575 5732 609
rect 5332 537 5732 575
rect 5332 503 5348 537
rect 5716 503 5732 537
rect 5332 456 5732 503
rect 5920 609 6320 656
rect 5920 575 5936 609
rect 6304 575 6320 609
rect 5920 537 6320 575
rect 5920 503 5936 537
rect 6304 503 6320 537
rect 5920 456 6320 503
rect 6508 609 6908 656
rect 6508 575 6524 609
rect 6892 575 6908 609
rect 6508 537 6908 575
rect 6508 503 6524 537
rect 6892 503 6908 537
rect 6508 456 6908 503
rect 7096 609 7496 656
rect 7096 575 7112 609
rect 7480 575 7496 609
rect 7096 537 7496 575
rect 7096 503 7112 537
rect 7480 503 7496 537
rect 7096 456 7496 503
rect 7684 609 8084 656
rect 7684 575 7700 609
rect 8068 575 8084 609
rect 7684 537 8084 575
rect 7684 503 7700 537
rect 8068 503 8084 537
rect 7684 456 8084 503
rect 8272 609 8672 656
rect 8272 575 8288 609
rect 8656 575 8672 609
rect 8272 537 8672 575
rect 8272 503 8288 537
rect 8656 503 8672 537
rect 8272 456 8672 503
rect 8860 609 9260 656
rect 8860 575 8876 609
rect 9244 575 9260 609
rect 8860 537 9260 575
rect 8860 503 8876 537
rect 9244 503 9260 537
rect 8860 456 9260 503
rect 9448 609 9848 656
rect 9448 575 9464 609
rect 9832 575 9848 609
rect 9448 537 9848 575
rect 9448 503 9464 537
rect 9832 503 9848 537
rect 9448 456 9848 503
rect 10036 609 10436 656
rect 10036 575 10052 609
rect 10420 575 10436 609
rect 10036 537 10436 575
rect 10036 503 10052 537
rect 10420 503 10436 537
rect 10036 456 10436 503
rect 10624 609 11024 656
rect 10624 575 10640 609
rect 11008 575 11024 609
rect 10624 537 11024 575
rect 10624 503 10640 537
rect 11008 503 11024 537
rect 10624 456 11024 503
rect 11212 609 11612 656
rect 11212 575 11228 609
rect 11596 575 11612 609
rect 11212 537 11612 575
rect 11212 503 11228 537
rect 11596 503 11612 537
rect 11212 456 11612 503
rect 11800 609 12200 656
rect 11800 575 11816 609
rect 12184 575 12200 609
rect 11800 537 12200 575
rect 11800 503 11816 537
rect 12184 503 12200 537
rect 11800 456 12200 503
rect 12388 609 12788 656
rect 12388 575 12404 609
rect 12772 575 12788 609
rect 12388 537 12788 575
rect 12388 503 12404 537
rect 12772 503 12788 537
rect 12388 456 12788 503
rect 12976 609 13376 656
rect 12976 575 12992 609
rect 13360 575 13376 609
rect 12976 537 13376 575
rect 12976 503 12992 537
rect 13360 503 13376 537
rect 12976 456 13376 503
rect 13564 609 13964 656
rect 13564 575 13580 609
rect 13948 575 13964 609
rect 13564 537 13964 575
rect 13564 503 13580 537
rect 13948 503 13964 537
rect 13564 456 13964 503
rect 14152 609 14552 656
rect 14152 575 14168 609
rect 14536 575 14552 609
rect 14152 537 14552 575
rect 14152 503 14168 537
rect 14536 503 14552 537
rect 14152 456 14552 503
rect 14740 609 15140 656
rect 14740 575 14756 609
rect 15124 575 15140 609
rect 14740 537 15140 575
rect 14740 503 14756 537
rect 15124 503 15140 537
rect 14740 456 15140 503
rect 15328 609 15728 656
rect 15328 575 15344 609
rect 15712 575 15728 609
rect 15328 537 15728 575
rect 15328 503 15344 537
rect 15712 503 15728 537
rect 15328 456 15728 503
rect 15916 609 16316 656
rect 15916 575 15932 609
rect 16300 575 16316 609
rect 15916 537 16316 575
rect 15916 503 15932 537
rect 16300 503 16316 537
rect 15916 456 16316 503
rect 16504 609 16904 656
rect 16504 575 16520 609
rect 16888 575 16904 609
rect 16504 537 16904 575
rect 16504 503 16520 537
rect 16888 503 16904 537
rect 16504 456 16904 503
rect 17092 609 17492 656
rect 17092 575 17108 609
rect 17476 575 17492 609
rect 17092 537 17492 575
rect 17092 503 17108 537
rect 17476 503 17492 537
rect 17092 456 17492 503
rect 17680 609 18080 656
rect 17680 575 17696 609
rect 18064 575 18080 609
rect 17680 537 18080 575
rect 17680 503 17696 537
rect 18064 503 18080 537
rect 17680 456 18080 503
rect 18268 609 18668 656
rect 18268 575 18284 609
rect 18652 575 18668 609
rect 18268 537 18668 575
rect 18268 503 18284 537
rect 18652 503 18668 537
rect 18268 456 18668 503
rect 18856 609 19256 656
rect 18856 575 18872 609
rect 19240 575 19256 609
rect 18856 537 19256 575
rect 18856 503 18872 537
rect 19240 503 19256 537
rect 18856 456 19256 503
rect 19444 609 19844 656
rect 19444 575 19460 609
rect 19828 575 19844 609
rect 19444 537 19844 575
rect 19444 503 19460 537
rect 19828 503 19844 537
rect 19444 456 19844 503
rect 20032 609 20432 656
rect 20032 575 20048 609
rect 20416 575 20432 609
rect 20032 537 20432 575
rect 20032 503 20048 537
rect 20416 503 20432 537
rect 20032 456 20432 503
rect 20620 609 21020 656
rect 20620 575 20636 609
rect 21004 575 21020 609
rect 20620 537 21020 575
rect 20620 503 20636 537
rect 21004 503 21020 537
rect 20620 456 21020 503
rect 21208 609 21608 656
rect 21208 575 21224 609
rect 21592 575 21608 609
rect 21208 537 21608 575
rect 21208 503 21224 537
rect 21592 503 21608 537
rect 21208 456 21608 503
rect -6428 -391 -6028 -344
rect -6428 -425 -6412 -391
rect -6044 -425 -6028 -391
rect -6428 -441 -6028 -425
rect -5840 -391 -5440 -344
rect -5840 -425 -5824 -391
rect -5456 -425 -5440 -391
rect -5840 -441 -5440 -425
rect -5252 -391 -4852 -344
rect -5252 -425 -5236 -391
rect -4868 -425 -4852 -391
rect -5252 -441 -4852 -425
rect -4664 -391 -4264 -344
rect -4664 -425 -4648 -391
rect -4280 -425 -4264 -391
rect -4664 -441 -4264 -425
rect -4076 -391 -3676 -344
rect -4076 -425 -4060 -391
rect -3692 -425 -3676 -391
rect -4076 -441 -3676 -425
rect -3488 -391 -3088 -344
rect -3488 -425 -3472 -391
rect -3104 -425 -3088 -391
rect -3488 -441 -3088 -425
rect -2900 -391 -2500 -344
rect -2900 -425 -2884 -391
rect -2516 -425 -2500 -391
rect -2900 -441 -2500 -425
rect -2312 -391 -1912 -344
rect -2312 -425 -2296 -391
rect -1928 -425 -1912 -391
rect -2312 -441 -1912 -425
rect -1724 -391 -1324 -344
rect -1724 -425 -1708 -391
rect -1340 -425 -1324 -391
rect -1724 -441 -1324 -425
rect -1136 -391 -736 -344
rect -1136 -425 -1120 -391
rect -752 -425 -736 -391
rect -1136 -441 -736 -425
rect -548 -391 -148 -344
rect -548 -425 -532 -391
rect -164 -425 -148 -391
rect -548 -441 -148 -425
rect 40 -391 440 -344
rect 40 -425 56 -391
rect 424 -425 440 -391
rect 40 -441 440 -425
rect 628 -391 1028 -344
rect 628 -425 644 -391
rect 1012 -425 1028 -391
rect 628 -441 1028 -425
rect 1216 -391 1616 -344
rect 1216 -425 1232 -391
rect 1600 -425 1616 -391
rect 1216 -441 1616 -425
rect 1804 -391 2204 -344
rect 1804 -425 1820 -391
rect 2188 -425 2204 -391
rect 1804 -441 2204 -425
rect 2392 -391 2792 -344
rect 2392 -425 2408 -391
rect 2776 -425 2792 -391
rect 2392 -441 2792 -425
rect 2980 -391 3380 -344
rect 2980 -425 2996 -391
rect 3364 -425 3380 -391
rect 2980 -441 3380 -425
rect 3568 -391 3968 -344
rect 3568 -425 3584 -391
rect 3952 -425 3968 -391
rect 3568 -441 3968 -425
rect 4156 -391 4556 -344
rect 4156 -425 4172 -391
rect 4540 -425 4556 -391
rect 4156 -441 4556 -425
rect 4744 -391 5144 -344
rect 4744 -425 4760 -391
rect 5128 -425 5144 -391
rect 4744 -441 5144 -425
rect 5332 -391 5732 -344
rect 5332 -425 5348 -391
rect 5716 -425 5732 -391
rect 5332 -441 5732 -425
rect 5920 -391 6320 -344
rect 5920 -425 5936 -391
rect 6304 -425 6320 -391
rect 5920 -441 6320 -425
rect 6508 -391 6908 -344
rect 6508 -425 6524 -391
rect 6892 -425 6908 -391
rect 6508 -441 6908 -425
rect 7096 -391 7496 -344
rect 7096 -425 7112 -391
rect 7480 -425 7496 -391
rect 7096 -441 7496 -425
rect 7684 -391 8084 -344
rect 7684 -425 7700 -391
rect 8068 -425 8084 -391
rect 7684 -441 8084 -425
rect 8272 -391 8672 -344
rect 8272 -425 8288 -391
rect 8656 -425 8672 -391
rect 8272 -441 8672 -425
rect 8860 -391 9260 -344
rect 8860 -425 8876 -391
rect 9244 -425 9260 -391
rect 8860 -441 9260 -425
rect 9448 -391 9848 -344
rect 9448 -425 9464 -391
rect 9832 -425 9848 -391
rect 9448 -441 9848 -425
rect 10036 -391 10436 -344
rect 10036 -425 10052 -391
rect 10420 -425 10436 -391
rect 10036 -441 10436 -425
rect 10624 -391 11024 -344
rect 10624 -425 10640 -391
rect 11008 -425 11024 -391
rect 10624 -441 11024 -425
rect 11212 -391 11612 -344
rect 11212 -425 11228 -391
rect 11596 -425 11612 -391
rect 11212 -441 11612 -425
rect 11800 -391 12200 -344
rect 11800 -425 11816 -391
rect 12184 -425 12200 -391
rect 11800 -441 12200 -425
rect 12388 -391 12788 -344
rect 12388 -425 12404 -391
rect 12772 -425 12788 -391
rect 12388 -441 12788 -425
rect 12976 -391 13376 -344
rect 12976 -425 12992 -391
rect 13360 -425 13376 -391
rect 12976 -441 13376 -425
rect 13564 -391 13964 -344
rect 13564 -425 13580 -391
rect 13948 -425 13964 -391
rect 13564 -441 13964 -425
rect 14152 -391 14552 -344
rect 14152 -425 14168 -391
rect 14536 -425 14552 -391
rect 14152 -441 14552 -425
rect 14740 -391 15140 -344
rect 14740 -425 14756 -391
rect 15124 -425 15140 -391
rect 14740 -441 15140 -425
rect 15328 -391 15728 -344
rect 15328 -425 15344 -391
rect 15712 -425 15728 -391
rect 15328 -441 15728 -425
rect 15916 -391 16316 -344
rect 15916 -425 15932 -391
rect 16300 -425 16316 -391
rect 15916 -441 16316 -425
rect 16504 -391 16904 -344
rect 16504 -425 16520 -391
rect 16888 -425 16904 -391
rect 16504 -441 16904 -425
rect 17092 -391 17492 -344
rect 17092 -425 17108 -391
rect 17476 -425 17492 -391
rect 17092 -441 17492 -425
rect 17680 -391 18080 -344
rect 17680 -425 17696 -391
rect 18064 -425 18080 -391
rect 17680 -441 18080 -425
rect 18268 -391 18668 -344
rect 18268 -425 18284 -391
rect 18652 -425 18668 -391
rect 18268 -441 18668 -425
rect 18856 -391 19256 -344
rect 18856 -425 18872 -391
rect 19240 -425 19256 -391
rect 18856 -441 19256 -425
rect 19444 -391 19844 -344
rect 19444 -425 19460 -391
rect 19828 -425 19844 -391
rect 19444 -441 19844 -425
rect 20032 -391 20432 -344
rect 20032 -425 20048 -391
rect 20416 -425 20432 -391
rect 20032 -441 20432 -425
rect 20620 -391 21020 -344
rect 20620 -425 20636 -391
rect 21004 -425 21020 -391
rect 20620 -441 21020 -425
rect 21208 -391 21608 -344
rect 21208 -425 21224 -391
rect 21592 -425 21608 -391
rect 21208 -441 21608 -425
rect 6624 -1820 6694 -1814
rect 6624 -1952 6640 -1820
rect 6678 -1952 6694 -1820
rect 6624 -1990 6694 -1952
rect 6890 -1820 6960 -1814
rect 6890 -1952 6906 -1820
rect 6944 -1952 6960 -1820
rect 6890 -1990 6960 -1952
rect 7156 -1820 7226 -1814
rect 7156 -1952 7172 -1820
rect 7210 -1952 7226 -1820
rect 7156 -1990 7226 -1952
rect 7422 -1820 7492 -1814
rect 7422 -1952 7438 -1820
rect 7476 -1952 7492 -1820
rect 7422 -1990 7492 -1952
rect 7688 -1820 7758 -1814
rect 7688 -1952 7704 -1820
rect 7742 -1952 7758 -1820
rect 7688 -1990 7758 -1952
rect 7954 -1820 8024 -1814
rect 7954 -1952 7970 -1820
rect 8008 -1952 8024 -1820
rect 7954 -1990 8024 -1952
rect 8220 -1820 8290 -1814
rect 8220 -1952 8236 -1820
rect 8274 -1952 8290 -1820
rect 8220 -1990 8290 -1952
rect 8486 -1820 8556 -1814
rect 8486 -1952 8502 -1820
rect 8540 -1952 8556 -1820
rect 8486 -1990 8556 -1952
rect 6624 -2830 6694 -2790
rect 6624 -2962 6640 -2830
rect 6678 -2962 6694 -2830
rect 6624 -3000 6694 -2962
rect 6890 -2830 6960 -2790
rect 6890 -2962 6906 -2830
rect 6944 -2962 6960 -2830
rect 6890 -3000 6960 -2962
rect 7156 -2830 7226 -2790
rect 7156 -2962 7172 -2830
rect 7210 -2962 7226 -2830
rect 7156 -3000 7226 -2962
rect 7422 -2830 7492 -2790
rect 7422 -2962 7438 -2830
rect 7476 -2962 7492 -2830
rect 7422 -3000 7492 -2962
rect 7688 -2830 7758 -2790
rect 7688 -2962 7704 -2830
rect 7742 -2962 7758 -2830
rect 7688 -3000 7758 -2962
rect 7954 -2830 8024 -2790
rect 7954 -2962 7970 -2830
rect 8008 -2962 8024 -2830
rect 7954 -3000 8024 -2962
rect 8220 -2830 8290 -2790
rect 8220 -2962 8236 -2830
rect 8274 -2962 8290 -2830
rect 8220 -3000 8290 -2962
rect 8486 -2830 8556 -2790
rect 8486 -2962 8502 -2830
rect 8540 -2962 8556 -2830
rect 8486 -3000 8556 -2962
rect 6624 -3840 6694 -3800
rect 6624 -3972 6640 -3840
rect 6678 -3972 6694 -3840
rect 6624 -4010 6694 -3972
rect 6890 -3840 6960 -3800
rect 6890 -3972 6906 -3840
rect 6944 -3972 6960 -3840
rect 6890 -4010 6960 -3972
rect 7156 -3840 7226 -3800
rect 7156 -3972 7172 -3840
rect 7210 -3972 7226 -3840
rect 7156 -4010 7226 -3972
rect 7422 -3840 7492 -3800
rect 7422 -3972 7438 -3840
rect 7476 -3972 7492 -3840
rect 7422 -4010 7492 -3972
rect 7688 -3840 7758 -3800
rect 7688 -3972 7704 -3840
rect 7742 -3972 7758 -3840
rect 7688 -4010 7758 -3972
rect 7954 -3840 8024 -3800
rect 7954 -3972 7970 -3840
rect 8008 -3972 8024 -3840
rect 7954 -4010 8024 -3972
rect 8220 -3840 8290 -3800
rect 8220 -3972 8236 -3840
rect 8274 -3972 8290 -3840
rect 8220 -4010 8290 -3972
rect 8486 -3840 8556 -3800
rect 8486 -3972 8502 -3840
rect 8540 -3972 8556 -3840
rect 8486 -4010 8556 -3972
rect 6624 -4850 6694 -4810
rect 6624 -4982 6640 -4850
rect 6678 -4982 6694 -4850
rect 6624 -4992 6694 -4982
rect 6890 -4850 6960 -4810
rect 6890 -4982 6906 -4850
rect 6944 -4982 6960 -4850
rect 6890 -4992 6960 -4982
rect 7156 -4850 7226 -4810
rect 7156 -4982 7172 -4850
rect 7210 -4982 7226 -4850
rect 7156 -4992 7226 -4982
rect 7422 -4850 7492 -4810
rect 7422 -4982 7438 -4850
rect 7476 -4982 7492 -4850
rect 7422 -4992 7492 -4982
rect 7688 -4850 7758 -4810
rect 7688 -4982 7704 -4850
rect 7742 -4982 7758 -4850
rect 7688 -4992 7758 -4982
rect 7954 -4850 8024 -4810
rect 7954 -4982 7970 -4850
rect 8008 -4982 8024 -4850
rect 7954 -4992 8024 -4982
rect 8220 -4850 8290 -4810
rect 8220 -4982 8236 -4850
rect 8274 -4982 8290 -4850
rect 8220 -4992 8290 -4982
rect 8486 -4850 8556 -4810
rect 8486 -4982 8502 -4850
rect 8540 -4982 8556 -4850
rect 8486 -4992 8556 -4982
rect 7196 -6018 7266 -6012
rect 7196 -6144 7212 -6018
rect 7250 -6144 7266 -6018
rect 7196 -6182 7266 -6144
rect 7436 -6018 7506 -6012
rect 7436 -6144 7452 -6018
rect 7490 -6144 7506 -6018
rect 7436 -6182 7506 -6144
rect 7676 -6018 7746 -6012
rect 7676 -6144 7692 -6018
rect 7730 -6144 7746 -6018
rect 7676 -6182 7746 -6144
rect 7916 -6018 7986 -6012
rect 7916 -6144 7932 -6018
rect 7970 -6144 7986 -6018
rect 7916 -6182 7986 -6144
rect 7196 -6820 7266 -6782
rect 7196 -6952 7212 -6820
rect 7250 -6952 7266 -6820
rect 7196 -6990 7266 -6952
rect 7436 -6820 7506 -6782
rect 7436 -6952 7452 -6820
rect 7490 -6952 7506 -6820
rect 7436 -6990 7506 -6952
rect 7676 -6820 7746 -6782
rect 7676 -6952 7692 -6820
rect 7730 -6952 7746 -6820
rect 7676 -6990 7746 -6952
rect 7916 -6820 7986 -6782
rect 7916 -6952 7932 -6820
rect 7970 -6952 7986 -6820
rect 7916 -6990 7986 -6952
rect 7196 -7628 7266 -7590
rect 7196 -7760 7212 -7628
rect 7250 -7760 7266 -7628
rect 7436 -7628 7506 -7590
rect 7436 -7760 7452 -7628
rect 7490 -7760 7506 -7628
rect 7676 -7628 7746 -7590
rect 7676 -7760 7692 -7628
rect 7730 -7760 7746 -7628
rect 7916 -7628 7986 -7590
rect 7916 -7760 7932 -7628
rect 7970 -7760 7986 -7628
<< polycont >>
rect 2892 6614 2930 6746
rect 3132 6614 3170 6746
rect 3372 6614 3410 6746
rect 3612 6614 3650 6746
rect 3852 6614 3890 6746
rect 4092 6614 4130 6746
rect 4332 6614 4370 6746
rect 4572 6614 4610 6746
rect 4812 6614 4850 6746
rect 5052 6614 5090 6746
rect 5292 6614 5330 6746
rect 5532 6614 5570 6746
rect 5772 6614 5810 6746
rect 6012 6614 6050 6746
rect 6252 6614 6290 6746
rect 6492 6614 6530 6746
rect 6732 6614 6770 6746
rect 6972 6614 7010 6746
rect 7212 6614 7250 6746
rect 7452 6614 7490 6746
rect 7692 6614 7730 6746
rect 7932 6614 7970 6746
rect 8172 6614 8210 6746
rect 8412 6614 8450 6746
rect 8652 6614 8690 6746
rect 8892 6614 8930 6746
rect 9132 6614 9170 6746
rect 9372 6614 9410 6746
rect 9612 6614 9650 6746
rect 9852 6614 9890 6746
rect 10092 6614 10130 6746
rect 10332 6614 10370 6746
rect 10572 6614 10610 6746
rect 10812 6614 10850 6746
rect 11052 6614 11090 6746
rect 11292 6614 11330 6746
rect 11532 6614 11570 6746
rect 11772 6614 11810 6746
rect 12012 6614 12050 6746
rect 12252 6614 12290 6746
rect 2892 5806 2930 5938
rect 3132 5806 3170 5938
rect 3372 5806 3410 5938
rect 3612 5806 3650 5938
rect 3852 5806 3890 5938
rect 4092 5806 4130 5938
rect 4332 5806 4370 5938
rect 4572 5806 4610 5938
rect 4812 5806 4850 5938
rect 5052 5806 5090 5938
rect 5292 5806 5330 5938
rect 5532 5806 5570 5938
rect 5772 5806 5810 5938
rect 6012 5806 6050 5938
rect 6252 5806 6290 5938
rect 6492 5806 6530 5938
rect 6732 5806 6770 5938
rect 6972 5806 7010 5938
rect 7212 5806 7250 5938
rect 7452 5806 7490 5938
rect 7692 5806 7730 5938
rect 7932 5806 7970 5938
rect 8172 5806 8210 5938
rect 8412 5806 8450 5938
rect 8652 5806 8690 5938
rect 8892 5806 8930 5938
rect 9132 5806 9170 5938
rect 9372 5806 9410 5938
rect 9612 5806 9650 5938
rect 9852 5806 9890 5938
rect 10092 5806 10130 5938
rect 10332 5806 10370 5938
rect 10572 5806 10610 5938
rect 10812 5806 10850 5938
rect 11052 5806 11090 5938
rect 11292 5806 11330 5938
rect 11532 5806 11570 5938
rect 11772 5806 11810 5938
rect 12012 5806 12050 5938
rect 12252 5806 12290 5938
rect 2892 4998 2930 5130
rect 3132 4998 3170 5130
rect 3372 4998 3410 5130
rect 3612 4998 3650 5130
rect 3852 4998 3890 5130
rect 4092 4998 4130 5130
rect 4332 4998 4370 5130
rect 4572 4998 4610 5130
rect 4812 4998 4850 5130
rect 5052 4998 5090 5130
rect 5292 4998 5330 5130
rect 5532 4998 5570 5130
rect 5772 4998 5810 5130
rect 6012 4998 6050 5130
rect 6252 4998 6290 5130
rect 6492 4998 6530 5130
rect 6732 4998 6770 5130
rect 6972 4998 7010 5130
rect 7212 4998 7250 5130
rect 7452 4998 7490 5130
rect 7692 4998 7730 5130
rect 7932 4998 7970 5130
rect 8172 4998 8210 5130
rect 8412 4998 8450 5130
rect 8652 4998 8690 5130
rect 8892 4998 8930 5130
rect 9132 4998 9170 5130
rect 9372 4998 9410 5130
rect 9612 4998 9650 5130
rect 9852 4998 9890 5130
rect 10092 4998 10130 5130
rect 10332 4998 10370 5130
rect 10572 4998 10610 5130
rect 10812 4998 10850 5130
rect 11052 4998 11090 5130
rect 11292 4998 11330 5130
rect 11532 4998 11570 5130
rect 11772 4998 11810 5130
rect 12012 4998 12050 5130
rect 12252 4998 12290 5130
rect -6412 2503 -6044 2537
rect -5824 2503 -5456 2537
rect -5236 2503 -4868 2537
rect -4648 2503 -4280 2537
rect -4060 2503 -3692 2537
rect -3472 2503 -3104 2537
rect -2884 2503 -2516 2537
rect -2296 2503 -1928 2537
rect -1708 2503 -1340 2537
rect -1120 2503 -752 2537
rect -532 2503 -164 2537
rect 56 2503 424 2537
rect 644 2503 1012 2537
rect 1232 2503 1600 2537
rect 1820 2503 2188 2537
rect 2408 2503 2776 2537
rect 2996 2503 3364 2537
rect 3584 2503 3952 2537
rect 4172 2503 4540 2537
rect 4760 2503 5128 2537
rect 5348 2503 5716 2537
rect 5936 2503 6304 2537
rect 6524 2503 6892 2537
rect 7112 2503 7480 2537
rect 7700 2503 8068 2537
rect 8288 2503 8656 2537
rect 8876 2503 9244 2537
rect 9464 2503 9832 2537
rect 10052 2503 10420 2537
rect 10640 2503 11008 2537
rect 11228 2503 11596 2537
rect 11816 2503 12184 2537
rect 12404 2503 12772 2537
rect 12992 2503 13360 2537
rect 13580 2503 13948 2537
rect 14168 2503 14536 2537
rect 14756 2503 15124 2537
rect 15344 2503 15712 2537
rect 15932 2503 16300 2537
rect 16520 2503 16888 2537
rect 17108 2503 17476 2537
rect 17696 2503 18064 2537
rect 18284 2503 18652 2537
rect 18872 2503 19240 2537
rect 19460 2503 19828 2537
rect 20048 2503 20416 2537
rect 20636 2503 21004 2537
rect 21224 2503 21592 2537
rect -6412 1575 -6044 1609
rect -6412 1503 -6044 1537
rect -5824 1575 -5456 1609
rect -5824 1503 -5456 1537
rect -5236 1575 -4868 1609
rect -5236 1503 -4868 1537
rect -4648 1575 -4280 1609
rect -4648 1503 -4280 1537
rect -4060 1575 -3692 1609
rect -4060 1503 -3692 1537
rect -3472 1575 -3104 1609
rect -3472 1503 -3104 1537
rect -2884 1575 -2516 1609
rect -2884 1503 -2516 1537
rect -2296 1575 -1928 1609
rect -2296 1503 -1928 1537
rect -1708 1575 -1340 1609
rect -1708 1503 -1340 1537
rect -1120 1575 -752 1609
rect -1120 1503 -752 1537
rect -532 1575 -164 1609
rect -532 1503 -164 1537
rect 56 1575 424 1609
rect 56 1503 424 1537
rect 644 1575 1012 1609
rect 644 1503 1012 1537
rect 1232 1575 1600 1609
rect 1232 1503 1600 1537
rect 1820 1575 2188 1609
rect 1820 1503 2188 1537
rect 2408 1575 2776 1609
rect 2408 1503 2776 1537
rect 2996 1575 3364 1609
rect 2996 1503 3364 1537
rect 3584 1575 3952 1609
rect 3584 1503 3952 1537
rect 4172 1575 4540 1609
rect 4172 1503 4540 1537
rect 4760 1575 5128 1609
rect 4760 1503 5128 1537
rect 5348 1575 5716 1609
rect 5348 1503 5716 1537
rect 5936 1575 6304 1609
rect 5936 1503 6304 1537
rect 6524 1575 6892 1609
rect 6524 1503 6892 1537
rect 7112 1575 7480 1609
rect 7112 1503 7480 1537
rect 7700 1575 8068 1609
rect 7700 1503 8068 1537
rect 8288 1575 8656 1609
rect 8288 1503 8656 1537
rect 8876 1575 9244 1609
rect 8876 1503 9244 1537
rect 9464 1575 9832 1609
rect 9464 1503 9832 1537
rect 10052 1575 10420 1609
rect 10052 1503 10420 1537
rect 10640 1575 11008 1609
rect 10640 1503 11008 1537
rect 11228 1575 11596 1609
rect 11228 1503 11596 1537
rect 11816 1575 12184 1609
rect 11816 1503 12184 1537
rect 12404 1575 12772 1609
rect 12404 1503 12772 1537
rect 12992 1575 13360 1609
rect 12992 1503 13360 1537
rect 13580 1575 13948 1609
rect 13580 1503 13948 1537
rect 14168 1575 14536 1609
rect 14168 1503 14536 1537
rect 14756 1575 15124 1609
rect 14756 1503 15124 1537
rect 15344 1575 15712 1609
rect 15344 1503 15712 1537
rect 15932 1575 16300 1609
rect 15932 1503 16300 1537
rect 16520 1575 16888 1609
rect 16520 1503 16888 1537
rect 17108 1575 17476 1609
rect 17108 1503 17476 1537
rect 17696 1575 18064 1609
rect 17696 1503 18064 1537
rect 18284 1575 18652 1609
rect 18284 1503 18652 1537
rect 18872 1575 19240 1609
rect 18872 1503 19240 1537
rect 19460 1575 19828 1609
rect 19460 1503 19828 1537
rect 20048 1575 20416 1609
rect 20048 1503 20416 1537
rect 20636 1575 21004 1609
rect 20636 1503 21004 1537
rect 21224 1575 21592 1609
rect 21224 1503 21592 1537
rect -6412 575 -6044 609
rect -6412 503 -6044 537
rect -5824 575 -5456 609
rect -5824 503 -5456 537
rect -5236 575 -4868 609
rect -5236 503 -4868 537
rect -4648 575 -4280 609
rect -4648 503 -4280 537
rect -4060 575 -3692 609
rect -4060 503 -3692 537
rect -3472 575 -3104 609
rect -3472 503 -3104 537
rect -2884 575 -2516 609
rect -2884 503 -2516 537
rect -2296 575 -1928 609
rect -2296 503 -1928 537
rect -1708 575 -1340 609
rect -1708 503 -1340 537
rect -1120 575 -752 609
rect -1120 503 -752 537
rect -532 575 -164 609
rect -532 503 -164 537
rect 56 575 424 609
rect 56 503 424 537
rect 644 575 1012 609
rect 644 503 1012 537
rect 1232 575 1600 609
rect 1232 503 1600 537
rect 1820 575 2188 609
rect 1820 503 2188 537
rect 2408 575 2776 609
rect 2408 503 2776 537
rect 2996 575 3364 609
rect 2996 503 3364 537
rect 3584 575 3952 609
rect 3584 503 3952 537
rect 4172 575 4540 609
rect 4172 503 4540 537
rect 4760 575 5128 609
rect 4760 503 5128 537
rect 5348 575 5716 609
rect 5348 503 5716 537
rect 5936 575 6304 609
rect 5936 503 6304 537
rect 6524 575 6892 609
rect 6524 503 6892 537
rect 7112 575 7480 609
rect 7112 503 7480 537
rect 7700 575 8068 609
rect 7700 503 8068 537
rect 8288 575 8656 609
rect 8288 503 8656 537
rect 8876 575 9244 609
rect 8876 503 9244 537
rect 9464 575 9832 609
rect 9464 503 9832 537
rect 10052 575 10420 609
rect 10052 503 10420 537
rect 10640 575 11008 609
rect 10640 503 11008 537
rect 11228 575 11596 609
rect 11228 503 11596 537
rect 11816 575 12184 609
rect 11816 503 12184 537
rect 12404 575 12772 609
rect 12404 503 12772 537
rect 12992 575 13360 609
rect 12992 503 13360 537
rect 13580 575 13948 609
rect 13580 503 13948 537
rect 14168 575 14536 609
rect 14168 503 14536 537
rect 14756 575 15124 609
rect 14756 503 15124 537
rect 15344 575 15712 609
rect 15344 503 15712 537
rect 15932 575 16300 609
rect 15932 503 16300 537
rect 16520 575 16888 609
rect 16520 503 16888 537
rect 17108 575 17476 609
rect 17108 503 17476 537
rect 17696 575 18064 609
rect 17696 503 18064 537
rect 18284 575 18652 609
rect 18284 503 18652 537
rect 18872 575 19240 609
rect 18872 503 19240 537
rect 19460 575 19828 609
rect 19460 503 19828 537
rect 20048 575 20416 609
rect 20048 503 20416 537
rect 20636 575 21004 609
rect 20636 503 21004 537
rect 21224 575 21592 609
rect 21224 503 21592 537
rect -6412 -425 -6044 -391
rect -5824 -425 -5456 -391
rect -5236 -425 -4868 -391
rect -4648 -425 -4280 -391
rect -4060 -425 -3692 -391
rect -3472 -425 -3104 -391
rect -2884 -425 -2516 -391
rect -2296 -425 -1928 -391
rect -1708 -425 -1340 -391
rect -1120 -425 -752 -391
rect -532 -425 -164 -391
rect 56 -425 424 -391
rect 644 -425 1012 -391
rect 1232 -425 1600 -391
rect 1820 -425 2188 -391
rect 2408 -425 2776 -391
rect 2996 -425 3364 -391
rect 3584 -425 3952 -391
rect 4172 -425 4540 -391
rect 4760 -425 5128 -391
rect 5348 -425 5716 -391
rect 5936 -425 6304 -391
rect 6524 -425 6892 -391
rect 7112 -425 7480 -391
rect 7700 -425 8068 -391
rect 8288 -425 8656 -391
rect 8876 -425 9244 -391
rect 9464 -425 9832 -391
rect 10052 -425 10420 -391
rect 10640 -425 11008 -391
rect 11228 -425 11596 -391
rect 11816 -425 12184 -391
rect 12404 -425 12772 -391
rect 12992 -425 13360 -391
rect 13580 -425 13948 -391
rect 14168 -425 14536 -391
rect 14756 -425 15124 -391
rect 15344 -425 15712 -391
rect 15932 -425 16300 -391
rect 16520 -425 16888 -391
rect 17108 -425 17476 -391
rect 17696 -425 18064 -391
rect 18284 -425 18652 -391
rect 18872 -425 19240 -391
rect 19460 -425 19828 -391
rect 20048 -425 20416 -391
rect 20636 -425 21004 -391
rect 21224 -425 21592 -391
rect 6640 -1952 6678 -1820
rect 6906 -1952 6944 -1820
rect 7172 -1952 7210 -1820
rect 7438 -1952 7476 -1820
rect 7704 -1952 7742 -1820
rect 7970 -1952 8008 -1820
rect 8236 -1952 8274 -1820
rect 8502 -1952 8540 -1820
rect 6640 -2962 6678 -2830
rect 6906 -2962 6944 -2830
rect 7172 -2962 7210 -2830
rect 7438 -2962 7476 -2830
rect 7704 -2962 7742 -2830
rect 7970 -2962 8008 -2830
rect 8236 -2962 8274 -2830
rect 8502 -2962 8540 -2830
rect 6640 -3972 6678 -3840
rect 6906 -3972 6944 -3840
rect 7172 -3972 7210 -3840
rect 7438 -3972 7476 -3840
rect 7704 -3972 7742 -3840
rect 7970 -3972 8008 -3840
rect 8236 -3972 8274 -3840
rect 8502 -3972 8540 -3840
rect 6640 -4982 6678 -4850
rect 6906 -4982 6944 -4850
rect 7172 -4982 7210 -4850
rect 7438 -4982 7476 -4850
rect 7704 -4982 7742 -4850
rect 7970 -4982 8008 -4850
rect 8236 -4982 8274 -4850
rect 8502 -4982 8540 -4850
rect 7212 -6144 7250 -6018
rect 7452 -6144 7490 -6018
rect 7692 -6144 7730 -6018
rect 7932 -6144 7970 -6018
rect 7212 -6952 7250 -6820
rect 7452 -6952 7490 -6820
rect 7692 -6952 7730 -6820
rect 7932 -6952 7970 -6820
rect 7212 -7760 7250 -7628
rect 7452 -7760 7490 -7628
rect 7692 -7760 7730 -7628
rect 7932 -7760 7970 -7628
<< xpolycontact >>
rect 13743 -3929 13813 -3497
rect 13743 -4921 13813 -4489
<< xpolyres >>
rect 13743 -4489 13813 -3929
<< locali >>
rect 2484 7056 2572 7090
rect 12610 7056 12698 7090
rect 2484 7022 2518 7056
rect 12664 7024 12698 7056
rect 2876 6614 2892 6746
rect 2930 6614 3132 6746
rect 3170 6614 3372 6746
rect 3410 6614 3612 6746
rect 3650 6614 3852 6746
rect 3890 6614 4092 6746
rect 4130 6614 4332 6746
rect 4370 6614 4572 6746
rect 4610 6614 4812 6746
rect 4850 6614 5052 6746
rect 5090 6614 5292 6746
rect 5330 6614 5532 6746
rect 5570 6614 5772 6746
rect 5810 6614 6012 6746
rect 6050 6614 6252 6746
rect 6290 6614 6492 6746
rect 6530 6614 6732 6746
rect 6770 6614 6972 6746
rect 7010 6614 7212 6746
rect 7250 6614 7452 6746
rect 7490 6614 7692 6746
rect 7730 6614 7932 6746
rect 7970 6614 8172 6746
rect 8210 6614 8412 6746
rect 8450 6614 8652 6746
rect 8690 6614 8892 6746
rect 8930 6614 9132 6746
rect 9170 6614 9372 6746
rect 9410 6614 9612 6746
rect 9650 6614 9852 6746
rect 9890 6614 10092 6746
rect 10130 6614 10332 6746
rect 10370 6614 10572 6746
rect 10610 6614 10812 6746
rect 10850 6614 11052 6746
rect 11090 6614 11292 6746
rect 11330 6614 11532 6746
rect 11570 6614 11772 6746
rect 11810 6614 12012 6746
rect 12050 6614 12252 6746
rect 12290 6614 12316 6746
rect 2830 6564 2864 6580
rect 2830 5972 2864 5988
rect 2958 6564 2992 6580
rect 2958 5972 2992 5988
rect 3070 6564 3104 6580
rect 3070 5972 3104 5988
rect 3198 6564 3232 6580
rect 3198 5972 3232 5988
rect 3310 6564 3344 6580
rect 3310 5972 3344 5988
rect 3438 6564 3472 6580
rect 3438 5972 3472 5988
rect 3550 6564 3584 6580
rect 3550 5972 3584 5988
rect 3678 6564 3712 6580
rect 3678 5972 3712 5988
rect 3790 6564 3824 6580
rect 3790 5972 3824 5988
rect 3918 6564 3952 6580
rect 3918 5972 3952 5988
rect 4030 6564 4064 6580
rect 4030 5972 4064 5988
rect 4158 6564 4192 6580
rect 4158 5972 4192 5988
rect 4270 6564 4304 6580
rect 4270 5972 4304 5988
rect 4398 6564 4432 6580
rect 4398 5972 4432 5988
rect 4510 6564 4544 6580
rect 4510 5972 4544 5988
rect 4638 6564 4672 6580
rect 4638 5972 4672 5988
rect 4750 6564 4784 6580
rect 4750 5972 4784 5988
rect 4878 6564 4912 6580
rect 4878 5972 4912 5988
rect 4990 6564 5024 6580
rect 4990 5972 5024 5988
rect 5118 6564 5152 6580
rect 5118 5972 5152 5988
rect 5230 6564 5264 6580
rect 5230 5972 5264 5988
rect 5358 6564 5392 6580
rect 5358 5972 5392 5988
rect 5470 6564 5504 6580
rect 5470 5972 5504 5988
rect 5598 6564 5632 6580
rect 5598 5972 5632 5988
rect 5710 6564 5744 6580
rect 5710 5972 5744 5988
rect 5838 6564 5872 6580
rect 5838 5972 5872 5988
rect 5950 6564 5984 6580
rect 5950 5972 5984 5988
rect 6078 6564 6112 6580
rect 6078 5972 6112 5988
rect 6190 6564 6224 6580
rect 6190 5972 6224 5988
rect 6318 6564 6352 6580
rect 6318 5972 6352 5988
rect 6430 6564 6464 6580
rect 6430 5972 6464 5988
rect 6558 6564 6592 6580
rect 6558 5972 6592 5988
rect 6670 6564 6704 6580
rect 6670 5972 6704 5988
rect 6798 6564 6832 6580
rect 6798 5972 6832 5988
rect 6910 6564 6944 6580
rect 6910 5972 6944 5988
rect 7038 6564 7072 6580
rect 7038 5972 7072 5988
rect 7150 6564 7184 6580
rect 7150 5972 7184 5988
rect 7278 6564 7312 6580
rect 7278 5972 7312 5988
rect 7390 6564 7424 6580
rect 7390 5972 7424 5988
rect 7518 6564 7552 6580
rect 7518 5972 7552 5988
rect 7630 6564 7664 6580
rect 7630 5972 7664 5988
rect 7758 6564 7792 6580
rect 7758 5972 7792 5988
rect 7870 6564 7904 6580
rect 7870 5972 7904 5988
rect 7998 6564 8032 6580
rect 7998 5972 8032 5988
rect 8110 6564 8144 6580
rect 8110 5972 8144 5988
rect 8238 6564 8272 6580
rect 8238 5972 8272 5988
rect 8350 6564 8384 6580
rect 8350 5972 8384 5988
rect 8478 6564 8512 6580
rect 8478 5972 8512 5988
rect 8590 6564 8624 6580
rect 8590 5972 8624 5988
rect 8718 6564 8752 6580
rect 8718 5972 8752 5988
rect 8830 6564 8864 6580
rect 8830 5972 8864 5988
rect 8958 6564 8992 6580
rect 8958 5972 8992 5988
rect 9070 6564 9104 6580
rect 9070 5972 9104 5988
rect 9198 6564 9232 6580
rect 9198 5972 9232 5988
rect 9310 6564 9344 6580
rect 9310 5972 9344 5988
rect 9438 6564 9472 6580
rect 9438 5972 9472 5988
rect 9550 6564 9584 6580
rect 9550 5972 9584 5988
rect 9678 6564 9712 6580
rect 9678 5972 9712 5988
rect 9790 6564 9824 6580
rect 9790 5972 9824 5988
rect 9918 6564 9952 6580
rect 9918 5972 9952 5988
rect 10030 6564 10064 6580
rect 10030 5972 10064 5988
rect 10158 6564 10192 6580
rect 10158 5972 10192 5988
rect 10270 6564 10304 6580
rect 10270 5972 10304 5988
rect 10398 6564 10432 6580
rect 10398 5972 10432 5988
rect 10510 6564 10544 6580
rect 10510 5972 10544 5988
rect 10638 6564 10672 6580
rect 10638 5972 10672 5988
rect 10750 6564 10784 6580
rect 10750 5972 10784 5988
rect 10878 6564 10912 6580
rect 10878 5972 10912 5988
rect 10990 6564 11024 6580
rect 10990 5972 11024 5988
rect 11118 6564 11152 6580
rect 11118 5972 11152 5988
rect 11230 6564 11264 6580
rect 11230 5972 11264 5988
rect 11358 6564 11392 6580
rect 11358 5972 11392 5988
rect 11470 6564 11504 6580
rect 11470 5972 11504 5988
rect 11598 6564 11632 6580
rect 11598 5972 11632 5988
rect 11710 6564 11744 6580
rect 11710 5972 11744 5988
rect 11838 6564 11872 6580
rect 11838 5972 11872 5988
rect 11950 6564 11984 6580
rect 11950 5972 11984 5988
rect 12078 6564 12112 6580
rect 12078 5972 12112 5988
rect 12190 6564 12224 6580
rect 12190 5972 12224 5988
rect 12318 6564 12352 6580
rect 12318 5972 12352 5988
rect 2876 5806 2892 5938
rect 2930 5806 3132 5938
rect 3170 5806 3372 5938
rect 3410 5806 3612 5938
rect 3650 5806 3852 5938
rect 3890 5806 4092 5938
rect 4130 5806 4332 5938
rect 4370 5806 4572 5938
rect 4610 5806 4812 5938
rect 4850 5806 5052 5938
rect 5090 5806 5292 5938
rect 5330 5806 5532 5938
rect 5570 5806 5772 5938
rect 5810 5806 6012 5938
rect 6050 5806 6252 5938
rect 6290 5806 6492 5938
rect 6530 5806 6732 5938
rect 6770 5806 6972 5938
rect 7010 5806 7212 5938
rect 7250 5806 7452 5938
rect 7490 5806 7692 5938
rect 7730 5806 7932 5938
rect 7970 5806 8172 5938
rect 8210 5806 8412 5938
rect 8450 5806 8652 5938
rect 8690 5806 8892 5938
rect 8930 5806 9132 5938
rect 9170 5806 9372 5938
rect 9410 5806 9612 5938
rect 9650 5806 9852 5938
rect 9890 5806 10092 5938
rect 10130 5806 10332 5938
rect 10370 5806 10572 5938
rect 10610 5806 10812 5938
rect 10850 5806 11052 5938
rect 11090 5806 11292 5938
rect 11330 5806 11532 5938
rect 11570 5806 11772 5938
rect 11810 5806 12012 5938
rect 12050 5806 12252 5938
rect 12290 5806 12316 5938
rect 2830 5756 2864 5772
rect 2830 5164 2864 5180
rect 2958 5756 2992 5772
rect 2958 5164 2992 5180
rect 3070 5756 3104 5772
rect 3070 5164 3104 5180
rect 3198 5756 3232 5772
rect 3198 5164 3232 5180
rect 3310 5756 3344 5772
rect 3310 5164 3344 5180
rect 3438 5756 3472 5772
rect 3438 5164 3472 5180
rect 3550 5756 3584 5772
rect 3550 5164 3584 5180
rect 3678 5756 3712 5772
rect 3678 5164 3712 5180
rect 3790 5756 3824 5772
rect 3790 5164 3824 5180
rect 3918 5756 3952 5772
rect 3918 5164 3952 5180
rect 4030 5756 4064 5772
rect 4030 5164 4064 5180
rect 4158 5756 4192 5772
rect 4158 5164 4192 5180
rect 4270 5756 4304 5772
rect 4270 5164 4304 5180
rect 4398 5756 4432 5772
rect 4398 5164 4432 5180
rect 4510 5756 4544 5772
rect 4510 5164 4544 5180
rect 4638 5756 4672 5772
rect 4638 5164 4672 5180
rect 4750 5756 4784 5772
rect 4750 5164 4784 5180
rect 4878 5756 4912 5772
rect 4878 5164 4912 5180
rect 4990 5756 5024 5772
rect 4990 5164 5024 5180
rect 5118 5756 5152 5772
rect 5118 5164 5152 5180
rect 5230 5756 5264 5772
rect 5230 5164 5264 5180
rect 5358 5756 5392 5772
rect 5358 5164 5392 5180
rect 5470 5756 5504 5772
rect 5470 5164 5504 5180
rect 5598 5756 5632 5772
rect 5598 5164 5632 5180
rect 5710 5756 5744 5772
rect 5710 5164 5744 5180
rect 5838 5756 5872 5772
rect 5838 5164 5872 5180
rect 5950 5756 5984 5772
rect 5950 5164 5984 5180
rect 6078 5756 6112 5772
rect 6078 5164 6112 5180
rect 6190 5756 6224 5772
rect 6190 5164 6224 5180
rect 6318 5756 6352 5772
rect 6318 5164 6352 5180
rect 6430 5756 6464 5772
rect 6430 5164 6464 5180
rect 6558 5756 6592 5772
rect 6558 5164 6592 5180
rect 6670 5756 6704 5772
rect 6670 5164 6704 5180
rect 6798 5756 6832 5772
rect 6798 5164 6832 5180
rect 6910 5756 6944 5772
rect 6910 5164 6944 5180
rect 7038 5756 7072 5772
rect 7038 5164 7072 5180
rect 7150 5756 7184 5772
rect 7150 5164 7184 5180
rect 7278 5756 7312 5772
rect 7278 5164 7312 5180
rect 7390 5756 7424 5772
rect 7390 5164 7424 5180
rect 7518 5756 7552 5772
rect 7518 5164 7552 5180
rect 7630 5756 7664 5772
rect 7630 5164 7664 5180
rect 7758 5756 7792 5772
rect 7758 5164 7792 5180
rect 7870 5756 7904 5772
rect 7870 5164 7904 5180
rect 7998 5756 8032 5772
rect 7998 5164 8032 5180
rect 8110 5756 8144 5772
rect 8110 5164 8144 5180
rect 8238 5756 8272 5772
rect 8238 5164 8272 5180
rect 8350 5756 8384 5772
rect 8350 5164 8384 5180
rect 8478 5756 8512 5772
rect 8478 5164 8512 5180
rect 8590 5756 8624 5772
rect 8590 5164 8624 5180
rect 8718 5756 8752 5772
rect 8718 5164 8752 5180
rect 8830 5756 8864 5772
rect 8830 5164 8864 5180
rect 8958 5756 8992 5772
rect 8958 5164 8992 5180
rect 9070 5756 9104 5772
rect 9070 5164 9104 5180
rect 9198 5756 9232 5772
rect 9198 5164 9232 5180
rect 9310 5756 9344 5772
rect 9310 5164 9344 5180
rect 9438 5756 9472 5772
rect 9438 5164 9472 5180
rect 9550 5756 9584 5772
rect 9550 5164 9584 5180
rect 9678 5756 9712 5772
rect 9678 5164 9712 5180
rect 9790 5756 9824 5772
rect 9790 5164 9824 5180
rect 9918 5756 9952 5772
rect 9918 5164 9952 5180
rect 10030 5756 10064 5772
rect 10030 5164 10064 5180
rect 10158 5756 10192 5772
rect 10158 5164 10192 5180
rect 10270 5756 10304 5772
rect 10270 5164 10304 5180
rect 10398 5756 10432 5772
rect 10398 5164 10432 5180
rect 10510 5756 10544 5772
rect 10510 5164 10544 5180
rect 10638 5756 10672 5772
rect 10638 5164 10672 5180
rect 10750 5756 10784 5772
rect 10750 5164 10784 5180
rect 10878 5756 10912 5772
rect 10878 5164 10912 5180
rect 10990 5756 11024 5772
rect 10990 5164 11024 5180
rect 11118 5756 11152 5772
rect 11118 5164 11152 5180
rect 11230 5756 11264 5772
rect 11230 5164 11264 5180
rect 11358 5756 11392 5772
rect 11358 5164 11392 5180
rect 11470 5756 11504 5772
rect 11470 5164 11504 5180
rect 11598 5756 11632 5772
rect 11598 5164 11632 5180
rect 11710 5756 11744 5772
rect 11710 5164 11744 5180
rect 11838 5756 11872 5772
rect 11838 5164 11872 5180
rect 11950 5756 11984 5772
rect 11950 5164 11984 5180
rect 12078 5756 12112 5772
rect 12078 5164 12112 5180
rect 12190 5756 12224 5772
rect 12190 5164 12224 5180
rect 12318 5756 12352 5772
rect 12318 5164 12352 5180
rect 2876 4998 2892 5130
rect 2930 4998 3132 5130
rect 3170 4998 3372 5130
rect 3410 4998 3612 5130
rect 3650 4998 3852 5130
rect 3890 4998 4092 5130
rect 4130 4998 4332 5130
rect 4370 4998 4572 5130
rect 4610 4998 4812 5130
rect 4850 4998 5052 5130
rect 5090 4998 5292 5130
rect 5330 4998 5532 5130
rect 5570 4998 5772 5130
rect 5810 4998 6012 5130
rect 6050 4998 6252 5130
rect 6290 4998 6492 5130
rect 6530 4998 6732 5130
rect 6770 4998 6972 5130
rect 7010 4998 7212 5130
rect 7250 4998 7452 5130
rect 7490 4998 7692 5130
rect 7730 4998 7932 5130
rect 7970 4998 8172 5130
rect 8210 4998 8412 5130
rect 8450 4998 8652 5130
rect 8690 4998 8892 5130
rect 8930 4998 9132 5130
rect 9170 4998 9372 5130
rect 9410 4998 9612 5130
rect 9650 4998 9852 5130
rect 9890 4998 10092 5130
rect 10130 4998 10332 5130
rect 10370 4998 10572 5130
rect 10610 4998 10812 5130
rect 10850 4998 11052 5130
rect 11090 4998 11292 5130
rect 11330 4998 11532 5130
rect 11570 4998 11772 5130
rect 11810 4998 12012 5130
rect 12050 4998 12252 5130
rect 12290 4998 12316 5130
rect 2484 4654 2518 4742
rect 12664 4654 12698 4742
rect -6820 2854 -6660 2888
rect 21862 2860 22000 2888
rect 21862 2854 21966 2860
rect -6820 2826 -6786 2854
rect -6428 2537 5332 2538
rect 5732 2537 5920 2538
rect 6320 2537 6508 2538
rect 6908 2537 7096 2538
rect 7496 2537 7684 2538
rect 8084 2537 8272 2538
rect 8672 2537 8860 2538
rect 9260 2537 9448 2538
rect 9848 2537 21608 2538
rect -6428 2503 -6412 2537
rect -6044 2503 -5824 2537
rect -5456 2503 -5236 2537
rect -4868 2503 -4648 2537
rect -4280 2503 -4060 2537
rect -3692 2503 -3472 2537
rect -3104 2503 -2884 2537
rect -2516 2503 -2296 2537
rect -1928 2503 -1708 2537
rect -1340 2503 -1120 2537
rect -752 2503 -532 2537
rect -164 2503 56 2537
rect 424 2503 644 2537
rect 1012 2503 1232 2537
rect 1600 2503 1820 2537
rect 2188 2503 2408 2537
rect 2776 2503 2996 2537
rect 3364 2503 3584 2537
rect 3952 2503 4172 2537
rect 4540 2503 4760 2537
rect 5128 2503 5348 2537
rect 5716 2503 5936 2537
rect 6304 2503 6524 2537
rect 6892 2503 7112 2537
rect 7480 2503 7700 2537
rect 8068 2503 8288 2537
rect 8656 2503 8876 2537
rect 9244 2503 9464 2537
rect 9832 2503 10052 2537
rect 10420 2503 10640 2537
rect 11008 2503 11228 2537
rect 11596 2503 11816 2537
rect 12184 2503 12404 2537
rect 12772 2503 12992 2537
rect 13360 2503 13580 2537
rect 13948 2503 14168 2537
rect 14536 2503 14756 2537
rect 15124 2503 15344 2537
rect 15712 2503 15932 2537
rect 16300 2503 16520 2537
rect 16888 2503 17108 2537
rect 17476 2503 17696 2537
rect 18064 2503 18284 2537
rect 18652 2503 18872 2537
rect 19240 2503 19460 2537
rect 19828 2503 20048 2537
rect 20416 2503 20636 2537
rect 21004 2503 21224 2537
rect 21592 2503 21608 2537
rect -6428 2502 5332 2503
rect 5732 2502 5920 2503
rect 6320 2502 6508 2503
rect 6908 2502 7096 2503
rect 5286 2460 5332 2502
rect 7496 2460 7684 2503
rect 8084 2502 8272 2503
rect 8672 2502 8860 2503
rect 9260 2502 9448 2503
rect 9848 2502 21608 2503
rect 9848 2460 9894 2502
rect -6474 2444 -6440 2460
rect -6474 1652 -6440 1668
rect -6016 2444 -5982 2460
rect -6016 1652 -5982 1668
rect -5886 2444 -5852 2460
rect -5886 1652 -5852 1668
rect -5428 2444 -5394 2460
rect -5428 1652 -5394 1668
rect -5298 2444 -5264 2460
rect -5298 1652 -5264 1668
rect -4840 2444 -4806 2460
rect -4840 1652 -4806 1668
rect -4710 2444 -4676 2460
rect -4710 1652 -4676 1668
rect -4252 2444 -4218 2460
rect -4252 1652 -4218 1668
rect -4122 2444 -4088 2460
rect -4122 1652 -4088 1668
rect -3664 2444 -3630 2460
rect -3664 1652 -3630 1668
rect -3534 2444 -3500 2460
rect -3534 1652 -3500 1668
rect -3076 2444 -3042 2460
rect -3076 1652 -3042 1668
rect -2946 2444 -2912 2460
rect -2946 1652 -2912 1668
rect -2488 2444 -2454 2460
rect -2488 1652 -2454 1668
rect -2358 2444 -2324 2460
rect -2358 1652 -2324 1668
rect -1900 2444 -1866 2460
rect -1900 1652 -1866 1668
rect -1770 2444 -1736 2460
rect -1770 1652 -1736 1668
rect -1312 2444 -1278 2460
rect -1312 1652 -1278 1668
rect -1182 2444 -1148 2460
rect -1182 1652 -1148 1668
rect -724 2444 -690 2460
rect -724 1652 -690 1668
rect -594 2444 -560 2460
rect -594 1652 -560 1668
rect -136 2444 -102 2460
rect -136 1652 -102 1668
rect -6 2444 28 2460
rect -6 1652 28 1668
rect 452 2444 486 2460
rect 452 1652 486 1668
rect 582 2444 616 2460
rect 582 1652 616 1668
rect 1040 2444 1074 2460
rect 1040 1652 1074 1668
rect 1170 2444 1204 2460
rect 1170 1652 1204 1668
rect 1628 2444 1662 2460
rect 1628 1652 1662 1668
rect 1758 2444 1792 2460
rect 1758 1652 1792 1668
rect 2216 2444 2250 2460
rect 2216 1652 2250 1668
rect 2346 2444 2380 2460
rect 2346 1652 2380 1668
rect 2804 2444 2838 2460
rect 2804 1652 2838 1668
rect 2934 2444 2968 2460
rect 2934 1652 2968 1668
rect 3392 2444 3426 2460
rect 3392 1652 3426 1668
rect 3522 2444 3556 2460
rect 3522 1652 3556 1668
rect 3980 2444 4014 2460
rect 3980 1652 4014 1668
rect 4110 2444 4144 2460
rect 4110 1652 4144 1668
rect 4568 2444 4602 2460
rect 4568 1652 4602 1668
rect 4698 2444 4732 2460
rect 4698 1652 4732 1668
rect 5156 2444 5190 2460
rect 5156 1652 5190 1668
rect 5286 2444 5320 2460
rect 5286 1610 5320 1668
rect 5744 2444 5778 2460
rect 5744 1652 5778 1668
rect 5874 2444 5908 2460
rect 5874 1652 5908 1668
rect 6332 2444 6366 2460
rect 6332 1652 6366 1668
rect 6462 2444 6496 2460
rect 6462 1652 6496 1668
rect 6920 2444 6954 2460
rect 6920 1652 6954 1668
rect 7050 2444 7084 2460
rect 7050 1652 7084 1668
rect 7508 2444 7672 2460
rect 7542 1668 7638 2444
rect 7508 1610 7672 1668
rect 8096 2444 8130 2460
rect 8096 1652 8130 1668
rect 8226 2444 8260 2460
rect 8226 1652 8260 1668
rect 8684 2444 8718 2460
rect 8684 1652 8718 1668
rect 8814 2444 8848 2460
rect 8814 1652 8848 1668
rect 9272 2444 9306 2460
rect 9272 1652 9306 1668
rect 9402 2444 9436 2460
rect 9402 1652 9436 1668
rect 9860 2444 9894 2460
rect 9860 1610 9894 1668
rect 9990 2444 10024 2460
rect 9990 1652 10024 1668
rect 10448 2444 10482 2460
rect 10448 1652 10482 1668
rect 10578 2444 10612 2460
rect 10578 1652 10612 1668
rect 11036 2444 11070 2460
rect 11036 1652 11070 1668
rect 11166 2444 11200 2460
rect 11166 1652 11200 1668
rect 11624 2444 11658 2460
rect 11624 1652 11658 1668
rect 11754 2444 11788 2460
rect 11754 1652 11788 1668
rect 12212 2444 12246 2460
rect 12212 1652 12246 1668
rect 12342 2444 12376 2460
rect 12342 1652 12376 1668
rect 12800 2444 12834 2460
rect 12800 1652 12834 1668
rect 12930 2444 12964 2460
rect 12930 1652 12964 1668
rect 13388 2444 13422 2460
rect 13388 1652 13422 1668
rect 13518 2444 13552 2460
rect 13518 1652 13552 1668
rect 13976 2444 14010 2460
rect 13976 1652 14010 1668
rect 14106 2444 14140 2460
rect 14106 1652 14140 1668
rect 14564 2444 14598 2460
rect 14564 1652 14598 1668
rect 14694 2444 14728 2460
rect 14694 1652 14728 1668
rect 15152 2444 15186 2460
rect 15152 1652 15186 1668
rect 15282 2444 15316 2460
rect 15282 1652 15316 1668
rect 15740 2444 15774 2460
rect 15740 1652 15774 1668
rect 15870 2444 15904 2460
rect 15870 1652 15904 1668
rect 16328 2444 16362 2460
rect 16328 1652 16362 1668
rect 16458 2444 16492 2460
rect 16458 1652 16492 1668
rect 16916 2444 16950 2460
rect 16916 1652 16950 1668
rect 17046 2444 17080 2460
rect 17046 1652 17080 1668
rect 17504 2444 17538 2460
rect 17504 1652 17538 1668
rect 17634 2444 17668 2460
rect 17634 1652 17668 1668
rect 18092 2444 18126 2460
rect 18092 1652 18126 1668
rect 18222 2444 18256 2460
rect 18222 1652 18256 1668
rect 18680 2444 18714 2460
rect 18680 1652 18714 1668
rect 18810 2444 18844 2460
rect 18810 1652 18844 1668
rect 19268 2444 19302 2460
rect 19268 1652 19302 1668
rect 19398 2444 19432 2460
rect 19398 1652 19432 1668
rect 19856 2444 19890 2460
rect 19856 1652 19890 1668
rect 19986 2444 20020 2460
rect 19986 1652 20020 1668
rect 20444 2444 20478 2460
rect 20444 1652 20478 1668
rect 20574 2444 20608 2460
rect 20574 1652 20608 1668
rect 21032 2444 21066 2460
rect 21032 1652 21066 1668
rect 21162 2444 21196 2460
rect 21162 1652 21196 1668
rect 21620 2444 21654 2460
rect 21620 1652 21654 1668
rect -6428 1609 5332 1610
rect 5732 1609 5920 1610
rect 6320 1609 6508 1610
rect 6908 1609 7096 1610
rect 7496 1609 7684 1610
rect 8084 1609 8272 1610
rect 8672 1609 8860 1610
rect 9260 1609 9448 1610
rect 9848 1609 21608 1610
rect -6428 1575 -6412 1609
rect -6044 1575 -5824 1609
rect -5456 1575 -5236 1609
rect -4868 1575 -4648 1609
rect -4280 1575 -4060 1609
rect -3692 1575 -3472 1609
rect -3104 1575 -2884 1609
rect -2516 1575 -2296 1609
rect -1928 1575 -1708 1609
rect -1340 1575 -1120 1609
rect -752 1575 -532 1609
rect -164 1575 56 1609
rect 424 1575 644 1609
rect 1012 1575 1232 1609
rect 1600 1575 1820 1609
rect 2188 1575 2408 1609
rect 2776 1575 2996 1609
rect 3364 1575 3584 1609
rect 3952 1575 4172 1609
rect 4540 1575 4760 1609
rect 5128 1575 5348 1609
rect 5716 1575 5936 1609
rect 6304 1575 6524 1609
rect 6892 1575 7112 1609
rect 7480 1575 7700 1609
rect 8068 1575 8288 1609
rect 8656 1575 8876 1609
rect 9244 1575 9464 1609
rect 9832 1575 10052 1609
rect 10420 1575 10640 1609
rect 11008 1575 11228 1609
rect 11596 1575 11816 1609
rect 12184 1575 12404 1609
rect 12772 1575 12992 1609
rect 13360 1575 13580 1609
rect 13948 1575 14168 1609
rect 14536 1575 14756 1609
rect 15124 1575 15344 1609
rect 15712 1575 15932 1609
rect 16300 1575 16520 1609
rect 16888 1575 17108 1609
rect 17476 1575 17696 1609
rect 18064 1575 18284 1609
rect 18652 1575 18872 1609
rect 19240 1575 19460 1609
rect 19828 1575 20048 1609
rect 20416 1575 20636 1609
rect 21004 1575 21224 1609
rect 21592 1575 21608 1609
rect -6428 1537 5332 1575
rect 5732 1537 5920 1575
rect 6320 1574 6508 1575
rect 6320 1537 6508 1538
rect 6908 1537 7096 1575
rect 7496 1537 7684 1575
rect 8084 1537 8272 1575
rect 8672 1574 8860 1575
rect 8672 1537 8860 1538
rect 9260 1537 9448 1575
rect 9848 1537 21608 1575
rect -6428 1503 -6412 1537
rect -6044 1503 -5824 1537
rect -5456 1503 -5236 1537
rect -4868 1503 -4648 1537
rect -4280 1503 -4060 1537
rect -3692 1503 -3472 1537
rect -3104 1503 -2884 1537
rect -2516 1503 -2296 1537
rect -1928 1503 -1708 1537
rect -1340 1503 -1120 1537
rect -752 1503 -532 1537
rect -164 1503 56 1537
rect 424 1503 644 1537
rect 1012 1503 1232 1537
rect 1600 1503 1820 1537
rect 2188 1503 2408 1537
rect 2776 1503 2996 1537
rect 3364 1503 3584 1537
rect 3952 1503 4172 1537
rect 4540 1503 4760 1537
rect 5128 1503 5348 1537
rect 5716 1503 5936 1537
rect 6304 1503 6524 1537
rect 6892 1503 7112 1537
rect 7480 1503 7700 1537
rect 8068 1503 8288 1537
rect 8656 1503 8876 1537
rect 9244 1503 9464 1537
rect 9832 1503 10052 1537
rect 10420 1503 10640 1537
rect 11008 1503 11228 1537
rect 11596 1503 11816 1537
rect 12184 1503 12404 1537
rect 12772 1503 12992 1537
rect 13360 1503 13580 1537
rect 13948 1503 14168 1537
rect 14536 1503 14756 1537
rect 15124 1503 15344 1537
rect 15712 1503 15932 1537
rect 16300 1503 16520 1537
rect 16888 1503 17108 1537
rect 17476 1503 17696 1537
rect 18064 1503 18284 1537
rect 18652 1503 18872 1537
rect 19240 1503 19460 1537
rect 19828 1503 20048 1537
rect 20416 1503 20636 1537
rect 21004 1503 21224 1537
rect 21592 1503 21608 1537
rect -6428 1502 5332 1503
rect 5732 1502 5920 1503
rect 6320 1502 6508 1503
rect 6908 1502 7096 1503
rect 7496 1502 7684 1503
rect 8084 1502 8272 1503
rect 8672 1502 8860 1503
rect 9260 1502 9448 1503
rect 9848 1502 21608 1503
rect -6474 1444 -6440 1460
rect -6474 652 -6440 668
rect -6016 1444 -5982 1460
rect -6016 652 -5982 668
rect -5886 1444 -5852 1460
rect -5886 652 -5852 668
rect -5428 1444 -5394 1460
rect -5428 652 -5394 668
rect -5298 1444 -5264 1460
rect -5298 652 -5264 668
rect -4840 1444 -4806 1460
rect -4840 652 -4806 668
rect -4710 1444 -4676 1460
rect -4710 652 -4676 668
rect -4252 1444 -4218 1460
rect -4252 652 -4218 668
rect -4122 1444 -4088 1460
rect -4122 652 -4088 668
rect -3664 1444 -3630 1460
rect -3664 652 -3630 668
rect -3534 1444 -3500 1460
rect -3534 652 -3500 668
rect -3076 1444 -3042 1460
rect -3076 652 -3042 668
rect -2946 1444 -2912 1460
rect -2946 652 -2912 668
rect -2488 1444 -2454 1460
rect -2488 652 -2454 668
rect -2358 1444 -2324 1460
rect -2358 652 -2324 668
rect -1900 1444 -1866 1460
rect -1900 652 -1866 668
rect -1770 1444 -1736 1460
rect -1770 652 -1736 668
rect -1312 1444 -1278 1460
rect -1312 652 -1278 668
rect -1182 1444 -1148 1460
rect -1182 652 -1148 668
rect -724 1444 -690 1460
rect -724 652 -690 668
rect -594 1444 -560 1460
rect -594 652 -560 668
rect -136 1444 -102 1460
rect -136 652 -102 668
rect -6 1444 28 1460
rect -6 652 28 668
rect 452 1444 486 1460
rect 452 652 486 668
rect 582 1444 616 1460
rect 582 652 616 668
rect 1040 1444 1074 1460
rect 1040 652 1074 668
rect 1170 1444 1204 1460
rect 1170 652 1204 668
rect 1628 1444 1662 1460
rect 1628 652 1662 668
rect 1758 1444 1792 1460
rect 1758 652 1792 668
rect 2216 1444 2250 1460
rect 2216 652 2250 668
rect 2346 1444 2380 1460
rect 2346 652 2380 668
rect 2804 1444 2838 1460
rect 2804 652 2838 668
rect 2934 1444 2968 1460
rect 2934 652 2968 668
rect 3392 1444 3426 1460
rect 3392 652 3426 668
rect 3522 1444 3556 1460
rect 3522 652 3556 668
rect 3980 1444 4014 1460
rect 3980 652 4014 668
rect 4110 1444 4144 1460
rect 4110 652 4144 668
rect 4568 1444 4602 1460
rect 4568 652 4602 668
rect 4698 1444 4732 1460
rect 4698 652 4732 668
rect 5156 1444 5190 1460
rect 5156 652 5190 668
rect 5286 1444 5320 1502
rect 5286 610 5320 668
rect 5744 1444 5778 1460
rect 5744 652 5778 668
rect 5874 1444 5908 1460
rect 5874 652 5908 668
rect 6332 1444 6366 1460
rect 6332 652 6366 668
rect 6462 1444 6496 1460
rect 6462 652 6496 668
rect 6920 1444 6954 1460
rect 6920 652 6954 668
rect 7050 1444 7084 1460
rect 7050 652 7084 668
rect 7508 1444 7672 1502
rect 7542 668 7638 1444
rect 7508 610 7672 668
rect 8096 1444 8130 1460
rect 8096 652 8130 668
rect 8226 1444 8260 1460
rect 8226 652 8260 668
rect 8684 1444 8718 1460
rect 8684 652 8718 668
rect 8814 1444 8848 1460
rect 8814 652 8848 668
rect 9272 1444 9306 1460
rect 9272 652 9306 668
rect 9402 1444 9436 1460
rect 9402 652 9436 668
rect 9860 1444 9894 1502
rect 9860 610 9894 668
rect 9990 1444 10024 1460
rect 9990 652 10024 668
rect 10448 1444 10482 1460
rect 10448 652 10482 668
rect 10578 1444 10612 1460
rect 10578 652 10612 668
rect 11036 1444 11070 1460
rect 11036 652 11070 668
rect 11166 1444 11200 1460
rect 11166 652 11200 668
rect 11624 1444 11658 1460
rect 11624 652 11658 668
rect 11754 1444 11788 1460
rect 11754 652 11788 668
rect 12212 1444 12246 1460
rect 12212 652 12246 668
rect 12342 1444 12376 1460
rect 12342 652 12376 668
rect 12800 1444 12834 1460
rect 12800 652 12834 668
rect 12930 1444 12964 1460
rect 12930 652 12964 668
rect 13388 1444 13422 1460
rect 13388 652 13422 668
rect 13518 1444 13552 1460
rect 13518 652 13552 668
rect 13976 1444 14010 1460
rect 13976 652 14010 668
rect 14106 1444 14140 1460
rect 14106 652 14140 668
rect 14564 1444 14598 1460
rect 14564 652 14598 668
rect 14694 1444 14728 1460
rect 14694 652 14728 668
rect 15152 1444 15186 1460
rect 15152 652 15186 668
rect 15282 1444 15316 1460
rect 15282 652 15316 668
rect 15740 1444 15774 1460
rect 15740 652 15774 668
rect 15870 1444 15904 1460
rect 15870 652 15904 668
rect 16328 1444 16362 1460
rect 16328 652 16362 668
rect 16458 1444 16492 1460
rect 16458 652 16492 668
rect 16916 1444 16950 1460
rect 16916 652 16950 668
rect 17046 1444 17080 1460
rect 17046 652 17080 668
rect 17504 1444 17538 1460
rect 17504 652 17538 668
rect 17634 1444 17668 1460
rect 17634 652 17668 668
rect 18092 1444 18126 1460
rect 18092 652 18126 668
rect 18222 1444 18256 1460
rect 18222 652 18256 668
rect 18680 1444 18714 1460
rect 18680 652 18714 668
rect 18810 1444 18844 1460
rect 18810 652 18844 668
rect 19268 1444 19302 1460
rect 19268 652 19302 668
rect 19398 1444 19432 1460
rect 19398 652 19432 668
rect 19856 1444 19890 1460
rect 19856 652 19890 668
rect 19986 1444 20020 1460
rect 19986 652 20020 668
rect 20444 1444 20478 1460
rect 20444 652 20478 668
rect 20574 1444 20608 1460
rect 20574 652 20608 668
rect 21032 1444 21066 1460
rect 21032 652 21066 668
rect 21162 1444 21196 1460
rect 21162 652 21196 668
rect 21620 1444 21654 1460
rect 21620 652 21654 668
rect -6428 609 5332 610
rect 5732 609 5920 610
rect 6320 609 6508 610
rect 6908 609 7096 610
rect 7496 609 7684 610
rect 8084 609 8272 610
rect 8672 609 8860 610
rect 9260 609 9448 610
rect 9848 609 21608 610
rect -6428 575 -6412 609
rect -6044 575 -5824 609
rect -5456 575 -5236 609
rect -4868 575 -4648 609
rect -4280 575 -4060 609
rect -3692 575 -3472 609
rect -3104 575 -2884 609
rect -2516 575 -2296 609
rect -1928 575 -1708 609
rect -1340 575 -1120 609
rect -752 575 -532 609
rect -164 575 56 609
rect 424 575 644 609
rect 1012 575 1232 609
rect 1600 575 1820 609
rect 2188 575 2408 609
rect 2776 575 2996 609
rect 3364 575 3584 609
rect 3952 575 4172 609
rect 4540 575 4760 609
rect 5128 575 5348 609
rect 5716 575 5936 609
rect 6304 575 6524 609
rect 6892 575 7112 609
rect 7480 575 7700 609
rect 8068 575 8288 609
rect 8656 575 8876 609
rect 9244 575 9464 609
rect 9832 575 10052 609
rect 10420 575 10640 609
rect 11008 575 11228 609
rect 11596 575 11816 609
rect 12184 575 12404 609
rect 12772 575 12992 609
rect 13360 575 13580 609
rect 13948 575 14168 609
rect 14536 575 14756 609
rect 15124 575 15344 609
rect 15712 575 15932 609
rect 16300 575 16520 609
rect 16888 575 17108 609
rect 17476 575 17696 609
rect 18064 575 18284 609
rect 18652 575 18872 609
rect 19240 575 19460 609
rect 19828 575 20048 609
rect 20416 575 20636 609
rect 21004 575 21224 609
rect 21592 575 21608 609
rect -6428 537 5332 575
rect 5732 537 5920 575
rect 6320 574 6508 575
rect 6320 537 6508 538
rect 6908 537 7096 575
rect 7496 537 7684 575
rect 8084 537 8272 575
rect 8672 574 8860 575
rect 8672 537 8860 538
rect 9260 537 9448 575
rect 9848 537 21608 575
rect -6428 503 -6412 537
rect -6044 503 -5824 537
rect -5456 503 -5236 537
rect -4868 503 -4648 537
rect -4280 503 -4060 537
rect -3692 503 -3472 537
rect -3104 503 -2884 537
rect -2516 503 -2296 537
rect -1928 503 -1708 537
rect -1340 503 -1120 537
rect -752 503 -532 537
rect -164 503 56 537
rect 424 503 644 537
rect 1012 503 1232 537
rect 1600 503 1820 537
rect 2188 503 2408 537
rect 2776 503 2996 537
rect 3364 503 3584 537
rect 3952 503 4172 537
rect 4540 503 4760 537
rect 5128 503 5348 537
rect 5716 503 5936 537
rect 6304 503 6524 537
rect 6892 503 7112 537
rect 7480 503 7700 537
rect 8068 503 8288 537
rect 8656 503 8876 537
rect 9244 503 9464 537
rect 9832 503 10052 537
rect 10420 503 10640 537
rect 11008 503 11228 537
rect 11596 503 11816 537
rect 12184 503 12404 537
rect 12772 503 12992 537
rect 13360 503 13580 537
rect 13948 503 14168 537
rect 14536 503 14756 537
rect 15124 503 15344 537
rect 15712 503 15932 537
rect 16300 503 16520 537
rect 16888 503 17108 537
rect 17476 503 17696 537
rect 18064 503 18284 537
rect 18652 503 18872 537
rect 19240 503 19460 537
rect 19828 503 20048 537
rect 20416 503 20636 537
rect 21004 503 21224 537
rect 21592 503 21608 537
rect -6428 502 5332 503
rect 5732 502 5920 503
rect 6320 502 6508 503
rect 6908 502 7096 503
rect 7496 502 7684 503
rect 8084 502 8272 503
rect 8672 502 8860 503
rect 9260 502 9448 503
rect 9848 502 21608 503
rect -6474 444 -6440 460
rect -6474 -348 -6440 -332
rect -6016 444 -5982 460
rect -6016 -348 -5982 -332
rect -5886 444 -5852 460
rect -5886 -348 -5852 -332
rect -5428 444 -5394 460
rect -5428 -348 -5394 -332
rect -5298 444 -5264 460
rect -5298 -348 -5264 -332
rect -4840 444 -4806 460
rect -4840 -348 -4806 -332
rect -4710 444 -4676 460
rect -4710 -348 -4676 -332
rect -4252 444 -4218 460
rect -4252 -348 -4218 -332
rect -4122 444 -4088 460
rect -4122 -348 -4088 -332
rect -3664 444 -3630 460
rect -3664 -348 -3630 -332
rect -3534 444 -3500 460
rect -3534 -348 -3500 -332
rect -3076 444 -3042 460
rect -3076 -348 -3042 -332
rect -2946 444 -2912 460
rect -2946 -348 -2912 -332
rect -2488 444 -2454 460
rect -2488 -348 -2454 -332
rect -2358 444 -2324 460
rect -2358 -348 -2324 -332
rect -1900 444 -1866 460
rect -1900 -348 -1866 -332
rect -1770 444 -1736 460
rect -1770 -348 -1736 -332
rect -1312 444 -1278 460
rect -1312 -348 -1278 -332
rect -1182 444 -1148 460
rect -1182 -348 -1148 -332
rect -724 444 -690 460
rect -724 -348 -690 -332
rect -594 444 -560 460
rect -594 -348 -560 -332
rect -136 444 -102 460
rect -136 -348 -102 -332
rect -6 444 28 460
rect -6 -348 28 -332
rect 452 444 486 460
rect 452 -348 486 -332
rect 582 444 616 460
rect 582 -348 616 -332
rect 1040 444 1074 460
rect 1040 -348 1074 -332
rect 1170 444 1204 460
rect 1170 -348 1204 -332
rect 1628 444 1662 460
rect 1628 -348 1662 -332
rect 1758 444 1792 460
rect 1758 -348 1792 -332
rect 2216 444 2250 460
rect 2216 -348 2250 -332
rect 2346 444 2380 460
rect 2346 -348 2380 -332
rect 2804 444 2838 460
rect 2804 -348 2838 -332
rect 2934 444 2968 460
rect 2934 -348 2968 -332
rect 3392 444 3426 460
rect 3392 -348 3426 -332
rect 3522 444 3556 460
rect 3522 -348 3556 -332
rect 3980 444 4014 460
rect 3980 -348 4014 -332
rect 4110 444 4144 460
rect 4110 -348 4144 -332
rect 4568 444 4602 460
rect 4568 -348 4602 -332
rect 4698 444 4732 460
rect 4698 -348 4732 -332
rect 5156 444 5190 460
rect 5156 -348 5190 -332
rect 5286 444 5320 502
rect 5286 -348 5320 -332
rect 5744 444 5778 460
rect 5744 -348 5778 -332
rect 5874 444 5908 460
rect 5874 -348 5908 -332
rect 6332 444 6366 460
rect 6332 -348 6366 -332
rect 6462 444 6496 460
rect 6462 -348 6496 -332
rect 6920 444 6954 460
rect 6920 -348 6954 -332
rect 7050 444 7084 460
rect 7050 -348 7084 -332
rect 7508 444 7672 502
rect 7542 -332 7638 444
rect 7508 -348 7672 -332
rect 8096 444 8130 460
rect 8096 -348 8130 -332
rect 8226 444 8260 460
rect 8226 -348 8260 -332
rect 8684 444 8718 460
rect 8684 -348 8718 -332
rect 8814 444 8848 460
rect 8814 -348 8848 -332
rect 9272 444 9306 460
rect 9272 -348 9306 -332
rect 9402 444 9436 460
rect 9402 -348 9436 -332
rect 9860 444 9894 502
rect 9860 -348 9894 -332
rect 9990 444 10024 460
rect 9990 -348 10024 -332
rect 10448 444 10482 460
rect 10448 -348 10482 -332
rect 10578 444 10612 460
rect 10578 -348 10612 -332
rect 11036 444 11070 460
rect 11036 -348 11070 -332
rect 11166 444 11200 460
rect 11166 -348 11200 -332
rect 11624 444 11658 460
rect 11624 -348 11658 -332
rect 11754 444 11788 460
rect 11754 -348 11788 -332
rect 12212 444 12246 460
rect 12212 -348 12246 -332
rect 12342 444 12376 460
rect 12342 -348 12376 -332
rect 12800 444 12834 460
rect 12800 -348 12834 -332
rect 12930 444 12964 460
rect 12930 -348 12964 -332
rect 13388 444 13422 460
rect 13388 -348 13422 -332
rect 13518 444 13552 460
rect 13518 -348 13552 -332
rect 13976 444 14010 460
rect 13976 -348 14010 -332
rect 14106 444 14140 460
rect 14106 -348 14140 -332
rect 14564 444 14598 460
rect 14564 -348 14598 -332
rect 14694 444 14728 460
rect 14694 -348 14728 -332
rect 15152 444 15186 460
rect 15152 -348 15186 -332
rect 15282 444 15316 460
rect 15282 -348 15316 -332
rect 15740 444 15774 460
rect 15740 -348 15774 -332
rect 15870 444 15904 460
rect 15870 -348 15904 -332
rect 16328 444 16362 460
rect 16328 -348 16362 -332
rect 16458 444 16492 460
rect 16458 -348 16492 -332
rect 16916 444 16950 460
rect 16916 -348 16950 -332
rect 17046 444 17080 460
rect 17046 -348 17080 -332
rect 17504 444 17538 460
rect 17504 -348 17538 -332
rect 17634 444 17668 460
rect 17634 -348 17668 -332
rect 18092 444 18126 460
rect 18092 -348 18126 -332
rect 18222 444 18256 460
rect 18222 -348 18256 -332
rect 18680 444 18714 460
rect 18680 -348 18714 -332
rect 18810 444 18844 460
rect 18810 -348 18844 -332
rect 19268 444 19302 460
rect 19268 -348 19302 -332
rect 19398 444 19432 460
rect 19398 -348 19432 -332
rect 19856 444 19890 460
rect 19856 -348 19890 -332
rect 19986 444 20020 460
rect 19986 -348 20020 -332
rect 20444 444 20478 460
rect 20444 -348 20478 -332
rect 20574 444 20608 460
rect 20574 -348 20608 -332
rect 21032 444 21066 460
rect 21032 -348 21066 -332
rect 21162 444 21196 460
rect 21162 -348 21196 -332
rect 21620 444 21654 460
rect 21620 -348 21654 -332
rect 5286 -390 5332 -348
rect -6428 -391 5332 -390
rect 5732 -391 5920 -390
rect 6320 -391 6508 -390
rect 6908 -391 7096 -390
rect 7496 -391 7684 -348
rect 9848 -390 9894 -348
rect 8084 -391 8272 -390
rect 8672 -391 8860 -390
rect 9260 -391 9448 -390
rect 9848 -391 21608 -390
rect -6428 -425 -6412 -391
rect -6044 -425 -5824 -391
rect -5456 -425 -5236 -391
rect -4868 -425 -4648 -391
rect -4280 -425 -4060 -391
rect -3692 -425 -3472 -391
rect -3104 -425 -2884 -391
rect -2516 -425 -2296 -391
rect -1928 -425 -1708 -391
rect -1340 -425 -1120 -391
rect -752 -425 -532 -391
rect -164 -425 56 -391
rect 424 -425 644 -391
rect 1012 -425 1232 -391
rect 1600 -425 1820 -391
rect 2188 -425 2408 -391
rect 2776 -425 2996 -391
rect 3364 -425 3584 -391
rect 3952 -425 4172 -391
rect 4540 -425 4760 -391
rect 5128 -425 5348 -391
rect 5716 -425 5936 -391
rect 6304 -425 6524 -391
rect 6892 -425 7112 -391
rect 7480 -425 7700 -391
rect 8068 -425 8288 -391
rect 8656 -425 8876 -391
rect 9244 -425 9464 -391
rect 9832 -425 10052 -391
rect 10420 -425 10640 -391
rect 11008 -425 11228 -391
rect 11596 -425 11816 -391
rect 12184 -425 12404 -391
rect 12772 -425 12992 -391
rect 13360 -425 13580 -391
rect 13948 -425 14168 -391
rect 14536 -425 14756 -391
rect 15124 -425 15344 -391
rect 15712 -425 15932 -391
rect 16300 -425 16520 -391
rect 16888 -425 17108 -391
rect 17476 -425 17696 -391
rect 18064 -425 18284 -391
rect 18652 -425 18872 -391
rect 19240 -425 19460 -391
rect 19828 -425 20048 -391
rect 20416 -425 20636 -391
rect 21004 -425 21224 -391
rect 21592 -425 21608 -391
rect -6428 -426 5332 -425
rect 5732 -426 5920 -425
rect 6320 -426 6508 -425
rect 6908 -426 7096 -425
rect 7496 -426 7684 -425
rect 8084 -426 8272 -425
rect 8672 -426 8860 -425
rect 9260 -426 9448 -425
rect 9848 -426 21608 -425
rect -6820 -742 -6786 -722
rect 21966 -742 22000 -688
rect -6820 -776 -6702 -742
rect 21912 -776 22000 -742
rect 6882 -804 6908 -776
rect 7096 -804 7126 -776
rect 6882 -1486 7126 -804
rect 8056 -804 8084 -776
rect 8272 -804 8300 -776
rect 8056 -1486 8300 -804
rect 6192 -1520 6226 -1486
rect 8954 -1520 8988 -1486
rect 6624 -1952 6640 -1820
rect 6678 -1952 6906 -1820
rect 6944 -1952 6962 -1820
rect 7156 -1952 7172 -1820
rect 7210 -1952 7438 -1820
rect 7476 -1952 7494 -1820
rect 7688 -1952 7704 -1820
rect 7742 -1952 7970 -1820
rect 8008 -1952 8026 -1820
rect 8220 -1952 8236 -1820
rect 8274 -1952 8502 -1820
rect 8540 -1952 8558 -1820
rect 6578 -2002 6612 -1986
rect 6578 -2794 6612 -2778
rect 6706 -2002 6740 -1986
rect 6706 -2794 6740 -2778
rect 6844 -2002 6878 -1986
rect 6844 -2794 6878 -2778
rect 6972 -2002 7006 -1986
rect 6972 -2794 7006 -2778
rect 7110 -2002 7144 -1986
rect 7110 -2794 7144 -2778
rect 7238 -2002 7272 -1986
rect 7238 -2794 7272 -2778
rect 7376 -2002 7410 -1986
rect 7376 -2794 7410 -2778
rect 7504 -2002 7538 -1986
rect 7504 -2794 7538 -2778
rect 7642 -2002 7676 -1986
rect 7642 -2794 7676 -2778
rect 7770 -2002 7804 -1986
rect 7770 -2794 7804 -2778
rect 7908 -2002 7942 -1986
rect 7908 -2794 7942 -2778
rect 8036 -2002 8070 -1986
rect 8036 -2794 8070 -2778
rect 8174 -2002 8208 -1986
rect 8174 -2794 8208 -2778
rect 8302 -2002 8336 -1986
rect 8302 -2794 8336 -2778
rect 8440 -2002 8474 -1986
rect 8440 -2794 8474 -2778
rect 8568 -2002 8602 -1986
rect 8568 -2794 8602 -2778
rect 6624 -2962 6640 -2830
rect 6678 -2962 6906 -2830
rect 6944 -2962 6962 -2830
rect 7156 -2962 7172 -2830
rect 7210 -2962 7438 -2830
rect 7476 -2962 7494 -2830
rect 7688 -2962 7704 -2830
rect 7742 -2962 7970 -2830
rect 8008 -2962 8026 -2830
rect 8220 -2962 8236 -2830
rect 8274 -2962 8502 -2830
rect 8540 -2962 8558 -2830
rect 6578 -3012 6612 -2996
rect 6578 -3804 6612 -3788
rect 6706 -3012 6740 -2996
rect 6706 -3804 6740 -3788
rect 6844 -3012 6878 -2996
rect 6844 -3804 6878 -3788
rect 6972 -3012 7006 -2996
rect 6972 -3804 7006 -3788
rect 7110 -3012 7144 -2996
rect 7110 -3804 7144 -3788
rect 7238 -3012 7272 -2996
rect 7238 -3804 7272 -3788
rect 7376 -3012 7410 -2996
rect 7376 -3804 7410 -3788
rect 7504 -3012 7538 -2996
rect 7504 -3804 7538 -3788
rect 7642 -3012 7676 -2996
rect 7642 -3804 7676 -3788
rect 7770 -3012 7804 -2996
rect 7770 -3804 7804 -3788
rect 7908 -3012 7942 -2996
rect 7908 -3804 7942 -3788
rect 8036 -3012 8070 -2996
rect 8036 -3804 8070 -3788
rect 8174 -3012 8208 -2996
rect 8174 -3804 8208 -3788
rect 8302 -3012 8336 -2996
rect 8302 -3804 8336 -3788
rect 8440 -3012 8474 -2996
rect 8440 -3804 8474 -3788
rect 8568 -3012 8602 -2996
rect 8568 -3804 8602 -3788
rect 6624 -3972 6640 -3840
rect 6678 -3972 6906 -3840
rect 6944 -3972 6962 -3840
rect 7156 -3972 7172 -3840
rect 7210 -3972 7438 -3840
rect 7476 -3972 7494 -3840
rect 7688 -3972 7704 -3840
rect 7742 -3972 7970 -3840
rect 8008 -3972 8026 -3840
rect 8220 -3972 8236 -3840
rect 8274 -3972 8502 -3840
rect 8540 -3972 8558 -3840
rect 6578 -4022 6612 -4006
rect 6578 -4814 6612 -4798
rect 6706 -4022 6740 -4006
rect 6706 -4814 6740 -4798
rect 6844 -4022 6878 -4006
rect 6844 -4814 6878 -4798
rect 6972 -4022 7006 -4006
rect 6972 -4814 7006 -4798
rect 7110 -4022 7144 -4006
rect 7110 -4814 7144 -4798
rect 7238 -4022 7272 -4006
rect 7238 -4814 7272 -4798
rect 7376 -4022 7410 -4006
rect 7376 -4814 7410 -4798
rect 7504 -4022 7538 -4006
rect 7504 -4814 7538 -4798
rect 7642 -4022 7676 -4006
rect 7642 -4814 7676 -4798
rect 7770 -4022 7804 -4006
rect 7770 -4814 7804 -4798
rect 7908 -4022 7942 -4006
rect 7908 -4814 7942 -4798
rect 8036 -4022 8070 -4006
rect 8036 -4814 8070 -4798
rect 8174 -4022 8208 -4006
rect 8174 -4814 8208 -4798
rect 8302 -4022 8336 -4006
rect 8302 -4814 8336 -4798
rect 8440 -4022 8474 -4006
rect 8440 -4814 8474 -4798
rect 8568 -4022 8602 -4006
rect 8568 -4814 8602 -4798
rect 6624 -4982 6640 -4850
rect 6678 -4982 6906 -4850
rect 6944 -4982 6962 -4850
rect 7156 -4982 7172 -4850
rect 7210 -4982 7438 -4850
rect 7476 -4982 7494 -4850
rect 7688 -4982 7704 -4850
rect 7742 -4982 7970 -4850
rect 8008 -4982 8026 -4850
rect 8220 -4982 8236 -4850
rect 8274 -4982 8502 -4850
rect 8540 -4982 8558 -4850
rect 13613 -3401 13709 -3367
rect 13847 -3401 13943 -3367
rect 13613 -3463 13647 -3401
rect 13909 -3463 13943 -3401
rect 13613 -5017 13647 -4955
rect 13943 -4122 14206 -4102
rect 13943 -4582 14048 -4122
rect 14188 -4582 14206 -4122
rect 13943 -4604 14206 -4582
rect 13909 -5017 13943 -4955
rect 13613 -5051 13709 -5017
rect 13847 -5051 13943 -5017
rect 6192 -5316 6226 -5282
rect 8954 -5316 8988 -5282
rect 6804 -5712 6950 -5678
rect 8160 -5712 8378 -5678
rect 7150 -6018 8032 -6012
rect 7150 -6144 7212 -6018
rect 7250 -6144 7452 -6018
rect 7490 -6144 7692 -6018
rect 7730 -6144 7932 -6018
rect 7970 -6144 8032 -6018
rect 7150 -6194 7184 -6144
rect 7150 -6820 7184 -6770
rect 7278 -6194 7312 -6178
rect 7278 -6786 7312 -6770
rect 7390 -6194 7424 -6178
rect 7390 -6786 7424 -6770
rect 7518 -6194 7552 -6178
rect 7518 -6786 7552 -6770
rect 7630 -6194 7664 -6178
rect 7630 -6786 7664 -6770
rect 7758 -6194 7792 -6178
rect 7758 -6786 7792 -6770
rect 7870 -6194 7904 -6178
rect 7870 -6786 7904 -6770
rect 7998 -6194 8032 -6144
rect 7998 -6820 8032 -6770
rect 7150 -6952 7212 -6820
rect 7250 -6952 7452 -6820
rect 7490 -6952 7692 -6820
rect 7730 -6952 7932 -6820
rect 7970 -6952 8032 -6820
rect 7150 -7002 7184 -6952
rect 7150 -7628 7184 -7578
rect 7278 -7002 7312 -6986
rect 7278 -7594 7312 -7578
rect 7390 -7002 7424 -6986
rect 7390 -7594 7424 -7578
rect 7518 -7002 7552 -6986
rect 7518 -7594 7552 -7578
rect 7630 -7002 7664 -6986
rect 7630 -7594 7664 -7578
rect 7758 -7002 7792 -6986
rect 7758 -7594 7792 -7578
rect 7870 -7002 7904 -6986
rect 7870 -7594 7904 -7578
rect 7998 -7002 8032 -6952
rect 7998 -7628 8032 -7578
rect 7150 -7760 7212 -7628
rect 7250 -7760 7452 -7628
rect 7490 -7760 7692 -7628
rect 7730 -7760 7932 -7628
rect 7970 -7760 8032 -7628
rect 6804 -8094 6902 -8060
rect 8254 -8094 8378 -8060
<< viali >>
rect 2976 7056 3086 7090
rect 3456 7056 3566 7090
rect 3936 7056 4046 7090
rect 4416 7056 4526 7090
rect 4896 7056 5006 7090
rect 5376 7056 5486 7090
rect 5856 7056 5966 7090
rect 6336 7056 6446 7090
rect 6816 7056 6926 7090
rect 7296 7056 7406 7090
rect 7776 7056 7886 7090
rect 8256 7056 8366 7090
rect 8736 7056 8846 7090
rect 9216 7056 9326 7090
rect 9696 7056 9806 7090
rect 10176 7056 10286 7090
rect 10656 7056 10766 7090
rect 11136 7056 11246 7090
rect 11616 7056 11726 7090
rect 12096 7056 12206 7090
rect 2976 7018 3086 7056
rect 3456 7018 3566 7056
rect 3936 7018 4046 7056
rect 4416 7018 4526 7056
rect 4896 7018 5006 7056
rect 5376 7018 5486 7056
rect 5856 7018 5966 7056
rect 6336 7018 6446 7056
rect 6816 7018 6926 7056
rect 7296 7018 7406 7056
rect 7776 7018 7886 7056
rect 8256 7018 8366 7056
rect 8736 7018 8846 7056
rect 9216 7018 9326 7056
rect 9696 7018 9806 7056
rect 10176 7018 10286 7056
rect 10656 7018 10766 7056
rect 11136 7018 11246 7056
rect 11616 7018 11726 7056
rect 12096 7018 12206 7056
rect 2892 6614 2930 6746
rect 3132 6614 3170 6746
rect 3372 6614 3410 6746
rect 3612 6614 3650 6746
rect 3852 6614 3890 6746
rect 4092 6614 4130 6746
rect 4332 6614 4370 6746
rect 4572 6614 4610 6746
rect 4812 6614 4850 6746
rect 5052 6614 5090 6746
rect 5292 6614 5330 6746
rect 5532 6614 5570 6746
rect 5772 6614 5810 6746
rect 6012 6614 6050 6746
rect 6252 6614 6290 6746
rect 6492 6614 6530 6746
rect 6732 6614 6770 6746
rect 6972 6614 7010 6746
rect 7212 6614 7250 6746
rect 7452 6614 7490 6746
rect 7692 6614 7730 6746
rect 7932 6614 7970 6746
rect 8172 6614 8210 6746
rect 8412 6614 8450 6746
rect 8652 6614 8690 6746
rect 8892 6614 8930 6746
rect 9132 6614 9170 6746
rect 9372 6614 9410 6746
rect 9612 6614 9650 6746
rect 9852 6614 9890 6746
rect 10092 6614 10130 6746
rect 10332 6614 10370 6746
rect 10572 6614 10610 6746
rect 10812 6614 10850 6746
rect 11052 6614 11090 6746
rect 11292 6614 11330 6746
rect 11532 6614 11570 6746
rect 11772 6614 11810 6746
rect 12012 6614 12050 6746
rect 12252 6614 12290 6746
rect 2830 5988 2864 6564
rect 2958 5988 2992 6564
rect 3070 5988 3104 6564
rect 3198 5988 3232 6564
rect 3310 5988 3344 6564
rect 3438 5988 3472 6564
rect 3550 5988 3584 6564
rect 3678 5988 3712 6564
rect 3790 5988 3824 6564
rect 3918 5988 3952 6564
rect 4030 5988 4064 6564
rect 4158 5988 4192 6564
rect 4270 5988 4304 6564
rect 4398 5988 4432 6564
rect 4510 5988 4544 6564
rect 4638 5988 4672 6564
rect 4750 5988 4784 6564
rect 4878 5988 4912 6564
rect 4990 5988 5024 6564
rect 5118 5988 5152 6564
rect 5230 5988 5264 6564
rect 5358 5988 5392 6564
rect 5470 5988 5504 6564
rect 5598 5988 5632 6564
rect 5710 5988 5744 6564
rect 5838 5988 5872 6564
rect 5950 5988 5984 6564
rect 6078 5988 6112 6564
rect 6190 5988 6224 6564
rect 6318 5988 6352 6564
rect 6430 5988 6464 6564
rect 6558 5988 6592 6564
rect 6670 5988 6704 6564
rect 6798 5988 6832 6564
rect 6910 5988 6944 6564
rect 7038 5988 7072 6564
rect 7150 5988 7184 6564
rect 7278 5988 7312 6564
rect 7390 5988 7424 6564
rect 7518 5988 7552 6564
rect 7630 5988 7664 6564
rect 7758 5988 7792 6564
rect 7870 5988 7904 6564
rect 7998 5988 8032 6564
rect 8110 5988 8144 6564
rect 8238 5988 8272 6564
rect 8350 5988 8384 6564
rect 8478 5988 8512 6564
rect 8590 5988 8624 6564
rect 8718 5988 8752 6564
rect 8830 5988 8864 6564
rect 8958 5988 8992 6564
rect 9070 5988 9104 6564
rect 9198 5988 9232 6564
rect 9310 5988 9344 6564
rect 9438 5988 9472 6564
rect 9550 5988 9584 6564
rect 9678 5988 9712 6564
rect 9790 5988 9824 6564
rect 9918 5988 9952 6564
rect 10030 5988 10064 6564
rect 10158 5988 10192 6564
rect 10270 5988 10304 6564
rect 10398 5988 10432 6564
rect 10510 5988 10544 6564
rect 10638 5988 10672 6564
rect 10750 5988 10784 6564
rect 10878 5988 10912 6564
rect 10990 5988 11024 6564
rect 11118 5988 11152 6564
rect 11230 5988 11264 6564
rect 11358 5988 11392 6564
rect 11470 5988 11504 6564
rect 11598 5988 11632 6564
rect 11710 5988 11744 6564
rect 11838 5988 11872 6564
rect 11950 5988 11984 6564
rect 12078 5988 12112 6564
rect 12190 5988 12224 6564
rect 12318 5988 12352 6564
rect 2892 5806 2930 5938
rect 3132 5806 3170 5938
rect 3372 5806 3410 5938
rect 3612 5806 3650 5938
rect 3852 5806 3890 5938
rect 4092 5806 4130 5938
rect 4332 5806 4370 5938
rect 4572 5806 4610 5938
rect 4812 5806 4850 5938
rect 5052 5806 5090 5938
rect 5292 5806 5330 5938
rect 5532 5806 5570 5938
rect 5772 5806 5810 5938
rect 6012 5806 6050 5938
rect 6252 5806 6290 5938
rect 6492 5806 6530 5938
rect 6732 5806 6770 5938
rect 6972 5806 7010 5938
rect 7212 5806 7250 5938
rect 7452 5806 7490 5938
rect 7692 5806 7730 5938
rect 7932 5806 7970 5938
rect 8172 5806 8210 5938
rect 8412 5806 8450 5938
rect 8652 5806 8690 5938
rect 8892 5806 8930 5938
rect 9132 5806 9170 5938
rect 9372 5806 9410 5938
rect 9612 5806 9650 5938
rect 9852 5806 9890 5938
rect 10092 5806 10130 5938
rect 10332 5806 10370 5938
rect 10572 5806 10610 5938
rect 10812 5806 10850 5938
rect 11052 5806 11090 5938
rect 11292 5806 11330 5938
rect 11532 5806 11570 5938
rect 11772 5806 11810 5938
rect 12012 5806 12050 5938
rect 12252 5806 12290 5938
rect 2830 5180 2864 5756
rect 2958 5180 2992 5756
rect 3070 5180 3104 5756
rect 3198 5180 3232 5756
rect 3310 5180 3344 5756
rect 3438 5180 3472 5756
rect 3550 5180 3584 5756
rect 3678 5180 3712 5756
rect 3790 5180 3824 5756
rect 3918 5180 3952 5756
rect 4030 5180 4064 5756
rect 4158 5180 4192 5756
rect 4270 5180 4304 5756
rect 4398 5180 4432 5756
rect 4510 5180 4544 5756
rect 4638 5180 4672 5756
rect 4750 5180 4784 5756
rect 4878 5180 4912 5756
rect 4990 5180 5024 5756
rect 5118 5180 5152 5756
rect 5230 5180 5264 5756
rect 5358 5180 5392 5756
rect 5470 5180 5504 5756
rect 5598 5180 5632 5756
rect 5710 5180 5744 5756
rect 5838 5180 5872 5756
rect 5950 5180 5984 5756
rect 6078 5180 6112 5756
rect 6190 5180 6224 5756
rect 6318 5180 6352 5756
rect 6430 5180 6464 5756
rect 6558 5180 6592 5756
rect 6670 5180 6704 5756
rect 6798 5180 6832 5756
rect 6910 5180 6944 5756
rect 7038 5180 7072 5756
rect 7150 5180 7184 5756
rect 7278 5180 7312 5756
rect 7390 5180 7424 5756
rect 7518 5180 7552 5756
rect 7630 5180 7664 5756
rect 7758 5180 7792 5756
rect 7870 5180 7904 5756
rect 7998 5180 8032 5756
rect 8110 5180 8144 5756
rect 8238 5180 8272 5756
rect 8350 5180 8384 5756
rect 8478 5180 8512 5756
rect 8590 5180 8624 5756
rect 8718 5180 8752 5756
rect 8830 5180 8864 5756
rect 8958 5180 8992 5756
rect 9070 5180 9104 5756
rect 9198 5180 9232 5756
rect 9310 5180 9344 5756
rect 9438 5180 9472 5756
rect 9550 5180 9584 5756
rect 9678 5180 9712 5756
rect 9790 5180 9824 5756
rect 9918 5180 9952 5756
rect 10030 5180 10064 5756
rect 10158 5180 10192 5756
rect 10270 5180 10304 5756
rect 10398 5180 10432 5756
rect 10510 5180 10544 5756
rect 10638 5180 10672 5756
rect 10750 5180 10784 5756
rect 10878 5180 10912 5756
rect 10990 5180 11024 5756
rect 11118 5180 11152 5756
rect 11230 5180 11264 5756
rect 11358 5180 11392 5756
rect 11470 5180 11504 5756
rect 11598 5180 11632 5756
rect 11710 5180 11744 5756
rect 11838 5180 11872 5756
rect 11950 5180 11984 5756
rect 12078 5180 12112 5756
rect 12190 5180 12224 5756
rect 12318 5180 12352 5756
rect 2892 4998 2930 5130
rect 3132 4998 3170 5130
rect 3372 4998 3410 5130
rect 3612 4998 3650 5130
rect 3852 4998 3890 5130
rect 4092 4998 4130 5130
rect 4332 4998 4370 5130
rect 4572 4998 4610 5130
rect 4812 4998 4850 5130
rect 5052 4998 5090 5130
rect 5292 4998 5330 5130
rect 5532 4998 5570 5130
rect 5772 4998 5810 5130
rect 6012 4998 6050 5130
rect 6252 4998 6290 5130
rect 6492 4998 6530 5130
rect 6732 4998 6770 5130
rect 6972 4998 7010 5130
rect 7212 4998 7250 5130
rect 7452 4998 7490 5130
rect 7692 4998 7730 5130
rect 7932 4998 7970 5130
rect 8172 4998 8210 5130
rect 8412 4998 8450 5130
rect 8652 4998 8690 5130
rect 8892 4998 8930 5130
rect 9132 4998 9170 5130
rect 9372 4998 9410 5130
rect 9612 4998 9650 5130
rect 9852 4998 9890 5130
rect 10092 4998 10130 5130
rect 10332 4998 10370 5130
rect 10572 4998 10610 5130
rect 10812 4998 10850 5130
rect 11052 4998 11090 5130
rect 11292 4998 11330 5130
rect 11532 4998 11570 5130
rect 11772 4998 11810 5130
rect 12012 4998 12050 5130
rect 12252 4998 12290 5130
rect -6412 2503 -6044 2537
rect -5824 2503 -5456 2537
rect -5236 2503 -4868 2537
rect -4648 2503 -4280 2537
rect -4060 2503 -3692 2537
rect -3472 2503 -3104 2537
rect -2884 2503 -2516 2537
rect -2296 2503 -1928 2537
rect -1708 2503 -1340 2537
rect -1120 2503 -752 2537
rect -532 2503 -164 2537
rect 56 2503 424 2537
rect 644 2503 1012 2537
rect 1232 2503 1600 2537
rect 1820 2503 2188 2537
rect 2408 2503 2776 2537
rect 2996 2503 3364 2537
rect 3584 2503 3952 2537
rect 4172 2503 4540 2537
rect 4760 2503 5128 2537
rect 5348 2503 5716 2537
rect 5936 2503 6304 2537
rect 6524 2503 6892 2537
rect 7112 2503 7480 2537
rect 7700 2503 8068 2537
rect 8288 2503 8656 2537
rect 8876 2503 9244 2537
rect 9464 2503 9832 2537
rect 10052 2503 10420 2537
rect 10640 2503 11008 2537
rect 11228 2503 11596 2537
rect 11816 2503 12184 2537
rect 12404 2503 12772 2537
rect 12992 2503 13360 2537
rect 13580 2503 13948 2537
rect 14168 2503 14536 2537
rect 14756 2503 15124 2537
rect 15344 2503 15712 2537
rect 15932 2503 16300 2537
rect 16520 2503 16888 2537
rect 17108 2503 17476 2537
rect 17696 2503 18064 2537
rect 18284 2503 18652 2537
rect 18872 2503 19240 2537
rect 19460 2503 19828 2537
rect 20048 2503 20416 2537
rect 20636 2503 21004 2537
rect 21224 2503 21592 2537
rect -6474 1668 -6440 2444
rect -6016 1668 -5982 2444
rect -5886 1668 -5852 2444
rect -5428 1668 -5394 2444
rect -5298 1668 -5264 2444
rect -4840 1668 -4806 2444
rect -4710 1668 -4676 2444
rect -4252 1668 -4218 2444
rect -4122 1668 -4088 2444
rect -3664 1668 -3630 2444
rect -3534 1668 -3500 2444
rect -3076 1668 -3042 2444
rect -2946 1668 -2912 2444
rect -2488 1668 -2454 2444
rect -2358 1668 -2324 2444
rect -1900 1668 -1866 2444
rect -1770 1668 -1736 2444
rect -1312 1668 -1278 2444
rect -1182 1668 -1148 2444
rect -724 1668 -690 2444
rect -594 1668 -560 2444
rect -136 1668 -102 2444
rect -6 1668 28 2444
rect 452 1668 486 2444
rect 582 1668 616 2444
rect 1040 1668 1074 2444
rect 1170 1668 1204 2444
rect 1628 1668 1662 2444
rect 1758 1668 1792 2444
rect 2216 1668 2250 2444
rect 2346 1668 2380 2444
rect 2804 1668 2838 2444
rect 2934 1668 2968 2444
rect 3392 1668 3426 2444
rect 3522 1668 3556 2444
rect 3980 1668 4014 2444
rect 4110 1668 4144 2444
rect 4568 1668 4602 2444
rect 4698 1668 4732 2444
rect 5156 1668 5190 2444
rect 5286 1668 5320 2444
rect 5744 1668 5778 2444
rect 5874 1668 5908 2444
rect 6332 1668 6366 2444
rect 6462 1668 6496 2444
rect 6920 1668 6954 2444
rect 7050 1668 7084 2444
rect 7508 1668 7542 2444
rect 7638 1668 7672 2444
rect 8096 1668 8130 2444
rect 8226 1668 8260 2444
rect 8684 1668 8718 2444
rect 8814 1668 8848 2444
rect 9272 1668 9306 2444
rect 9402 1668 9436 2444
rect 9860 1668 9894 2444
rect 9990 1668 10024 2444
rect 10448 1668 10482 2444
rect 10578 1668 10612 2444
rect 11036 1668 11070 2444
rect 11166 1668 11200 2444
rect 11624 1668 11658 2444
rect 11754 1668 11788 2444
rect 12212 1668 12246 2444
rect 12342 1668 12376 2444
rect 12800 1668 12834 2444
rect 12930 1668 12964 2444
rect 13388 1668 13422 2444
rect 13518 1668 13552 2444
rect 13976 1668 14010 2444
rect 14106 1668 14140 2444
rect 14564 1668 14598 2444
rect 14694 1668 14728 2444
rect 15152 1668 15186 2444
rect 15282 1668 15316 2444
rect 15740 1668 15774 2444
rect 15870 1668 15904 2444
rect 16328 1668 16362 2444
rect 16458 1668 16492 2444
rect 16916 1668 16950 2444
rect 17046 1668 17080 2444
rect 17504 1668 17538 2444
rect 17634 1668 17668 2444
rect 18092 1668 18126 2444
rect 18222 1668 18256 2444
rect 18680 1668 18714 2444
rect 18810 1668 18844 2444
rect 19268 1668 19302 2444
rect 19398 1668 19432 2444
rect 19856 1668 19890 2444
rect 19986 1668 20020 2444
rect 20444 1668 20478 2444
rect 20574 1668 20608 2444
rect 21032 1668 21066 2444
rect 21162 1668 21196 2444
rect 21620 1668 21654 2444
rect -6412 1575 -6044 1609
rect -5824 1575 -5456 1609
rect -5236 1575 -4868 1609
rect -4648 1575 -4280 1609
rect -4060 1575 -3692 1609
rect -3472 1575 -3104 1609
rect -2884 1575 -2516 1609
rect -2296 1575 -1928 1609
rect -1708 1575 -1340 1609
rect -1120 1575 -752 1609
rect -532 1575 -164 1609
rect 56 1575 424 1609
rect 644 1575 1012 1609
rect 1232 1575 1600 1609
rect 1820 1575 2188 1609
rect 2408 1575 2776 1609
rect 2996 1575 3364 1609
rect 3584 1575 3952 1609
rect 4172 1575 4540 1609
rect 4760 1575 5128 1609
rect 5348 1575 5716 1609
rect 5936 1575 6304 1609
rect 6524 1575 6892 1609
rect 7112 1575 7480 1609
rect 7700 1575 8068 1609
rect 8288 1575 8656 1609
rect 8876 1575 9244 1609
rect 9464 1575 9832 1609
rect 10052 1575 10420 1609
rect 10640 1575 11008 1609
rect 11228 1575 11596 1609
rect 11816 1575 12184 1609
rect 12404 1575 12772 1609
rect 12992 1575 13360 1609
rect 13580 1575 13948 1609
rect 14168 1575 14536 1609
rect 14756 1575 15124 1609
rect 15344 1575 15712 1609
rect 15932 1575 16300 1609
rect 16520 1575 16888 1609
rect 17108 1575 17476 1609
rect 17696 1575 18064 1609
rect 18284 1575 18652 1609
rect 18872 1575 19240 1609
rect 19460 1575 19828 1609
rect 20048 1575 20416 1609
rect 20636 1575 21004 1609
rect 21224 1575 21592 1609
rect -6412 1503 -6044 1537
rect -5824 1503 -5456 1537
rect -5236 1503 -4868 1537
rect -4648 1503 -4280 1537
rect -4060 1503 -3692 1537
rect -3472 1503 -3104 1537
rect -2884 1503 -2516 1537
rect -2296 1503 -1928 1537
rect -1708 1503 -1340 1537
rect -1120 1503 -752 1537
rect -532 1503 -164 1537
rect 56 1503 424 1537
rect 644 1503 1012 1537
rect 1232 1503 1600 1537
rect 1820 1503 2188 1537
rect 2408 1503 2776 1537
rect 2996 1503 3364 1537
rect 3584 1503 3952 1537
rect 4172 1503 4540 1537
rect 4760 1503 5128 1537
rect 5348 1503 5716 1537
rect 5936 1503 6304 1537
rect 6524 1503 6892 1537
rect 7112 1503 7480 1537
rect 7700 1503 8068 1537
rect 8288 1503 8656 1537
rect 8876 1503 9244 1537
rect 9464 1503 9832 1537
rect 10052 1503 10420 1537
rect 10640 1503 11008 1537
rect 11228 1503 11596 1537
rect 11816 1503 12184 1537
rect 12404 1503 12772 1537
rect 12992 1503 13360 1537
rect 13580 1503 13948 1537
rect 14168 1503 14536 1537
rect 14756 1503 15124 1537
rect 15344 1503 15712 1537
rect 15932 1503 16300 1537
rect 16520 1503 16888 1537
rect 17108 1503 17476 1537
rect 17696 1503 18064 1537
rect 18284 1503 18652 1537
rect 18872 1503 19240 1537
rect 19460 1503 19828 1537
rect 20048 1503 20416 1537
rect 20636 1503 21004 1537
rect 21224 1503 21592 1537
rect -6474 668 -6440 1444
rect -6016 668 -5982 1444
rect -5886 668 -5852 1444
rect -5428 668 -5394 1444
rect -5298 668 -5264 1444
rect -4840 668 -4806 1444
rect -4710 668 -4676 1444
rect -4252 668 -4218 1444
rect -4122 668 -4088 1444
rect -3664 668 -3630 1444
rect -3534 668 -3500 1444
rect -3076 668 -3042 1444
rect -2946 668 -2912 1444
rect -2488 668 -2454 1444
rect -2358 668 -2324 1444
rect -1900 668 -1866 1444
rect -1770 668 -1736 1444
rect -1312 668 -1278 1444
rect -1182 668 -1148 1444
rect -724 668 -690 1444
rect -594 668 -560 1444
rect -136 668 -102 1444
rect -6 668 28 1444
rect 452 668 486 1444
rect 582 668 616 1444
rect 1040 668 1074 1444
rect 1170 668 1204 1444
rect 1628 668 1662 1444
rect 1758 668 1792 1444
rect 2216 668 2250 1444
rect 2346 668 2380 1444
rect 2804 668 2838 1444
rect 2934 668 2968 1444
rect 3392 668 3426 1444
rect 3522 668 3556 1444
rect 3980 668 4014 1444
rect 4110 668 4144 1444
rect 4568 668 4602 1444
rect 4698 668 4732 1444
rect 5156 668 5190 1444
rect 5286 668 5320 1444
rect 5744 668 5778 1444
rect 5874 668 5908 1444
rect 6332 668 6366 1444
rect 6462 668 6496 1444
rect 6920 668 6954 1444
rect 7050 668 7084 1444
rect 7508 668 7542 1444
rect 7638 668 7672 1444
rect 8096 668 8130 1444
rect 8226 668 8260 1444
rect 8684 668 8718 1444
rect 8814 668 8848 1444
rect 9272 668 9306 1444
rect 9402 668 9436 1444
rect 9860 668 9894 1444
rect 9990 668 10024 1444
rect 10448 668 10482 1444
rect 10578 668 10612 1444
rect 11036 668 11070 1444
rect 11166 668 11200 1444
rect 11624 668 11658 1444
rect 11754 668 11788 1444
rect 12212 668 12246 1444
rect 12342 668 12376 1444
rect 12800 668 12834 1444
rect 12930 668 12964 1444
rect 13388 668 13422 1444
rect 13518 668 13552 1444
rect 13976 668 14010 1444
rect 14106 668 14140 1444
rect 14564 668 14598 1444
rect 14694 668 14728 1444
rect 15152 668 15186 1444
rect 15282 668 15316 1444
rect 15740 668 15774 1444
rect 15870 668 15904 1444
rect 16328 668 16362 1444
rect 16458 668 16492 1444
rect 16916 668 16950 1444
rect 17046 668 17080 1444
rect 17504 668 17538 1444
rect 17634 668 17668 1444
rect 18092 668 18126 1444
rect 18222 668 18256 1444
rect 18680 668 18714 1444
rect 18810 668 18844 1444
rect 19268 668 19302 1444
rect 19398 668 19432 1444
rect 19856 668 19890 1444
rect 19986 668 20020 1444
rect 20444 668 20478 1444
rect 20574 668 20608 1444
rect 21032 668 21066 1444
rect 21162 668 21196 1444
rect 21620 668 21654 1444
rect -6412 575 -6044 609
rect -5824 575 -5456 609
rect -5236 575 -4868 609
rect -4648 575 -4280 609
rect -4060 575 -3692 609
rect -3472 575 -3104 609
rect -2884 575 -2516 609
rect -2296 575 -1928 609
rect -1708 575 -1340 609
rect -1120 575 -752 609
rect -532 575 -164 609
rect 56 575 424 609
rect 644 575 1012 609
rect 1232 575 1600 609
rect 1820 575 2188 609
rect 2408 575 2776 609
rect 2996 575 3364 609
rect 3584 575 3952 609
rect 4172 575 4540 609
rect 4760 575 5128 609
rect 5348 575 5716 609
rect 5936 575 6304 609
rect 6524 575 6892 609
rect 7112 575 7480 609
rect 7700 575 8068 609
rect 8288 575 8656 609
rect 8876 575 9244 609
rect 9464 575 9832 609
rect 10052 575 10420 609
rect 10640 575 11008 609
rect 11228 575 11596 609
rect 11816 575 12184 609
rect 12404 575 12772 609
rect 12992 575 13360 609
rect 13580 575 13948 609
rect 14168 575 14536 609
rect 14756 575 15124 609
rect 15344 575 15712 609
rect 15932 575 16300 609
rect 16520 575 16888 609
rect 17108 575 17476 609
rect 17696 575 18064 609
rect 18284 575 18652 609
rect 18872 575 19240 609
rect 19460 575 19828 609
rect 20048 575 20416 609
rect 20636 575 21004 609
rect 21224 575 21592 609
rect -6412 503 -6044 537
rect -5824 503 -5456 537
rect -5236 503 -4868 537
rect -4648 503 -4280 537
rect -4060 503 -3692 537
rect -3472 503 -3104 537
rect -2884 503 -2516 537
rect -2296 503 -1928 537
rect -1708 503 -1340 537
rect -1120 503 -752 537
rect -532 503 -164 537
rect 56 503 424 537
rect 644 503 1012 537
rect 1232 503 1600 537
rect 1820 503 2188 537
rect 2408 503 2776 537
rect 2996 503 3364 537
rect 3584 503 3952 537
rect 4172 503 4540 537
rect 4760 503 5128 537
rect 5348 503 5716 537
rect 5936 503 6304 537
rect 6524 503 6892 537
rect 7112 503 7480 537
rect 7700 503 8068 537
rect 8288 503 8656 537
rect 8876 503 9244 537
rect 9464 503 9832 537
rect 10052 503 10420 537
rect 10640 503 11008 537
rect 11228 503 11596 537
rect 11816 503 12184 537
rect 12404 503 12772 537
rect 12992 503 13360 537
rect 13580 503 13948 537
rect 14168 503 14536 537
rect 14756 503 15124 537
rect 15344 503 15712 537
rect 15932 503 16300 537
rect 16520 503 16888 537
rect 17108 503 17476 537
rect 17696 503 18064 537
rect 18284 503 18652 537
rect 18872 503 19240 537
rect 19460 503 19828 537
rect 20048 503 20416 537
rect 20636 503 21004 537
rect 21224 503 21592 537
rect -6474 -332 -6440 444
rect -6016 -332 -5982 444
rect -5886 -332 -5852 444
rect -5428 -332 -5394 444
rect -5298 -332 -5264 444
rect -4840 -332 -4806 444
rect -4710 -332 -4676 444
rect -4252 -332 -4218 444
rect -4122 -332 -4088 444
rect -3664 -332 -3630 444
rect -3534 -332 -3500 444
rect -3076 -332 -3042 444
rect -2946 -332 -2912 444
rect -2488 -332 -2454 444
rect -2358 -332 -2324 444
rect -1900 -332 -1866 444
rect -1770 -332 -1736 444
rect -1312 -332 -1278 444
rect -1182 -332 -1148 444
rect -724 -332 -690 444
rect -594 -332 -560 444
rect -136 -332 -102 444
rect -6 -332 28 444
rect 452 -332 486 444
rect 582 -332 616 444
rect 1040 -332 1074 444
rect 1170 -332 1204 444
rect 1628 -332 1662 444
rect 1758 -332 1792 444
rect 2216 -332 2250 444
rect 2346 -332 2380 444
rect 2804 -332 2838 444
rect 2934 -332 2968 444
rect 3392 -332 3426 444
rect 3522 -332 3556 444
rect 3980 -332 4014 444
rect 4110 -332 4144 444
rect 4568 -332 4602 444
rect 4698 -332 4732 444
rect 5156 -332 5190 444
rect 5286 -332 5320 444
rect 5744 -332 5778 444
rect 5874 -332 5908 444
rect 6332 -332 6366 444
rect 6462 -332 6496 444
rect 6920 -332 6954 444
rect 7050 -332 7084 444
rect 7508 -332 7542 444
rect 7638 -332 7672 444
rect 8096 -332 8130 444
rect 8226 -332 8260 444
rect 8684 -332 8718 444
rect 8814 -332 8848 444
rect 9272 -332 9306 444
rect 9402 -332 9436 444
rect 9860 -332 9894 444
rect 9990 -332 10024 444
rect 10448 -332 10482 444
rect 10578 -332 10612 444
rect 11036 -332 11070 444
rect 11166 -332 11200 444
rect 11624 -332 11658 444
rect 11754 -332 11788 444
rect 12212 -332 12246 444
rect 12342 -332 12376 444
rect 12800 -332 12834 444
rect 12930 -332 12964 444
rect 13388 -332 13422 444
rect 13518 -332 13552 444
rect 13976 -332 14010 444
rect 14106 -332 14140 444
rect 14564 -332 14598 444
rect 14694 -332 14728 444
rect 15152 -332 15186 444
rect 15282 -332 15316 444
rect 15740 -332 15774 444
rect 15870 -332 15904 444
rect 16328 -332 16362 444
rect 16458 -332 16492 444
rect 16916 -332 16950 444
rect 17046 -332 17080 444
rect 17504 -332 17538 444
rect 17634 -332 17668 444
rect 18092 -332 18126 444
rect 18222 -332 18256 444
rect 18680 -332 18714 444
rect 18810 -332 18844 444
rect 19268 -332 19302 444
rect 19398 -332 19432 444
rect 19856 -332 19890 444
rect 19986 -332 20020 444
rect 20444 -332 20478 444
rect 20574 -332 20608 444
rect 21032 -332 21066 444
rect 21162 -332 21196 444
rect 21620 -332 21654 444
rect -6412 -425 -6044 -391
rect -5824 -425 -5456 -391
rect -5236 -425 -4868 -391
rect -4648 -425 -4280 -391
rect -4060 -425 -3692 -391
rect -3472 -425 -3104 -391
rect -2884 -425 -2516 -391
rect -2296 -425 -1928 -391
rect -1708 -425 -1340 -391
rect -1120 -425 -752 -391
rect -532 -425 -164 -391
rect 56 -425 424 -391
rect 644 -425 1012 -391
rect 1232 -425 1600 -391
rect 1820 -425 2188 -391
rect 2408 -425 2776 -391
rect 2996 -425 3364 -391
rect 3584 -425 3952 -391
rect 4172 -425 4540 -391
rect 4760 -425 5128 -391
rect 5348 -425 5716 -391
rect 5936 -425 6304 -391
rect 6524 -425 6892 -391
rect 7112 -425 7480 -391
rect 7700 -425 8068 -391
rect 8288 -425 8656 -391
rect 8876 -425 9244 -391
rect 9464 -425 9832 -391
rect 10052 -425 10420 -391
rect 10640 -425 11008 -391
rect 11228 -425 11596 -391
rect 11816 -425 12184 -391
rect 12404 -425 12772 -391
rect 12992 -425 13360 -391
rect 13580 -425 13948 -391
rect 14168 -425 14536 -391
rect 14756 -425 15124 -391
rect 15344 -425 15712 -391
rect 15932 -425 16300 -391
rect 16520 -425 16888 -391
rect 17108 -425 17476 -391
rect 17696 -425 18064 -391
rect 18284 -425 18652 -391
rect 18872 -425 19240 -391
rect 19460 -425 19828 -391
rect 20048 -425 20416 -391
rect 20636 -425 21004 -391
rect 21224 -425 21592 -391
rect -6028 -742 -5840 -694
rect -4852 -742 -4664 -694
rect -3676 -742 -3488 -694
rect -2500 -742 -2312 -694
rect -1324 -742 -1136 -694
rect -148 -742 40 -694
rect 1028 -742 1216 -694
rect 2204 -742 2392 -694
rect 3380 -742 3568 -694
rect 4556 -742 4744 -694
rect 5732 -742 5920 -694
rect 6908 -742 7096 -694
rect 8084 -742 8272 -694
rect 9260 -742 9448 -694
rect 10436 -742 10624 -694
rect 11612 -742 11800 -694
rect 12788 -742 12976 -684
rect 13964 -742 14152 -694
rect 15140 -742 15328 -694
rect 16316 -742 16504 -694
rect 17478 -742 17690 -684
rect 18668 -742 18856 -694
rect 19844 -742 20032 -694
rect 21020 -742 21208 -694
rect -6028 -776 -5840 -742
rect -4852 -776 -4664 -742
rect -3676 -776 -3488 -742
rect -2500 -776 -2312 -742
rect -1324 -776 -1136 -742
rect -148 -776 40 -742
rect 1028 -776 1216 -742
rect 2204 -776 2392 -742
rect 3380 -776 3568 -742
rect 4556 -776 4744 -742
rect 5732 -776 5920 -742
rect 6908 -776 7096 -742
rect 8084 -776 8272 -742
rect 9260 -776 9448 -742
rect 10436 -776 10624 -742
rect 11612 -776 11800 -742
rect 12788 -776 12976 -742
rect 13964 -776 14152 -742
rect 15140 -776 15328 -742
rect 16316 -776 16504 -742
rect 17478 -776 17690 -742
rect 18668 -776 18856 -742
rect 19844 -776 20032 -742
rect 21020 -776 21208 -742
rect -6028 -804 -5840 -776
rect -4852 -804 -4664 -776
rect -3676 -804 -3488 -776
rect -2500 -804 -2312 -776
rect -1324 -804 -1136 -776
rect -148 -804 40 -776
rect 1028 -804 1216 -776
rect 2204 -804 2392 -776
rect 3380 -804 3568 -776
rect 4556 -804 4744 -776
rect 5732 -804 5920 -776
rect 6908 -804 7096 -776
rect 8084 -804 8272 -776
rect 9260 -804 9448 -776
rect 10436 -804 10624 -776
rect 11612 -804 11800 -776
rect 12788 -794 12976 -776
rect 13964 -804 14152 -776
rect 15140 -804 15328 -776
rect 16316 -804 16504 -776
rect 17478 -806 17690 -776
rect 18668 -804 18856 -776
rect 19844 -804 20032 -776
rect 21020 -804 21208 -776
rect 6640 -1952 6678 -1820
rect 6906 -1952 6944 -1820
rect 7172 -1952 7210 -1820
rect 7438 -1952 7476 -1820
rect 7704 -1952 7742 -1820
rect 7970 -1952 8008 -1820
rect 8236 -1952 8274 -1820
rect 8502 -1952 8540 -1820
rect 6578 -2778 6612 -2002
rect 6706 -2778 6740 -2002
rect 6844 -2778 6878 -2002
rect 6972 -2778 7006 -2002
rect 7110 -2778 7144 -2002
rect 7238 -2778 7272 -2002
rect 7376 -2778 7410 -2002
rect 7504 -2778 7538 -2002
rect 7642 -2778 7676 -2002
rect 7770 -2778 7804 -2002
rect 7908 -2778 7942 -2002
rect 8036 -2778 8070 -2002
rect 8174 -2778 8208 -2002
rect 8302 -2778 8336 -2002
rect 8440 -2778 8474 -2002
rect 8568 -2778 8602 -2002
rect 6640 -2962 6678 -2830
rect 6906 -2962 6944 -2830
rect 7172 -2962 7210 -2830
rect 7438 -2962 7476 -2830
rect 7704 -2962 7742 -2830
rect 7970 -2962 8008 -2830
rect 8236 -2962 8274 -2830
rect 8502 -2962 8540 -2830
rect 6578 -3788 6612 -3012
rect 6706 -3788 6740 -3012
rect 6844 -3788 6878 -3012
rect 6972 -3788 7006 -3012
rect 7110 -3788 7144 -3012
rect 7238 -3788 7272 -3012
rect 7376 -3788 7410 -3012
rect 7504 -3788 7538 -3012
rect 7642 -3788 7676 -3012
rect 7770 -3788 7804 -3012
rect 7908 -3788 7942 -3012
rect 8036 -3788 8070 -3012
rect 8174 -3788 8208 -3012
rect 8302 -3788 8336 -3012
rect 8440 -3788 8474 -3012
rect 8568 -3788 8602 -3012
rect 6640 -3972 6678 -3840
rect 6906 -3972 6944 -3840
rect 7172 -3972 7210 -3840
rect 7438 -3972 7476 -3840
rect 7704 -3972 7742 -3840
rect 7970 -3972 8008 -3840
rect 8236 -3972 8274 -3840
rect 8502 -3972 8540 -3840
rect 6578 -4798 6612 -4022
rect 6706 -4798 6740 -4022
rect 6844 -4798 6878 -4022
rect 6972 -4798 7006 -4022
rect 7110 -4798 7144 -4022
rect 7238 -4798 7272 -4022
rect 7376 -4798 7410 -4022
rect 7504 -4798 7538 -4022
rect 7642 -4798 7676 -4022
rect 7770 -4798 7804 -4022
rect 7908 -4798 7942 -4022
rect 8036 -4798 8070 -4022
rect 8174 -4798 8208 -4022
rect 8302 -4798 8336 -4022
rect 8440 -4798 8474 -4022
rect 8568 -4798 8602 -4022
rect 6640 -4982 6678 -4850
rect 6906 -4982 6944 -4850
rect 7172 -4982 7210 -4850
rect 7438 -4982 7476 -4850
rect 7704 -4982 7742 -4850
rect 7970 -4982 8008 -4850
rect 8236 -4982 8274 -4850
rect 8502 -4982 8540 -4850
rect 13759 -3912 13797 -3515
rect 13759 -4903 13797 -4506
rect 14048 -4582 14188 -4122
rect 7212 -6144 7250 -6018
rect 7452 -6144 7490 -6018
rect 7692 -6144 7730 -6018
rect 7932 -6144 7970 -6018
rect 7150 -6770 7184 -6194
rect 7278 -6770 7312 -6194
rect 7390 -6770 7424 -6194
rect 7518 -6770 7552 -6194
rect 7630 -6770 7664 -6194
rect 7758 -6770 7792 -6194
rect 7870 -6770 7904 -6194
rect 7998 -6770 8032 -6194
rect 7212 -6952 7250 -6820
rect 7452 -6952 7490 -6820
rect 7692 -6952 7730 -6820
rect 7932 -6952 7970 -6820
rect 7150 -7578 7184 -7002
rect 7278 -7578 7312 -7002
rect 7390 -7578 7424 -7002
rect 7518 -7578 7552 -7002
rect 7630 -7578 7664 -7002
rect 7758 -7578 7792 -7002
rect 7870 -7578 7904 -7002
rect 7998 -7578 8032 -7002
rect 7212 -7760 7250 -7628
rect 7452 -7760 7490 -7628
rect 7692 -7760 7730 -7628
rect 7932 -7760 7970 -7628
rect 6902 -8060 8254 -8012
rect 6902 -8094 6962 -8060
rect 6962 -8094 8172 -8060
rect 8172 -8094 8254 -8060
rect 6902 -8124 8254 -8094
<< metal1 >>
rect 2964 7090 3098 7096
rect 2964 7018 2976 7090
rect 3086 7018 3098 7090
rect 2964 7012 3098 7018
rect 3444 7090 3578 7096
rect 3444 7018 3456 7090
rect 3566 7018 3578 7090
rect 3444 7012 3578 7018
rect 3924 7090 4058 7096
rect 3924 7018 3936 7090
rect 4046 7018 4058 7090
rect 3924 7012 4058 7018
rect 4404 7090 4538 7096
rect 4404 7018 4416 7090
rect 4526 7018 4538 7090
rect 4404 7012 4538 7018
rect 4884 7090 5018 7096
rect 4884 7018 4896 7090
rect 5006 7018 5018 7090
rect 4884 7012 5018 7018
rect 5364 7090 5498 7096
rect 5364 7018 5376 7090
rect 5486 7018 5498 7090
rect 5364 7012 5498 7018
rect 5844 7090 5978 7096
rect 5844 7018 5856 7090
rect 5966 7018 5978 7090
rect 5844 7012 5978 7018
rect 6324 7090 6458 7096
rect 6324 7018 6336 7090
rect 6446 7018 6458 7090
rect 6324 7012 6458 7018
rect 6804 7090 6938 7096
rect 6804 7018 6816 7090
rect 6926 7018 6938 7090
rect 6804 7012 6938 7018
rect 7284 7090 7418 7096
rect 7284 7018 7296 7090
rect 7406 7018 7418 7090
rect 7284 7012 7418 7018
rect 7764 7090 7898 7096
rect 7764 7018 7776 7090
rect 7886 7018 7898 7090
rect 7764 7012 7898 7018
rect 8244 7090 8378 7096
rect 8244 7018 8256 7090
rect 8366 7018 8378 7090
rect 8244 7012 8378 7018
rect 8724 7090 8858 7096
rect 8724 7018 8736 7090
rect 8846 7018 8858 7090
rect 8724 7012 8858 7018
rect 9204 7090 9338 7096
rect 9204 7018 9216 7090
rect 9326 7018 9338 7090
rect 9204 7012 9338 7018
rect 9684 7090 9818 7096
rect 9684 7018 9696 7090
rect 9806 7018 9818 7090
rect 9684 7012 9818 7018
rect 10164 7090 10298 7096
rect 10164 7018 10176 7090
rect 10286 7018 10298 7090
rect 10164 7012 10298 7018
rect 10644 7090 10778 7096
rect 10644 7018 10656 7090
rect 10766 7018 10778 7090
rect 10644 7012 10778 7018
rect 11124 7090 11258 7096
rect 11124 7018 11136 7090
rect 11246 7018 11258 7090
rect 11124 7012 11258 7018
rect 11604 7090 11738 7096
rect 11604 7018 11616 7090
rect 11726 7018 11738 7090
rect 11604 7012 11738 7018
rect 12084 7090 12218 7096
rect 12084 7018 12096 7090
rect 12206 7018 12218 7090
rect 12084 7012 12218 7018
rect 2876 6746 2946 6752
rect 2866 6614 2876 6746
rect 2946 6614 2956 6746
rect 2876 6608 2946 6614
rect 3004 6576 3058 7012
rect 3116 6746 3186 6752
rect 3106 6614 3116 6746
rect 3186 6614 3196 6746
rect 3116 6608 3186 6614
rect 3244 6604 3298 6756
rect 3356 6746 3426 6752
rect 3346 6614 3356 6746
rect 3426 6614 3436 6746
rect 3356 6608 3426 6614
rect 3484 6576 3538 7012
rect 3596 6746 3666 6752
rect 3586 6614 3596 6746
rect 3666 6614 3676 6746
rect 3596 6608 3666 6614
rect 3724 6604 3778 6756
rect 3836 6746 3906 6752
rect 3826 6614 3836 6746
rect 3906 6614 3916 6746
rect 3836 6608 3906 6614
rect 3964 6576 4018 7012
rect 4076 6746 4146 6752
rect 4066 6614 4076 6746
rect 4146 6614 4156 6746
rect 4076 6608 4146 6614
rect 4204 6604 4258 6756
rect 4316 6746 4386 6752
rect 4306 6614 4316 6746
rect 4386 6614 4396 6746
rect 4316 6608 4386 6614
rect 4444 6576 4498 7012
rect 4556 6746 4626 6752
rect 4546 6614 4556 6746
rect 4626 6614 4636 6746
rect 4556 6608 4626 6614
rect 4684 6604 4738 6756
rect 4796 6746 4866 6752
rect 4786 6614 4796 6746
rect 4866 6614 4876 6746
rect 4796 6608 4866 6614
rect 4924 6576 4978 7012
rect 5036 6746 5106 6752
rect 5026 6614 5036 6746
rect 5106 6614 5116 6746
rect 5036 6608 5106 6614
rect 5164 6604 5218 6756
rect 5276 6746 5346 6752
rect 5266 6614 5276 6746
rect 5346 6614 5356 6746
rect 5276 6608 5346 6614
rect 5404 6576 5458 7012
rect 5516 6746 5586 6752
rect 5506 6614 5516 6746
rect 5586 6614 5596 6746
rect 5516 6608 5586 6614
rect 5644 6604 5698 6756
rect 5756 6746 5826 6752
rect 5746 6614 5756 6746
rect 5826 6614 5836 6746
rect 5756 6608 5826 6614
rect 5884 6576 5938 7012
rect 5996 6746 6066 6752
rect 5986 6614 5996 6746
rect 6066 6614 6076 6746
rect 5996 6608 6066 6614
rect 6124 6604 6178 6756
rect 6236 6746 6306 6752
rect 6226 6614 6236 6746
rect 6306 6614 6316 6746
rect 6236 6608 6306 6614
rect 6364 6576 6418 7012
rect 6476 6746 6546 6752
rect 6466 6614 6476 6746
rect 6546 6614 6556 6746
rect 6476 6608 6546 6614
rect 6604 6604 6658 6756
rect 6716 6746 6786 6752
rect 6706 6614 6716 6746
rect 6786 6614 6796 6746
rect 6716 6608 6786 6614
rect 6844 6576 6898 7012
rect 6956 6746 7026 6752
rect 6946 6614 6956 6746
rect 7026 6614 7036 6746
rect 6956 6608 7026 6614
rect 7084 6604 7138 6756
rect 7196 6746 7266 6752
rect 7186 6614 7196 6746
rect 7266 6614 7276 6746
rect 7196 6608 7266 6614
rect 7324 6576 7378 7012
rect 7436 6746 7506 6752
rect 7426 6614 7436 6746
rect 7506 6614 7516 6746
rect 7436 6608 7506 6614
rect 7564 6604 7618 6756
rect 7676 6746 7746 6752
rect 7666 6614 7676 6746
rect 7746 6614 7756 6746
rect 7676 6608 7746 6614
rect 7804 6576 7858 7012
rect 7916 6746 7986 6752
rect 7906 6614 7916 6746
rect 7986 6614 7996 6746
rect 7916 6608 7986 6614
rect 8044 6604 8098 6756
rect 8156 6746 8226 6752
rect 8146 6614 8156 6746
rect 8226 6614 8236 6746
rect 8156 6608 8226 6614
rect 8284 6576 8338 7012
rect 8396 6746 8466 6752
rect 8386 6614 8396 6746
rect 8466 6614 8476 6746
rect 8396 6608 8466 6614
rect 8524 6604 8578 6756
rect 8636 6746 8706 6752
rect 8626 6614 8636 6746
rect 8706 6614 8716 6746
rect 8636 6608 8706 6614
rect 8764 6576 8818 7012
rect 8876 6746 8946 6752
rect 8866 6614 8876 6746
rect 8946 6614 8956 6746
rect 8876 6608 8946 6614
rect 9004 6604 9058 6756
rect 9116 6746 9186 6752
rect 9106 6614 9116 6746
rect 9186 6614 9196 6746
rect 9116 6608 9186 6614
rect 9244 6576 9298 7012
rect 9356 6746 9426 6752
rect 9346 6614 9356 6746
rect 9426 6614 9436 6746
rect 9356 6608 9426 6614
rect 9484 6604 9538 6756
rect 9596 6746 9666 6752
rect 9586 6614 9596 6746
rect 9666 6614 9676 6746
rect 9596 6608 9666 6614
rect 9724 6576 9778 7012
rect 9836 6746 9906 6752
rect 9826 6614 9836 6746
rect 9906 6614 9916 6746
rect 9836 6608 9906 6614
rect 9964 6604 10018 6756
rect 10076 6746 10146 6752
rect 10066 6614 10076 6746
rect 10146 6614 10156 6746
rect 10076 6608 10146 6614
rect 10204 6576 10258 7012
rect 10316 6746 10386 6752
rect 10306 6614 10316 6746
rect 10386 6614 10396 6746
rect 10316 6608 10386 6614
rect 10444 6604 10498 6756
rect 10556 6746 10626 6752
rect 10546 6614 10556 6746
rect 10626 6614 10636 6746
rect 10556 6608 10626 6614
rect 10684 6576 10738 7012
rect 10796 6746 10866 6752
rect 10786 6614 10796 6746
rect 10866 6614 10876 6746
rect 10796 6608 10866 6614
rect 10924 6604 10978 6756
rect 11036 6746 11106 6752
rect 11026 6614 11036 6746
rect 11106 6614 11116 6746
rect 11036 6608 11106 6614
rect 11164 6576 11218 7012
rect 11276 6746 11346 6752
rect 11266 6614 11276 6746
rect 11346 6614 11356 6746
rect 11276 6608 11346 6614
rect 11404 6604 11458 6756
rect 11516 6746 11586 6752
rect 11506 6614 11516 6746
rect 11586 6614 11596 6746
rect 11516 6608 11586 6614
rect 11644 6576 11698 7012
rect 11756 6746 11826 6752
rect 11746 6614 11756 6746
rect 11826 6614 11836 6746
rect 11756 6608 11826 6614
rect 11884 6604 11938 6756
rect 11996 6746 12066 6752
rect 11986 6614 11996 6746
rect 12066 6614 12076 6746
rect 11996 6608 12066 6614
rect 12124 6576 12178 7012
rect 12236 6746 12306 6752
rect 12226 6614 12236 6746
rect 12306 6614 12316 6746
rect 12236 6608 12306 6614
rect 2752 6564 2870 6576
rect 2752 5988 2830 6564
rect 2864 5988 2870 6564
rect 2752 5976 2870 5988
rect 2952 6564 3110 6576
rect 2952 5988 2958 6564
rect 2992 5988 3070 6564
rect 3104 5988 3110 6564
rect 2952 5976 3110 5988
rect 3192 6564 3350 6576
rect 3192 5988 3198 6564
rect 3232 5988 3310 6564
rect 3344 5988 3350 6564
rect 3192 5976 3350 5988
rect 3432 6564 3590 6576
rect 3432 5988 3438 6564
rect 3472 5988 3550 6564
rect 3584 5988 3590 6564
rect 3432 5976 3590 5988
rect 3672 6564 3830 6576
rect 3672 5988 3678 6564
rect 3712 5988 3790 6564
rect 3824 5988 3830 6564
rect 3672 5976 3830 5988
rect 3912 6564 4070 6576
rect 3912 5988 3918 6564
rect 3952 5988 4030 6564
rect 4064 5988 4070 6564
rect 3912 5976 4070 5988
rect 4152 6564 4310 6576
rect 4152 5988 4158 6564
rect 4192 5988 4270 6564
rect 4304 5988 4310 6564
rect 4152 5976 4310 5988
rect 4392 6564 4550 6576
rect 4392 5988 4398 6564
rect 4432 5988 4510 6564
rect 4544 5988 4550 6564
rect 4392 5976 4550 5988
rect 4632 6564 4790 6576
rect 4632 5988 4638 6564
rect 4672 5988 4750 6564
rect 4784 5988 4790 6564
rect 4632 5976 4790 5988
rect 4872 6564 5030 6576
rect 4872 5988 4878 6564
rect 4912 5988 4990 6564
rect 5024 5988 5030 6564
rect 4872 5976 5030 5988
rect 5112 6564 5270 6576
rect 5112 5988 5118 6564
rect 5152 5988 5230 6564
rect 5264 5988 5270 6564
rect 5112 5976 5270 5988
rect 5352 6564 5510 6576
rect 5352 5988 5358 6564
rect 5392 5988 5470 6564
rect 5504 5988 5510 6564
rect 5352 5976 5510 5988
rect 5592 6564 5750 6576
rect 5592 5988 5598 6564
rect 5632 5988 5710 6564
rect 5744 5988 5750 6564
rect 5592 5976 5750 5988
rect 5832 6564 5990 6576
rect 5832 5988 5838 6564
rect 5872 5988 5950 6564
rect 5984 5988 5990 6564
rect 5832 5976 5990 5988
rect 6072 6564 6230 6576
rect 6072 5988 6078 6564
rect 6112 5988 6190 6564
rect 6224 5988 6230 6564
rect 6072 5976 6230 5988
rect 6312 6564 6470 6576
rect 6312 5988 6318 6564
rect 6352 5988 6430 6564
rect 6464 5988 6470 6564
rect 6312 5976 6470 5988
rect 6552 6564 6710 6576
rect 6552 5988 6558 6564
rect 6592 5988 6670 6564
rect 6704 5988 6710 6564
rect 6552 5976 6710 5988
rect 6792 6564 6950 6576
rect 6792 5988 6798 6564
rect 6832 5988 6910 6564
rect 6944 5988 6950 6564
rect 6792 5976 6950 5988
rect 7032 6564 7190 6576
rect 7032 5988 7038 6564
rect 7072 5988 7150 6564
rect 7184 5988 7190 6564
rect 7032 5976 7190 5988
rect 7272 6564 7430 6576
rect 7272 5988 7278 6564
rect 7312 5988 7390 6564
rect 7424 5988 7430 6564
rect 7272 5976 7430 5988
rect 7512 6564 7670 6576
rect 7512 5988 7518 6564
rect 7552 5988 7630 6564
rect 7664 5988 7670 6564
rect 7512 5976 7670 5988
rect 7752 6564 7910 6576
rect 7752 5988 7758 6564
rect 7792 5988 7870 6564
rect 7904 5988 7910 6564
rect 7752 5976 7910 5988
rect 7992 6564 8150 6576
rect 7992 5988 7998 6564
rect 8032 5988 8110 6564
rect 8144 5988 8150 6564
rect 7992 5976 8150 5988
rect 8232 6564 8390 6576
rect 8232 5988 8238 6564
rect 8272 5988 8350 6564
rect 8384 5988 8390 6564
rect 8232 5976 8390 5988
rect 8472 6564 8630 6576
rect 8472 5988 8478 6564
rect 8512 5988 8590 6564
rect 8624 5988 8630 6564
rect 8472 5976 8630 5988
rect 8712 6564 8870 6576
rect 8712 5988 8718 6564
rect 8752 5988 8830 6564
rect 8864 5988 8870 6564
rect 8712 5976 8870 5988
rect 8952 6564 9110 6576
rect 8952 5988 8958 6564
rect 8992 5988 9070 6564
rect 9104 5988 9110 6564
rect 8952 5976 9110 5988
rect 9192 6564 9350 6576
rect 9192 5988 9198 6564
rect 9232 5988 9310 6564
rect 9344 5988 9350 6564
rect 9192 5976 9350 5988
rect 9432 6564 9590 6576
rect 9432 5988 9438 6564
rect 9472 5988 9550 6564
rect 9584 5988 9590 6564
rect 9432 5976 9590 5988
rect 9672 6564 9830 6576
rect 9672 5988 9678 6564
rect 9712 5988 9790 6564
rect 9824 5988 9830 6564
rect 9672 5976 9830 5988
rect 9912 6564 10070 6576
rect 9912 5988 9918 6564
rect 9952 5988 10030 6564
rect 10064 5988 10070 6564
rect 9912 5976 10070 5988
rect 10152 6564 10310 6576
rect 10152 5988 10158 6564
rect 10192 5988 10270 6564
rect 10304 5988 10310 6564
rect 10152 5976 10310 5988
rect 10392 6564 10550 6576
rect 10392 5988 10398 6564
rect 10432 5988 10510 6564
rect 10544 5988 10550 6564
rect 10392 5976 10550 5988
rect 10632 6564 10790 6576
rect 10632 5988 10638 6564
rect 10672 5988 10750 6564
rect 10784 5988 10790 6564
rect 10632 5976 10790 5988
rect 10872 6564 11030 6576
rect 10872 5988 10878 6564
rect 10912 5988 10990 6564
rect 11024 5988 11030 6564
rect 10872 5976 11030 5988
rect 11112 6564 11270 6576
rect 11112 5988 11118 6564
rect 11152 5988 11230 6564
rect 11264 5988 11270 6564
rect 11112 5976 11270 5988
rect 11352 6564 11510 6576
rect 11352 5988 11358 6564
rect 11392 5988 11470 6564
rect 11504 5988 11510 6564
rect 11352 5976 11510 5988
rect 11592 6564 11750 6576
rect 11592 5988 11598 6564
rect 11632 5988 11710 6564
rect 11744 5988 11750 6564
rect 11592 5976 11750 5988
rect 11832 6564 11990 6576
rect 11832 5988 11838 6564
rect 11872 5988 11950 6564
rect 11984 5988 11990 6564
rect 11832 5976 11990 5988
rect 12072 6564 12230 6576
rect 12072 5988 12078 6564
rect 12112 5988 12190 6564
rect 12224 5988 12230 6564
rect 12072 5976 12230 5988
rect 12312 6564 12430 6576
rect 12312 5988 12318 6564
rect 12352 5988 12430 6564
rect 12312 5976 12430 5988
rect 2752 5768 2830 5976
rect 2876 5938 2946 5944
rect 2866 5806 2876 5938
rect 2946 5806 2956 5938
rect 2876 5800 2946 5806
rect 2998 5768 3064 5976
rect 3116 5938 3186 5944
rect 3106 5806 3116 5938
rect 3186 5806 3196 5938
rect 3116 5800 3186 5806
rect 3238 5768 3304 5976
rect 3356 5938 3426 5944
rect 3346 5806 3356 5938
rect 3426 5806 3436 5938
rect 3356 5800 3426 5806
rect 3478 5768 3544 5976
rect 3596 5938 3666 5944
rect 3586 5806 3596 5938
rect 3666 5806 3676 5938
rect 3596 5800 3666 5806
rect 3712 5768 3790 5976
rect 3836 5938 3906 5944
rect 3826 5806 3836 5938
rect 3906 5806 3916 5938
rect 3836 5800 3906 5806
rect 3958 5768 4024 5976
rect 4076 5938 4146 5944
rect 4066 5806 4076 5938
rect 4146 5806 4156 5938
rect 4076 5800 4146 5806
rect 4198 5768 4264 5976
rect 4316 5938 4386 5944
rect 4306 5806 4316 5938
rect 4386 5806 4396 5938
rect 4316 5800 4386 5806
rect 4438 5768 4504 5976
rect 4556 5938 4626 5944
rect 4546 5806 4556 5938
rect 4626 5806 4636 5938
rect 4556 5800 4626 5806
rect 4672 5768 4750 5976
rect 4796 5938 4866 5944
rect 4786 5806 4796 5938
rect 4866 5806 4876 5938
rect 4796 5800 4866 5806
rect 4918 5768 4984 5976
rect 5036 5938 5106 5944
rect 5026 5806 5036 5938
rect 5106 5806 5116 5938
rect 5036 5800 5106 5806
rect 5158 5768 5224 5976
rect 5276 5938 5346 5944
rect 5266 5806 5276 5938
rect 5346 5806 5356 5938
rect 5276 5800 5346 5806
rect 5398 5768 5464 5976
rect 5516 5938 5586 5944
rect 5506 5806 5516 5938
rect 5586 5806 5596 5938
rect 5516 5800 5586 5806
rect 5632 5768 5710 5976
rect 5756 5938 5826 5944
rect 5746 5806 5756 5938
rect 5826 5806 5836 5938
rect 5756 5800 5826 5806
rect 5878 5768 5944 5976
rect 5996 5938 6066 5944
rect 5986 5806 5996 5938
rect 6066 5806 6076 5938
rect 5996 5800 6066 5806
rect 6118 5768 6184 5976
rect 6236 5938 6306 5944
rect 6226 5806 6236 5938
rect 6306 5806 6316 5938
rect 6236 5800 6306 5806
rect 6358 5768 6424 5976
rect 6476 5938 6546 5944
rect 6466 5806 6476 5938
rect 6546 5806 6556 5938
rect 6476 5800 6546 5806
rect 6592 5768 6670 5976
rect 6716 5938 6786 5944
rect 6706 5806 6716 5938
rect 6786 5806 6796 5938
rect 6716 5800 6786 5806
rect 6838 5768 6904 5976
rect 6956 5938 7026 5944
rect 6946 5806 6956 5938
rect 7026 5806 7036 5938
rect 6956 5800 7026 5806
rect 7078 5768 7144 5976
rect 7196 5938 7266 5944
rect 7186 5806 7196 5938
rect 7266 5806 7276 5938
rect 7196 5800 7266 5806
rect 7318 5768 7384 5976
rect 7436 5938 7506 5944
rect 7426 5806 7436 5938
rect 7506 5806 7516 5938
rect 7436 5800 7506 5806
rect 7552 5768 7630 5976
rect 7676 5938 7746 5944
rect 7666 5806 7676 5938
rect 7746 5806 7756 5938
rect 7676 5800 7746 5806
rect 7798 5768 7864 5976
rect 7916 5938 7986 5944
rect 7906 5806 7916 5938
rect 7986 5806 7996 5938
rect 7916 5800 7986 5806
rect 8038 5768 8104 5976
rect 8156 5938 8226 5944
rect 8146 5806 8156 5938
rect 8226 5806 8236 5938
rect 8156 5800 8226 5806
rect 8278 5768 8344 5976
rect 8396 5938 8466 5944
rect 8386 5806 8396 5938
rect 8466 5806 8476 5938
rect 8396 5800 8466 5806
rect 8512 5768 8590 5976
rect 8636 5938 8706 5944
rect 8626 5806 8636 5938
rect 8706 5806 8716 5938
rect 8636 5800 8706 5806
rect 8758 5768 8824 5976
rect 8876 5938 8946 5944
rect 8866 5806 8876 5938
rect 8946 5806 8956 5938
rect 8876 5800 8946 5806
rect 8998 5768 9064 5976
rect 9116 5938 9186 5944
rect 9106 5806 9116 5938
rect 9186 5806 9196 5938
rect 9116 5800 9186 5806
rect 9238 5768 9304 5976
rect 9356 5938 9426 5944
rect 9346 5806 9356 5938
rect 9426 5806 9436 5938
rect 9356 5800 9426 5806
rect 9472 5768 9550 5976
rect 9596 5938 9666 5944
rect 9586 5806 9596 5938
rect 9666 5806 9676 5938
rect 9596 5800 9666 5806
rect 9718 5768 9784 5976
rect 9836 5938 9906 5944
rect 9826 5806 9836 5938
rect 9906 5806 9916 5938
rect 9836 5800 9906 5806
rect 9958 5768 10024 5976
rect 10076 5938 10146 5944
rect 10066 5806 10076 5938
rect 10146 5806 10156 5938
rect 10076 5800 10146 5806
rect 10198 5768 10264 5976
rect 10316 5938 10386 5944
rect 10306 5806 10316 5938
rect 10386 5806 10396 5938
rect 10316 5800 10386 5806
rect 10432 5768 10510 5976
rect 10556 5938 10626 5944
rect 10546 5806 10556 5938
rect 10626 5806 10636 5938
rect 10556 5800 10626 5806
rect 10678 5768 10744 5976
rect 10796 5938 10866 5944
rect 10786 5806 10796 5938
rect 10866 5806 10876 5938
rect 10796 5800 10866 5806
rect 10918 5768 10984 5976
rect 11036 5938 11106 5944
rect 11026 5806 11036 5938
rect 11106 5806 11116 5938
rect 11036 5800 11106 5806
rect 11158 5768 11224 5976
rect 11276 5938 11346 5944
rect 11266 5806 11276 5938
rect 11346 5806 11356 5938
rect 11276 5800 11346 5806
rect 11392 5768 11470 5976
rect 11516 5938 11586 5944
rect 11506 5806 11516 5938
rect 11586 5806 11596 5938
rect 11516 5800 11586 5806
rect 11638 5768 11704 5976
rect 11756 5938 11826 5944
rect 11746 5806 11756 5938
rect 11826 5806 11836 5938
rect 11756 5800 11826 5806
rect 11878 5768 11944 5976
rect 11996 5938 12066 5944
rect 11986 5806 11996 5938
rect 12066 5806 12076 5938
rect 11996 5800 12066 5806
rect 12118 5768 12184 5976
rect 12236 5938 12306 5944
rect 12226 5806 12236 5938
rect 12306 5806 12316 5938
rect 12236 5800 12306 5806
rect 12352 5768 12430 5976
rect 2752 5756 2870 5768
rect 2752 5180 2830 5756
rect 2864 5180 2870 5756
rect 2752 5168 2870 5180
rect 2952 5756 3110 5768
rect 2952 5180 2958 5756
rect 2992 5180 3070 5756
rect 3104 5180 3110 5756
rect 2952 5168 3110 5180
rect 3192 5756 3350 5768
rect 3192 5180 3198 5756
rect 3232 5180 3310 5756
rect 3344 5180 3350 5756
rect 3192 5168 3350 5180
rect 3432 5756 3590 5768
rect 3432 5180 3438 5756
rect 3472 5180 3550 5756
rect 3584 5180 3590 5756
rect 3432 5168 3590 5180
rect 3672 5756 3830 5768
rect 3672 5180 3678 5756
rect 3712 5180 3790 5756
rect 3824 5180 3830 5756
rect 3672 5168 3830 5180
rect 3912 5756 4070 5768
rect 3912 5180 3918 5756
rect 3952 5180 4030 5756
rect 4064 5180 4070 5756
rect 3912 5168 4070 5180
rect 4152 5756 4310 5768
rect 4152 5180 4158 5756
rect 4192 5180 4270 5756
rect 4304 5180 4310 5756
rect 4152 5168 4310 5180
rect 4392 5756 4550 5768
rect 4392 5180 4398 5756
rect 4432 5180 4510 5756
rect 4544 5180 4550 5756
rect 4392 5168 4550 5180
rect 4632 5756 4790 5768
rect 4632 5180 4638 5756
rect 4672 5180 4750 5756
rect 4784 5180 4790 5756
rect 4632 5168 4790 5180
rect 4872 5756 5030 5768
rect 4872 5180 4878 5756
rect 4912 5180 4990 5756
rect 5024 5180 5030 5756
rect 4872 5168 5030 5180
rect 5112 5756 5270 5768
rect 5112 5180 5118 5756
rect 5152 5180 5230 5756
rect 5264 5180 5270 5756
rect 5112 5168 5270 5180
rect 5352 5756 5510 5768
rect 5352 5180 5358 5756
rect 5392 5180 5470 5756
rect 5504 5180 5510 5756
rect 5352 5168 5510 5180
rect 5592 5756 5750 5768
rect 5592 5180 5598 5756
rect 5632 5180 5710 5756
rect 5744 5180 5750 5756
rect 5592 5168 5750 5180
rect 5832 5756 5990 5768
rect 5832 5180 5838 5756
rect 5872 5180 5950 5756
rect 5984 5180 5990 5756
rect 5832 5168 5990 5180
rect 6072 5756 6230 5768
rect 6072 5180 6078 5756
rect 6112 5180 6190 5756
rect 6224 5180 6230 5756
rect 6072 5168 6230 5180
rect 6312 5756 6470 5768
rect 6312 5180 6318 5756
rect 6352 5180 6430 5756
rect 6464 5180 6470 5756
rect 6312 5168 6470 5180
rect 6552 5756 6710 5768
rect 6552 5180 6558 5756
rect 6592 5180 6670 5756
rect 6704 5180 6710 5756
rect 6552 5168 6710 5180
rect 6792 5756 6950 5768
rect 6792 5180 6798 5756
rect 6832 5180 6910 5756
rect 6944 5180 6950 5756
rect 6792 5168 6950 5180
rect 7032 5756 7190 5768
rect 7032 5180 7038 5756
rect 7072 5180 7150 5756
rect 7184 5180 7190 5756
rect 7032 5168 7190 5180
rect 7272 5756 7430 5768
rect 7272 5180 7278 5756
rect 7312 5180 7390 5756
rect 7424 5180 7430 5756
rect 7272 5168 7430 5180
rect 7512 5756 7670 5768
rect 7512 5180 7518 5756
rect 7552 5180 7630 5756
rect 7664 5180 7670 5756
rect 7512 5168 7670 5180
rect 7752 5756 7910 5768
rect 7752 5180 7758 5756
rect 7792 5180 7870 5756
rect 7904 5180 7910 5756
rect 7752 5168 7910 5180
rect 7992 5756 8150 5768
rect 7992 5180 7998 5756
rect 8032 5180 8110 5756
rect 8144 5180 8150 5756
rect 7992 5168 8150 5180
rect 8232 5756 8390 5768
rect 8232 5180 8238 5756
rect 8272 5180 8350 5756
rect 8384 5180 8390 5756
rect 8232 5168 8390 5180
rect 8472 5756 8630 5768
rect 8472 5180 8478 5756
rect 8512 5180 8590 5756
rect 8624 5180 8630 5756
rect 8472 5168 8630 5180
rect 8712 5756 8870 5768
rect 8712 5180 8718 5756
rect 8752 5180 8830 5756
rect 8864 5180 8870 5756
rect 8712 5168 8870 5180
rect 8952 5756 9110 5768
rect 8952 5180 8958 5756
rect 8992 5180 9070 5756
rect 9104 5180 9110 5756
rect 8952 5168 9110 5180
rect 9192 5756 9350 5768
rect 9192 5180 9198 5756
rect 9232 5180 9310 5756
rect 9344 5180 9350 5756
rect 9192 5168 9350 5180
rect 9432 5756 9590 5768
rect 9432 5180 9438 5756
rect 9472 5180 9550 5756
rect 9584 5180 9590 5756
rect 9432 5168 9590 5180
rect 9672 5756 9830 5768
rect 9672 5180 9678 5756
rect 9712 5180 9790 5756
rect 9824 5180 9830 5756
rect 9672 5168 9830 5180
rect 9912 5756 10070 5768
rect 9912 5180 9918 5756
rect 9952 5180 10030 5756
rect 10064 5180 10070 5756
rect 9912 5168 10070 5180
rect 10152 5756 10310 5768
rect 10152 5180 10158 5756
rect 10192 5180 10270 5756
rect 10304 5180 10310 5756
rect 10152 5168 10310 5180
rect 10392 5756 10550 5768
rect 10392 5180 10398 5756
rect 10432 5180 10510 5756
rect 10544 5180 10550 5756
rect 10392 5168 10550 5180
rect 10632 5756 10790 5768
rect 10632 5180 10638 5756
rect 10672 5180 10750 5756
rect 10784 5180 10790 5756
rect 10632 5168 10790 5180
rect 10872 5756 11030 5768
rect 10872 5180 10878 5756
rect 10912 5180 10990 5756
rect 11024 5180 11030 5756
rect 10872 5168 11030 5180
rect 11112 5756 11270 5768
rect 11112 5180 11118 5756
rect 11152 5180 11230 5756
rect 11264 5180 11270 5756
rect 11112 5168 11270 5180
rect 11352 5756 11510 5768
rect 11352 5180 11358 5756
rect 11392 5180 11470 5756
rect 11504 5180 11510 5756
rect 11352 5168 11510 5180
rect 11592 5756 11750 5768
rect 11592 5180 11598 5756
rect 11632 5180 11710 5756
rect 11744 5180 11750 5756
rect 11592 5168 11750 5180
rect 11832 5756 11990 5768
rect 11832 5180 11838 5756
rect 11872 5180 11950 5756
rect 11984 5180 11990 5756
rect 11832 5168 11990 5180
rect 12072 5756 12230 5768
rect 12072 5180 12078 5756
rect 12112 5180 12190 5756
rect 12224 5180 12230 5756
rect 12072 5168 12230 5180
rect 12312 5756 12430 5768
rect 12312 5180 12318 5756
rect 12352 5180 12430 5756
rect 12312 5168 12430 5180
rect 2752 4302 2818 5168
rect 2876 5130 2946 5136
rect 3116 5130 3186 5136
rect 2866 4998 2876 5130
rect 2946 4998 2956 5130
rect 3106 4998 3116 5130
rect 3186 4998 3196 5130
rect 2876 4992 2946 4998
rect 3116 4992 3186 4998
rect 3244 4302 3298 5168
rect 3356 5130 3426 5136
rect 3596 5130 3666 5136
rect 3346 4998 3356 5130
rect 3426 4998 3436 5130
rect 3586 4998 3596 5130
rect 3666 4998 3676 5130
rect 3356 4992 3426 4998
rect 3596 4992 3666 4998
rect 3724 4302 3778 5168
rect 3836 5130 3906 5136
rect 4076 5130 4146 5136
rect 3826 4998 3836 5130
rect 3906 4998 3916 5130
rect 4066 4998 4076 5130
rect 4146 4998 4156 5130
rect 3836 4992 3906 4998
rect 4076 4992 4146 4998
rect 4204 4302 4258 5168
rect 4316 5130 4386 5136
rect 4556 5130 4626 5136
rect 4306 4998 4316 5130
rect 4386 4998 4396 5130
rect 4546 4998 4556 5130
rect 4626 4998 4636 5130
rect 4316 4992 4386 4998
rect 4556 4992 4626 4998
rect 4684 4302 4738 5168
rect 4796 5130 4866 5136
rect 5036 5130 5106 5136
rect 4786 4998 4796 5130
rect 4866 4998 4876 5130
rect 5026 4998 5036 5130
rect 5106 4998 5116 5130
rect 4796 4992 4866 4998
rect 5036 4992 5106 4998
rect 5164 4302 5218 5168
rect 5276 5130 5346 5136
rect 5516 5130 5586 5136
rect 5266 4998 5276 5130
rect 5346 4998 5356 5130
rect 5506 4998 5516 5130
rect 5586 4998 5596 5130
rect 5276 4992 5346 4998
rect 5516 4992 5586 4998
rect 5644 4302 5698 5168
rect 5756 5130 5826 5136
rect 5996 5130 6066 5136
rect 5746 4998 5756 5130
rect 5826 4998 5836 5130
rect 5986 4998 5996 5130
rect 6066 4998 6076 5130
rect 5756 4992 5826 4998
rect 5996 4992 6066 4998
rect 6124 4302 6178 5168
rect 6236 5130 6306 5136
rect 6476 5130 6546 5136
rect 6226 4998 6236 5130
rect 6306 4998 6316 5130
rect 6466 4998 6476 5130
rect 6546 4998 6556 5130
rect 6236 4992 6306 4998
rect 6476 4992 6546 4998
rect 6604 4302 6658 5168
rect 6716 5130 6786 5136
rect 6956 5130 7026 5136
rect 6706 4998 6716 5130
rect 6786 4998 6796 5130
rect 6946 4998 6956 5130
rect 7026 4998 7036 5130
rect 6716 4992 6786 4998
rect 6956 4992 7026 4998
rect 7084 4302 7138 5168
rect 7196 5130 7266 5136
rect 7436 5130 7506 5136
rect 7186 4998 7196 5130
rect 7266 4998 7276 5130
rect 7426 4998 7436 5130
rect 7506 4998 7516 5130
rect 7196 4992 7266 4998
rect 7436 4992 7506 4998
rect 7564 4302 7618 5168
rect 7676 5130 7746 5136
rect 7916 5130 7986 5136
rect 7666 4998 7676 5130
rect 7746 4998 7756 5130
rect 7906 4998 7916 5130
rect 7986 4998 7996 5130
rect 7676 4992 7746 4998
rect 7916 4992 7986 4998
rect 8044 4302 8098 5168
rect 8156 5130 8226 5136
rect 8396 5130 8466 5136
rect 8146 4998 8156 5130
rect 8226 4998 8236 5130
rect 8386 4998 8396 5130
rect 8466 4998 8476 5130
rect 8156 4992 8226 4998
rect 8396 4992 8466 4998
rect 8524 4302 8578 5168
rect 8636 5130 8706 5136
rect 8876 5130 8946 5136
rect 8626 4998 8636 5130
rect 8706 4998 8716 5130
rect 8866 4998 8876 5130
rect 8946 4998 8956 5130
rect 8636 4992 8706 4998
rect 8876 4992 8946 4998
rect 9004 4302 9058 5168
rect 9116 5130 9186 5136
rect 9356 5130 9426 5136
rect 9106 4998 9116 5130
rect 9186 4998 9196 5130
rect 9346 4998 9356 5130
rect 9426 4998 9436 5130
rect 9116 4992 9186 4998
rect 9356 4992 9426 4998
rect 9484 4302 9538 5168
rect 9596 5130 9666 5136
rect 9836 5130 9906 5136
rect 9586 4998 9596 5130
rect 9666 4998 9676 5130
rect 9826 4998 9836 5130
rect 9906 4998 9916 5130
rect 9596 4992 9666 4998
rect 9836 4992 9906 4998
rect 9964 4302 10018 5168
rect 10076 5130 10146 5136
rect 10316 5130 10386 5136
rect 10066 4998 10076 5130
rect 10146 4998 10156 5130
rect 10306 4998 10316 5130
rect 10386 4998 10396 5130
rect 10076 4992 10146 4998
rect 10316 4992 10386 4998
rect 10444 4302 10498 5168
rect 10556 5130 10626 5136
rect 10796 5130 10866 5136
rect 10546 4998 10556 5130
rect 10626 4998 10636 5130
rect 10786 4998 10796 5130
rect 10866 4998 10876 5130
rect 10556 4992 10626 4998
rect 10796 4992 10866 4998
rect 10924 4302 10978 5168
rect 11036 5130 11106 5136
rect 11276 5130 11346 5136
rect 11026 4998 11036 5130
rect 11106 4998 11116 5130
rect 11266 4998 11276 5130
rect 11346 4998 11356 5130
rect 11036 4992 11106 4998
rect 11276 4992 11346 4998
rect 11404 4302 11458 5168
rect 11516 5130 11586 5136
rect 11756 5130 11826 5136
rect 11506 4998 11516 5130
rect 11586 4998 11596 5130
rect 11746 4998 11756 5130
rect 11826 4998 11836 5130
rect 11516 4992 11586 4998
rect 11756 4992 11826 4998
rect 11884 4302 11938 5168
rect 11996 5130 12066 5136
rect 12236 5130 12306 5136
rect 11986 4998 11996 5130
rect 12066 4998 12076 5130
rect 12226 4998 12236 5130
rect 12306 4998 12316 5130
rect 11996 4992 12066 4998
rect 12236 4992 12306 4998
rect 12364 4302 12430 5168
rect -6564 4104 21744 4302
rect -6564 3560 16818 4104
rect 17718 3560 21744 4104
rect -6564 3394 21744 3560
rect -6564 2456 -6486 3394
rect -6424 2537 -6032 2543
rect -6424 2503 -6412 2537
rect -6044 2503 -6032 2537
rect -6424 2497 -6032 2503
rect -5836 2537 -5444 2543
rect -5836 2503 -5824 2537
rect -5456 2503 -5444 2537
rect -5836 2497 -5444 2503
rect -5382 2456 -5310 3394
rect -5248 2537 -4856 2543
rect -5248 2503 -5236 2537
rect -4868 2503 -4856 2537
rect -5248 2497 -4856 2503
rect -4660 2537 -4268 2543
rect -4660 2503 -4648 2537
rect -4280 2503 -4268 2537
rect -4660 2497 -4268 2503
rect -4206 2456 -4134 3394
rect -4072 2537 -3680 2543
rect -4072 2503 -4060 2537
rect -3692 2503 -3680 2537
rect -4072 2497 -3680 2503
rect -3484 2537 -3092 2543
rect -3484 2503 -3472 2537
rect -3104 2503 -3092 2537
rect -3484 2497 -3092 2503
rect -3030 2456 -2958 3394
rect -2896 2537 -2504 2543
rect -2896 2503 -2884 2537
rect -2516 2503 -2504 2537
rect -2896 2497 -2504 2503
rect -2308 2537 -1916 2543
rect -2308 2503 -2296 2537
rect -1928 2503 -1916 2537
rect -2308 2497 -1916 2503
rect -1854 2456 -1782 3394
rect -1720 2537 -1328 2543
rect -1720 2503 -1708 2537
rect -1340 2503 -1328 2537
rect -1720 2497 -1328 2503
rect -1132 2537 -740 2543
rect -1132 2503 -1120 2537
rect -752 2503 -740 2537
rect -1132 2497 -740 2503
rect -678 2456 -606 3394
rect -544 2537 -152 2543
rect -544 2503 -532 2537
rect -164 2503 -152 2537
rect -544 2497 -152 2503
rect 44 2537 436 2543
rect 44 2503 56 2537
rect 424 2503 436 2537
rect 44 2497 436 2503
rect 498 2456 570 3394
rect 632 2537 1024 2543
rect 632 2503 644 2537
rect 1012 2503 1024 2537
rect 632 2497 1024 2503
rect 1220 2537 1612 2543
rect 1220 2503 1232 2537
rect 1600 2503 1612 2537
rect 1220 2497 1612 2503
rect 1674 2456 1746 3394
rect 1808 2537 2200 2543
rect 1808 2503 1820 2537
rect 2188 2503 2200 2537
rect 1808 2497 2200 2503
rect 2396 2537 2788 2543
rect 2396 2503 2408 2537
rect 2776 2503 2788 2537
rect 2396 2497 2788 2503
rect 2850 2456 2922 3394
rect 2984 2537 3376 2543
rect 2984 2503 2996 2537
rect 3364 2503 3376 2537
rect 2984 2497 3376 2503
rect 3572 2537 3964 2543
rect 3572 2503 3584 2537
rect 3952 2503 3964 2537
rect 3572 2497 3964 2503
rect 4026 2456 4098 3394
rect 4160 2537 4552 2543
rect 4160 2503 4172 2537
rect 4540 2503 4552 2537
rect 4160 2497 4552 2503
rect 4748 2537 5140 2543
rect 4748 2503 4760 2537
rect 5128 2503 5140 2537
rect 4748 2497 5140 2503
rect 5174 2456 5246 3394
rect 5336 2537 5728 2543
rect 5336 2503 5348 2537
rect 5716 2503 5728 2537
rect 5336 2497 5728 2503
rect 5924 2537 6316 2543
rect 5924 2503 5936 2537
rect 6304 2503 6316 2537
rect 5924 2497 6316 2503
rect 6512 2537 6904 2543
rect 6512 2503 6524 2537
rect 6892 2503 6904 2537
rect 6512 2497 6904 2503
rect 7100 2537 7492 2543
rect 7100 2503 7112 2537
rect 7480 2503 7492 2537
rect 7100 2497 7492 2503
rect 7688 2537 8080 2543
rect 7688 2503 7700 2537
rect 8068 2503 8080 2537
rect 7688 2497 8080 2503
rect 8276 2537 8668 2543
rect 8276 2503 8288 2537
rect 8656 2503 8668 2537
rect 8276 2497 8668 2503
rect 8864 2537 9256 2543
rect 8864 2503 8876 2537
rect 9244 2503 9256 2537
rect 8864 2497 9256 2503
rect 9452 2537 9844 2543
rect 9452 2503 9464 2537
rect 9832 2503 9844 2537
rect 9452 2497 9844 2503
rect 9934 2456 10006 3394
rect 10040 2537 10432 2543
rect 10040 2503 10052 2537
rect 10420 2503 10432 2537
rect 10040 2497 10432 2503
rect 10628 2537 11020 2543
rect 10628 2503 10640 2537
rect 11008 2503 11020 2537
rect 10628 2497 11020 2503
rect 11082 2456 11154 3394
rect 11216 2537 11608 2543
rect 11216 2503 11228 2537
rect 11596 2503 11608 2537
rect 11216 2497 11608 2503
rect 11804 2537 12196 2543
rect 11804 2503 11816 2537
rect 12184 2503 12196 2537
rect 11804 2497 12196 2503
rect 12258 2456 12330 3394
rect 12392 2537 12784 2543
rect 12392 2503 12404 2537
rect 12772 2503 12784 2537
rect 12392 2497 12784 2503
rect 12980 2537 13372 2543
rect 12980 2503 12992 2537
rect 13360 2503 13372 2537
rect 12980 2497 13372 2503
rect 13434 2456 13506 3394
rect 13568 2537 13960 2543
rect 13568 2503 13580 2537
rect 13948 2503 13960 2537
rect 13568 2497 13960 2503
rect 14156 2537 14548 2543
rect 14156 2503 14168 2537
rect 14536 2503 14548 2537
rect 14156 2497 14548 2503
rect 14610 2456 14682 3394
rect 14744 2537 15136 2543
rect 14744 2503 14756 2537
rect 15124 2503 15136 2537
rect 14744 2497 15136 2503
rect 15332 2537 15724 2543
rect 15332 2503 15344 2537
rect 15712 2503 15724 2537
rect 15332 2497 15724 2503
rect 15786 2456 15858 3394
rect 15920 2537 16312 2543
rect 15920 2503 15932 2537
rect 16300 2503 16312 2537
rect 15920 2497 16312 2503
rect 16508 2537 16900 2543
rect 16508 2503 16520 2537
rect 16888 2503 16900 2537
rect 16508 2497 16900 2503
rect 16962 2456 17034 3394
rect 17096 2537 17488 2543
rect 17096 2503 17108 2537
rect 17476 2503 17488 2537
rect 17096 2497 17488 2503
rect 17684 2537 18076 2543
rect 17684 2503 17696 2537
rect 18064 2503 18076 2537
rect 17684 2497 18076 2503
rect 18138 2456 18210 3394
rect 18272 2537 18664 2543
rect 18272 2503 18284 2537
rect 18652 2503 18664 2537
rect 18272 2497 18664 2503
rect 18860 2537 19252 2543
rect 18860 2503 18872 2537
rect 19240 2503 19252 2537
rect 18860 2497 19252 2503
rect 19314 2456 19386 3394
rect 19448 2537 19840 2543
rect 19448 2503 19460 2537
rect 19828 2503 19840 2537
rect 19448 2497 19840 2503
rect 20036 2537 20428 2543
rect 20036 2503 20048 2537
rect 20416 2503 20428 2537
rect 20036 2497 20428 2503
rect 20490 2456 20562 3394
rect 20624 2537 21016 2543
rect 20624 2503 20636 2537
rect 21004 2503 21016 2537
rect 20624 2497 21016 2503
rect 21212 2537 21604 2543
rect 21212 2503 21224 2537
rect 21592 2503 21604 2537
rect 21212 2497 21604 2503
rect 21666 2456 21744 3394
rect -6564 2444 -6434 2456
rect -6564 1668 -6474 2444
rect -6440 1668 -6434 2444
rect -6564 1656 -6434 1668
rect -6022 2444 -5846 2456
rect -6022 1668 -6016 2444
rect -5982 1668 -5886 2444
rect -5852 1668 -5846 2444
rect -6022 1656 -5846 1668
rect -5434 2444 -5258 2456
rect -5434 1668 -5428 2444
rect -5394 1668 -5298 2444
rect -5264 1668 -5258 2444
rect -5434 1656 -5258 1668
rect -4846 2444 -4670 2456
rect -4846 1668 -4840 2444
rect -4806 1668 -4710 2444
rect -4676 1668 -4670 2444
rect -4846 1656 -4670 1668
rect -4258 2444 -4082 2456
rect -4258 1668 -4252 2444
rect -4218 1668 -4122 2444
rect -4088 1668 -4082 2444
rect -4258 1656 -4082 1668
rect -3670 2444 -3494 2456
rect -3670 1668 -3664 2444
rect -3630 1668 -3534 2444
rect -3500 1668 -3494 2444
rect -3670 1656 -3494 1668
rect -3082 2444 -2906 2456
rect -3082 1668 -3076 2444
rect -3042 1668 -2946 2444
rect -2912 1668 -2906 2444
rect -3082 1656 -2906 1668
rect -2494 2444 -2318 2456
rect -2494 1668 -2488 2444
rect -2454 1668 -2358 2444
rect -2324 1668 -2318 2444
rect -2494 1656 -2318 1668
rect -1906 2444 -1730 2456
rect -1906 1668 -1900 2444
rect -1866 1668 -1770 2444
rect -1736 1668 -1730 2444
rect -1906 1656 -1730 1668
rect -1318 2444 -1142 2456
rect -1318 1668 -1312 2444
rect -1278 1668 -1182 2444
rect -1148 1668 -1142 2444
rect -1318 1656 -1142 1668
rect -730 2444 -554 2456
rect -730 1668 -724 2444
rect -690 1668 -594 2444
rect -560 1668 -554 2444
rect -730 1656 -554 1668
rect -142 2444 34 2456
rect -142 1668 -136 2444
rect -102 1668 -6 2444
rect 28 1668 34 2444
rect -142 1656 34 1668
rect 446 2444 622 2456
rect 446 1668 452 2444
rect 486 1668 582 2444
rect 616 1668 622 2444
rect 446 1656 622 1668
rect 1034 2444 1210 2456
rect 1034 1668 1040 2444
rect 1074 1668 1170 2444
rect 1204 1668 1210 2444
rect 1034 1656 1210 1668
rect 1622 2444 1798 2456
rect 1622 1668 1628 2444
rect 1662 1668 1758 2444
rect 1792 1668 1798 2444
rect 1622 1656 1798 1668
rect 2210 2444 2386 2456
rect 2210 1668 2216 2444
rect 2250 1668 2346 2444
rect 2380 1668 2386 2444
rect 2210 1656 2386 1668
rect 2798 2444 2974 2456
rect 2798 1668 2804 2444
rect 2838 1668 2934 2444
rect 2968 1668 2974 2444
rect 2798 1656 2974 1668
rect 3386 2444 3562 2456
rect 3386 1668 3392 2444
rect 3426 1668 3522 2444
rect 3556 1668 3562 2444
rect 3386 1656 3562 1668
rect 3974 2444 4150 2456
rect 3974 1668 3980 2444
rect 4014 1668 4110 2444
rect 4144 1668 4150 2444
rect 3974 1656 4150 1668
rect 4562 2444 4738 2456
rect 4562 1668 4568 2444
rect 4602 1668 4698 2444
rect 4732 1668 4738 2444
rect 4562 1656 4738 1668
rect 5150 2444 5246 2456
rect 5150 1668 5156 2444
rect 5190 1720 5246 2444
rect 5280 2444 5326 2456
rect 5190 1668 5248 1720
rect 5150 1656 5248 1668
rect 5280 1668 5286 2444
rect 5320 1668 5326 2444
rect 5280 1656 5326 1668
rect 5738 2444 5914 2456
rect 5738 1668 5744 2444
rect 5778 1668 5874 2444
rect 5908 1668 5914 2444
rect 5738 1656 5914 1668
rect 6326 2444 6502 2456
rect 6326 1668 6332 2444
rect 6366 1668 6462 2444
rect 6496 1668 6502 2444
rect 6326 1656 6502 1668
rect 6914 2444 7090 2456
rect 6914 1668 6920 2444
rect 6954 1668 7050 2444
rect 7084 1668 7090 2444
rect 6914 1656 7090 1668
rect 7502 2444 7548 2456
rect 7502 1668 7508 2444
rect 7542 1668 7548 2444
rect 7502 1656 7548 1668
rect 7632 2444 7678 2456
rect 7632 1668 7638 2444
rect 7672 1668 7678 2444
rect 7632 1656 7678 1668
rect 8090 2444 8266 2456
rect 8090 1668 8096 2444
rect 8130 1668 8226 2444
rect 8260 1668 8266 2444
rect 8090 1656 8266 1668
rect 8678 2444 8854 2456
rect 8678 1668 8684 2444
rect 8718 1668 8814 2444
rect 8848 1668 8854 2444
rect 8678 1656 8854 1668
rect 9266 2444 9442 2456
rect 9266 1668 9272 2444
rect 9306 1668 9402 2444
rect 9436 1668 9442 2444
rect 9266 1656 9442 1668
rect 9854 2444 9900 2456
rect 9854 1668 9860 2444
rect 9894 1668 9900 2444
rect 9854 1656 9900 1668
rect 9934 2444 10030 2456
rect 9934 1668 9990 2444
rect 10024 1668 10030 2444
rect 9934 1656 10030 1668
rect 10442 2444 10618 2456
rect 10442 1668 10448 2444
rect 10482 1668 10578 2444
rect 10612 1668 10618 2444
rect 10442 1656 10618 1668
rect 11030 2444 11206 2456
rect 11030 1668 11036 2444
rect 11070 1668 11166 2444
rect 11200 1668 11206 2444
rect 11030 1656 11206 1668
rect 11618 2444 11794 2456
rect 11618 1668 11624 2444
rect 11658 1668 11754 2444
rect 11788 1668 11794 2444
rect 11618 1656 11794 1668
rect 12206 2444 12382 2456
rect 12206 1668 12212 2444
rect 12246 1668 12342 2444
rect 12376 1668 12382 2444
rect 12206 1656 12382 1668
rect 12794 2444 12970 2456
rect 12794 1668 12800 2444
rect 12834 1668 12930 2444
rect 12964 1668 12970 2444
rect 12794 1656 12970 1668
rect 13382 2444 13558 2456
rect 13382 1668 13388 2444
rect 13422 1668 13518 2444
rect 13552 1668 13558 2444
rect 13382 1656 13558 1668
rect 13970 2444 14146 2456
rect 13970 1668 13976 2444
rect 14010 1668 14106 2444
rect 14140 1668 14146 2444
rect 13970 1656 14146 1668
rect 14558 2444 14734 2456
rect 14558 1668 14564 2444
rect 14598 1668 14694 2444
rect 14728 1668 14734 2444
rect 14558 1656 14734 1668
rect 15146 2444 15322 2456
rect 15146 1668 15152 2444
rect 15186 1668 15282 2444
rect 15316 1668 15322 2444
rect 15146 1656 15322 1668
rect 15734 2444 15910 2456
rect 15734 1668 15740 2444
rect 15774 1668 15870 2444
rect 15904 1668 15910 2444
rect 15734 1656 15910 1668
rect 16322 2444 16498 2456
rect 16322 1668 16328 2444
rect 16362 1668 16458 2444
rect 16492 1668 16498 2444
rect 16322 1656 16498 1668
rect 16910 2444 17086 2456
rect 16910 1668 16916 2444
rect 16950 1668 17046 2444
rect 17080 1668 17086 2444
rect 16910 1656 17086 1668
rect 17498 2444 17674 2456
rect 17498 1668 17504 2444
rect 17538 1668 17634 2444
rect 17668 1668 17674 2444
rect 17498 1656 17674 1668
rect 18086 2444 18262 2456
rect 18086 1668 18092 2444
rect 18126 1668 18222 2444
rect 18256 1668 18262 2444
rect 18086 1656 18262 1668
rect 18674 2444 18850 2456
rect 18674 1668 18680 2444
rect 18714 1668 18810 2444
rect 18844 1668 18850 2444
rect 18674 1656 18850 1668
rect 19262 2444 19438 2456
rect 19262 1668 19268 2444
rect 19302 1668 19398 2444
rect 19432 1668 19438 2444
rect 19262 1656 19438 1668
rect 19850 2444 20026 2456
rect 19850 1668 19856 2444
rect 19890 1668 19986 2444
rect 20020 1668 20026 2444
rect 19850 1656 20026 1668
rect 20438 2444 20614 2456
rect 20438 1668 20444 2444
rect 20478 1668 20574 2444
rect 20608 1668 20614 2444
rect 20438 1656 20614 1668
rect 21026 2444 21202 2456
rect 21026 1668 21032 2444
rect 21066 1668 21162 2444
rect 21196 1668 21202 2444
rect 21026 1656 21202 1668
rect 21614 2444 21744 2456
rect 21614 1668 21620 2444
rect 21654 1668 21744 2444
rect 21614 1656 21744 1668
rect -6564 1456 -6480 1656
rect -6424 1609 -6032 1615
rect -6424 1575 -6412 1609
rect -6044 1575 -6032 1609
rect -6424 1537 -6032 1575
rect -6424 1503 -6412 1537
rect -6044 1503 -6032 1537
rect -6424 1497 -6032 1503
rect -5976 1456 -5892 1656
rect -5836 1609 -5444 1615
rect -5836 1575 -5824 1609
rect -5456 1575 -5444 1609
rect -5836 1537 -5444 1575
rect -5836 1503 -5824 1537
rect -5456 1503 -5444 1537
rect -5836 1497 -5444 1503
rect -5388 1456 -5304 1656
rect -5248 1609 -4856 1615
rect -5248 1575 -5236 1609
rect -4868 1575 -4856 1609
rect -5248 1537 -4856 1575
rect -5248 1503 -5236 1537
rect -4868 1503 -4856 1537
rect -5248 1497 -4856 1503
rect -4800 1456 -4716 1656
rect -4660 1609 -4268 1615
rect -4660 1575 -4648 1609
rect -4280 1575 -4268 1609
rect -4660 1537 -4268 1575
rect -4660 1503 -4648 1537
rect -4280 1503 -4268 1537
rect -4660 1497 -4268 1503
rect -4212 1456 -4128 1656
rect -4072 1609 -3680 1615
rect -4072 1575 -4060 1609
rect -3692 1575 -3680 1609
rect -4072 1537 -3680 1575
rect -4072 1503 -4060 1537
rect -3692 1503 -3680 1537
rect -4072 1497 -3680 1503
rect -3624 1456 -3540 1656
rect -3484 1609 -3092 1615
rect -3484 1575 -3472 1609
rect -3104 1575 -3092 1609
rect -3484 1537 -3092 1575
rect -3484 1503 -3472 1537
rect -3104 1503 -3092 1537
rect -3484 1497 -3092 1503
rect -3036 1456 -2952 1656
rect -2896 1609 -2504 1615
rect -2896 1575 -2884 1609
rect -2516 1575 -2504 1609
rect -2896 1537 -2504 1575
rect -2896 1503 -2884 1537
rect -2516 1503 -2504 1537
rect -2896 1497 -2504 1503
rect -2448 1456 -2364 1656
rect -2308 1609 -1916 1615
rect -2308 1575 -2296 1609
rect -1928 1575 -1916 1609
rect -2308 1537 -1916 1575
rect -2308 1503 -2296 1537
rect -1928 1503 -1916 1537
rect -2308 1497 -1916 1503
rect -1860 1456 -1776 1656
rect -1720 1609 -1328 1615
rect -1720 1575 -1708 1609
rect -1340 1575 -1328 1609
rect -1720 1537 -1328 1575
rect -1720 1503 -1708 1537
rect -1340 1503 -1328 1537
rect -1720 1497 -1328 1503
rect -1272 1456 -1188 1656
rect -1132 1609 -740 1615
rect -1132 1575 -1120 1609
rect -752 1575 -740 1609
rect -1132 1537 -740 1575
rect -1132 1503 -1120 1537
rect -752 1503 -740 1537
rect -1132 1497 -740 1503
rect -684 1456 -600 1656
rect -544 1609 -152 1615
rect -544 1575 -532 1609
rect -164 1575 -152 1609
rect -544 1537 -152 1575
rect -544 1503 -532 1537
rect -164 1503 -152 1537
rect -544 1497 -152 1503
rect -96 1456 -12 1656
rect 44 1609 436 1615
rect 44 1575 56 1609
rect 424 1575 436 1609
rect 44 1537 436 1575
rect 44 1503 56 1537
rect 424 1503 436 1537
rect 44 1497 436 1503
rect 492 1456 576 1656
rect 632 1609 1024 1615
rect 632 1575 644 1609
rect 1012 1575 1024 1609
rect 632 1537 1024 1575
rect 632 1503 644 1537
rect 1012 1503 1024 1537
rect 632 1497 1024 1503
rect 1080 1456 1164 1656
rect 1220 1609 1612 1615
rect 1220 1575 1232 1609
rect 1600 1575 1612 1609
rect 1220 1537 1612 1575
rect 1220 1503 1232 1537
rect 1600 1503 1612 1537
rect 1220 1497 1612 1503
rect 1668 1456 1752 1656
rect 1808 1609 2200 1615
rect 1808 1575 1820 1609
rect 2188 1575 2200 1609
rect 1808 1537 2200 1575
rect 1808 1503 1820 1537
rect 2188 1503 2200 1537
rect 1808 1497 2200 1503
rect 2256 1456 2340 1656
rect 2396 1609 2788 1615
rect 2396 1575 2408 1609
rect 2776 1575 2788 1609
rect 2396 1537 2788 1575
rect 2396 1503 2408 1537
rect 2776 1503 2788 1537
rect 2396 1497 2788 1503
rect 2844 1456 2928 1656
rect 2984 1609 3376 1615
rect 2984 1575 2996 1609
rect 3364 1575 3376 1609
rect 2984 1537 3376 1575
rect 2984 1503 2996 1537
rect 3364 1503 3376 1537
rect 2984 1497 3376 1503
rect 3432 1456 3516 1656
rect 3572 1609 3964 1615
rect 3572 1575 3584 1609
rect 3952 1575 3964 1609
rect 3572 1537 3964 1575
rect 3572 1503 3584 1537
rect 3952 1503 3964 1537
rect 3572 1497 3964 1503
rect 4020 1456 4104 1656
rect 4160 1609 4552 1615
rect 4160 1575 4172 1609
rect 4540 1575 4552 1609
rect 4160 1537 4552 1575
rect 4160 1503 4172 1537
rect 4540 1503 4552 1537
rect 4160 1497 4552 1503
rect 4608 1456 4692 1656
rect 4748 1609 5140 1615
rect 4748 1575 4760 1609
rect 5128 1575 5140 1609
rect 4748 1537 5140 1575
rect 4748 1503 4760 1537
rect 5128 1503 5140 1537
rect 4748 1497 5140 1503
rect 5190 1456 5248 1656
rect 5336 1609 5728 1615
rect 5336 1575 5348 1609
rect 5716 1575 5728 1609
rect 5336 1537 5728 1575
rect 5336 1503 5348 1537
rect 5716 1503 5728 1537
rect 5336 1497 5728 1503
rect 5784 1456 5868 1656
rect 5924 1609 6316 1615
rect 5924 1575 5936 1609
rect 6304 1575 6316 1609
rect 5924 1537 6316 1575
rect 5924 1503 5936 1537
rect 6304 1503 6316 1537
rect 5924 1497 6316 1503
rect 6372 1456 6456 1656
rect 6512 1609 6904 1615
rect 6512 1575 6524 1609
rect 6892 1575 6904 1609
rect 6512 1537 6904 1575
rect 6512 1503 6524 1537
rect 6892 1503 6904 1537
rect 6512 1497 6904 1503
rect 6960 1456 7044 1656
rect 7100 1609 7492 1615
rect 7100 1575 7112 1609
rect 7480 1575 7492 1609
rect 7100 1537 7492 1575
rect 7100 1503 7112 1537
rect 7480 1503 7492 1537
rect 7100 1497 7492 1503
rect 7688 1609 8080 1615
rect 7688 1575 7700 1609
rect 8068 1575 8080 1609
rect 7688 1537 8080 1575
rect 7688 1503 7700 1537
rect 8068 1503 8080 1537
rect 7688 1497 8080 1503
rect 8136 1456 8220 1656
rect 8276 1609 8668 1615
rect 8276 1575 8288 1609
rect 8656 1575 8668 1609
rect 8276 1537 8668 1575
rect 8276 1503 8288 1537
rect 8656 1503 8668 1537
rect 8276 1497 8668 1503
rect 8724 1456 8808 1656
rect 8864 1609 9256 1615
rect 8864 1575 8876 1609
rect 9244 1575 9256 1609
rect 8864 1537 9256 1575
rect 8864 1503 8876 1537
rect 9244 1503 9256 1537
rect 8864 1497 9256 1503
rect 9312 1456 9396 1656
rect 9452 1609 9844 1615
rect 9452 1575 9464 1609
rect 9832 1575 9844 1609
rect 9452 1537 9844 1575
rect 9452 1503 9464 1537
rect 9832 1503 9844 1537
rect 9452 1497 9844 1503
rect 9934 1456 9990 1656
rect 10040 1609 10432 1615
rect 10040 1575 10052 1609
rect 10420 1575 10432 1609
rect 10040 1537 10432 1575
rect 10040 1503 10052 1537
rect 10420 1503 10432 1537
rect 10040 1497 10432 1503
rect 10488 1456 10572 1656
rect 10628 1609 11020 1615
rect 10628 1575 10640 1609
rect 11008 1575 11020 1609
rect 10628 1537 11020 1575
rect 10628 1503 10640 1537
rect 11008 1503 11020 1537
rect 10628 1497 11020 1503
rect 11076 1456 11160 1656
rect 11216 1609 11608 1615
rect 11216 1575 11228 1609
rect 11596 1575 11608 1609
rect 11216 1537 11608 1575
rect 11216 1503 11228 1537
rect 11596 1503 11608 1537
rect 11216 1497 11608 1503
rect 11664 1456 11748 1656
rect 11804 1609 12196 1615
rect 11804 1575 11816 1609
rect 12184 1575 12196 1609
rect 11804 1537 12196 1575
rect 11804 1503 11816 1537
rect 12184 1503 12196 1537
rect 11804 1497 12196 1503
rect 12252 1456 12336 1656
rect 12392 1609 12784 1615
rect 12392 1575 12404 1609
rect 12772 1575 12784 1609
rect 12392 1537 12784 1575
rect 12392 1503 12404 1537
rect 12772 1503 12784 1537
rect 12392 1497 12784 1503
rect 12840 1456 12924 1656
rect 12980 1609 13372 1615
rect 12980 1575 12992 1609
rect 13360 1575 13372 1609
rect 12980 1537 13372 1575
rect 12980 1503 12992 1537
rect 13360 1503 13372 1537
rect 12980 1497 13372 1503
rect 13428 1456 13512 1656
rect 13568 1609 13960 1615
rect 13568 1575 13580 1609
rect 13948 1575 13960 1609
rect 13568 1537 13960 1575
rect 13568 1503 13580 1537
rect 13948 1503 13960 1537
rect 13568 1497 13960 1503
rect 14016 1456 14100 1656
rect 14156 1609 14548 1615
rect 14156 1575 14168 1609
rect 14536 1575 14548 1609
rect 14156 1537 14548 1575
rect 14156 1503 14168 1537
rect 14536 1503 14548 1537
rect 14156 1497 14548 1503
rect 14604 1456 14688 1656
rect 14744 1609 15136 1615
rect 14744 1575 14756 1609
rect 15124 1575 15136 1609
rect 14744 1537 15136 1575
rect 14744 1503 14756 1537
rect 15124 1503 15136 1537
rect 14744 1497 15136 1503
rect 15192 1456 15276 1656
rect 15332 1609 15724 1615
rect 15332 1575 15344 1609
rect 15712 1575 15724 1609
rect 15332 1537 15724 1575
rect 15332 1503 15344 1537
rect 15712 1503 15724 1537
rect 15332 1497 15724 1503
rect 15780 1456 15864 1656
rect 15920 1609 16312 1615
rect 15920 1575 15932 1609
rect 16300 1575 16312 1609
rect 15920 1537 16312 1575
rect 15920 1503 15932 1537
rect 16300 1503 16312 1537
rect 15920 1497 16312 1503
rect 16368 1456 16452 1656
rect 16508 1609 16900 1615
rect 16508 1575 16520 1609
rect 16888 1575 16900 1609
rect 16508 1537 16900 1575
rect 16508 1503 16520 1537
rect 16888 1503 16900 1537
rect 16508 1497 16900 1503
rect 16956 1456 17040 1656
rect 17096 1609 17488 1615
rect 17096 1575 17108 1609
rect 17476 1575 17488 1609
rect 17096 1537 17488 1575
rect 17096 1503 17108 1537
rect 17476 1503 17488 1537
rect 17096 1497 17488 1503
rect 17544 1456 17628 1656
rect 17684 1609 18076 1615
rect 17684 1575 17696 1609
rect 18064 1575 18076 1609
rect 17684 1537 18076 1575
rect 17684 1503 17696 1537
rect 18064 1503 18076 1537
rect 17684 1497 18076 1503
rect 18132 1456 18216 1656
rect 18272 1609 18664 1615
rect 18272 1575 18284 1609
rect 18652 1575 18664 1609
rect 18272 1537 18664 1575
rect 18272 1503 18284 1537
rect 18652 1503 18664 1537
rect 18272 1497 18664 1503
rect 18720 1456 18804 1656
rect 18860 1609 19252 1615
rect 18860 1575 18872 1609
rect 19240 1575 19252 1609
rect 18860 1537 19252 1575
rect 18860 1503 18872 1537
rect 19240 1503 19252 1537
rect 18860 1497 19252 1503
rect 19308 1456 19392 1656
rect 19448 1609 19840 1615
rect 19448 1575 19460 1609
rect 19828 1575 19840 1609
rect 19448 1537 19840 1575
rect 19448 1503 19460 1537
rect 19828 1503 19840 1537
rect 19448 1497 19840 1503
rect 19896 1456 19980 1656
rect 20036 1609 20428 1615
rect 20036 1575 20048 1609
rect 20416 1575 20428 1609
rect 20036 1537 20428 1575
rect 20036 1503 20048 1537
rect 20416 1503 20428 1537
rect 20036 1497 20428 1503
rect 20484 1456 20568 1656
rect 20624 1609 21016 1615
rect 20624 1575 20636 1609
rect 21004 1575 21016 1609
rect 20624 1537 21016 1575
rect 20624 1503 20636 1537
rect 21004 1503 21016 1537
rect 20624 1497 21016 1503
rect 21072 1456 21156 1656
rect 21212 1609 21604 1615
rect 21212 1575 21224 1609
rect 21592 1575 21604 1609
rect 21212 1537 21604 1575
rect 21212 1503 21224 1537
rect 21592 1503 21604 1537
rect 21212 1497 21604 1503
rect 21660 1456 21744 1656
rect -6564 1444 -6434 1456
rect -6564 668 -6474 1444
rect -6440 668 -6434 1444
rect -6564 656 -6434 668
rect -6022 1444 -5846 1456
rect -6022 668 -6016 1444
rect -5982 668 -5886 1444
rect -5852 668 -5846 1444
rect -6022 656 -5846 668
rect -5434 1444 -5258 1456
rect -5434 668 -5428 1444
rect -5394 668 -5298 1444
rect -5264 668 -5258 1444
rect -5434 656 -5258 668
rect -4846 1444 -4670 1456
rect -4846 668 -4840 1444
rect -4806 668 -4710 1444
rect -4676 668 -4670 1444
rect -4846 656 -4670 668
rect -4258 1444 -4082 1456
rect -4258 668 -4252 1444
rect -4218 668 -4122 1444
rect -4088 668 -4082 1444
rect -4258 656 -4082 668
rect -3670 1444 -3494 1456
rect -3670 668 -3664 1444
rect -3630 668 -3534 1444
rect -3500 668 -3494 1444
rect -3670 656 -3494 668
rect -3082 1444 -2906 1456
rect -3082 668 -3076 1444
rect -3042 668 -2946 1444
rect -2912 668 -2906 1444
rect -3082 656 -2906 668
rect -2494 1444 -2318 1456
rect -2494 668 -2488 1444
rect -2454 668 -2358 1444
rect -2324 668 -2318 1444
rect -2494 656 -2318 668
rect -1906 1444 -1730 1456
rect -1906 668 -1900 1444
rect -1866 668 -1770 1444
rect -1736 668 -1730 1444
rect -1906 656 -1730 668
rect -1318 1444 -1142 1456
rect -1318 668 -1312 1444
rect -1278 668 -1182 1444
rect -1148 668 -1142 1444
rect -1318 656 -1142 668
rect -730 1444 -554 1456
rect -730 668 -724 1444
rect -690 668 -594 1444
rect -560 668 -554 1444
rect -730 656 -554 668
rect -142 1444 34 1456
rect -142 668 -136 1444
rect -102 668 -6 1444
rect 28 668 34 1444
rect -142 656 34 668
rect 446 1444 622 1456
rect 446 668 452 1444
rect 486 668 582 1444
rect 616 668 622 1444
rect 446 656 622 668
rect 1034 1444 1210 1456
rect 1034 668 1040 1444
rect 1074 668 1170 1444
rect 1204 668 1210 1444
rect 1034 656 1210 668
rect 1622 1444 1798 1456
rect 1622 668 1628 1444
rect 1662 668 1758 1444
rect 1792 668 1798 1444
rect 1622 656 1798 668
rect 2210 1444 2386 1456
rect 2210 668 2216 1444
rect 2250 668 2346 1444
rect 2380 668 2386 1444
rect 2210 656 2386 668
rect 2798 1444 2974 1456
rect 2798 668 2804 1444
rect 2838 668 2934 1444
rect 2968 668 2974 1444
rect 2798 656 2974 668
rect 3386 1444 3562 1456
rect 3386 668 3392 1444
rect 3426 668 3522 1444
rect 3556 668 3562 1444
rect 3386 656 3562 668
rect 3974 1444 4150 1456
rect 3974 668 3980 1444
rect 4014 668 4110 1444
rect 4144 668 4150 1444
rect 3974 656 4150 668
rect 4562 1444 4738 1456
rect 4562 668 4568 1444
rect 4602 668 4698 1444
rect 4732 668 4738 1444
rect 4562 656 4738 668
rect 5150 1444 5248 1456
rect 5150 668 5156 1444
rect 5190 668 5248 1444
rect 5150 656 5248 668
rect 5280 1444 5326 1456
rect 5280 668 5286 1444
rect 5320 668 5326 1444
rect 5280 656 5326 668
rect 5738 1444 5914 1456
rect 5738 668 5744 1444
rect 5778 668 5874 1444
rect 5908 668 5914 1444
rect 5738 656 5914 668
rect 6326 1444 6502 1456
rect 6326 668 6332 1444
rect 6366 668 6462 1444
rect 6496 668 6502 1444
rect 6326 656 6502 668
rect 6914 1444 7090 1456
rect 6914 668 6920 1444
rect 6954 668 7050 1444
rect 7084 668 7090 1444
rect 6914 656 7090 668
rect 7502 1444 7548 1456
rect 7502 668 7508 1444
rect 7542 668 7548 1444
rect 7502 656 7548 668
rect 7632 1444 7678 1456
rect 7632 668 7638 1444
rect 7672 668 7678 1444
rect 7632 656 7678 668
rect 8090 1444 8266 1456
rect 8090 668 8096 1444
rect 8130 668 8226 1444
rect 8260 668 8266 1444
rect 8090 656 8266 668
rect 8678 1444 8854 1456
rect 8678 668 8684 1444
rect 8718 668 8814 1444
rect 8848 668 8854 1444
rect 8678 656 8854 668
rect 9266 1444 9442 1456
rect 9266 668 9272 1444
rect 9306 668 9402 1444
rect 9436 668 9442 1444
rect 9266 656 9442 668
rect 9854 1444 9900 1456
rect 9854 668 9860 1444
rect 9894 668 9900 1444
rect 9854 656 9900 668
rect 9934 1444 10030 1456
rect 9934 668 9990 1444
rect 10024 668 10030 1444
rect 9934 656 10030 668
rect 10442 1444 10618 1456
rect 10442 668 10448 1444
rect 10482 668 10578 1444
rect 10612 668 10618 1444
rect 10442 656 10618 668
rect 11030 1444 11206 1456
rect 11030 668 11036 1444
rect 11070 668 11166 1444
rect 11200 668 11206 1444
rect 11030 656 11206 668
rect 11618 1444 11794 1456
rect 11618 668 11624 1444
rect 11658 668 11754 1444
rect 11788 668 11794 1444
rect 11618 656 11794 668
rect 12206 1444 12382 1456
rect 12206 668 12212 1444
rect 12246 668 12342 1444
rect 12376 668 12382 1444
rect 12206 656 12382 668
rect 12794 1444 12970 1456
rect 12794 668 12800 1444
rect 12834 668 12930 1444
rect 12964 668 12970 1444
rect 12794 656 12970 668
rect 13382 1444 13558 1456
rect 13382 668 13388 1444
rect 13422 668 13518 1444
rect 13552 668 13558 1444
rect 13382 656 13558 668
rect 13970 1444 14146 1456
rect 13970 668 13976 1444
rect 14010 668 14106 1444
rect 14140 668 14146 1444
rect 13970 656 14146 668
rect 14558 1444 14734 1456
rect 14558 668 14564 1444
rect 14598 668 14694 1444
rect 14728 668 14734 1444
rect 14558 656 14734 668
rect 15146 1444 15322 1456
rect 15146 668 15152 1444
rect 15186 668 15282 1444
rect 15316 668 15322 1444
rect 15146 656 15322 668
rect 15734 1444 15910 1456
rect 15734 668 15740 1444
rect 15774 668 15870 1444
rect 15904 668 15910 1444
rect 15734 656 15910 668
rect 16322 1444 16498 1456
rect 16322 668 16328 1444
rect 16362 668 16458 1444
rect 16492 668 16498 1444
rect 16322 656 16498 668
rect 16910 1444 17086 1456
rect 16910 668 16916 1444
rect 16950 668 17046 1444
rect 17080 668 17086 1444
rect 16910 656 17086 668
rect 17498 1444 17674 1456
rect 17498 668 17504 1444
rect 17538 668 17634 1444
rect 17668 668 17674 1444
rect 17498 656 17674 668
rect 18086 1444 18262 1456
rect 18086 668 18092 1444
rect 18126 668 18222 1444
rect 18256 668 18262 1444
rect 18086 656 18262 668
rect 18674 1444 18850 1456
rect 18674 668 18680 1444
rect 18714 668 18810 1444
rect 18844 668 18850 1444
rect 18674 656 18850 668
rect 19262 1444 19438 1456
rect 19262 668 19268 1444
rect 19302 668 19398 1444
rect 19432 668 19438 1444
rect 19262 656 19438 668
rect 19850 1444 20026 1456
rect 19850 668 19856 1444
rect 19890 668 19986 1444
rect 20020 668 20026 1444
rect 19850 656 20026 668
rect 20438 1444 20614 1456
rect 20438 668 20444 1444
rect 20478 668 20574 1444
rect 20608 668 20614 1444
rect 20438 656 20614 668
rect 21026 1444 21202 1456
rect 21026 668 21032 1444
rect 21066 668 21162 1444
rect 21196 668 21202 1444
rect 21026 656 21202 668
rect 21614 1444 21744 1456
rect 21614 668 21620 1444
rect 21654 668 21744 1444
rect 21614 656 21744 668
rect -6564 456 -6480 656
rect -6424 609 -6032 615
rect -6424 575 -6412 609
rect -6044 575 -6032 609
rect -6424 537 -6032 575
rect -6424 503 -6412 537
rect -6044 503 -6032 537
rect -6424 497 -6032 503
rect -5976 456 -5892 656
rect -5836 609 -5444 615
rect -5836 575 -5824 609
rect -5456 575 -5444 609
rect -5836 537 -5444 575
rect -5836 503 -5824 537
rect -5456 503 -5444 537
rect -5836 497 -5444 503
rect -5388 456 -5304 656
rect -5248 609 -4856 615
rect -5248 575 -5236 609
rect -4868 575 -4856 609
rect -5248 537 -4856 575
rect -5248 503 -5236 537
rect -4868 503 -4856 537
rect -5248 497 -4856 503
rect -4800 456 -4716 656
rect -4660 609 -4268 615
rect -4660 575 -4648 609
rect -4280 575 -4268 609
rect -4660 537 -4268 575
rect -4660 503 -4648 537
rect -4280 503 -4268 537
rect -4660 497 -4268 503
rect -4212 456 -4128 656
rect -4072 609 -3680 615
rect -4072 575 -4060 609
rect -3692 575 -3680 609
rect -4072 537 -3680 575
rect -4072 503 -4060 537
rect -3692 503 -3680 537
rect -4072 497 -3680 503
rect -3624 456 -3540 656
rect -3484 609 -3092 615
rect -3484 575 -3472 609
rect -3104 575 -3092 609
rect -3484 537 -3092 575
rect -3484 503 -3472 537
rect -3104 503 -3092 537
rect -3484 497 -3092 503
rect -3036 456 -2952 656
rect -2896 609 -2504 615
rect -2896 575 -2884 609
rect -2516 575 -2504 609
rect -2896 537 -2504 575
rect -2896 503 -2884 537
rect -2516 503 -2504 537
rect -2896 497 -2504 503
rect -2448 456 -2364 656
rect -2308 609 -1916 615
rect -2308 575 -2296 609
rect -1928 575 -1916 609
rect -2308 537 -1916 575
rect -2308 503 -2296 537
rect -1928 503 -1916 537
rect -2308 497 -1916 503
rect -1860 456 -1776 656
rect -1720 609 -1328 615
rect -1720 575 -1708 609
rect -1340 575 -1328 609
rect -1720 537 -1328 575
rect -1720 503 -1708 537
rect -1340 503 -1328 537
rect -1720 497 -1328 503
rect -1272 456 -1188 656
rect -1132 609 -740 615
rect -1132 575 -1120 609
rect -752 575 -740 609
rect -1132 537 -740 575
rect -1132 503 -1120 537
rect -752 503 -740 537
rect -1132 497 -740 503
rect -684 456 -600 656
rect -544 609 -152 615
rect -544 575 -532 609
rect -164 575 -152 609
rect -544 537 -152 575
rect -544 503 -532 537
rect -164 503 -152 537
rect -544 497 -152 503
rect -96 456 -12 656
rect 44 609 436 615
rect 44 575 56 609
rect 424 575 436 609
rect 44 537 436 575
rect 44 503 56 537
rect 424 503 436 537
rect 44 497 436 503
rect 492 456 576 656
rect 632 609 1024 615
rect 632 575 644 609
rect 1012 575 1024 609
rect 632 537 1024 575
rect 632 503 644 537
rect 1012 503 1024 537
rect 632 497 1024 503
rect 1080 456 1164 656
rect 1220 609 1612 615
rect 1220 575 1232 609
rect 1600 575 1612 609
rect 1220 537 1612 575
rect 1220 503 1232 537
rect 1600 503 1612 537
rect 1220 497 1612 503
rect 1668 456 1752 656
rect 1808 609 2200 615
rect 1808 575 1820 609
rect 2188 575 2200 609
rect 1808 537 2200 575
rect 1808 503 1820 537
rect 2188 503 2200 537
rect 1808 497 2200 503
rect 2256 456 2340 656
rect 2396 609 2788 615
rect 2396 575 2408 609
rect 2776 575 2788 609
rect 2396 537 2788 575
rect 2396 503 2408 537
rect 2776 503 2788 537
rect 2396 497 2788 503
rect 2844 456 2928 656
rect 2984 609 3376 615
rect 2984 575 2996 609
rect 3364 575 3376 609
rect 2984 537 3376 575
rect 2984 503 2996 537
rect 3364 503 3376 537
rect 2984 497 3376 503
rect 3432 456 3516 656
rect 3572 609 3964 615
rect 3572 575 3584 609
rect 3952 575 3964 609
rect 3572 537 3964 575
rect 3572 503 3584 537
rect 3952 503 3964 537
rect 3572 497 3964 503
rect 4020 456 4104 656
rect 4160 609 4552 615
rect 4160 575 4172 609
rect 4540 575 4552 609
rect 4160 537 4552 575
rect 4160 503 4172 537
rect 4540 503 4552 537
rect 4160 497 4552 503
rect 4608 456 4692 656
rect 4748 609 5140 615
rect 4748 575 4760 609
rect 5128 575 5140 609
rect 4748 537 5140 575
rect 4748 503 4760 537
rect 5128 503 5140 537
rect 4748 497 5140 503
rect 5190 456 5248 656
rect 5336 609 5728 615
rect 5336 575 5348 609
rect 5716 575 5728 609
rect 5336 537 5728 575
rect 5336 503 5348 537
rect 5716 503 5728 537
rect 5336 497 5728 503
rect 5784 456 5868 656
rect 5924 609 6316 615
rect 5924 575 5936 609
rect 6304 575 6316 609
rect 5924 537 6316 575
rect 5924 503 5936 537
rect 6304 503 6316 537
rect 5924 497 6316 503
rect 6372 456 6456 656
rect 6512 609 6904 615
rect 6512 575 6524 609
rect 6892 575 6904 609
rect 6512 537 6904 575
rect 6512 503 6524 537
rect 6892 503 6904 537
rect 6512 497 6904 503
rect 6960 456 7044 656
rect 7100 609 7492 615
rect 7100 575 7112 609
rect 7480 575 7492 609
rect 7100 537 7492 575
rect 7100 503 7112 537
rect 7480 503 7492 537
rect 7100 497 7492 503
rect 7688 609 8080 615
rect 7688 575 7700 609
rect 8068 575 8080 609
rect 7688 537 8080 575
rect 7688 503 7700 537
rect 8068 503 8080 537
rect 7688 497 8080 503
rect 8136 456 8220 656
rect 8276 609 8668 615
rect 8276 575 8288 609
rect 8656 575 8668 609
rect 8276 537 8668 575
rect 8276 503 8288 537
rect 8656 503 8668 537
rect 8276 497 8668 503
rect 8724 456 8808 656
rect 8864 609 9256 615
rect 8864 575 8876 609
rect 9244 575 9256 609
rect 8864 537 9256 575
rect 8864 503 8876 537
rect 9244 503 9256 537
rect 8864 497 9256 503
rect 9312 456 9396 656
rect 9452 609 9844 615
rect 9452 575 9464 609
rect 9832 575 9844 609
rect 9452 537 9844 575
rect 9452 503 9464 537
rect 9832 503 9844 537
rect 9452 497 9844 503
rect 9934 456 9990 656
rect 10040 609 10432 615
rect 10040 575 10052 609
rect 10420 575 10432 609
rect 10040 537 10432 575
rect 10040 503 10052 537
rect 10420 503 10432 537
rect 10040 497 10432 503
rect 10488 456 10572 656
rect 10628 609 11020 615
rect 10628 575 10640 609
rect 11008 575 11020 609
rect 10628 537 11020 575
rect 10628 503 10640 537
rect 11008 503 11020 537
rect 10628 497 11020 503
rect 11076 456 11160 656
rect 11216 609 11608 615
rect 11216 575 11228 609
rect 11596 575 11608 609
rect 11216 537 11608 575
rect 11216 503 11228 537
rect 11596 503 11608 537
rect 11216 497 11608 503
rect 11664 456 11748 656
rect 11804 609 12196 615
rect 11804 575 11816 609
rect 12184 575 12196 609
rect 11804 537 12196 575
rect 11804 503 11816 537
rect 12184 503 12196 537
rect 11804 497 12196 503
rect 12252 456 12336 656
rect 12392 609 12784 615
rect 12392 575 12404 609
rect 12772 575 12784 609
rect 12392 537 12784 575
rect 12392 503 12404 537
rect 12772 503 12784 537
rect 12392 497 12784 503
rect 12840 456 12924 656
rect 12980 609 13372 615
rect 12980 575 12992 609
rect 13360 575 13372 609
rect 12980 537 13372 575
rect 12980 503 12992 537
rect 13360 503 13372 537
rect 12980 497 13372 503
rect 13428 456 13512 656
rect 13568 609 13960 615
rect 13568 575 13580 609
rect 13948 575 13960 609
rect 13568 537 13960 575
rect 13568 503 13580 537
rect 13948 503 13960 537
rect 13568 497 13960 503
rect 14016 456 14100 656
rect 14156 609 14548 615
rect 14156 575 14168 609
rect 14536 575 14548 609
rect 14156 537 14548 575
rect 14156 503 14168 537
rect 14536 503 14548 537
rect 14156 497 14548 503
rect 14604 456 14688 656
rect 14744 609 15136 615
rect 14744 575 14756 609
rect 15124 575 15136 609
rect 14744 537 15136 575
rect 14744 503 14756 537
rect 15124 503 15136 537
rect 14744 497 15136 503
rect 15192 456 15276 656
rect 15332 609 15724 615
rect 15332 575 15344 609
rect 15712 575 15724 609
rect 15332 537 15724 575
rect 15332 503 15344 537
rect 15712 503 15724 537
rect 15332 497 15724 503
rect 15780 456 15864 656
rect 15920 609 16312 615
rect 15920 575 15932 609
rect 16300 575 16312 609
rect 15920 537 16312 575
rect 15920 503 15932 537
rect 16300 503 16312 537
rect 15920 497 16312 503
rect 16368 456 16452 656
rect 16508 609 16900 615
rect 16508 575 16520 609
rect 16888 575 16900 609
rect 16508 537 16900 575
rect 16508 503 16520 537
rect 16888 503 16900 537
rect 16508 497 16900 503
rect 16956 456 17040 656
rect 17096 609 17488 615
rect 17096 575 17108 609
rect 17476 575 17488 609
rect 17096 537 17488 575
rect 17096 503 17108 537
rect 17476 503 17488 537
rect 17096 497 17488 503
rect 17544 456 17628 656
rect 17684 609 18076 615
rect 17684 575 17696 609
rect 18064 575 18076 609
rect 17684 537 18076 575
rect 17684 503 17696 537
rect 18064 503 18076 537
rect 17684 497 18076 503
rect 18132 456 18216 656
rect 18272 609 18664 615
rect 18272 575 18284 609
rect 18652 575 18664 609
rect 18272 537 18664 575
rect 18272 503 18284 537
rect 18652 503 18664 537
rect 18272 497 18664 503
rect 18720 456 18804 656
rect 18860 609 19252 615
rect 18860 575 18872 609
rect 19240 575 19252 609
rect 18860 537 19252 575
rect 18860 503 18872 537
rect 19240 503 19252 537
rect 18860 497 19252 503
rect 19308 456 19392 656
rect 19448 609 19840 615
rect 19448 575 19460 609
rect 19828 575 19840 609
rect 19448 537 19840 575
rect 19448 503 19460 537
rect 19828 503 19840 537
rect 19448 497 19840 503
rect 19896 456 19980 656
rect 20036 609 20428 615
rect 20036 575 20048 609
rect 20416 575 20428 609
rect 20036 537 20428 575
rect 20036 503 20048 537
rect 20416 503 20428 537
rect 20036 497 20428 503
rect 20484 456 20568 656
rect 20624 609 21016 615
rect 20624 575 20636 609
rect 21004 575 21016 609
rect 20624 537 21016 575
rect 20624 503 20636 537
rect 21004 503 21016 537
rect 20624 497 21016 503
rect 21072 456 21156 656
rect 21212 609 21604 615
rect 21212 575 21224 609
rect 21592 575 21604 609
rect 21212 537 21604 575
rect 21212 503 21224 537
rect 21592 503 21604 537
rect 21212 497 21604 503
rect 21660 456 21744 656
rect -6564 444 -6434 456
rect -6564 -332 -6474 444
rect -6440 -332 -6434 444
rect -6564 -344 -6434 -332
rect -6022 444 -5846 456
rect -6022 -332 -6016 444
rect -5982 -332 -5886 444
rect -5852 -332 -5846 444
rect -6022 -344 -5846 -332
rect -5434 444 -5258 456
rect -5434 -332 -5428 444
rect -5394 -332 -5298 444
rect -5264 -332 -5258 444
rect -5434 -344 -5258 -332
rect -4846 444 -4670 456
rect -4846 -332 -4840 444
rect -4806 -332 -4710 444
rect -4676 -332 -4670 444
rect -4846 -344 -4670 -332
rect -4258 444 -4082 456
rect -4258 -332 -4252 444
rect -4218 -332 -4122 444
rect -4088 -332 -4082 444
rect -4258 -344 -4082 -332
rect -3670 444 -3494 456
rect -3670 -332 -3664 444
rect -3630 -332 -3534 444
rect -3500 -332 -3494 444
rect -3670 -344 -3494 -332
rect -3082 444 -2906 456
rect -3082 -332 -3076 444
rect -3042 -332 -2946 444
rect -2912 -332 -2906 444
rect -3082 -344 -2906 -332
rect -2494 444 -2318 456
rect -2494 -332 -2488 444
rect -2454 -332 -2358 444
rect -2324 -332 -2318 444
rect -2494 -344 -2318 -332
rect -1906 444 -1730 456
rect -1906 -332 -1900 444
rect -1866 -332 -1770 444
rect -1736 -332 -1730 444
rect -1906 -344 -1730 -332
rect -1318 444 -1142 456
rect -1318 -332 -1312 444
rect -1278 -332 -1182 444
rect -1148 -332 -1142 444
rect -1318 -344 -1142 -332
rect -730 444 -554 456
rect -730 -332 -724 444
rect -690 -332 -594 444
rect -560 -332 -554 444
rect -730 -344 -554 -332
rect -142 444 34 456
rect -142 -332 -136 444
rect -102 -332 -6 444
rect 28 -332 34 444
rect -142 -344 34 -332
rect 446 444 622 456
rect 446 -332 452 444
rect 486 -332 582 444
rect 616 -332 622 444
rect 446 -344 622 -332
rect 1034 444 1210 456
rect 1034 -332 1040 444
rect 1074 -332 1170 444
rect 1204 -332 1210 444
rect 1034 -344 1210 -332
rect 1622 444 1798 456
rect 1622 -332 1628 444
rect 1662 -332 1758 444
rect 1792 -332 1798 444
rect 1622 -344 1798 -332
rect 2210 444 2386 456
rect 2210 -332 2216 444
rect 2250 -332 2346 444
rect 2380 -332 2386 444
rect 2210 -344 2386 -332
rect 2798 444 2974 456
rect 2798 -332 2804 444
rect 2838 -332 2934 444
rect 2968 -332 2974 444
rect 2798 -344 2974 -332
rect 3386 444 3562 456
rect 3386 -332 3392 444
rect 3426 -332 3522 444
rect 3556 -332 3562 444
rect 3386 -344 3562 -332
rect 3974 444 4150 456
rect 3974 -332 3980 444
rect 4014 -332 4110 444
rect 4144 -332 4150 444
rect 3974 -344 4150 -332
rect 4562 444 4738 456
rect 4562 -332 4568 444
rect 4602 -332 4698 444
rect 4732 -332 4738 444
rect 4562 -344 4738 -332
rect 5150 444 5248 456
rect 5150 -332 5156 444
rect 5190 -332 5248 444
rect 5150 -344 5248 -332
rect 5280 444 5326 456
rect 5280 -332 5286 444
rect 5320 -332 5326 444
rect 5280 -344 5326 -332
rect 5738 444 5914 456
rect 5738 -332 5744 444
rect 5778 -332 5874 444
rect 5908 -332 5914 444
rect 5738 -344 5914 -332
rect 6326 444 6502 456
rect 6326 -332 6332 444
rect 6366 -332 6462 444
rect 6496 -332 6502 444
rect 6326 -344 6502 -332
rect 6914 444 7090 456
rect 6914 -332 6920 444
rect 6954 -332 7050 444
rect 7084 -332 7090 444
rect 6914 -344 7090 -332
rect 7502 444 7548 456
rect 7502 -332 7508 444
rect 7542 -332 7548 444
rect 7502 -344 7548 -332
rect 7632 444 7678 456
rect 7632 -332 7638 444
rect 7672 -332 7678 444
rect 7632 -344 7678 -332
rect 8090 444 8266 456
rect 8090 -332 8096 444
rect 8130 -332 8226 444
rect 8260 -332 8266 444
rect 8090 -344 8266 -332
rect 8678 444 8854 456
rect 8678 -332 8684 444
rect 8718 -332 8814 444
rect 8848 -332 8854 444
rect 8678 -344 8854 -332
rect 9266 444 9442 456
rect 9266 -332 9272 444
rect 9306 -332 9402 444
rect 9436 -332 9442 444
rect 9266 -344 9442 -332
rect 9854 444 9900 456
rect 9854 -332 9860 444
rect 9894 -332 9900 444
rect 9854 -344 9900 -332
rect 9934 444 10030 456
rect 9934 -332 9990 444
rect 10024 -332 10030 444
rect 9934 -344 10030 -332
rect 10442 444 10618 456
rect 10442 -332 10448 444
rect 10482 -332 10578 444
rect 10612 -332 10618 444
rect 10442 -344 10618 -332
rect 11030 444 11206 456
rect 11030 -332 11036 444
rect 11070 -332 11166 444
rect 11200 -332 11206 444
rect 11030 -344 11206 -332
rect 11618 444 11794 456
rect 11618 -332 11624 444
rect 11658 -332 11754 444
rect 11788 -332 11794 444
rect 11618 -344 11794 -332
rect 12206 444 12382 456
rect 12206 -332 12212 444
rect 12246 -332 12342 444
rect 12376 -332 12382 444
rect 12206 -344 12382 -332
rect 12794 444 12970 456
rect 12794 -332 12800 444
rect 12834 -332 12930 444
rect 12964 -332 12970 444
rect 12794 -344 12970 -332
rect 13382 444 13558 456
rect 13382 -332 13388 444
rect 13422 -332 13518 444
rect 13552 -332 13558 444
rect 13382 -344 13558 -332
rect 13970 444 14146 456
rect 13970 -332 13976 444
rect 14010 -332 14106 444
rect 14140 -332 14146 444
rect 13970 -344 14146 -332
rect 14558 444 14734 456
rect 14558 -332 14564 444
rect 14598 -332 14694 444
rect 14728 -332 14734 444
rect 14558 -344 14734 -332
rect 15146 444 15322 456
rect 15146 -332 15152 444
rect 15186 -332 15282 444
rect 15316 -332 15322 444
rect 15146 -344 15322 -332
rect 15734 444 15910 456
rect 15734 -332 15740 444
rect 15774 -332 15870 444
rect 15904 -332 15910 444
rect 15734 -344 15910 -332
rect 16322 444 16498 456
rect 16322 -332 16328 444
rect 16362 -332 16458 444
rect 16492 -332 16498 444
rect 16322 -344 16498 -332
rect 16910 444 17086 456
rect 16910 -332 16916 444
rect 16950 -332 17046 444
rect 17080 -332 17086 444
rect 16910 -344 17086 -332
rect 17498 444 17674 456
rect 17498 -332 17504 444
rect 17538 -332 17634 444
rect 17668 -332 17674 444
rect 17498 -344 17674 -332
rect 18086 444 18262 456
rect 18086 -332 18092 444
rect 18126 -332 18222 444
rect 18256 -332 18262 444
rect 18086 -344 18262 -332
rect 18674 444 18850 456
rect 18674 -332 18680 444
rect 18714 -332 18810 444
rect 18844 -332 18850 444
rect 18674 -344 18850 -332
rect 19262 444 19438 456
rect 19262 -332 19268 444
rect 19302 -332 19398 444
rect 19432 -332 19438 444
rect 19262 -344 19438 -332
rect 19850 444 20026 456
rect 19850 -332 19856 444
rect 19890 -332 19986 444
rect 20020 -332 20026 444
rect 19850 -344 20026 -332
rect 20438 444 20614 456
rect 20438 -332 20444 444
rect 20478 -332 20574 444
rect 20608 -332 20614 444
rect 20438 -344 20614 -332
rect 21026 444 21202 456
rect 21026 -332 21032 444
rect 21066 -332 21162 444
rect 21196 -332 21202 444
rect 21026 -344 21202 -332
rect 21614 444 21744 456
rect 21614 -332 21620 444
rect 21654 -332 21744 444
rect 21614 -344 21744 -332
rect -6424 -391 -6032 -385
rect -6424 -425 -6412 -391
rect -6044 -425 -6032 -391
rect -6424 -431 -6032 -425
rect -5970 -688 -5898 -344
rect -5836 -391 -5444 -385
rect -5836 -425 -5824 -391
rect -5456 -425 -5444 -391
rect -5836 -431 -5444 -425
rect -5248 -391 -4856 -385
rect -5248 -425 -5236 -391
rect -4868 -425 -4856 -391
rect -5248 -431 -4856 -425
rect -4794 -688 -4722 -344
rect -4660 -391 -4268 -385
rect -4660 -425 -4648 -391
rect -4280 -425 -4268 -391
rect -4660 -431 -4268 -425
rect -4072 -391 -3680 -385
rect -4072 -425 -4060 -391
rect -3692 -425 -3680 -391
rect -4072 -431 -3680 -425
rect -3618 -688 -3546 -344
rect -3484 -391 -3092 -385
rect -3484 -425 -3472 -391
rect -3104 -425 -3092 -391
rect -3484 -431 -3092 -425
rect -2896 -391 -2504 -385
rect -2896 -425 -2884 -391
rect -2516 -425 -2504 -391
rect -2896 -431 -2504 -425
rect -2442 -688 -2370 -344
rect -2308 -391 -1916 -385
rect -2308 -425 -2296 -391
rect -1928 -425 -1916 -391
rect -2308 -431 -1916 -425
rect -1720 -391 -1328 -385
rect -1720 -425 -1708 -391
rect -1340 -425 -1328 -391
rect -1720 -431 -1328 -425
rect -1266 -688 -1194 -344
rect -1132 -391 -740 -385
rect -1132 -425 -1120 -391
rect -752 -425 -740 -391
rect -1132 -431 -740 -425
rect -544 -391 -152 -385
rect -544 -425 -532 -391
rect -164 -425 -152 -391
rect -544 -431 -152 -425
rect -90 -688 -18 -344
rect 44 -391 436 -385
rect 44 -425 56 -391
rect 424 -425 436 -391
rect 44 -431 436 -425
rect 632 -391 1024 -385
rect 632 -425 644 -391
rect 1012 -425 1024 -391
rect 632 -431 1024 -425
rect 1086 -688 1158 -344
rect 1220 -391 1612 -385
rect 1220 -425 1232 -391
rect 1600 -425 1612 -391
rect 1220 -431 1612 -425
rect 1808 -391 2200 -385
rect 1808 -425 1820 -391
rect 2188 -425 2200 -391
rect 1808 -431 2200 -425
rect 2262 -688 2334 -344
rect 2396 -391 2788 -385
rect 2396 -425 2408 -391
rect 2776 -425 2788 -391
rect 2396 -431 2788 -425
rect 2984 -391 3376 -385
rect 2984 -425 2996 -391
rect 3364 -425 3376 -391
rect 2984 -431 3376 -425
rect 3438 -688 3510 -344
rect 3572 -391 3964 -385
rect 3572 -425 3584 -391
rect 3952 -425 3964 -391
rect 3572 -431 3964 -425
rect 4160 -391 4552 -385
rect 4160 -425 4172 -391
rect 4540 -425 4552 -391
rect 4160 -431 4552 -425
rect 4614 -688 4686 -344
rect 4748 -391 5140 -385
rect 4748 -425 4760 -391
rect 5128 -425 5140 -391
rect 4748 -431 5140 -425
rect 5336 -391 5728 -385
rect 5336 -425 5348 -391
rect 5716 -425 5728 -391
rect 5336 -431 5728 -425
rect 5790 -688 5862 -344
rect 5924 -391 6316 -385
rect 5924 -425 5936 -391
rect 6304 -425 6316 -391
rect 5924 -431 6316 -425
rect -6040 -694 -5828 -688
rect -6040 -804 -6028 -694
rect -5840 -804 -5828 -694
rect -6040 -810 -5828 -804
rect -4864 -694 -4652 -688
rect -4864 -804 -4852 -694
rect -4664 -804 -4652 -694
rect -4864 -810 -4652 -804
rect -3688 -694 -3476 -688
rect -3688 -804 -3676 -694
rect -3488 -804 -3476 -694
rect -3688 -810 -3476 -804
rect -2512 -694 -2300 -688
rect -2512 -804 -2500 -694
rect -2312 -804 -2300 -694
rect -2512 -810 -2300 -804
rect -1336 -694 -1124 -688
rect -1336 -804 -1324 -694
rect -1136 -804 -1124 -694
rect -1336 -810 -1124 -804
rect -160 -694 52 -688
rect -160 -804 -148 -694
rect 40 -804 52 -694
rect -160 -810 52 -804
rect 1016 -694 1228 -688
rect 1016 -804 1028 -694
rect 1216 -804 1228 -694
rect 1016 -810 1228 -804
rect 2192 -694 2404 -688
rect 2192 -804 2204 -694
rect 2392 -804 2404 -694
rect 2192 -810 2404 -804
rect 3368 -694 3580 -688
rect 3368 -804 3380 -694
rect 3568 -804 3580 -694
rect 3368 -810 3580 -804
rect 4544 -694 4756 -688
rect 4544 -804 4556 -694
rect 4744 -804 4756 -694
rect 4544 -810 4756 -804
rect 5720 -694 5932 -688
rect 5720 -804 5732 -694
rect 5920 -804 5932 -694
rect 5720 -810 5932 -804
rect 6378 -1196 6450 -344
rect 6512 -391 6904 -385
rect 6512 -425 6524 -391
rect 6892 -425 6904 -391
rect 6512 -431 6904 -425
rect 6966 -688 7038 -344
rect 7100 -391 7492 -385
rect 7100 -425 7112 -391
rect 7480 -425 7492 -391
rect 7100 -431 7492 -425
rect 7688 -391 8080 -385
rect 7688 -425 7700 -391
rect 8068 -425 8080 -391
rect 7688 -431 8080 -425
rect 8142 -688 8214 -344
rect 8276 -391 8668 -385
rect 8276 -425 8288 -391
rect 8656 -425 8668 -391
rect 8276 -431 8668 -425
rect 6896 -694 7108 -688
rect 6896 -804 6908 -694
rect 7096 -804 7108 -694
rect 6896 -810 7108 -804
rect 8072 -694 8284 -688
rect 8072 -804 8084 -694
rect 8272 -804 8284 -694
rect 8072 -810 8284 -804
rect 8730 -1196 8802 -344
rect 8864 -391 9256 -385
rect 8864 -425 8876 -391
rect 9244 -425 9256 -391
rect 8864 -431 9256 -425
rect 9318 -688 9390 -344
rect 9452 -391 9844 -385
rect 9452 -425 9464 -391
rect 9832 -425 9844 -391
rect 9452 -431 9844 -425
rect 10040 -391 10432 -385
rect 10040 -425 10052 -391
rect 10420 -425 10432 -391
rect 10040 -431 10432 -425
rect 10494 -688 10566 -344
rect 10628 -391 11020 -385
rect 10628 -425 10640 -391
rect 11008 -425 11020 -391
rect 10628 -431 11020 -425
rect 11216 -391 11608 -385
rect 11216 -425 11228 -391
rect 11596 -425 11608 -391
rect 11216 -431 11608 -425
rect 11670 -688 11742 -344
rect 11804 -391 12196 -385
rect 11804 -425 11816 -391
rect 12184 -425 12196 -391
rect 11804 -431 12196 -425
rect 12392 -391 12784 -385
rect 12392 -425 12404 -391
rect 12772 -425 12784 -391
rect 12392 -431 12784 -425
rect 12846 -678 12918 -344
rect 12980 -391 13372 -385
rect 12980 -425 12992 -391
rect 13360 -425 13372 -391
rect 12980 -431 13372 -425
rect 13568 -391 13960 -385
rect 13568 -425 13580 -391
rect 13948 -425 13960 -391
rect 13568 -431 13960 -425
rect 12776 -684 12988 -678
rect 9248 -694 9460 -688
rect 9248 -804 9260 -694
rect 9448 -804 9460 -694
rect 9248 -810 9460 -804
rect 10424 -694 10636 -688
rect 10424 -804 10436 -694
rect 10624 -804 10636 -694
rect 10424 -810 10636 -804
rect 11600 -694 11812 -688
rect 11600 -804 11612 -694
rect 11800 -804 11812 -694
rect 12776 -794 12788 -684
rect 12976 -794 12988 -684
rect 14022 -688 14094 -344
rect 14156 -391 14548 -385
rect 14156 -425 14168 -391
rect 14536 -425 14548 -391
rect 14156 -431 14548 -425
rect 14744 -391 15136 -385
rect 14744 -425 14756 -391
rect 15124 -425 15136 -391
rect 14744 -431 15136 -425
rect 15198 -688 15270 -344
rect 15332 -391 15724 -385
rect 15332 -425 15344 -391
rect 15712 -425 15724 -391
rect 15332 -431 15724 -425
rect 15920 -391 16312 -385
rect 15920 -425 15932 -391
rect 16300 -425 16312 -391
rect 15920 -431 16312 -425
rect 16374 -688 16446 -344
rect 16508 -391 16900 -385
rect 16508 -425 16520 -391
rect 16888 -425 16900 -391
rect 16508 -431 16900 -425
rect 17096 -391 17488 -385
rect 17096 -425 17108 -391
rect 17476 -425 17488 -391
rect 17096 -431 17488 -425
rect 17550 -678 17622 -344
rect 17684 -391 18076 -385
rect 17684 -425 17696 -391
rect 18064 -425 18076 -391
rect 17684 -431 18076 -425
rect 18272 -391 18664 -385
rect 18272 -425 18284 -391
rect 18652 -425 18664 -391
rect 18272 -431 18664 -425
rect 17466 -684 17702 -678
rect 12776 -800 12988 -794
rect 13952 -694 14164 -688
rect 11600 -810 11812 -804
rect 13952 -804 13964 -694
rect 14152 -804 14164 -694
rect 13952 -810 14164 -804
rect 15128 -694 15340 -688
rect 15128 -804 15140 -694
rect 15328 -804 15340 -694
rect 15128 -810 15340 -804
rect 16304 -694 16516 -688
rect 16304 -804 16316 -694
rect 16504 -804 16516 -694
rect 16304 -810 16516 -804
rect 17466 -806 17478 -684
rect 17690 -806 17702 -684
rect 18726 -688 18798 -344
rect 18860 -391 19252 -385
rect 18860 -425 18872 -391
rect 19240 -425 19252 -391
rect 18860 -431 19252 -425
rect 19448 -391 19840 -385
rect 19448 -425 19460 -391
rect 19828 -425 19840 -391
rect 19448 -431 19840 -425
rect 19902 -688 19974 -344
rect 20036 -391 20428 -385
rect 20036 -425 20048 -391
rect 20416 -425 20428 -391
rect 20036 -431 20428 -425
rect 20624 -391 21016 -385
rect 20624 -425 20636 -391
rect 21004 -425 21016 -391
rect 20624 -431 21016 -425
rect 21078 -688 21150 -344
rect 21212 -391 21604 -385
rect 21212 -425 21224 -391
rect 21592 -425 21604 -391
rect 21212 -431 21604 -425
rect 17466 -812 17702 -806
rect 18656 -694 18868 -688
rect 18656 -804 18668 -694
rect 18856 -804 18868 -694
rect 18656 -810 18868 -804
rect 19832 -694 20044 -688
rect 19832 -804 19844 -694
rect 20032 -804 20044 -694
rect 19832 -810 20044 -804
rect 21008 -694 21220 -688
rect 21008 -804 21020 -694
rect 21208 -804 21220 -694
rect 21008 -810 21220 -804
rect 6378 -1276 8802 -1196
rect 6486 -1990 6566 -1276
rect 6622 -1820 6696 -1814
rect 6622 -1952 6632 -1820
rect 6686 -1952 6696 -1820
rect 6622 -1958 6696 -1952
rect 6888 -1820 6962 -1814
rect 6888 -1952 6898 -1820
rect 6952 -1952 6962 -1820
rect 6888 -1958 6962 -1952
rect 7018 -1990 7098 -1276
rect 7154 -1820 7228 -1814
rect 7154 -1952 7164 -1820
rect 7218 -1952 7228 -1820
rect 7154 -1958 7228 -1952
rect 7420 -1820 7494 -1814
rect 7420 -1952 7430 -1820
rect 7484 -1952 7494 -1820
rect 7420 -1958 7494 -1952
rect 7550 -1990 7630 -1276
rect 7686 -1820 7760 -1814
rect 7686 -1952 7696 -1820
rect 7750 -1952 7760 -1820
rect 7686 -1958 7760 -1952
rect 7952 -1820 8026 -1814
rect 7952 -1952 7962 -1820
rect 8016 -1952 8026 -1820
rect 7952 -1958 8026 -1952
rect 8082 -1990 8162 -1276
rect 8218 -1820 8292 -1814
rect 8218 -1952 8228 -1820
rect 8282 -1952 8292 -1820
rect 8218 -1958 8292 -1952
rect 8484 -1820 8558 -1814
rect 8484 -1952 8494 -1820
rect 8548 -1952 8558 -1820
rect 8484 -1958 8558 -1952
rect 8614 -1990 8694 -1276
rect 6486 -2002 6618 -1990
rect 6486 -2778 6578 -2002
rect 6612 -2778 6618 -2002
rect 6486 -2790 6618 -2778
rect 6700 -2002 6884 -1990
rect 6700 -2778 6706 -2002
rect 6740 -2778 6844 -2002
rect 6878 -2778 6884 -2002
rect 6700 -2790 6884 -2778
rect 6966 -2002 7150 -1990
rect 6966 -2778 6972 -2002
rect 7006 -2778 7110 -2002
rect 7144 -2778 7150 -2002
rect 6966 -2790 7150 -2778
rect 7232 -2002 7416 -1990
rect 7232 -2778 7238 -2002
rect 7272 -2778 7376 -2002
rect 7410 -2778 7416 -2002
rect 7232 -2790 7416 -2778
rect 7498 -2002 7682 -1990
rect 7498 -2778 7504 -2002
rect 7538 -2778 7642 -2002
rect 7676 -2778 7682 -2002
rect 7498 -2790 7682 -2778
rect 7764 -2002 7948 -1990
rect 7764 -2778 7770 -2002
rect 7804 -2778 7908 -2002
rect 7942 -2778 7948 -2002
rect 7764 -2790 7948 -2778
rect 8030 -2002 8214 -1990
rect 8030 -2778 8036 -2002
rect 8070 -2778 8174 -2002
rect 8208 -2778 8214 -2002
rect 8030 -2790 8214 -2778
rect 8296 -2002 8480 -1990
rect 8296 -2778 8302 -2002
rect 8336 -2778 8440 -2002
rect 8474 -2778 8480 -2002
rect 8296 -2790 8480 -2778
rect 8562 -2002 8694 -1990
rect 8562 -2778 8568 -2002
rect 8602 -2778 8694 -2002
rect 8562 -2790 8694 -2778
rect 6486 -3000 6572 -2790
rect 6622 -2830 6696 -2824
rect 6622 -2962 6632 -2830
rect 6686 -2962 6696 -2830
rect 6622 -2968 6696 -2962
rect 6746 -3000 6838 -2790
rect 6888 -2830 6962 -2824
rect 6888 -2962 6898 -2830
rect 6952 -2962 6962 -2830
rect 6888 -2968 6962 -2962
rect 7012 -3000 7104 -2790
rect 7154 -2830 7228 -2824
rect 7154 -2962 7164 -2830
rect 7218 -2962 7228 -2830
rect 7154 -2968 7228 -2962
rect 7278 -3000 7370 -2790
rect 7420 -2830 7494 -2824
rect 7420 -2962 7430 -2830
rect 7484 -2962 7494 -2830
rect 7420 -2968 7494 -2962
rect 7544 -3000 7636 -2790
rect 7686 -2830 7760 -2824
rect 7686 -2962 7696 -2830
rect 7750 -2962 7760 -2830
rect 7686 -2968 7760 -2962
rect 7810 -3000 7902 -2790
rect 7952 -2830 8026 -2824
rect 7952 -2962 7962 -2830
rect 8016 -2962 8026 -2830
rect 7952 -2968 8026 -2962
rect 8076 -3000 8168 -2790
rect 8218 -2830 8292 -2824
rect 8218 -2962 8228 -2830
rect 8282 -2962 8292 -2830
rect 8218 -2968 8292 -2962
rect 8342 -3000 8434 -2790
rect 8484 -2830 8558 -2824
rect 8484 -2962 8494 -2830
rect 8548 -2962 8558 -2830
rect 8484 -2968 8558 -2962
rect 8608 -3000 8694 -2790
rect 6486 -3012 6618 -3000
rect 6486 -3788 6578 -3012
rect 6612 -3788 6618 -3012
rect 6486 -3800 6618 -3788
rect 6700 -3012 6884 -3000
rect 6700 -3788 6706 -3012
rect 6740 -3788 6844 -3012
rect 6878 -3788 6884 -3012
rect 6700 -3800 6884 -3788
rect 6966 -3012 7150 -3000
rect 6966 -3788 6972 -3012
rect 7006 -3788 7110 -3012
rect 7144 -3788 7150 -3012
rect 6966 -3800 7150 -3788
rect 7232 -3012 7416 -3000
rect 7232 -3788 7238 -3012
rect 7272 -3788 7376 -3012
rect 7410 -3788 7416 -3012
rect 7232 -3800 7416 -3788
rect 7498 -3012 7682 -3000
rect 7498 -3788 7504 -3012
rect 7538 -3788 7642 -3012
rect 7676 -3788 7682 -3012
rect 7498 -3800 7682 -3788
rect 7764 -3012 7948 -3000
rect 7764 -3788 7770 -3012
rect 7804 -3788 7908 -3012
rect 7942 -3788 7948 -3012
rect 7764 -3800 7948 -3788
rect 8030 -3012 8214 -3000
rect 8030 -3788 8036 -3012
rect 8070 -3788 8174 -3012
rect 8208 -3788 8214 -3012
rect 8030 -3800 8214 -3788
rect 8296 -3012 8480 -3000
rect 8296 -3788 8302 -3012
rect 8336 -3788 8440 -3012
rect 8474 -3788 8480 -3012
rect 8296 -3800 8480 -3788
rect 8562 -3012 8694 -3000
rect 8562 -3788 8568 -3012
rect 8602 -3788 8694 -3012
rect 8562 -3800 8694 -3788
rect 6486 -4010 6572 -3800
rect 6622 -3840 6696 -3834
rect 6622 -3972 6632 -3840
rect 6686 -3972 6696 -3840
rect 6622 -3978 6696 -3972
rect 6746 -4010 6838 -3800
rect 6888 -3840 6962 -3834
rect 6888 -3972 6898 -3840
rect 6952 -3972 6962 -3840
rect 6888 -3978 6962 -3972
rect 7012 -4010 7104 -3800
rect 7154 -3840 7228 -3834
rect 7154 -3972 7164 -3840
rect 7218 -3972 7228 -3840
rect 7154 -3978 7228 -3972
rect 7278 -4010 7370 -3800
rect 7420 -3840 7494 -3834
rect 7420 -3972 7430 -3840
rect 7484 -3972 7494 -3840
rect 7420 -3978 7494 -3972
rect 7544 -4010 7636 -3800
rect 7686 -3840 7760 -3834
rect 7686 -3972 7696 -3840
rect 7750 -3972 7760 -3840
rect 7686 -3978 7760 -3972
rect 7810 -4010 7902 -3800
rect 7952 -3840 8026 -3834
rect 7952 -3972 7962 -3840
rect 8016 -3972 8026 -3840
rect 7952 -3978 8026 -3972
rect 8076 -4010 8168 -3800
rect 8218 -3840 8292 -3834
rect 8218 -3972 8228 -3840
rect 8282 -3972 8292 -3840
rect 8218 -3978 8292 -3972
rect 8342 -4010 8434 -3800
rect 8484 -3840 8558 -3834
rect 8484 -3972 8494 -3840
rect 8548 -3972 8558 -3840
rect 8484 -3978 8558 -3972
rect 8608 -4010 8694 -3800
rect 13532 -3854 13542 -3316
rect 14024 -3854 14034 -3316
rect 13753 -3912 13759 -3854
rect 13797 -3912 13803 -3854
rect 13753 -3924 13803 -3912
rect 6486 -4022 6618 -4010
rect 6486 -4798 6578 -4022
rect 6612 -4798 6618 -4022
rect 6486 -4810 6618 -4798
rect 6700 -4022 6884 -4010
rect 6700 -4798 6706 -4022
rect 6740 -4798 6844 -4022
rect 6878 -4798 6884 -4022
rect 6700 -4810 6884 -4798
rect 6966 -4022 7150 -4010
rect 6966 -4798 6972 -4022
rect 7006 -4798 7110 -4022
rect 7144 -4798 7150 -4022
rect 6966 -4810 7150 -4798
rect 7232 -4022 7416 -4010
rect 7232 -4798 7238 -4022
rect 7272 -4798 7376 -4022
rect 7410 -4798 7416 -4022
rect 7232 -4810 7416 -4798
rect 7498 -4022 7682 -4010
rect 7498 -4798 7504 -4022
rect 7538 -4798 7642 -4022
rect 7676 -4798 7682 -4022
rect 7498 -4810 7682 -4798
rect 7764 -4022 7948 -4010
rect 7764 -4798 7770 -4022
rect 7804 -4798 7908 -4022
rect 7942 -4798 7948 -4022
rect 7764 -4810 7948 -4798
rect 8030 -4022 8214 -4010
rect 8030 -4798 8036 -4022
rect 8070 -4798 8174 -4022
rect 8208 -4798 8214 -4022
rect 8030 -4810 8214 -4798
rect 8296 -4022 8480 -4010
rect 8296 -4798 8302 -4022
rect 8336 -4798 8440 -4022
rect 8474 -4798 8480 -4022
rect 8296 -4810 8480 -4798
rect 8562 -4022 8694 -4010
rect 8562 -4798 8568 -4022
rect 8602 -4798 8694 -4022
rect 14032 -4122 14206 -4102
rect 8562 -4810 8694 -4798
rect 13753 -4506 13803 -4494
rect 6622 -4850 6696 -4844
rect 6622 -4982 6632 -4850
rect 6686 -4982 6696 -4850
rect 6622 -4988 6696 -4982
rect 6752 -6182 6832 -4810
rect 6888 -4850 6962 -4844
rect 6888 -4982 6898 -4850
rect 6952 -4982 6962 -4850
rect 6888 -4988 6962 -4982
rect 7154 -4850 7228 -4844
rect 7154 -4982 7164 -4850
rect 7218 -4982 7228 -4850
rect 7154 -4988 7228 -4982
rect 7284 -5366 7364 -4810
rect 7420 -4850 7494 -4844
rect 7420 -4982 7430 -4850
rect 7484 -4982 7494 -4850
rect 7420 -4988 7494 -4982
rect 7686 -4850 7760 -4844
rect 7686 -4982 7696 -4850
rect 7750 -4982 7760 -4850
rect 7686 -4988 7760 -4982
rect 7816 -5366 7896 -4810
rect 7952 -4850 8026 -4844
rect 7952 -4982 7962 -4850
rect 8016 -4982 8026 -4850
rect 7952 -4988 8026 -4982
rect 8218 -4850 8292 -4844
rect 8218 -4982 8228 -4850
rect 8282 -4982 8292 -4850
rect 8218 -4988 8292 -4982
rect 7284 -5398 7896 -5366
rect 7284 -5526 7330 -5398
rect 7824 -5526 7896 -5398
rect 7284 -5556 7896 -5526
rect 7196 -6018 7506 -6012
rect 7196 -6144 7212 -6018
rect 7250 -6144 7452 -6018
rect 7490 -6144 7506 -6018
rect 7196 -6150 7266 -6144
rect 7436 -6150 7506 -6144
rect 7564 -6182 7618 -5556
rect 7676 -6018 7986 -6012
rect 7676 -6144 7692 -6018
rect 7730 -6144 7932 -6018
rect 7970 -6144 7986 -6018
rect 7676 -6150 7746 -6144
rect 7916 -6150 7986 -6144
rect 8348 -6182 8428 -4810
rect 8484 -4850 8558 -4844
rect 8484 -4982 8494 -4850
rect 8548 -4982 8558 -4850
rect 13753 -4890 13759 -4506
rect 8484 -4988 8558 -4982
rect 13742 -4903 13759 -4890
rect 13797 -4890 13803 -4506
rect 14032 -4582 14048 -4122
rect 14188 -4582 14206 -4122
rect 13797 -4903 13814 -4890
rect 13742 -5332 13814 -4903
rect 13618 -5698 13628 -5332
rect 13910 -5698 13920 -5332
rect 6752 -6194 7190 -6182
rect 6752 -6252 7150 -6194
rect 7100 -6770 7150 -6252
rect 7184 -6770 7190 -6194
rect 7100 -6782 7190 -6770
rect 7272 -6194 7430 -6182
rect 7272 -6770 7278 -6194
rect 7312 -6770 7390 -6194
rect 7424 -6770 7430 -6194
rect 7272 -6782 7430 -6770
rect 7512 -6194 7670 -6182
rect 7512 -6770 7518 -6194
rect 7552 -6770 7630 -6194
rect 7664 -6770 7670 -6194
rect 7512 -6782 7670 -6770
rect 7752 -6194 7910 -6182
rect 7752 -6770 7758 -6194
rect 7792 -6770 7870 -6194
rect 7904 -6770 7910 -6194
rect 7752 -6782 7910 -6770
rect 7992 -6194 8428 -6182
rect 7992 -6770 7998 -6194
rect 8032 -6252 8428 -6194
rect 8032 -6770 8088 -6252
rect 7992 -6782 8088 -6770
rect 7100 -6990 7150 -6782
rect 7196 -6820 7266 -6814
rect 7196 -6952 7212 -6820
rect 7250 -6952 7266 -6820
rect 7196 -6958 7266 -6952
rect 7318 -6990 7384 -6782
rect 7436 -6820 7506 -6814
rect 7436 -6952 7452 -6820
rect 7490 -6952 7506 -6820
rect 7436 -6958 7506 -6952
rect 7558 -6990 7624 -6782
rect 7676 -6820 7746 -6814
rect 7676 -6952 7692 -6820
rect 7730 -6952 7746 -6820
rect 7676 -6958 7746 -6952
rect 7798 -6990 7864 -6782
rect 7916 -6820 7986 -6814
rect 7916 -6952 7932 -6820
rect 7970 -6952 7986 -6820
rect 7916 -6958 7986 -6952
rect 8038 -6990 8088 -6782
rect 7100 -7002 7190 -6990
rect 7100 -7578 7150 -7002
rect 7184 -7578 7190 -7002
rect 7100 -7590 7190 -7578
rect 7272 -7002 7430 -6990
rect 7272 -7578 7278 -7002
rect 7312 -7578 7390 -7002
rect 7424 -7578 7430 -7002
rect 7272 -7590 7430 -7578
rect 7512 -7002 7670 -6990
rect 7512 -7578 7518 -7002
rect 7552 -7578 7630 -7002
rect 7664 -7578 7670 -7002
rect 7512 -7590 7670 -7578
rect 7752 -7002 7910 -6990
rect 7752 -7578 7758 -7002
rect 7792 -7578 7870 -7002
rect 7904 -7578 7910 -7002
rect 7752 -7590 7910 -7578
rect 7992 -7002 8088 -6990
rect 7992 -7578 7998 -7002
rect 8032 -7578 8088 -7002
rect 14032 -7432 14206 -4582
rect 7992 -7590 8088 -7578
rect 7196 -7628 7266 -7622
rect 7196 -7760 7212 -7628
rect 7250 -7760 7266 -7628
rect 7196 -7766 7266 -7760
rect 7324 -8006 7378 -7590
rect 7436 -7628 7506 -7622
rect 7436 -7760 7452 -7628
rect 7490 -7760 7506 -7628
rect 7436 -7766 7506 -7760
rect 7676 -7628 7746 -7622
rect 7676 -7760 7692 -7628
rect 7730 -7760 7746 -7628
rect 7676 -7766 7746 -7760
rect 7804 -8006 7858 -7590
rect 7916 -7628 7986 -7622
rect 7916 -7760 7932 -7628
rect 7970 -7760 7986 -7628
rect 7916 -7766 7986 -7760
rect 6890 -8012 8266 -8006
rect 6890 -8124 6902 -8012
rect 8254 -8124 8266 -8012
rect 13744 -8098 13754 -7432
rect 14510 -8098 14520 -7432
rect 6890 -8130 8266 -8124
<< via1 >>
rect 2976 7018 3086 7090
rect 3456 7018 3566 7090
rect 3936 7018 4046 7090
rect 4416 7018 4526 7090
rect 4896 7018 5006 7090
rect 5376 7018 5486 7090
rect 5856 7018 5966 7090
rect 6336 7018 6446 7090
rect 6816 7018 6926 7090
rect 7296 7018 7406 7090
rect 7776 7018 7886 7090
rect 8256 7018 8366 7090
rect 8736 7018 8846 7090
rect 9216 7018 9326 7090
rect 9696 7018 9806 7090
rect 10176 7018 10286 7090
rect 10656 7018 10766 7090
rect 11136 7018 11246 7090
rect 11616 7018 11726 7090
rect 12096 7018 12206 7090
rect 2876 6614 2892 6746
rect 2892 6614 2930 6746
rect 2930 6614 2946 6746
rect 3116 6614 3132 6746
rect 3132 6614 3170 6746
rect 3170 6614 3186 6746
rect 3356 6614 3372 6746
rect 3372 6614 3410 6746
rect 3410 6614 3426 6746
rect 3596 6614 3612 6746
rect 3612 6614 3650 6746
rect 3650 6614 3666 6746
rect 3836 6614 3852 6746
rect 3852 6614 3890 6746
rect 3890 6614 3906 6746
rect 4076 6614 4092 6746
rect 4092 6614 4130 6746
rect 4130 6614 4146 6746
rect 4316 6614 4332 6746
rect 4332 6614 4370 6746
rect 4370 6614 4386 6746
rect 4556 6614 4572 6746
rect 4572 6614 4610 6746
rect 4610 6614 4626 6746
rect 4796 6614 4812 6746
rect 4812 6614 4850 6746
rect 4850 6614 4866 6746
rect 5036 6614 5052 6746
rect 5052 6614 5090 6746
rect 5090 6614 5106 6746
rect 5276 6614 5292 6746
rect 5292 6614 5330 6746
rect 5330 6614 5346 6746
rect 5516 6614 5532 6746
rect 5532 6614 5570 6746
rect 5570 6614 5586 6746
rect 5756 6614 5772 6746
rect 5772 6614 5810 6746
rect 5810 6614 5826 6746
rect 5996 6614 6012 6746
rect 6012 6614 6050 6746
rect 6050 6614 6066 6746
rect 6236 6614 6252 6746
rect 6252 6614 6290 6746
rect 6290 6614 6306 6746
rect 6476 6614 6492 6746
rect 6492 6614 6530 6746
rect 6530 6614 6546 6746
rect 6716 6614 6732 6746
rect 6732 6614 6770 6746
rect 6770 6614 6786 6746
rect 6956 6614 6972 6746
rect 6972 6614 7010 6746
rect 7010 6614 7026 6746
rect 7196 6614 7212 6746
rect 7212 6614 7250 6746
rect 7250 6614 7266 6746
rect 7436 6614 7452 6746
rect 7452 6614 7490 6746
rect 7490 6614 7506 6746
rect 7676 6614 7692 6746
rect 7692 6614 7730 6746
rect 7730 6614 7746 6746
rect 7916 6614 7932 6746
rect 7932 6614 7970 6746
rect 7970 6614 7986 6746
rect 8156 6614 8172 6746
rect 8172 6614 8210 6746
rect 8210 6614 8226 6746
rect 8396 6614 8412 6746
rect 8412 6614 8450 6746
rect 8450 6614 8466 6746
rect 8636 6614 8652 6746
rect 8652 6614 8690 6746
rect 8690 6614 8706 6746
rect 8876 6614 8892 6746
rect 8892 6614 8930 6746
rect 8930 6614 8946 6746
rect 9116 6614 9132 6746
rect 9132 6614 9170 6746
rect 9170 6614 9186 6746
rect 9356 6614 9372 6746
rect 9372 6614 9410 6746
rect 9410 6614 9426 6746
rect 9596 6614 9612 6746
rect 9612 6614 9650 6746
rect 9650 6614 9666 6746
rect 9836 6614 9852 6746
rect 9852 6614 9890 6746
rect 9890 6614 9906 6746
rect 10076 6614 10092 6746
rect 10092 6614 10130 6746
rect 10130 6614 10146 6746
rect 10316 6614 10332 6746
rect 10332 6614 10370 6746
rect 10370 6614 10386 6746
rect 10556 6614 10572 6746
rect 10572 6614 10610 6746
rect 10610 6614 10626 6746
rect 10796 6614 10812 6746
rect 10812 6614 10850 6746
rect 10850 6614 10866 6746
rect 11036 6614 11052 6746
rect 11052 6614 11090 6746
rect 11090 6614 11106 6746
rect 11276 6614 11292 6746
rect 11292 6614 11330 6746
rect 11330 6614 11346 6746
rect 11516 6614 11532 6746
rect 11532 6614 11570 6746
rect 11570 6614 11586 6746
rect 11756 6614 11772 6746
rect 11772 6614 11810 6746
rect 11810 6614 11826 6746
rect 11996 6614 12012 6746
rect 12012 6614 12050 6746
rect 12050 6614 12066 6746
rect 12236 6614 12252 6746
rect 12252 6614 12290 6746
rect 12290 6614 12306 6746
rect 2876 5806 2892 5938
rect 2892 5806 2930 5938
rect 2930 5806 2946 5938
rect 3116 5806 3132 5938
rect 3132 5806 3170 5938
rect 3170 5806 3186 5938
rect 3356 5806 3372 5938
rect 3372 5806 3410 5938
rect 3410 5806 3426 5938
rect 3596 5806 3612 5938
rect 3612 5806 3650 5938
rect 3650 5806 3666 5938
rect 3836 5806 3852 5938
rect 3852 5806 3890 5938
rect 3890 5806 3906 5938
rect 4076 5806 4092 5938
rect 4092 5806 4130 5938
rect 4130 5806 4146 5938
rect 4316 5806 4332 5938
rect 4332 5806 4370 5938
rect 4370 5806 4386 5938
rect 4556 5806 4572 5938
rect 4572 5806 4610 5938
rect 4610 5806 4626 5938
rect 4796 5806 4812 5938
rect 4812 5806 4850 5938
rect 4850 5806 4866 5938
rect 5036 5806 5052 5938
rect 5052 5806 5090 5938
rect 5090 5806 5106 5938
rect 5276 5806 5292 5938
rect 5292 5806 5330 5938
rect 5330 5806 5346 5938
rect 5516 5806 5532 5938
rect 5532 5806 5570 5938
rect 5570 5806 5586 5938
rect 5756 5806 5772 5938
rect 5772 5806 5810 5938
rect 5810 5806 5826 5938
rect 5996 5806 6012 5938
rect 6012 5806 6050 5938
rect 6050 5806 6066 5938
rect 6236 5806 6252 5938
rect 6252 5806 6290 5938
rect 6290 5806 6306 5938
rect 6476 5806 6492 5938
rect 6492 5806 6530 5938
rect 6530 5806 6546 5938
rect 6716 5806 6732 5938
rect 6732 5806 6770 5938
rect 6770 5806 6786 5938
rect 6956 5806 6972 5938
rect 6972 5806 7010 5938
rect 7010 5806 7026 5938
rect 7196 5806 7212 5938
rect 7212 5806 7250 5938
rect 7250 5806 7266 5938
rect 7436 5806 7452 5938
rect 7452 5806 7490 5938
rect 7490 5806 7506 5938
rect 7676 5806 7692 5938
rect 7692 5806 7730 5938
rect 7730 5806 7746 5938
rect 7916 5806 7932 5938
rect 7932 5806 7970 5938
rect 7970 5806 7986 5938
rect 8156 5806 8172 5938
rect 8172 5806 8210 5938
rect 8210 5806 8226 5938
rect 8396 5806 8412 5938
rect 8412 5806 8450 5938
rect 8450 5806 8466 5938
rect 8636 5806 8652 5938
rect 8652 5806 8690 5938
rect 8690 5806 8706 5938
rect 8876 5806 8892 5938
rect 8892 5806 8930 5938
rect 8930 5806 8946 5938
rect 9116 5806 9132 5938
rect 9132 5806 9170 5938
rect 9170 5806 9186 5938
rect 9356 5806 9372 5938
rect 9372 5806 9410 5938
rect 9410 5806 9426 5938
rect 9596 5806 9612 5938
rect 9612 5806 9650 5938
rect 9650 5806 9666 5938
rect 9836 5806 9852 5938
rect 9852 5806 9890 5938
rect 9890 5806 9906 5938
rect 10076 5806 10092 5938
rect 10092 5806 10130 5938
rect 10130 5806 10146 5938
rect 10316 5806 10332 5938
rect 10332 5806 10370 5938
rect 10370 5806 10386 5938
rect 10556 5806 10572 5938
rect 10572 5806 10610 5938
rect 10610 5806 10626 5938
rect 10796 5806 10812 5938
rect 10812 5806 10850 5938
rect 10850 5806 10866 5938
rect 11036 5806 11052 5938
rect 11052 5806 11090 5938
rect 11090 5806 11106 5938
rect 11276 5806 11292 5938
rect 11292 5806 11330 5938
rect 11330 5806 11346 5938
rect 11516 5806 11532 5938
rect 11532 5806 11570 5938
rect 11570 5806 11586 5938
rect 11756 5806 11772 5938
rect 11772 5806 11810 5938
rect 11810 5806 11826 5938
rect 11996 5806 12012 5938
rect 12012 5806 12050 5938
rect 12050 5806 12066 5938
rect 12236 5806 12252 5938
rect 12252 5806 12290 5938
rect 12290 5806 12306 5938
rect 2876 4998 2892 5130
rect 2892 4998 2930 5130
rect 2930 4998 2946 5130
rect 3116 4998 3132 5130
rect 3132 4998 3170 5130
rect 3170 4998 3186 5130
rect 3356 4998 3372 5130
rect 3372 4998 3410 5130
rect 3410 4998 3426 5130
rect 3596 4998 3612 5130
rect 3612 4998 3650 5130
rect 3650 4998 3666 5130
rect 3836 4998 3852 5130
rect 3852 4998 3890 5130
rect 3890 4998 3906 5130
rect 4076 4998 4092 5130
rect 4092 4998 4130 5130
rect 4130 4998 4146 5130
rect 4316 4998 4332 5130
rect 4332 4998 4370 5130
rect 4370 4998 4386 5130
rect 4556 4998 4572 5130
rect 4572 4998 4610 5130
rect 4610 4998 4626 5130
rect 4796 4998 4812 5130
rect 4812 4998 4850 5130
rect 4850 4998 4866 5130
rect 5036 4998 5052 5130
rect 5052 4998 5090 5130
rect 5090 4998 5106 5130
rect 5276 4998 5292 5130
rect 5292 4998 5330 5130
rect 5330 4998 5346 5130
rect 5516 4998 5532 5130
rect 5532 4998 5570 5130
rect 5570 4998 5586 5130
rect 5756 4998 5772 5130
rect 5772 4998 5810 5130
rect 5810 4998 5826 5130
rect 5996 4998 6012 5130
rect 6012 4998 6050 5130
rect 6050 4998 6066 5130
rect 6236 4998 6252 5130
rect 6252 4998 6290 5130
rect 6290 4998 6306 5130
rect 6476 4998 6492 5130
rect 6492 4998 6530 5130
rect 6530 4998 6546 5130
rect 6716 4998 6732 5130
rect 6732 4998 6770 5130
rect 6770 4998 6786 5130
rect 6956 4998 6972 5130
rect 6972 4998 7010 5130
rect 7010 4998 7026 5130
rect 7196 4998 7212 5130
rect 7212 4998 7250 5130
rect 7250 4998 7266 5130
rect 7436 4998 7452 5130
rect 7452 4998 7490 5130
rect 7490 4998 7506 5130
rect 7676 4998 7692 5130
rect 7692 4998 7730 5130
rect 7730 4998 7746 5130
rect 7916 4998 7932 5130
rect 7932 4998 7970 5130
rect 7970 4998 7986 5130
rect 8156 4998 8172 5130
rect 8172 4998 8210 5130
rect 8210 4998 8226 5130
rect 8396 4998 8412 5130
rect 8412 4998 8450 5130
rect 8450 4998 8466 5130
rect 8636 4998 8652 5130
rect 8652 4998 8690 5130
rect 8690 4998 8706 5130
rect 8876 4998 8892 5130
rect 8892 4998 8930 5130
rect 8930 4998 8946 5130
rect 9116 4998 9132 5130
rect 9132 4998 9170 5130
rect 9170 4998 9186 5130
rect 9356 4998 9372 5130
rect 9372 4998 9410 5130
rect 9410 4998 9426 5130
rect 9596 4998 9612 5130
rect 9612 4998 9650 5130
rect 9650 4998 9666 5130
rect 9836 4998 9852 5130
rect 9852 4998 9890 5130
rect 9890 4998 9906 5130
rect 10076 4998 10092 5130
rect 10092 4998 10130 5130
rect 10130 4998 10146 5130
rect 10316 4998 10332 5130
rect 10332 4998 10370 5130
rect 10370 4998 10386 5130
rect 10556 4998 10572 5130
rect 10572 4998 10610 5130
rect 10610 4998 10626 5130
rect 10796 4998 10812 5130
rect 10812 4998 10850 5130
rect 10850 4998 10866 5130
rect 11036 4998 11052 5130
rect 11052 4998 11090 5130
rect 11090 4998 11106 5130
rect 11276 4998 11292 5130
rect 11292 4998 11330 5130
rect 11330 4998 11346 5130
rect 11516 4998 11532 5130
rect 11532 4998 11570 5130
rect 11570 4998 11586 5130
rect 11756 4998 11772 5130
rect 11772 4998 11810 5130
rect 11810 4998 11826 5130
rect 11996 4998 12012 5130
rect 12012 4998 12050 5130
rect 12050 4998 12066 5130
rect 12236 4998 12252 5130
rect 12252 4998 12290 5130
rect 12290 4998 12306 5130
rect 16818 3560 17718 4104
rect -6028 -804 -5840 -694
rect -4852 -804 -4664 -694
rect -3676 -804 -3488 -694
rect -2500 -804 -2312 -694
rect -1324 -804 -1136 -694
rect -148 -804 40 -694
rect 1028 -804 1216 -694
rect 2204 -804 2392 -694
rect 3380 -804 3568 -694
rect 4556 -804 4744 -694
rect 5732 -804 5920 -694
rect 6908 -804 7096 -694
rect 8084 -804 8272 -694
rect 9260 -804 9448 -694
rect 10436 -804 10624 -694
rect 11612 -804 11800 -694
rect 13964 -804 14152 -694
rect 15140 -804 15328 -694
rect 16316 -804 16504 -694
rect 18668 -804 18856 -694
rect 19844 -804 20032 -694
rect 21020 -804 21208 -694
rect 6632 -1952 6640 -1820
rect 6640 -1952 6678 -1820
rect 6678 -1952 6686 -1820
rect 6898 -1952 6906 -1820
rect 6906 -1952 6944 -1820
rect 6944 -1952 6952 -1820
rect 7164 -1952 7172 -1820
rect 7172 -1952 7210 -1820
rect 7210 -1952 7218 -1820
rect 7430 -1952 7438 -1820
rect 7438 -1952 7476 -1820
rect 7476 -1952 7484 -1820
rect 7696 -1952 7704 -1820
rect 7704 -1952 7742 -1820
rect 7742 -1952 7750 -1820
rect 7962 -1952 7970 -1820
rect 7970 -1952 8008 -1820
rect 8008 -1952 8016 -1820
rect 8228 -1952 8236 -1820
rect 8236 -1952 8274 -1820
rect 8274 -1952 8282 -1820
rect 8494 -1952 8502 -1820
rect 8502 -1952 8540 -1820
rect 8540 -1952 8548 -1820
rect 6632 -2962 6640 -2830
rect 6640 -2962 6678 -2830
rect 6678 -2962 6686 -2830
rect 6898 -2962 6906 -2830
rect 6906 -2962 6944 -2830
rect 6944 -2962 6952 -2830
rect 7164 -2962 7172 -2830
rect 7172 -2962 7210 -2830
rect 7210 -2962 7218 -2830
rect 7430 -2962 7438 -2830
rect 7438 -2962 7476 -2830
rect 7476 -2962 7484 -2830
rect 7696 -2962 7704 -2830
rect 7704 -2962 7742 -2830
rect 7742 -2962 7750 -2830
rect 7962 -2962 7970 -2830
rect 7970 -2962 8008 -2830
rect 8008 -2962 8016 -2830
rect 8228 -2962 8236 -2830
rect 8236 -2962 8274 -2830
rect 8274 -2962 8282 -2830
rect 8494 -2962 8502 -2830
rect 8502 -2962 8540 -2830
rect 8540 -2962 8548 -2830
rect 6632 -3972 6640 -3840
rect 6640 -3972 6678 -3840
rect 6678 -3972 6686 -3840
rect 6898 -3972 6906 -3840
rect 6906 -3972 6944 -3840
rect 6944 -3972 6952 -3840
rect 7164 -3972 7172 -3840
rect 7172 -3972 7210 -3840
rect 7210 -3972 7218 -3840
rect 7430 -3972 7438 -3840
rect 7438 -3972 7476 -3840
rect 7476 -3972 7484 -3840
rect 7696 -3972 7704 -3840
rect 7704 -3972 7742 -3840
rect 7742 -3972 7750 -3840
rect 7962 -3972 7970 -3840
rect 7970 -3972 8008 -3840
rect 8008 -3972 8016 -3840
rect 8228 -3972 8236 -3840
rect 8236 -3972 8274 -3840
rect 8274 -3972 8282 -3840
rect 8494 -3972 8502 -3840
rect 8502 -3972 8540 -3840
rect 8540 -3972 8548 -3840
rect 13542 -3515 14024 -3316
rect 13542 -3854 13759 -3515
rect 13759 -3854 13797 -3515
rect 13797 -3854 14024 -3515
rect 6632 -4982 6640 -4850
rect 6640 -4982 6678 -4850
rect 6678 -4982 6686 -4850
rect 6898 -4982 6906 -4850
rect 6906 -4982 6944 -4850
rect 6944 -4982 6952 -4850
rect 7164 -4982 7172 -4850
rect 7172 -4982 7210 -4850
rect 7210 -4982 7218 -4850
rect 7430 -4982 7438 -4850
rect 7438 -4982 7476 -4850
rect 7476 -4982 7484 -4850
rect 7696 -4982 7704 -4850
rect 7704 -4982 7742 -4850
rect 7742 -4982 7750 -4850
rect 7962 -4982 7970 -4850
rect 7970 -4982 8008 -4850
rect 8008 -4982 8016 -4850
rect 8228 -4982 8236 -4850
rect 8236 -4982 8274 -4850
rect 8274 -4982 8282 -4850
rect 7330 -5526 7824 -5398
rect 8494 -4982 8502 -4850
rect 8502 -4982 8540 -4850
rect 8540 -4982 8548 -4850
rect 13628 -5698 13910 -5332
rect 6902 -8124 8254 -8012
rect 13754 -8098 14510 -7432
<< metal2 >>
rect 2976 7090 3086 7100
rect 2976 7008 3086 7018
rect 3456 7090 3566 7100
rect 3456 7008 3566 7018
rect 3936 7090 4046 7100
rect 3936 7008 4046 7018
rect 4416 7090 4526 7100
rect 4416 7008 4526 7018
rect 4896 7090 5006 7100
rect 4896 7008 5006 7018
rect 5376 7090 5486 7100
rect 5376 7008 5486 7018
rect 5856 7090 5966 7100
rect 5856 7008 5966 7018
rect 6336 7090 6446 7100
rect 6336 7008 6446 7018
rect 6816 7090 6926 7100
rect 6816 7008 6926 7018
rect 7296 7090 7406 7100
rect 7296 7008 7406 7018
rect 7776 7090 7886 7100
rect 7776 7008 7886 7018
rect 8256 7090 8366 7100
rect 8256 7008 8366 7018
rect 8736 7090 8846 7100
rect 8736 7008 8846 7018
rect 9216 7090 9326 7100
rect 9216 7008 9326 7018
rect 9696 7090 9806 7100
rect 9696 7008 9806 7018
rect 10176 7090 10286 7100
rect 10176 7008 10286 7018
rect 10656 7090 10766 7100
rect 10656 7008 10766 7018
rect 11136 7090 11246 7100
rect 11136 7008 11246 7018
rect 11616 7090 11726 7100
rect 11616 7008 11726 7018
rect 12096 7090 12206 7100
rect 12096 7008 12206 7018
rect 12914 6904 13214 6914
rect 2866 6746 12914 6756
rect 2866 6614 2876 6746
rect 2946 6614 3116 6746
rect 3186 6614 3356 6746
rect 3426 6614 3596 6746
rect 3666 6614 3836 6746
rect 3906 6614 4076 6746
rect 4146 6614 4316 6746
rect 4386 6614 4556 6746
rect 4626 6614 4796 6746
rect 4866 6614 5036 6746
rect 5106 6614 5276 6746
rect 5346 6614 5516 6746
rect 5586 6614 5756 6746
rect 5826 6614 5996 6746
rect 6066 6614 6236 6746
rect 6306 6614 6476 6746
rect 6546 6614 6716 6746
rect 6786 6614 6956 6746
rect 7026 6614 7196 6746
rect 7266 6614 7436 6746
rect 7506 6614 7676 6746
rect 7746 6614 7916 6746
rect 7986 6614 8156 6746
rect 8226 6614 8396 6746
rect 8466 6614 8636 6746
rect 8706 6614 8876 6746
rect 8946 6614 9116 6746
rect 9186 6614 9356 6746
rect 9426 6614 9596 6746
rect 9666 6614 9836 6746
rect 9906 6614 10076 6746
rect 10146 6614 10316 6746
rect 10386 6614 10556 6746
rect 10626 6614 10796 6746
rect 10866 6614 11036 6746
rect 11106 6614 11276 6746
rect 11346 6614 11516 6746
rect 11586 6614 11756 6746
rect 11826 6614 11996 6746
rect 12066 6614 12236 6746
rect 12306 6614 12914 6746
rect 2866 6604 12914 6614
rect 12914 6594 13214 6604
rect 12914 6096 13214 6106
rect 2866 5938 12914 5948
rect 2866 5806 2876 5938
rect 2946 5806 3116 5938
rect 3186 5806 3356 5938
rect 3426 5806 3596 5938
rect 3666 5806 3836 5938
rect 3906 5806 4076 5938
rect 4146 5806 4316 5938
rect 4386 5806 4556 5938
rect 4626 5806 4796 5938
rect 4866 5806 5036 5938
rect 5106 5806 5276 5938
rect 5346 5806 5516 5938
rect 5586 5806 5756 5938
rect 5826 5806 5996 5938
rect 6066 5806 6236 5938
rect 6306 5806 6476 5938
rect 6546 5806 6716 5938
rect 6786 5806 6956 5938
rect 7026 5806 7196 5938
rect 7266 5806 7436 5938
rect 7506 5806 7676 5938
rect 7746 5806 7916 5938
rect 7986 5806 8156 5938
rect 8226 5806 8396 5938
rect 8466 5806 8636 5938
rect 8706 5806 8876 5938
rect 8946 5806 9116 5938
rect 9186 5806 9356 5938
rect 9426 5806 9596 5938
rect 9666 5806 9836 5938
rect 9906 5806 10076 5938
rect 10146 5806 10316 5938
rect 10386 5806 10556 5938
rect 10626 5806 10796 5938
rect 10866 5806 11036 5938
rect 11106 5806 11276 5938
rect 11346 5806 11516 5938
rect 11586 5806 11756 5938
rect 11826 5806 11996 5938
rect 12066 5806 12236 5938
rect 12306 5806 12914 5938
rect 2866 5796 12914 5806
rect 12914 5786 13214 5796
rect 12914 5288 13214 5298
rect 2866 5130 12914 5140
rect 2866 4998 2876 5130
rect 2946 4998 3116 5130
rect 3186 4998 3356 5130
rect 3426 4998 3596 5130
rect 3666 4998 3836 5130
rect 3906 4998 4076 5130
rect 4146 4998 4316 5130
rect 4386 4998 4556 5130
rect 4626 4998 4796 5130
rect 4866 4998 5036 5130
rect 5106 4998 5276 5130
rect 5346 4998 5516 5130
rect 5586 4998 5756 5130
rect 5826 4998 5996 5130
rect 6066 4998 6236 5130
rect 6306 4998 6476 5130
rect 6546 4998 6716 5130
rect 6786 4998 6956 5130
rect 7026 4998 7196 5130
rect 7266 4998 7436 5130
rect 7506 4998 7676 5130
rect 7746 4998 7916 5130
rect 7986 4998 8156 5130
rect 8226 4998 8396 5130
rect 8466 4998 8636 5130
rect 8706 4998 8876 5130
rect 8946 4998 9116 5130
rect 9186 4998 9356 5130
rect 9426 4998 9596 5130
rect 9666 4998 9836 5130
rect 9906 4998 10076 5130
rect 10146 4998 10316 5130
rect 10386 4998 10556 5130
rect 10626 4998 10796 5130
rect 10866 4998 11036 5130
rect 11106 4998 11276 5130
rect 11346 4998 11516 5130
rect 11586 4998 11756 5130
rect 11826 4998 11996 5130
rect 12066 4998 12236 5130
rect 12306 4998 12914 5130
rect 2866 4988 12914 4998
rect 12914 4978 13214 4988
rect 16818 4104 17718 4114
rect 16818 3550 17718 3560
rect -6028 -694 -5840 -684
rect -6028 -814 -5840 -804
rect -4852 -694 -4664 -684
rect -4852 -814 -4664 -804
rect -3676 -694 -3488 -684
rect -3676 -814 -3488 -804
rect -2500 -694 -2312 -684
rect -2500 -814 -2312 -804
rect -1324 -694 -1136 -684
rect -1324 -814 -1136 -804
rect -148 -694 40 -684
rect -148 -814 40 -804
rect 1028 -694 1216 -684
rect 1028 -814 1216 -804
rect 2204 -694 2392 -684
rect 2204 -814 2392 -804
rect 3380 -694 3568 -684
rect 3380 -814 3568 -804
rect 4556 -694 4744 -684
rect 4556 -814 4744 -804
rect 5732 -694 5920 -684
rect 5732 -814 5920 -804
rect 6908 -694 7096 -684
rect 6908 -814 7096 -804
rect 8084 -694 8272 -684
rect 8084 -814 8272 -804
rect 9260 -694 9448 -684
rect 9260 -814 9448 -804
rect 10436 -694 10624 -684
rect 10436 -814 10624 -804
rect 11612 -694 11800 -684
rect 11612 -814 11800 -804
rect 13964 -694 14152 -684
rect 13964 -814 14152 -804
rect 15140 -694 15328 -684
rect 15140 -814 15328 -804
rect 16316 -694 16504 -684
rect 16316 -814 16504 -804
rect 18668 -694 18856 -684
rect 18668 -814 18856 -804
rect 19844 -694 20032 -684
rect 19844 -814 20032 -804
rect 21020 -694 21208 -684
rect 21020 -814 21208 -804
rect 7164 -1696 9204 -1570
rect 7164 -1810 7484 -1696
rect 6632 -1820 6952 -1810
rect 6686 -1952 6898 -1820
rect 6632 -2076 6952 -1952
rect 7164 -1820 7218 -1810
rect 7164 -1962 7218 -1952
rect 7430 -1820 7484 -1810
rect 7430 -1962 7484 -1952
rect 7696 -1820 8016 -1696
rect 7750 -1952 7962 -1820
rect 7696 -1958 8016 -1952
rect 8228 -1820 8282 -1810
rect 8228 -1958 8282 -1952
rect 8494 -1820 8548 -1810
rect 8494 -1958 8548 -1952
rect 8228 -2076 8548 -1958
rect 5976 -2202 8548 -2076
rect 5976 -3086 6086 -2202
rect 9094 -2580 9204 -1696
rect 7164 -2706 9204 -2580
rect 7164 -2820 7484 -2706
rect 7704 -2820 8024 -2706
rect 6632 -2830 6686 -2820
rect 6632 -2972 6686 -2962
rect 6898 -2830 6952 -2820
rect 6898 -2972 6952 -2962
rect 7164 -2830 7218 -2820
rect 7164 -2972 7218 -2962
rect 7430 -2830 7484 -2820
rect 7430 -2972 7484 -2962
rect 7696 -2830 7750 -2820
rect 7696 -2972 7750 -2962
rect 7962 -2830 8016 -2820
rect 7962 -2972 8016 -2962
rect 8228 -2830 8282 -2820
rect 8228 -2972 8282 -2962
rect 8494 -2830 8548 -2820
rect 8494 -2972 8548 -2962
rect 6632 -3086 6952 -2972
rect 8228 -3086 8548 -2972
rect 5976 -3212 8548 -3086
rect 5976 -4096 6086 -3212
rect 9094 -3590 9204 -2706
rect 7164 -3716 9204 -3590
rect 7164 -3830 7484 -3716
rect 6632 -3840 6686 -3830
rect 6632 -3982 6686 -3972
rect 6898 -3840 6952 -3830
rect 6898 -3982 6952 -3972
rect 7164 -3840 7218 -3830
rect 7164 -3982 7218 -3972
rect 7430 -3840 7484 -3830
rect 7430 -3982 7484 -3972
rect 7696 -3834 8016 -3716
rect 7696 -3840 7750 -3834
rect 7696 -3982 7750 -3972
rect 7962 -3840 8016 -3834
rect 7962 -3982 8016 -3972
rect 8228 -3840 8282 -3830
rect 8228 -3982 8282 -3972
rect 8494 -3840 8548 -3830
rect 8494 -3982 8548 -3972
rect 6632 -4096 6952 -3982
rect 8228 -4096 8548 -3982
rect 5976 -4222 8548 -4096
rect 5976 -5106 6086 -4222
rect 9094 -4600 9204 -3716
rect 13542 -3316 14024 -3306
rect 14848 -3352 15436 -3342
rect 14024 -3672 14848 -3506
rect 13542 -3864 14024 -3854
rect 14848 -3910 15436 -3900
rect 7164 -4726 9204 -4600
rect 7164 -4840 7484 -4726
rect 6632 -4850 6686 -4840
rect 6632 -4992 6686 -4982
rect 6898 -4850 6952 -4840
rect 6898 -4992 6952 -4982
rect 7164 -4850 7218 -4840
rect 7164 -4992 7218 -4982
rect 7430 -4850 7484 -4840
rect 7430 -4992 7484 -4982
rect 7696 -4840 8016 -4726
rect 7696 -4850 7750 -4840
rect 7696 -4992 7750 -4982
rect 7962 -4850 8016 -4840
rect 7962 -4992 8016 -4982
rect 8228 -4850 8282 -4840
rect 8228 -4992 8282 -4982
rect 8494 -4850 8548 -4840
rect 8494 -4992 8548 -4982
rect 6632 -5106 6952 -4992
rect 8228 -5106 8548 -4992
rect 5976 -5232 8548 -5106
rect 12686 -4944 13466 -4934
rect 7330 -5398 12686 -5388
rect 7824 -5526 12686 -5398
rect 7330 -5536 12686 -5526
rect 13628 -5332 13910 -5322
rect 13466 -5536 13628 -5388
rect 13628 -5708 13910 -5698
rect 12686 -5764 13466 -5754
rect 13754 -7432 14510 -7422
rect 6902 -8012 8254 -8002
rect 13754 -8108 14510 -8098
rect 6902 -8134 8254 -8124
<< via2 >>
rect 2976 7018 3086 7090
rect 3456 7018 3566 7090
rect 3936 7018 4046 7090
rect 4416 7018 4526 7090
rect 4896 7018 5006 7090
rect 5376 7018 5486 7090
rect 5856 7018 5966 7090
rect 6336 7018 6446 7090
rect 6816 7018 6926 7090
rect 7296 7018 7406 7090
rect 7776 7018 7886 7090
rect 8256 7018 8366 7090
rect 8736 7018 8846 7090
rect 9216 7018 9326 7090
rect 9696 7018 9806 7090
rect 10176 7018 10286 7090
rect 10656 7018 10766 7090
rect 11136 7018 11246 7090
rect 11616 7018 11726 7090
rect 12096 7018 12206 7090
rect 12914 6604 13214 6904
rect 12914 5796 13214 6096
rect 12914 4988 13214 5288
rect 16818 3560 17718 4104
rect -6028 -804 -5840 -694
rect -4852 -804 -4664 -694
rect -3676 -804 -3488 -694
rect -2500 -804 -2312 -694
rect -1324 -804 -1136 -694
rect -148 -804 40 -694
rect 1028 -804 1216 -694
rect 2204 -804 2392 -694
rect 3380 -804 3568 -694
rect 4556 -804 4744 -694
rect 5732 -804 5920 -694
rect 6908 -804 7096 -694
rect 8084 -804 8272 -694
rect 9260 -804 9448 -694
rect 10436 -804 10624 -694
rect 11612 -804 11800 -694
rect 13964 -804 14152 -694
rect 15140 -804 15328 -694
rect 16316 -804 16504 -694
rect 18668 -804 18856 -694
rect 19844 -804 20032 -694
rect 21020 -804 21208 -694
rect 14848 -3900 15436 -3352
rect 12686 -5754 13466 -4944
rect 6902 -8124 8254 -8012
rect 13754 -8098 14510 -7432
<< metal3 >>
rect 2966 7090 3096 7095
rect 2966 7018 2976 7090
rect 3086 7018 3096 7090
rect 2966 7013 3096 7018
rect 3446 7090 3576 7095
rect 3446 7018 3456 7090
rect 3566 7018 3576 7090
rect 3446 7013 3576 7018
rect 3926 7090 4056 7095
rect 3926 7018 3936 7090
rect 4046 7018 4056 7090
rect 3926 7013 4056 7018
rect 4406 7090 4536 7095
rect 4406 7018 4416 7090
rect 4526 7018 4536 7090
rect 4406 7013 4536 7018
rect 4886 7090 5016 7095
rect 4886 7018 4896 7090
rect 5006 7018 5016 7090
rect 4886 7013 5016 7018
rect 5366 7090 5496 7095
rect 5366 7018 5376 7090
rect 5486 7018 5496 7090
rect 5366 7013 5496 7018
rect 5846 7090 5976 7095
rect 5846 7018 5856 7090
rect 5966 7018 5976 7090
rect 5846 7013 5976 7018
rect 6326 7090 6456 7095
rect 6326 7018 6336 7090
rect 6446 7018 6456 7090
rect 6326 7013 6456 7018
rect 6806 7090 6936 7095
rect 6806 7018 6816 7090
rect 6926 7018 6936 7090
rect 6806 7013 6936 7018
rect 7286 7090 7416 7095
rect 7286 7018 7296 7090
rect 7406 7018 7416 7090
rect 7286 7013 7416 7018
rect 7766 7090 7896 7095
rect 7766 7018 7776 7090
rect 7886 7018 7896 7090
rect 7766 7013 7896 7018
rect 8246 7090 8376 7095
rect 8246 7018 8256 7090
rect 8366 7018 8376 7090
rect 8246 7013 8376 7018
rect 8726 7090 8856 7095
rect 8726 7018 8736 7090
rect 8846 7018 8856 7090
rect 8726 7013 8856 7018
rect 9206 7090 9336 7095
rect 9206 7018 9216 7090
rect 9326 7018 9336 7090
rect 9206 7013 9336 7018
rect 9686 7090 9816 7095
rect 9686 7018 9696 7090
rect 9806 7018 9816 7090
rect 9686 7013 9816 7018
rect 10166 7090 10296 7095
rect 10166 7018 10176 7090
rect 10286 7018 10296 7090
rect 10166 7013 10296 7018
rect 10646 7090 10776 7095
rect 10646 7018 10656 7090
rect 10766 7018 10776 7090
rect 10646 7013 10776 7018
rect 11126 7090 11256 7095
rect 11126 7018 11136 7090
rect 11246 7018 11256 7090
rect 11126 7013 11256 7018
rect 11606 7090 11736 7095
rect 11606 7018 11616 7090
rect 11726 7018 11736 7090
rect 11606 7013 11736 7018
rect 12086 7090 12216 7095
rect 12086 7018 12096 7090
rect 12206 7018 12216 7090
rect 12086 7013 12216 7018
rect 12904 6908 13224 6909
rect 12904 6904 13234 6908
rect 12904 6604 12914 6904
rect 13214 6604 13234 6904
rect 12904 6599 13234 6604
rect 12914 6101 13234 6599
rect 12904 6096 13234 6101
rect 12904 5796 12914 6096
rect 13214 5796 13234 6096
rect 12904 5791 13234 5796
rect 12914 5293 13234 5791
rect 12904 5288 13234 5293
rect 12904 4988 12914 5288
rect 13214 4988 13234 5288
rect 12904 4983 13234 4988
rect -6038 -694 -5830 -689
rect -6038 -804 -6028 -694
rect -5840 -804 -5830 -694
rect -6038 -809 -5830 -804
rect -4862 -694 -4654 -689
rect -4862 -804 -4852 -694
rect -4664 -804 -4654 -694
rect -4862 -809 -4654 -804
rect -3686 -694 -3478 -689
rect -3686 -804 -3676 -694
rect -3488 -804 -3478 -694
rect -3686 -809 -3478 -804
rect -2510 -694 -2302 -689
rect -2510 -804 -2500 -694
rect -2312 -804 -2302 -694
rect -2510 -809 -2302 -804
rect -1334 -694 -1126 -689
rect -1334 -804 -1324 -694
rect -1136 -804 -1126 -694
rect -1334 -809 -1126 -804
rect -158 -694 50 -689
rect -158 -804 -148 -694
rect 40 -804 50 -694
rect -158 -809 50 -804
rect 1018 -694 1226 -689
rect 1018 -804 1028 -694
rect 1216 -804 1226 -694
rect 1018 -809 1226 -804
rect 2194 -694 2402 -689
rect 2194 -804 2204 -694
rect 2392 -804 2402 -694
rect 2194 -809 2402 -804
rect 3370 -694 3578 -689
rect 3370 -804 3380 -694
rect 3568 -804 3578 -694
rect 3370 -809 3578 -804
rect 4546 -694 4754 -689
rect 4546 -804 4556 -694
rect 4744 -804 4754 -694
rect 4546 -809 4754 -804
rect 5722 -694 5930 -689
rect 5722 -804 5732 -694
rect 5920 -804 5930 -694
rect 5722 -809 5930 -804
rect 6898 -694 7106 -689
rect 6898 -804 6908 -694
rect 7096 -804 7106 -694
rect 6898 -809 7106 -804
rect 8074 -694 8282 -689
rect 8074 -804 8084 -694
rect 8272 -804 8282 -694
rect 8074 -809 8282 -804
rect 9250 -694 9458 -689
rect 9250 -804 9260 -694
rect 9448 -804 9458 -694
rect 9250 -809 9458 -804
rect 10426 -694 10634 -689
rect 10426 -804 10436 -694
rect 10624 -804 10634 -694
rect 10426 -809 10634 -804
rect 11602 -694 11810 -689
rect 11602 -804 11612 -694
rect 11800 -804 11810 -694
rect 11602 -809 11810 -804
rect 12914 -4939 13234 4983
rect 16808 4104 17728 4109
rect 16808 3560 16818 4104
rect 17718 3560 17728 4104
rect 16808 3555 17728 3560
rect 13954 -694 14162 -689
rect 13954 -804 13964 -694
rect 14152 -804 14162 -694
rect 13954 -809 14162 -804
rect 15130 -694 15338 -689
rect 15130 -804 15140 -694
rect 15328 -804 15338 -694
rect 15130 -809 15338 -804
rect 16306 -694 16514 -689
rect 16306 -804 16316 -694
rect 16504 -804 16514 -694
rect 16306 -809 16514 -804
rect 16862 -1564 17700 3555
rect 18658 -694 18866 -689
rect 18658 -804 18668 -694
rect 18856 -804 18866 -694
rect 18658 -809 18866 -804
rect 19834 -694 20042 -689
rect 19834 -804 19844 -694
rect 20032 -804 20042 -694
rect 19834 -809 20042 -804
rect 21010 -694 21218 -689
rect 21010 -804 21020 -694
rect 21208 -804 21218 -694
rect 21010 -809 21218 -804
rect 16824 -2464 16834 -1564
rect 17734 -2464 17744 -1564
rect 14838 -3352 15446 -3347
rect 14838 -3900 14848 -3352
rect 15436 -3508 15446 -3352
rect 16026 -3508 21990 -2592
rect 15436 -3820 21990 -3508
rect 15436 -3900 15446 -3820
rect 14838 -3905 15446 -3900
rect 12676 -4944 13476 -4939
rect 12676 -5754 12686 -4944
rect 13466 -5754 13476 -4944
rect 12676 -5759 13476 -5754
rect 13744 -7432 14520 -7427
rect 6892 -8012 8264 -8007
rect 6892 -8124 6902 -8012
rect 8254 -8124 8264 -8012
rect 13744 -8098 13754 -7432
rect 14510 -8098 14520 -7432
rect 13744 -8103 14520 -8098
rect 6892 -8129 8264 -8124
rect 16026 -8592 21990 -3820
<< via3 >>
rect 2976 7018 3086 7090
rect 3456 7018 3566 7090
rect 3936 7018 4046 7090
rect 4416 7018 4526 7090
rect 4896 7018 5006 7090
rect 5376 7018 5486 7090
rect 5856 7018 5966 7090
rect 6336 7018 6446 7090
rect 6816 7018 6926 7090
rect 7296 7018 7406 7090
rect 7776 7018 7886 7090
rect 8256 7018 8366 7090
rect 8736 7018 8846 7090
rect 9216 7018 9326 7090
rect 9696 7018 9806 7090
rect 10176 7018 10286 7090
rect 10656 7018 10766 7090
rect 11136 7018 11246 7090
rect 11616 7018 11726 7090
rect 12096 7018 12206 7090
rect -6028 -804 -5840 -694
rect -4852 -804 -4664 -694
rect -3676 -804 -3488 -694
rect -2500 -804 -2312 -694
rect -1324 -804 -1136 -694
rect -148 -804 40 -694
rect 1028 -804 1216 -694
rect 2204 -804 2392 -694
rect 3380 -804 3568 -694
rect 4556 -804 4744 -694
rect 5732 -804 5920 -694
rect 6908 -804 7096 -694
rect 8084 -804 8272 -694
rect 9260 -804 9448 -694
rect 10436 -804 10624 -694
rect 11612 -804 11800 -694
rect 13964 -804 14152 -694
rect 15140 -804 15328 -694
rect 16316 -804 16504 -694
rect 18668 -804 18856 -694
rect 19844 -804 20032 -694
rect 21020 -804 21208 -694
rect 16834 -2464 17734 -1564
rect 6902 -8124 8254 -8012
rect 13754 -8098 14510 -7432
<< mimcap >>
rect 16126 -2732 21926 -2692
rect 16126 -8452 16166 -2732
rect 21886 -8452 21926 -2732
rect 16126 -8492 21926 -8452
<< mimcapcontact >>
rect 16166 -8452 21886 -2732
<< metal4 >>
rect -17050 7090 18658 7796
rect -17050 7018 2976 7090
rect 3086 7018 3456 7090
rect 3566 7018 3936 7090
rect 4046 7018 4416 7090
rect 4526 7018 4896 7090
rect 5006 7018 5376 7090
rect 5486 7018 5856 7090
rect 5966 7018 6336 7090
rect 6446 7018 6816 7090
rect 6926 7018 7296 7090
rect 7406 7018 7776 7090
rect 7886 7018 8256 7090
rect 8366 7018 8736 7090
rect 8846 7018 9216 7090
rect 9326 7018 9696 7090
rect 9806 7018 10176 7090
rect 10286 7018 10656 7090
rect 10766 7018 11136 7090
rect 11246 7018 11616 7090
rect 11726 7018 12096 7090
rect 12206 7018 18658 7090
rect -17050 6796 18658 7018
rect -17048 6532 18658 6796
rect -17048 6530 -3176 6532
rect -17048 -7118 -15438 6530
rect -8052 -694 22432 170
rect -8052 -804 -6028 -694
rect -5840 -804 -4852 -694
rect -4664 -804 -3676 -694
rect -3488 -804 -2500 -694
rect -2312 -804 -1324 -694
rect -1136 -804 -148 -694
rect 40 -804 1028 -694
rect 1216 -804 2204 -694
rect 2392 -804 3380 -694
rect 3568 -804 4556 -694
rect 4744 -804 5732 -694
rect 5920 -804 6908 -694
rect 7096 -804 8084 -694
rect 8272 -804 9260 -694
rect 9448 -804 10436 -694
rect 10624 -804 11612 -694
rect 11800 -804 13964 -694
rect 14152 -804 15140 -694
rect 15328 -804 16316 -694
rect 16504 -804 18668 -694
rect 18856 -804 19844 -694
rect 20032 -804 21020 -694
rect 21208 -804 22432 -694
rect -8052 -1362 22432 -804
rect 16833 -1564 17735 -1563
rect 16833 -2464 16834 -1564
rect 17734 -2464 17735 -1564
rect 16833 -2465 17735 -2464
rect 16890 -2731 17692 -2465
rect 16165 -2732 21887 -2731
rect -17048 -7432 14920 -7118
rect -17048 -8012 13754 -7432
rect -17048 -8124 6902 -8012
rect 8254 -8098 13754 -8012
rect 14510 -8098 14920 -7432
rect 8254 -8124 14920 -8098
rect -17048 -8650 14920 -8124
rect 16165 -8452 16166 -2732
rect 21886 -8452 21887 -2732
rect 16165 -8453 21887 -8452
<< labels >>
flabel metal4 -7878 -506 -7878 -506 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal4 -7394 -8256 -7394 -8256 0 FreeSans 1600 0 0 0 vss
port 4 nsew
flabel metal1 20222 3748 20222 3748 0 FreeSans 1600 0 0 0 vout
port 5 nsew
flabel metal1 -6254 552 -6254 552 0 FreeSans 1600 0 0 0 vbias
port 3 nsew
flabel metal2 6022 -2964 6022 -2964 0 FreeSans 1600 0 0 0 vn
port 2 nsew
flabel metal2 9132 -2620 9132 -2620 0 FreeSans 1600 0 0 0 vp
port 1 nsew
<< end >>
