* NGSPICE file created from OTA_int_revised_post.ext - technology: sky130A

.subckt OTA_int_revised_post vdd vp vn vbias vss vout
X0 vdd.t95 vbias.t48 vout.t66 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1 vss.t63 a_21167_3051.t33 vout.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2 vss.t62 a_21167_3051.t34 vout.t108 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3 vss.t61 a_21167_3051.t35 vout.t109 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4 vout.t2 a_21167_3051.t36 vss.t60 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5 w_20027_5063.t17 vn.t0 a_20223_2963.t0 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6 a_21167_3051.t0 vp.t0 w_20027_5063.t0 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7 a_21167_3051.t11 a_20223_2963.t48 vss.t85 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8 vdd.t94 vbias.t40 vbias.t41 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9 w_20027_5063.t50 vp.t1 a_21167_3051.t23 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10 vss.t78 a_20223_2963.t49 a_21167_3051.t9 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X11 a_20223_2963.t13 vn.t1 w_20027_5063.t16 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X12 vout.t3 a_21167_3051.t37 vss.t59 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X13 w_20027_5063.t41 vbias.t49 vdd.t93 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14 a_20223_2963.t47 a_20223_2963.t46 vss.t75 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X15 vdd.t92 vbias.t2 vbias.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X16 w_20027_5063.t40 vbias.t50 vdd.t91 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X17 vdd.t90 vbias.t51 vout.t61 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X18 vss.t58 a_21167_3051.t38 vout.t106 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X19 vout.t107 a_21167_3051.t39 vss.t57 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X20 vss.t56 a_21167_3051.t40 vout.t31 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X21 vout.t49 vbias.t52 vdd.t89 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X22 vss.t55 a_21167_3051.t41 vout.t32 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X23 vout.t11 a_21167_3051.t42 vss.t54 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X24 w_20027_5063.t15 vn.t2 a_20223_2963.t14 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X25 vdd.t88 vbias.t53 vout.t63 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X26 vdd.t87 vbias.t10 vbias.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X27 w_20027_5063.t39 vbias.t54 vdd.t86 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X28 vout.t50 vbias.t55 vdd.t85 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X29 vdd.t84 vbias.t56 w_20027_5063.t38 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X30 a_20223_2963.t9 vn.t3 w_20027_5063.t14 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X31 vss.t53 a_21167_3051.t43 vout.t12 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X32 a_21167_3051.t8 a_20223_2963.t50 vss.t76 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X33 vdd.t83 vbias.t57 w_20027_5063.t37 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X34 vdd.t82 vbias.t58 vout.t67 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X35 vout.t104 a_21167_3051.t44 vss.t52 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X36 vout.t105 a_21167_3051.t45 vss.t51 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X37 vss.t70 a_20223_2963.t44 a_20223_2963.t45 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X38 vout.t37 vbias.t59 vdd.t81 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X39 vss.t50 a_21167_3051.t46 vout.t92 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X40 vdd.t80 vbias.t60 vout.t52 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X41 w_20027_5063.t36 vbias.t61 vdd.t79 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X42 vout.t93 a_21167_3051.t47 vss.t49 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X43 vdd.t78 vbias.t62 w_20027_5063.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X44 vout.t79 vbias.t63 vdd.t77 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X45 w_20027_5063.t13 vn.t4 a_20223_2963.t10 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X46 w_20027_5063.t49 vp.t2 a_21167_3051.t22 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X47 vss.t82 a_20223_2963.t42 a_20223_2963.t43 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X48 vbias.t45 vbias.t44 vdd.t76 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X49 a_21167_3051.t21 vp.t3 w_20027_5063.t48 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X50 vss.t48 a_21167_3051.t48 vout.t25 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X51 vbias.t7 vbias.t6 vdd.t75 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X52 vout.t26 a_21167_3051.t49 vss.t47 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X53 vss.t80 a_20223_2963.t40 a_20223_2963.t41 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X54 vout.t102 a_21167_3051.t50 vss.t46 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X55 vdd.t74 vbias.t64 w_20027_5063.t34 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X56 vout.t38 vbias.t65 vdd.t73 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X57 vss.t45 a_21167_3051.t51 vout.t103 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X58 vout.t96 a_21167_3051.t52 vss.t44 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X59 vout.t97 a_21167_3051.t53 vss.t43 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X60 vout.t80 vbias.t66 vdd.t72 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X61 vdd.t71 vbias.t67 vout.t81 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X62 a_21167_3051.t20 vp.t4 w_20027_5063.t47 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X63 vout.t90 a_21167_3051.t54 vss.t42 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X64 w_20027_5063.t46 vp.t5 a_21167_3051.t19 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X65 vdd.t70 vbias.t28 vbias.t29 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X66 vdd.t69 vbias.t68 vout.t68 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X67 vbias.t31 vbias.t30 vdd.t68 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X68 vdd.t67 vbias.t69 vout.t39 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X69 a_20223_2963.t11 vn.t5 w_20027_5063.t12 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X70 vdd.t66 vbias.t14 vbias.t15 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X71 vout.t91 a_21167_3051.t55 vss.t41 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X72 vss.t40 a_21167_3051.t56 vout.t23 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X73 vout.t69 vbias.t70 vdd.t65 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X74 a_21167_3051.t12 a_20223_2963.t51 vss.t88 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X75 vout.t40 vbias.t71 vdd.t64 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X76 vss.t89 a_20223_2963.t52 a_21167_3051.t13 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X77 vout.t24 a_21167_3051.t57 vss.t39 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X78 vout.t29 a_21167_3051.t58 vss.t38 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X79 vdd.t63 vbias.t72 vout.t53 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X80 vbias.t23 vbias.t22 vdd.t62 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X81 vout.t51 vbias.t73 vdd.t61 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X82 w_20027_5063.t55 vp.t6 a_21167_3051.t32 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X83 vss.t72 a_20223_2963.t53 a_21167_3051.t7 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X84 a_20223_2963.t1 vn.t6 w_20027_5063.t11 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X85 vout.t41 vbias.t74 vdd.t60 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X86 vbias.t47 vbias.t46 vdd.t59 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X87 vdd.t58 vbias.t8 vbias.t9 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X88 vout.t30 a_21167_3051.t59 vss.t37 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X89 a_23819_6897# vout sky130_fd_pr__cap_mim_m3_1 l=1.4e+07u w=3e+07u
X90 a_21167_3051.t15 a_20223_2963.t54 vss.t91 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X91 vss.t93 a_20223_2963.t55 a_21167_3051.t25 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X92 vss.t83 a_20223_2963.t38 a_20223_2963.t39 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X93 w_20027_5063.t33 vbias.t75 vdd.t57 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X94 vbias.t13 vbias.t12 vdd.t56 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X95 vout.t70 vbias.t76 vdd.t55 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X96 vout.t9 a_21167_3051.t60 vss.t36 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X97 vout.t10 a_21167_3051.t61 vss.t35 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X98 vss.t34 a_21167_3051.t62 vout.t100 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X99 vout.t48 vbias.t77 vdd.t54 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X100 w_20027_5063.t10 vn.t7 a_20223_2963.t6 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X101 vout.t101 a_21167_3051.t63 vss.t33 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X102 w_20027_5063.t32 vbias.t78 vdd.t53 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X103 vdd.t52 vbias.t32 vbias.t33 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X104 a_21167_3051.t14 vp.t7 w_20027_5063.t42 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X105 a_21167_3051.t2 a_23819_6897# vss sky130_fd_pr__res_xhigh_po w=350000u l=2.8e+06u
X106 a_20223_2963.t12 vn.t8 w_20027_5063.t9 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X107 a_20223_2963.t37 a_20223_2963.t36 vss.t73 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X108 vdd.t51 vbias.t79 vout.t36 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X109 w_20027_5063.t8 vn.t9 a_20223_2963.t2 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X110 w_20027_5063.t31 vbias.t80 vdd.t50 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X111 vdd.t49 vbias.t81 w_20027_5063.t30 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X112 vss.t64 a_20223_2963.t34 a_20223_2963.t35 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X113 vss.t32 a_21167_3051.t64 vout.t88 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X114 vss.t31 a_21167_3051.t65 vout.t89 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X115 vdd.t48 vbias.t82 vout.t54 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X116 vout.t47 vbias.t83 vdd.t47 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X117 vout.t21 a_21167_3051.t66 vss.t30 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X118 vdd.t46 vbias.t84 vout.t71 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X119 vss.t29 a_21167_3051.t67 vout.t22 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X120 vout.t42 vbias.t85 vdd.t45 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X121 vout.t98 a_21167_3051.t68 vss.t28 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X122 a_20223_2963.t7 vn.t10 w_20027_5063.t7 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X123 a_20223_2963.t33 a_20223_2963.t32 vss.t79 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X124 vdd.t44 vbias.t16 vbias.t17 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X125 a_23819_6897# vout sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=1.4e+07u
X126 vss.t27 a_21167_3051.t69 vout.t99 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X127 vdd.t43 vbias.t86 w_20027_5063.t29 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X128 w_20027_5063.t28 vbias.t87 vdd.t42 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X129 vss.t77 a_20223_2963.t30 a_20223_2963.t31 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X130 vout.t43 vbias.t88 vdd.t41 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X131 vss.t26 a_21167_3051.t70 vout.t94 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X132 vss.t25 a_21167_3051.t71 vout.t95 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X133 vss.t95 a_20223_2963.t56 a_21167_3051.t31 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X134 a_21167_3051.t6 a_20223_2963.t57 vss.t69 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X135 vdd.t40 vbias.t89 vout.t55 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X136 vout.t72 vbias.t90 vdd.t39 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X137 vout.t86 a_21167_3051.t72 vss.t24 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X138 vout.t87 a_21167_3051.t73 vss.t23 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X139 w_20027_5063.t54 vp.t8 a_21167_3051.t29 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X140 vbias.t25 vbias.t24 vdd.t38 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X141 vdd.t37 vbias.t91 vout.t56 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X142 vss.t22 a_21167_3051.t74 vout.t19 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X143 a_21167_3051.t28 vp.t9 w_20027_5063.t53 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X144 a_21167_3051.t30 a_20223_2963.t58 vss.t94 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X145 vdd.t36 vbias.t92 w_20027_5063.t27 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X146 vout.t60 vbias.t93 vdd.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X147 vdd.t34 vbias.t94 vout.t44 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X148 a_21167_3051.t18 vp.t10 w_20027_5063.t45 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X149 w_20027_5063.t44 vp.t11 a_21167_3051.t17 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X150 vss.t21 a_21167_3051.t75 vout.t20 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X151 vbias.t19 vbias.t18 vdd.t33 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X152 vss.t66 a_20223_2963.t59 a_21167_3051.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X153 vdd.t32 vbias.t95 vout.t73 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X154 vbias.t27 vbias.t26 vdd.t31 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X155 vss.t20 a_21167_3051.t76 vout.t34 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X156 vss.t19 a_21167_3051.t77 vout.t35 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X157 vout.t27 a_21167_3051.t78 vss.t18 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X158 vout.t57 vbias.t96 vdd.t30 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X159 a_20223_2963.t8 vn.t11 w_20027_5063.t6 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X160 vout.t74 vbias.t97 vdd.t29 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X161 w_20027_5063.t26 vbias.t98 vdd.t28 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X162 w_20027_5063.t5 vn.t12 a_20223_2963.t5 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X163 vss.t84 a_20223_2963.t60 a_21167_3051.t10 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X164 vss.t17 a_21167_3051.t79 vout.t28 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X165 w_20027_5063.t25 vbias.t99 vdd.t27 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X166 vss.t67 a_20223_2963.t28 a_20223_2963.t29 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X167 vout.t84 a_21167_3051.t80 vss.t16 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X168 vdd.t26 vbias.t100 w_20027_5063.t24 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X169 vdd.t25 vbias.t101 vout.t45 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X170 vout.t58 vbias.t102 vdd.t24 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X171 vout.t85 a_21167_3051.t81 vss.t15 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X172 a_20223_2963.t27 a_20223_2963.t26 vss.t87 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X173 vdd.t23 vbias.t34 vbias.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X174 vout.t17 a_21167_3051.t82 vss.t14 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X175 vss.t13 a_21167_3051.t83 vout.t18 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X176 vdd.t22 vbias.t20 vbias.t21 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X177 a_20223_2963.t3 vn.t13 w_20027_5063.t4 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X178 vss.t12 a_21167_3051.t84 vout.t110 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X179 vdd.t21 vbias.t103 vout.t46 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X180 w_20027_5063.t23 vbias.t104 vdd.t20 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X181 vdd.t19 vbias.t105 vout.t75 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X182 vdd.t18 vbias.t4 vbias.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X183 w_20027_5063.t3 vn.t14 a_20223_2963.t15 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X184 vdd.t17 vbias.t106 vout.t59 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X185 vout.t111 a_21167_3051.t85 vss.t11 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X186 vout.t76 vbias.t107 vdd.t16 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X187 a_20223_2963.t25 a_20223_2963.t24 vss.t81 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X188 a_20223_2963.t23 a_20223_2963.t22 vss.t74 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X189 vdd.t15 vbias.t108 vout.t62 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X190 vss.t10 a_21167_3051.t86 vout.t13 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X191 vdd.t14 vbias.t109 w_20027_5063.t22 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X192 a_21167_3051.t27 vp.t12 w_20027_5063.t52 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X193 vss.t9 a_21167_3051.t87 vout.t14 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X194 vss.t8 a_21167_3051.t88 vout.t15 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X195 vss.t7 a_21167_3051.t89 vout.t16 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X196 w_20027_5063.t21 vbias.t110 vdd.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X197 w_20027_5063.t2 vn.t15 a_20223_2963.t4 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X198 vbias.t43 vbias.t42 vdd.t12 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X199 vout.t112 a_21167_3051.t90 vss.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X200 vss.t71 a_20223_2963.t20 a_20223_2963.t21 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X201 vdd.t11 vbias.t111 w_20027_5063.t20 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X202 a_21167_3051.t1 vp.t13 w_20027_5063.t1 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X203 w_20027_5063.t43 vp.t14 a_21167_3051.t16 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X204 vout.t64 vbias.t112 vdd.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X205 vout.t82 vbias.t113 vdd.t9 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X206 a_20223_2963.t19 a_20223_2963.t18 vss.t90 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X207 vss.t65 a_20223_2963.t61 a_21167_3051.t3 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X208 vbias.t37 vbias.t36 vdd.t8 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X209 vss.t5 a_21167_3051.t91 vout.t113 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X210 vout.t0 a_21167_3051.t92 vss.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X211 a_21167_3051.t24 a_20223_2963.t62 vss.t92 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X212 vdd.t7 vbias.t114 vout.t77 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X213 vout.t1 a_21167_3051.t93 vss.t3 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X214 vss.t2 a_21167_3051.t94 vout.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X215 vss.t1 a_21167_3051.t95 vout.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X216 vout.t78 vbias.t115 vdd.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X217 vdd.t5 vbias.t116 w_20027_5063.t19 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X218 vbias.t1 vbias.t0 vdd.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X219 vdd.t3 vbias.t38 vbias.t39 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X220 vdd.t2 vbias.t117 vout.t65 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X221 w_20027_5063.t51 vp.t15 a_21167_3051.t26 w_20027_5063# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X222 vout.t33 a_21167_3051.t96 vss.t0 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X223 vdd.t1 vbias.t118 w_20027_5063.t18 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X224 a_21167_3051.t5 a_20223_2963.t63 vss.t68 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X225 vdd.t0 vbias.t119 vout.t83 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X226 a_20223_2963.t17 a_20223_2963.t16 vss.t86 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
C0 a_23819_6897# vout 80.16fF
C1 vdd vbias 34.89fF
C2 vdd vout 13.17fF
C3 vbias vout 9.70fF
C4 vn vp 1.91fF
R0 vbias.n128 vbias.t8 63.632
R1 vbias.n195 vbias.t20 63.63
R2 vbias.n87 vbias.t2 63.63
R3 vbias.n194 vbias.t75 63.63
R4 vbias.n19 vbias.t97 63.63
R5 vbias.n105 vbias.t74 63.63
R6 vbias.n105 vbias.t59 63.63
R7 vbias.n20 vbias.t68 63.63
R8 vbias.n106 vbias.t117 63.63
R9 vbias.n106 vbias.t84 63.63
R10 vbias.n18 vbias.t103 63.63
R11 vbias.n104 vbias.t79 63.63
R12 vbias.n104 vbias.t106 63.63
R13 vbias.n21 vbias.t85 63.63
R14 vbias.n107 vbias.t63 63.63
R15 vbias.n107 vbias.t52 63.63
R16 vbias.n23 vbias.t96 63.63
R17 vbias.n109 vbias.t73 63.63
R18 vbias.n109 vbias.t76 63.63
R19 vbias.n24 vbias.t114 63.63
R20 vbias.n110 vbias.t91 63.63
R21 vbias.n110 vbias.t48 63.63
R22 vbias.n22 vbias.t53 63.63
R23 vbias.n108 vbias.t105 63.63
R24 vbias.n108 vbias.t51 63.63
R25 vbias.n25 vbias.t66 63.63
R26 vbias.n111 vbias.t115 63.63
R27 vbias.n111 vbias.t65 63.63
R28 vbias.n27 vbias.t77 63.63
R29 vbias.n113 vbias.t55 63.63
R30 vbias.n113 vbias.t88 63.63
R31 vbias.n28 vbias.t95 63.63
R32 vbias.n114 vbias.t72 63.63
R33 vbias.n114 vbias.t58 63.63
R34 vbias.n26 vbias.t82 63.63
R35 vbias.n112 vbias.t60 63.63
R36 vbias.n112 vbias.t108 63.63
R37 vbias.n29 vbias.t112 63.63
R38 vbias.n115 vbias.t90 63.63
R39 vbias.n115 vbias.t102 63.63
R40 vbias.n31 vbias.t107 63.63
R41 vbias.n117 vbias.t83 63.63
R42 vbias.n117 vbias.t70 63.63
R43 vbias.n32 vbias.t69 63.63
R44 vbias.n118 vbias.t119 63.63
R45 vbias.n118 vbias.t94 63.63
R46 vbias.n30 vbias.t89 63.63
R47 vbias.n116 vbias.t67 63.63
R48 vbias.n116 vbias.t101 63.63
R49 vbias.n63 vbias.t104 63.63
R50 vbias.n126 vbias.t80 63.63
R51 vbias.n126 vbias.t49 63.63
R52 vbias.n159 vbias.t46 63.63
R53 vbias.n159 vbias.t18 63.63
R54 vbias.n77 vbias.t0 63.63
R55 vbias.n64 vbias.t28 63.63
R56 vbias.n103 vbias.t38 63.63
R57 vbias.n62 vbias.t86 63.63
R58 vbias.n125 vbias.t64 63.63
R59 vbias.n125 vbias.t81 63.63
R60 vbias.n33 vbias.t93 63.63
R61 vbias.n119 vbias.t71 63.63
R62 vbias.n119 vbias.t113 63.63
R63 vbias.n123 vbias.t6 63.63
R64 vbias.n35 vbias.t44 63.63
R65 vbias.n123 vbias.t36 63.63
R66 vbias.n78 vbias.t62 63.63
R67 vbias.n161 vbias.t111 63.63
R68 vbias.n161 vbias.t118 63.63
R69 vbias.n83 vbias.t116 63.63
R70 vbias.n188 vbias.t92 63.63
R71 vbias.n188 vbias.t56 63.63
R72 vbias.n189 vbias.t98 63.63
R73 vbias.n190 vbias.t40 63.63
R74 vbias.n192 vbias.t12 63.63
R75 vbias.n192 vbias.t22 63.63
R76 vbias.n85 vbias.t34 63.63
R77 vbias.n190 vbias.t32 63.63
R78 vbias.n163 vbias.t4 63.63
R79 vbias.n80 vbias.t10 63.63
R80 vbias.n82 vbias.t24 63.63
R81 vbias.n186 vbias.t30 63.63
R82 vbias.n163 vbias.t16 63.63
R83 vbias.n186 vbias.t42 63.63
R84 vbias.n79 vbias.t78 63.63
R85 vbias.n162 vbias.t54 63.63
R86 vbias.n162 vbias.t87 63.63
R87 vbias.n90 vbias.t57 63.63
R88 vbias.n193 vbias.t109 63.63
R89 vbias.n193 vbias.t100 63.63
R90 vbias.n194 vbias.t50 63.63
R91 vbias.n189 vbias.t110 63.63
R92 vbias.n84 vbias.t61 63.63
R93 vbias.n91 vbias.t26 63.63
R94 vbias.n89 vbias.t99 63.63
R95 vbias.n195 vbias.t14 63.63
R96 vbias.n0 vbias.t21 14.295
R97 vbias.n9 vbias.t3 14.295
R98 vbias.n156 vbias.t47 14.295
R99 vbias.n156 vbias.t9 14.295
R100 vbias.n132 vbias.t39 14.295
R101 vbias.n132 vbias.t19 14.295
R102 vbias.n74 vbias.t29 14.295
R103 vbias.n74 vbias.t1 14.295
R104 vbias.n134 vbias.t7 14.295
R105 vbias.n53 vbias.t45 14.295
R106 vbias.n56 vbias.t37 14.295
R107 vbias.n101 vbias.t13 14.295
R108 vbias.n101 vbias.t41 14.295
R109 vbias.n94 vbias.t33 14.295
R110 vbias.n94 vbias.t23 14.295
R111 vbias.n17 vbias.t35 14.295
R112 vbias.n17 vbias.t27 14.295
R113 vbias.n183 vbias.t17 14.295
R114 vbias.n183 vbias.t43 14.295
R115 vbias.n173 vbias.t5 14.295
R116 vbias.n173 vbias.t31 14.295
R117 vbias.n171 vbias.t25 14.295
R118 vbias.n171 vbias.t11 14.295
R119 vbias.n3 vbias.t15 14.295
R120 vbias.n196 vbias.n0 3.25
R121 vbias.n196 vbias.n3 1.139
R122 vbias.n3 vbias.n2 0.874
R123 vbias.n10 vbias.n9 0.87
R124 vbias.n53 vbias.n52 0.823
R125 vbias.n150 vbias.n134 0.823
R126 vbias.n54 vbias.n53 0.594
R127 vbias.n57 vbias.n56 0.58
R128 vbias.n13 vbias.n12 0.577
R129 vbias.n37 vbias.n36 0.575
R130 vbias.n38 vbias.n37 0.575
R131 vbias.n39 vbias.n38 0.575
R132 vbias.n41 vbias.n40 0.575
R133 vbias.n42 vbias.n41 0.575
R134 vbias.n40 vbias.n39 0.575
R135 vbias.n43 vbias.n42 0.575
R136 vbias.n45 vbias.n44 0.575
R137 vbias.n46 vbias.n45 0.575
R138 vbias.n44 vbias.n43 0.575
R139 vbias.n47 vbias.n46 0.575
R140 vbias.n49 vbias.n48 0.575
R141 vbias.n50 vbias.n49 0.575
R142 vbias.n48 vbias.n47 0.575
R143 vbias.n66 vbias.n65 0.575
R144 vbias.n152 vbias.n151 0.575
R145 vbias.n167 vbias.n166 0.575
R146 vbias.n5 vbias.n4 0.575
R147 vbias.n2 vbias.n1 0.575
R148 vbias.n138 vbias.n137 0.574
R149 vbias.n139 vbias.n138 0.574
R150 vbias.n142 vbias.n141 0.574
R151 vbias.n143 vbias.n142 0.574
R152 vbias.n146 vbias.n145 0.574
R153 vbias.n147 vbias.n146 0.574
R154 vbias.n67 vbias.n66 0.574
R155 vbias.n153 vbias.n152 0.574
R156 vbias.n96 vbias.n95 0.574
R157 vbias.n168 vbias.n167 0.574
R158 vbias.n175 vbias.n174 0.574
R159 vbias.n176 vbias.n175 0.574
R160 vbias.n12 vbias.n11 0.574
R161 vbias.n6 vbias.n5 0.574
R162 vbias.n11 vbias.n10 0.574
R163 vbias.n137 vbias.n136 0.574
R164 vbias.n141 vbias.n140 0.574
R165 vbias.n145 vbias.n144 0.574
R166 vbias.n149 vbias.n148 0.574
R167 vbias.n136 vbias.n135 0.573
R168 vbias.n140 vbias.n139 0.573
R169 vbias.n144 vbias.n143 0.573
R170 vbias.n148 vbias.n147 0.573
R171 vbias.n154 vbias.n153 0.573
R172 vbias.n98 vbias.n97 0.573
R173 vbias.n99 vbias.n98 0.573
R174 vbias.n52 vbias.n50 0.57
R175 vbias.n150 vbias.n149 0.569
R176 vbias.n73 vbias.n68 0.376
R177 vbias.n16 vbias.n7 0.376
R178 vbias.n182 vbias.n177 0.376
R179 vbias.n156 vbias.n155 0.337
R180 vbias.n171 vbias.n170 0.337
R181 vbias.n101 vbias.n100 0.332
R182 vbias.n188 vbias.n187 0.284
R183 vbias.n161 vbias.n160 0.284
R184 vbias.n125 vbias.n124 0.284
R185 vbias.n78 vbias.n77 0.281
R186 vbias.n193 vbias.n192 0.281
R187 vbias.n83 vbias.n82 0.281
R188 vbias.n20 vbias.n19 0.281
R189 vbias.n106 vbias.n105 0.281
R190 vbias.n21 vbias.n20 0.281
R191 vbias.n107 vbias.n106 0.281
R192 vbias.n19 vbias.n18 0.281
R193 vbias.n105 vbias.n104 0.281
R194 vbias.n22 vbias.n21 0.281
R195 vbias.n108 vbias.n107 0.281
R196 vbias.n24 vbias.n23 0.281
R197 vbias.n110 vbias.n109 0.281
R198 vbias.n25 vbias.n24 0.281
R199 vbias.n111 vbias.n110 0.281
R200 vbias.n23 vbias.n22 0.281
R201 vbias.n109 vbias.n108 0.281
R202 vbias.n26 vbias.n25 0.281
R203 vbias.n112 vbias.n111 0.281
R204 vbias.n28 vbias.n27 0.281
R205 vbias.n114 vbias.n113 0.281
R206 vbias.n29 vbias.n28 0.281
R207 vbias.n115 vbias.n114 0.281
R208 vbias.n27 vbias.n26 0.281
R209 vbias.n113 vbias.n112 0.281
R210 vbias.n30 vbias.n29 0.281
R211 vbias.n116 vbias.n115 0.281
R212 vbias.n32 vbias.n31 0.281
R213 vbias.n118 vbias.n117 0.281
R214 vbias.n33 vbias.n32 0.281
R215 vbias.n119 vbias.n118 0.281
R216 vbias.n31 vbias.n30 0.281
R217 vbias.n117 vbias.n116 0.281
R218 vbias.n63 vbias.n62 0.281
R219 vbias.n126 vbias.n125 0.281
R220 vbias.n79 vbias.n78 0.281
R221 vbias.n162 vbias.n161 0.281
R222 vbias.n84 vbias.n83 0.281
R223 vbias.n189 vbias.n188 0.281
R224 vbias.n91 vbias.n90 0.281
R225 vbias.n194 vbias.n193 0.281
R226 vbias.n85 vbias.n84 0.281
R227 vbias.n90 vbias.n89 0.281
R228 vbias.n64 vbias.n63 0.281
R229 vbias.n89 vbias.n88 0.281
R230 vbias.n62 vbias.n61 0.281
R231 vbias.n190 vbias.n189 0.28
R232 vbias.n163 vbias.n162 0.28
R233 vbias.n80 vbias.n79 0.28
R234 vbias.n195 vbias.n194 0.28
R235 vbias.n102 vbias.n94 0.234
R236 vbias.n94 vbias.n93 0.231
R237 vbias.n93 vbias.n17 0.231
R238 vbias.n74 vbias.n73 0.229
R239 vbias.n17 vbias.n16 0.229
R240 vbias.n183 vbias.n182 0.229
R241 vbias.n157 vbias.n132 0.227
R242 vbias.n75 vbias.n74 0.227
R243 vbias.n157 vbias.n156 0.227
R244 vbias.n102 vbias.n101 0.227
R245 vbias.n184 vbias.n173 0.227
R246 vbias.n173 vbias.n172 0.227
R247 vbias.n172 vbias.n171 0.227
R248 vbias.n184 vbias.n183 0.227
R249 vbias.n127 vbias.n126 0.217
R250 vbias.n34 vbias.n33 0.217
R251 vbias.n120 vbias.n119 0.217
R252 vbias.n131 vbias.n130 0.215
R253 vbias.n165 vbias.n164 0.215
R254 vbias.n73 vbias.n72 0.212
R255 vbias.n16 vbias.n15 0.212
R256 vbias.n182 vbias.n181 0.212
R257 vbias.n72 vbias.n71 0.175
R258 vbias.n15 vbias.n14 0.175
R259 vbias.n181 vbias.n180 0.175
R260 vbias.n155 vbias.n133 0.167
R261 vbias.n170 vbias.n169 0.167
R262 vbias.n155 vbias.n154 0.167
R263 vbias.n170 vbias.n168 0.167
R264 vbias.n100 vbias.n96 0.165
R265 vbias.n100 vbias.n99 0.164
R266 vbias.n179 vbias.n178 0.132
R267 vbias.n70 vbias.n69 0.132
R268 vbias.n13 vbias.n8 0.132
R269 vbias.n88 vbias.n86 0.09
R270 vbias.n196 vbias.n195 0.085
R271 vbias.n158 vbias.n157 0.081
R272 vbias.n185 vbias.n184 0.081
R273 vbias.n92 vbias.n91 0.074
R274 vbias.n192 vbias.n191 0.074
R275 vbias.n191 vbias.n190 0.074
R276 vbias.n92 vbias.n85 0.074
R277 vbias.n77 vbias.n76 0.073
R278 vbias.n82 vbias.n81 0.073
R279 vbias.n76 vbias.n64 0.073
R280 vbias.n81 vbias.n80 0.073
R281 vbias.n123 vbias.n122 0.068
R282 vbias.n159 vbias.n158 0.067
R283 vbias.n186 vbias.n185 0.067
R284 vbias.n124 vbias.n120 0.065
R285 vbias.n160 vbias.n131 0.065
R286 vbias.n187 vbias.n165 0.065
R287 vbias.n128 vbias.n127 0.064
R288 vbias.n55 vbias.n34 0.064
R289 vbias.n93 vbias.n92 0.039
R290 vbias.n191 vbias.n102 0.038
R291 vbias.n76 vbias.n75 0.038
R292 vbias vbias.n196 0.021
R293 vbias.n58 vbias.n57 0.014
R294 vbias.n177 vbias.n176 0.005
R295 vbias.n68 vbias.n67 0.005
R296 vbias.n7 vbias.n6 0.005
R297 vbias.n151 vbias.n150 0.005
R298 vbias.n52 vbias.n51 0.005
R299 vbias.n164 vbias.n163 0.002
R300 vbias.n130 vbias.n129 0.002
R301 vbias.n55 vbias.n54 0.001
R302 vbias.n59 vbias.n58 0.001
R303 vbias.n180 vbias.n179 0.001
R304 vbias.n129 vbias.n128 0.001
R305 vbias.n122 vbias.n121 0.001
R306 vbias.n61 vbias.n60 0.001
R307 vbias.n88 vbias.n87 0.001
R308 vbias.n129 vbias.n103 0.001
R309 vbias.n54 vbias.n35 0.001
R310 vbias.n160 vbias.n159 0.001
R311 vbias.n71 vbias.n70 0.001
R312 vbias.n124 vbias.n123 0.001
R313 vbias.n14 vbias.n13 0.001
R314 vbias.n187 vbias.n186 0.001
R315 vbias.n60 vbias.n59 0.001
R316 vbias.n59 vbias.n55 0.001
R317 vout.n70 vout.t16 17.43
R318 vout.n70 vout.t93 17.43
R319 vout.n69 vout.t94 17.43
R320 vout.n69 vout.t0 17.43
R321 vout.n68 vout.t32 17.43
R322 vout.n68 vout.t101 17.43
R323 vout.n67 vout.t5 17.43
R324 vout.n67 vout.t97 17.43
R325 vout.n64 vout.t110 17.43
R326 vout.n64 vout.t2 17.43
R327 vout.n63 vout.t89 17.43
R328 vout.n63 vout.t84 17.43
R329 vout.n62 vout.t109 17.43
R330 vout.n62 vout.t90 17.43
R331 vout.n61 vout.t14 17.43
R332 vout.n61 vout.t107 17.43
R333 vout.n58 vout.t19 17.43
R334 vout.n58 vout.t29 17.43
R335 vout.n57 vout.t23 17.43
R336 vout.n57 vout.t3 17.43
R337 vout.n56 vout.t15 17.43
R338 vout.n56 vout.t87 17.43
R339 vout.n55 vout.t34 17.43
R340 vout.n55 vout.t9 17.43
R341 vout.n33 vout.t6 17.43
R342 vout.n33 vout.t98 17.43
R343 vout.n32 vout.t20 17.43
R344 vout.n32 vout.t102 17.43
R345 vout.n31 vout.t92 17.43
R346 vout.n31 vout.t17 17.43
R347 vout.n30 vout.t4 17.43
R348 vout.n30 vout.t86 17.43
R349 vout.n37 vout.t22 17.43
R350 vout.n37 vout.t11 17.43
R351 vout.n36 vout.t25 17.43
R352 vout.n36 vout.t111 17.43
R353 vout.n35 vout.t18 17.43
R354 vout.n35 vout.t24 17.43
R355 vout.n34 vout.t95 17.43
R356 vout.n34 vout.t104 17.43
R357 vout.n41 vout.t100 17.43
R358 vout.n41 vout.t27 17.43
R359 vout.n40 vout.t12 17.43
R360 vout.n40 vout.t30 17.43
R361 vout.n39 vout.t35 17.43
R362 vout.n39 vout.t1 17.43
R363 vout.n38 vout.t88 17.43
R364 vout.n38 vout.t85 17.43
R365 vout.n45 vout.t108 17.43
R366 vout.n45 vout.t96 17.43
R367 vout.n44 vout.t28 17.43
R368 vout.n44 vout.t33 17.43
R369 vout.n43 vout.t103 17.43
R370 vout.n43 vout.t21 17.43
R371 vout.n42 vout.t106 17.43
R372 vout.n42 vout.t91 17.43
R373 vout.n49 vout.t13 17.43
R374 vout.n49 vout.t105 17.43
R375 vout.n48 vout.t99 17.43
R376 vout.n48 vout.t112 17.43
R377 vout.n47 vout.t31 17.43
R378 vout.n47 vout.t10 17.43
R379 vout.n46 vout.t113 17.43
R380 vout.n46 vout.t26 17.43
R381 vout.n24 vout.t44 14.295
R382 vout.n24 vout.t82 14.295
R383 vout.n23 vout.t83 14.295
R384 vout.n23 vout.t40 14.295
R385 vout.n22 vout.t60 14.295
R386 vout.n22 vout.t39 14.295
R387 vout.n21 vout.t69 14.295
R388 vout.n21 vout.t45 14.295
R389 vout.n20 vout.t47 14.295
R390 vout.n20 vout.t81 14.295
R391 vout.n19 vout.t76 14.295
R392 vout.n19 vout.t55 14.295
R393 vout.n17 vout.t43 14.295
R394 vout.n17 vout.t62 14.295
R395 vout.n16 vout.t50 14.295
R396 vout.n16 vout.t52 14.295
R397 vout.n15 vout.t48 14.295
R398 vout.n15 vout.t54 14.295
R399 vout.n13 vout.t38 14.295
R400 vout.n13 vout.t66 14.295
R401 vout.n12 vout.t78 14.295
R402 vout.n12 vout.t56 14.295
R403 vout.n11 vout.t80 14.295
R404 vout.n11 vout.t77 14.295
R405 vout.n2 vout.t70 14.295
R406 vout.n2 vout.t61 14.295
R407 vout.n1 vout.t51 14.295
R408 vout.n1 vout.t75 14.295
R409 vout.n0 vout.t57 14.295
R410 vout.n0 vout.t63 14.295
R411 vout.n5 vout.t49 14.295
R412 vout.n5 vout.t71 14.295
R413 vout.n4 vout.t79 14.295
R414 vout.n4 vout.t65 14.295
R415 vout.n3 vout.t42 14.295
R416 vout.n3 vout.t68 14.295
R417 vout.n8 vout.t37 14.295
R418 vout.n8 vout.t59 14.295
R419 vout.n7 vout.t41 14.295
R420 vout.n7 vout.t36 14.295
R421 vout.n6 vout.t74 14.295
R422 vout.n6 vout.t46 14.295
R423 vout.n28 vout.t58 14.295
R424 vout.n28 vout.t67 14.295
R425 vout.n27 vout.t72 14.295
R426 vout.n27 vout.t53 14.295
R427 vout.n26 vout.t64 14.295
R428 vout.n26 vout.t73 14.295
R429 vout.n50 vout.n49 1.558
R430 vout.n25 vout.n24 1.247
R431 vout.n9 vout.n8 1.247
R432 vout.n71 vout.n70 1.107
R433 vout.n65 vout.n64 1.107
R434 vout.n59 vout.n58 1.107
R435 vout.n53 vout.n33 1.107
R436 vout.n52 vout.n37 1.107
R437 vout.n51 vout.n41 1.107
R438 vout.n50 vout.n45 1.107
R439 vout.n25 vout.n21 0.929
R440 vout.n18 vout.n17 0.929
R441 vout.n14 vout.n13 0.929
R442 vout.n10 vout.n2 0.929
R443 vout.n9 vout.n5 0.929
R444 vout.n29 vout.n28 0.929
R445 vout.n23 vout.n22 0.733
R446 vout.n24 vout.n23 0.733
R447 vout.n20 vout.n19 0.733
R448 vout.n21 vout.n20 0.733
R449 vout.n16 vout.n15 0.733
R450 vout.n17 vout.n16 0.733
R451 vout.n12 vout.n11 0.733
R452 vout.n13 vout.n12 0.733
R453 vout.n1 vout.n0 0.733
R454 vout.n2 vout.n1 0.733
R455 vout.n4 vout.n3 0.733
R456 vout.n5 vout.n4 0.733
R457 vout.n7 vout.n6 0.733
R458 vout.n8 vout.n7 0.733
R459 vout.n27 vout.n26 0.733
R460 vout.n28 vout.n27 0.733
R461 vout.n68 vout.n67 0.545
R462 vout.n69 vout.n68 0.545
R463 vout.n70 vout.n69 0.545
R464 vout.n62 vout.n61 0.545
R465 vout.n63 vout.n62 0.545
R466 vout.n64 vout.n63 0.545
R467 vout.n56 vout.n55 0.545
R468 vout.n57 vout.n56 0.545
R469 vout.n58 vout.n57 0.545
R470 vout.n31 vout.n30 0.545
R471 vout.n32 vout.n31 0.545
R472 vout.n33 vout.n32 0.545
R473 vout.n35 vout.n34 0.545
R474 vout.n36 vout.n35 0.545
R475 vout.n37 vout.n36 0.545
R476 vout.n39 vout.n38 0.545
R477 vout.n40 vout.n39 0.545
R478 vout.n41 vout.n40 0.545
R479 vout.n43 vout.n42 0.545
R480 vout.n44 vout.n43 0.545
R481 vout.n45 vout.n44 0.545
R482 vout.n47 vout.n46 0.545
R483 vout.n48 vout.n47 0.545
R484 vout.n49 vout.n48 0.545
R485 vout.n51 vout.n50 0.451
R486 vout.n52 vout.n51 0.451
R487 vout.n53 vout.n52 0.451
R488 vout.n10 vout.n9 0.318
R489 vout.n29 vout.n25 0.318
R490 vout.n66 vout.n65 0.13
R491 vout.n60 vout.n59 0.13
R492 vout.n54 vout.n53 0.13
R493 vout.n72 vout.n71 0.13
R494 vout vout.n72 0.098
R495 vout.n60 vout.n18 0.053
R496 vout.n66 vout.n14 0.053
R497 vout.n72 vout.n10 0.053
R498 vout.n54 vout.n29 0.053
R499 vout.n72 vout.n66 0.011
R500 vout.n66 vout.n60 0.011
R501 vout.n60 vout.n54 0.011
R502 vdd.n118 vdd.n117 386.601
R503 vdd.n103 vdd.n101 127.023
R504 vdd.n98 vdd.n96 127.023
R505 vdd.n87 vdd.n85 127.023
R506 vdd.n82 vdd.n80 127.023
R507 vdd.n71 vdd.n69 127.023
R508 vdd.n66 vdd.n64 127.023
R509 vdd.n45 vdd.n43 127.023
R510 vdd.n40 vdd.n38 127.023
R511 vdd.n29 vdd.n27 127.023
R512 vdd.n24 vdd.n22 127.023
R513 vdd.n13 vdd.n11 127.023
R514 vdd.n8 vdd.n4 127.023
R515 vdd.n8 vdd.n6 127.023
R516 vdd.n122 vdd.n120 116.986
R517 vdd.n57 vdd.t9 15.566
R518 vdd.n114 vdd.t17 15.351
R519 vdd.n144 vdd.t27 14.295
R520 vdd.n144 vdd.t92 14.295
R521 vdd.n143 vdd.t57 14.295
R522 vdd.n143 vdd.t22 14.295
R523 vdd.n142 vdd.t91 14.295
R524 vdd.n142 vdd.t66 14.295
R525 vdd.n2 vdd.t31 14.295
R526 vdd.n2 vdd.t83 14.295
R527 vdd.n1 vdd.t62 14.295
R528 vdd.n1 vdd.t14 14.295
R529 vdd.n0 vdd.t56 14.295
R530 vdd.n0 vdd.t26 14.295
R531 vdd.n16 vdd.t79 14.295
R532 vdd.n16 vdd.t23 14.295
R533 vdd.n15 vdd.t13 14.295
R534 vdd.n15 vdd.t52 14.295
R535 vdd.n14 vdd.t28 14.295
R536 vdd.n14 vdd.t94 14.295
R537 vdd.n20 vdd.t38 14.295
R538 vdd.n20 vdd.t5 14.295
R539 vdd.n19 vdd.t68 14.295
R540 vdd.n19 vdd.t36 14.295
R541 vdd.n18 vdd.t12 14.295
R542 vdd.n18 vdd.t84 14.295
R543 vdd.n32 vdd.t53 14.295
R544 vdd.n32 vdd.t87 14.295
R545 vdd.n31 vdd.t86 14.295
R546 vdd.n31 vdd.t18 14.295
R547 vdd.n30 vdd.t42 14.295
R548 vdd.n30 vdd.t44 14.295
R549 vdd.n36 vdd.t4 14.295
R550 vdd.n36 vdd.t78 14.295
R551 vdd.n35 vdd.t33 14.295
R552 vdd.n35 vdd.t11 14.295
R553 vdd.n34 vdd.t59 14.295
R554 vdd.n34 vdd.t1 14.295
R555 vdd.n48 vdd.t20 14.295
R556 vdd.n48 vdd.t70 14.295
R557 vdd.n47 vdd.t50 14.295
R558 vdd.n47 vdd.t3 14.295
R559 vdd.n46 vdd.t93 14.295
R560 vdd.n46 vdd.t58 14.295
R561 vdd.n52 vdd.t76 14.295
R562 vdd.n52 vdd.t43 14.295
R563 vdd.n51 vdd.t8 14.295
R564 vdd.n51 vdd.t74 14.295
R565 vdd.n50 vdd.t75 14.295
R566 vdd.n50 vdd.t49 14.295
R567 vdd.n58 vdd.t35 14.295
R568 vdd.n57 vdd.t64 14.295
R569 vdd.n62 vdd.t16 14.295
R570 vdd.n62 vdd.t67 14.295
R571 vdd.n61 vdd.t47 14.295
R572 vdd.n61 vdd.t0 14.295
R573 vdd.n60 vdd.t65 14.295
R574 vdd.n60 vdd.t34 14.295
R575 vdd.n74 vdd.t10 14.295
R576 vdd.n74 vdd.t40 14.295
R577 vdd.n73 vdd.t39 14.295
R578 vdd.n73 vdd.t71 14.295
R579 vdd.n72 vdd.t24 14.295
R580 vdd.n72 vdd.t25 14.295
R581 vdd.n78 vdd.t54 14.295
R582 vdd.n78 vdd.t32 14.295
R583 vdd.n77 vdd.t85 14.295
R584 vdd.n77 vdd.t63 14.295
R585 vdd.n76 vdd.t41 14.295
R586 vdd.n76 vdd.t82 14.295
R587 vdd.n90 vdd.t72 14.295
R588 vdd.n90 vdd.t48 14.295
R589 vdd.n89 vdd.t6 14.295
R590 vdd.n89 vdd.t80 14.295
R591 vdd.n88 vdd.t73 14.295
R592 vdd.n88 vdd.t15 14.295
R593 vdd.n94 vdd.t30 14.295
R594 vdd.n94 vdd.t7 14.295
R595 vdd.n93 vdd.t61 14.295
R596 vdd.n93 vdd.t37 14.295
R597 vdd.n92 vdd.t55 14.295
R598 vdd.n92 vdd.t95 14.295
R599 vdd.n106 vdd.t45 14.295
R600 vdd.n106 vdd.t88 14.295
R601 vdd.n105 vdd.t77 14.295
R602 vdd.n105 vdd.t19 14.295
R603 vdd.n104 vdd.t89 14.295
R604 vdd.n104 vdd.t90 14.295
R605 vdd.n110 vdd.t29 14.295
R606 vdd.n110 vdd.t69 14.295
R607 vdd.n109 vdd.t60 14.295
R608 vdd.n109 vdd.t2 14.295
R609 vdd.n108 vdd.t81 14.295
R610 vdd.n108 vdd.t46 14.295
R611 vdd.n115 vdd.t21 14.295
R612 vdd.n114 vdd.t51 14.295
R613 vdd.n58 vdd.n57 1.271
R614 vdd.n115 vdd.n114 1.056
R615 vdd.n143 vdd.n142 0.733
R616 vdd.n144 vdd.n143 0.733
R617 vdd.n1 vdd.n0 0.733
R618 vdd.n2 vdd.n1 0.733
R619 vdd.n15 vdd.n14 0.733
R620 vdd.n16 vdd.n15 0.733
R621 vdd.n19 vdd.n18 0.733
R622 vdd.n20 vdd.n19 0.733
R623 vdd.n31 vdd.n30 0.733
R624 vdd.n32 vdd.n31 0.733
R625 vdd.n35 vdd.n34 0.733
R626 vdd.n36 vdd.n35 0.733
R627 vdd.n47 vdd.n46 0.733
R628 vdd.n48 vdd.n47 0.733
R629 vdd.n51 vdd.n50 0.733
R630 vdd.n52 vdd.n51 0.733
R631 vdd.n61 vdd.n60 0.733
R632 vdd.n62 vdd.n61 0.733
R633 vdd.n73 vdd.n72 0.733
R634 vdd.n74 vdd.n73 0.733
R635 vdd.n77 vdd.n76 0.733
R636 vdd.n78 vdd.n77 0.733
R637 vdd.n89 vdd.n88 0.733
R638 vdd.n90 vdd.n89 0.733
R639 vdd.n93 vdd.n92 0.733
R640 vdd.n94 vdd.n93 0.733
R641 vdd.n105 vdd.n104 0.733
R642 vdd.n106 vdd.n105 0.733
R643 vdd.n109 vdd.n108 0.733
R644 vdd.n110 vdd.n109 0.733
R645 vdd.n59 vdd.n58 0.698
R646 vdd.n116 vdd.n115 0.586
R647 vdd.n145 vdd.n144 0.477
R648 vdd.n17 vdd.n16 0.477
R649 vdd.n33 vdd.n32 0.477
R650 vdd.n49 vdd.n48 0.477
R651 vdd.n75 vdd.n74 0.477
R652 vdd.n91 vdd.n90 0.477
R653 vdd.n107 vdd.n106 0.477
R654 vdd.n113 vdd.n110 0.477
R655 vdd.n99 vdd.n94 0.477
R656 vdd.n83 vdd.n78 0.477
R657 vdd.n67 vdd.n62 0.477
R658 vdd.n55 vdd.n52 0.477
R659 vdd.n41 vdd.n36 0.477
R660 vdd.n25 vdd.n20 0.477
R661 vdd.n9 vdd.n2 0.477
R662 vdd.n133 vdd.n55 0.378
R663 vdd vdd.n145 0.296
R664 vdd.n132 vdd.n59 0.286
R665 vdd.n139 vdd.n9 0.274
R666 vdd.n137 vdd.n25 0.274
R667 vdd.n135 vdd.n41 0.274
R668 vdd.n131 vdd.n67 0.274
R669 vdd.n129 vdd.n83 0.274
R670 vdd.n127 vdd.n99 0.274
R671 vdd.n125 vdd.n113 0.274
R672 vdd.n126 vdd.n107 0.274
R673 vdd.n128 vdd.n91 0.274
R674 vdd.n130 vdd.n75 0.274
R675 vdd.n134 vdd.n49 0.274
R676 vdd.n136 vdd.n33 0.274
R677 vdd.n138 vdd.n17 0.274
R678 vdd.n125 vdd.n124 0.261
R679 vdd.n123 vdd.n122 0.212
R680 vdd.n122 vdd.n121 0.212
R681 vdd.n112 vdd.n111 0.195
R682 vdd.n103 vdd.n102 0.195
R683 vdd.n98 vdd.n97 0.195
R684 vdd.n87 vdd.n86 0.195
R685 vdd.n82 vdd.n81 0.195
R686 vdd.n71 vdd.n70 0.195
R687 vdd.n45 vdd.n44 0.195
R688 vdd.n40 vdd.n39 0.195
R689 vdd.n29 vdd.n28 0.195
R690 vdd.n24 vdd.n23 0.195
R691 vdd.n13 vdd.n12 0.195
R692 vdd.n8 vdd.n7 0.195
R693 vdd.n126 vdd.n125 0.034
R694 vdd.n127 vdd.n126 0.034
R695 vdd.n128 vdd.n127 0.034
R696 vdd.n129 vdd.n128 0.034
R697 vdd.n130 vdd.n129 0.034
R698 vdd.n131 vdd.n130 0.034
R699 vdd.n132 vdd.n131 0.034
R700 vdd.n134 vdd.n133 0.034
R701 vdd.n135 vdd.n134 0.034
R702 vdd.n136 vdd.n135 0.034
R703 vdd.n137 vdd.n136 0.034
R704 vdd.n138 vdd.n137 0.034
R705 vdd.n139 vdd.n138 0.034
R706 vdd.n124 vdd.n123 0.027
R707 vdd.n66 vdd.n65 0.018
R708 vdd.n133 vdd.n132 0.017
R709 vdd.n141 vdd.n140 0.017
R710 vdd.n54 vdd.n53 0.017
R711 vdd vdd.n139 0.011
R712 vdd.n123 vdd.n118 0.001
R713 vdd.n120 vdd.n119 0.001
R714 vdd.n101 vdd.n100 0.001
R715 vdd.n96 vdd.n95 0.001
R716 vdd.n85 vdd.n84 0.001
R717 vdd.n80 vdd.n79 0.001
R718 vdd.n69 vdd.n68 0.001
R719 vdd.n64 vdd.n63 0.001
R720 vdd.n43 vdd.n42 0.001
R721 vdd.n38 vdd.n37 0.001
R722 vdd.n27 vdd.n26 0.001
R723 vdd.n22 vdd.n21 0.001
R724 vdd.n11 vdd.n10 0.001
R725 vdd.n4 vdd.n3 0.001
R726 vdd.n6 vdd.n5 0.001
R727 vdd.n59 vdd.n56 0.001
R728 vdd.n113 vdd.n112 0.001
R729 vdd.n107 vdd.n103 0.001
R730 vdd.n99 vdd.n98 0.001
R731 vdd.n91 vdd.n87 0.001
R732 vdd.n83 vdd.n82 0.001
R733 vdd.n75 vdd.n71 0.001
R734 vdd.n67 vdd.n66 0.001
R735 vdd.n55 vdd.n54 0.001
R736 vdd.n49 vdd.n45 0.001
R737 vdd.n41 vdd.n40 0.001
R738 vdd.n33 vdd.n29 0.001
R739 vdd.n25 vdd.n24 0.001
R740 vdd.n17 vdd.n13 0.001
R741 vdd.n9 vdd.n8 0.001
R742 vdd.n145 vdd.n141 0.001
R743 vdd.n118 vdd.n116 0.001
R744 a_21167_3051.n4 a_21167_3051.t2 154.596
R745 a_21167_3051.n2 a_21167_3051.t53 37.361
R746 a_21167_3051.n7 a_21167_3051.t63 37.361
R747 a_21167_3051.n5 a_21167_3051.t92 37.361
R748 a_21167_3051.n2 a_21167_3051.t87 37.361
R749 a_21167_3051.n7 a_21167_3051.t35 37.361
R750 a_21167_3051.n5 a_21167_3051.t65 37.361
R751 a_21167_3051.n2 a_21167_3051.t39 37.361
R752 a_21167_3051.n7 a_21167_3051.t54 37.361
R753 a_21167_3051.n5 a_21167_3051.t80 37.361
R754 a_21167_3051.n2 a_21167_3051.t76 37.361
R755 a_21167_3051.n7 a_21167_3051.t88 37.361
R756 a_21167_3051.n5 a_21167_3051.t56 37.361
R757 a_21167_3051.n2 a_21167_3051.t60 37.361
R758 a_21167_3051.n4 a_21167_3051.t73 37.361
R759 a_21167_3051.n5 a_21167_3051.t37 37.361
R760 a_21167_3051.n2 a_21167_3051.t33 37.361
R761 a_21167_3051.n4 a_21167_3051.t46 37.361
R762 a_21167_3051.n5 a_21167_3051.t75 37.361
R763 a_21167_3051.n2 a_21167_3051.t72 37.361
R764 a_21167_3051.n4 a_21167_3051.t82 37.361
R765 a_21167_3051.n5 a_21167_3051.t50 37.361
R766 a_21167_3051.n2 a_21167_3051.t71 37.361
R767 a_21167_3051.n4 a_21167_3051.t83 37.361
R768 a_21167_3051.n5 a_21167_3051.t48 37.361
R769 a_21167_3051.n4 a_21167_3051.t44 37.361
R770 a_21167_3051.n4 a_21167_3051.t57 37.361
R771 a_21167_3051.n5 a_21167_3051.t85 37.361
R772 a_21167_3051.n4 a_21167_3051.t64 37.361
R773 a_21167_3051.n4 a_21167_3051.t77 37.361
R774 a_21167_3051.n5 a_21167_3051.t43 37.361
R775 a_21167_3051.n4 a_21167_3051.t81 37.361
R776 a_21167_3051.n4 a_21167_3051.t93 37.361
R777 a_21167_3051.n5 a_21167_3051.t59 37.361
R778 a_21167_3051.n4 a_21167_3051.t38 37.361
R779 a_21167_3051.n4 a_21167_3051.t51 37.361
R780 a_21167_3051.n5 a_21167_3051.t79 37.361
R781 a_21167_3051.n4 a_21167_3051.t55 37.361
R782 a_21167_3051.n4 a_21167_3051.t66 37.361
R783 a_21167_3051.n4 a_21167_3051.t96 37.361
R784 a_21167_3051.n4 a_21167_3051.t91 37.361
R785 a_21167_3051.n4 a_21167_3051.t40 37.361
R786 a_21167_3051.n4 a_21167_3051.t69 37.361
R787 a_21167_3051.n4 a_21167_3051.t49 37.361
R788 a_21167_3051.n4 a_21167_3051.t61 37.361
R789 a_21167_3051.n4 a_21167_3051.t90 37.361
R790 a_21167_3051.n4 a_21167_3051.t45 37.361
R791 a_21167_3051.n5 a_21167_3051.t89 37.361
R792 a_21167_3051.n4 a_21167_3051.t52 37.361
R793 a_21167_3051.n4 a_21167_3051.t86 37.361
R794 a_21167_3051.n5 a_21167_3051.t62 37.361
R795 a_21167_3051.n5 a_21167_3051.t78 37.361
R796 a_21167_3051.n5 a_21167_3051.t68 37.361
R797 a_21167_3051.n5 a_21167_3051.t67 37.361
R798 a_21167_3051.n5 a_21167_3051.t74 37.361
R799 a_21167_3051.n5 a_21167_3051.t58 37.361
R800 a_21167_3051.n5 a_21167_3051.t47 37.361
R801 a_21167_3051.n5 a_21167_3051.t84 37.361
R802 a_21167_3051.n5 a_21167_3051.t36 37.361
R803 a_21167_3051.n5 a_21167_3051.t95 37.361
R804 a_21167_3051.n5 a_21167_3051.t42 37.361
R805 a_21167_3051.n5 a_21167_3051.t34 37.361
R806 a_21167_3051.n5 a_21167_3051.t70 37.361
R807 a_21167_3051.n7 a_21167_3051.t41 37.361
R808 a_21167_3051.n2 a_21167_3051.t94 37.361
R809 a_21167_3051.n1 a_21167_3051.t13 17.43
R810 a_21167_3051.n1 a_21167_3051.t12 17.43
R811 a_21167_3051.n1 a_21167_3051.t9 17.43
R812 a_21167_3051.n1 a_21167_3051.t11 17.43
R813 a_21167_3051.n1 a_21167_3051.t31 17.43
R814 a_21167_3051.n1 a_21167_3051.t6 17.43
R815 a_21167_3051.n1 a_21167_3051.t25 17.43
R816 a_21167_3051.n1 a_21167_3051.t15 17.43
R817 a_21167_3051.n4 a_21167_3051.t4 17.43
R818 a_21167_3051.n4 a_21167_3051.t24 17.43
R819 a_21167_3051.n4 a_21167_3051.t7 17.43
R820 a_21167_3051.n4 a_21167_3051.t30 17.43
R821 a_21167_3051.n6 a_21167_3051.t3 17.43
R822 a_21167_3051.n6 a_21167_3051.t8 17.43
R823 a_21167_3051.n6 a_21167_3051.t10 17.43
R824 a_21167_3051.n6 a_21167_3051.t5 17.43
R825 a_21167_3051.n4 a_21167_3051.n9 8.457
R826 a_21167_3051.n1 a_21167_3051.t23 7.146
R827 a_21167_3051.n1 a_21167_3051.t1 7.146
R828 a_21167_3051.n1 a_21167_3051.t16 7.146
R829 a_21167_3051.n1 a_21167_3051.t20 7.146
R830 a_21167_3051.n1 a_21167_3051.t19 7.146
R831 a_21167_3051.n0 a_21167_3051.t18 7.146
R832 a_21167_3051.n0 a_21167_3051.t17 7.146
R833 a_21167_3051.n3 a_21167_3051.t32 7.146
R834 a_21167_3051.n3 a_21167_3051.t28 7.146
R835 a_21167_3051.n3 a_21167_3051.t22 7.146
R836 a_21167_3051.n3 a_21167_3051.t14 7.146
R837 a_21167_3051.n8 a_21167_3051.t29 7.146
R838 a_21167_3051.n8 a_21167_3051.t27 7.146
R839 a_21167_3051.n8 a_21167_3051.t21 7.146
R840 a_21167_3051.n8 a_21167_3051.t26 7.146
R841 a_21167_3051.t0 a_21167_3051.n1 7.146
R842 a_21167_3051.n4 a_21167_3051.n5 4.284
R843 a_21167_3051.n1 a_21167_3051.n0 4.152
R844 a_21167_3051.n4 a_21167_3051.n2 3.928
R845 a_21167_3051.n4 a_21167_3051.n3 3.818
R846 a_21167_3051.n3 a_21167_3051.n8 3.135
R847 a_21167_3051.n4 a_21167_3051.n6 3.082
R848 a_21167_3051.n1 a_21167_3051.n4 3.061
R849 a_21167_3051.n4 a_21167_3051.n7 2.806
R850 vss.n87 vss.n85 127.023
R851 vss.n78 vss.n76 127.023
R852 vss.n69 vss.n67 127.023
R853 vss.n60 vss.n58 127.023
R854 vss.n38 vss.n36 127.023
R855 vss.n29 vss.n27 127.023
R856 vss.n20 vss.n18 127.023
R857 vss.n11 vss.n9 127.023
R858 vss.n6 vss.n4 113.388
R859 vss.n106 vss.n104 112.311
R860 vss.n0 vss.t74 18.06
R861 vss.n100 vss.t7 18.06
R862 vss.n2 vss.t90 17.43
R863 vss.n1 vss.t75 17.43
R864 vss.n0 vss.t79 17.43
R865 vss.n15 vss.t77 17.43
R866 vss.n15 vss.t68 17.43
R867 vss.n14 vss.t67 17.43
R868 vss.n14 vss.t76 17.43
R869 vss.n13 vss.t82 17.43
R870 vss.n13 vss.t94 17.43
R871 vss.n12 vss.t64 17.43
R872 vss.n12 vss.t92 17.43
R873 vss.n24 vss.t84 17.43
R874 vss.n24 vss.t91 17.43
R875 vss.n23 vss.t65 17.43
R876 vss.n23 vss.t69 17.43
R877 vss.n22 vss.t72 17.43
R878 vss.n22 vss.t85 17.43
R879 vss.n21 vss.t66 17.43
R880 vss.n21 vss.t88 17.43
R881 vss.n33 vss.t93 17.43
R882 vss.n33 vss.t81 17.43
R883 vss.n32 vss.t95 17.43
R884 vss.n32 vss.t86 17.43
R885 vss.n31 vss.t78 17.43
R886 vss.n31 vss.t73 17.43
R887 vss.n30 vss.t89 17.43
R888 vss.n30 vss.t87 17.43
R889 vss.n42 vss.t80 17.43
R890 vss.n42 vss.t47 17.43
R891 vss.n41 vss.t83 17.43
R892 vss.n41 vss.t35 17.43
R893 vss.n40 vss.t71 17.43
R894 vss.n40 vss.t6 17.43
R895 vss.n39 vss.t70 17.43
R896 vss.n39 vss.t51 17.43
R897 vss.n49 vss.t5 17.43
R898 vss.n49 vss.t41 17.43
R899 vss.n48 vss.t56 17.43
R900 vss.n48 vss.t30 17.43
R901 vss.n47 vss.t27 17.43
R902 vss.n47 vss.t0 17.43
R903 vss.n46 vss.t10 17.43
R904 vss.n46 vss.t44 17.43
R905 vss.n55 vss.t58 17.43
R906 vss.n55 vss.t15 17.43
R907 vss.n54 vss.t45 17.43
R908 vss.n54 vss.t3 17.43
R909 vss.n53 vss.t17 17.43
R910 vss.n53 vss.t37 17.43
R911 vss.n52 vss.t62 17.43
R912 vss.n52 vss.t18 17.43
R913 vss.n64 vss.t32 17.43
R914 vss.n64 vss.t52 17.43
R915 vss.n63 vss.t19 17.43
R916 vss.n63 vss.t39 17.43
R917 vss.n62 vss.t53 17.43
R918 vss.n62 vss.t11 17.43
R919 vss.n61 vss.t34 17.43
R920 vss.n61 vss.t54 17.43
R921 vss.n73 vss.t25 17.43
R922 vss.n73 vss.t24 17.43
R923 vss.n72 vss.t13 17.43
R924 vss.n72 vss.t14 17.43
R925 vss.n71 vss.t48 17.43
R926 vss.n71 vss.t46 17.43
R927 vss.n70 vss.t29 17.43
R928 vss.n70 vss.t28 17.43
R929 vss.n82 vss.t63 17.43
R930 vss.n82 vss.t36 17.43
R931 vss.n81 vss.t50 17.43
R932 vss.n81 vss.t23 17.43
R933 vss.n80 vss.t21 17.43
R934 vss.n80 vss.t59 17.43
R935 vss.n79 vss.t1 17.43
R936 vss.n79 vss.t38 17.43
R937 vss.n91 vss.t20 17.43
R938 vss.n91 vss.t57 17.43
R939 vss.n90 vss.t8 17.43
R940 vss.n90 vss.t42 17.43
R941 vss.n89 vss.t40 17.43
R942 vss.n89 vss.t16 17.43
R943 vss.n88 vss.t22 17.43
R944 vss.n88 vss.t60 17.43
R945 vss.n98 vss.t9 17.43
R946 vss.n98 vss.t43 17.43
R947 vss.n97 vss.t61 17.43
R948 vss.n97 vss.t33 17.43
R949 vss.n96 vss.t31 17.43
R950 vss.n96 vss.t4 17.43
R951 vss.n95 vss.t12 17.43
R952 vss.n95 vss.t49 17.43
R953 vss.n102 vss.t2 17.43
R954 vss.n101 vss.t55 17.43
R955 vss.n100 vss.t26 17.43
R956 vss.n1 vss.n0 0.63
R957 vss.n2 vss.n1 0.63
R958 vss.n101 vss.n100 0.63
R959 vss.n102 vss.n101 0.63
R960 vss.n13 vss.n12 0.545
R961 vss.n14 vss.n13 0.545
R962 vss.n15 vss.n14 0.545
R963 vss.n22 vss.n21 0.545
R964 vss.n23 vss.n22 0.545
R965 vss.n24 vss.n23 0.545
R966 vss.n31 vss.n30 0.545
R967 vss.n32 vss.n31 0.545
R968 vss.n33 vss.n32 0.545
R969 vss.n40 vss.n39 0.545
R970 vss.n41 vss.n40 0.545
R971 vss.n42 vss.n41 0.545
R972 vss.n47 vss.n46 0.545
R973 vss.n48 vss.n47 0.545
R974 vss.n49 vss.n48 0.545
R975 vss.n53 vss.n52 0.545
R976 vss.n54 vss.n53 0.545
R977 vss.n55 vss.n54 0.545
R978 vss.n62 vss.n61 0.545
R979 vss.n63 vss.n62 0.545
R980 vss.n64 vss.n63 0.545
R981 vss.n71 vss.n70 0.545
R982 vss.n72 vss.n71 0.545
R983 vss.n73 vss.n72 0.545
R984 vss.n80 vss.n79 0.545
R985 vss.n81 vss.n80 0.545
R986 vss.n82 vss.n81 0.545
R987 vss.n89 vss.n88 0.545
R988 vss.n90 vss.n89 0.545
R989 vss.n91 vss.n90 0.545
R990 vss.n96 vss.n95 0.545
R991 vss.n97 vss.n96 0.545
R992 vss.n98 vss.n97 0.545
R993 vss.n16 vss.n15 0.379
R994 vss.n25 vss.n24 0.379
R995 vss.n34 vss.n33 0.379
R996 vss.n43 vss.n42 0.379
R997 vss.n50 vss.n49 0.379
R998 vss.n56 vss.n55 0.379
R999 vss.n65 vss.n64 0.379
R1000 vss.n74 vss.n73 0.379
R1001 vss.n83 vss.n82 0.379
R1002 vss.n92 vss.n91 0.379
R1003 vss.n99 vss.n98 0.379
R1004 vss.n7 vss.n2 0.375
R1005 vss.n106 vss.n102 0.367
R1006 vss.n117 vss.n16 0.197
R1007 vss.n115 vss.n34 0.197
R1008 vss.n113 vss.n50 0.197
R1009 vss.n111 vss.n65 0.197
R1010 vss.n109 vss.n83 0.197
R1011 vss.n107 vss.n99 0.197
R1012 vss.n108 vss.n92 0.197
R1013 vss.n110 vss.n74 0.197
R1014 vss.n112 vss.n56 0.197
R1015 vss.n114 vss.n43 0.197
R1016 vss.n116 vss.n25 0.197
R1017 vss.n94 vss.n93 0.195
R1018 vss.n87 vss.n86 0.195
R1019 vss.n78 vss.n77 0.195
R1020 vss.n69 vss.n68 0.195
R1021 vss.n38 vss.n37 0.195
R1022 vss.n29 vss.n28 0.195
R1023 vss.n20 vss.n19 0.195
R1024 vss.n11 vss.n10 0.195
R1025 vss.n107 vss.n106 0.181
R1026 vss.n118 vss.n7 0.147
R1027 vss vss.n118 0.05
R1028 vss.n108 vss.n107 0.034
R1029 vss.n109 vss.n108 0.034
R1030 vss.n110 vss.n109 0.034
R1031 vss.n111 vss.n110 0.034
R1032 vss.n112 vss.n111 0.034
R1033 vss.n113 vss.n112 0.034
R1034 vss.n114 vss.n113 0.034
R1035 vss.n115 vss.n114 0.034
R1036 vss.n116 vss.n115 0.034
R1037 vss.n117 vss.n116 0.034
R1038 vss.n118 vss.n117 0.033
R1039 vss.n60 vss.n59 0.011
R1040 vss.n45 vss.n44 0.011
R1041 vss.n106 vss.n105 0.008
R1042 vss.n6 vss.n5 0.008
R1043 vss.n104 vss.n103 0.001
R1044 vss.n85 vss.n84 0.001
R1045 vss.n76 vss.n75 0.001
R1046 vss.n67 vss.n66 0.001
R1047 vss.n58 vss.n57 0.001
R1048 vss.n36 vss.n35 0.001
R1049 vss.n27 vss.n26 0.001
R1050 vss.n18 vss.n17 0.001
R1051 vss.n9 vss.n8 0.001
R1052 vss.n4 vss.n3 0.001
R1053 vss.n99 vss.n94 0.001
R1054 vss.n92 vss.n87 0.001
R1055 vss.n83 vss.n78 0.001
R1056 vss.n74 vss.n69 0.001
R1057 vss.n65 vss.n60 0.001
R1058 vss.n56 vss.n51 0.001
R1059 vss.n50 vss.n45 0.001
R1060 vss.n43 vss.n38 0.001
R1061 vss.n34 vss.n29 0.001
R1062 vss.n25 vss.n20 0.001
R1063 vss.n16 vss.n11 0.001
R1064 vss.n7 vss.n6 0.001
R1065 vn.n10 vn.t1 111.977
R1066 vn.n21 vn.t3 111.977
R1067 vn.n10 vn.t9 111.975
R1068 vn.n21 vn.t14 111.975
R1069 vn.n1 vn.t15 111.83
R1070 vn.n7 vn.t2 111.83
R1071 vn.n12 vn.t4 111.83
R1072 vn.n18 vn.t7 111.83
R1073 vn.n8 vn.t11 111.83
R1074 vn.n5 vn.t5 111.83
R1075 vn.n2 vn.t8 111.83
R1076 vn.n4 vn.t12 111.83
R1077 vn.n19 vn.t13 111.83
R1078 vn.n16 vn.t6 111.83
R1079 vn.n13 vn.t10 111.83
R1080 vn.n15 vn.t0 111.83
R1081 vn.n22 vn.n10 2.763
R1082 vn.n9 vn.n6 2.018
R1083 vn.n6 vn.n3 2.018
R1084 vn.n20 vn.n17 2.018
R1085 vn.n17 vn.n14 2.018
R1086 vn.n10 vn.n9 2.016
R1087 vn.n21 vn.n20 2.016
R1088 vn.n3 vn.n0 1.995
R1089 vn.n14 vn.n11 1.995
R1090 vn vn.n22 0.811
R1091 vn.n9 vn.n8 0.14
R1092 vn.n6 vn.n5 0.14
R1093 vn.n3 vn.n2 0.14
R1094 vn.n20 vn.n19 0.14
R1095 vn.n17 vn.n16 0.14
R1096 vn.n14 vn.n13 0.14
R1097 vn.n3 vn.n1 0.139
R1098 vn.n6 vn.n4 0.139
R1099 vn.n9 vn.n7 0.139
R1100 vn.n14 vn.n12 0.139
R1101 vn.n17 vn.n15 0.139
R1102 vn.n20 vn.n18 0.139
R1103 vn.n22 vn.n21 0.133
R1104 a_20223_2963.n0 a_20223_2963.t55 37.361
R1105 a_20223_2963.n2 a_20223_2963.t56 37.361
R1106 a_20223_2963.n7 a_20223_2963.t52 37.361
R1107 a_20223_2963.n4 a_20223_2963.t53 37.361
R1108 a_20223_2963.n1 a_20223_2963.t54 37.361
R1109 a_20223_2963.n4 a_20223_2963.t57 37.361
R1110 a_20223_2963.n4 a_20223_2963.t48 37.361
R1111 a_20223_2963.n6 a_20223_2963.t51 37.361
R1112 a_20223_2963.n7 a_20223_2963.t44 37.361
R1113 a_20223_2963.n7 a_20223_2963.t26 37.361
R1114 a_20223_2963.n2 a_20223_2963.t20 37.361
R1115 a_20223_2963.n0 a_20223_2963.t24 37.361
R1116 a_20223_2963.n8 a_20223_2963.t40 37.361
R1117 a_20223_2963.n2 a_20223_2963.t38 37.361
R1118 a_20223_2963.n2 a_20223_2963.t16 37.361
R1119 a_20223_2963.n3 a_20223_2963.t34 37.361
R1120 a_20223_2963.n3 a_20223_2963.t22 37.361
R1121 a_20223_2963.n3 a_20223_2963.t28 37.361
R1122 a_20223_2963.n3 a_20223_2963.t42 37.361
R1123 a_20223_2963.n3 a_20223_2963.t46 37.361
R1124 a_20223_2963.n3 a_20223_2963.t32 37.361
R1125 a_20223_2963.n3 a_20223_2963.t62 37.361
R1126 a_20223_2963.n6 a_20223_2963.t59 37.361
R1127 a_20223_2963.n3 a_20223_2963.t58 37.361
R1128 a_20223_2963.n3 a_20223_2963.t50 37.361
R1129 a_20223_2963.n2 a_20223_2963.t36 37.361
R1130 a_20223_2963.n2 a_20223_2963.t49 37.361
R1131 a_20223_2963.n4 a_20223_2963.t61 37.361
R1132 a_20223_2963.n1 a_20223_2963.t60 37.361
R1133 a_20223_2963.n1 a_20223_2963.t63 37.361
R1134 a_20223_2963.n1 a_20223_2963.t18 37.361
R1135 a_20223_2963.n1 a_20223_2963.t30 37.361
R1136 a_20223_2963.n1 a_20223_2963.t29 17.43
R1137 a_20223_2963.n7 a_20223_2963.t45 17.43
R1138 a_20223_2963.n7 a_20223_2963.t27 17.43
R1139 a_20223_2963.n2 a_20223_2963.t17 17.43
R1140 a_20223_2963.n2 a_20223_2963.t39 17.43
R1141 a_20223_2963.n0 a_20223_2963.t25 17.43
R1142 a_20223_2963.n0 a_20223_2963.t41 17.43
R1143 a_20223_2963.n2 a_20223_2963.t37 17.43
R1144 a_20223_2963.n2 a_20223_2963.t21 17.43
R1145 a_20223_2963.n3 a_20223_2963.t23 17.43
R1146 a_20223_2963.n3 a_20223_2963.t35 17.43
R1147 a_20223_2963.n3 a_20223_2963.t43 17.43
R1148 a_20223_2963.n3 a_20223_2963.t33 17.43
R1149 a_20223_2963.n1 a_20223_2963.t31 17.43
R1150 a_20223_2963.n1 a_20223_2963.t19 17.43
R1151 a_20223_2963.t47 a_20223_2963.n1 17.43
R1152 a_20223_2963.n12 a_20223_2963.t12 7.146
R1153 a_20223_2963.n12 a_20223_2963.t4 7.146
R1154 a_20223_2963.n11 a_20223_2963.t11 7.146
R1155 a_20223_2963.n11 a_20223_2963.t5 7.146
R1156 a_20223_2963.n10 a_20223_2963.t8 7.146
R1157 a_20223_2963.n10 a_20223_2963.t14 7.146
R1158 a_20223_2963.n9 a_20223_2963.t13 7.146
R1159 a_20223_2963.n9 a_20223_2963.t2 7.146
R1160 a_20223_2963.n19 a_20223_2963.t10 7.146
R1161 a_20223_2963.n19 a_20223_2963.t7 7.146
R1162 a_20223_2963.n18 a_20223_2963.t0 7.146
R1163 a_20223_2963.n18 a_20223_2963.t1 7.146
R1164 a_20223_2963.n17 a_20223_2963.t6 7.146
R1165 a_20223_2963.n17 a_20223_2963.t3 7.146
R1166 a_20223_2963.n16 a_20223_2963.t9 7.146
R1167 a_20223_2963.n16 a_20223_2963.t15 7.146
R1168 a_20223_2963.n7 a_20223_2963.n12 1.777
R1169 a_20223_2963.n5 a_20223_2963.n19 1.583
R1170 a_20223_2963.n1 a_20223_2963.n0 1.406
R1171 a_20223_2963.n1 a_20223_2963.n22 1.076
R1172 a_20223_2963.n5 a_20223_2963.n15 1.048
R1173 a_20223_2963.n10 a_20223_2963.n9 1.045
R1174 a_20223_2963.n11 a_20223_2963.n10 1.045
R1175 a_20223_2963.n12 a_20223_2963.n11 1.045
R1176 a_20223_2963.n17 a_20223_2963.n16 1.045
R1177 a_20223_2963.n18 a_20223_2963.n17 1.045
R1178 a_20223_2963.n19 a_20223_2963.n18 1.045
R1179 a_20223_2963.n4 a_20223_2963.n2 1.012
R1180 a_20223_2963.n6 a_20223_2963.n7 0.878
R1181 a_20223_2963.n1 a_20223_2963.n3 0.849
R1182 a_20223_2963.n3 a_20223_2963.n6 0.841
R1183 a_20223_2963.n3 a_20223_2963.n4 0.841
R1184 a_20223_2963.n3 a_20223_2963.n5 0.696
R1185 a_20223_2963.n15 a_20223_2963.n14 0.604
R1186 a_20223_2963.n21 a_20223_2963.n20 0.603
R1187 a_20223_2963.n22 a_20223_2963.n21 0.603
R1188 a_20223_2963.n14 a_20223_2963.n13 0.603
R1189 a_20223_2963.n0 a_20223_2963.n8 0.564
R1190 w_20027_5063.n36 w_20027_5063.n35 779.876
R1191 w_20027_5063.n10 w_20027_5063.n51 60.285
R1192 w_20027_5063.n5 w_20027_5063.t26 14.295
R1193 w_20027_5063.n5 w_20027_5063.t38 14.295
R1194 w_20027_5063.n4 w_20027_5063.t21 14.295
R1195 w_20027_5063.n4 w_20027_5063.t27 14.295
R1196 w_20027_5063.n3 w_20027_5063.t36 14.295
R1197 w_20027_5063.n3 w_20027_5063.t19 14.295
R1198 w_20027_5063.n14 w_20027_5063.t28 14.295
R1199 w_20027_5063.n14 w_20027_5063.t18 14.295
R1200 w_20027_5063.n13 w_20027_5063.t39 14.295
R1201 w_20027_5063.n13 w_20027_5063.t20 14.295
R1202 w_20027_5063.n12 w_20027_5063.t32 14.295
R1203 w_20027_5063.n12 w_20027_5063.t35 14.295
R1204 w_20027_5063.n23 w_20027_5063.t41 14.295
R1205 w_20027_5063.n23 w_20027_5063.t30 14.295
R1206 w_20027_5063.n22 w_20027_5063.t31 14.295
R1207 w_20027_5063.n22 w_20027_5063.t34 14.295
R1208 w_20027_5063.n21 w_20027_5063.t23 14.295
R1209 w_20027_5063.n21 w_20027_5063.t29 14.295
R1210 w_20027_5063.n34 w_20027_5063.t24 14.295
R1211 w_20027_5063.n34 w_20027_5063.t40 14.295
R1212 w_20027_5063.n33 w_20027_5063.t22 14.295
R1213 w_20027_5063.n33 w_20027_5063.t33 14.295
R1214 w_20027_5063.n32 w_20027_5063.t25 14.295
R1215 w_20027_5063.n32 w_20027_5063.t37 14.295
R1216 w_20027_5063.n37 w_20027_5063.t7 8.834
R1217 w_20027_5063.n24 w_20027_5063.t2 8.766
R1218 w_20027_5063.n50 w_20027_5063.t42 7.146
R1219 w_20027_5063.n48 w_20027_5063.t52 7.146
R1220 w_20027_5063.n48 w_20027_5063.t10 7.146
R1221 w_20027_5063.n47 w_20027_5063.t48 7.146
R1222 w_20027_5063.n47 w_20027_5063.t3 7.146
R1223 w_20027_5063.n9 w_20027_5063.t45 7.146
R1224 w_20027_5063.n9 w_20027_5063.t51 7.146
R1225 w_20027_5063.n8 w_20027_5063.t47 7.146
R1226 w_20027_5063.n8 w_20027_5063.t54 7.146
R1227 w_20027_5063.n7 w_20027_5063.t1 7.146
R1228 w_20027_5063.n7 w_20027_5063.t49 7.146
R1229 w_20027_5063.n6 w_20027_5063.t0 7.146
R1230 w_20027_5063.n6 w_20027_5063.t55 7.146
R1231 w_20027_5063.n19 w_20027_5063.t16 7.146
R1232 w_20027_5063.n19 w_20027_5063.t44 7.146
R1233 w_20027_5063.n18 w_20027_5063.t6 7.146
R1234 w_20027_5063.n18 w_20027_5063.t46 7.146
R1235 w_20027_5063.n17 w_20027_5063.t12 7.146
R1236 w_20027_5063.n17 w_20027_5063.t43 7.146
R1237 w_20027_5063.n16 w_20027_5063.t9 7.146
R1238 w_20027_5063.n16 w_20027_5063.t50 7.146
R1239 w_20027_5063.n26 w_20027_5063.t8 7.146
R1240 w_20027_5063.n25 w_20027_5063.t15 7.146
R1241 w_20027_5063.n24 w_20027_5063.t5 7.146
R1242 w_20027_5063.n39 w_20027_5063.t14 7.146
R1243 w_20027_5063.n38 w_20027_5063.t4 7.146
R1244 w_20027_5063.n37 w_20027_5063.t11 7.146
R1245 w_20027_5063.n49 w_20027_5063.t53 7.146
R1246 w_20027_5063.n49 w_20027_5063.t13 7.146
R1247 w_20027_5063.t17 w_20027_5063.n50 7.146
R1248 w_20027_5063.n0 w_20027_5063.n36 5.228
R1249 w_20027_5063.n27 w_20027_5063.n23 2.373
R1250 w_20027_5063.n42 w_20027_5063.n34 2.373
R1251 w_20027_5063.n38 w_20027_5063.n37 1.688
R1252 w_20027_5063.n39 w_20027_5063.n38 1.688
R1253 w_20027_5063.n25 w_20027_5063.n24 1.62
R1254 w_20027_5063.n26 w_20027_5063.n25 1.62
R1255 w_20027_5063.n27 w_20027_5063.n26 1.149
R1256 w_20027_5063.n7 w_20027_5063.n6 1.045
R1257 w_20027_5063.n8 w_20027_5063.n7 1.045
R1258 w_20027_5063.n9 w_20027_5063.n8 1.045
R1259 w_20027_5063.n17 w_20027_5063.n16 1.045
R1260 w_20027_5063.n18 w_20027_5063.n17 1.045
R1261 w_20027_5063.n19 w_20027_5063.n18 1.045
R1262 w_20027_5063.n48 w_20027_5063.n47 1.045
R1263 w_20027_5063.n50 w_20027_5063.n48 1.045
R1264 w_20027_5063.n50 w_20027_5063.n49 1.045
R1265 w_20027_5063.n45 w_20027_5063.n5 0.893
R1266 w_20027_5063.n29 w_20027_5063.n14 0.893
R1267 w_20027_5063.n0 w_20027_5063.n39 0.871
R1268 w_20027_5063.n31 w_20027_5063.n30 0.748
R1269 w_20027_5063.n29 w_20027_5063.n28 0.748
R1270 w_20027_5063.n4 w_20027_5063.n3 0.733
R1271 w_20027_5063.n5 w_20027_5063.n4 0.733
R1272 w_20027_5063.n13 w_20027_5063.n12 0.733
R1273 w_20027_5063.n14 w_20027_5063.n13 0.733
R1274 w_20027_5063.n22 w_20027_5063.n21 0.733
R1275 w_20027_5063.n23 w_20027_5063.n22 0.733
R1276 w_20027_5063.n33 w_20027_5063.n32 0.733
R1277 w_20027_5063.n34 w_20027_5063.n33 0.733
R1278 w_20027_5063.n44 w_20027_5063.n42 0.72
R1279 w_20027_5063.n10 w_20027_5063.n9 0.621
R1280 w_20027_5063.n1 w_20027_5063.n19 0.621
R1281 w_20027_5063.n47 w_20027_5063.n2 0.621
R1282 w_20027_5063.n45 w_20027_5063.n31 1.316
R1283 w_20027_5063.n30 w_20027_5063.n29 0.568
R1284 w_20027_5063.n45 w_20027_5063.n44 0.568
R1285 w_20027_5063.n28 w_20027_5063.n27 0.541
R1286 w_20027_5063.n44 w_20027_5063.n43 0.491
R1287 w_20027_5063.n28 w_20027_5063.n20 0.491
R1288 w_20027_5063.n30 w_20027_5063.n11 0.491
R1289 w_20027_5063.n42 w_20027_5063.n0 0.288
R1290 w_20027_5063.n0 w_20027_5063.n41 0.28
R1291 w_20027_5063.n41 w_20027_5063.n40 0.28
R1292 w_20027_5063.n29 w_20027_5063.n1 0.267
R1293 w_20027_5063.n31 w_20027_5063.n10 0.267
R1294 w_20027_5063.n2 w_20027_5063.n45 0.267
R1295 w_20027_5063.n2 w_20027_5063.n46 0.196
R1296 w_20027_5063.n1 w_20027_5063.n15 0.196
R1297 vp.n0 vp.t1 111.996
R1298 vp.n25 vp.t9 111.994
R1299 vp.n6 vp.t10 111.83
R1300 vp.n10 vp.t4 111.83
R1301 vp.n21 vp.t13 111.83
R1302 vp.n1 vp.t0 111.83
R1303 vp.n15 vp.t11 111.83
R1304 vp.n17 vp.t5 111.83
R1305 vp.n19 vp.t14 111.83
R1306 vp.n8 vp.t3 111.83
R1307 vp.n12 vp.t12 111.83
R1308 vp.n23 vp.t7 111.83
R1309 vp.n2 vp.t6 111.83
R1310 vp.n22 vp.t2 111.83
R1311 vp.n11 vp.t8 111.83
R1312 vp.n7 vp.t15 111.83
R1313 vp.n25 vp.n24 2.022
R1314 vp.n18 vp.n16 2.018
R1315 vp.n13 vp.n9 2.018
R1316 vp.n24 vp.n13 2.018
R1317 vp.n20 vp.n18 2.018
R1318 vp.n9 vp.n5 1.986
R1319 vp.n16 vp.n14 1.986
R1320 vp vp.n26 1.714
R1321 vp.n26 vp.n0 0.868
R1322 vp.n2 vp.n1 0.619
R1323 vp.n4 vp.n3 0.547
R1324 vp.n7 vp.n6 0.281
R1325 vp.n11 vp.n10 0.281
R1326 vp.n22 vp.n21 0.281
R1327 vp.n5 vp.n4 0.273
R1328 vp.n25 vp.n2 0.167
R1329 vp.n21 vp.n20 0.14
R1330 vp.n24 vp.n23 0.14
R1331 vp.n13 vp.n12 0.14
R1332 vp.n9 vp.n8 0.14
R1333 vp.n16 vp.n15 0.139
R1334 vp.n18 vp.n17 0.139
R1335 vp.n20 vp.n19 0.139
R1336 vp.n24 vp.n22 0.139
R1337 vp.n13 vp.n11 0.139
R1338 vp.n9 vp.n7 0.139
R1339 vp.n26 vp.n25 0.136
C5 vp vss 7.41fF
C6 vn vss 6.69fF
C7 vout vss 53.03fF
C8 vbias vss 43.40fF
C9 vdd vss 123.73fF
C10 a_23819_6897# vss 1.85fF
C11 w_20027_5063.n3 vss 1.58fF $ **FLOATING
C12 w_20027_5063.n4 vss 1.68fF $ **FLOATING
C13 w_20027_5063.n5 vss 1.65fF $ **FLOATING
C14 w_20027_5063.n6 vss 3.06fF $ **FLOATING
C15 w_20027_5063.n7 vss 3.16fF $ **FLOATING
C16 w_20027_5063.n8 vss 3.16fF $ **FLOATING
C17 w_20027_5063.n9 vss 2.90fF $ **FLOATING
C18 w_20027_5063.n12 vss 1.58fF $ **FLOATING
C19 w_20027_5063.n13 vss 1.68fF $ **FLOATING
C20 w_20027_5063.n14 vss 1.65fF $ **FLOATING
C21 w_20027_5063.n16 vss 3.06fF $ **FLOATING
C22 w_20027_5063.n17 vss 3.16fF $ **FLOATING
C23 w_20027_5063.n18 vss 3.16fF $ **FLOATING
C24 w_20027_5063.n19 vss 2.90fF $ **FLOATING
C25 w_20027_5063.n21 vss 1.58fF $ **FLOATING
C26 w_20027_5063.n22 vss 1.68fF $ **FLOATING
C27 w_20027_5063.n23 vss 1.94fF $ **FLOATING
C28 w_20027_5063.n24 vss 3.12fF $ **FLOATING
C29 w_20027_5063.n25 vss 1.76fF $ **FLOATING
C30 w_20027_5063.n26 vss 2.61fF $ **FLOATING
C31 w_20027_5063.n27 vss 3.82fF $ **FLOATING
C32 w_20027_5063.n32 vss 1.58fF $ **FLOATING
C33 w_20027_5063.n33 vss 1.68fF $ **FLOATING
C34 w_20027_5063.n34 vss 1.94fF $ **FLOATING
C35 w_20027_5063.n35 vss 4.69fF $ **FLOATING
C36 w_20027_5063.n37 vss 3.09fF $ **FLOATING
C37 w_20027_5063.n38 vss 1.74fF $ **FLOATING
C38 w_20027_5063.n39 vss 1.56fF $ **FLOATING
C39 w_20027_5063.n47 vss 2.90fF $ **FLOATING
C40 w_20027_5063.n48 vss 3.16fF $ **FLOATING
C41 w_20027_5063.n49 vss 3.06fF $ **FLOATING
C42 w_20027_5063.n50 vss 3.16fF $ **FLOATING
C43 a_20223_2963.n0 vss 3.31fF $ **FLOATING
C44 a_20223_2963.n1 vss 5.30fF $ **FLOATING
C45 a_20223_2963.n2 vss 3.15fF $ **FLOATING
C46 a_20223_2963.n3 vss 5.70fF $ **FLOATING
C47 a_20223_2963.n4 vss 1.60fF $ **FLOATING
C48 a_20223_2963.n6 vss 1.60fF $ **FLOATING
C49 a_20223_2963.n7 vss 4.07fF $ **FLOATING
C50 a_20223_2963.n9 vss 1.41fF $ **FLOATING
C51 a_20223_2963.n10 vss 1.46fF $ **FLOATING
C52 a_20223_2963.n11 vss 1.46fF $ **FLOATING
C53 a_20223_2963.n12 vss 1.63fF $ **FLOATING
C54 a_20223_2963.n16 vss 1.41fF $ **FLOATING
C55 a_20223_2963.n17 vss 1.46fF $ **FLOATING
C56 a_20223_2963.n18 vss 1.46fF $ **FLOATING
C57 a_20223_2963.n19 vss 1.49fF $ **FLOATING
C58 vn.n10 vss 1.27fF $ **FLOATING
C59 a_21167_3051.n0 vss 1.49fF $ **FLOATING
C60 a_21167_3051.n1 vss 6.75fF $ **FLOATING
C61 a_21167_3051.n2 vss 7.51fF $ **FLOATING
C62 a_21167_3051.n3 vss 3.02fF $ **FLOATING
C63 a_21167_3051.n4 vss 33.49fF $ **FLOATING
C64 a_21167_3051.n5 vss 10.89fF $ **FLOATING
C65 a_21167_3051.n7 vss 4.13fF $ **FLOATING
C66 a_21167_3051.n8 vss 3.03fF $ **FLOATING
C67 a_21167_3051.n9 vss 3.24fF $ **FLOATING
C68 vdd.n114 vss 1.05fF $ **FLOATING
C69 vdd.n117 vss 3.91fF $ **FLOATING
C70 vdd.n125 vss 10.94fF $ **FLOATING
C71 vdd.n126 vss 6.13fF $ **FLOATING
C72 vdd.n127 vss 6.13fF $ **FLOATING
C73 vdd.n128 vss 6.13fF $ **FLOATING
C74 vdd.n129 vss 6.13fF $ **FLOATING
C75 vdd.n130 vss 6.13fF $ **FLOATING
C76 vdd.n131 vss 6.13fF $ **FLOATING
C77 vdd.n132 vss 4.83fF $ **FLOATING
C78 vdd.n133 vss 4.84fF $ **FLOATING
C79 vdd.n134 vss 6.13fF $ **FLOATING
C80 vdd.n135 vss 6.13fF $ **FLOATING
C81 vdd.n136 vss 6.13fF $ **FLOATING
C82 vdd.n137 vss 6.13fF $ **FLOATING
C83 vdd.n138 vss 6.13fF $ **FLOATING
C84 vdd.n139 vss 4.42fF $ **FLOATING
C85 vdd.n140 vss 3.68fF $ **FLOATING
C86 vout.n8 vss 1.11fF $ **FLOATING
C87 vout.n9 vss 2.66fF $ **FLOATING
C88 vout.n10 vss 2.18fF $ **FLOATING
C89 vout.n14 vss 2.18fF $ **FLOATING
C90 vout.n18 vss 2.18fF $ **FLOATING
C91 vout.n24 vss 1.11fF $ **FLOATING
C92 vout.n25 vss 2.66fF $ **FLOATING
C93 vout.n29 vss 2.18fF $ **FLOATING
C94 vout.n50 vss 2.24fF $ **FLOATING
C95 vout.n51 vss 1.40fF $ **FLOATING
C96 vout.n52 vss 1.40fF $ **FLOATING
C97 vout.n53 vss 2.30fF $ **FLOATING
C98 vout.n54 vss 38.33fF $ **FLOATING
C99 vout.n59 vss 2.30fF $ **FLOATING
C100 vout.n60 vss 12.77fF $ **FLOATING
C101 vout.n65 vss 2.30fF $ **FLOATING
C102 vout.n66 vss 12.77fF $ **FLOATING
C103 vout.n71 vss 2.07fF $ **FLOATING
C104 vout.n72 vss 32.48fF $ **FLOATING
.ends
