magic
tech sky130A
magscale 1 2
timestamp 1627023135
<< nwell >>
rect 10118 7780 39138 11644
rect 23130 3240 26126 7270
<< pwell >>
rect 19422 13108 29836 15744
rect 30615 3569 31017 5325
rect 23742 462 25516 3078
<< pmoslvt >>
rect 10610 10312 11010 11112
rect 11198 10312 11598 11112
rect 11786 10312 12186 11112
rect 12374 10312 12774 11112
rect 12962 10312 13362 11112
rect 13550 10312 13950 11112
rect 14138 10312 14538 11112
rect 14726 10312 15126 11112
rect 15314 10312 15714 11112
rect 15902 10312 16302 11112
rect 16490 10312 16890 11112
rect 17078 10312 17478 11112
rect 17666 10312 18066 11112
rect 18254 10312 18654 11112
rect 18842 10312 19242 11112
rect 19430 10312 19830 11112
rect 20018 10312 20418 11112
rect 20606 10312 21006 11112
rect 21194 10312 21594 11112
rect 21782 10312 22182 11112
rect 22370 10312 22770 11112
rect 22958 10312 23358 11112
rect 23546 10312 23946 11112
rect 24134 10312 24534 11112
rect 24722 10312 25122 11112
rect 25310 10312 25710 11112
rect 25898 10312 26298 11112
rect 26486 10312 26886 11112
rect 27074 10312 27474 11112
rect 27662 10312 28062 11112
rect 28250 10312 28650 11112
rect 28838 10312 29238 11112
rect 29426 10312 29826 11112
rect 30014 10312 30414 11112
rect 30602 10312 31002 11112
rect 31190 10312 31590 11112
rect 31778 10312 32178 11112
rect 32366 10312 32766 11112
rect 32954 10312 33354 11112
rect 33542 10312 33942 11112
rect 34130 10312 34530 11112
rect 34718 10312 35118 11112
rect 35306 10312 35706 11112
rect 35894 10312 36294 11112
rect 36482 10312 36882 11112
rect 37070 10312 37470 11112
rect 37658 10312 38058 11112
rect 38246 10312 38646 11112
rect 10610 9312 11010 10112
rect 11198 9312 11598 10112
rect 11786 9312 12186 10112
rect 12374 9312 12774 10112
rect 12962 9312 13362 10112
rect 13550 9312 13950 10112
rect 14138 9312 14538 10112
rect 14726 9312 15126 10112
rect 15314 9312 15714 10112
rect 15902 9312 16302 10112
rect 16490 9312 16890 10112
rect 17078 9312 17478 10112
rect 17666 9312 18066 10112
rect 18254 9312 18654 10112
rect 18842 9312 19242 10112
rect 19430 9312 19830 10112
rect 20018 9312 20418 10112
rect 20606 9312 21006 10112
rect 21194 9312 21594 10112
rect 21782 9312 22182 10112
rect 22370 9312 22770 10112
rect 22958 9312 23358 10112
rect 23546 9312 23946 10112
rect 24134 9312 24534 10112
rect 24722 9312 25122 10112
rect 25310 9312 25710 10112
rect 25898 9312 26298 10112
rect 26486 9312 26886 10112
rect 27074 9312 27474 10112
rect 27662 9312 28062 10112
rect 28250 9312 28650 10112
rect 28838 9312 29238 10112
rect 29426 9312 29826 10112
rect 30014 9312 30414 10112
rect 30602 9312 31002 10112
rect 31190 9312 31590 10112
rect 31778 9312 32178 10112
rect 32366 9312 32766 10112
rect 32954 9312 33354 10112
rect 33542 9312 33942 10112
rect 34130 9312 34530 10112
rect 34718 9312 35118 10112
rect 35306 9312 35706 10112
rect 35894 9312 36294 10112
rect 36482 9312 36882 10112
rect 37070 9312 37470 10112
rect 37658 9312 38058 10112
rect 38246 9312 38646 10112
rect 10610 8312 11010 9112
rect 11198 8312 11598 9112
rect 11786 8312 12186 9112
rect 12374 8312 12774 9112
rect 12962 8312 13362 9112
rect 13550 8312 13950 9112
rect 14138 8312 14538 9112
rect 14726 8312 15126 9112
rect 15314 8312 15714 9112
rect 15902 8312 16302 9112
rect 16490 8312 16890 9112
rect 17078 8312 17478 9112
rect 17666 8312 18066 9112
rect 18254 8312 18654 9112
rect 18842 8312 19242 9112
rect 19430 8312 19830 9112
rect 20018 8312 20418 9112
rect 20606 8312 21006 9112
rect 21194 8312 21594 9112
rect 21782 8312 22182 9112
rect 22370 8312 22770 9112
rect 22958 8312 23358 9112
rect 23546 8312 23946 9112
rect 24134 8312 24534 9112
rect 24722 8312 25122 9112
rect 25310 8312 25710 9112
rect 25898 8312 26298 9112
rect 26486 8312 26886 9112
rect 27074 8312 27474 9112
rect 27662 8312 28062 9112
rect 28250 8312 28650 9112
rect 28838 8312 29238 9112
rect 29426 8312 29826 9112
rect 30014 8312 30414 9112
rect 30602 8312 31002 9112
rect 31190 8312 31590 9112
rect 31778 8312 32178 9112
rect 32366 8312 32766 9112
rect 32954 8312 33354 9112
rect 33542 8312 33942 9112
rect 34130 8312 34530 9112
rect 34718 8312 35118 9112
rect 35306 8312 35706 9112
rect 35894 8312 36294 9112
rect 36482 8312 36882 9112
rect 37070 8312 37470 9112
rect 37658 8312 38058 9112
rect 38246 8312 38646 9112
rect 23662 5866 23732 6666
rect 23928 5866 23998 6666
rect 24194 5866 24264 6666
rect 24460 5866 24530 6666
rect 24726 5866 24796 6666
rect 24992 5866 25062 6666
rect 25258 5866 25328 6666
rect 25524 5866 25594 6666
rect 23662 4856 23732 5656
rect 23928 4856 23998 5656
rect 24194 4856 24264 5656
rect 24460 4856 24530 5656
rect 24726 4856 24796 5656
rect 24992 4856 25062 5656
rect 25258 4856 25328 5656
rect 25524 4856 25594 5656
rect 23662 3846 23732 4646
rect 23928 3846 23998 4646
rect 24194 3846 24264 4646
rect 24460 3846 24530 4646
rect 24726 3846 24796 4646
rect 24992 3846 25062 4646
rect 25258 3846 25328 4646
rect 25524 3846 25594 4646
<< nmoslvt >>
rect 19914 14530 19984 15130
rect 20154 14530 20224 15130
rect 20394 14530 20464 15130
rect 20634 14530 20704 15130
rect 20874 14530 20944 15130
rect 21114 14530 21184 15130
rect 21354 14530 21424 15130
rect 21594 14530 21664 15130
rect 21834 14530 21904 15130
rect 22074 14530 22144 15130
rect 22314 14530 22384 15130
rect 22554 14530 22624 15130
rect 22794 14530 22864 15130
rect 23034 14530 23104 15130
rect 23274 14530 23344 15130
rect 23514 14530 23584 15130
rect 23754 14530 23824 15130
rect 23994 14530 24064 15130
rect 24234 14530 24304 15130
rect 24474 14530 24544 15130
rect 24714 14530 24784 15130
rect 24954 14530 25024 15130
rect 25194 14530 25264 15130
rect 25434 14530 25504 15130
rect 25674 14530 25744 15130
rect 25914 14530 25984 15130
rect 26154 14530 26224 15130
rect 26394 14530 26464 15130
rect 26634 14530 26704 15130
rect 26874 14530 26944 15130
rect 27114 14530 27184 15130
rect 27354 14530 27424 15130
rect 27594 14530 27664 15130
rect 27834 14530 27904 15130
rect 28074 14530 28144 15130
rect 28314 14530 28384 15130
rect 28554 14530 28624 15130
rect 28794 14530 28864 15130
rect 29034 14530 29104 15130
rect 29274 14530 29344 15130
rect 19914 13722 19984 14322
rect 20154 13722 20224 14322
rect 20394 13722 20464 14322
rect 20634 13722 20704 14322
rect 20874 13722 20944 14322
rect 21114 13722 21184 14322
rect 21354 13722 21424 14322
rect 21594 13722 21664 14322
rect 21834 13722 21904 14322
rect 22074 13722 22144 14322
rect 22314 13722 22384 14322
rect 22554 13722 22624 14322
rect 22794 13722 22864 14322
rect 23034 13722 23104 14322
rect 23274 13722 23344 14322
rect 23514 13722 23584 14322
rect 23754 13722 23824 14322
rect 23994 13722 24064 14322
rect 24234 13722 24304 14322
rect 24474 13722 24544 14322
rect 24714 13722 24784 14322
rect 24954 13722 25024 14322
rect 25194 13722 25264 14322
rect 25434 13722 25504 14322
rect 25674 13722 25744 14322
rect 25914 13722 25984 14322
rect 26154 13722 26224 14322
rect 26394 13722 26464 14322
rect 26634 13722 26704 14322
rect 26874 13722 26944 14322
rect 27114 13722 27184 14322
rect 27354 13722 27424 14322
rect 27594 13722 27664 14322
rect 27834 13722 27904 14322
rect 28074 13722 28144 14322
rect 28314 13722 28384 14322
rect 28554 13722 28624 14322
rect 28794 13722 28864 14322
rect 29034 13722 29104 14322
rect 29274 13722 29344 14322
rect 24234 1874 24304 2474
rect 24474 1874 24544 2474
rect 24714 1874 24784 2474
rect 24954 1874 25024 2474
rect 24234 1066 24304 1666
rect 24474 1066 24544 1666
rect 24714 1066 24784 1666
rect 24954 1066 25024 1666
<< ndiff >>
rect 19856 15118 19914 15130
rect 19856 14542 19868 15118
rect 19902 14542 19914 15118
rect 19856 14530 19914 14542
rect 19984 15118 20042 15130
rect 19984 14542 19996 15118
rect 20030 14542 20042 15118
rect 19984 14530 20042 14542
rect 20096 15118 20154 15130
rect 20096 14542 20108 15118
rect 20142 14542 20154 15118
rect 20096 14530 20154 14542
rect 20224 15118 20282 15130
rect 20224 14542 20236 15118
rect 20270 14542 20282 15118
rect 20224 14530 20282 14542
rect 20336 15118 20394 15130
rect 20336 14542 20348 15118
rect 20382 14542 20394 15118
rect 20336 14530 20394 14542
rect 20464 15118 20522 15130
rect 20464 14542 20476 15118
rect 20510 14542 20522 15118
rect 20464 14530 20522 14542
rect 20576 15118 20634 15130
rect 20576 14542 20588 15118
rect 20622 14542 20634 15118
rect 20576 14530 20634 14542
rect 20704 15118 20762 15130
rect 20704 14542 20716 15118
rect 20750 14542 20762 15118
rect 20704 14530 20762 14542
rect 20816 15118 20874 15130
rect 20816 14542 20828 15118
rect 20862 14542 20874 15118
rect 20816 14530 20874 14542
rect 20944 15118 21002 15130
rect 20944 14542 20956 15118
rect 20990 14542 21002 15118
rect 20944 14530 21002 14542
rect 21056 15118 21114 15130
rect 21056 14542 21068 15118
rect 21102 14542 21114 15118
rect 21056 14530 21114 14542
rect 21184 15118 21242 15130
rect 21184 14542 21196 15118
rect 21230 14542 21242 15118
rect 21184 14530 21242 14542
rect 21296 15118 21354 15130
rect 21296 14542 21308 15118
rect 21342 14542 21354 15118
rect 21296 14530 21354 14542
rect 21424 15118 21482 15130
rect 21424 14542 21436 15118
rect 21470 14542 21482 15118
rect 21424 14530 21482 14542
rect 21536 15118 21594 15130
rect 21536 14542 21548 15118
rect 21582 14542 21594 15118
rect 21536 14530 21594 14542
rect 21664 15118 21722 15130
rect 21664 14542 21676 15118
rect 21710 14542 21722 15118
rect 21664 14530 21722 14542
rect 21776 15118 21834 15130
rect 21776 14542 21788 15118
rect 21822 14542 21834 15118
rect 21776 14530 21834 14542
rect 21904 15118 21962 15130
rect 21904 14542 21916 15118
rect 21950 14542 21962 15118
rect 21904 14530 21962 14542
rect 22016 15118 22074 15130
rect 22016 14542 22028 15118
rect 22062 14542 22074 15118
rect 22016 14530 22074 14542
rect 22144 15118 22202 15130
rect 22144 14542 22156 15118
rect 22190 14542 22202 15118
rect 22144 14530 22202 14542
rect 22256 15118 22314 15130
rect 22256 14542 22268 15118
rect 22302 14542 22314 15118
rect 22256 14530 22314 14542
rect 22384 15118 22442 15130
rect 22384 14542 22396 15118
rect 22430 14542 22442 15118
rect 22384 14530 22442 14542
rect 22496 15118 22554 15130
rect 22496 14542 22508 15118
rect 22542 14542 22554 15118
rect 22496 14530 22554 14542
rect 22624 15118 22682 15130
rect 22624 14542 22636 15118
rect 22670 14542 22682 15118
rect 22624 14530 22682 14542
rect 22736 15118 22794 15130
rect 22736 14542 22748 15118
rect 22782 14542 22794 15118
rect 22736 14530 22794 14542
rect 22864 15118 22922 15130
rect 22864 14542 22876 15118
rect 22910 14542 22922 15118
rect 22864 14530 22922 14542
rect 22976 15118 23034 15130
rect 22976 14542 22988 15118
rect 23022 14542 23034 15118
rect 22976 14530 23034 14542
rect 23104 15118 23162 15130
rect 23104 14542 23116 15118
rect 23150 14542 23162 15118
rect 23104 14530 23162 14542
rect 23216 15118 23274 15130
rect 23216 14542 23228 15118
rect 23262 14542 23274 15118
rect 23216 14530 23274 14542
rect 23344 15118 23402 15130
rect 23344 14542 23356 15118
rect 23390 14542 23402 15118
rect 23344 14530 23402 14542
rect 23456 15118 23514 15130
rect 23456 14542 23468 15118
rect 23502 14542 23514 15118
rect 23456 14530 23514 14542
rect 23584 15118 23642 15130
rect 23584 14542 23596 15118
rect 23630 14542 23642 15118
rect 23584 14530 23642 14542
rect 23696 15118 23754 15130
rect 23696 14542 23708 15118
rect 23742 14542 23754 15118
rect 23696 14530 23754 14542
rect 23824 15118 23882 15130
rect 23824 14542 23836 15118
rect 23870 14542 23882 15118
rect 23824 14530 23882 14542
rect 23936 15118 23994 15130
rect 23936 14542 23948 15118
rect 23982 14542 23994 15118
rect 23936 14530 23994 14542
rect 24064 15118 24122 15130
rect 24064 14542 24076 15118
rect 24110 14542 24122 15118
rect 24064 14530 24122 14542
rect 24176 15118 24234 15130
rect 24176 14542 24188 15118
rect 24222 14542 24234 15118
rect 24176 14530 24234 14542
rect 24304 15118 24362 15130
rect 24304 14542 24316 15118
rect 24350 14542 24362 15118
rect 24304 14530 24362 14542
rect 24416 15118 24474 15130
rect 24416 14542 24428 15118
rect 24462 14542 24474 15118
rect 24416 14530 24474 14542
rect 24544 15118 24602 15130
rect 24544 14542 24556 15118
rect 24590 14542 24602 15118
rect 24544 14530 24602 14542
rect 24656 15118 24714 15130
rect 24656 14542 24668 15118
rect 24702 14542 24714 15118
rect 24656 14530 24714 14542
rect 24784 15118 24842 15130
rect 24784 14542 24796 15118
rect 24830 14542 24842 15118
rect 24784 14530 24842 14542
rect 24896 15118 24954 15130
rect 24896 14542 24908 15118
rect 24942 14542 24954 15118
rect 24896 14530 24954 14542
rect 25024 15118 25082 15130
rect 25024 14542 25036 15118
rect 25070 14542 25082 15118
rect 25024 14530 25082 14542
rect 25136 15118 25194 15130
rect 25136 14542 25148 15118
rect 25182 14542 25194 15118
rect 25136 14530 25194 14542
rect 25264 15118 25322 15130
rect 25264 14542 25276 15118
rect 25310 14542 25322 15118
rect 25264 14530 25322 14542
rect 25376 15118 25434 15130
rect 25376 14542 25388 15118
rect 25422 14542 25434 15118
rect 25376 14530 25434 14542
rect 25504 15118 25562 15130
rect 25504 14542 25516 15118
rect 25550 14542 25562 15118
rect 25504 14530 25562 14542
rect 25616 15118 25674 15130
rect 25616 14542 25628 15118
rect 25662 14542 25674 15118
rect 25616 14530 25674 14542
rect 25744 15118 25802 15130
rect 25744 14542 25756 15118
rect 25790 14542 25802 15118
rect 25744 14530 25802 14542
rect 25856 15118 25914 15130
rect 25856 14542 25868 15118
rect 25902 14542 25914 15118
rect 25856 14530 25914 14542
rect 25984 15118 26042 15130
rect 25984 14542 25996 15118
rect 26030 14542 26042 15118
rect 25984 14530 26042 14542
rect 26096 15118 26154 15130
rect 26096 14542 26108 15118
rect 26142 14542 26154 15118
rect 26096 14530 26154 14542
rect 26224 15118 26282 15130
rect 26224 14542 26236 15118
rect 26270 14542 26282 15118
rect 26224 14530 26282 14542
rect 26336 15118 26394 15130
rect 26336 14542 26348 15118
rect 26382 14542 26394 15118
rect 26336 14530 26394 14542
rect 26464 15118 26522 15130
rect 26464 14542 26476 15118
rect 26510 14542 26522 15118
rect 26464 14530 26522 14542
rect 26576 15118 26634 15130
rect 26576 14542 26588 15118
rect 26622 14542 26634 15118
rect 26576 14530 26634 14542
rect 26704 15118 26762 15130
rect 26704 14542 26716 15118
rect 26750 14542 26762 15118
rect 26704 14530 26762 14542
rect 26816 15118 26874 15130
rect 26816 14542 26828 15118
rect 26862 14542 26874 15118
rect 26816 14530 26874 14542
rect 26944 15118 27002 15130
rect 26944 14542 26956 15118
rect 26990 14542 27002 15118
rect 26944 14530 27002 14542
rect 27056 15118 27114 15130
rect 27056 14542 27068 15118
rect 27102 14542 27114 15118
rect 27056 14530 27114 14542
rect 27184 15118 27242 15130
rect 27184 14542 27196 15118
rect 27230 14542 27242 15118
rect 27184 14530 27242 14542
rect 27296 15118 27354 15130
rect 27296 14542 27308 15118
rect 27342 14542 27354 15118
rect 27296 14530 27354 14542
rect 27424 15118 27482 15130
rect 27424 14542 27436 15118
rect 27470 14542 27482 15118
rect 27424 14530 27482 14542
rect 27536 15118 27594 15130
rect 27536 14542 27548 15118
rect 27582 14542 27594 15118
rect 27536 14530 27594 14542
rect 27664 15118 27722 15130
rect 27664 14542 27676 15118
rect 27710 14542 27722 15118
rect 27664 14530 27722 14542
rect 27776 15118 27834 15130
rect 27776 14542 27788 15118
rect 27822 14542 27834 15118
rect 27776 14530 27834 14542
rect 27904 15118 27962 15130
rect 27904 14542 27916 15118
rect 27950 14542 27962 15118
rect 27904 14530 27962 14542
rect 28016 15118 28074 15130
rect 28016 14542 28028 15118
rect 28062 14542 28074 15118
rect 28016 14530 28074 14542
rect 28144 15118 28202 15130
rect 28144 14542 28156 15118
rect 28190 14542 28202 15118
rect 28144 14530 28202 14542
rect 28256 15118 28314 15130
rect 28256 14542 28268 15118
rect 28302 14542 28314 15118
rect 28256 14530 28314 14542
rect 28384 15118 28442 15130
rect 28384 14542 28396 15118
rect 28430 14542 28442 15118
rect 28384 14530 28442 14542
rect 28496 15118 28554 15130
rect 28496 14542 28508 15118
rect 28542 14542 28554 15118
rect 28496 14530 28554 14542
rect 28624 15118 28682 15130
rect 28624 14542 28636 15118
rect 28670 14542 28682 15118
rect 28624 14530 28682 14542
rect 28736 15118 28794 15130
rect 28736 14542 28748 15118
rect 28782 14542 28794 15118
rect 28736 14530 28794 14542
rect 28864 15118 28922 15130
rect 28864 14542 28876 15118
rect 28910 14542 28922 15118
rect 28864 14530 28922 14542
rect 28976 15118 29034 15130
rect 28976 14542 28988 15118
rect 29022 14542 29034 15118
rect 28976 14530 29034 14542
rect 29104 15118 29162 15130
rect 29104 14542 29116 15118
rect 29150 14542 29162 15118
rect 29104 14530 29162 14542
rect 29216 15118 29274 15130
rect 29216 14542 29228 15118
rect 29262 14542 29274 15118
rect 29216 14530 29274 14542
rect 29344 15118 29402 15130
rect 29344 14542 29356 15118
rect 29390 14542 29402 15118
rect 29344 14530 29402 14542
rect 19856 14310 19914 14322
rect 19856 13734 19868 14310
rect 19902 13734 19914 14310
rect 19856 13722 19914 13734
rect 19984 14310 20042 14322
rect 19984 13734 19996 14310
rect 20030 13734 20042 14310
rect 19984 13722 20042 13734
rect 20096 14310 20154 14322
rect 20096 13734 20108 14310
rect 20142 13734 20154 14310
rect 20096 13722 20154 13734
rect 20224 14310 20282 14322
rect 20224 13734 20236 14310
rect 20270 13734 20282 14310
rect 20224 13722 20282 13734
rect 20336 14310 20394 14322
rect 20336 13734 20348 14310
rect 20382 13734 20394 14310
rect 20336 13722 20394 13734
rect 20464 14310 20522 14322
rect 20464 13734 20476 14310
rect 20510 13734 20522 14310
rect 20464 13722 20522 13734
rect 20576 14310 20634 14322
rect 20576 13734 20588 14310
rect 20622 13734 20634 14310
rect 20576 13722 20634 13734
rect 20704 14310 20762 14322
rect 20704 13734 20716 14310
rect 20750 13734 20762 14310
rect 20704 13722 20762 13734
rect 20816 14310 20874 14322
rect 20816 13734 20828 14310
rect 20862 13734 20874 14310
rect 20816 13722 20874 13734
rect 20944 14310 21002 14322
rect 20944 13734 20956 14310
rect 20990 13734 21002 14310
rect 20944 13722 21002 13734
rect 21056 14310 21114 14322
rect 21056 13734 21068 14310
rect 21102 13734 21114 14310
rect 21056 13722 21114 13734
rect 21184 14310 21242 14322
rect 21184 13734 21196 14310
rect 21230 13734 21242 14310
rect 21184 13722 21242 13734
rect 21296 14310 21354 14322
rect 21296 13734 21308 14310
rect 21342 13734 21354 14310
rect 21296 13722 21354 13734
rect 21424 14310 21482 14322
rect 21424 13734 21436 14310
rect 21470 13734 21482 14310
rect 21424 13722 21482 13734
rect 21536 14310 21594 14322
rect 21536 13734 21548 14310
rect 21582 13734 21594 14310
rect 21536 13722 21594 13734
rect 21664 14310 21722 14322
rect 21664 13734 21676 14310
rect 21710 13734 21722 14310
rect 21664 13722 21722 13734
rect 21776 14310 21834 14322
rect 21776 13734 21788 14310
rect 21822 13734 21834 14310
rect 21776 13722 21834 13734
rect 21904 14310 21962 14322
rect 21904 13734 21916 14310
rect 21950 13734 21962 14310
rect 21904 13722 21962 13734
rect 22016 14310 22074 14322
rect 22016 13734 22028 14310
rect 22062 13734 22074 14310
rect 22016 13722 22074 13734
rect 22144 14310 22202 14322
rect 22144 13734 22156 14310
rect 22190 13734 22202 14310
rect 22144 13722 22202 13734
rect 22256 14310 22314 14322
rect 22256 13734 22268 14310
rect 22302 13734 22314 14310
rect 22256 13722 22314 13734
rect 22384 14310 22442 14322
rect 22384 13734 22396 14310
rect 22430 13734 22442 14310
rect 22384 13722 22442 13734
rect 22496 14310 22554 14322
rect 22496 13734 22508 14310
rect 22542 13734 22554 14310
rect 22496 13722 22554 13734
rect 22624 14310 22682 14322
rect 22624 13734 22636 14310
rect 22670 13734 22682 14310
rect 22624 13722 22682 13734
rect 22736 14310 22794 14322
rect 22736 13734 22748 14310
rect 22782 13734 22794 14310
rect 22736 13722 22794 13734
rect 22864 14310 22922 14322
rect 22864 13734 22876 14310
rect 22910 13734 22922 14310
rect 22864 13722 22922 13734
rect 22976 14310 23034 14322
rect 22976 13734 22988 14310
rect 23022 13734 23034 14310
rect 22976 13722 23034 13734
rect 23104 14310 23162 14322
rect 23104 13734 23116 14310
rect 23150 13734 23162 14310
rect 23104 13722 23162 13734
rect 23216 14310 23274 14322
rect 23216 13734 23228 14310
rect 23262 13734 23274 14310
rect 23216 13722 23274 13734
rect 23344 14310 23402 14322
rect 23344 13734 23356 14310
rect 23390 13734 23402 14310
rect 23344 13722 23402 13734
rect 23456 14310 23514 14322
rect 23456 13734 23468 14310
rect 23502 13734 23514 14310
rect 23456 13722 23514 13734
rect 23584 14310 23642 14322
rect 23584 13734 23596 14310
rect 23630 13734 23642 14310
rect 23584 13722 23642 13734
rect 23696 14310 23754 14322
rect 23696 13734 23708 14310
rect 23742 13734 23754 14310
rect 23696 13722 23754 13734
rect 23824 14310 23882 14322
rect 23824 13734 23836 14310
rect 23870 13734 23882 14310
rect 23824 13722 23882 13734
rect 23936 14310 23994 14322
rect 23936 13734 23948 14310
rect 23982 13734 23994 14310
rect 23936 13722 23994 13734
rect 24064 14310 24122 14322
rect 24064 13734 24076 14310
rect 24110 13734 24122 14310
rect 24064 13722 24122 13734
rect 24176 14310 24234 14322
rect 24176 13734 24188 14310
rect 24222 13734 24234 14310
rect 24176 13722 24234 13734
rect 24304 14310 24362 14322
rect 24304 13734 24316 14310
rect 24350 13734 24362 14310
rect 24304 13722 24362 13734
rect 24416 14310 24474 14322
rect 24416 13734 24428 14310
rect 24462 13734 24474 14310
rect 24416 13722 24474 13734
rect 24544 14310 24602 14322
rect 24544 13734 24556 14310
rect 24590 13734 24602 14310
rect 24544 13722 24602 13734
rect 24656 14310 24714 14322
rect 24656 13734 24668 14310
rect 24702 13734 24714 14310
rect 24656 13722 24714 13734
rect 24784 14310 24842 14322
rect 24784 13734 24796 14310
rect 24830 13734 24842 14310
rect 24784 13722 24842 13734
rect 24896 14310 24954 14322
rect 24896 13734 24908 14310
rect 24942 13734 24954 14310
rect 24896 13722 24954 13734
rect 25024 14310 25082 14322
rect 25024 13734 25036 14310
rect 25070 13734 25082 14310
rect 25024 13722 25082 13734
rect 25136 14310 25194 14322
rect 25136 13734 25148 14310
rect 25182 13734 25194 14310
rect 25136 13722 25194 13734
rect 25264 14310 25322 14322
rect 25264 13734 25276 14310
rect 25310 13734 25322 14310
rect 25264 13722 25322 13734
rect 25376 14310 25434 14322
rect 25376 13734 25388 14310
rect 25422 13734 25434 14310
rect 25376 13722 25434 13734
rect 25504 14310 25562 14322
rect 25504 13734 25516 14310
rect 25550 13734 25562 14310
rect 25504 13722 25562 13734
rect 25616 14310 25674 14322
rect 25616 13734 25628 14310
rect 25662 13734 25674 14310
rect 25616 13722 25674 13734
rect 25744 14310 25802 14322
rect 25744 13734 25756 14310
rect 25790 13734 25802 14310
rect 25744 13722 25802 13734
rect 25856 14310 25914 14322
rect 25856 13734 25868 14310
rect 25902 13734 25914 14310
rect 25856 13722 25914 13734
rect 25984 14310 26042 14322
rect 25984 13734 25996 14310
rect 26030 13734 26042 14310
rect 25984 13722 26042 13734
rect 26096 14310 26154 14322
rect 26096 13734 26108 14310
rect 26142 13734 26154 14310
rect 26096 13722 26154 13734
rect 26224 14310 26282 14322
rect 26224 13734 26236 14310
rect 26270 13734 26282 14310
rect 26224 13722 26282 13734
rect 26336 14310 26394 14322
rect 26336 13734 26348 14310
rect 26382 13734 26394 14310
rect 26336 13722 26394 13734
rect 26464 14310 26522 14322
rect 26464 13734 26476 14310
rect 26510 13734 26522 14310
rect 26464 13722 26522 13734
rect 26576 14310 26634 14322
rect 26576 13734 26588 14310
rect 26622 13734 26634 14310
rect 26576 13722 26634 13734
rect 26704 14310 26762 14322
rect 26704 13734 26716 14310
rect 26750 13734 26762 14310
rect 26704 13722 26762 13734
rect 26816 14310 26874 14322
rect 26816 13734 26828 14310
rect 26862 13734 26874 14310
rect 26816 13722 26874 13734
rect 26944 14310 27002 14322
rect 26944 13734 26956 14310
rect 26990 13734 27002 14310
rect 26944 13722 27002 13734
rect 27056 14310 27114 14322
rect 27056 13734 27068 14310
rect 27102 13734 27114 14310
rect 27056 13722 27114 13734
rect 27184 14310 27242 14322
rect 27184 13734 27196 14310
rect 27230 13734 27242 14310
rect 27184 13722 27242 13734
rect 27296 14310 27354 14322
rect 27296 13734 27308 14310
rect 27342 13734 27354 14310
rect 27296 13722 27354 13734
rect 27424 14310 27482 14322
rect 27424 13734 27436 14310
rect 27470 13734 27482 14310
rect 27424 13722 27482 13734
rect 27536 14310 27594 14322
rect 27536 13734 27548 14310
rect 27582 13734 27594 14310
rect 27536 13722 27594 13734
rect 27664 14310 27722 14322
rect 27664 13734 27676 14310
rect 27710 13734 27722 14310
rect 27664 13722 27722 13734
rect 27776 14310 27834 14322
rect 27776 13734 27788 14310
rect 27822 13734 27834 14310
rect 27776 13722 27834 13734
rect 27904 14310 27962 14322
rect 27904 13734 27916 14310
rect 27950 13734 27962 14310
rect 27904 13722 27962 13734
rect 28016 14310 28074 14322
rect 28016 13734 28028 14310
rect 28062 13734 28074 14310
rect 28016 13722 28074 13734
rect 28144 14310 28202 14322
rect 28144 13734 28156 14310
rect 28190 13734 28202 14310
rect 28144 13722 28202 13734
rect 28256 14310 28314 14322
rect 28256 13734 28268 14310
rect 28302 13734 28314 14310
rect 28256 13722 28314 13734
rect 28384 14310 28442 14322
rect 28384 13734 28396 14310
rect 28430 13734 28442 14310
rect 28384 13722 28442 13734
rect 28496 14310 28554 14322
rect 28496 13734 28508 14310
rect 28542 13734 28554 14310
rect 28496 13722 28554 13734
rect 28624 14310 28682 14322
rect 28624 13734 28636 14310
rect 28670 13734 28682 14310
rect 28624 13722 28682 13734
rect 28736 14310 28794 14322
rect 28736 13734 28748 14310
rect 28782 13734 28794 14310
rect 28736 13722 28794 13734
rect 28864 14310 28922 14322
rect 28864 13734 28876 14310
rect 28910 13734 28922 14310
rect 28864 13722 28922 13734
rect 28976 14310 29034 14322
rect 28976 13734 28988 14310
rect 29022 13734 29034 14310
rect 28976 13722 29034 13734
rect 29104 14310 29162 14322
rect 29104 13734 29116 14310
rect 29150 13734 29162 14310
rect 29104 13722 29162 13734
rect 29216 14310 29274 14322
rect 29216 13734 29228 14310
rect 29262 13734 29274 14310
rect 29216 13722 29274 13734
rect 29344 14310 29402 14322
rect 29344 13734 29356 14310
rect 29390 13734 29402 14310
rect 29344 13722 29402 13734
rect 24176 2462 24234 2474
rect 24176 1886 24188 2462
rect 24222 1886 24234 2462
rect 24176 1874 24234 1886
rect 24304 2462 24362 2474
rect 24304 1886 24316 2462
rect 24350 1886 24362 2462
rect 24304 1874 24362 1886
rect 24416 2462 24474 2474
rect 24416 1886 24428 2462
rect 24462 1886 24474 2462
rect 24416 1874 24474 1886
rect 24544 2462 24602 2474
rect 24544 1886 24556 2462
rect 24590 1886 24602 2462
rect 24544 1874 24602 1886
rect 24656 2462 24714 2474
rect 24656 1886 24668 2462
rect 24702 1886 24714 2462
rect 24656 1874 24714 1886
rect 24784 2462 24842 2474
rect 24784 1886 24796 2462
rect 24830 1886 24842 2462
rect 24784 1874 24842 1886
rect 24896 2462 24954 2474
rect 24896 1886 24908 2462
rect 24942 1886 24954 2462
rect 24896 1874 24954 1886
rect 25024 2462 25082 2474
rect 25024 1886 25036 2462
rect 25070 1886 25082 2462
rect 25024 1874 25082 1886
rect 24176 1654 24234 1666
rect 24176 1078 24188 1654
rect 24222 1078 24234 1654
rect 24176 1066 24234 1078
rect 24304 1654 24362 1666
rect 24304 1078 24316 1654
rect 24350 1078 24362 1654
rect 24304 1066 24362 1078
rect 24416 1654 24474 1666
rect 24416 1078 24428 1654
rect 24462 1078 24474 1654
rect 24416 1066 24474 1078
rect 24544 1654 24602 1666
rect 24544 1078 24556 1654
rect 24590 1078 24602 1654
rect 24544 1066 24602 1078
rect 24656 1654 24714 1666
rect 24656 1078 24668 1654
rect 24702 1078 24714 1654
rect 24656 1066 24714 1078
rect 24784 1654 24842 1666
rect 24784 1078 24796 1654
rect 24830 1078 24842 1654
rect 24784 1066 24842 1078
rect 24896 1654 24954 1666
rect 24896 1078 24908 1654
rect 24942 1078 24954 1654
rect 24896 1066 24954 1078
rect 25024 1654 25082 1666
rect 25024 1078 25036 1654
rect 25070 1078 25082 1654
rect 25024 1066 25082 1078
<< pdiff >>
rect 10552 11100 10610 11112
rect 10552 10324 10564 11100
rect 10598 10324 10610 11100
rect 10552 10312 10610 10324
rect 11010 11100 11068 11112
rect 11010 10324 11022 11100
rect 11056 10324 11068 11100
rect 11010 10312 11068 10324
rect 11140 11100 11198 11112
rect 11140 10324 11152 11100
rect 11186 10324 11198 11100
rect 11140 10312 11198 10324
rect 11598 11100 11656 11112
rect 11598 10324 11610 11100
rect 11644 10324 11656 11100
rect 11598 10312 11656 10324
rect 11728 11100 11786 11112
rect 11728 10324 11740 11100
rect 11774 10324 11786 11100
rect 11728 10312 11786 10324
rect 12186 11100 12244 11112
rect 12186 10324 12198 11100
rect 12232 10324 12244 11100
rect 12186 10312 12244 10324
rect 12316 11100 12374 11112
rect 12316 10324 12328 11100
rect 12362 10324 12374 11100
rect 12316 10312 12374 10324
rect 12774 11100 12832 11112
rect 12774 10324 12786 11100
rect 12820 10324 12832 11100
rect 12774 10312 12832 10324
rect 12904 11100 12962 11112
rect 12904 10324 12916 11100
rect 12950 10324 12962 11100
rect 12904 10312 12962 10324
rect 13362 11100 13420 11112
rect 13362 10324 13374 11100
rect 13408 10324 13420 11100
rect 13362 10312 13420 10324
rect 13492 11100 13550 11112
rect 13492 10324 13504 11100
rect 13538 10324 13550 11100
rect 13492 10312 13550 10324
rect 13950 11100 14008 11112
rect 13950 10324 13962 11100
rect 13996 10324 14008 11100
rect 13950 10312 14008 10324
rect 14080 11100 14138 11112
rect 14080 10324 14092 11100
rect 14126 10324 14138 11100
rect 14080 10312 14138 10324
rect 14538 11100 14596 11112
rect 14538 10324 14550 11100
rect 14584 10324 14596 11100
rect 14538 10312 14596 10324
rect 14668 11100 14726 11112
rect 14668 10324 14680 11100
rect 14714 10324 14726 11100
rect 14668 10312 14726 10324
rect 15126 11100 15184 11112
rect 15126 10324 15138 11100
rect 15172 10324 15184 11100
rect 15126 10312 15184 10324
rect 15256 11100 15314 11112
rect 15256 10324 15268 11100
rect 15302 10324 15314 11100
rect 15256 10312 15314 10324
rect 15714 11100 15772 11112
rect 15714 10324 15726 11100
rect 15760 10324 15772 11100
rect 15714 10312 15772 10324
rect 15844 11100 15902 11112
rect 15844 10324 15856 11100
rect 15890 10324 15902 11100
rect 15844 10312 15902 10324
rect 16302 11100 16360 11112
rect 16302 10324 16314 11100
rect 16348 10324 16360 11100
rect 16302 10312 16360 10324
rect 16432 11100 16490 11112
rect 16432 10324 16444 11100
rect 16478 10324 16490 11100
rect 16432 10312 16490 10324
rect 16890 11100 16948 11112
rect 16890 10324 16902 11100
rect 16936 10324 16948 11100
rect 16890 10312 16948 10324
rect 17020 11100 17078 11112
rect 17020 10324 17032 11100
rect 17066 10324 17078 11100
rect 17020 10312 17078 10324
rect 17478 11100 17536 11112
rect 17478 10324 17490 11100
rect 17524 10324 17536 11100
rect 17478 10312 17536 10324
rect 17608 11100 17666 11112
rect 17608 10324 17620 11100
rect 17654 10324 17666 11100
rect 17608 10312 17666 10324
rect 18066 11100 18124 11112
rect 18066 10324 18078 11100
rect 18112 10324 18124 11100
rect 18066 10312 18124 10324
rect 18196 11100 18254 11112
rect 18196 10324 18208 11100
rect 18242 10324 18254 11100
rect 18196 10312 18254 10324
rect 18654 11100 18712 11112
rect 18654 10324 18666 11100
rect 18700 10324 18712 11100
rect 18654 10312 18712 10324
rect 18784 11100 18842 11112
rect 18784 10324 18796 11100
rect 18830 10324 18842 11100
rect 18784 10312 18842 10324
rect 19242 11100 19300 11112
rect 19242 10324 19254 11100
rect 19288 10324 19300 11100
rect 19242 10312 19300 10324
rect 19372 11100 19430 11112
rect 19372 10324 19384 11100
rect 19418 10324 19430 11100
rect 19372 10312 19430 10324
rect 19830 11100 19888 11112
rect 19830 10324 19842 11100
rect 19876 10324 19888 11100
rect 19830 10312 19888 10324
rect 19960 11100 20018 11112
rect 19960 10324 19972 11100
rect 20006 10324 20018 11100
rect 19960 10312 20018 10324
rect 20418 11100 20476 11112
rect 20418 10324 20430 11100
rect 20464 10324 20476 11100
rect 20418 10312 20476 10324
rect 20548 11100 20606 11112
rect 20548 10324 20560 11100
rect 20594 10324 20606 11100
rect 20548 10312 20606 10324
rect 21006 11100 21064 11112
rect 21006 10324 21018 11100
rect 21052 10324 21064 11100
rect 21006 10312 21064 10324
rect 21136 11100 21194 11112
rect 21136 10324 21148 11100
rect 21182 10324 21194 11100
rect 21136 10312 21194 10324
rect 21594 11100 21652 11112
rect 21594 10324 21606 11100
rect 21640 10324 21652 11100
rect 21594 10312 21652 10324
rect 21724 11100 21782 11112
rect 21724 10324 21736 11100
rect 21770 10324 21782 11100
rect 21724 10312 21782 10324
rect 22182 11100 22240 11112
rect 22182 10324 22194 11100
rect 22228 10324 22240 11100
rect 22182 10312 22240 10324
rect 22312 11100 22370 11112
rect 22312 10324 22324 11100
rect 22358 10324 22370 11100
rect 22312 10312 22370 10324
rect 22770 11100 22828 11112
rect 22770 10324 22782 11100
rect 22816 10324 22828 11100
rect 22770 10312 22828 10324
rect 22900 11100 22958 11112
rect 22900 10324 22912 11100
rect 22946 10324 22958 11100
rect 22900 10312 22958 10324
rect 23358 11100 23416 11112
rect 23358 10324 23370 11100
rect 23404 10324 23416 11100
rect 23358 10312 23416 10324
rect 23488 11100 23546 11112
rect 23488 10324 23500 11100
rect 23534 10324 23546 11100
rect 23488 10312 23546 10324
rect 23946 11100 24004 11112
rect 23946 10324 23958 11100
rect 23992 10324 24004 11100
rect 23946 10312 24004 10324
rect 24076 11100 24134 11112
rect 24076 10324 24088 11100
rect 24122 10324 24134 11100
rect 24076 10312 24134 10324
rect 24534 11100 24592 11112
rect 24534 10324 24546 11100
rect 24580 10324 24592 11100
rect 24534 10312 24592 10324
rect 24664 11100 24722 11112
rect 24664 10324 24676 11100
rect 24710 10324 24722 11100
rect 24664 10312 24722 10324
rect 25122 11100 25180 11112
rect 25122 10324 25134 11100
rect 25168 10324 25180 11100
rect 25122 10312 25180 10324
rect 25252 11100 25310 11112
rect 25252 10324 25264 11100
rect 25298 10324 25310 11100
rect 25252 10312 25310 10324
rect 25710 11100 25768 11112
rect 25710 10324 25722 11100
rect 25756 10324 25768 11100
rect 25710 10312 25768 10324
rect 25840 11100 25898 11112
rect 25840 10324 25852 11100
rect 25886 10324 25898 11100
rect 25840 10312 25898 10324
rect 26298 11100 26356 11112
rect 26298 10324 26310 11100
rect 26344 10324 26356 11100
rect 26298 10312 26356 10324
rect 26428 11100 26486 11112
rect 26428 10324 26440 11100
rect 26474 10324 26486 11100
rect 26428 10312 26486 10324
rect 26886 11100 26944 11112
rect 26886 10324 26898 11100
rect 26932 10324 26944 11100
rect 26886 10312 26944 10324
rect 27016 11100 27074 11112
rect 27016 10324 27028 11100
rect 27062 10324 27074 11100
rect 27016 10312 27074 10324
rect 27474 11100 27532 11112
rect 27474 10324 27486 11100
rect 27520 10324 27532 11100
rect 27474 10312 27532 10324
rect 27604 11100 27662 11112
rect 27604 10324 27616 11100
rect 27650 10324 27662 11100
rect 27604 10312 27662 10324
rect 28062 11100 28120 11112
rect 28062 10324 28074 11100
rect 28108 10324 28120 11100
rect 28062 10312 28120 10324
rect 28192 11100 28250 11112
rect 28192 10324 28204 11100
rect 28238 10324 28250 11100
rect 28192 10312 28250 10324
rect 28650 11100 28708 11112
rect 28650 10324 28662 11100
rect 28696 10324 28708 11100
rect 28650 10312 28708 10324
rect 28780 11100 28838 11112
rect 28780 10324 28792 11100
rect 28826 10324 28838 11100
rect 28780 10312 28838 10324
rect 29238 11100 29296 11112
rect 29238 10324 29250 11100
rect 29284 10324 29296 11100
rect 29238 10312 29296 10324
rect 29368 11100 29426 11112
rect 29368 10324 29380 11100
rect 29414 10324 29426 11100
rect 29368 10312 29426 10324
rect 29826 11100 29884 11112
rect 29826 10324 29838 11100
rect 29872 10324 29884 11100
rect 29826 10312 29884 10324
rect 29956 11100 30014 11112
rect 29956 10324 29968 11100
rect 30002 10324 30014 11100
rect 29956 10312 30014 10324
rect 30414 11100 30472 11112
rect 30414 10324 30426 11100
rect 30460 10324 30472 11100
rect 30414 10312 30472 10324
rect 30544 11100 30602 11112
rect 30544 10324 30556 11100
rect 30590 10324 30602 11100
rect 30544 10312 30602 10324
rect 31002 11100 31060 11112
rect 31002 10324 31014 11100
rect 31048 10324 31060 11100
rect 31002 10312 31060 10324
rect 31132 11100 31190 11112
rect 31132 10324 31144 11100
rect 31178 10324 31190 11100
rect 31132 10312 31190 10324
rect 31590 11100 31648 11112
rect 31590 10324 31602 11100
rect 31636 10324 31648 11100
rect 31590 10312 31648 10324
rect 31720 11100 31778 11112
rect 31720 10324 31732 11100
rect 31766 10324 31778 11100
rect 31720 10312 31778 10324
rect 32178 11100 32236 11112
rect 32178 10324 32190 11100
rect 32224 10324 32236 11100
rect 32178 10312 32236 10324
rect 32308 11100 32366 11112
rect 32308 10324 32320 11100
rect 32354 10324 32366 11100
rect 32308 10312 32366 10324
rect 32766 11100 32824 11112
rect 32766 10324 32778 11100
rect 32812 10324 32824 11100
rect 32766 10312 32824 10324
rect 32896 11100 32954 11112
rect 32896 10324 32908 11100
rect 32942 10324 32954 11100
rect 32896 10312 32954 10324
rect 33354 11100 33412 11112
rect 33354 10324 33366 11100
rect 33400 10324 33412 11100
rect 33354 10312 33412 10324
rect 33484 11100 33542 11112
rect 33484 10324 33496 11100
rect 33530 10324 33542 11100
rect 33484 10312 33542 10324
rect 33942 11100 34000 11112
rect 33942 10324 33954 11100
rect 33988 10324 34000 11100
rect 33942 10312 34000 10324
rect 34072 11100 34130 11112
rect 34072 10324 34084 11100
rect 34118 10324 34130 11100
rect 34072 10312 34130 10324
rect 34530 11100 34588 11112
rect 34530 10324 34542 11100
rect 34576 10324 34588 11100
rect 34530 10312 34588 10324
rect 34660 11100 34718 11112
rect 34660 10324 34672 11100
rect 34706 10324 34718 11100
rect 34660 10312 34718 10324
rect 35118 11100 35176 11112
rect 35118 10324 35130 11100
rect 35164 10324 35176 11100
rect 35118 10312 35176 10324
rect 35248 11100 35306 11112
rect 35248 10324 35260 11100
rect 35294 10324 35306 11100
rect 35248 10312 35306 10324
rect 35706 11100 35764 11112
rect 35706 10324 35718 11100
rect 35752 10324 35764 11100
rect 35706 10312 35764 10324
rect 35836 11100 35894 11112
rect 35836 10324 35848 11100
rect 35882 10324 35894 11100
rect 35836 10312 35894 10324
rect 36294 11100 36352 11112
rect 36294 10324 36306 11100
rect 36340 10324 36352 11100
rect 36294 10312 36352 10324
rect 36424 11100 36482 11112
rect 36424 10324 36436 11100
rect 36470 10324 36482 11100
rect 36424 10312 36482 10324
rect 36882 11100 36940 11112
rect 36882 10324 36894 11100
rect 36928 10324 36940 11100
rect 36882 10312 36940 10324
rect 37012 11100 37070 11112
rect 37012 10324 37024 11100
rect 37058 10324 37070 11100
rect 37012 10312 37070 10324
rect 37470 11100 37528 11112
rect 37470 10324 37482 11100
rect 37516 10324 37528 11100
rect 37470 10312 37528 10324
rect 37600 11100 37658 11112
rect 37600 10324 37612 11100
rect 37646 10324 37658 11100
rect 37600 10312 37658 10324
rect 38058 11100 38116 11112
rect 38058 10324 38070 11100
rect 38104 10324 38116 11100
rect 38058 10312 38116 10324
rect 38188 11100 38246 11112
rect 38188 10324 38200 11100
rect 38234 10324 38246 11100
rect 38188 10312 38246 10324
rect 38646 11100 38704 11112
rect 38646 10324 38658 11100
rect 38692 10324 38704 11100
rect 38646 10312 38704 10324
rect 10552 10100 10610 10112
rect 10552 9324 10564 10100
rect 10598 9324 10610 10100
rect 10552 9312 10610 9324
rect 11010 10100 11068 10112
rect 11010 9324 11022 10100
rect 11056 9324 11068 10100
rect 11010 9312 11068 9324
rect 11140 10100 11198 10112
rect 11140 9324 11152 10100
rect 11186 9324 11198 10100
rect 11140 9312 11198 9324
rect 11598 10100 11656 10112
rect 11598 9324 11610 10100
rect 11644 9324 11656 10100
rect 11598 9312 11656 9324
rect 11728 10100 11786 10112
rect 11728 9324 11740 10100
rect 11774 9324 11786 10100
rect 11728 9312 11786 9324
rect 12186 10100 12244 10112
rect 12186 9324 12198 10100
rect 12232 9324 12244 10100
rect 12186 9312 12244 9324
rect 12316 10100 12374 10112
rect 12316 9324 12328 10100
rect 12362 9324 12374 10100
rect 12316 9312 12374 9324
rect 12774 10100 12832 10112
rect 12774 9324 12786 10100
rect 12820 9324 12832 10100
rect 12774 9312 12832 9324
rect 12904 10100 12962 10112
rect 12904 9324 12916 10100
rect 12950 9324 12962 10100
rect 12904 9312 12962 9324
rect 13362 10100 13420 10112
rect 13362 9324 13374 10100
rect 13408 9324 13420 10100
rect 13362 9312 13420 9324
rect 13492 10100 13550 10112
rect 13492 9324 13504 10100
rect 13538 9324 13550 10100
rect 13492 9312 13550 9324
rect 13950 10100 14008 10112
rect 13950 9324 13962 10100
rect 13996 9324 14008 10100
rect 13950 9312 14008 9324
rect 14080 10100 14138 10112
rect 14080 9324 14092 10100
rect 14126 9324 14138 10100
rect 14080 9312 14138 9324
rect 14538 10100 14596 10112
rect 14538 9324 14550 10100
rect 14584 9324 14596 10100
rect 14538 9312 14596 9324
rect 14668 10100 14726 10112
rect 14668 9324 14680 10100
rect 14714 9324 14726 10100
rect 14668 9312 14726 9324
rect 15126 10100 15184 10112
rect 15126 9324 15138 10100
rect 15172 9324 15184 10100
rect 15126 9312 15184 9324
rect 15256 10100 15314 10112
rect 15256 9324 15268 10100
rect 15302 9324 15314 10100
rect 15256 9312 15314 9324
rect 15714 10100 15772 10112
rect 15714 9324 15726 10100
rect 15760 9324 15772 10100
rect 15714 9312 15772 9324
rect 15844 10100 15902 10112
rect 15844 9324 15856 10100
rect 15890 9324 15902 10100
rect 15844 9312 15902 9324
rect 16302 10100 16360 10112
rect 16302 9324 16314 10100
rect 16348 9324 16360 10100
rect 16302 9312 16360 9324
rect 16432 10100 16490 10112
rect 16432 9324 16444 10100
rect 16478 9324 16490 10100
rect 16432 9312 16490 9324
rect 16890 10100 16948 10112
rect 16890 9324 16902 10100
rect 16936 9324 16948 10100
rect 16890 9312 16948 9324
rect 17020 10100 17078 10112
rect 17020 9324 17032 10100
rect 17066 9324 17078 10100
rect 17020 9312 17078 9324
rect 17478 10100 17536 10112
rect 17478 9324 17490 10100
rect 17524 9324 17536 10100
rect 17478 9312 17536 9324
rect 17608 10100 17666 10112
rect 17608 9324 17620 10100
rect 17654 9324 17666 10100
rect 17608 9312 17666 9324
rect 18066 10100 18124 10112
rect 18066 9324 18078 10100
rect 18112 9324 18124 10100
rect 18066 9312 18124 9324
rect 18196 10100 18254 10112
rect 18196 9324 18208 10100
rect 18242 9324 18254 10100
rect 18196 9312 18254 9324
rect 18654 10100 18712 10112
rect 18654 9324 18666 10100
rect 18700 9324 18712 10100
rect 18654 9312 18712 9324
rect 18784 10100 18842 10112
rect 18784 9324 18796 10100
rect 18830 9324 18842 10100
rect 18784 9312 18842 9324
rect 19242 10100 19300 10112
rect 19242 9324 19254 10100
rect 19288 9324 19300 10100
rect 19242 9312 19300 9324
rect 19372 10100 19430 10112
rect 19372 9324 19384 10100
rect 19418 9324 19430 10100
rect 19372 9312 19430 9324
rect 19830 10100 19888 10112
rect 19830 9324 19842 10100
rect 19876 9324 19888 10100
rect 19830 9312 19888 9324
rect 19960 10100 20018 10112
rect 19960 9324 19972 10100
rect 20006 9324 20018 10100
rect 19960 9312 20018 9324
rect 20418 10100 20476 10112
rect 20418 9324 20430 10100
rect 20464 9324 20476 10100
rect 20418 9312 20476 9324
rect 20548 10100 20606 10112
rect 20548 9324 20560 10100
rect 20594 9324 20606 10100
rect 20548 9312 20606 9324
rect 21006 10100 21064 10112
rect 21006 9324 21018 10100
rect 21052 9324 21064 10100
rect 21006 9312 21064 9324
rect 21136 10100 21194 10112
rect 21136 9324 21148 10100
rect 21182 9324 21194 10100
rect 21136 9312 21194 9324
rect 21594 10100 21652 10112
rect 21594 9324 21606 10100
rect 21640 9324 21652 10100
rect 21594 9312 21652 9324
rect 21724 10100 21782 10112
rect 21724 9324 21736 10100
rect 21770 9324 21782 10100
rect 21724 9312 21782 9324
rect 22182 10100 22240 10112
rect 22182 9324 22194 10100
rect 22228 9324 22240 10100
rect 22182 9312 22240 9324
rect 22312 10100 22370 10112
rect 22312 9324 22324 10100
rect 22358 9324 22370 10100
rect 22312 9312 22370 9324
rect 22770 10100 22828 10112
rect 22770 9324 22782 10100
rect 22816 9324 22828 10100
rect 22770 9312 22828 9324
rect 22900 10100 22958 10112
rect 22900 9324 22912 10100
rect 22946 9324 22958 10100
rect 22900 9312 22958 9324
rect 23358 10100 23416 10112
rect 23358 9324 23370 10100
rect 23404 9324 23416 10100
rect 23358 9312 23416 9324
rect 23488 10100 23546 10112
rect 23488 9324 23500 10100
rect 23534 9324 23546 10100
rect 23488 9312 23546 9324
rect 23946 10100 24004 10112
rect 23946 9324 23958 10100
rect 23992 9324 24004 10100
rect 23946 9312 24004 9324
rect 24076 10100 24134 10112
rect 24076 9324 24088 10100
rect 24122 9324 24134 10100
rect 24076 9312 24134 9324
rect 24534 10100 24592 10112
rect 24534 9324 24546 10100
rect 24580 9324 24592 10100
rect 24534 9312 24592 9324
rect 24664 10100 24722 10112
rect 24664 9324 24676 10100
rect 24710 9324 24722 10100
rect 24664 9312 24722 9324
rect 25122 10100 25180 10112
rect 25122 9324 25134 10100
rect 25168 9324 25180 10100
rect 25122 9312 25180 9324
rect 25252 10100 25310 10112
rect 25252 9324 25264 10100
rect 25298 9324 25310 10100
rect 25252 9312 25310 9324
rect 25710 10100 25768 10112
rect 25710 9324 25722 10100
rect 25756 9324 25768 10100
rect 25710 9312 25768 9324
rect 25840 10100 25898 10112
rect 25840 9324 25852 10100
rect 25886 9324 25898 10100
rect 25840 9312 25898 9324
rect 26298 10100 26356 10112
rect 26298 9324 26310 10100
rect 26344 9324 26356 10100
rect 26298 9312 26356 9324
rect 26428 10100 26486 10112
rect 26428 9324 26440 10100
rect 26474 9324 26486 10100
rect 26428 9312 26486 9324
rect 26886 10100 26944 10112
rect 26886 9324 26898 10100
rect 26932 9324 26944 10100
rect 26886 9312 26944 9324
rect 27016 10100 27074 10112
rect 27016 9324 27028 10100
rect 27062 9324 27074 10100
rect 27016 9312 27074 9324
rect 27474 10100 27532 10112
rect 27474 9324 27486 10100
rect 27520 9324 27532 10100
rect 27474 9312 27532 9324
rect 27604 10100 27662 10112
rect 27604 9324 27616 10100
rect 27650 9324 27662 10100
rect 27604 9312 27662 9324
rect 28062 10100 28120 10112
rect 28062 9324 28074 10100
rect 28108 9324 28120 10100
rect 28062 9312 28120 9324
rect 28192 10100 28250 10112
rect 28192 9324 28204 10100
rect 28238 9324 28250 10100
rect 28192 9312 28250 9324
rect 28650 10100 28708 10112
rect 28650 9324 28662 10100
rect 28696 9324 28708 10100
rect 28650 9312 28708 9324
rect 28780 10100 28838 10112
rect 28780 9324 28792 10100
rect 28826 9324 28838 10100
rect 28780 9312 28838 9324
rect 29238 10100 29296 10112
rect 29238 9324 29250 10100
rect 29284 9324 29296 10100
rect 29238 9312 29296 9324
rect 29368 10100 29426 10112
rect 29368 9324 29380 10100
rect 29414 9324 29426 10100
rect 29368 9312 29426 9324
rect 29826 10100 29884 10112
rect 29826 9324 29838 10100
rect 29872 9324 29884 10100
rect 29826 9312 29884 9324
rect 29956 10100 30014 10112
rect 29956 9324 29968 10100
rect 30002 9324 30014 10100
rect 29956 9312 30014 9324
rect 30414 10100 30472 10112
rect 30414 9324 30426 10100
rect 30460 9324 30472 10100
rect 30414 9312 30472 9324
rect 30544 10100 30602 10112
rect 30544 9324 30556 10100
rect 30590 9324 30602 10100
rect 30544 9312 30602 9324
rect 31002 10100 31060 10112
rect 31002 9324 31014 10100
rect 31048 9324 31060 10100
rect 31002 9312 31060 9324
rect 31132 10100 31190 10112
rect 31132 9324 31144 10100
rect 31178 9324 31190 10100
rect 31132 9312 31190 9324
rect 31590 10100 31648 10112
rect 31590 9324 31602 10100
rect 31636 9324 31648 10100
rect 31590 9312 31648 9324
rect 31720 10100 31778 10112
rect 31720 9324 31732 10100
rect 31766 9324 31778 10100
rect 31720 9312 31778 9324
rect 32178 10100 32236 10112
rect 32178 9324 32190 10100
rect 32224 9324 32236 10100
rect 32178 9312 32236 9324
rect 32308 10100 32366 10112
rect 32308 9324 32320 10100
rect 32354 9324 32366 10100
rect 32308 9312 32366 9324
rect 32766 10100 32824 10112
rect 32766 9324 32778 10100
rect 32812 9324 32824 10100
rect 32766 9312 32824 9324
rect 32896 10100 32954 10112
rect 32896 9324 32908 10100
rect 32942 9324 32954 10100
rect 32896 9312 32954 9324
rect 33354 10100 33412 10112
rect 33354 9324 33366 10100
rect 33400 9324 33412 10100
rect 33354 9312 33412 9324
rect 33484 10100 33542 10112
rect 33484 9324 33496 10100
rect 33530 9324 33542 10100
rect 33484 9312 33542 9324
rect 33942 10100 34000 10112
rect 33942 9324 33954 10100
rect 33988 9324 34000 10100
rect 33942 9312 34000 9324
rect 34072 10100 34130 10112
rect 34072 9324 34084 10100
rect 34118 9324 34130 10100
rect 34072 9312 34130 9324
rect 34530 10100 34588 10112
rect 34530 9324 34542 10100
rect 34576 9324 34588 10100
rect 34530 9312 34588 9324
rect 34660 10100 34718 10112
rect 34660 9324 34672 10100
rect 34706 9324 34718 10100
rect 34660 9312 34718 9324
rect 35118 10100 35176 10112
rect 35118 9324 35130 10100
rect 35164 9324 35176 10100
rect 35118 9312 35176 9324
rect 35248 10100 35306 10112
rect 35248 9324 35260 10100
rect 35294 9324 35306 10100
rect 35248 9312 35306 9324
rect 35706 10100 35764 10112
rect 35706 9324 35718 10100
rect 35752 9324 35764 10100
rect 35706 9312 35764 9324
rect 35836 10100 35894 10112
rect 35836 9324 35848 10100
rect 35882 9324 35894 10100
rect 35836 9312 35894 9324
rect 36294 10100 36352 10112
rect 36294 9324 36306 10100
rect 36340 9324 36352 10100
rect 36294 9312 36352 9324
rect 36424 10100 36482 10112
rect 36424 9324 36436 10100
rect 36470 9324 36482 10100
rect 36424 9312 36482 9324
rect 36882 10100 36940 10112
rect 36882 9324 36894 10100
rect 36928 9324 36940 10100
rect 36882 9312 36940 9324
rect 37012 10100 37070 10112
rect 37012 9324 37024 10100
rect 37058 9324 37070 10100
rect 37012 9312 37070 9324
rect 37470 10100 37528 10112
rect 37470 9324 37482 10100
rect 37516 9324 37528 10100
rect 37470 9312 37528 9324
rect 37600 10100 37658 10112
rect 37600 9324 37612 10100
rect 37646 9324 37658 10100
rect 37600 9312 37658 9324
rect 38058 10100 38116 10112
rect 38058 9324 38070 10100
rect 38104 9324 38116 10100
rect 38058 9312 38116 9324
rect 38188 10100 38246 10112
rect 38188 9324 38200 10100
rect 38234 9324 38246 10100
rect 38188 9312 38246 9324
rect 38646 10100 38704 10112
rect 38646 9324 38658 10100
rect 38692 9324 38704 10100
rect 38646 9312 38704 9324
rect 10552 9100 10610 9112
rect 10552 8324 10564 9100
rect 10598 8324 10610 9100
rect 10552 8312 10610 8324
rect 11010 9100 11068 9112
rect 11010 8324 11022 9100
rect 11056 8324 11068 9100
rect 11010 8312 11068 8324
rect 11140 9100 11198 9112
rect 11140 8324 11152 9100
rect 11186 8324 11198 9100
rect 11140 8312 11198 8324
rect 11598 9100 11656 9112
rect 11598 8324 11610 9100
rect 11644 8324 11656 9100
rect 11598 8312 11656 8324
rect 11728 9100 11786 9112
rect 11728 8324 11740 9100
rect 11774 8324 11786 9100
rect 11728 8312 11786 8324
rect 12186 9100 12244 9112
rect 12186 8324 12198 9100
rect 12232 8324 12244 9100
rect 12186 8312 12244 8324
rect 12316 9100 12374 9112
rect 12316 8324 12328 9100
rect 12362 8324 12374 9100
rect 12316 8312 12374 8324
rect 12774 9100 12832 9112
rect 12774 8324 12786 9100
rect 12820 8324 12832 9100
rect 12774 8312 12832 8324
rect 12904 9100 12962 9112
rect 12904 8324 12916 9100
rect 12950 8324 12962 9100
rect 12904 8312 12962 8324
rect 13362 9100 13420 9112
rect 13362 8324 13374 9100
rect 13408 8324 13420 9100
rect 13362 8312 13420 8324
rect 13492 9100 13550 9112
rect 13492 8324 13504 9100
rect 13538 8324 13550 9100
rect 13492 8312 13550 8324
rect 13950 9100 14008 9112
rect 13950 8324 13962 9100
rect 13996 8324 14008 9100
rect 13950 8312 14008 8324
rect 14080 9100 14138 9112
rect 14080 8324 14092 9100
rect 14126 8324 14138 9100
rect 14080 8312 14138 8324
rect 14538 9100 14596 9112
rect 14538 8324 14550 9100
rect 14584 8324 14596 9100
rect 14538 8312 14596 8324
rect 14668 9100 14726 9112
rect 14668 8324 14680 9100
rect 14714 8324 14726 9100
rect 14668 8312 14726 8324
rect 15126 9100 15184 9112
rect 15126 8324 15138 9100
rect 15172 8324 15184 9100
rect 15126 8312 15184 8324
rect 15256 9100 15314 9112
rect 15256 8324 15268 9100
rect 15302 8324 15314 9100
rect 15256 8312 15314 8324
rect 15714 9100 15772 9112
rect 15714 8324 15726 9100
rect 15760 8324 15772 9100
rect 15714 8312 15772 8324
rect 15844 9100 15902 9112
rect 15844 8324 15856 9100
rect 15890 8324 15902 9100
rect 15844 8312 15902 8324
rect 16302 9100 16360 9112
rect 16302 8324 16314 9100
rect 16348 8324 16360 9100
rect 16302 8312 16360 8324
rect 16432 9100 16490 9112
rect 16432 8324 16444 9100
rect 16478 8324 16490 9100
rect 16432 8312 16490 8324
rect 16890 9100 16948 9112
rect 16890 8324 16902 9100
rect 16936 8324 16948 9100
rect 16890 8312 16948 8324
rect 17020 9100 17078 9112
rect 17020 8324 17032 9100
rect 17066 8324 17078 9100
rect 17020 8312 17078 8324
rect 17478 9100 17536 9112
rect 17478 8324 17490 9100
rect 17524 8324 17536 9100
rect 17478 8312 17536 8324
rect 17608 9100 17666 9112
rect 17608 8324 17620 9100
rect 17654 8324 17666 9100
rect 17608 8312 17666 8324
rect 18066 9100 18124 9112
rect 18066 8324 18078 9100
rect 18112 8324 18124 9100
rect 18066 8312 18124 8324
rect 18196 9100 18254 9112
rect 18196 8324 18208 9100
rect 18242 8324 18254 9100
rect 18196 8312 18254 8324
rect 18654 9100 18712 9112
rect 18654 8324 18666 9100
rect 18700 8324 18712 9100
rect 18654 8312 18712 8324
rect 18784 9100 18842 9112
rect 18784 8324 18796 9100
rect 18830 8324 18842 9100
rect 18784 8312 18842 8324
rect 19242 9100 19300 9112
rect 19242 8324 19254 9100
rect 19288 8324 19300 9100
rect 19242 8312 19300 8324
rect 19372 9100 19430 9112
rect 19372 8324 19384 9100
rect 19418 8324 19430 9100
rect 19372 8312 19430 8324
rect 19830 9100 19888 9112
rect 19830 8324 19842 9100
rect 19876 8324 19888 9100
rect 19830 8312 19888 8324
rect 19960 9100 20018 9112
rect 19960 8324 19972 9100
rect 20006 8324 20018 9100
rect 19960 8312 20018 8324
rect 20418 9100 20476 9112
rect 20418 8324 20430 9100
rect 20464 8324 20476 9100
rect 20418 8312 20476 8324
rect 20548 9100 20606 9112
rect 20548 8324 20560 9100
rect 20594 8324 20606 9100
rect 20548 8312 20606 8324
rect 21006 9100 21064 9112
rect 21006 8324 21018 9100
rect 21052 8324 21064 9100
rect 21006 8312 21064 8324
rect 21136 9100 21194 9112
rect 21136 8324 21148 9100
rect 21182 8324 21194 9100
rect 21136 8312 21194 8324
rect 21594 9100 21652 9112
rect 21594 8324 21606 9100
rect 21640 8324 21652 9100
rect 21594 8312 21652 8324
rect 21724 9100 21782 9112
rect 21724 8324 21736 9100
rect 21770 8324 21782 9100
rect 21724 8312 21782 8324
rect 22182 9100 22240 9112
rect 22182 8324 22194 9100
rect 22228 8324 22240 9100
rect 22182 8312 22240 8324
rect 22312 9100 22370 9112
rect 22312 8324 22324 9100
rect 22358 8324 22370 9100
rect 22312 8312 22370 8324
rect 22770 9100 22828 9112
rect 22770 8324 22782 9100
rect 22816 8324 22828 9100
rect 22770 8312 22828 8324
rect 22900 9100 22958 9112
rect 22900 8324 22912 9100
rect 22946 8324 22958 9100
rect 22900 8312 22958 8324
rect 23358 9100 23416 9112
rect 23358 8324 23370 9100
rect 23404 8324 23416 9100
rect 23358 8312 23416 8324
rect 23488 9100 23546 9112
rect 23488 8324 23500 9100
rect 23534 8324 23546 9100
rect 23488 8312 23546 8324
rect 23946 9100 24004 9112
rect 23946 8324 23958 9100
rect 23992 8324 24004 9100
rect 23946 8312 24004 8324
rect 24076 9100 24134 9112
rect 24076 8324 24088 9100
rect 24122 8324 24134 9100
rect 24076 8312 24134 8324
rect 24534 9100 24592 9112
rect 24534 8324 24546 9100
rect 24580 8324 24592 9100
rect 24534 8312 24592 8324
rect 24664 9100 24722 9112
rect 24664 8324 24676 9100
rect 24710 8324 24722 9100
rect 24664 8312 24722 8324
rect 25122 9100 25180 9112
rect 25122 8324 25134 9100
rect 25168 8324 25180 9100
rect 25122 8312 25180 8324
rect 25252 9100 25310 9112
rect 25252 8324 25264 9100
rect 25298 8324 25310 9100
rect 25252 8312 25310 8324
rect 25710 9100 25768 9112
rect 25710 8324 25722 9100
rect 25756 8324 25768 9100
rect 25710 8312 25768 8324
rect 25840 9100 25898 9112
rect 25840 8324 25852 9100
rect 25886 8324 25898 9100
rect 25840 8312 25898 8324
rect 26298 9100 26356 9112
rect 26298 8324 26310 9100
rect 26344 8324 26356 9100
rect 26298 8312 26356 8324
rect 26428 9100 26486 9112
rect 26428 8324 26440 9100
rect 26474 8324 26486 9100
rect 26428 8312 26486 8324
rect 26886 9100 26944 9112
rect 26886 8324 26898 9100
rect 26932 8324 26944 9100
rect 26886 8312 26944 8324
rect 27016 9100 27074 9112
rect 27016 8324 27028 9100
rect 27062 8324 27074 9100
rect 27016 8312 27074 8324
rect 27474 9100 27532 9112
rect 27474 8324 27486 9100
rect 27520 8324 27532 9100
rect 27474 8312 27532 8324
rect 27604 9100 27662 9112
rect 27604 8324 27616 9100
rect 27650 8324 27662 9100
rect 27604 8312 27662 8324
rect 28062 9100 28120 9112
rect 28062 8324 28074 9100
rect 28108 8324 28120 9100
rect 28062 8312 28120 8324
rect 28192 9100 28250 9112
rect 28192 8324 28204 9100
rect 28238 8324 28250 9100
rect 28192 8312 28250 8324
rect 28650 9100 28708 9112
rect 28650 8324 28662 9100
rect 28696 8324 28708 9100
rect 28650 8312 28708 8324
rect 28780 9100 28838 9112
rect 28780 8324 28792 9100
rect 28826 8324 28838 9100
rect 28780 8312 28838 8324
rect 29238 9100 29296 9112
rect 29238 8324 29250 9100
rect 29284 8324 29296 9100
rect 29238 8312 29296 8324
rect 29368 9100 29426 9112
rect 29368 8324 29380 9100
rect 29414 8324 29426 9100
rect 29368 8312 29426 8324
rect 29826 9100 29884 9112
rect 29826 8324 29838 9100
rect 29872 8324 29884 9100
rect 29826 8312 29884 8324
rect 29956 9100 30014 9112
rect 29956 8324 29968 9100
rect 30002 8324 30014 9100
rect 29956 8312 30014 8324
rect 30414 9100 30472 9112
rect 30414 8324 30426 9100
rect 30460 8324 30472 9100
rect 30414 8312 30472 8324
rect 30544 9100 30602 9112
rect 30544 8324 30556 9100
rect 30590 8324 30602 9100
rect 30544 8312 30602 8324
rect 31002 9100 31060 9112
rect 31002 8324 31014 9100
rect 31048 8324 31060 9100
rect 31002 8312 31060 8324
rect 31132 9100 31190 9112
rect 31132 8324 31144 9100
rect 31178 8324 31190 9100
rect 31132 8312 31190 8324
rect 31590 9100 31648 9112
rect 31590 8324 31602 9100
rect 31636 8324 31648 9100
rect 31590 8312 31648 8324
rect 31720 9100 31778 9112
rect 31720 8324 31732 9100
rect 31766 8324 31778 9100
rect 31720 8312 31778 8324
rect 32178 9100 32236 9112
rect 32178 8324 32190 9100
rect 32224 8324 32236 9100
rect 32178 8312 32236 8324
rect 32308 9100 32366 9112
rect 32308 8324 32320 9100
rect 32354 8324 32366 9100
rect 32308 8312 32366 8324
rect 32766 9100 32824 9112
rect 32766 8324 32778 9100
rect 32812 8324 32824 9100
rect 32766 8312 32824 8324
rect 32896 9100 32954 9112
rect 32896 8324 32908 9100
rect 32942 8324 32954 9100
rect 32896 8312 32954 8324
rect 33354 9100 33412 9112
rect 33354 8324 33366 9100
rect 33400 8324 33412 9100
rect 33354 8312 33412 8324
rect 33484 9100 33542 9112
rect 33484 8324 33496 9100
rect 33530 8324 33542 9100
rect 33484 8312 33542 8324
rect 33942 9100 34000 9112
rect 33942 8324 33954 9100
rect 33988 8324 34000 9100
rect 33942 8312 34000 8324
rect 34072 9100 34130 9112
rect 34072 8324 34084 9100
rect 34118 8324 34130 9100
rect 34072 8312 34130 8324
rect 34530 9100 34588 9112
rect 34530 8324 34542 9100
rect 34576 8324 34588 9100
rect 34530 8312 34588 8324
rect 34660 9100 34718 9112
rect 34660 8324 34672 9100
rect 34706 8324 34718 9100
rect 34660 8312 34718 8324
rect 35118 9100 35176 9112
rect 35118 8324 35130 9100
rect 35164 8324 35176 9100
rect 35118 8312 35176 8324
rect 35248 9100 35306 9112
rect 35248 8324 35260 9100
rect 35294 8324 35306 9100
rect 35248 8312 35306 8324
rect 35706 9100 35764 9112
rect 35706 8324 35718 9100
rect 35752 8324 35764 9100
rect 35706 8312 35764 8324
rect 35836 9100 35894 9112
rect 35836 8324 35848 9100
rect 35882 8324 35894 9100
rect 35836 8312 35894 8324
rect 36294 9100 36352 9112
rect 36294 8324 36306 9100
rect 36340 8324 36352 9100
rect 36294 8312 36352 8324
rect 36424 9100 36482 9112
rect 36424 8324 36436 9100
rect 36470 8324 36482 9100
rect 36424 8312 36482 8324
rect 36882 9100 36940 9112
rect 36882 8324 36894 9100
rect 36928 8324 36940 9100
rect 36882 8312 36940 8324
rect 37012 9100 37070 9112
rect 37012 8324 37024 9100
rect 37058 8324 37070 9100
rect 37012 8312 37070 8324
rect 37470 9100 37528 9112
rect 37470 8324 37482 9100
rect 37516 8324 37528 9100
rect 37470 8312 37528 8324
rect 37600 9100 37658 9112
rect 37600 8324 37612 9100
rect 37646 8324 37658 9100
rect 37600 8312 37658 8324
rect 38058 9100 38116 9112
rect 38058 8324 38070 9100
rect 38104 8324 38116 9100
rect 38058 8312 38116 8324
rect 38188 9100 38246 9112
rect 38188 8324 38200 9100
rect 38234 8324 38246 9100
rect 38188 8312 38246 8324
rect 38646 9100 38704 9112
rect 38646 8324 38658 9100
rect 38692 8324 38704 9100
rect 38646 8312 38704 8324
rect 23604 6654 23662 6666
rect 23604 5878 23616 6654
rect 23650 5878 23662 6654
rect 23604 5866 23662 5878
rect 23732 6654 23790 6666
rect 23732 5878 23744 6654
rect 23778 5878 23790 6654
rect 23732 5866 23790 5878
rect 23870 6654 23928 6666
rect 23870 5878 23882 6654
rect 23916 5878 23928 6654
rect 23870 5866 23928 5878
rect 23998 6654 24056 6666
rect 23998 5878 24010 6654
rect 24044 5878 24056 6654
rect 23998 5866 24056 5878
rect 24136 6654 24194 6666
rect 24136 5878 24148 6654
rect 24182 5878 24194 6654
rect 24136 5866 24194 5878
rect 24264 6654 24322 6666
rect 24264 5878 24276 6654
rect 24310 5878 24322 6654
rect 24264 5866 24322 5878
rect 24402 6654 24460 6666
rect 24402 5878 24414 6654
rect 24448 5878 24460 6654
rect 24402 5866 24460 5878
rect 24530 6654 24588 6666
rect 24530 5878 24542 6654
rect 24576 5878 24588 6654
rect 24530 5866 24588 5878
rect 24668 6654 24726 6666
rect 24668 5878 24680 6654
rect 24714 5878 24726 6654
rect 24668 5866 24726 5878
rect 24796 6654 24854 6666
rect 24796 5878 24808 6654
rect 24842 5878 24854 6654
rect 24796 5866 24854 5878
rect 24934 6654 24992 6666
rect 24934 5878 24946 6654
rect 24980 5878 24992 6654
rect 24934 5866 24992 5878
rect 25062 6654 25120 6666
rect 25062 5878 25074 6654
rect 25108 5878 25120 6654
rect 25062 5866 25120 5878
rect 25200 6654 25258 6666
rect 25200 5878 25212 6654
rect 25246 5878 25258 6654
rect 25200 5866 25258 5878
rect 25328 6654 25386 6666
rect 25328 5878 25340 6654
rect 25374 5878 25386 6654
rect 25328 5866 25386 5878
rect 25466 6654 25524 6666
rect 25466 5878 25478 6654
rect 25512 5878 25524 6654
rect 25466 5866 25524 5878
rect 25594 6654 25652 6666
rect 25594 5878 25606 6654
rect 25640 5878 25652 6654
rect 25594 5866 25652 5878
rect 23604 5644 23662 5656
rect 23604 4868 23616 5644
rect 23650 4868 23662 5644
rect 23604 4856 23662 4868
rect 23732 5644 23790 5656
rect 23732 4868 23744 5644
rect 23778 4868 23790 5644
rect 23732 4856 23790 4868
rect 23870 5644 23928 5656
rect 23870 4868 23882 5644
rect 23916 4868 23928 5644
rect 23870 4856 23928 4868
rect 23998 5644 24056 5656
rect 23998 4868 24010 5644
rect 24044 4868 24056 5644
rect 23998 4856 24056 4868
rect 24136 5644 24194 5656
rect 24136 4868 24148 5644
rect 24182 4868 24194 5644
rect 24136 4856 24194 4868
rect 24264 5644 24322 5656
rect 24264 4868 24276 5644
rect 24310 4868 24322 5644
rect 24264 4856 24322 4868
rect 24402 5644 24460 5656
rect 24402 4868 24414 5644
rect 24448 4868 24460 5644
rect 24402 4856 24460 4868
rect 24530 5644 24588 5656
rect 24530 4868 24542 5644
rect 24576 4868 24588 5644
rect 24530 4856 24588 4868
rect 24668 5644 24726 5656
rect 24668 4868 24680 5644
rect 24714 4868 24726 5644
rect 24668 4856 24726 4868
rect 24796 5644 24854 5656
rect 24796 4868 24808 5644
rect 24842 4868 24854 5644
rect 24796 4856 24854 4868
rect 24934 5644 24992 5656
rect 24934 4868 24946 5644
rect 24980 4868 24992 5644
rect 24934 4856 24992 4868
rect 25062 5644 25120 5656
rect 25062 4868 25074 5644
rect 25108 4868 25120 5644
rect 25062 4856 25120 4868
rect 25200 5644 25258 5656
rect 25200 4868 25212 5644
rect 25246 4868 25258 5644
rect 25200 4856 25258 4868
rect 25328 5644 25386 5656
rect 25328 4868 25340 5644
rect 25374 4868 25386 5644
rect 25328 4856 25386 4868
rect 25466 5644 25524 5656
rect 25466 4868 25478 5644
rect 25512 4868 25524 5644
rect 25466 4856 25524 4868
rect 25594 5644 25652 5656
rect 25594 4868 25606 5644
rect 25640 4868 25652 5644
rect 25594 4856 25652 4868
rect 23604 4634 23662 4646
rect 23604 3858 23616 4634
rect 23650 3858 23662 4634
rect 23604 3846 23662 3858
rect 23732 4634 23790 4646
rect 23732 3858 23744 4634
rect 23778 3858 23790 4634
rect 23732 3846 23790 3858
rect 23870 4634 23928 4646
rect 23870 3858 23882 4634
rect 23916 3858 23928 4634
rect 23870 3846 23928 3858
rect 23998 4634 24056 4646
rect 23998 3858 24010 4634
rect 24044 3858 24056 4634
rect 23998 3846 24056 3858
rect 24136 4634 24194 4646
rect 24136 3858 24148 4634
rect 24182 3858 24194 4634
rect 24136 3846 24194 3858
rect 24264 4634 24322 4646
rect 24264 3858 24276 4634
rect 24310 3858 24322 4634
rect 24264 3846 24322 3858
rect 24402 4634 24460 4646
rect 24402 3858 24414 4634
rect 24448 3858 24460 4634
rect 24402 3846 24460 3858
rect 24530 4634 24588 4646
rect 24530 3858 24542 4634
rect 24576 3858 24588 4634
rect 24530 3846 24588 3858
rect 24668 4634 24726 4646
rect 24668 3858 24680 4634
rect 24714 3858 24726 4634
rect 24668 3846 24726 3858
rect 24796 4634 24854 4646
rect 24796 3858 24808 4634
rect 24842 3858 24854 4634
rect 24796 3846 24854 3858
rect 24934 4634 24992 4646
rect 24934 3858 24946 4634
rect 24980 3858 24992 4634
rect 24934 3846 24992 3858
rect 25062 4634 25120 4646
rect 25062 3858 25074 4634
rect 25108 3858 25120 4634
rect 25062 3846 25120 3858
rect 25200 4634 25258 4646
rect 25200 3858 25212 4634
rect 25246 3858 25258 4634
rect 25200 3846 25258 3858
rect 25328 4634 25386 4646
rect 25328 3858 25340 4634
rect 25374 3858 25386 4634
rect 25328 3846 25386 3858
rect 25466 4634 25524 4646
rect 25466 3858 25478 4634
rect 25512 3858 25524 4634
rect 25466 3846 25524 3858
rect 25594 4634 25652 4646
rect 25594 3858 25606 4634
rect 25640 3858 25652 4634
rect 25594 3846 25652 3858
<< ndiffc >>
rect 19868 14542 19902 15118
rect 19996 14542 20030 15118
rect 20108 14542 20142 15118
rect 20236 14542 20270 15118
rect 20348 14542 20382 15118
rect 20476 14542 20510 15118
rect 20588 14542 20622 15118
rect 20716 14542 20750 15118
rect 20828 14542 20862 15118
rect 20956 14542 20990 15118
rect 21068 14542 21102 15118
rect 21196 14542 21230 15118
rect 21308 14542 21342 15118
rect 21436 14542 21470 15118
rect 21548 14542 21582 15118
rect 21676 14542 21710 15118
rect 21788 14542 21822 15118
rect 21916 14542 21950 15118
rect 22028 14542 22062 15118
rect 22156 14542 22190 15118
rect 22268 14542 22302 15118
rect 22396 14542 22430 15118
rect 22508 14542 22542 15118
rect 22636 14542 22670 15118
rect 22748 14542 22782 15118
rect 22876 14542 22910 15118
rect 22988 14542 23022 15118
rect 23116 14542 23150 15118
rect 23228 14542 23262 15118
rect 23356 14542 23390 15118
rect 23468 14542 23502 15118
rect 23596 14542 23630 15118
rect 23708 14542 23742 15118
rect 23836 14542 23870 15118
rect 23948 14542 23982 15118
rect 24076 14542 24110 15118
rect 24188 14542 24222 15118
rect 24316 14542 24350 15118
rect 24428 14542 24462 15118
rect 24556 14542 24590 15118
rect 24668 14542 24702 15118
rect 24796 14542 24830 15118
rect 24908 14542 24942 15118
rect 25036 14542 25070 15118
rect 25148 14542 25182 15118
rect 25276 14542 25310 15118
rect 25388 14542 25422 15118
rect 25516 14542 25550 15118
rect 25628 14542 25662 15118
rect 25756 14542 25790 15118
rect 25868 14542 25902 15118
rect 25996 14542 26030 15118
rect 26108 14542 26142 15118
rect 26236 14542 26270 15118
rect 26348 14542 26382 15118
rect 26476 14542 26510 15118
rect 26588 14542 26622 15118
rect 26716 14542 26750 15118
rect 26828 14542 26862 15118
rect 26956 14542 26990 15118
rect 27068 14542 27102 15118
rect 27196 14542 27230 15118
rect 27308 14542 27342 15118
rect 27436 14542 27470 15118
rect 27548 14542 27582 15118
rect 27676 14542 27710 15118
rect 27788 14542 27822 15118
rect 27916 14542 27950 15118
rect 28028 14542 28062 15118
rect 28156 14542 28190 15118
rect 28268 14542 28302 15118
rect 28396 14542 28430 15118
rect 28508 14542 28542 15118
rect 28636 14542 28670 15118
rect 28748 14542 28782 15118
rect 28876 14542 28910 15118
rect 28988 14542 29022 15118
rect 29116 14542 29150 15118
rect 29228 14542 29262 15118
rect 29356 14542 29390 15118
rect 19868 13734 19902 14310
rect 19996 13734 20030 14310
rect 20108 13734 20142 14310
rect 20236 13734 20270 14310
rect 20348 13734 20382 14310
rect 20476 13734 20510 14310
rect 20588 13734 20622 14310
rect 20716 13734 20750 14310
rect 20828 13734 20862 14310
rect 20956 13734 20990 14310
rect 21068 13734 21102 14310
rect 21196 13734 21230 14310
rect 21308 13734 21342 14310
rect 21436 13734 21470 14310
rect 21548 13734 21582 14310
rect 21676 13734 21710 14310
rect 21788 13734 21822 14310
rect 21916 13734 21950 14310
rect 22028 13734 22062 14310
rect 22156 13734 22190 14310
rect 22268 13734 22302 14310
rect 22396 13734 22430 14310
rect 22508 13734 22542 14310
rect 22636 13734 22670 14310
rect 22748 13734 22782 14310
rect 22876 13734 22910 14310
rect 22988 13734 23022 14310
rect 23116 13734 23150 14310
rect 23228 13734 23262 14310
rect 23356 13734 23390 14310
rect 23468 13734 23502 14310
rect 23596 13734 23630 14310
rect 23708 13734 23742 14310
rect 23836 13734 23870 14310
rect 23948 13734 23982 14310
rect 24076 13734 24110 14310
rect 24188 13734 24222 14310
rect 24316 13734 24350 14310
rect 24428 13734 24462 14310
rect 24556 13734 24590 14310
rect 24668 13734 24702 14310
rect 24796 13734 24830 14310
rect 24908 13734 24942 14310
rect 25036 13734 25070 14310
rect 25148 13734 25182 14310
rect 25276 13734 25310 14310
rect 25388 13734 25422 14310
rect 25516 13734 25550 14310
rect 25628 13734 25662 14310
rect 25756 13734 25790 14310
rect 25868 13734 25902 14310
rect 25996 13734 26030 14310
rect 26108 13734 26142 14310
rect 26236 13734 26270 14310
rect 26348 13734 26382 14310
rect 26476 13734 26510 14310
rect 26588 13734 26622 14310
rect 26716 13734 26750 14310
rect 26828 13734 26862 14310
rect 26956 13734 26990 14310
rect 27068 13734 27102 14310
rect 27196 13734 27230 14310
rect 27308 13734 27342 14310
rect 27436 13734 27470 14310
rect 27548 13734 27582 14310
rect 27676 13734 27710 14310
rect 27788 13734 27822 14310
rect 27916 13734 27950 14310
rect 28028 13734 28062 14310
rect 28156 13734 28190 14310
rect 28268 13734 28302 14310
rect 28396 13734 28430 14310
rect 28508 13734 28542 14310
rect 28636 13734 28670 14310
rect 28748 13734 28782 14310
rect 28876 13734 28910 14310
rect 28988 13734 29022 14310
rect 29116 13734 29150 14310
rect 29228 13734 29262 14310
rect 29356 13734 29390 14310
rect 24188 1886 24222 2462
rect 24316 1886 24350 2462
rect 24428 1886 24462 2462
rect 24556 1886 24590 2462
rect 24668 1886 24702 2462
rect 24796 1886 24830 2462
rect 24908 1886 24942 2462
rect 25036 1886 25070 2462
rect 24188 1078 24222 1654
rect 24316 1078 24350 1654
rect 24428 1078 24462 1654
rect 24556 1078 24590 1654
rect 24668 1078 24702 1654
rect 24796 1078 24830 1654
rect 24908 1078 24942 1654
rect 25036 1078 25070 1654
<< pdiffc >>
rect 10564 10324 10598 11100
rect 11022 10324 11056 11100
rect 11152 10324 11186 11100
rect 11610 10324 11644 11100
rect 11740 10324 11774 11100
rect 12198 10324 12232 11100
rect 12328 10324 12362 11100
rect 12786 10324 12820 11100
rect 12916 10324 12950 11100
rect 13374 10324 13408 11100
rect 13504 10324 13538 11100
rect 13962 10324 13996 11100
rect 14092 10324 14126 11100
rect 14550 10324 14584 11100
rect 14680 10324 14714 11100
rect 15138 10324 15172 11100
rect 15268 10324 15302 11100
rect 15726 10324 15760 11100
rect 15856 10324 15890 11100
rect 16314 10324 16348 11100
rect 16444 10324 16478 11100
rect 16902 10324 16936 11100
rect 17032 10324 17066 11100
rect 17490 10324 17524 11100
rect 17620 10324 17654 11100
rect 18078 10324 18112 11100
rect 18208 10324 18242 11100
rect 18666 10324 18700 11100
rect 18796 10324 18830 11100
rect 19254 10324 19288 11100
rect 19384 10324 19418 11100
rect 19842 10324 19876 11100
rect 19972 10324 20006 11100
rect 20430 10324 20464 11100
rect 20560 10324 20594 11100
rect 21018 10324 21052 11100
rect 21148 10324 21182 11100
rect 21606 10324 21640 11100
rect 21736 10324 21770 11100
rect 22194 10324 22228 11100
rect 22324 10324 22358 11100
rect 22782 10324 22816 11100
rect 22912 10324 22946 11100
rect 23370 10324 23404 11100
rect 23500 10324 23534 11100
rect 23958 10324 23992 11100
rect 24088 10324 24122 11100
rect 24546 10324 24580 11100
rect 24676 10324 24710 11100
rect 25134 10324 25168 11100
rect 25264 10324 25298 11100
rect 25722 10324 25756 11100
rect 25852 10324 25886 11100
rect 26310 10324 26344 11100
rect 26440 10324 26474 11100
rect 26898 10324 26932 11100
rect 27028 10324 27062 11100
rect 27486 10324 27520 11100
rect 27616 10324 27650 11100
rect 28074 10324 28108 11100
rect 28204 10324 28238 11100
rect 28662 10324 28696 11100
rect 28792 10324 28826 11100
rect 29250 10324 29284 11100
rect 29380 10324 29414 11100
rect 29838 10324 29872 11100
rect 29968 10324 30002 11100
rect 30426 10324 30460 11100
rect 30556 10324 30590 11100
rect 31014 10324 31048 11100
rect 31144 10324 31178 11100
rect 31602 10324 31636 11100
rect 31732 10324 31766 11100
rect 32190 10324 32224 11100
rect 32320 10324 32354 11100
rect 32778 10324 32812 11100
rect 32908 10324 32942 11100
rect 33366 10324 33400 11100
rect 33496 10324 33530 11100
rect 33954 10324 33988 11100
rect 34084 10324 34118 11100
rect 34542 10324 34576 11100
rect 34672 10324 34706 11100
rect 35130 10324 35164 11100
rect 35260 10324 35294 11100
rect 35718 10324 35752 11100
rect 35848 10324 35882 11100
rect 36306 10324 36340 11100
rect 36436 10324 36470 11100
rect 36894 10324 36928 11100
rect 37024 10324 37058 11100
rect 37482 10324 37516 11100
rect 37612 10324 37646 11100
rect 38070 10324 38104 11100
rect 38200 10324 38234 11100
rect 38658 10324 38692 11100
rect 10564 9324 10598 10100
rect 11022 9324 11056 10100
rect 11152 9324 11186 10100
rect 11610 9324 11644 10100
rect 11740 9324 11774 10100
rect 12198 9324 12232 10100
rect 12328 9324 12362 10100
rect 12786 9324 12820 10100
rect 12916 9324 12950 10100
rect 13374 9324 13408 10100
rect 13504 9324 13538 10100
rect 13962 9324 13996 10100
rect 14092 9324 14126 10100
rect 14550 9324 14584 10100
rect 14680 9324 14714 10100
rect 15138 9324 15172 10100
rect 15268 9324 15302 10100
rect 15726 9324 15760 10100
rect 15856 9324 15890 10100
rect 16314 9324 16348 10100
rect 16444 9324 16478 10100
rect 16902 9324 16936 10100
rect 17032 9324 17066 10100
rect 17490 9324 17524 10100
rect 17620 9324 17654 10100
rect 18078 9324 18112 10100
rect 18208 9324 18242 10100
rect 18666 9324 18700 10100
rect 18796 9324 18830 10100
rect 19254 9324 19288 10100
rect 19384 9324 19418 10100
rect 19842 9324 19876 10100
rect 19972 9324 20006 10100
rect 20430 9324 20464 10100
rect 20560 9324 20594 10100
rect 21018 9324 21052 10100
rect 21148 9324 21182 10100
rect 21606 9324 21640 10100
rect 21736 9324 21770 10100
rect 22194 9324 22228 10100
rect 22324 9324 22358 10100
rect 22782 9324 22816 10100
rect 22912 9324 22946 10100
rect 23370 9324 23404 10100
rect 23500 9324 23534 10100
rect 23958 9324 23992 10100
rect 24088 9324 24122 10100
rect 24546 9324 24580 10100
rect 24676 9324 24710 10100
rect 25134 9324 25168 10100
rect 25264 9324 25298 10100
rect 25722 9324 25756 10100
rect 25852 9324 25886 10100
rect 26310 9324 26344 10100
rect 26440 9324 26474 10100
rect 26898 9324 26932 10100
rect 27028 9324 27062 10100
rect 27486 9324 27520 10100
rect 27616 9324 27650 10100
rect 28074 9324 28108 10100
rect 28204 9324 28238 10100
rect 28662 9324 28696 10100
rect 28792 9324 28826 10100
rect 29250 9324 29284 10100
rect 29380 9324 29414 10100
rect 29838 9324 29872 10100
rect 29968 9324 30002 10100
rect 30426 9324 30460 10100
rect 30556 9324 30590 10100
rect 31014 9324 31048 10100
rect 31144 9324 31178 10100
rect 31602 9324 31636 10100
rect 31732 9324 31766 10100
rect 32190 9324 32224 10100
rect 32320 9324 32354 10100
rect 32778 9324 32812 10100
rect 32908 9324 32942 10100
rect 33366 9324 33400 10100
rect 33496 9324 33530 10100
rect 33954 9324 33988 10100
rect 34084 9324 34118 10100
rect 34542 9324 34576 10100
rect 34672 9324 34706 10100
rect 35130 9324 35164 10100
rect 35260 9324 35294 10100
rect 35718 9324 35752 10100
rect 35848 9324 35882 10100
rect 36306 9324 36340 10100
rect 36436 9324 36470 10100
rect 36894 9324 36928 10100
rect 37024 9324 37058 10100
rect 37482 9324 37516 10100
rect 37612 9324 37646 10100
rect 38070 9324 38104 10100
rect 38200 9324 38234 10100
rect 38658 9324 38692 10100
rect 10564 8324 10598 9100
rect 11022 8324 11056 9100
rect 11152 8324 11186 9100
rect 11610 8324 11644 9100
rect 11740 8324 11774 9100
rect 12198 8324 12232 9100
rect 12328 8324 12362 9100
rect 12786 8324 12820 9100
rect 12916 8324 12950 9100
rect 13374 8324 13408 9100
rect 13504 8324 13538 9100
rect 13962 8324 13996 9100
rect 14092 8324 14126 9100
rect 14550 8324 14584 9100
rect 14680 8324 14714 9100
rect 15138 8324 15172 9100
rect 15268 8324 15302 9100
rect 15726 8324 15760 9100
rect 15856 8324 15890 9100
rect 16314 8324 16348 9100
rect 16444 8324 16478 9100
rect 16902 8324 16936 9100
rect 17032 8324 17066 9100
rect 17490 8324 17524 9100
rect 17620 8324 17654 9100
rect 18078 8324 18112 9100
rect 18208 8324 18242 9100
rect 18666 8324 18700 9100
rect 18796 8324 18830 9100
rect 19254 8324 19288 9100
rect 19384 8324 19418 9100
rect 19842 8324 19876 9100
rect 19972 8324 20006 9100
rect 20430 8324 20464 9100
rect 20560 8324 20594 9100
rect 21018 8324 21052 9100
rect 21148 8324 21182 9100
rect 21606 8324 21640 9100
rect 21736 8324 21770 9100
rect 22194 8324 22228 9100
rect 22324 8324 22358 9100
rect 22782 8324 22816 9100
rect 22912 8324 22946 9100
rect 23370 8324 23404 9100
rect 23500 8324 23534 9100
rect 23958 8324 23992 9100
rect 24088 8324 24122 9100
rect 24546 8324 24580 9100
rect 24676 8324 24710 9100
rect 25134 8324 25168 9100
rect 25264 8324 25298 9100
rect 25722 8324 25756 9100
rect 25852 8324 25886 9100
rect 26310 8324 26344 9100
rect 26440 8324 26474 9100
rect 26898 8324 26932 9100
rect 27028 8324 27062 9100
rect 27486 8324 27520 9100
rect 27616 8324 27650 9100
rect 28074 8324 28108 9100
rect 28204 8324 28238 9100
rect 28662 8324 28696 9100
rect 28792 8324 28826 9100
rect 29250 8324 29284 9100
rect 29380 8324 29414 9100
rect 29838 8324 29872 9100
rect 29968 8324 30002 9100
rect 30426 8324 30460 9100
rect 30556 8324 30590 9100
rect 31014 8324 31048 9100
rect 31144 8324 31178 9100
rect 31602 8324 31636 9100
rect 31732 8324 31766 9100
rect 32190 8324 32224 9100
rect 32320 8324 32354 9100
rect 32778 8324 32812 9100
rect 32908 8324 32942 9100
rect 33366 8324 33400 9100
rect 33496 8324 33530 9100
rect 33954 8324 33988 9100
rect 34084 8324 34118 9100
rect 34542 8324 34576 9100
rect 34672 8324 34706 9100
rect 35130 8324 35164 9100
rect 35260 8324 35294 9100
rect 35718 8324 35752 9100
rect 35848 8324 35882 9100
rect 36306 8324 36340 9100
rect 36436 8324 36470 9100
rect 36894 8324 36928 9100
rect 37024 8324 37058 9100
rect 37482 8324 37516 9100
rect 37612 8324 37646 9100
rect 38070 8324 38104 9100
rect 38200 8324 38234 9100
rect 38658 8324 38692 9100
rect 23616 5878 23650 6654
rect 23744 5878 23778 6654
rect 23882 5878 23916 6654
rect 24010 5878 24044 6654
rect 24148 5878 24182 6654
rect 24276 5878 24310 6654
rect 24414 5878 24448 6654
rect 24542 5878 24576 6654
rect 24680 5878 24714 6654
rect 24808 5878 24842 6654
rect 24946 5878 24980 6654
rect 25074 5878 25108 6654
rect 25212 5878 25246 6654
rect 25340 5878 25374 6654
rect 25478 5878 25512 6654
rect 25606 5878 25640 6654
rect 23616 4868 23650 5644
rect 23744 4868 23778 5644
rect 23882 4868 23916 5644
rect 24010 4868 24044 5644
rect 24148 4868 24182 5644
rect 24276 4868 24310 5644
rect 24414 4868 24448 5644
rect 24542 4868 24576 5644
rect 24680 4868 24714 5644
rect 24808 4868 24842 5644
rect 24946 4868 24980 5644
rect 25074 4868 25108 5644
rect 25212 4868 25246 5644
rect 25340 4868 25374 5644
rect 25478 4868 25512 5644
rect 25606 4868 25640 5644
rect 23616 3858 23650 4634
rect 23744 3858 23778 4634
rect 23882 3858 23916 4634
rect 24010 3858 24044 4634
rect 24148 3858 24182 4634
rect 24276 3858 24310 4634
rect 24414 3858 24448 4634
rect 24542 3858 24576 4634
rect 24680 3858 24714 4634
rect 24808 3858 24842 4634
rect 24946 3858 24980 4634
rect 25074 3858 25108 4634
rect 25212 3858 25246 4634
rect 25340 3858 25374 4634
rect 25478 3858 25512 4634
rect 25606 3858 25640 4634
<< psubdiff >>
rect 30651 5255 30747 5289
rect 30885 5255 30981 5289
rect 30651 5193 30685 5255
rect 30947 5193 30981 5255
rect 30651 3639 30685 3701
rect 30947 3639 30981 3701
rect 30651 3605 30747 3639
rect 30885 3605 30981 3639
<< nsubdiff >>
rect 23230 7136 23264 7170
rect 25992 7136 26026 7170
rect 23230 3340 23264 3374
rect 25992 3340 26026 3374
<< psubdiffcont >>
rect 19610 15610 29648 15644
rect 19522 13296 19556 15576
rect 29702 13296 29736 15578
rect 19556 13208 29702 13242
rect 30747 5255 30885 5289
rect 30651 3701 30685 5193
rect 30947 3701 30981 5193
rect 30747 3605 30885 3639
rect 23988 2944 25198 2978
rect 23842 596 23876 2944
rect 25382 596 25416 2944
rect 24000 562 25210 596
<< nsubdiffcont >>
rect 10378 11510 38900 11544
rect 10218 7934 10252 11482
rect 39004 7968 39038 11516
rect 10336 7880 38950 7914
rect 23264 7136 25992 7170
rect 23230 3374 23264 7136
rect 25992 3374 26026 7136
rect 23264 3340 25992 3374
<< poly >>
rect 19914 15300 19984 15310
rect 19914 15168 19930 15300
rect 19968 15168 19984 15300
rect 19914 15130 19984 15168
rect 20154 15300 20224 15310
rect 20154 15168 20170 15300
rect 20208 15168 20224 15300
rect 20154 15130 20224 15168
rect 20394 15300 20464 15310
rect 20394 15168 20410 15300
rect 20448 15168 20464 15300
rect 20394 15130 20464 15168
rect 20634 15300 20704 15310
rect 20634 15168 20650 15300
rect 20688 15168 20704 15300
rect 20634 15130 20704 15168
rect 20874 15300 20944 15310
rect 20874 15168 20890 15300
rect 20928 15168 20944 15300
rect 20874 15130 20944 15168
rect 21114 15300 21184 15310
rect 21114 15168 21130 15300
rect 21168 15168 21184 15300
rect 21114 15130 21184 15168
rect 21354 15300 21424 15310
rect 21354 15168 21370 15300
rect 21408 15168 21424 15300
rect 21354 15130 21424 15168
rect 21594 15300 21664 15310
rect 21594 15168 21610 15300
rect 21648 15168 21664 15300
rect 21594 15130 21664 15168
rect 21834 15300 21904 15310
rect 21834 15168 21850 15300
rect 21888 15168 21904 15300
rect 21834 15130 21904 15168
rect 22074 15300 22144 15310
rect 22074 15168 22090 15300
rect 22128 15168 22144 15300
rect 22074 15130 22144 15168
rect 22314 15300 22384 15310
rect 22314 15168 22330 15300
rect 22368 15168 22384 15300
rect 22314 15130 22384 15168
rect 22554 15300 22624 15310
rect 22554 15168 22570 15300
rect 22608 15168 22624 15300
rect 22554 15130 22624 15168
rect 22794 15300 22864 15310
rect 22794 15168 22810 15300
rect 22848 15168 22864 15300
rect 22794 15130 22864 15168
rect 23034 15300 23104 15310
rect 23034 15168 23050 15300
rect 23088 15168 23104 15300
rect 23034 15130 23104 15168
rect 23274 15300 23344 15310
rect 23274 15168 23290 15300
rect 23328 15168 23344 15300
rect 23274 15130 23344 15168
rect 23514 15300 23584 15310
rect 23514 15168 23530 15300
rect 23568 15168 23584 15300
rect 23514 15130 23584 15168
rect 23754 15300 23824 15310
rect 23754 15168 23770 15300
rect 23808 15168 23824 15300
rect 23754 15130 23824 15168
rect 23994 15300 24064 15310
rect 23994 15168 24010 15300
rect 24048 15168 24064 15300
rect 23994 15130 24064 15168
rect 24234 15300 24304 15310
rect 24234 15168 24250 15300
rect 24288 15168 24304 15300
rect 24234 15130 24304 15168
rect 24474 15300 24544 15310
rect 24474 15168 24490 15300
rect 24528 15168 24544 15300
rect 24474 15130 24544 15168
rect 24714 15300 24784 15310
rect 24714 15168 24730 15300
rect 24768 15168 24784 15300
rect 24714 15130 24784 15168
rect 24954 15300 25024 15310
rect 24954 15168 24970 15300
rect 25008 15168 25024 15300
rect 24954 15130 25024 15168
rect 25194 15300 25264 15310
rect 25194 15168 25210 15300
rect 25248 15168 25264 15300
rect 25194 15130 25264 15168
rect 25434 15300 25504 15310
rect 25434 15168 25450 15300
rect 25488 15168 25504 15300
rect 25434 15130 25504 15168
rect 25674 15300 25744 15310
rect 25674 15168 25690 15300
rect 25728 15168 25744 15300
rect 25674 15130 25744 15168
rect 25914 15300 25984 15310
rect 25914 15168 25930 15300
rect 25968 15168 25984 15300
rect 25914 15130 25984 15168
rect 26154 15300 26224 15310
rect 26154 15168 26170 15300
rect 26208 15168 26224 15300
rect 26154 15130 26224 15168
rect 26394 15300 26464 15310
rect 26394 15168 26410 15300
rect 26448 15168 26464 15300
rect 26394 15130 26464 15168
rect 26634 15300 26704 15310
rect 26634 15168 26650 15300
rect 26688 15168 26704 15300
rect 26634 15130 26704 15168
rect 26874 15300 26944 15310
rect 26874 15168 26890 15300
rect 26928 15168 26944 15300
rect 26874 15130 26944 15168
rect 27114 15300 27184 15310
rect 27114 15168 27130 15300
rect 27168 15168 27184 15300
rect 27114 15130 27184 15168
rect 27354 15300 27424 15310
rect 27354 15168 27370 15300
rect 27408 15168 27424 15300
rect 27354 15130 27424 15168
rect 27594 15300 27664 15310
rect 27594 15168 27610 15300
rect 27648 15168 27664 15300
rect 27594 15130 27664 15168
rect 27834 15300 27904 15310
rect 27834 15168 27850 15300
rect 27888 15168 27904 15300
rect 27834 15130 27904 15168
rect 28074 15300 28144 15310
rect 28074 15168 28090 15300
rect 28128 15168 28144 15300
rect 28074 15130 28144 15168
rect 28314 15300 28384 15310
rect 28314 15168 28330 15300
rect 28368 15168 28384 15300
rect 28314 15130 28384 15168
rect 28554 15300 28624 15310
rect 28554 15168 28570 15300
rect 28608 15168 28624 15300
rect 28554 15130 28624 15168
rect 28794 15300 28864 15310
rect 28794 15168 28810 15300
rect 28848 15168 28864 15300
rect 28794 15130 28864 15168
rect 29034 15300 29104 15310
rect 29034 15168 29050 15300
rect 29088 15168 29104 15300
rect 29034 15130 29104 15168
rect 29274 15300 29344 15310
rect 29274 15168 29290 15300
rect 29328 15168 29344 15300
rect 29274 15130 29344 15168
rect 19914 14492 19984 14530
rect 19914 14360 19930 14492
rect 19968 14360 19984 14492
rect 19914 14322 19984 14360
rect 20154 14492 20224 14530
rect 20154 14360 20170 14492
rect 20208 14360 20224 14492
rect 20154 14322 20224 14360
rect 20394 14492 20464 14530
rect 20394 14360 20410 14492
rect 20448 14360 20464 14492
rect 20394 14322 20464 14360
rect 20634 14492 20704 14530
rect 20634 14360 20650 14492
rect 20688 14360 20704 14492
rect 20634 14322 20704 14360
rect 20874 14492 20944 14530
rect 20874 14360 20890 14492
rect 20928 14360 20944 14492
rect 20874 14322 20944 14360
rect 21114 14492 21184 14530
rect 21114 14360 21130 14492
rect 21168 14360 21184 14492
rect 21114 14322 21184 14360
rect 21354 14492 21424 14530
rect 21354 14360 21370 14492
rect 21408 14360 21424 14492
rect 21354 14322 21424 14360
rect 21594 14492 21664 14530
rect 21594 14360 21610 14492
rect 21648 14360 21664 14492
rect 21594 14322 21664 14360
rect 21834 14492 21904 14530
rect 21834 14360 21850 14492
rect 21888 14360 21904 14492
rect 21834 14322 21904 14360
rect 22074 14492 22144 14530
rect 22074 14360 22090 14492
rect 22128 14360 22144 14492
rect 22074 14322 22144 14360
rect 22314 14492 22384 14530
rect 22314 14360 22330 14492
rect 22368 14360 22384 14492
rect 22314 14322 22384 14360
rect 22554 14492 22624 14530
rect 22554 14360 22570 14492
rect 22608 14360 22624 14492
rect 22554 14322 22624 14360
rect 22794 14492 22864 14530
rect 22794 14360 22810 14492
rect 22848 14360 22864 14492
rect 22794 14322 22864 14360
rect 23034 14492 23104 14530
rect 23034 14360 23050 14492
rect 23088 14360 23104 14492
rect 23034 14322 23104 14360
rect 23274 14492 23344 14530
rect 23274 14360 23290 14492
rect 23328 14360 23344 14492
rect 23274 14322 23344 14360
rect 23514 14492 23584 14530
rect 23514 14360 23530 14492
rect 23568 14360 23584 14492
rect 23514 14322 23584 14360
rect 23754 14492 23824 14530
rect 23754 14360 23770 14492
rect 23808 14360 23824 14492
rect 23754 14322 23824 14360
rect 23994 14492 24064 14530
rect 23994 14360 24010 14492
rect 24048 14360 24064 14492
rect 23994 14322 24064 14360
rect 24234 14492 24304 14530
rect 24234 14360 24250 14492
rect 24288 14360 24304 14492
rect 24234 14322 24304 14360
rect 24474 14492 24544 14530
rect 24474 14360 24490 14492
rect 24528 14360 24544 14492
rect 24474 14322 24544 14360
rect 24714 14492 24784 14530
rect 24714 14360 24730 14492
rect 24768 14360 24784 14492
rect 24714 14322 24784 14360
rect 24954 14492 25024 14530
rect 24954 14360 24970 14492
rect 25008 14360 25024 14492
rect 24954 14322 25024 14360
rect 25194 14492 25264 14530
rect 25194 14360 25210 14492
rect 25248 14360 25264 14492
rect 25194 14322 25264 14360
rect 25434 14492 25504 14530
rect 25434 14360 25450 14492
rect 25488 14360 25504 14492
rect 25434 14322 25504 14360
rect 25674 14492 25744 14530
rect 25674 14360 25690 14492
rect 25728 14360 25744 14492
rect 25674 14322 25744 14360
rect 25914 14492 25984 14530
rect 25914 14360 25930 14492
rect 25968 14360 25984 14492
rect 25914 14322 25984 14360
rect 26154 14492 26224 14530
rect 26154 14360 26170 14492
rect 26208 14360 26224 14492
rect 26154 14322 26224 14360
rect 26394 14492 26464 14530
rect 26394 14360 26410 14492
rect 26448 14360 26464 14492
rect 26394 14322 26464 14360
rect 26634 14492 26704 14530
rect 26634 14360 26650 14492
rect 26688 14360 26704 14492
rect 26634 14322 26704 14360
rect 26874 14492 26944 14530
rect 26874 14360 26890 14492
rect 26928 14360 26944 14492
rect 26874 14322 26944 14360
rect 27114 14492 27184 14530
rect 27114 14360 27130 14492
rect 27168 14360 27184 14492
rect 27114 14322 27184 14360
rect 27354 14492 27424 14530
rect 27354 14360 27370 14492
rect 27408 14360 27424 14492
rect 27354 14322 27424 14360
rect 27594 14492 27664 14530
rect 27594 14360 27610 14492
rect 27648 14360 27664 14492
rect 27594 14322 27664 14360
rect 27834 14492 27904 14530
rect 27834 14360 27850 14492
rect 27888 14360 27904 14492
rect 27834 14322 27904 14360
rect 28074 14492 28144 14530
rect 28074 14360 28090 14492
rect 28128 14360 28144 14492
rect 28074 14322 28144 14360
rect 28314 14492 28384 14530
rect 28314 14360 28330 14492
rect 28368 14360 28384 14492
rect 28314 14322 28384 14360
rect 28554 14492 28624 14530
rect 28554 14360 28570 14492
rect 28608 14360 28624 14492
rect 28554 14322 28624 14360
rect 28794 14492 28864 14530
rect 28794 14360 28810 14492
rect 28848 14360 28864 14492
rect 28794 14322 28864 14360
rect 29034 14492 29104 14530
rect 29034 14360 29050 14492
rect 29088 14360 29104 14492
rect 29034 14322 29104 14360
rect 29274 14492 29344 14530
rect 29274 14360 29290 14492
rect 29328 14360 29344 14492
rect 29274 14322 29344 14360
rect 19914 13684 19984 13722
rect 19914 13552 19930 13684
rect 19968 13552 19984 13684
rect 19914 13542 19984 13552
rect 20154 13684 20224 13722
rect 20154 13552 20170 13684
rect 20208 13552 20224 13684
rect 20154 13542 20224 13552
rect 20394 13684 20464 13722
rect 20394 13552 20410 13684
rect 20448 13552 20464 13684
rect 20394 13542 20464 13552
rect 20634 13684 20704 13722
rect 20634 13552 20650 13684
rect 20688 13552 20704 13684
rect 20634 13542 20704 13552
rect 20874 13684 20944 13722
rect 20874 13552 20890 13684
rect 20928 13552 20944 13684
rect 20874 13542 20944 13552
rect 21114 13684 21184 13722
rect 21114 13552 21130 13684
rect 21168 13552 21184 13684
rect 21114 13542 21184 13552
rect 21354 13684 21424 13722
rect 21354 13552 21370 13684
rect 21408 13552 21424 13684
rect 21354 13542 21424 13552
rect 21594 13684 21664 13722
rect 21594 13552 21610 13684
rect 21648 13552 21664 13684
rect 21594 13542 21664 13552
rect 21834 13684 21904 13722
rect 21834 13552 21850 13684
rect 21888 13552 21904 13684
rect 21834 13542 21904 13552
rect 22074 13684 22144 13722
rect 22074 13552 22090 13684
rect 22128 13552 22144 13684
rect 22074 13542 22144 13552
rect 22314 13684 22384 13722
rect 22314 13552 22330 13684
rect 22368 13552 22384 13684
rect 22314 13542 22384 13552
rect 22554 13684 22624 13722
rect 22554 13552 22570 13684
rect 22608 13552 22624 13684
rect 22554 13542 22624 13552
rect 22794 13684 22864 13722
rect 22794 13552 22810 13684
rect 22848 13552 22864 13684
rect 22794 13542 22864 13552
rect 23034 13684 23104 13722
rect 23034 13552 23050 13684
rect 23088 13552 23104 13684
rect 23034 13542 23104 13552
rect 23274 13684 23344 13722
rect 23274 13552 23290 13684
rect 23328 13552 23344 13684
rect 23274 13542 23344 13552
rect 23514 13684 23584 13722
rect 23514 13552 23530 13684
rect 23568 13552 23584 13684
rect 23514 13542 23584 13552
rect 23754 13684 23824 13722
rect 23754 13552 23770 13684
rect 23808 13552 23824 13684
rect 23754 13542 23824 13552
rect 23994 13684 24064 13722
rect 23994 13552 24010 13684
rect 24048 13552 24064 13684
rect 23994 13542 24064 13552
rect 24234 13684 24304 13722
rect 24234 13552 24250 13684
rect 24288 13552 24304 13684
rect 24234 13542 24304 13552
rect 24474 13684 24544 13722
rect 24474 13552 24490 13684
rect 24528 13552 24544 13684
rect 24474 13542 24544 13552
rect 24714 13684 24784 13722
rect 24714 13552 24730 13684
rect 24768 13552 24784 13684
rect 24714 13542 24784 13552
rect 24954 13684 25024 13722
rect 24954 13552 24970 13684
rect 25008 13552 25024 13684
rect 24954 13542 25024 13552
rect 25194 13684 25264 13722
rect 25194 13552 25210 13684
rect 25248 13552 25264 13684
rect 25194 13542 25264 13552
rect 25434 13684 25504 13722
rect 25434 13552 25450 13684
rect 25488 13552 25504 13684
rect 25434 13542 25504 13552
rect 25674 13684 25744 13722
rect 25674 13552 25690 13684
rect 25728 13552 25744 13684
rect 25674 13542 25744 13552
rect 25914 13684 25984 13722
rect 25914 13552 25930 13684
rect 25968 13552 25984 13684
rect 25914 13542 25984 13552
rect 26154 13684 26224 13722
rect 26154 13552 26170 13684
rect 26208 13552 26224 13684
rect 26154 13542 26224 13552
rect 26394 13684 26464 13722
rect 26394 13552 26410 13684
rect 26448 13552 26464 13684
rect 26394 13542 26464 13552
rect 26634 13684 26704 13722
rect 26634 13552 26650 13684
rect 26688 13552 26704 13684
rect 26634 13542 26704 13552
rect 26874 13684 26944 13722
rect 26874 13552 26890 13684
rect 26928 13552 26944 13684
rect 26874 13542 26944 13552
rect 27114 13684 27184 13722
rect 27114 13552 27130 13684
rect 27168 13552 27184 13684
rect 27114 13542 27184 13552
rect 27354 13684 27424 13722
rect 27354 13552 27370 13684
rect 27408 13552 27424 13684
rect 27354 13542 27424 13552
rect 27594 13684 27664 13722
rect 27594 13552 27610 13684
rect 27648 13552 27664 13684
rect 27594 13542 27664 13552
rect 27834 13684 27904 13722
rect 27834 13552 27850 13684
rect 27888 13552 27904 13684
rect 27834 13542 27904 13552
rect 28074 13684 28144 13722
rect 28074 13552 28090 13684
rect 28128 13552 28144 13684
rect 28074 13542 28144 13552
rect 28314 13684 28384 13722
rect 28314 13552 28330 13684
rect 28368 13552 28384 13684
rect 28314 13542 28384 13552
rect 28554 13684 28624 13722
rect 28554 13552 28570 13684
rect 28608 13552 28624 13684
rect 28554 13542 28624 13552
rect 28794 13684 28864 13722
rect 28794 13552 28810 13684
rect 28848 13552 28864 13684
rect 28794 13542 28864 13552
rect 29034 13684 29104 13722
rect 29034 13552 29050 13684
rect 29088 13552 29104 13684
rect 29034 13542 29104 13552
rect 29274 13684 29344 13722
rect 29274 13552 29290 13684
rect 29328 13552 29344 13684
rect 29274 13542 29344 13552
rect 10610 11193 11010 11209
rect 10610 11159 10626 11193
rect 10994 11159 11010 11193
rect 10610 11112 11010 11159
rect 11198 11193 11598 11209
rect 11198 11159 11214 11193
rect 11582 11159 11598 11193
rect 11198 11112 11598 11159
rect 11786 11193 12186 11209
rect 11786 11159 11802 11193
rect 12170 11159 12186 11193
rect 11786 11112 12186 11159
rect 12374 11193 12774 11209
rect 12374 11159 12390 11193
rect 12758 11159 12774 11193
rect 12374 11112 12774 11159
rect 12962 11193 13362 11209
rect 12962 11159 12978 11193
rect 13346 11159 13362 11193
rect 12962 11112 13362 11159
rect 13550 11193 13950 11209
rect 13550 11159 13566 11193
rect 13934 11159 13950 11193
rect 13550 11112 13950 11159
rect 14138 11193 14538 11209
rect 14138 11159 14154 11193
rect 14522 11159 14538 11193
rect 14138 11112 14538 11159
rect 14726 11193 15126 11209
rect 14726 11159 14742 11193
rect 15110 11159 15126 11193
rect 14726 11112 15126 11159
rect 15314 11193 15714 11209
rect 15314 11159 15330 11193
rect 15698 11159 15714 11193
rect 15314 11112 15714 11159
rect 15902 11193 16302 11209
rect 15902 11159 15918 11193
rect 16286 11159 16302 11193
rect 15902 11112 16302 11159
rect 16490 11193 16890 11209
rect 16490 11159 16506 11193
rect 16874 11159 16890 11193
rect 16490 11112 16890 11159
rect 17078 11193 17478 11209
rect 17078 11159 17094 11193
rect 17462 11159 17478 11193
rect 17078 11112 17478 11159
rect 17666 11193 18066 11209
rect 17666 11159 17682 11193
rect 18050 11159 18066 11193
rect 17666 11112 18066 11159
rect 18254 11193 18654 11209
rect 18254 11159 18270 11193
rect 18638 11159 18654 11193
rect 18254 11112 18654 11159
rect 18842 11193 19242 11209
rect 18842 11159 18858 11193
rect 19226 11159 19242 11193
rect 18842 11112 19242 11159
rect 19430 11193 19830 11209
rect 19430 11159 19446 11193
rect 19814 11159 19830 11193
rect 19430 11112 19830 11159
rect 20018 11193 20418 11209
rect 20018 11159 20034 11193
rect 20402 11159 20418 11193
rect 20018 11112 20418 11159
rect 20606 11193 21006 11209
rect 20606 11159 20622 11193
rect 20990 11159 21006 11193
rect 20606 11112 21006 11159
rect 21194 11193 21594 11209
rect 21194 11159 21210 11193
rect 21578 11159 21594 11193
rect 21194 11112 21594 11159
rect 21782 11193 22182 11209
rect 21782 11159 21798 11193
rect 22166 11159 22182 11193
rect 21782 11112 22182 11159
rect 22370 11193 22770 11209
rect 22370 11159 22386 11193
rect 22754 11159 22770 11193
rect 22370 11112 22770 11159
rect 22958 11193 23358 11209
rect 22958 11159 22974 11193
rect 23342 11159 23358 11193
rect 22958 11112 23358 11159
rect 23546 11193 23946 11209
rect 23546 11159 23562 11193
rect 23930 11159 23946 11193
rect 23546 11112 23946 11159
rect 24134 11193 24534 11209
rect 24134 11159 24150 11193
rect 24518 11159 24534 11193
rect 24134 11112 24534 11159
rect 24722 11193 25122 11209
rect 24722 11159 24738 11193
rect 25106 11159 25122 11193
rect 24722 11112 25122 11159
rect 25310 11193 25710 11209
rect 25310 11159 25326 11193
rect 25694 11159 25710 11193
rect 25310 11112 25710 11159
rect 25898 11193 26298 11209
rect 25898 11159 25914 11193
rect 26282 11159 26298 11193
rect 25898 11112 26298 11159
rect 26486 11193 26886 11209
rect 26486 11159 26502 11193
rect 26870 11159 26886 11193
rect 26486 11112 26886 11159
rect 27074 11193 27474 11209
rect 27074 11159 27090 11193
rect 27458 11159 27474 11193
rect 27074 11112 27474 11159
rect 27662 11193 28062 11209
rect 27662 11159 27678 11193
rect 28046 11159 28062 11193
rect 27662 11112 28062 11159
rect 28250 11193 28650 11209
rect 28250 11159 28266 11193
rect 28634 11159 28650 11193
rect 28250 11112 28650 11159
rect 28838 11193 29238 11209
rect 28838 11159 28854 11193
rect 29222 11159 29238 11193
rect 28838 11112 29238 11159
rect 29426 11193 29826 11209
rect 29426 11159 29442 11193
rect 29810 11159 29826 11193
rect 29426 11112 29826 11159
rect 30014 11193 30414 11209
rect 30014 11159 30030 11193
rect 30398 11159 30414 11193
rect 30014 11112 30414 11159
rect 30602 11193 31002 11209
rect 30602 11159 30618 11193
rect 30986 11159 31002 11193
rect 30602 11112 31002 11159
rect 31190 11193 31590 11209
rect 31190 11159 31206 11193
rect 31574 11159 31590 11193
rect 31190 11112 31590 11159
rect 31778 11193 32178 11209
rect 31778 11159 31794 11193
rect 32162 11159 32178 11193
rect 31778 11112 32178 11159
rect 32366 11193 32766 11209
rect 32366 11159 32382 11193
rect 32750 11159 32766 11193
rect 32366 11112 32766 11159
rect 32954 11193 33354 11209
rect 32954 11159 32970 11193
rect 33338 11159 33354 11193
rect 32954 11112 33354 11159
rect 33542 11193 33942 11209
rect 33542 11159 33558 11193
rect 33926 11159 33942 11193
rect 33542 11112 33942 11159
rect 34130 11193 34530 11209
rect 34130 11159 34146 11193
rect 34514 11159 34530 11193
rect 34130 11112 34530 11159
rect 34718 11193 35118 11209
rect 34718 11159 34734 11193
rect 35102 11159 35118 11193
rect 34718 11112 35118 11159
rect 35306 11193 35706 11209
rect 35306 11159 35322 11193
rect 35690 11159 35706 11193
rect 35306 11112 35706 11159
rect 35894 11193 36294 11209
rect 35894 11159 35910 11193
rect 36278 11159 36294 11193
rect 35894 11112 36294 11159
rect 36482 11193 36882 11209
rect 36482 11159 36498 11193
rect 36866 11159 36882 11193
rect 36482 11112 36882 11159
rect 37070 11193 37470 11209
rect 37070 11159 37086 11193
rect 37454 11159 37470 11193
rect 37070 11112 37470 11159
rect 37658 11193 38058 11209
rect 37658 11159 37674 11193
rect 38042 11159 38058 11193
rect 37658 11112 38058 11159
rect 38246 11193 38646 11209
rect 38246 11159 38262 11193
rect 38630 11159 38646 11193
rect 38246 11112 38646 11159
rect 10610 10265 11010 10312
rect 10610 10231 10626 10265
rect 10994 10231 11010 10265
rect 10610 10193 11010 10231
rect 10610 10159 10626 10193
rect 10994 10159 11010 10193
rect 10610 10112 11010 10159
rect 11198 10265 11598 10312
rect 11198 10231 11214 10265
rect 11582 10231 11598 10265
rect 11198 10193 11598 10231
rect 11198 10159 11214 10193
rect 11582 10159 11598 10193
rect 11198 10112 11598 10159
rect 11786 10265 12186 10312
rect 11786 10231 11802 10265
rect 12170 10231 12186 10265
rect 11786 10193 12186 10231
rect 11786 10159 11802 10193
rect 12170 10159 12186 10193
rect 11786 10112 12186 10159
rect 12374 10265 12774 10312
rect 12374 10231 12390 10265
rect 12758 10231 12774 10265
rect 12374 10193 12774 10231
rect 12374 10159 12390 10193
rect 12758 10159 12774 10193
rect 12374 10112 12774 10159
rect 12962 10265 13362 10312
rect 12962 10231 12978 10265
rect 13346 10231 13362 10265
rect 12962 10193 13362 10231
rect 12962 10159 12978 10193
rect 13346 10159 13362 10193
rect 12962 10112 13362 10159
rect 13550 10265 13950 10312
rect 13550 10231 13566 10265
rect 13934 10231 13950 10265
rect 13550 10193 13950 10231
rect 13550 10159 13566 10193
rect 13934 10159 13950 10193
rect 13550 10112 13950 10159
rect 14138 10265 14538 10312
rect 14138 10231 14154 10265
rect 14522 10231 14538 10265
rect 14138 10193 14538 10231
rect 14138 10159 14154 10193
rect 14522 10159 14538 10193
rect 14138 10112 14538 10159
rect 14726 10265 15126 10312
rect 14726 10231 14742 10265
rect 15110 10231 15126 10265
rect 14726 10193 15126 10231
rect 14726 10159 14742 10193
rect 15110 10159 15126 10193
rect 14726 10112 15126 10159
rect 15314 10265 15714 10312
rect 15314 10231 15330 10265
rect 15698 10231 15714 10265
rect 15314 10193 15714 10231
rect 15314 10159 15330 10193
rect 15698 10159 15714 10193
rect 15314 10112 15714 10159
rect 15902 10265 16302 10312
rect 15902 10231 15918 10265
rect 16286 10231 16302 10265
rect 15902 10193 16302 10231
rect 15902 10159 15918 10193
rect 16286 10159 16302 10193
rect 15902 10112 16302 10159
rect 16490 10265 16890 10312
rect 16490 10231 16506 10265
rect 16874 10231 16890 10265
rect 16490 10193 16890 10231
rect 16490 10159 16506 10193
rect 16874 10159 16890 10193
rect 16490 10112 16890 10159
rect 17078 10265 17478 10312
rect 17078 10231 17094 10265
rect 17462 10231 17478 10265
rect 17078 10193 17478 10231
rect 17078 10159 17094 10193
rect 17462 10159 17478 10193
rect 17078 10112 17478 10159
rect 17666 10265 18066 10312
rect 17666 10231 17682 10265
rect 18050 10231 18066 10265
rect 17666 10193 18066 10231
rect 17666 10159 17682 10193
rect 18050 10159 18066 10193
rect 17666 10112 18066 10159
rect 18254 10265 18654 10312
rect 18254 10231 18270 10265
rect 18638 10231 18654 10265
rect 18254 10193 18654 10231
rect 18254 10159 18270 10193
rect 18638 10159 18654 10193
rect 18254 10112 18654 10159
rect 18842 10265 19242 10312
rect 18842 10231 18858 10265
rect 19226 10231 19242 10265
rect 18842 10193 19242 10231
rect 18842 10159 18858 10193
rect 19226 10159 19242 10193
rect 18842 10112 19242 10159
rect 19430 10265 19830 10312
rect 19430 10231 19446 10265
rect 19814 10231 19830 10265
rect 19430 10193 19830 10231
rect 19430 10159 19446 10193
rect 19814 10159 19830 10193
rect 19430 10112 19830 10159
rect 20018 10265 20418 10312
rect 20018 10231 20034 10265
rect 20402 10231 20418 10265
rect 20018 10193 20418 10231
rect 20018 10159 20034 10193
rect 20402 10159 20418 10193
rect 20018 10112 20418 10159
rect 20606 10265 21006 10312
rect 20606 10231 20622 10265
rect 20990 10231 21006 10265
rect 20606 10193 21006 10231
rect 20606 10159 20622 10193
rect 20990 10159 21006 10193
rect 20606 10112 21006 10159
rect 21194 10265 21594 10312
rect 21194 10231 21210 10265
rect 21578 10231 21594 10265
rect 21194 10193 21594 10231
rect 21194 10159 21210 10193
rect 21578 10159 21594 10193
rect 21194 10112 21594 10159
rect 21782 10265 22182 10312
rect 21782 10231 21798 10265
rect 22166 10231 22182 10265
rect 21782 10193 22182 10231
rect 21782 10159 21798 10193
rect 22166 10159 22182 10193
rect 21782 10112 22182 10159
rect 22370 10265 22770 10312
rect 22370 10231 22386 10265
rect 22754 10231 22770 10265
rect 22370 10193 22770 10231
rect 22370 10159 22386 10193
rect 22754 10159 22770 10193
rect 22370 10112 22770 10159
rect 22958 10265 23358 10312
rect 22958 10231 22974 10265
rect 23342 10231 23358 10265
rect 22958 10193 23358 10231
rect 22958 10159 22974 10193
rect 23342 10159 23358 10193
rect 22958 10112 23358 10159
rect 23546 10265 23946 10312
rect 23546 10231 23562 10265
rect 23930 10231 23946 10265
rect 23546 10193 23946 10231
rect 23546 10159 23562 10193
rect 23930 10159 23946 10193
rect 23546 10112 23946 10159
rect 24134 10265 24534 10312
rect 24134 10231 24150 10265
rect 24518 10231 24534 10265
rect 24134 10193 24534 10231
rect 24134 10159 24150 10193
rect 24518 10159 24534 10193
rect 24134 10112 24534 10159
rect 24722 10265 25122 10312
rect 24722 10231 24738 10265
rect 25106 10231 25122 10265
rect 24722 10193 25122 10231
rect 24722 10159 24738 10193
rect 25106 10159 25122 10193
rect 24722 10112 25122 10159
rect 25310 10265 25710 10312
rect 25310 10231 25326 10265
rect 25694 10231 25710 10265
rect 25310 10193 25710 10231
rect 25310 10159 25326 10193
rect 25694 10159 25710 10193
rect 25310 10112 25710 10159
rect 25898 10265 26298 10312
rect 25898 10231 25914 10265
rect 26282 10231 26298 10265
rect 25898 10193 26298 10231
rect 25898 10159 25914 10193
rect 26282 10159 26298 10193
rect 25898 10112 26298 10159
rect 26486 10265 26886 10312
rect 26486 10231 26502 10265
rect 26870 10231 26886 10265
rect 26486 10193 26886 10231
rect 26486 10159 26502 10193
rect 26870 10159 26886 10193
rect 26486 10112 26886 10159
rect 27074 10265 27474 10312
rect 27074 10231 27090 10265
rect 27458 10231 27474 10265
rect 27074 10193 27474 10231
rect 27074 10159 27090 10193
rect 27458 10159 27474 10193
rect 27074 10112 27474 10159
rect 27662 10265 28062 10312
rect 27662 10231 27678 10265
rect 28046 10231 28062 10265
rect 27662 10193 28062 10231
rect 27662 10159 27678 10193
rect 28046 10159 28062 10193
rect 27662 10112 28062 10159
rect 28250 10265 28650 10312
rect 28250 10231 28266 10265
rect 28634 10231 28650 10265
rect 28250 10193 28650 10231
rect 28250 10159 28266 10193
rect 28634 10159 28650 10193
rect 28250 10112 28650 10159
rect 28838 10265 29238 10312
rect 28838 10231 28854 10265
rect 29222 10231 29238 10265
rect 28838 10193 29238 10231
rect 28838 10159 28854 10193
rect 29222 10159 29238 10193
rect 28838 10112 29238 10159
rect 29426 10265 29826 10312
rect 29426 10231 29442 10265
rect 29810 10231 29826 10265
rect 29426 10193 29826 10231
rect 29426 10159 29442 10193
rect 29810 10159 29826 10193
rect 29426 10112 29826 10159
rect 30014 10265 30414 10312
rect 30014 10231 30030 10265
rect 30398 10231 30414 10265
rect 30014 10193 30414 10231
rect 30014 10159 30030 10193
rect 30398 10159 30414 10193
rect 30014 10112 30414 10159
rect 30602 10265 31002 10312
rect 30602 10231 30618 10265
rect 30986 10231 31002 10265
rect 30602 10193 31002 10231
rect 30602 10159 30618 10193
rect 30986 10159 31002 10193
rect 30602 10112 31002 10159
rect 31190 10265 31590 10312
rect 31190 10231 31206 10265
rect 31574 10231 31590 10265
rect 31190 10193 31590 10231
rect 31190 10159 31206 10193
rect 31574 10159 31590 10193
rect 31190 10112 31590 10159
rect 31778 10265 32178 10312
rect 31778 10231 31794 10265
rect 32162 10231 32178 10265
rect 31778 10193 32178 10231
rect 31778 10159 31794 10193
rect 32162 10159 32178 10193
rect 31778 10112 32178 10159
rect 32366 10265 32766 10312
rect 32366 10231 32382 10265
rect 32750 10231 32766 10265
rect 32366 10193 32766 10231
rect 32366 10159 32382 10193
rect 32750 10159 32766 10193
rect 32366 10112 32766 10159
rect 32954 10265 33354 10312
rect 32954 10231 32970 10265
rect 33338 10231 33354 10265
rect 32954 10193 33354 10231
rect 32954 10159 32970 10193
rect 33338 10159 33354 10193
rect 32954 10112 33354 10159
rect 33542 10265 33942 10312
rect 33542 10231 33558 10265
rect 33926 10231 33942 10265
rect 33542 10193 33942 10231
rect 33542 10159 33558 10193
rect 33926 10159 33942 10193
rect 33542 10112 33942 10159
rect 34130 10265 34530 10312
rect 34130 10231 34146 10265
rect 34514 10231 34530 10265
rect 34130 10193 34530 10231
rect 34130 10159 34146 10193
rect 34514 10159 34530 10193
rect 34130 10112 34530 10159
rect 34718 10265 35118 10312
rect 34718 10231 34734 10265
rect 35102 10231 35118 10265
rect 34718 10193 35118 10231
rect 34718 10159 34734 10193
rect 35102 10159 35118 10193
rect 34718 10112 35118 10159
rect 35306 10265 35706 10312
rect 35306 10231 35322 10265
rect 35690 10231 35706 10265
rect 35306 10193 35706 10231
rect 35306 10159 35322 10193
rect 35690 10159 35706 10193
rect 35306 10112 35706 10159
rect 35894 10265 36294 10312
rect 35894 10231 35910 10265
rect 36278 10231 36294 10265
rect 35894 10193 36294 10231
rect 35894 10159 35910 10193
rect 36278 10159 36294 10193
rect 35894 10112 36294 10159
rect 36482 10265 36882 10312
rect 36482 10231 36498 10265
rect 36866 10231 36882 10265
rect 36482 10193 36882 10231
rect 36482 10159 36498 10193
rect 36866 10159 36882 10193
rect 36482 10112 36882 10159
rect 37070 10265 37470 10312
rect 37070 10231 37086 10265
rect 37454 10231 37470 10265
rect 37070 10193 37470 10231
rect 37070 10159 37086 10193
rect 37454 10159 37470 10193
rect 37070 10112 37470 10159
rect 37658 10265 38058 10312
rect 37658 10231 37674 10265
rect 38042 10231 38058 10265
rect 37658 10193 38058 10231
rect 37658 10159 37674 10193
rect 38042 10159 38058 10193
rect 37658 10112 38058 10159
rect 38246 10265 38646 10312
rect 38246 10231 38262 10265
rect 38630 10231 38646 10265
rect 38246 10193 38646 10231
rect 38246 10159 38262 10193
rect 38630 10159 38646 10193
rect 38246 10112 38646 10159
rect 10610 9265 11010 9312
rect 10610 9231 10626 9265
rect 10994 9231 11010 9265
rect 10610 9193 11010 9231
rect 10610 9159 10626 9193
rect 10994 9159 11010 9193
rect 10610 9112 11010 9159
rect 11198 9265 11598 9312
rect 11198 9231 11214 9265
rect 11582 9231 11598 9265
rect 11198 9193 11598 9231
rect 11198 9159 11214 9193
rect 11582 9159 11598 9193
rect 11198 9112 11598 9159
rect 11786 9265 12186 9312
rect 11786 9231 11802 9265
rect 12170 9231 12186 9265
rect 11786 9193 12186 9231
rect 11786 9159 11802 9193
rect 12170 9159 12186 9193
rect 11786 9112 12186 9159
rect 12374 9265 12774 9312
rect 12374 9231 12390 9265
rect 12758 9231 12774 9265
rect 12374 9193 12774 9231
rect 12374 9159 12390 9193
rect 12758 9159 12774 9193
rect 12374 9112 12774 9159
rect 12962 9265 13362 9312
rect 12962 9231 12978 9265
rect 13346 9231 13362 9265
rect 12962 9193 13362 9231
rect 12962 9159 12978 9193
rect 13346 9159 13362 9193
rect 12962 9112 13362 9159
rect 13550 9265 13950 9312
rect 13550 9231 13566 9265
rect 13934 9231 13950 9265
rect 13550 9193 13950 9231
rect 13550 9159 13566 9193
rect 13934 9159 13950 9193
rect 13550 9112 13950 9159
rect 14138 9265 14538 9312
rect 14138 9231 14154 9265
rect 14522 9231 14538 9265
rect 14138 9193 14538 9231
rect 14138 9159 14154 9193
rect 14522 9159 14538 9193
rect 14138 9112 14538 9159
rect 14726 9265 15126 9312
rect 14726 9231 14742 9265
rect 15110 9231 15126 9265
rect 14726 9193 15126 9231
rect 14726 9159 14742 9193
rect 15110 9159 15126 9193
rect 14726 9112 15126 9159
rect 15314 9265 15714 9312
rect 15314 9231 15330 9265
rect 15698 9231 15714 9265
rect 15314 9193 15714 9231
rect 15314 9159 15330 9193
rect 15698 9159 15714 9193
rect 15314 9112 15714 9159
rect 15902 9265 16302 9312
rect 15902 9231 15918 9265
rect 16286 9231 16302 9265
rect 15902 9193 16302 9231
rect 15902 9159 15918 9193
rect 16286 9159 16302 9193
rect 15902 9112 16302 9159
rect 16490 9265 16890 9312
rect 16490 9231 16506 9265
rect 16874 9231 16890 9265
rect 16490 9193 16890 9231
rect 16490 9159 16506 9193
rect 16874 9159 16890 9193
rect 16490 9112 16890 9159
rect 17078 9265 17478 9312
rect 17078 9231 17094 9265
rect 17462 9231 17478 9265
rect 17078 9193 17478 9231
rect 17078 9159 17094 9193
rect 17462 9159 17478 9193
rect 17078 9112 17478 9159
rect 17666 9265 18066 9312
rect 17666 9231 17682 9265
rect 18050 9231 18066 9265
rect 17666 9193 18066 9231
rect 17666 9159 17682 9193
rect 18050 9159 18066 9193
rect 17666 9112 18066 9159
rect 18254 9265 18654 9312
rect 18254 9231 18270 9265
rect 18638 9231 18654 9265
rect 18254 9193 18654 9231
rect 18254 9159 18270 9193
rect 18638 9159 18654 9193
rect 18254 9112 18654 9159
rect 18842 9265 19242 9312
rect 18842 9231 18858 9265
rect 19226 9231 19242 9265
rect 18842 9193 19242 9231
rect 18842 9159 18858 9193
rect 19226 9159 19242 9193
rect 18842 9112 19242 9159
rect 19430 9265 19830 9312
rect 19430 9231 19446 9265
rect 19814 9231 19830 9265
rect 19430 9193 19830 9231
rect 19430 9159 19446 9193
rect 19814 9159 19830 9193
rect 19430 9112 19830 9159
rect 20018 9265 20418 9312
rect 20018 9231 20034 9265
rect 20402 9231 20418 9265
rect 20018 9193 20418 9231
rect 20018 9159 20034 9193
rect 20402 9159 20418 9193
rect 20018 9112 20418 9159
rect 20606 9265 21006 9312
rect 20606 9231 20622 9265
rect 20990 9231 21006 9265
rect 20606 9193 21006 9231
rect 20606 9159 20622 9193
rect 20990 9159 21006 9193
rect 20606 9112 21006 9159
rect 21194 9265 21594 9312
rect 21194 9231 21210 9265
rect 21578 9231 21594 9265
rect 21194 9193 21594 9231
rect 21194 9159 21210 9193
rect 21578 9159 21594 9193
rect 21194 9112 21594 9159
rect 21782 9265 22182 9312
rect 21782 9231 21798 9265
rect 22166 9231 22182 9265
rect 21782 9193 22182 9231
rect 21782 9159 21798 9193
rect 22166 9159 22182 9193
rect 21782 9112 22182 9159
rect 22370 9265 22770 9312
rect 22370 9231 22386 9265
rect 22754 9231 22770 9265
rect 22370 9193 22770 9231
rect 22370 9159 22386 9193
rect 22754 9159 22770 9193
rect 22370 9112 22770 9159
rect 22958 9265 23358 9312
rect 22958 9231 22974 9265
rect 23342 9231 23358 9265
rect 22958 9193 23358 9231
rect 22958 9159 22974 9193
rect 23342 9159 23358 9193
rect 22958 9112 23358 9159
rect 23546 9265 23946 9312
rect 23546 9231 23562 9265
rect 23930 9231 23946 9265
rect 23546 9193 23946 9231
rect 23546 9159 23562 9193
rect 23930 9159 23946 9193
rect 23546 9112 23946 9159
rect 24134 9265 24534 9312
rect 24134 9231 24150 9265
rect 24518 9231 24534 9265
rect 24134 9193 24534 9231
rect 24134 9159 24150 9193
rect 24518 9159 24534 9193
rect 24134 9112 24534 9159
rect 24722 9265 25122 9312
rect 24722 9231 24738 9265
rect 25106 9231 25122 9265
rect 24722 9193 25122 9231
rect 24722 9159 24738 9193
rect 25106 9159 25122 9193
rect 24722 9112 25122 9159
rect 25310 9265 25710 9312
rect 25310 9231 25326 9265
rect 25694 9231 25710 9265
rect 25310 9193 25710 9231
rect 25310 9159 25326 9193
rect 25694 9159 25710 9193
rect 25310 9112 25710 9159
rect 25898 9265 26298 9312
rect 25898 9231 25914 9265
rect 26282 9231 26298 9265
rect 25898 9193 26298 9231
rect 25898 9159 25914 9193
rect 26282 9159 26298 9193
rect 25898 9112 26298 9159
rect 26486 9265 26886 9312
rect 26486 9231 26502 9265
rect 26870 9231 26886 9265
rect 26486 9193 26886 9231
rect 26486 9159 26502 9193
rect 26870 9159 26886 9193
rect 26486 9112 26886 9159
rect 27074 9265 27474 9312
rect 27074 9231 27090 9265
rect 27458 9231 27474 9265
rect 27074 9193 27474 9231
rect 27074 9159 27090 9193
rect 27458 9159 27474 9193
rect 27074 9112 27474 9159
rect 27662 9265 28062 9312
rect 27662 9231 27678 9265
rect 28046 9231 28062 9265
rect 27662 9193 28062 9231
rect 27662 9159 27678 9193
rect 28046 9159 28062 9193
rect 27662 9112 28062 9159
rect 28250 9265 28650 9312
rect 28250 9231 28266 9265
rect 28634 9231 28650 9265
rect 28250 9193 28650 9231
rect 28250 9159 28266 9193
rect 28634 9159 28650 9193
rect 28250 9112 28650 9159
rect 28838 9265 29238 9312
rect 28838 9231 28854 9265
rect 29222 9231 29238 9265
rect 28838 9193 29238 9231
rect 28838 9159 28854 9193
rect 29222 9159 29238 9193
rect 28838 9112 29238 9159
rect 29426 9265 29826 9312
rect 29426 9231 29442 9265
rect 29810 9231 29826 9265
rect 29426 9193 29826 9231
rect 29426 9159 29442 9193
rect 29810 9159 29826 9193
rect 29426 9112 29826 9159
rect 30014 9265 30414 9312
rect 30014 9231 30030 9265
rect 30398 9231 30414 9265
rect 30014 9193 30414 9231
rect 30014 9159 30030 9193
rect 30398 9159 30414 9193
rect 30014 9112 30414 9159
rect 30602 9265 31002 9312
rect 30602 9231 30618 9265
rect 30986 9231 31002 9265
rect 30602 9193 31002 9231
rect 30602 9159 30618 9193
rect 30986 9159 31002 9193
rect 30602 9112 31002 9159
rect 31190 9265 31590 9312
rect 31190 9231 31206 9265
rect 31574 9231 31590 9265
rect 31190 9193 31590 9231
rect 31190 9159 31206 9193
rect 31574 9159 31590 9193
rect 31190 9112 31590 9159
rect 31778 9265 32178 9312
rect 31778 9231 31794 9265
rect 32162 9231 32178 9265
rect 31778 9193 32178 9231
rect 31778 9159 31794 9193
rect 32162 9159 32178 9193
rect 31778 9112 32178 9159
rect 32366 9265 32766 9312
rect 32366 9231 32382 9265
rect 32750 9231 32766 9265
rect 32366 9193 32766 9231
rect 32366 9159 32382 9193
rect 32750 9159 32766 9193
rect 32366 9112 32766 9159
rect 32954 9265 33354 9312
rect 32954 9231 32970 9265
rect 33338 9231 33354 9265
rect 32954 9193 33354 9231
rect 32954 9159 32970 9193
rect 33338 9159 33354 9193
rect 32954 9112 33354 9159
rect 33542 9265 33942 9312
rect 33542 9231 33558 9265
rect 33926 9231 33942 9265
rect 33542 9193 33942 9231
rect 33542 9159 33558 9193
rect 33926 9159 33942 9193
rect 33542 9112 33942 9159
rect 34130 9265 34530 9312
rect 34130 9231 34146 9265
rect 34514 9231 34530 9265
rect 34130 9193 34530 9231
rect 34130 9159 34146 9193
rect 34514 9159 34530 9193
rect 34130 9112 34530 9159
rect 34718 9265 35118 9312
rect 34718 9231 34734 9265
rect 35102 9231 35118 9265
rect 34718 9193 35118 9231
rect 34718 9159 34734 9193
rect 35102 9159 35118 9193
rect 34718 9112 35118 9159
rect 35306 9265 35706 9312
rect 35306 9231 35322 9265
rect 35690 9231 35706 9265
rect 35306 9193 35706 9231
rect 35306 9159 35322 9193
rect 35690 9159 35706 9193
rect 35306 9112 35706 9159
rect 35894 9265 36294 9312
rect 35894 9231 35910 9265
rect 36278 9231 36294 9265
rect 35894 9193 36294 9231
rect 35894 9159 35910 9193
rect 36278 9159 36294 9193
rect 35894 9112 36294 9159
rect 36482 9265 36882 9312
rect 36482 9231 36498 9265
rect 36866 9231 36882 9265
rect 36482 9193 36882 9231
rect 36482 9159 36498 9193
rect 36866 9159 36882 9193
rect 36482 9112 36882 9159
rect 37070 9265 37470 9312
rect 37070 9231 37086 9265
rect 37454 9231 37470 9265
rect 37070 9193 37470 9231
rect 37070 9159 37086 9193
rect 37454 9159 37470 9193
rect 37070 9112 37470 9159
rect 37658 9265 38058 9312
rect 37658 9231 37674 9265
rect 38042 9231 38058 9265
rect 37658 9193 38058 9231
rect 37658 9159 37674 9193
rect 38042 9159 38058 9193
rect 37658 9112 38058 9159
rect 38246 9265 38646 9312
rect 38246 9231 38262 9265
rect 38630 9231 38646 9265
rect 38246 9193 38646 9231
rect 38246 9159 38262 9193
rect 38630 9159 38646 9193
rect 38246 9112 38646 9159
rect 10610 8265 11010 8312
rect 10610 8231 10626 8265
rect 10994 8231 11010 8265
rect 10610 8215 11010 8231
rect 11198 8265 11598 8312
rect 11198 8231 11214 8265
rect 11582 8231 11598 8265
rect 11198 8215 11598 8231
rect 11786 8265 12186 8312
rect 11786 8231 11802 8265
rect 12170 8231 12186 8265
rect 11786 8215 12186 8231
rect 12374 8265 12774 8312
rect 12374 8231 12390 8265
rect 12758 8231 12774 8265
rect 12374 8215 12774 8231
rect 12962 8265 13362 8312
rect 12962 8231 12978 8265
rect 13346 8231 13362 8265
rect 12962 8215 13362 8231
rect 13550 8265 13950 8312
rect 13550 8231 13566 8265
rect 13934 8231 13950 8265
rect 13550 8215 13950 8231
rect 14138 8265 14538 8312
rect 14138 8231 14154 8265
rect 14522 8231 14538 8265
rect 14138 8215 14538 8231
rect 14726 8265 15126 8312
rect 14726 8231 14742 8265
rect 15110 8231 15126 8265
rect 14726 8215 15126 8231
rect 15314 8265 15714 8312
rect 15314 8231 15330 8265
rect 15698 8231 15714 8265
rect 15314 8215 15714 8231
rect 15902 8265 16302 8312
rect 15902 8231 15918 8265
rect 16286 8231 16302 8265
rect 15902 8215 16302 8231
rect 16490 8265 16890 8312
rect 16490 8231 16506 8265
rect 16874 8231 16890 8265
rect 16490 8215 16890 8231
rect 17078 8265 17478 8312
rect 17078 8231 17094 8265
rect 17462 8231 17478 8265
rect 17078 8215 17478 8231
rect 17666 8265 18066 8312
rect 17666 8231 17682 8265
rect 18050 8231 18066 8265
rect 17666 8215 18066 8231
rect 18254 8265 18654 8312
rect 18254 8231 18270 8265
rect 18638 8231 18654 8265
rect 18254 8215 18654 8231
rect 18842 8265 19242 8312
rect 18842 8231 18858 8265
rect 19226 8231 19242 8265
rect 18842 8215 19242 8231
rect 19430 8265 19830 8312
rect 19430 8231 19446 8265
rect 19814 8231 19830 8265
rect 19430 8215 19830 8231
rect 20018 8265 20418 8312
rect 20018 8231 20034 8265
rect 20402 8231 20418 8265
rect 20018 8215 20418 8231
rect 20606 8265 21006 8312
rect 20606 8231 20622 8265
rect 20990 8231 21006 8265
rect 20606 8215 21006 8231
rect 21194 8265 21594 8312
rect 21194 8231 21210 8265
rect 21578 8231 21594 8265
rect 21194 8215 21594 8231
rect 21782 8265 22182 8312
rect 21782 8231 21798 8265
rect 22166 8231 22182 8265
rect 21782 8215 22182 8231
rect 22370 8265 22770 8312
rect 22370 8231 22386 8265
rect 22754 8231 22770 8265
rect 22370 8215 22770 8231
rect 22958 8265 23358 8312
rect 22958 8231 22974 8265
rect 23342 8231 23358 8265
rect 22958 8215 23358 8231
rect 23546 8265 23946 8312
rect 23546 8231 23562 8265
rect 23930 8231 23946 8265
rect 23546 8215 23946 8231
rect 24134 8265 24534 8312
rect 24134 8231 24150 8265
rect 24518 8231 24534 8265
rect 24134 8215 24534 8231
rect 24722 8265 25122 8312
rect 24722 8231 24738 8265
rect 25106 8231 25122 8265
rect 24722 8215 25122 8231
rect 25310 8265 25710 8312
rect 25310 8231 25326 8265
rect 25694 8231 25710 8265
rect 25310 8215 25710 8231
rect 25898 8265 26298 8312
rect 25898 8231 25914 8265
rect 26282 8231 26298 8265
rect 25898 8215 26298 8231
rect 26486 8265 26886 8312
rect 26486 8231 26502 8265
rect 26870 8231 26886 8265
rect 26486 8215 26886 8231
rect 27074 8265 27474 8312
rect 27074 8231 27090 8265
rect 27458 8231 27474 8265
rect 27074 8215 27474 8231
rect 27662 8265 28062 8312
rect 27662 8231 27678 8265
rect 28046 8231 28062 8265
rect 27662 8215 28062 8231
rect 28250 8265 28650 8312
rect 28250 8231 28266 8265
rect 28634 8231 28650 8265
rect 28250 8215 28650 8231
rect 28838 8265 29238 8312
rect 28838 8231 28854 8265
rect 29222 8231 29238 8265
rect 28838 8215 29238 8231
rect 29426 8265 29826 8312
rect 29426 8231 29442 8265
rect 29810 8231 29826 8265
rect 29426 8215 29826 8231
rect 30014 8265 30414 8312
rect 30014 8231 30030 8265
rect 30398 8231 30414 8265
rect 30014 8215 30414 8231
rect 30602 8265 31002 8312
rect 30602 8231 30618 8265
rect 30986 8231 31002 8265
rect 30602 8215 31002 8231
rect 31190 8265 31590 8312
rect 31190 8231 31206 8265
rect 31574 8231 31590 8265
rect 31190 8215 31590 8231
rect 31778 8265 32178 8312
rect 31778 8231 31794 8265
rect 32162 8231 32178 8265
rect 31778 8215 32178 8231
rect 32366 8265 32766 8312
rect 32366 8231 32382 8265
rect 32750 8231 32766 8265
rect 32366 8215 32766 8231
rect 32954 8265 33354 8312
rect 32954 8231 32970 8265
rect 33338 8231 33354 8265
rect 32954 8215 33354 8231
rect 33542 8265 33942 8312
rect 33542 8231 33558 8265
rect 33926 8231 33942 8265
rect 33542 8215 33942 8231
rect 34130 8265 34530 8312
rect 34130 8231 34146 8265
rect 34514 8231 34530 8265
rect 34130 8215 34530 8231
rect 34718 8265 35118 8312
rect 34718 8231 34734 8265
rect 35102 8231 35118 8265
rect 34718 8215 35118 8231
rect 35306 8265 35706 8312
rect 35306 8231 35322 8265
rect 35690 8231 35706 8265
rect 35306 8215 35706 8231
rect 35894 8265 36294 8312
rect 35894 8231 35910 8265
rect 36278 8231 36294 8265
rect 35894 8215 36294 8231
rect 36482 8265 36882 8312
rect 36482 8231 36498 8265
rect 36866 8231 36882 8265
rect 36482 8215 36882 8231
rect 37070 8265 37470 8312
rect 37070 8231 37086 8265
rect 37454 8231 37470 8265
rect 37070 8215 37470 8231
rect 37658 8265 38058 8312
rect 37658 8231 37674 8265
rect 38042 8231 38058 8265
rect 37658 8215 38058 8231
rect 38246 8265 38646 8312
rect 38246 8231 38262 8265
rect 38630 8231 38646 8265
rect 38246 8215 38646 8231
rect 23662 6836 23732 6842
rect 23662 6704 23678 6836
rect 23716 6704 23732 6836
rect 23662 6666 23732 6704
rect 23928 6836 23998 6842
rect 23928 6704 23944 6836
rect 23982 6704 23998 6836
rect 23928 6666 23998 6704
rect 24194 6836 24264 6842
rect 24194 6704 24210 6836
rect 24248 6704 24264 6836
rect 24194 6666 24264 6704
rect 24460 6836 24530 6842
rect 24460 6704 24476 6836
rect 24514 6704 24530 6836
rect 24460 6666 24530 6704
rect 24726 6836 24796 6842
rect 24726 6704 24742 6836
rect 24780 6704 24796 6836
rect 24726 6666 24796 6704
rect 24992 6836 25062 6842
rect 24992 6704 25008 6836
rect 25046 6704 25062 6836
rect 24992 6666 25062 6704
rect 25258 6836 25328 6842
rect 25258 6704 25274 6836
rect 25312 6704 25328 6836
rect 25258 6666 25328 6704
rect 25524 6836 25594 6842
rect 25524 6704 25540 6836
rect 25578 6704 25594 6836
rect 25524 6666 25594 6704
rect 23662 5826 23732 5866
rect 23662 5694 23678 5826
rect 23716 5694 23732 5826
rect 23662 5656 23732 5694
rect 23928 5826 23998 5866
rect 23928 5694 23944 5826
rect 23982 5694 23998 5826
rect 23928 5656 23998 5694
rect 24194 5826 24264 5866
rect 24194 5694 24210 5826
rect 24248 5694 24264 5826
rect 24194 5656 24264 5694
rect 24460 5826 24530 5866
rect 24460 5694 24476 5826
rect 24514 5694 24530 5826
rect 24460 5656 24530 5694
rect 24726 5826 24796 5866
rect 24726 5694 24742 5826
rect 24780 5694 24796 5826
rect 24726 5656 24796 5694
rect 24992 5826 25062 5866
rect 24992 5694 25008 5826
rect 25046 5694 25062 5826
rect 24992 5656 25062 5694
rect 25258 5826 25328 5866
rect 25258 5694 25274 5826
rect 25312 5694 25328 5826
rect 25258 5656 25328 5694
rect 25524 5826 25594 5866
rect 25524 5694 25540 5826
rect 25578 5694 25594 5826
rect 25524 5656 25594 5694
rect 23662 4816 23732 4856
rect 23662 4684 23678 4816
rect 23716 4684 23732 4816
rect 23662 4646 23732 4684
rect 23928 4816 23998 4856
rect 23928 4684 23944 4816
rect 23982 4684 23998 4816
rect 23928 4646 23998 4684
rect 24194 4816 24264 4856
rect 24194 4684 24210 4816
rect 24248 4684 24264 4816
rect 24194 4646 24264 4684
rect 24460 4816 24530 4856
rect 24460 4684 24476 4816
rect 24514 4684 24530 4816
rect 24460 4646 24530 4684
rect 24726 4816 24796 4856
rect 24726 4684 24742 4816
rect 24780 4684 24796 4816
rect 24726 4646 24796 4684
rect 24992 4816 25062 4856
rect 24992 4684 25008 4816
rect 25046 4684 25062 4816
rect 24992 4646 25062 4684
rect 25258 4816 25328 4856
rect 25258 4684 25274 4816
rect 25312 4684 25328 4816
rect 25258 4646 25328 4684
rect 25524 4816 25594 4856
rect 25524 4684 25540 4816
rect 25578 4684 25594 4816
rect 25524 4646 25594 4684
rect 23662 3806 23732 3846
rect 23662 3674 23678 3806
rect 23716 3674 23732 3806
rect 23662 3664 23732 3674
rect 23928 3806 23998 3846
rect 23928 3674 23944 3806
rect 23982 3674 23998 3806
rect 23928 3664 23998 3674
rect 24194 3806 24264 3846
rect 24194 3674 24210 3806
rect 24248 3674 24264 3806
rect 24194 3664 24264 3674
rect 24460 3806 24530 3846
rect 24460 3674 24476 3806
rect 24514 3674 24530 3806
rect 24460 3664 24530 3674
rect 24726 3806 24796 3846
rect 24726 3674 24742 3806
rect 24780 3674 24796 3806
rect 24726 3664 24796 3674
rect 24992 3806 25062 3846
rect 24992 3674 25008 3806
rect 25046 3674 25062 3806
rect 24992 3664 25062 3674
rect 25258 3806 25328 3846
rect 25258 3674 25274 3806
rect 25312 3674 25328 3806
rect 25258 3664 25328 3674
rect 25524 3806 25594 3846
rect 25524 3674 25540 3806
rect 25578 3674 25594 3806
rect 25524 3664 25594 3674
rect 24234 2638 24304 2644
rect 24234 2512 24250 2638
rect 24288 2512 24304 2638
rect 24234 2474 24304 2512
rect 24474 2638 24544 2644
rect 24474 2512 24490 2638
rect 24528 2512 24544 2638
rect 24474 2474 24544 2512
rect 24714 2638 24784 2644
rect 24714 2512 24730 2638
rect 24768 2512 24784 2638
rect 24714 2474 24784 2512
rect 24954 2638 25024 2644
rect 24954 2512 24970 2638
rect 25008 2512 25024 2638
rect 24954 2474 25024 2512
rect 24234 1836 24304 1874
rect 24234 1704 24250 1836
rect 24288 1704 24304 1836
rect 24234 1666 24304 1704
rect 24474 1836 24544 1874
rect 24474 1704 24490 1836
rect 24528 1704 24544 1836
rect 24474 1666 24544 1704
rect 24714 1836 24784 1874
rect 24714 1704 24730 1836
rect 24768 1704 24784 1836
rect 24714 1666 24784 1704
rect 24954 1836 25024 1874
rect 24954 1704 24970 1836
rect 25008 1704 25024 1836
rect 24954 1666 25024 1704
rect 24234 1028 24304 1066
rect 24234 896 24250 1028
rect 24288 896 24304 1028
rect 24474 1028 24544 1066
rect 24474 896 24490 1028
rect 24528 896 24544 1028
rect 24714 1028 24784 1066
rect 24714 896 24730 1028
rect 24768 896 24784 1028
rect 24954 1028 25024 1066
rect 24954 896 24970 1028
rect 25008 896 25024 1028
<< polycont >>
rect 19930 15168 19968 15300
rect 20170 15168 20208 15300
rect 20410 15168 20448 15300
rect 20650 15168 20688 15300
rect 20890 15168 20928 15300
rect 21130 15168 21168 15300
rect 21370 15168 21408 15300
rect 21610 15168 21648 15300
rect 21850 15168 21888 15300
rect 22090 15168 22128 15300
rect 22330 15168 22368 15300
rect 22570 15168 22608 15300
rect 22810 15168 22848 15300
rect 23050 15168 23088 15300
rect 23290 15168 23328 15300
rect 23530 15168 23568 15300
rect 23770 15168 23808 15300
rect 24010 15168 24048 15300
rect 24250 15168 24288 15300
rect 24490 15168 24528 15300
rect 24730 15168 24768 15300
rect 24970 15168 25008 15300
rect 25210 15168 25248 15300
rect 25450 15168 25488 15300
rect 25690 15168 25728 15300
rect 25930 15168 25968 15300
rect 26170 15168 26208 15300
rect 26410 15168 26448 15300
rect 26650 15168 26688 15300
rect 26890 15168 26928 15300
rect 27130 15168 27168 15300
rect 27370 15168 27408 15300
rect 27610 15168 27648 15300
rect 27850 15168 27888 15300
rect 28090 15168 28128 15300
rect 28330 15168 28368 15300
rect 28570 15168 28608 15300
rect 28810 15168 28848 15300
rect 29050 15168 29088 15300
rect 29290 15168 29328 15300
rect 19930 14360 19968 14492
rect 20170 14360 20208 14492
rect 20410 14360 20448 14492
rect 20650 14360 20688 14492
rect 20890 14360 20928 14492
rect 21130 14360 21168 14492
rect 21370 14360 21408 14492
rect 21610 14360 21648 14492
rect 21850 14360 21888 14492
rect 22090 14360 22128 14492
rect 22330 14360 22368 14492
rect 22570 14360 22608 14492
rect 22810 14360 22848 14492
rect 23050 14360 23088 14492
rect 23290 14360 23328 14492
rect 23530 14360 23568 14492
rect 23770 14360 23808 14492
rect 24010 14360 24048 14492
rect 24250 14360 24288 14492
rect 24490 14360 24528 14492
rect 24730 14360 24768 14492
rect 24970 14360 25008 14492
rect 25210 14360 25248 14492
rect 25450 14360 25488 14492
rect 25690 14360 25728 14492
rect 25930 14360 25968 14492
rect 26170 14360 26208 14492
rect 26410 14360 26448 14492
rect 26650 14360 26688 14492
rect 26890 14360 26928 14492
rect 27130 14360 27168 14492
rect 27370 14360 27408 14492
rect 27610 14360 27648 14492
rect 27850 14360 27888 14492
rect 28090 14360 28128 14492
rect 28330 14360 28368 14492
rect 28570 14360 28608 14492
rect 28810 14360 28848 14492
rect 29050 14360 29088 14492
rect 29290 14360 29328 14492
rect 19930 13552 19968 13684
rect 20170 13552 20208 13684
rect 20410 13552 20448 13684
rect 20650 13552 20688 13684
rect 20890 13552 20928 13684
rect 21130 13552 21168 13684
rect 21370 13552 21408 13684
rect 21610 13552 21648 13684
rect 21850 13552 21888 13684
rect 22090 13552 22128 13684
rect 22330 13552 22368 13684
rect 22570 13552 22608 13684
rect 22810 13552 22848 13684
rect 23050 13552 23088 13684
rect 23290 13552 23328 13684
rect 23530 13552 23568 13684
rect 23770 13552 23808 13684
rect 24010 13552 24048 13684
rect 24250 13552 24288 13684
rect 24490 13552 24528 13684
rect 24730 13552 24768 13684
rect 24970 13552 25008 13684
rect 25210 13552 25248 13684
rect 25450 13552 25488 13684
rect 25690 13552 25728 13684
rect 25930 13552 25968 13684
rect 26170 13552 26208 13684
rect 26410 13552 26448 13684
rect 26650 13552 26688 13684
rect 26890 13552 26928 13684
rect 27130 13552 27168 13684
rect 27370 13552 27408 13684
rect 27610 13552 27648 13684
rect 27850 13552 27888 13684
rect 28090 13552 28128 13684
rect 28330 13552 28368 13684
rect 28570 13552 28608 13684
rect 28810 13552 28848 13684
rect 29050 13552 29088 13684
rect 29290 13552 29328 13684
rect 10626 11159 10994 11193
rect 11214 11159 11582 11193
rect 11802 11159 12170 11193
rect 12390 11159 12758 11193
rect 12978 11159 13346 11193
rect 13566 11159 13934 11193
rect 14154 11159 14522 11193
rect 14742 11159 15110 11193
rect 15330 11159 15698 11193
rect 15918 11159 16286 11193
rect 16506 11159 16874 11193
rect 17094 11159 17462 11193
rect 17682 11159 18050 11193
rect 18270 11159 18638 11193
rect 18858 11159 19226 11193
rect 19446 11159 19814 11193
rect 20034 11159 20402 11193
rect 20622 11159 20990 11193
rect 21210 11159 21578 11193
rect 21798 11159 22166 11193
rect 22386 11159 22754 11193
rect 22974 11159 23342 11193
rect 23562 11159 23930 11193
rect 24150 11159 24518 11193
rect 24738 11159 25106 11193
rect 25326 11159 25694 11193
rect 25914 11159 26282 11193
rect 26502 11159 26870 11193
rect 27090 11159 27458 11193
rect 27678 11159 28046 11193
rect 28266 11159 28634 11193
rect 28854 11159 29222 11193
rect 29442 11159 29810 11193
rect 30030 11159 30398 11193
rect 30618 11159 30986 11193
rect 31206 11159 31574 11193
rect 31794 11159 32162 11193
rect 32382 11159 32750 11193
rect 32970 11159 33338 11193
rect 33558 11159 33926 11193
rect 34146 11159 34514 11193
rect 34734 11159 35102 11193
rect 35322 11159 35690 11193
rect 35910 11159 36278 11193
rect 36498 11159 36866 11193
rect 37086 11159 37454 11193
rect 37674 11159 38042 11193
rect 38262 11159 38630 11193
rect 10626 10231 10994 10265
rect 10626 10159 10994 10193
rect 11214 10231 11582 10265
rect 11214 10159 11582 10193
rect 11802 10231 12170 10265
rect 11802 10159 12170 10193
rect 12390 10231 12758 10265
rect 12390 10159 12758 10193
rect 12978 10231 13346 10265
rect 12978 10159 13346 10193
rect 13566 10231 13934 10265
rect 13566 10159 13934 10193
rect 14154 10231 14522 10265
rect 14154 10159 14522 10193
rect 14742 10231 15110 10265
rect 14742 10159 15110 10193
rect 15330 10231 15698 10265
rect 15330 10159 15698 10193
rect 15918 10231 16286 10265
rect 15918 10159 16286 10193
rect 16506 10231 16874 10265
rect 16506 10159 16874 10193
rect 17094 10231 17462 10265
rect 17094 10159 17462 10193
rect 17682 10231 18050 10265
rect 17682 10159 18050 10193
rect 18270 10231 18638 10265
rect 18270 10159 18638 10193
rect 18858 10231 19226 10265
rect 18858 10159 19226 10193
rect 19446 10231 19814 10265
rect 19446 10159 19814 10193
rect 20034 10231 20402 10265
rect 20034 10159 20402 10193
rect 20622 10231 20990 10265
rect 20622 10159 20990 10193
rect 21210 10231 21578 10265
rect 21210 10159 21578 10193
rect 21798 10231 22166 10265
rect 21798 10159 22166 10193
rect 22386 10231 22754 10265
rect 22386 10159 22754 10193
rect 22974 10231 23342 10265
rect 22974 10159 23342 10193
rect 23562 10231 23930 10265
rect 23562 10159 23930 10193
rect 24150 10231 24518 10265
rect 24150 10159 24518 10193
rect 24738 10231 25106 10265
rect 24738 10159 25106 10193
rect 25326 10231 25694 10265
rect 25326 10159 25694 10193
rect 25914 10231 26282 10265
rect 25914 10159 26282 10193
rect 26502 10231 26870 10265
rect 26502 10159 26870 10193
rect 27090 10231 27458 10265
rect 27090 10159 27458 10193
rect 27678 10231 28046 10265
rect 27678 10159 28046 10193
rect 28266 10231 28634 10265
rect 28266 10159 28634 10193
rect 28854 10231 29222 10265
rect 28854 10159 29222 10193
rect 29442 10231 29810 10265
rect 29442 10159 29810 10193
rect 30030 10231 30398 10265
rect 30030 10159 30398 10193
rect 30618 10231 30986 10265
rect 30618 10159 30986 10193
rect 31206 10231 31574 10265
rect 31206 10159 31574 10193
rect 31794 10231 32162 10265
rect 31794 10159 32162 10193
rect 32382 10231 32750 10265
rect 32382 10159 32750 10193
rect 32970 10231 33338 10265
rect 32970 10159 33338 10193
rect 33558 10231 33926 10265
rect 33558 10159 33926 10193
rect 34146 10231 34514 10265
rect 34146 10159 34514 10193
rect 34734 10231 35102 10265
rect 34734 10159 35102 10193
rect 35322 10231 35690 10265
rect 35322 10159 35690 10193
rect 35910 10231 36278 10265
rect 35910 10159 36278 10193
rect 36498 10231 36866 10265
rect 36498 10159 36866 10193
rect 37086 10231 37454 10265
rect 37086 10159 37454 10193
rect 37674 10231 38042 10265
rect 37674 10159 38042 10193
rect 38262 10231 38630 10265
rect 38262 10159 38630 10193
rect 10626 9231 10994 9265
rect 10626 9159 10994 9193
rect 11214 9231 11582 9265
rect 11214 9159 11582 9193
rect 11802 9231 12170 9265
rect 11802 9159 12170 9193
rect 12390 9231 12758 9265
rect 12390 9159 12758 9193
rect 12978 9231 13346 9265
rect 12978 9159 13346 9193
rect 13566 9231 13934 9265
rect 13566 9159 13934 9193
rect 14154 9231 14522 9265
rect 14154 9159 14522 9193
rect 14742 9231 15110 9265
rect 14742 9159 15110 9193
rect 15330 9231 15698 9265
rect 15330 9159 15698 9193
rect 15918 9231 16286 9265
rect 15918 9159 16286 9193
rect 16506 9231 16874 9265
rect 16506 9159 16874 9193
rect 17094 9231 17462 9265
rect 17094 9159 17462 9193
rect 17682 9231 18050 9265
rect 17682 9159 18050 9193
rect 18270 9231 18638 9265
rect 18270 9159 18638 9193
rect 18858 9231 19226 9265
rect 18858 9159 19226 9193
rect 19446 9231 19814 9265
rect 19446 9159 19814 9193
rect 20034 9231 20402 9265
rect 20034 9159 20402 9193
rect 20622 9231 20990 9265
rect 20622 9159 20990 9193
rect 21210 9231 21578 9265
rect 21210 9159 21578 9193
rect 21798 9231 22166 9265
rect 21798 9159 22166 9193
rect 22386 9231 22754 9265
rect 22386 9159 22754 9193
rect 22974 9231 23342 9265
rect 22974 9159 23342 9193
rect 23562 9231 23930 9265
rect 23562 9159 23930 9193
rect 24150 9231 24518 9265
rect 24150 9159 24518 9193
rect 24738 9231 25106 9265
rect 24738 9159 25106 9193
rect 25326 9231 25694 9265
rect 25326 9159 25694 9193
rect 25914 9231 26282 9265
rect 25914 9159 26282 9193
rect 26502 9231 26870 9265
rect 26502 9159 26870 9193
rect 27090 9231 27458 9265
rect 27090 9159 27458 9193
rect 27678 9231 28046 9265
rect 27678 9159 28046 9193
rect 28266 9231 28634 9265
rect 28266 9159 28634 9193
rect 28854 9231 29222 9265
rect 28854 9159 29222 9193
rect 29442 9231 29810 9265
rect 29442 9159 29810 9193
rect 30030 9231 30398 9265
rect 30030 9159 30398 9193
rect 30618 9231 30986 9265
rect 30618 9159 30986 9193
rect 31206 9231 31574 9265
rect 31206 9159 31574 9193
rect 31794 9231 32162 9265
rect 31794 9159 32162 9193
rect 32382 9231 32750 9265
rect 32382 9159 32750 9193
rect 32970 9231 33338 9265
rect 32970 9159 33338 9193
rect 33558 9231 33926 9265
rect 33558 9159 33926 9193
rect 34146 9231 34514 9265
rect 34146 9159 34514 9193
rect 34734 9231 35102 9265
rect 34734 9159 35102 9193
rect 35322 9231 35690 9265
rect 35322 9159 35690 9193
rect 35910 9231 36278 9265
rect 35910 9159 36278 9193
rect 36498 9231 36866 9265
rect 36498 9159 36866 9193
rect 37086 9231 37454 9265
rect 37086 9159 37454 9193
rect 37674 9231 38042 9265
rect 37674 9159 38042 9193
rect 38262 9231 38630 9265
rect 38262 9159 38630 9193
rect 10626 8231 10994 8265
rect 11214 8231 11582 8265
rect 11802 8231 12170 8265
rect 12390 8231 12758 8265
rect 12978 8231 13346 8265
rect 13566 8231 13934 8265
rect 14154 8231 14522 8265
rect 14742 8231 15110 8265
rect 15330 8231 15698 8265
rect 15918 8231 16286 8265
rect 16506 8231 16874 8265
rect 17094 8231 17462 8265
rect 17682 8231 18050 8265
rect 18270 8231 18638 8265
rect 18858 8231 19226 8265
rect 19446 8231 19814 8265
rect 20034 8231 20402 8265
rect 20622 8231 20990 8265
rect 21210 8231 21578 8265
rect 21798 8231 22166 8265
rect 22386 8231 22754 8265
rect 22974 8231 23342 8265
rect 23562 8231 23930 8265
rect 24150 8231 24518 8265
rect 24738 8231 25106 8265
rect 25326 8231 25694 8265
rect 25914 8231 26282 8265
rect 26502 8231 26870 8265
rect 27090 8231 27458 8265
rect 27678 8231 28046 8265
rect 28266 8231 28634 8265
rect 28854 8231 29222 8265
rect 29442 8231 29810 8265
rect 30030 8231 30398 8265
rect 30618 8231 30986 8265
rect 31206 8231 31574 8265
rect 31794 8231 32162 8265
rect 32382 8231 32750 8265
rect 32970 8231 33338 8265
rect 33558 8231 33926 8265
rect 34146 8231 34514 8265
rect 34734 8231 35102 8265
rect 35322 8231 35690 8265
rect 35910 8231 36278 8265
rect 36498 8231 36866 8265
rect 37086 8231 37454 8265
rect 37674 8231 38042 8265
rect 38262 8231 38630 8265
rect 23678 6704 23716 6836
rect 23944 6704 23982 6836
rect 24210 6704 24248 6836
rect 24476 6704 24514 6836
rect 24742 6704 24780 6836
rect 25008 6704 25046 6836
rect 25274 6704 25312 6836
rect 25540 6704 25578 6836
rect 23678 5694 23716 5826
rect 23944 5694 23982 5826
rect 24210 5694 24248 5826
rect 24476 5694 24514 5826
rect 24742 5694 24780 5826
rect 25008 5694 25046 5826
rect 25274 5694 25312 5826
rect 25540 5694 25578 5826
rect 23678 4684 23716 4816
rect 23944 4684 23982 4816
rect 24210 4684 24248 4816
rect 24476 4684 24514 4816
rect 24742 4684 24780 4816
rect 25008 4684 25046 4816
rect 25274 4684 25312 4816
rect 25540 4684 25578 4816
rect 23678 3674 23716 3806
rect 23944 3674 23982 3806
rect 24210 3674 24248 3806
rect 24476 3674 24514 3806
rect 24742 3674 24780 3806
rect 25008 3674 25046 3806
rect 25274 3674 25312 3806
rect 25540 3674 25578 3806
rect 24250 2512 24288 2638
rect 24490 2512 24528 2638
rect 24730 2512 24768 2638
rect 24970 2512 25008 2638
rect 24250 1704 24288 1836
rect 24490 1704 24528 1836
rect 24730 1704 24768 1836
rect 24970 1704 25008 1836
rect 24250 896 24288 1028
rect 24490 896 24528 1028
rect 24730 896 24768 1028
rect 24970 896 25008 1028
<< xpolycontact >>
rect 30781 4727 30851 5159
rect 30781 3735 30851 4167
<< xpolyres >>
rect 30781 4167 30851 4727
<< locali >>
rect 19522 15610 19610 15644
rect 29648 15610 29736 15644
rect 19522 15576 19556 15610
rect 29702 15578 29736 15610
rect 19914 15168 19930 15300
rect 19968 15168 20170 15300
rect 20208 15168 20410 15300
rect 20448 15168 20650 15300
rect 20688 15168 20890 15300
rect 20928 15168 21130 15300
rect 21168 15168 21370 15300
rect 21408 15168 21610 15300
rect 21648 15168 21850 15300
rect 21888 15168 22090 15300
rect 22128 15168 22330 15300
rect 22368 15168 22570 15300
rect 22608 15168 22810 15300
rect 22848 15168 23050 15300
rect 23088 15168 23290 15300
rect 23328 15168 23530 15300
rect 23568 15168 23770 15300
rect 23808 15168 24010 15300
rect 24048 15168 24250 15300
rect 24288 15168 24490 15300
rect 24528 15168 24730 15300
rect 24768 15168 24970 15300
rect 25008 15168 25210 15300
rect 25248 15168 25450 15300
rect 25488 15168 25690 15300
rect 25728 15168 25930 15300
rect 25968 15168 26170 15300
rect 26208 15168 26410 15300
rect 26448 15168 26650 15300
rect 26688 15168 26890 15300
rect 26928 15168 27130 15300
rect 27168 15168 27370 15300
rect 27408 15168 27610 15300
rect 27648 15168 27850 15300
rect 27888 15168 28090 15300
rect 28128 15168 28330 15300
rect 28368 15168 28570 15300
rect 28608 15168 28810 15300
rect 28848 15168 29050 15300
rect 29088 15168 29290 15300
rect 29328 15168 29354 15300
rect 19868 15118 19902 15134
rect 19868 14526 19902 14542
rect 19996 15118 20030 15134
rect 19996 14526 20030 14542
rect 20108 15118 20142 15134
rect 20108 14526 20142 14542
rect 20236 15118 20270 15134
rect 20236 14526 20270 14542
rect 20348 15118 20382 15134
rect 20348 14526 20382 14542
rect 20476 15118 20510 15134
rect 20476 14526 20510 14542
rect 20588 15118 20622 15134
rect 20588 14526 20622 14542
rect 20716 15118 20750 15134
rect 20716 14526 20750 14542
rect 20828 15118 20862 15134
rect 20828 14526 20862 14542
rect 20956 15118 20990 15134
rect 20956 14526 20990 14542
rect 21068 15118 21102 15134
rect 21068 14526 21102 14542
rect 21196 15118 21230 15134
rect 21196 14526 21230 14542
rect 21308 15118 21342 15134
rect 21308 14526 21342 14542
rect 21436 15118 21470 15134
rect 21436 14526 21470 14542
rect 21548 15118 21582 15134
rect 21548 14526 21582 14542
rect 21676 15118 21710 15134
rect 21676 14526 21710 14542
rect 21788 15118 21822 15134
rect 21788 14526 21822 14542
rect 21916 15118 21950 15134
rect 21916 14526 21950 14542
rect 22028 15118 22062 15134
rect 22028 14526 22062 14542
rect 22156 15118 22190 15134
rect 22156 14526 22190 14542
rect 22268 15118 22302 15134
rect 22268 14526 22302 14542
rect 22396 15118 22430 15134
rect 22396 14526 22430 14542
rect 22508 15118 22542 15134
rect 22508 14526 22542 14542
rect 22636 15118 22670 15134
rect 22636 14526 22670 14542
rect 22748 15118 22782 15134
rect 22748 14526 22782 14542
rect 22876 15118 22910 15134
rect 22876 14526 22910 14542
rect 22988 15118 23022 15134
rect 22988 14526 23022 14542
rect 23116 15118 23150 15134
rect 23116 14526 23150 14542
rect 23228 15118 23262 15134
rect 23228 14526 23262 14542
rect 23356 15118 23390 15134
rect 23356 14526 23390 14542
rect 23468 15118 23502 15134
rect 23468 14526 23502 14542
rect 23596 15118 23630 15134
rect 23596 14526 23630 14542
rect 23708 15118 23742 15134
rect 23708 14526 23742 14542
rect 23836 15118 23870 15134
rect 23836 14526 23870 14542
rect 23948 15118 23982 15134
rect 23948 14526 23982 14542
rect 24076 15118 24110 15134
rect 24076 14526 24110 14542
rect 24188 15118 24222 15134
rect 24188 14526 24222 14542
rect 24316 15118 24350 15134
rect 24316 14526 24350 14542
rect 24428 15118 24462 15134
rect 24428 14526 24462 14542
rect 24556 15118 24590 15134
rect 24556 14526 24590 14542
rect 24668 15118 24702 15134
rect 24668 14526 24702 14542
rect 24796 15118 24830 15134
rect 24796 14526 24830 14542
rect 24908 15118 24942 15134
rect 24908 14526 24942 14542
rect 25036 15118 25070 15134
rect 25036 14526 25070 14542
rect 25148 15118 25182 15134
rect 25148 14526 25182 14542
rect 25276 15118 25310 15134
rect 25276 14526 25310 14542
rect 25388 15118 25422 15134
rect 25388 14526 25422 14542
rect 25516 15118 25550 15134
rect 25516 14526 25550 14542
rect 25628 15118 25662 15134
rect 25628 14526 25662 14542
rect 25756 15118 25790 15134
rect 25756 14526 25790 14542
rect 25868 15118 25902 15134
rect 25868 14526 25902 14542
rect 25996 15118 26030 15134
rect 25996 14526 26030 14542
rect 26108 15118 26142 15134
rect 26108 14526 26142 14542
rect 26236 15118 26270 15134
rect 26236 14526 26270 14542
rect 26348 15118 26382 15134
rect 26348 14526 26382 14542
rect 26476 15118 26510 15134
rect 26476 14526 26510 14542
rect 26588 15118 26622 15134
rect 26588 14526 26622 14542
rect 26716 15118 26750 15134
rect 26716 14526 26750 14542
rect 26828 15118 26862 15134
rect 26828 14526 26862 14542
rect 26956 15118 26990 15134
rect 26956 14526 26990 14542
rect 27068 15118 27102 15134
rect 27068 14526 27102 14542
rect 27196 15118 27230 15134
rect 27196 14526 27230 14542
rect 27308 15118 27342 15134
rect 27308 14526 27342 14542
rect 27436 15118 27470 15134
rect 27436 14526 27470 14542
rect 27548 15118 27582 15134
rect 27548 14526 27582 14542
rect 27676 15118 27710 15134
rect 27676 14526 27710 14542
rect 27788 15118 27822 15134
rect 27788 14526 27822 14542
rect 27916 15118 27950 15134
rect 27916 14526 27950 14542
rect 28028 15118 28062 15134
rect 28028 14526 28062 14542
rect 28156 15118 28190 15134
rect 28156 14526 28190 14542
rect 28268 15118 28302 15134
rect 28268 14526 28302 14542
rect 28396 15118 28430 15134
rect 28396 14526 28430 14542
rect 28508 15118 28542 15134
rect 28508 14526 28542 14542
rect 28636 15118 28670 15134
rect 28636 14526 28670 14542
rect 28748 15118 28782 15134
rect 28748 14526 28782 14542
rect 28876 15118 28910 15134
rect 28876 14526 28910 14542
rect 28988 15118 29022 15134
rect 28988 14526 29022 14542
rect 29116 15118 29150 15134
rect 29116 14526 29150 14542
rect 29228 15118 29262 15134
rect 29228 14526 29262 14542
rect 29356 15118 29390 15134
rect 29356 14526 29390 14542
rect 19914 14360 19930 14492
rect 19968 14360 20170 14492
rect 20208 14360 20410 14492
rect 20448 14360 20650 14492
rect 20688 14360 20890 14492
rect 20928 14360 21130 14492
rect 21168 14360 21370 14492
rect 21408 14360 21610 14492
rect 21648 14360 21850 14492
rect 21888 14360 22090 14492
rect 22128 14360 22330 14492
rect 22368 14360 22570 14492
rect 22608 14360 22810 14492
rect 22848 14360 23050 14492
rect 23088 14360 23290 14492
rect 23328 14360 23530 14492
rect 23568 14360 23770 14492
rect 23808 14360 24010 14492
rect 24048 14360 24250 14492
rect 24288 14360 24490 14492
rect 24528 14360 24730 14492
rect 24768 14360 24970 14492
rect 25008 14360 25210 14492
rect 25248 14360 25450 14492
rect 25488 14360 25690 14492
rect 25728 14360 25930 14492
rect 25968 14360 26170 14492
rect 26208 14360 26410 14492
rect 26448 14360 26650 14492
rect 26688 14360 26890 14492
rect 26928 14360 27130 14492
rect 27168 14360 27370 14492
rect 27408 14360 27610 14492
rect 27648 14360 27850 14492
rect 27888 14360 28090 14492
rect 28128 14360 28330 14492
rect 28368 14360 28570 14492
rect 28608 14360 28810 14492
rect 28848 14360 29050 14492
rect 29088 14360 29290 14492
rect 29328 14360 29354 14492
rect 19868 14310 19902 14326
rect 19868 13718 19902 13734
rect 19996 14310 20030 14326
rect 19996 13718 20030 13734
rect 20108 14310 20142 14326
rect 20108 13718 20142 13734
rect 20236 14310 20270 14326
rect 20236 13718 20270 13734
rect 20348 14310 20382 14326
rect 20348 13718 20382 13734
rect 20476 14310 20510 14326
rect 20476 13718 20510 13734
rect 20588 14310 20622 14326
rect 20588 13718 20622 13734
rect 20716 14310 20750 14326
rect 20716 13718 20750 13734
rect 20828 14310 20862 14326
rect 20828 13718 20862 13734
rect 20956 14310 20990 14326
rect 20956 13718 20990 13734
rect 21068 14310 21102 14326
rect 21068 13718 21102 13734
rect 21196 14310 21230 14326
rect 21196 13718 21230 13734
rect 21308 14310 21342 14326
rect 21308 13718 21342 13734
rect 21436 14310 21470 14326
rect 21436 13718 21470 13734
rect 21548 14310 21582 14326
rect 21548 13718 21582 13734
rect 21676 14310 21710 14326
rect 21676 13718 21710 13734
rect 21788 14310 21822 14326
rect 21788 13718 21822 13734
rect 21916 14310 21950 14326
rect 21916 13718 21950 13734
rect 22028 14310 22062 14326
rect 22028 13718 22062 13734
rect 22156 14310 22190 14326
rect 22156 13718 22190 13734
rect 22268 14310 22302 14326
rect 22268 13718 22302 13734
rect 22396 14310 22430 14326
rect 22396 13718 22430 13734
rect 22508 14310 22542 14326
rect 22508 13718 22542 13734
rect 22636 14310 22670 14326
rect 22636 13718 22670 13734
rect 22748 14310 22782 14326
rect 22748 13718 22782 13734
rect 22876 14310 22910 14326
rect 22876 13718 22910 13734
rect 22988 14310 23022 14326
rect 22988 13718 23022 13734
rect 23116 14310 23150 14326
rect 23116 13718 23150 13734
rect 23228 14310 23262 14326
rect 23228 13718 23262 13734
rect 23356 14310 23390 14326
rect 23356 13718 23390 13734
rect 23468 14310 23502 14326
rect 23468 13718 23502 13734
rect 23596 14310 23630 14326
rect 23596 13718 23630 13734
rect 23708 14310 23742 14326
rect 23708 13718 23742 13734
rect 23836 14310 23870 14326
rect 23836 13718 23870 13734
rect 23948 14310 23982 14326
rect 23948 13718 23982 13734
rect 24076 14310 24110 14326
rect 24076 13718 24110 13734
rect 24188 14310 24222 14326
rect 24188 13718 24222 13734
rect 24316 14310 24350 14326
rect 24316 13718 24350 13734
rect 24428 14310 24462 14326
rect 24428 13718 24462 13734
rect 24556 14310 24590 14326
rect 24556 13718 24590 13734
rect 24668 14310 24702 14326
rect 24668 13718 24702 13734
rect 24796 14310 24830 14326
rect 24796 13718 24830 13734
rect 24908 14310 24942 14326
rect 24908 13718 24942 13734
rect 25036 14310 25070 14326
rect 25036 13718 25070 13734
rect 25148 14310 25182 14326
rect 25148 13718 25182 13734
rect 25276 14310 25310 14326
rect 25276 13718 25310 13734
rect 25388 14310 25422 14326
rect 25388 13718 25422 13734
rect 25516 14310 25550 14326
rect 25516 13718 25550 13734
rect 25628 14310 25662 14326
rect 25628 13718 25662 13734
rect 25756 14310 25790 14326
rect 25756 13718 25790 13734
rect 25868 14310 25902 14326
rect 25868 13718 25902 13734
rect 25996 14310 26030 14326
rect 25996 13718 26030 13734
rect 26108 14310 26142 14326
rect 26108 13718 26142 13734
rect 26236 14310 26270 14326
rect 26236 13718 26270 13734
rect 26348 14310 26382 14326
rect 26348 13718 26382 13734
rect 26476 14310 26510 14326
rect 26476 13718 26510 13734
rect 26588 14310 26622 14326
rect 26588 13718 26622 13734
rect 26716 14310 26750 14326
rect 26716 13718 26750 13734
rect 26828 14310 26862 14326
rect 26828 13718 26862 13734
rect 26956 14310 26990 14326
rect 26956 13718 26990 13734
rect 27068 14310 27102 14326
rect 27068 13718 27102 13734
rect 27196 14310 27230 14326
rect 27196 13718 27230 13734
rect 27308 14310 27342 14326
rect 27308 13718 27342 13734
rect 27436 14310 27470 14326
rect 27436 13718 27470 13734
rect 27548 14310 27582 14326
rect 27548 13718 27582 13734
rect 27676 14310 27710 14326
rect 27676 13718 27710 13734
rect 27788 14310 27822 14326
rect 27788 13718 27822 13734
rect 27916 14310 27950 14326
rect 27916 13718 27950 13734
rect 28028 14310 28062 14326
rect 28028 13718 28062 13734
rect 28156 14310 28190 14326
rect 28156 13718 28190 13734
rect 28268 14310 28302 14326
rect 28268 13718 28302 13734
rect 28396 14310 28430 14326
rect 28396 13718 28430 13734
rect 28508 14310 28542 14326
rect 28508 13718 28542 13734
rect 28636 14310 28670 14326
rect 28636 13718 28670 13734
rect 28748 14310 28782 14326
rect 28748 13718 28782 13734
rect 28876 14310 28910 14326
rect 28876 13718 28910 13734
rect 28988 14310 29022 14326
rect 28988 13718 29022 13734
rect 29116 14310 29150 14326
rect 29116 13718 29150 13734
rect 29228 14310 29262 14326
rect 29228 13718 29262 13734
rect 29356 14310 29390 14326
rect 29356 13718 29390 13734
rect 19914 13552 19930 13684
rect 19968 13552 20170 13684
rect 20208 13552 20410 13684
rect 20448 13552 20650 13684
rect 20688 13552 20890 13684
rect 20928 13552 21130 13684
rect 21168 13552 21370 13684
rect 21408 13552 21610 13684
rect 21648 13552 21850 13684
rect 21888 13552 22090 13684
rect 22128 13552 22330 13684
rect 22368 13552 22570 13684
rect 22608 13552 22810 13684
rect 22848 13552 23050 13684
rect 23088 13552 23290 13684
rect 23328 13552 23530 13684
rect 23568 13552 23770 13684
rect 23808 13552 24010 13684
rect 24048 13552 24250 13684
rect 24288 13552 24490 13684
rect 24528 13552 24730 13684
rect 24768 13552 24970 13684
rect 25008 13552 25210 13684
rect 25248 13552 25450 13684
rect 25488 13552 25690 13684
rect 25728 13552 25930 13684
rect 25968 13552 26170 13684
rect 26208 13552 26410 13684
rect 26448 13552 26650 13684
rect 26688 13552 26890 13684
rect 26928 13552 27130 13684
rect 27168 13552 27370 13684
rect 27408 13552 27610 13684
rect 27648 13552 27850 13684
rect 27888 13552 28090 13684
rect 28128 13552 28330 13684
rect 28368 13552 28570 13684
rect 28608 13552 28810 13684
rect 28848 13552 29050 13684
rect 29088 13552 29290 13684
rect 29328 13552 29354 13684
rect 19522 13208 19556 13296
rect 29702 13208 29736 13296
rect 10218 11510 10378 11544
rect 38900 11516 39038 11544
rect 38900 11510 39004 11516
rect 10218 11482 10252 11510
rect 10610 11193 22370 11194
rect 22770 11193 22958 11194
rect 23358 11193 23546 11194
rect 23946 11193 24134 11194
rect 24534 11193 24722 11194
rect 25122 11193 25310 11194
rect 25710 11193 25898 11194
rect 26298 11193 26486 11194
rect 26886 11193 38646 11194
rect 10610 11159 10626 11193
rect 10994 11159 11214 11193
rect 11582 11159 11802 11193
rect 12170 11159 12390 11193
rect 12758 11159 12978 11193
rect 13346 11159 13566 11193
rect 13934 11159 14154 11193
rect 14522 11159 14742 11193
rect 15110 11159 15330 11193
rect 15698 11159 15918 11193
rect 16286 11159 16506 11193
rect 16874 11159 17094 11193
rect 17462 11159 17682 11193
rect 18050 11159 18270 11193
rect 18638 11159 18858 11193
rect 19226 11159 19446 11193
rect 19814 11159 20034 11193
rect 20402 11159 20622 11193
rect 20990 11159 21210 11193
rect 21578 11159 21798 11193
rect 22166 11159 22386 11193
rect 22754 11159 22974 11193
rect 23342 11159 23562 11193
rect 23930 11159 24150 11193
rect 24518 11159 24738 11193
rect 25106 11159 25326 11193
rect 25694 11159 25914 11193
rect 26282 11159 26502 11193
rect 26870 11159 27090 11193
rect 27458 11159 27678 11193
rect 28046 11159 28266 11193
rect 28634 11159 28854 11193
rect 29222 11159 29442 11193
rect 29810 11159 30030 11193
rect 30398 11159 30618 11193
rect 30986 11159 31206 11193
rect 31574 11159 31794 11193
rect 32162 11159 32382 11193
rect 32750 11159 32970 11193
rect 33338 11159 33558 11193
rect 33926 11159 34146 11193
rect 34514 11159 34734 11193
rect 35102 11159 35322 11193
rect 35690 11159 35910 11193
rect 36278 11159 36498 11193
rect 36866 11159 37086 11193
rect 37454 11159 37674 11193
rect 38042 11159 38262 11193
rect 38630 11159 38646 11193
rect 10610 11158 22370 11159
rect 22770 11158 22958 11159
rect 23358 11158 23546 11159
rect 23946 11158 24134 11159
rect 22324 11116 22370 11158
rect 24534 11116 24722 11159
rect 25122 11158 25310 11159
rect 25710 11158 25898 11159
rect 26298 11158 26486 11159
rect 26886 11158 38646 11159
rect 26886 11116 26932 11158
rect 10564 11100 10598 11116
rect 10564 10308 10598 10324
rect 11022 11100 11056 11116
rect 11022 10308 11056 10324
rect 11152 11100 11186 11116
rect 11152 10308 11186 10324
rect 11610 11100 11644 11116
rect 11610 10308 11644 10324
rect 11740 11100 11774 11116
rect 11740 10308 11774 10324
rect 12198 11100 12232 11116
rect 12198 10308 12232 10324
rect 12328 11100 12362 11116
rect 12328 10308 12362 10324
rect 12786 11100 12820 11116
rect 12786 10308 12820 10324
rect 12916 11100 12950 11116
rect 12916 10308 12950 10324
rect 13374 11100 13408 11116
rect 13374 10308 13408 10324
rect 13504 11100 13538 11116
rect 13504 10308 13538 10324
rect 13962 11100 13996 11116
rect 13962 10308 13996 10324
rect 14092 11100 14126 11116
rect 14092 10308 14126 10324
rect 14550 11100 14584 11116
rect 14550 10308 14584 10324
rect 14680 11100 14714 11116
rect 14680 10308 14714 10324
rect 15138 11100 15172 11116
rect 15138 10308 15172 10324
rect 15268 11100 15302 11116
rect 15268 10308 15302 10324
rect 15726 11100 15760 11116
rect 15726 10308 15760 10324
rect 15856 11100 15890 11116
rect 15856 10308 15890 10324
rect 16314 11100 16348 11116
rect 16314 10308 16348 10324
rect 16444 11100 16478 11116
rect 16444 10308 16478 10324
rect 16902 11100 16936 11116
rect 16902 10308 16936 10324
rect 17032 11100 17066 11116
rect 17032 10308 17066 10324
rect 17490 11100 17524 11116
rect 17490 10308 17524 10324
rect 17620 11100 17654 11116
rect 17620 10308 17654 10324
rect 18078 11100 18112 11116
rect 18078 10308 18112 10324
rect 18208 11100 18242 11116
rect 18208 10308 18242 10324
rect 18666 11100 18700 11116
rect 18666 10308 18700 10324
rect 18796 11100 18830 11116
rect 18796 10308 18830 10324
rect 19254 11100 19288 11116
rect 19254 10308 19288 10324
rect 19384 11100 19418 11116
rect 19384 10308 19418 10324
rect 19842 11100 19876 11116
rect 19842 10308 19876 10324
rect 19972 11100 20006 11116
rect 19972 10308 20006 10324
rect 20430 11100 20464 11116
rect 20430 10308 20464 10324
rect 20560 11100 20594 11116
rect 20560 10308 20594 10324
rect 21018 11100 21052 11116
rect 21018 10308 21052 10324
rect 21148 11100 21182 11116
rect 21148 10308 21182 10324
rect 21606 11100 21640 11116
rect 21606 10308 21640 10324
rect 21736 11100 21770 11116
rect 21736 10308 21770 10324
rect 22194 11100 22228 11116
rect 22194 10308 22228 10324
rect 22324 11100 22358 11116
rect 22324 10266 22358 10324
rect 22782 11100 22816 11116
rect 22782 10308 22816 10324
rect 22912 11100 22946 11116
rect 22912 10308 22946 10324
rect 23370 11100 23404 11116
rect 23370 10308 23404 10324
rect 23500 11100 23534 11116
rect 23500 10308 23534 10324
rect 23958 11100 23992 11116
rect 23958 10308 23992 10324
rect 24088 11100 24122 11116
rect 24088 10308 24122 10324
rect 24546 11100 24710 11116
rect 24580 10324 24676 11100
rect 24546 10266 24710 10324
rect 25134 11100 25168 11116
rect 25134 10308 25168 10324
rect 25264 11100 25298 11116
rect 25264 10308 25298 10324
rect 25722 11100 25756 11116
rect 25722 10308 25756 10324
rect 25852 11100 25886 11116
rect 25852 10308 25886 10324
rect 26310 11100 26344 11116
rect 26310 10308 26344 10324
rect 26440 11100 26474 11116
rect 26440 10308 26474 10324
rect 26898 11100 26932 11116
rect 26898 10266 26932 10324
rect 27028 11100 27062 11116
rect 27028 10308 27062 10324
rect 27486 11100 27520 11116
rect 27486 10308 27520 10324
rect 27616 11100 27650 11116
rect 27616 10308 27650 10324
rect 28074 11100 28108 11116
rect 28074 10308 28108 10324
rect 28204 11100 28238 11116
rect 28204 10308 28238 10324
rect 28662 11100 28696 11116
rect 28662 10308 28696 10324
rect 28792 11100 28826 11116
rect 28792 10308 28826 10324
rect 29250 11100 29284 11116
rect 29250 10308 29284 10324
rect 29380 11100 29414 11116
rect 29380 10308 29414 10324
rect 29838 11100 29872 11116
rect 29838 10308 29872 10324
rect 29968 11100 30002 11116
rect 29968 10308 30002 10324
rect 30426 11100 30460 11116
rect 30426 10308 30460 10324
rect 30556 11100 30590 11116
rect 30556 10308 30590 10324
rect 31014 11100 31048 11116
rect 31014 10308 31048 10324
rect 31144 11100 31178 11116
rect 31144 10308 31178 10324
rect 31602 11100 31636 11116
rect 31602 10308 31636 10324
rect 31732 11100 31766 11116
rect 31732 10308 31766 10324
rect 32190 11100 32224 11116
rect 32190 10308 32224 10324
rect 32320 11100 32354 11116
rect 32320 10308 32354 10324
rect 32778 11100 32812 11116
rect 32778 10308 32812 10324
rect 32908 11100 32942 11116
rect 32908 10308 32942 10324
rect 33366 11100 33400 11116
rect 33366 10308 33400 10324
rect 33496 11100 33530 11116
rect 33496 10308 33530 10324
rect 33954 11100 33988 11116
rect 33954 10308 33988 10324
rect 34084 11100 34118 11116
rect 34084 10308 34118 10324
rect 34542 11100 34576 11116
rect 34542 10308 34576 10324
rect 34672 11100 34706 11116
rect 34672 10308 34706 10324
rect 35130 11100 35164 11116
rect 35130 10308 35164 10324
rect 35260 11100 35294 11116
rect 35260 10308 35294 10324
rect 35718 11100 35752 11116
rect 35718 10308 35752 10324
rect 35848 11100 35882 11116
rect 35848 10308 35882 10324
rect 36306 11100 36340 11116
rect 36306 10308 36340 10324
rect 36436 11100 36470 11116
rect 36436 10308 36470 10324
rect 36894 11100 36928 11116
rect 36894 10308 36928 10324
rect 37024 11100 37058 11116
rect 37024 10308 37058 10324
rect 37482 11100 37516 11116
rect 37482 10308 37516 10324
rect 37612 11100 37646 11116
rect 37612 10308 37646 10324
rect 38070 11100 38104 11116
rect 38070 10308 38104 10324
rect 38200 11100 38234 11116
rect 38200 10308 38234 10324
rect 38658 11100 38692 11116
rect 38658 10308 38692 10324
rect 10610 10265 22370 10266
rect 22770 10265 22958 10266
rect 23358 10265 23546 10266
rect 23946 10265 24134 10266
rect 24534 10265 24722 10266
rect 25122 10265 25310 10266
rect 25710 10265 25898 10266
rect 26298 10265 26486 10266
rect 26886 10265 38646 10266
rect 10610 10231 10626 10265
rect 10994 10231 11214 10265
rect 11582 10231 11802 10265
rect 12170 10231 12390 10265
rect 12758 10231 12978 10265
rect 13346 10231 13566 10265
rect 13934 10231 14154 10265
rect 14522 10231 14742 10265
rect 15110 10231 15330 10265
rect 15698 10231 15918 10265
rect 16286 10231 16506 10265
rect 16874 10231 17094 10265
rect 17462 10231 17682 10265
rect 18050 10231 18270 10265
rect 18638 10231 18858 10265
rect 19226 10231 19446 10265
rect 19814 10231 20034 10265
rect 20402 10231 20622 10265
rect 20990 10231 21210 10265
rect 21578 10231 21798 10265
rect 22166 10231 22386 10265
rect 22754 10231 22974 10265
rect 23342 10231 23562 10265
rect 23930 10231 24150 10265
rect 24518 10231 24738 10265
rect 25106 10231 25326 10265
rect 25694 10231 25914 10265
rect 26282 10231 26502 10265
rect 26870 10231 27090 10265
rect 27458 10231 27678 10265
rect 28046 10231 28266 10265
rect 28634 10231 28854 10265
rect 29222 10231 29442 10265
rect 29810 10231 30030 10265
rect 30398 10231 30618 10265
rect 30986 10231 31206 10265
rect 31574 10231 31794 10265
rect 32162 10231 32382 10265
rect 32750 10231 32970 10265
rect 33338 10231 33558 10265
rect 33926 10231 34146 10265
rect 34514 10231 34734 10265
rect 35102 10231 35322 10265
rect 35690 10231 35910 10265
rect 36278 10231 36498 10265
rect 36866 10231 37086 10265
rect 37454 10231 37674 10265
rect 38042 10231 38262 10265
rect 38630 10231 38646 10265
rect 10610 10193 22370 10231
rect 22770 10193 22958 10231
rect 23358 10230 23546 10231
rect 23358 10193 23546 10194
rect 23946 10193 24134 10231
rect 24534 10193 24722 10231
rect 25122 10193 25310 10231
rect 25710 10230 25898 10231
rect 25710 10193 25898 10194
rect 26298 10193 26486 10231
rect 26886 10193 38646 10231
rect 10610 10159 10626 10193
rect 10994 10159 11214 10193
rect 11582 10159 11802 10193
rect 12170 10159 12390 10193
rect 12758 10159 12978 10193
rect 13346 10159 13566 10193
rect 13934 10159 14154 10193
rect 14522 10159 14742 10193
rect 15110 10159 15330 10193
rect 15698 10159 15918 10193
rect 16286 10159 16506 10193
rect 16874 10159 17094 10193
rect 17462 10159 17682 10193
rect 18050 10159 18270 10193
rect 18638 10159 18858 10193
rect 19226 10159 19446 10193
rect 19814 10159 20034 10193
rect 20402 10159 20622 10193
rect 20990 10159 21210 10193
rect 21578 10159 21798 10193
rect 22166 10159 22386 10193
rect 22754 10159 22974 10193
rect 23342 10159 23562 10193
rect 23930 10159 24150 10193
rect 24518 10159 24738 10193
rect 25106 10159 25326 10193
rect 25694 10159 25914 10193
rect 26282 10159 26502 10193
rect 26870 10159 27090 10193
rect 27458 10159 27678 10193
rect 28046 10159 28266 10193
rect 28634 10159 28854 10193
rect 29222 10159 29442 10193
rect 29810 10159 30030 10193
rect 30398 10159 30618 10193
rect 30986 10159 31206 10193
rect 31574 10159 31794 10193
rect 32162 10159 32382 10193
rect 32750 10159 32970 10193
rect 33338 10159 33558 10193
rect 33926 10159 34146 10193
rect 34514 10159 34734 10193
rect 35102 10159 35322 10193
rect 35690 10159 35910 10193
rect 36278 10159 36498 10193
rect 36866 10159 37086 10193
rect 37454 10159 37674 10193
rect 38042 10159 38262 10193
rect 38630 10159 38646 10193
rect 10610 10158 22370 10159
rect 22770 10158 22958 10159
rect 23358 10158 23546 10159
rect 23946 10158 24134 10159
rect 24534 10158 24722 10159
rect 25122 10158 25310 10159
rect 25710 10158 25898 10159
rect 26298 10158 26486 10159
rect 26886 10158 38646 10159
rect 10564 10100 10598 10116
rect 10564 9308 10598 9324
rect 11022 10100 11056 10116
rect 11022 9308 11056 9324
rect 11152 10100 11186 10116
rect 11152 9308 11186 9324
rect 11610 10100 11644 10116
rect 11610 9308 11644 9324
rect 11740 10100 11774 10116
rect 11740 9308 11774 9324
rect 12198 10100 12232 10116
rect 12198 9308 12232 9324
rect 12328 10100 12362 10116
rect 12328 9308 12362 9324
rect 12786 10100 12820 10116
rect 12786 9308 12820 9324
rect 12916 10100 12950 10116
rect 12916 9308 12950 9324
rect 13374 10100 13408 10116
rect 13374 9308 13408 9324
rect 13504 10100 13538 10116
rect 13504 9308 13538 9324
rect 13962 10100 13996 10116
rect 13962 9308 13996 9324
rect 14092 10100 14126 10116
rect 14092 9308 14126 9324
rect 14550 10100 14584 10116
rect 14550 9308 14584 9324
rect 14680 10100 14714 10116
rect 14680 9308 14714 9324
rect 15138 10100 15172 10116
rect 15138 9308 15172 9324
rect 15268 10100 15302 10116
rect 15268 9308 15302 9324
rect 15726 10100 15760 10116
rect 15726 9308 15760 9324
rect 15856 10100 15890 10116
rect 15856 9308 15890 9324
rect 16314 10100 16348 10116
rect 16314 9308 16348 9324
rect 16444 10100 16478 10116
rect 16444 9308 16478 9324
rect 16902 10100 16936 10116
rect 16902 9308 16936 9324
rect 17032 10100 17066 10116
rect 17032 9308 17066 9324
rect 17490 10100 17524 10116
rect 17490 9308 17524 9324
rect 17620 10100 17654 10116
rect 17620 9308 17654 9324
rect 18078 10100 18112 10116
rect 18078 9308 18112 9324
rect 18208 10100 18242 10116
rect 18208 9308 18242 9324
rect 18666 10100 18700 10116
rect 18666 9308 18700 9324
rect 18796 10100 18830 10116
rect 18796 9308 18830 9324
rect 19254 10100 19288 10116
rect 19254 9308 19288 9324
rect 19384 10100 19418 10116
rect 19384 9308 19418 9324
rect 19842 10100 19876 10116
rect 19842 9308 19876 9324
rect 19972 10100 20006 10116
rect 19972 9308 20006 9324
rect 20430 10100 20464 10116
rect 20430 9308 20464 9324
rect 20560 10100 20594 10116
rect 20560 9308 20594 9324
rect 21018 10100 21052 10116
rect 21018 9308 21052 9324
rect 21148 10100 21182 10116
rect 21148 9308 21182 9324
rect 21606 10100 21640 10116
rect 21606 9308 21640 9324
rect 21736 10100 21770 10116
rect 21736 9308 21770 9324
rect 22194 10100 22228 10116
rect 22194 9308 22228 9324
rect 22324 10100 22358 10158
rect 22324 9266 22358 9324
rect 22782 10100 22816 10116
rect 22782 9308 22816 9324
rect 22912 10100 22946 10116
rect 22912 9308 22946 9324
rect 23370 10100 23404 10116
rect 23370 9308 23404 9324
rect 23500 10100 23534 10116
rect 23500 9308 23534 9324
rect 23958 10100 23992 10116
rect 23958 9308 23992 9324
rect 24088 10100 24122 10116
rect 24088 9308 24122 9324
rect 24546 10100 24710 10158
rect 24580 9324 24676 10100
rect 24546 9266 24710 9324
rect 25134 10100 25168 10116
rect 25134 9308 25168 9324
rect 25264 10100 25298 10116
rect 25264 9308 25298 9324
rect 25722 10100 25756 10116
rect 25722 9308 25756 9324
rect 25852 10100 25886 10116
rect 25852 9308 25886 9324
rect 26310 10100 26344 10116
rect 26310 9308 26344 9324
rect 26440 10100 26474 10116
rect 26440 9308 26474 9324
rect 26898 10100 26932 10158
rect 26898 9266 26932 9324
rect 27028 10100 27062 10116
rect 27028 9308 27062 9324
rect 27486 10100 27520 10116
rect 27486 9308 27520 9324
rect 27616 10100 27650 10116
rect 27616 9308 27650 9324
rect 28074 10100 28108 10116
rect 28074 9308 28108 9324
rect 28204 10100 28238 10116
rect 28204 9308 28238 9324
rect 28662 10100 28696 10116
rect 28662 9308 28696 9324
rect 28792 10100 28826 10116
rect 28792 9308 28826 9324
rect 29250 10100 29284 10116
rect 29250 9308 29284 9324
rect 29380 10100 29414 10116
rect 29380 9308 29414 9324
rect 29838 10100 29872 10116
rect 29838 9308 29872 9324
rect 29968 10100 30002 10116
rect 29968 9308 30002 9324
rect 30426 10100 30460 10116
rect 30426 9308 30460 9324
rect 30556 10100 30590 10116
rect 30556 9308 30590 9324
rect 31014 10100 31048 10116
rect 31014 9308 31048 9324
rect 31144 10100 31178 10116
rect 31144 9308 31178 9324
rect 31602 10100 31636 10116
rect 31602 9308 31636 9324
rect 31732 10100 31766 10116
rect 31732 9308 31766 9324
rect 32190 10100 32224 10116
rect 32190 9308 32224 9324
rect 32320 10100 32354 10116
rect 32320 9308 32354 9324
rect 32778 10100 32812 10116
rect 32778 9308 32812 9324
rect 32908 10100 32942 10116
rect 32908 9308 32942 9324
rect 33366 10100 33400 10116
rect 33366 9308 33400 9324
rect 33496 10100 33530 10116
rect 33496 9308 33530 9324
rect 33954 10100 33988 10116
rect 33954 9308 33988 9324
rect 34084 10100 34118 10116
rect 34084 9308 34118 9324
rect 34542 10100 34576 10116
rect 34542 9308 34576 9324
rect 34672 10100 34706 10116
rect 34672 9308 34706 9324
rect 35130 10100 35164 10116
rect 35130 9308 35164 9324
rect 35260 10100 35294 10116
rect 35260 9308 35294 9324
rect 35718 10100 35752 10116
rect 35718 9308 35752 9324
rect 35848 10100 35882 10116
rect 35848 9308 35882 9324
rect 36306 10100 36340 10116
rect 36306 9308 36340 9324
rect 36436 10100 36470 10116
rect 36436 9308 36470 9324
rect 36894 10100 36928 10116
rect 36894 9308 36928 9324
rect 37024 10100 37058 10116
rect 37024 9308 37058 9324
rect 37482 10100 37516 10116
rect 37482 9308 37516 9324
rect 37612 10100 37646 10116
rect 37612 9308 37646 9324
rect 38070 10100 38104 10116
rect 38070 9308 38104 9324
rect 38200 10100 38234 10116
rect 38200 9308 38234 9324
rect 38658 10100 38692 10116
rect 38658 9308 38692 9324
rect 10610 9265 22370 9266
rect 22770 9265 22958 9266
rect 23358 9265 23546 9266
rect 23946 9265 24134 9266
rect 24534 9265 24722 9266
rect 25122 9265 25310 9266
rect 25710 9265 25898 9266
rect 26298 9265 26486 9266
rect 26886 9265 38646 9266
rect 10610 9231 10626 9265
rect 10994 9231 11214 9265
rect 11582 9231 11802 9265
rect 12170 9231 12390 9265
rect 12758 9231 12978 9265
rect 13346 9231 13566 9265
rect 13934 9231 14154 9265
rect 14522 9231 14742 9265
rect 15110 9231 15330 9265
rect 15698 9231 15918 9265
rect 16286 9231 16506 9265
rect 16874 9231 17094 9265
rect 17462 9231 17682 9265
rect 18050 9231 18270 9265
rect 18638 9231 18858 9265
rect 19226 9231 19446 9265
rect 19814 9231 20034 9265
rect 20402 9231 20622 9265
rect 20990 9231 21210 9265
rect 21578 9231 21798 9265
rect 22166 9231 22386 9265
rect 22754 9231 22974 9265
rect 23342 9231 23562 9265
rect 23930 9231 24150 9265
rect 24518 9231 24738 9265
rect 25106 9231 25326 9265
rect 25694 9231 25914 9265
rect 26282 9231 26502 9265
rect 26870 9231 27090 9265
rect 27458 9231 27678 9265
rect 28046 9231 28266 9265
rect 28634 9231 28854 9265
rect 29222 9231 29442 9265
rect 29810 9231 30030 9265
rect 30398 9231 30618 9265
rect 30986 9231 31206 9265
rect 31574 9231 31794 9265
rect 32162 9231 32382 9265
rect 32750 9231 32970 9265
rect 33338 9231 33558 9265
rect 33926 9231 34146 9265
rect 34514 9231 34734 9265
rect 35102 9231 35322 9265
rect 35690 9231 35910 9265
rect 36278 9231 36498 9265
rect 36866 9231 37086 9265
rect 37454 9231 37674 9265
rect 38042 9231 38262 9265
rect 38630 9231 38646 9265
rect 10610 9193 22370 9231
rect 22770 9193 22958 9231
rect 23358 9230 23546 9231
rect 23358 9193 23546 9194
rect 23946 9193 24134 9231
rect 24534 9193 24722 9231
rect 25122 9193 25310 9231
rect 25710 9230 25898 9231
rect 25710 9193 25898 9194
rect 26298 9193 26486 9231
rect 26886 9193 38646 9231
rect 10610 9159 10626 9193
rect 10994 9159 11214 9193
rect 11582 9159 11802 9193
rect 12170 9159 12390 9193
rect 12758 9159 12978 9193
rect 13346 9159 13566 9193
rect 13934 9159 14154 9193
rect 14522 9159 14742 9193
rect 15110 9159 15330 9193
rect 15698 9159 15918 9193
rect 16286 9159 16506 9193
rect 16874 9159 17094 9193
rect 17462 9159 17682 9193
rect 18050 9159 18270 9193
rect 18638 9159 18858 9193
rect 19226 9159 19446 9193
rect 19814 9159 20034 9193
rect 20402 9159 20622 9193
rect 20990 9159 21210 9193
rect 21578 9159 21798 9193
rect 22166 9159 22386 9193
rect 22754 9159 22974 9193
rect 23342 9159 23562 9193
rect 23930 9159 24150 9193
rect 24518 9159 24738 9193
rect 25106 9159 25326 9193
rect 25694 9159 25914 9193
rect 26282 9159 26502 9193
rect 26870 9159 27090 9193
rect 27458 9159 27678 9193
rect 28046 9159 28266 9193
rect 28634 9159 28854 9193
rect 29222 9159 29442 9193
rect 29810 9159 30030 9193
rect 30398 9159 30618 9193
rect 30986 9159 31206 9193
rect 31574 9159 31794 9193
rect 32162 9159 32382 9193
rect 32750 9159 32970 9193
rect 33338 9159 33558 9193
rect 33926 9159 34146 9193
rect 34514 9159 34734 9193
rect 35102 9159 35322 9193
rect 35690 9159 35910 9193
rect 36278 9159 36498 9193
rect 36866 9159 37086 9193
rect 37454 9159 37674 9193
rect 38042 9159 38262 9193
rect 38630 9159 38646 9193
rect 10610 9158 22370 9159
rect 22770 9158 22958 9159
rect 23358 9158 23546 9159
rect 23946 9158 24134 9159
rect 24534 9158 24722 9159
rect 25122 9158 25310 9159
rect 25710 9158 25898 9159
rect 26298 9158 26486 9159
rect 26886 9158 38646 9159
rect 10564 9100 10598 9116
rect 10564 8308 10598 8324
rect 11022 9100 11056 9116
rect 11022 8308 11056 8324
rect 11152 9100 11186 9116
rect 11152 8308 11186 8324
rect 11610 9100 11644 9116
rect 11610 8308 11644 8324
rect 11740 9100 11774 9116
rect 11740 8308 11774 8324
rect 12198 9100 12232 9116
rect 12198 8308 12232 8324
rect 12328 9100 12362 9116
rect 12328 8308 12362 8324
rect 12786 9100 12820 9116
rect 12786 8308 12820 8324
rect 12916 9100 12950 9116
rect 12916 8308 12950 8324
rect 13374 9100 13408 9116
rect 13374 8308 13408 8324
rect 13504 9100 13538 9116
rect 13504 8308 13538 8324
rect 13962 9100 13996 9116
rect 13962 8308 13996 8324
rect 14092 9100 14126 9116
rect 14092 8308 14126 8324
rect 14550 9100 14584 9116
rect 14550 8308 14584 8324
rect 14680 9100 14714 9116
rect 14680 8308 14714 8324
rect 15138 9100 15172 9116
rect 15138 8308 15172 8324
rect 15268 9100 15302 9116
rect 15268 8308 15302 8324
rect 15726 9100 15760 9116
rect 15726 8308 15760 8324
rect 15856 9100 15890 9116
rect 15856 8308 15890 8324
rect 16314 9100 16348 9116
rect 16314 8308 16348 8324
rect 16444 9100 16478 9116
rect 16444 8308 16478 8324
rect 16902 9100 16936 9116
rect 16902 8308 16936 8324
rect 17032 9100 17066 9116
rect 17032 8308 17066 8324
rect 17490 9100 17524 9116
rect 17490 8308 17524 8324
rect 17620 9100 17654 9116
rect 17620 8308 17654 8324
rect 18078 9100 18112 9116
rect 18078 8308 18112 8324
rect 18208 9100 18242 9116
rect 18208 8308 18242 8324
rect 18666 9100 18700 9116
rect 18666 8308 18700 8324
rect 18796 9100 18830 9116
rect 18796 8308 18830 8324
rect 19254 9100 19288 9116
rect 19254 8308 19288 8324
rect 19384 9100 19418 9116
rect 19384 8308 19418 8324
rect 19842 9100 19876 9116
rect 19842 8308 19876 8324
rect 19972 9100 20006 9116
rect 19972 8308 20006 8324
rect 20430 9100 20464 9116
rect 20430 8308 20464 8324
rect 20560 9100 20594 9116
rect 20560 8308 20594 8324
rect 21018 9100 21052 9116
rect 21018 8308 21052 8324
rect 21148 9100 21182 9116
rect 21148 8308 21182 8324
rect 21606 9100 21640 9116
rect 21606 8308 21640 8324
rect 21736 9100 21770 9116
rect 21736 8308 21770 8324
rect 22194 9100 22228 9116
rect 22194 8308 22228 8324
rect 22324 9100 22358 9158
rect 22324 8308 22358 8324
rect 22782 9100 22816 9116
rect 22782 8308 22816 8324
rect 22912 9100 22946 9116
rect 22912 8308 22946 8324
rect 23370 9100 23404 9116
rect 23370 8308 23404 8324
rect 23500 9100 23534 9116
rect 23500 8308 23534 8324
rect 23958 9100 23992 9116
rect 23958 8308 23992 8324
rect 24088 9100 24122 9116
rect 24088 8308 24122 8324
rect 24546 9100 24710 9158
rect 24580 8324 24676 9100
rect 24546 8308 24710 8324
rect 25134 9100 25168 9116
rect 25134 8308 25168 8324
rect 25264 9100 25298 9116
rect 25264 8308 25298 8324
rect 25722 9100 25756 9116
rect 25722 8308 25756 8324
rect 25852 9100 25886 9116
rect 25852 8308 25886 8324
rect 26310 9100 26344 9116
rect 26310 8308 26344 8324
rect 26440 9100 26474 9116
rect 26440 8308 26474 8324
rect 26898 9100 26932 9158
rect 26898 8308 26932 8324
rect 27028 9100 27062 9116
rect 27028 8308 27062 8324
rect 27486 9100 27520 9116
rect 27486 8308 27520 8324
rect 27616 9100 27650 9116
rect 27616 8308 27650 8324
rect 28074 9100 28108 9116
rect 28074 8308 28108 8324
rect 28204 9100 28238 9116
rect 28204 8308 28238 8324
rect 28662 9100 28696 9116
rect 28662 8308 28696 8324
rect 28792 9100 28826 9116
rect 28792 8308 28826 8324
rect 29250 9100 29284 9116
rect 29250 8308 29284 8324
rect 29380 9100 29414 9116
rect 29380 8308 29414 8324
rect 29838 9100 29872 9116
rect 29838 8308 29872 8324
rect 29968 9100 30002 9116
rect 29968 8308 30002 8324
rect 30426 9100 30460 9116
rect 30426 8308 30460 8324
rect 30556 9100 30590 9116
rect 30556 8308 30590 8324
rect 31014 9100 31048 9116
rect 31014 8308 31048 8324
rect 31144 9100 31178 9116
rect 31144 8308 31178 8324
rect 31602 9100 31636 9116
rect 31602 8308 31636 8324
rect 31732 9100 31766 9116
rect 31732 8308 31766 8324
rect 32190 9100 32224 9116
rect 32190 8308 32224 8324
rect 32320 9100 32354 9116
rect 32320 8308 32354 8324
rect 32778 9100 32812 9116
rect 32778 8308 32812 8324
rect 32908 9100 32942 9116
rect 32908 8308 32942 8324
rect 33366 9100 33400 9116
rect 33366 8308 33400 8324
rect 33496 9100 33530 9116
rect 33496 8308 33530 8324
rect 33954 9100 33988 9116
rect 33954 8308 33988 8324
rect 34084 9100 34118 9116
rect 34084 8308 34118 8324
rect 34542 9100 34576 9116
rect 34542 8308 34576 8324
rect 34672 9100 34706 9116
rect 34672 8308 34706 8324
rect 35130 9100 35164 9116
rect 35130 8308 35164 8324
rect 35260 9100 35294 9116
rect 35260 8308 35294 8324
rect 35718 9100 35752 9116
rect 35718 8308 35752 8324
rect 35848 9100 35882 9116
rect 35848 8308 35882 8324
rect 36306 9100 36340 9116
rect 36306 8308 36340 8324
rect 36436 9100 36470 9116
rect 36436 8308 36470 8324
rect 36894 9100 36928 9116
rect 36894 8308 36928 8324
rect 37024 9100 37058 9116
rect 37024 8308 37058 8324
rect 37482 9100 37516 9116
rect 37482 8308 37516 8324
rect 37612 9100 37646 9116
rect 37612 8308 37646 8324
rect 38070 9100 38104 9116
rect 38070 8308 38104 8324
rect 38200 9100 38234 9116
rect 38200 8308 38234 8324
rect 38658 9100 38692 9116
rect 38658 8308 38692 8324
rect 22324 8266 22370 8308
rect 10610 8265 22370 8266
rect 22770 8265 22958 8266
rect 23358 8265 23546 8266
rect 23946 8265 24134 8266
rect 24534 8265 24722 8308
rect 26886 8266 26932 8308
rect 25122 8265 25310 8266
rect 25710 8265 25898 8266
rect 26298 8265 26486 8266
rect 26886 8265 38646 8266
rect 10610 8231 10626 8265
rect 10994 8231 11214 8265
rect 11582 8231 11802 8265
rect 12170 8231 12390 8265
rect 12758 8231 12978 8265
rect 13346 8231 13566 8265
rect 13934 8231 14154 8265
rect 14522 8231 14742 8265
rect 15110 8231 15330 8265
rect 15698 8231 15918 8265
rect 16286 8231 16506 8265
rect 16874 8231 17094 8265
rect 17462 8231 17682 8265
rect 18050 8231 18270 8265
rect 18638 8231 18858 8265
rect 19226 8231 19446 8265
rect 19814 8231 20034 8265
rect 20402 8231 20622 8265
rect 20990 8231 21210 8265
rect 21578 8231 21798 8265
rect 22166 8231 22386 8265
rect 22754 8231 22974 8265
rect 23342 8231 23562 8265
rect 23930 8231 24150 8265
rect 24518 8231 24738 8265
rect 25106 8231 25326 8265
rect 25694 8231 25914 8265
rect 26282 8231 26502 8265
rect 26870 8231 27090 8265
rect 27458 8231 27678 8265
rect 28046 8231 28266 8265
rect 28634 8231 28854 8265
rect 29222 8231 29442 8265
rect 29810 8231 30030 8265
rect 30398 8231 30618 8265
rect 30986 8231 31206 8265
rect 31574 8231 31794 8265
rect 32162 8231 32382 8265
rect 32750 8231 32970 8265
rect 33338 8231 33558 8265
rect 33926 8231 34146 8265
rect 34514 8231 34734 8265
rect 35102 8231 35322 8265
rect 35690 8231 35910 8265
rect 36278 8231 36498 8265
rect 36866 8231 37086 8265
rect 37454 8231 37674 8265
rect 38042 8231 38262 8265
rect 38630 8231 38646 8265
rect 10610 8230 22370 8231
rect 22770 8230 22958 8231
rect 23358 8230 23546 8231
rect 23946 8230 24134 8231
rect 24534 8230 24722 8231
rect 25122 8230 25310 8231
rect 25710 8230 25898 8231
rect 26298 8230 26486 8231
rect 26886 8230 38646 8231
rect 10218 7914 10252 7934
rect 39004 7914 39038 7968
rect 10218 7880 10336 7914
rect 38950 7880 39038 7914
rect 23920 7852 23946 7880
rect 24134 7852 24164 7880
rect 23920 7170 24164 7852
rect 25094 7852 25122 7880
rect 25310 7852 25338 7880
rect 25094 7170 25338 7852
rect 23230 7136 23264 7170
rect 25992 7136 26026 7170
rect 23662 6704 23678 6836
rect 23716 6704 23944 6836
rect 23982 6704 24000 6836
rect 24194 6704 24210 6836
rect 24248 6704 24476 6836
rect 24514 6704 24532 6836
rect 24726 6704 24742 6836
rect 24780 6704 25008 6836
rect 25046 6704 25064 6836
rect 25258 6704 25274 6836
rect 25312 6704 25540 6836
rect 25578 6704 25596 6836
rect 23616 6654 23650 6670
rect 23616 5862 23650 5878
rect 23744 6654 23778 6670
rect 23744 5862 23778 5878
rect 23882 6654 23916 6670
rect 23882 5862 23916 5878
rect 24010 6654 24044 6670
rect 24010 5862 24044 5878
rect 24148 6654 24182 6670
rect 24148 5862 24182 5878
rect 24276 6654 24310 6670
rect 24276 5862 24310 5878
rect 24414 6654 24448 6670
rect 24414 5862 24448 5878
rect 24542 6654 24576 6670
rect 24542 5862 24576 5878
rect 24680 6654 24714 6670
rect 24680 5862 24714 5878
rect 24808 6654 24842 6670
rect 24808 5862 24842 5878
rect 24946 6654 24980 6670
rect 24946 5862 24980 5878
rect 25074 6654 25108 6670
rect 25074 5862 25108 5878
rect 25212 6654 25246 6670
rect 25212 5862 25246 5878
rect 25340 6654 25374 6670
rect 25340 5862 25374 5878
rect 25478 6654 25512 6670
rect 25478 5862 25512 5878
rect 25606 6654 25640 6670
rect 25606 5862 25640 5878
rect 23662 5694 23678 5826
rect 23716 5694 23944 5826
rect 23982 5694 24000 5826
rect 24194 5694 24210 5826
rect 24248 5694 24476 5826
rect 24514 5694 24532 5826
rect 24726 5694 24742 5826
rect 24780 5694 25008 5826
rect 25046 5694 25064 5826
rect 25258 5694 25274 5826
rect 25312 5694 25540 5826
rect 25578 5694 25596 5826
rect 23616 5644 23650 5660
rect 23616 4852 23650 4868
rect 23744 5644 23778 5660
rect 23744 4852 23778 4868
rect 23882 5644 23916 5660
rect 23882 4852 23916 4868
rect 24010 5644 24044 5660
rect 24010 4852 24044 4868
rect 24148 5644 24182 5660
rect 24148 4852 24182 4868
rect 24276 5644 24310 5660
rect 24276 4852 24310 4868
rect 24414 5644 24448 5660
rect 24414 4852 24448 4868
rect 24542 5644 24576 5660
rect 24542 4852 24576 4868
rect 24680 5644 24714 5660
rect 24680 4852 24714 4868
rect 24808 5644 24842 5660
rect 24808 4852 24842 4868
rect 24946 5644 24980 5660
rect 24946 4852 24980 4868
rect 25074 5644 25108 5660
rect 25074 4852 25108 4868
rect 25212 5644 25246 5660
rect 25212 4852 25246 4868
rect 25340 5644 25374 5660
rect 25340 4852 25374 4868
rect 25478 5644 25512 5660
rect 25478 4852 25512 4868
rect 25606 5644 25640 5660
rect 25606 4852 25640 4868
rect 23662 4684 23678 4816
rect 23716 4684 23944 4816
rect 23982 4684 24000 4816
rect 24194 4684 24210 4816
rect 24248 4684 24476 4816
rect 24514 4684 24532 4816
rect 24726 4684 24742 4816
rect 24780 4684 25008 4816
rect 25046 4684 25064 4816
rect 25258 4684 25274 4816
rect 25312 4684 25540 4816
rect 25578 4684 25596 4816
rect 23616 4634 23650 4650
rect 23616 3842 23650 3858
rect 23744 4634 23778 4650
rect 23744 3842 23778 3858
rect 23882 4634 23916 4650
rect 23882 3842 23916 3858
rect 24010 4634 24044 4650
rect 24010 3842 24044 3858
rect 24148 4634 24182 4650
rect 24148 3842 24182 3858
rect 24276 4634 24310 4650
rect 24276 3842 24310 3858
rect 24414 4634 24448 4650
rect 24414 3842 24448 3858
rect 24542 4634 24576 4650
rect 24542 3842 24576 3858
rect 24680 4634 24714 4650
rect 24680 3842 24714 3858
rect 24808 4634 24842 4650
rect 24808 3842 24842 3858
rect 24946 4634 24980 4650
rect 24946 3842 24980 3858
rect 25074 4634 25108 4650
rect 25074 3842 25108 3858
rect 25212 4634 25246 4650
rect 25212 3842 25246 3858
rect 25340 4634 25374 4650
rect 25340 3842 25374 3858
rect 25478 4634 25512 4650
rect 25478 3842 25512 3858
rect 25606 4634 25640 4650
rect 25606 3842 25640 3858
rect 23662 3674 23678 3806
rect 23716 3674 23944 3806
rect 23982 3674 24000 3806
rect 24194 3674 24210 3806
rect 24248 3674 24476 3806
rect 24514 3674 24532 3806
rect 24726 3674 24742 3806
rect 24780 3674 25008 3806
rect 25046 3674 25064 3806
rect 25258 3674 25274 3806
rect 25312 3674 25540 3806
rect 25578 3674 25596 3806
rect 30651 5255 30747 5289
rect 30885 5255 30981 5289
rect 30651 5193 30685 5255
rect 30947 5193 30981 5255
rect 30651 3639 30685 3701
rect 30981 4534 31244 4554
rect 30981 4074 31086 4534
rect 31226 4074 31244 4534
rect 30981 4052 31244 4074
rect 30947 3639 30981 3701
rect 30651 3605 30747 3639
rect 30885 3605 30981 3639
rect 23230 3340 23264 3374
rect 25992 3340 26026 3374
rect 23842 2944 23988 2978
rect 25198 2944 25416 2978
rect 24188 2638 25070 2644
rect 24188 2512 24250 2638
rect 24288 2512 24490 2638
rect 24528 2512 24730 2638
rect 24768 2512 24970 2638
rect 25008 2512 25070 2638
rect 24188 2462 24222 2512
rect 24188 1836 24222 1886
rect 24316 2462 24350 2478
rect 24316 1870 24350 1886
rect 24428 2462 24462 2478
rect 24428 1870 24462 1886
rect 24556 2462 24590 2478
rect 24556 1870 24590 1886
rect 24668 2462 24702 2478
rect 24668 1870 24702 1886
rect 24796 2462 24830 2478
rect 24796 1870 24830 1886
rect 24908 2462 24942 2478
rect 24908 1870 24942 1886
rect 25036 2462 25070 2512
rect 25036 1836 25070 1886
rect 24188 1704 24250 1836
rect 24288 1704 24490 1836
rect 24528 1704 24730 1836
rect 24768 1704 24970 1836
rect 25008 1704 25070 1836
rect 24188 1654 24222 1704
rect 24188 1028 24222 1078
rect 24316 1654 24350 1670
rect 24316 1062 24350 1078
rect 24428 1654 24462 1670
rect 24428 1062 24462 1078
rect 24556 1654 24590 1670
rect 24556 1062 24590 1078
rect 24668 1654 24702 1670
rect 24668 1062 24702 1078
rect 24796 1654 24830 1670
rect 24796 1062 24830 1078
rect 24908 1654 24942 1670
rect 24908 1062 24942 1078
rect 25036 1654 25070 1704
rect 25036 1028 25070 1078
rect 24188 896 24250 1028
rect 24288 896 24490 1028
rect 24528 896 24730 1028
rect 24768 896 24970 1028
rect 25008 896 25070 1028
rect 23842 562 23940 596
rect 25292 562 25416 596
<< viali >>
rect 20014 15610 20124 15644
rect 20494 15610 20604 15644
rect 20974 15610 21084 15644
rect 21454 15610 21564 15644
rect 21934 15610 22044 15644
rect 22414 15610 22524 15644
rect 22894 15610 23004 15644
rect 23374 15610 23484 15644
rect 23854 15610 23964 15644
rect 24334 15610 24444 15644
rect 24814 15610 24924 15644
rect 25294 15610 25404 15644
rect 25774 15610 25884 15644
rect 26254 15610 26364 15644
rect 26734 15610 26844 15644
rect 27214 15610 27324 15644
rect 27694 15610 27804 15644
rect 28174 15610 28284 15644
rect 28654 15610 28764 15644
rect 29134 15610 29244 15644
rect 20014 15572 20124 15610
rect 20494 15572 20604 15610
rect 20974 15572 21084 15610
rect 21454 15572 21564 15610
rect 21934 15572 22044 15610
rect 22414 15572 22524 15610
rect 22894 15572 23004 15610
rect 23374 15572 23484 15610
rect 23854 15572 23964 15610
rect 24334 15572 24444 15610
rect 24814 15572 24924 15610
rect 25294 15572 25404 15610
rect 25774 15572 25884 15610
rect 26254 15572 26364 15610
rect 26734 15572 26844 15610
rect 27214 15572 27324 15610
rect 27694 15572 27804 15610
rect 28174 15572 28284 15610
rect 28654 15572 28764 15610
rect 29134 15572 29244 15610
rect 19930 15168 19968 15300
rect 20170 15168 20208 15300
rect 20410 15168 20448 15300
rect 20650 15168 20688 15300
rect 20890 15168 20928 15300
rect 21130 15168 21168 15300
rect 21370 15168 21408 15300
rect 21610 15168 21648 15300
rect 21850 15168 21888 15300
rect 22090 15168 22128 15300
rect 22330 15168 22368 15300
rect 22570 15168 22608 15300
rect 22810 15168 22848 15300
rect 23050 15168 23088 15300
rect 23290 15168 23328 15300
rect 23530 15168 23568 15300
rect 23770 15168 23808 15300
rect 24010 15168 24048 15300
rect 24250 15168 24288 15300
rect 24490 15168 24528 15300
rect 24730 15168 24768 15300
rect 24970 15168 25008 15300
rect 25210 15168 25248 15300
rect 25450 15168 25488 15300
rect 25690 15168 25728 15300
rect 25930 15168 25968 15300
rect 26170 15168 26208 15300
rect 26410 15168 26448 15300
rect 26650 15168 26688 15300
rect 26890 15168 26928 15300
rect 27130 15168 27168 15300
rect 27370 15168 27408 15300
rect 27610 15168 27648 15300
rect 27850 15168 27888 15300
rect 28090 15168 28128 15300
rect 28330 15168 28368 15300
rect 28570 15168 28608 15300
rect 28810 15168 28848 15300
rect 29050 15168 29088 15300
rect 29290 15168 29328 15300
rect 19868 14542 19902 15118
rect 19996 14542 20030 15118
rect 20108 14542 20142 15118
rect 20236 14542 20270 15118
rect 20348 14542 20382 15118
rect 20476 14542 20510 15118
rect 20588 14542 20622 15118
rect 20716 14542 20750 15118
rect 20828 14542 20862 15118
rect 20956 14542 20990 15118
rect 21068 14542 21102 15118
rect 21196 14542 21230 15118
rect 21308 14542 21342 15118
rect 21436 14542 21470 15118
rect 21548 14542 21582 15118
rect 21676 14542 21710 15118
rect 21788 14542 21822 15118
rect 21916 14542 21950 15118
rect 22028 14542 22062 15118
rect 22156 14542 22190 15118
rect 22268 14542 22302 15118
rect 22396 14542 22430 15118
rect 22508 14542 22542 15118
rect 22636 14542 22670 15118
rect 22748 14542 22782 15118
rect 22876 14542 22910 15118
rect 22988 14542 23022 15118
rect 23116 14542 23150 15118
rect 23228 14542 23262 15118
rect 23356 14542 23390 15118
rect 23468 14542 23502 15118
rect 23596 14542 23630 15118
rect 23708 14542 23742 15118
rect 23836 14542 23870 15118
rect 23948 14542 23982 15118
rect 24076 14542 24110 15118
rect 24188 14542 24222 15118
rect 24316 14542 24350 15118
rect 24428 14542 24462 15118
rect 24556 14542 24590 15118
rect 24668 14542 24702 15118
rect 24796 14542 24830 15118
rect 24908 14542 24942 15118
rect 25036 14542 25070 15118
rect 25148 14542 25182 15118
rect 25276 14542 25310 15118
rect 25388 14542 25422 15118
rect 25516 14542 25550 15118
rect 25628 14542 25662 15118
rect 25756 14542 25790 15118
rect 25868 14542 25902 15118
rect 25996 14542 26030 15118
rect 26108 14542 26142 15118
rect 26236 14542 26270 15118
rect 26348 14542 26382 15118
rect 26476 14542 26510 15118
rect 26588 14542 26622 15118
rect 26716 14542 26750 15118
rect 26828 14542 26862 15118
rect 26956 14542 26990 15118
rect 27068 14542 27102 15118
rect 27196 14542 27230 15118
rect 27308 14542 27342 15118
rect 27436 14542 27470 15118
rect 27548 14542 27582 15118
rect 27676 14542 27710 15118
rect 27788 14542 27822 15118
rect 27916 14542 27950 15118
rect 28028 14542 28062 15118
rect 28156 14542 28190 15118
rect 28268 14542 28302 15118
rect 28396 14542 28430 15118
rect 28508 14542 28542 15118
rect 28636 14542 28670 15118
rect 28748 14542 28782 15118
rect 28876 14542 28910 15118
rect 28988 14542 29022 15118
rect 29116 14542 29150 15118
rect 29228 14542 29262 15118
rect 29356 14542 29390 15118
rect 19930 14360 19968 14492
rect 20170 14360 20208 14492
rect 20410 14360 20448 14492
rect 20650 14360 20688 14492
rect 20890 14360 20928 14492
rect 21130 14360 21168 14492
rect 21370 14360 21408 14492
rect 21610 14360 21648 14492
rect 21850 14360 21888 14492
rect 22090 14360 22128 14492
rect 22330 14360 22368 14492
rect 22570 14360 22608 14492
rect 22810 14360 22848 14492
rect 23050 14360 23088 14492
rect 23290 14360 23328 14492
rect 23530 14360 23568 14492
rect 23770 14360 23808 14492
rect 24010 14360 24048 14492
rect 24250 14360 24288 14492
rect 24490 14360 24528 14492
rect 24730 14360 24768 14492
rect 24970 14360 25008 14492
rect 25210 14360 25248 14492
rect 25450 14360 25488 14492
rect 25690 14360 25728 14492
rect 25930 14360 25968 14492
rect 26170 14360 26208 14492
rect 26410 14360 26448 14492
rect 26650 14360 26688 14492
rect 26890 14360 26928 14492
rect 27130 14360 27168 14492
rect 27370 14360 27408 14492
rect 27610 14360 27648 14492
rect 27850 14360 27888 14492
rect 28090 14360 28128 14492
rect 28330 14360 28368 14492
rect 28570 14360 28608 14492
rect 28810 14360 28848 14492
rect 29050 14360 29088 14492
rect 29290 14360 29328 14492
rect 19868 13734 19902 14310
rect 19996 13734 20030 14310
rect 20108 13734 20142 14310
rect 20236 13734 20270 14310
rect 20348 13734 20382 14310
rect 20476 13734 20510 14310
rect 20588 13734 20622 14310
rect 20716 13734 20750 14310
rect 20828 13734 20862 14310
rect 20956 13734 20990 14310
rect 21068 13734 21102 14310
rect 21196 13734 21230 14310
rect 21308 13734 21342 14310
rect 21436 13734 21470 14310
rect 21548 13734 21582 14310
rect 21676 13734 21710 14310
rect 21788 13734 21822 14310
rect 21916 13734 21950 14310
rect 22028 13734 22062 14310
rect 22156 13734 22190 14310
rect 22268 13734 22302 14310
rect 22396 13734 22430 14310
rect 22508 13734 22542 14310
rect 22636 13734 22670 14310
rect 22748 13734 22782 14310
rect 22876 13734 22910 14310
rect 22988 13734 23022 14310
rect 23116 13734 23150 14310
rect 23228 13734 23262 14310
rect 23356 13734 23390 14310
rect 23468 13734 23502 14310
rect 23596 13734 23630 14310
rect 23708 13734 23742 14310
rect 23836 13734 23870 14310
rect 23948 13734 23982 14310
rect 24076 13734 24110 14310
rect 24188 13734 24222 14310
rect 24316 13734 24350 14310
rect 24428 13734 24462 14310
rect 24556 13734 24590 14310
rect 24668 13734 24702 14310
rect 24796 13734 24830 14310
rect 24908 13734 24942 14310
rect 25036 13734 25070 14310
rect 25148 13734 25182 14310
rect 25276 13734 25310 14310
rect 25388 13734 25422 14310
rect 25516 13734 25550 14310
rect 25628 13734 25662 14310
rect 25756 13734 25790 14310
rect 25868 13734 25902 14310
rect 25996 13734 26030 14310
rect 26108 13734 26142 14310
rect 26236 13734 26270 14310
rect 26348 13734 26382 14310
rect 26476 13734 26510 14310
rect 26588 13734 26622 14310
rect 26716 13734 26750 14310
rect 26828 13734 26862 14310
rect 26956 13734 26990 14310
rect 27068 13734 27102 14310
rect 27196 13734 27230 14310
rect 27308 13734 27342 14310
rect 27436 13734 27470 14310
rect 27548 13734 27582 14310
rect 27676 13734 27710 14310
rect 27788 13734 27822 14310
rect 27916 13734 27950 14310
rect 28028 13734 28062 14310
rect 28156 13734 28190 14310
rect 28268 13734 28302 14310
rect 28396 13734 28430 14310
rect 28508 13734 28542 14310
rect 28636 13734 28670 14310
rect 28748 13734 28782 14310
rect 28876 13734 28910 14310
rect 28988 13734 29022 14310
rect 29116 13734 29150 14310
rect 29228 13734 29262 14310
rect 29356 13734 29390 14310
rect 19930 13552 19968 13684
rect 20170 13552 20208 13684
rect 20410 13552 20448 13684
rect 20650 13552 20688 13684
rect 20890 13552 20928 13684
rect 21130 13552 21168 13684
rect 21370 13552 21408 13684
rect 21610 13552 21648 13684
rect 21850 13552 21888 13684
rect 22090 13552 22128 13684
rect 22330 13552 22368 13684
rect 22570 13552 22608 13684
rect 22810 13552 22848 13684
rect 23050 13552 23088 13684
rect 23290 13552 23328 13684
rect 23530 13552 23568 13684
rect 23770 13552 23808 13684
rect 24010 13552 24048 13684
rect 24250 13552 24288 13684
rect 24490 13552 24528 13684
rect 24730 13552 24768 13684
rect 24970 13552 25008 13684
rect 25210 13552 25248 13684
rect 25450 13552 25488 13684
rect 25690 13552 25728 13684
rect 25930 13552 25968 13684
rect 26170 13552 26208 13684
rect 26410 13552 26448 13684
rect 26650 13552 26688 13684
rect 26890 13552 26928 13684
rect 27130 13552 27168 13684
rect 27370 13552 27408 13684
rect 27610 13552 27648 13684
rect 27850 13552 27888 13684
rect 28090 13552 28128 13684
rect 28330 13552 28368 13684
rect 28570 13552 28608 13684
rect 28810 13552 28848 13684
rect 29050 13552 29088 13684
rect 29290 13552 29328 13684
rect 10626 11159 10994 11193
rect 11214 11159 11582 11193
rect 11802 11159 12170 11193
rect 12390 11159 12758 11193
rect 12978 11159 13346 11193
rect 13566 11159 13934 11193
rect 14154 11159 14522 11193
rect 14742 11159 15110 11193
rect 15330 11159 15698 11193
rect 15918 11159 16286 11193
rect 16506 11159 16874 11193
rect 17094 11159 17462 11193
rect 17682 11159 18050 11193
rect 18270 11159 18638 11193
rect 18858 11159 19226 11193
rect 19446 11159 19814 11193
rect 20034 11159 20402 11193
rect 20622 11159 20990 11193
rect 21210 11159 21578 11193
rect 21798 11159 22166 11193
rect 22386 11159 22754 11193
rect 22974 11159 23342 11193
rect 23562 11159 23930 11193
rect 24150 11159 24518 11193
rect 24738 11159 25106 11193
rect 25326 11159 25694 11193
rect 25914 11159 26282 11193
rect 26502 11159 26870 11193
rect 27090 11159 27458 11193
rect 27678 11159 28046 11193
rect 28266 11159 28634 11193
rect 28854 11159 29222 11193
rect 29442 11159 29810 11193
rect 30030 11159 30398 11193
rect 30618 11159 30986 11193
rect 31206 11159 31574 11193
rect 31794 11159 32162 11193
rect 32382 11159 32750 11193
rect 32970 11159 33338 11193
rect 33558 11159 33926 11193
rect 34146 11159 34514 11193
rect 34734 11159 35102 11193
rect 35322 11159 35690 11193
rect 35910 11159 36278 11193
rect 36498 11159 36866 11193
rect 37086 11159 37454 11193
rect 37674 11159 38042 11193
rect 38262 11159 38630 11193
rect 10564 10324 10598 11100
rect 11022 10324 11056 11100
rect 11152 10324 11186 11100
rect 11610 10324 11644 11100
rect 11740 10324 11774 11100
rect 12198 10324 12232 11100
rect 12328 10324 12362 11100
rect 12786 10324 12820 11100
rect 12916 10324 12950 11100
rect 13374 10324 13408 11100
rect 13504 10324 13538 11100
rect 13962 10324 13996 11100
rect 14092 10324 14126 11100
rect 14550 10324 14584 11100
rect 14680 10324 14714 11100
rect 15138 10324 15172 11100
rect 15268 10324 15302 11100
rect 15726 10324 15760 11100
rect 15856 10324 15890 11100
rect 16314 10324 16348 11100
rect 16444 10324 16478 11100
rect 16902 10324 16936 11100
rect 17032 10324 17066 11100
rect 17490 10324 17524 11100
rect 17620 10324 17654 11100
rect 18078 10324 18112 11100
rect 18208 10324 18242 11100
rect 18666 10324 18700 11100
rect 18796 10324 18830 11100
rect 19254 10324 19288 11100
rect 19384 10324 19418 11100
rect 19842 10324 19876 11100
rect 19972 10324 20006 11100
rect 20430 10324 20464 11100
rect 20560 10324 20594 11100
rect 21018 10324 21052 11100
rect 21148 10324 21182 11100
rect 21606 10324 21640 11100
rect 21736 10324 21770 11100
rect 22194 10324 22228 11100
rect 22324 10324 22358 11100
rect 22782 10324 22816 11100
rect 22912 10324 22946 11100
rect 23370 10324 23404 11100
rect 23500 10324 23534 11100
rect 23958 10324 23992 11100
rect 24088 10324 24122 11100
rect 24546 10324 24580 11100
rect 24676 10324 24710 11100
rect 25134 10324 25168 11100
rect 25264 10324 25298 11100
rect 25722 10324 25756 11100
rect 25852 10324 25886 11100
rect 26310 10324 26344 11100
rect 26440 10324 26474 11100
rect 26898 10324 26932 11100
rect 27028 10324 27062 11100
rect 27486 10324 27520 11100
rect 27616 10324 27650 11100
rect 28074 10324 28108 11100
rect 28204 10324 28238 11100
rect 28662 10324 28696 11100
rect 28792 10324 28826 11100
rect 29250 10324 29284 11100
rect 29380 10324 29414 11100
rect 29838 10324 29872 11100
rect 29968 10324 30002 11100
rect 30426 10324 30460 11100
rect 30556 10324 30590 11100
rect 31014 10324 31048 11100
rect 31144 10324 31178 11100
rect 31602 10324 31636 11100
rect 31732 10324 31766 11100
rect 32190 10324 32224 11100
rect 32320 10324 32354 11100
rect 32778 10324 32812 11100
rect 32908 10324 32942 11100
rect 33366 10324 33400 11100
rect 33496 10324 33530 11100
rect 33954 10324 33988 11100
rect 34084 10324 34118 11100
rect 34542 10324 34576 11100
rect 34672 10324 34706 11100
rect 35130 10324 35164 11100
rect 35260 10324 35294 11100
rect 35718 10324 35752 11100
rect 35848 10324 35882 11100
rect 36306 10324 36340 11100
rect 36436 10324 36470 11100
rect 36894 10324 36928 11100
rect 37024 10324 37058 11100
rect 37482 10324 37516 11100
rect 37612 10324 37646 11100
rect 38070 10324 38104 11100
rect 38200 10324 38234 11100
rect 38658 10324 38692 11100
rect 10626 10231 10994 10265
rect 11214 10231 11582 10265
rect 11802 10231 12170 10265
rect 12390 10231 12758 10265
rect 12978 10231 13346 10265
rect 13566 10231 13934 10265
rect 14154 10231 14522 10265
rect 14742 10231 15110 10265
rect 15330 10231 15698 10265
rect 15918 10231 16286 10265
rect 16506 10231 16874 10265
rect 17094 10231 17462 10265
rect 17682 10231 18050 10265
rect 18270 10231 18638 10265
rect 18858 10231 19226 10265
rect 19446 10231 19814 10265
rect 20034 10231 20402 10265
rect 20622 10231 20990 10265
rect 21210 10231 21578 10265
rect 21798 10231 22166 10265
rect 22386 10231 22754 10265
rect 22974 10231 23342 10265
rect 23562 10231 23930 10265
rect 24150 10231 24518 10265
rect 24738 10231 25106 10265
rect 25326 10231 25694 10265
rect 25914 10231 26282 10265
rect 26502 10231 26870 10265
rect 27090 10231 27458 10265
rect 27678 10231 28046 10265
rect 28266 10231 28634 10265
rect 28854 10231 29222 10265
rect 29442 10231 29810 10265
rect 30030 10231 30398 10265
rect 30618 10231 30986 10265
rect 31206 10231 31574 10265
rect 31794 10231 32162 10265
rect 32382 10231 32750 10265
rect 32970 10231 33338 10265
rect 33558 10231 33926 10265
rect 34146 10231 34514 10265
rect 34734 10231 35102 10265
rect 35322 10231 35690 10265
rect 35910 10231 36278 10265
rect 36498 10231 36866 10265
rect 37086 10231 37454 10265
rect 37674 10231 38042 10265
rect 38262 10231 38630 10265
rect 10626 10159 10994 10193
rect 11214 10159 11582 10193
rect 11802 10159 12170 10193
rect 12390 10159 12758 10193
rect 12978 10159 13346 10193
rect 13566 10159 13934 10193
rect 14154 10159 14522 10193
rect 14742 10159 15110 10193
rect 15330 10159 15698 10193
rect 15918 10159 16286 10193
rect 16506 10159 16874 10193
rect 17094 10159 17462 10193
rect 17682 10159 18050 10193
rect 18270 10159 18638 10193
rect 18858 10159 19226 10193
rect 19446 10159 19814 10193
rect 20034 10159 20402 10193
rect 20622 10159 20990 10193
rect 21210 10159 21578 10193
rect 21798 10159 22166 10193
rect 22386 10159 22754 10193
rect 22974 10159 23342 10193
rect 23562 10159 23930 10193
rect 24150 10159 24518 10193
rect 24738 10159 25106 10193
rect 25326 10159 25694 10193
rect 25914 10159 26282 10193
rect 26502 10159 26870 10193
rect 27090 10159 27458 10193
rect 27678 10159 28046 10193
rect 28266 10159 28634 10193
rect 28854 10159 29222 10193
rect 29442 10159 29810 10193
rect 30030 10159 30398 10193
rect 30618 10159 30986 10193
rect 31206 10159 31574 10193
rect 31794 10159 32162 10193
rect 32382 10159 32750 10193
rect 32970 10159 33338 10193
rect 33558 10159 33926 10193
rect 34146 10159 34514 10193
rect 34734 10159 35102 10193
rect 35322 10159 35690 10193
rect 35910 10159 36278 10193
rect 36498 10159 36866 10193
rect 37086 10159 37454 10193
rect 37674 10159 38042 10193
rect 38262 10159 38630 10193
rect 10564 9324 10598 10100
rect 11022 9324 11056 10100
rect 11152 9324 11186 10100
rect 11610 9324 11644 10100
rect 11740 9324 11774 10100
rect 12198 9324 12232 10100
rect 12328 9324 12362 10100
rect 12786 9324 12820 10100
rect 12916 9324 12950 10100
rect 13374 9324 13408 10100
rect 13504 9324 13538 10100
rect 13962 9324 13996 10100
rect 14092 9324 14126 10100
rect 14550 9324 14584 10100
rect 14680 9324 14714 10100
rect 15138 9324 15172 10100
rect 15268 9324 15302 10100
rect 15726 9324 15760 10100
rect 15856 9324 15890 10100
rect 16314 9324 16348 10100
rect 16444 9324 16478 10100
rect 16902 9324 16936 10100
rect 17032 9324 17066 10100
rect 17490 9324 17524 10100
rect 17620 9324 17654 10100
rect 18078 9324 18112 10100
rect 18208 9324 18242 10100
rect 18666 9324 18700 10100
rect 18796 9324 18830 10100
rect 19254 9324 19288 10100
rect 19384 9324 19418 10100
rect 19842 9324 19876 10100
rect 19972 9324 20006 10100
rect 20430 9324 20464 10100
rect 20560 9324 20594 10100
rect 21018 9324 21052 10100
rect 21148 9324 21182 10100
rect 21606 9324 21640 10100
rect 21736 9324 21770 10100
rect 22194 9324 22228 10100
rect 22324 9324 22358 10100
rect 22782 9324 22816 10100
rect 22912 9324 22946 10100
rect 23370 9324 23404 10100
rect 23500 9324 23534 10100
rect 23958 9324 23992 10100
rect 24088 9324 24122 10100
rect 24546 9324 24580 10100
rect 24676 9324 24710 10100
rect 25134 9324 25168 10100
rect 25264 9324 25298 10100
rect 25722 9324 25756 10100
rect 25852 9324 25886 10100
rect 26310 9324 26344 10100
rect 26440 9324 26474 10100
rect 26898 9324 26932 10100
rect 27028 9324 27062 10100
rect 27486 9324 27520 10100
rect 27616 9324 27650 10100
rect 28074 9324 28108 10100
rect 28204 9324 28238 10100
rect 28662 9324 28696 10100
rect 28792 9324 28826 10100
rect 29250 9324 29284 10100
rect 29380 9324 29414 10100
rect 29838 9324 29872 10100
rect 29968 9324 30002 10100
rect 30426 9324 30460 10100
rect 30556 9324 30590 10100
rect 31014 9324 31048 10100
rect 31144 9324 31178 10100
rect 31602 9324 31636 10100
rect 31732 9324 31766 10100
rect 32190 9324 32224 10100
rect 32320 9324 32354 10100
rect 32778 9324 32812 10100
rect 32908 9324 32942 10100
rect 33366 9324 33400 10100
rect 33496 9324 33530 10100
rect 33954 9324 33988 10100
rect 34084 9324 34118 10100
rect 34542 9324 34576 10100
rect 34672 9324 34706 10100
rect 35130 9324 35164 10100
rect 35260 9324 35294 10100
rect 35718 9324 35752 10100
rect 35848 9324 35882 10100
rect 36306 9324 36340 10100
rect 36436 9324 36470 10100
rect 36894 9324 36928 10100
rect 37024 9324 37058 10100
rect 37482 9324 37516 10100
rect 37612 9324 37646 10100
rect 38070 9324 38104 10100
rect 38200 9324 38234 10100
rect 38658 9324 38692 10100
rect 10626 9231 10994 9265
rect 11214 9231 11582 9265
rect 11802 9231 12170 9265
rect 12390 9231 12758 9265
rect 12978 9231 13346 9265
rect 13566 9231 13934 9265
rect 14154 9231 14522 9265
rect 14742 9231 15110 9265
rect 15330 9231 15698 9265
rect 15918 9231 16286 9265
rect 16506 9231 16874 9265
rect 17094 9231 17462 9265
rect 17682 9231 18050 9265
rect 18270 9231 18638 9265
rect 18858 9231 19226 9265
rect 19446 9231 19814 9265
rect 20034 9231 20402 9265
rect 20622 9231 20990 9265
rect 21210 9231 21578 9265
rect 21798 9231 22166 9265
rect 22386 9231 22754 9265
rect 22974 9231 23342 9265
rect 23562 9231 23930 9265
rect 24150 9231 24518 9265
rect 24738 9231 25106 9265
rect 25326 9231 25694 9265
rect 25914 9231 26282 9265
rect 26502 9231 26870 9265
rect 27090 9231 27458 9265
rect 27678 9231 28046 9265
rect 28266 9231 28634 9265
rect 28854 9231 29222 9265
rect 29442 9231 29810 9265
rect 30030 9231 30398 9265
rect 30618 9231 30986 9265
rect 31206 9231 31574 9265
rect 31794 9231 32162 9265
rect 32382 9231 32750 9265
rect 32970 9231 33338 9265
rect 33558 9231 33926 9265
rect 34146 9231 34514 9265
rect 34734 9231 35102 9265
rect 35322 9231 35690 9265
rect 35910 9231 36278 9265
rect 36498 9231 36866 9265
rect 37086 9231 37454 9265
rect 37674 9231 38042 9265
rect 38262 9231 38630 9265
rect 10626 9159 10994 9193
rect 11214 9159 11582 9193
rect 11802 9159 12170 9193
rect 12390 9159 12758 9193
rect 12978 9159 13346 9193
rect 13566 9159 13934 9193
rect 14154 9159 14522 9193
rect 14742 9159 15110 9193
rect 15330 9159 15698 9193
rect 15918 9159 16286 9193
rect 16506 9159 16874 9193
rect 17094 9159 17462 9193
rect 17682 9159 18050 9193
rect 18270 9159 18638 9193
rect 18858 9159 19226 9193
rect 19446 9159 19814 9193
rect 20034 9159 20402 9193
rect 20622 9159 20990 9193
rect 21210 9159 21578 9193
rect 21798 9159 22166 9193
rect 22386 9159 22754 9193
rect 22974 9159 23342 9193
rect 23562 9159 23930 9193
rect 24150 9159 24518 9193
rect 24738 9159 25106 9193
rect 25326 9159 25694 9193
rect 25914 9159 26282 9193
rect 26502 9159 26870 9193
rect 27090 9159 27458 9193
rect 27678 9159 28046 9193
rect 28266 9159 28634 9193
rect 28854 9159 29222 9193
rect 29442 9159 29810 9193
rect 30030 9159 30398 9193
rect 30618 9159 30986 9193
rect 31206 9159 31574 9193
rect 31794 9159 32162 9193
rect 32382 9159 32750 9193
rect 32970 9159 33338 9193
rect 33558 9159 33926 9193
rect 34146 9159 34514 9193
rect 34734 9159 35102 9193
rect 35322 9159 35690 9193
rect 35910 9159 36278 9193
rect 36498 9159 36866 9193
rect 37086 9159 37454 9193
rect 37674 9159 38042 9193
rect 38262 9159 38630 9193
rect 10564 8324 10598 9100
rect 11022 8324 11056 9100
rect 11152 8324 11186 9100
rect 11610 8324 11644 9100
rect 11740 8324 11774 9100
rect 12198 8324 12232 9100
rect 12328 8324 12362 9100
rect 12786 8324 12820 9100
rect 12916 8324 12950 9100
rect 13374 8324 13408 9100
rect 13504 8324 13538 9100
rect 13962 8324 13996 9100
rect 14092 8324 14126 9100
rect 14550 8324 14584 9100
rect 14680 8324 14714 9100
rect 15138 8324 15172 9100
rect 15268 8324 15302 9100
rect 15726 8324 15760 9100
rect 15856 8324 15890 9100
rect 16314 8324 16348 9100
rect 16444 8324 16478 9100
rect 16902 8324 16936 9100
rect 17032 8324 17066 9100
rect 17490 8324 17524 9100
rect 17620 8324 17654 9100
rect 18078 8324 18112 9100
rect 18208 8324 18242 9100
rect 18666 8324 18700 9100
rect 18796 8324 18830 9100
rect 19254 8324 19288 9100
rect 19384 8324 19418 9100
rect 19842 8324 19876 9100
rect 19972 8324 20006 9100
rect 20430 8324 20464 9100
rect 20560 8324 20594 9100
rect 21018 8324 21052 9100
rect 21148 8324 21182 9100
rect 21606 8324 21640 9100
rect 21736 8324 21770 9100
rect 22194 8324 22228 9100
rect 22324 8324 22358 9100
rect 22782 8324 22816 9100
rect 22912 8324 22946 9100
rect 23370 8324 23404 9100
rect 23500 8324 23534 9100
rect 23958 8324 23992 9100
rect 24088 8324 24122 9100
rect 24546 8324 24580 9100
rect 24676 8324 24710 9100
rect 25134 8324 25168 9100
rect 25264 8324 25298 9100
rect 25722 8324 25756 9100
rect 25852 8324 25886 9100
rect 26310 8324 26344 9100
rect 26440 8324 26474 9100
rect 26898 8324 26932 9100
rect 27028 8324 27062 9100
rect 27486 8324 27520 9100
rect 27616 8324 27650 9100
rect 28074 8324 28108 9100
rect 28204 8324 28238 9100
rect 28662 8324 28696 9100
rect 28792 8324 28826 9100
rect 29250 8324 29284 9100
rect 29380 8324 29414 9100
rect 29838 8324 29872 9100
rect 29968 8324 30002 9100
rect 30426 8324 30460 9100
rect 30556 8324 30590 9100
rect 31014 8324 31048 9100
rect 31144 8324 31178 9100
rect 31602 8324 31636 9100
rect 31732 8324 31766 9100
rect 32190 8324 32224 9100
rect 32320 8324 32354 9100
rect 32778 8324 32812 9100
rect 32908 8324 32942 9100
rect 33366 8324 33400 9100
rect 33496 8324 33530 9100
rect 33954 8324 33988 9100
rect 34084 8324 34118 9100
rect 34542 8324 34576 9100
rect 34672 8324 34706 9100
rect 35130 8324 35164 9100
rect 35260 8324 35294 9100
rect 35718 8324 35752 9100
rect 35848 8324 35882 9100
rect 36306 8324 36340 9100
rect 36436 8324 36470 9100
rect 36894 8324 36928 9100
rect 37024 8324 37058 9100
rect 37482 8324 37516 9100
rect 37612 8324 37646 9100
rect 38070 8324 38104 9100
rect 38200 8324 38234 9100
rect 38658 8324 38692 9100
rect 10626 8231 10994 8265
rect 11214 8231 11582 8265
rect 11802 8231 12170 8265
rect 12390 8231 12758 8265
rect 12978 8231 13346 8265
rect 13566 8231 13934 8265
rect 14154 8231 14522 8265
rect 14742 8231 15110 8265
rect 15330 8231 15698 8265
rect 15918 8231 16286 8265
rect 16506 8231 16874 8265
rect 17094 8231 17462 8265
rect 17682 8231 18050 8265
rect 18270 8231 18638 8265
rect 18858 8231 19226 8265
rect 19446 8231 19814 8265
rect 20034 8231 20402 8265
rect 20622 8231 20990 8265
rect 21210 8231 21578 8265
rect 21798 8231 22166 8265
rect 22386 8231 22754 8265
rect 22974 8231 23342 8265
rect 23562 8231 23930 8265
rect 24150 8231 24518 8265
rect 24738 8231 25106 8265
rect 25326 8231 25694 8265
rect 25914 8231 26282 8265
rect 26502 8231 26870 8265
rect 27090 8231 27458 8265
rect 27678 8231 28046 8265
rect 28266 8231 28634 8265
rect 28854 8231 29222 8265
rect 29442 8231 29810 8265
rect 30030 8231 30398 8265
rect 30618 8231 30986 8265
rect 31206 8231 31574 8265
rect 31794 8231 32162 8265
rect 32382 8231 32750 8265
rect 32970 8231 33338 8265
rect 33558 8231 33926 8265
rect 34146 8231 34514 8265
rect 34734 8231 35102 8265
rect 35322 8231 35690 8265
rect 35910 8231 36278 8265
rect 36498 8231 36866 8265
rect 37086 8231 37454 8265
rect 37674 8231 38042 8265
rect 38262 8231 38630 8265
rect 11010 7914 11198 7962
rect 12186 7914 12374 7962
rect 13362 7914 13550 7962
rect 14538 7914 14726 7962
rect 15714 7914 15902 7962
rect 16890 7914 17078 7962
rect 18066 7914 18254 7962
rect 19242 7914 19430 7962
rect 20418 7914 20606 7962
rect 21594 7914 21782 7962
rect 22770 7914 22958 7962
rect 23946 7914 24134 7962
rect 25122 7914 25310 7962
rect 26298 7914 26486 7962
rect 27474 7914 27662 7962
rect 28650 7914 28838 7962
rect 29826 7914 30014 7972
rect 31002 7914 31190 7962
rect 32178 7914 32366 7962
rect 33354 7914 33542 7962
rect 34516 7914 34728 7972
rect 35706 7914 35894 7962
rect 36882 7914 37070 7962
rect 38058 7914 38246 7962
rect 11010 7880 11198 7914
rect 12186 7880 12374 7914
rect 13362 7880 13550 7914
rect 14538 7880 14726 7914
rect 15714 7880 15902 7914
rect 16890 7880 17078 7914
rect 18066 7880 18254 7914
rect 19242 7880 19430 7914
rect 20418 7880 20606 7914
rect 21594 7880 21782 7914
rect 22770 7880 22958 7914
rect 23946 7880 24134 7914
rect 25122 7880 25310 7914
rect 26298 7880 26486 7914
rect 27474 7880 27662 7914
rect 28650 7880 28838 7914
rect 29826 7880 30014 7914
rect 31002 7880 31190 7914
rect 32178 7880 32366 7914
rect 33354 7880 33542 7914
rect 34516 7880 34728 7914
rect 35706 7880 35894 7914
rect 36882 7880 37070 7914
rect 38058 7880 38246 7914
rect 11010 7852 11198 7880
rect 12186 7852 12374 7880
rect 13362 7852 13550 7880
rect 14538 7852 14726 7880
rect 15714 7852 15902 7880
rect 16890 7852 17078 7880
rect 18066 7852 18254 7880
rect 19242 7852 19430 7880
rect 20418 7852 20606 7880
rect 21594 7852 21782 7880
rect 22770 7852 22958 7880
rect 23946 7852 24134 7880
rect 25122 7852 25310 7880
rect 26298 7852 26486 7880
rect 27474 7852 27662 7880
rect 28650 7852 28838 7880
rect 29826 7862 30014 7880
rect 31002 7852 31190 7880
rect 32178 7852 32366 7880
rect 33354 7852 33542 7880
rect 34516 7850 34728 7880
rect 35706 7852 35894 7880
rect 36882 7852 37070 7880
rect 38058 7852 38246 7880
rect 23678 6704 23716 6836
rect 23944 6704 23982 6836
rect 24210 6704 24248 6836
rect 24476 6704 24514 6836
rect 24742 6704 24780 6836
rect 25008 6704 25046 6836
rect 25274 6704 25312 6836
rect 25540 6704 25578 6836
rect 23616 5878 23650 6654
rect 23744 5878 23778 6654
rect 23882 5878 23916 6654
rect 24010 5878 24044 6654
rect 24148 5878 24182 6654
rect 24276 5878 24310 6654
rect 24414 5878 24448 6654
rect 24542 5878 24576 6654
rect 24680 5878 24714 6654
rect 24808 5878 24842 6654
rect 24946 5878 24980 6654
rect 25074 5878 25108 6654
rect 25212 5878 25246 6654
rect 25340 5878 25374 6654
rect 25478 5878 25512 6654
rect 25606 5878 25640 6654
rect 23678 5694 23716 5826
rect 23944 5694 23982 5826
rect 24210 5694 24248 5826
rect 24476 5694 24514 5826
rect 24742 5694 24780 5826
rect 25008 5694 25046 5826
rect 25274 5694 25312 5826
rect 25540 5694 25578 5826
rect 23616 4868 23650 5644
rect 23744 4868 23778 5644
rect 23882 4868 23916 5644
rect 24010 4868 24044 5644
rect 24148 4868 24182 5644
rect 24276 4868 24310 5644
rect 24414 4868 24448 5644
rect 24542 4868 24576 5644
rect 24680 4868 24714 5644
rect 24808 4868 24842 5644
rect 24946 4868 24980 5644
rect 25074 4868 25108 5644
rect 25212 4868 25246 5644
rect 25340 4868 25374 5644
rect 25478 4868 25512 5644
rect 25606 4868 25640 5644
rect 23678 4684 23716 4816
rect 23944 4684 23982 4816
rect 24210 4684 24248 4816
rect 24476 4684 24514 4816
rect 24742 4684 24780 4816
rect 25008 4684 25046 4816
rect 25274 4684 25312 4816
rect 25540 4684 25578 4816
rect 23616 3858 23650 4634
rect 23744 3858 23778 4634
rect 23882 3858 23916 4634
rect 24010 3858 24044 4634
rect 24148 3858 24182 4634
rect 24276 3858 24310 4634
rect 24414 3858 24448 4634
rect 24542 3858 24576 4634
rect 24680 3858 24714 4634
rect 24808 3858 24842 4634
rect 24946 3858 24980 4634
rect 25074 3858 25108 4634
rect 25212 3858 25246 4634
rect 25340 3858 25374 4634
rect 25478 3858 25512 4634
rect 25606 3858 25640 4634
rect 23678 3674 23716 3806
rect 23944 3674 23982 3806
rect 24210 3674 24248 3806
rect 24476 3674 24514 3806
rect 24742 3674 24780 3806
rect 25008 3674 25046 3806
rect 25274 3674 25312 3806
rect 25540 3674 25578 3806
rect 30797 4744 30835 5141
rect 30797 3753 30835 4150
rect 31086 4074 31226 4534
rect 24250 2512 24288 2638
rect 24490 2512 24528 2638
rect 24730 2512 24768 2638
rect 24970 2512 25008 2638
rect 24188 1886 24222 2462
rect 24316 1886 24350 2462
rect 24428 1886 24462 2462
rect 24556 1886 24590 2462
rect 24668 1886 24702 2462
rect 24796 1886 24830 2462
rect 24908 1886 24942 2462
rect 25036 1886 25070 2462
rect 24250 1704 24288 1836
rect 24490 1704 24528 1836
rect 24730 1704 24768 1836
rect 24970 1704 25008 1836
rect 24188 1078 24222 1654
rect 24316 1078 24350 1654
rect 24428 1078 24462 1654
rect 24556 1078 24590 1654
rect 24668 1078 24702 1654
rect 24796 1078 24830 1654
rect 24908 1078 24942 1654
rect 25036 1078 25070 1654
rect 24250 896 24288 1028
rect 24490 896 24528 1028
rect 24730 896 24768 1028
rect 24970 896 25008 1028
rect 23940 596 25292 644
rect 23940 562 24000 596
rect 24000 562 25210 596
rect 25210 562 25292 596
rect 23940 532 25292 562
<< metal1 >>
rect 20002 15644 20136 15650
rect 20002 15572 20014 15644
rect 20124 15572 20136 15644
rect 20002 15566 20136 15572
rect 20482 15644 20616 15650
rect 20482 15572 20494 15644
rect 20604 15572 20616 15644
rect 20482 15566 20616 15572
rect 20962 15644 21096 15650
rect 20962 15572 20974 15644
rect 21084 15572 21096 15644
rect 20962 15566 21096 15572
rect 21442 15644 21576 15650
rect 21442 15572 21454 15644
rect 21564 15572 21576 15644
rect 21442 15566 21576 15572
rect 21922 15644 22056 15650
rect 21922 15572 21934 15644
rect 22044 15572 22056 15644
rect 21922 15566 22056 15572
rect 22402 15644 22536 15650
rect 22402 15572 22414 15644
rect 22524 15572 22536 15644
rect 22402 15566 22536 15572
rect 22882 15644 23016 15650
rect 22882 15572 22894 15644
rect 23004 15572 23016 15644
rect 22882 15566 23016 15572
rect 23362 15644 23496 15650
rect 23362 15572 23374 15644
rect 23484 15572 23496 15644
rect 23362 15566 23496 15572
rect 23842 15644 23976 15650
rect 23842 15572 23854 15644
rect 23964 15572 23976 15644
rect 23842 15566 23976 15572
rect 24322 15644 24456 15650
rect 24322 15572 24334 15644
rect 24444 15572 24456 15644
rect 24322 15566 24456 15572
rect 24802 15644 24936 15650
rect 24802 15572 24814 15644
rect 24924 15572 24936 15644
rect 24802 15566 24936 15572
rect 25282 15644 25416 15650
rect 25282 15572 25294 15644
rect 25404 15572 25416 15644
rect 25282 15566 25416 15572
rect 25762 15644 25896 15650
rect 25762 15572 25774 15644
rect 25884 15572 25896 15644
rect 25762 15566 25896 15572
rect 26242 15644 26376 15650
rect 26242 15572 26254 15644
rect 26364 15572 26376 15644
rect 26242 15566 26376 15572
rect 26722 15644 26856 15650
rect 26722 15572 26734 15644
rect 26844 15572 26856 15644
rect 26722 15566 26856 15572
rect 27202 15644 27336 15650
rect 27202 15572 27214 15644
rect 27324 15572 27336 15644
rect 27202 15566 27336 15572
rect 27682 15644 27816 15650
rect 27682 15572 27694 15644
rect 27804 15572 27816 15644
rect 27682 15566 27816 15572
rect 28162 15644 28296 15650
rect 28162 15572 28174 15644
rect 28284 15572 28296 15644
rect 28162 15566 28296 15572
rect 28642 15644 28776 15650
rect 28642 15572 28654 15644
rect 28764 15572 28776 15644
rect 28642 15566 28776 15572
rect 29122 15644 29256 15650
rect 29122 15572 29134 15644
rect 29244 15572 29256 15644
rect 29122 15566 29256 15572
rect 19914 15300 19984 15306
rect 19904 15168 19914 15300
rect 19984 15168 19994 15300
rect 19914 15162 19984 15168
rect 20042 15130 20096 15566
rect 20154 15300 20224 15306
rect 20144 15168 20154 15300
rect 20224 15168 20234 15300
rect 20154 15162 20224 15168
rect 20282 15158 20336 15310
rect 20394 15300 20464 15306
rect 20384 15168 20394 15300
rect 20464 15168 20474 15300
rect 20394 15162 20464 15168
rect 20522 15130 20576 15566
rect 20634 15300 20704 15306
rect 20624 15168 20634 15300
rect 20704 15168 20714 15300
rect 20634 15162 20704 15168
rect 20762 15158 20816 15310
rect 20874 15300 20944 15306
rect 20864 15168 20874 15300
rect 20944 15168 20954 15300
rect 20874 15162 20944 15168
rect 21002 15130 21056 15566
rect 21114 15300 21184 15306
rect 21104 15168 21114 15300
rect 21184 15168 21194 15300
rect 21114 15162 21184 15168
rect 21242 15158 21296 15310
rect 21354 15300 21424 15306
rect 21344 15168 21354 15300
rect 21424 15168 21434 15300
rect 21354 15162 21424 15168
rect 21482 15130 21536 15566
rect 21594 15300 21664 15306
rect 21584 15168 21594 15300
rect 21664 15168 21674 15300
rect 21594 15162 21664 15168
rect 21722 15158 21776 15310
rect 21834 15300 21904 15306
rect 21824 15168 21834 15300
rect 21904 15168 21914 15300
rect 21834 15162 21904 15168
rect 21962 15130 22016 15566
rect 22074 15300 22144 15306
rect 22064 15168 22074 15300
rect 22144 15168 22154 15300
rect 22074 15162 22144 15168
rect 22202 15158 22256 15310
rect 22314 15300 22384 15306
rect 22304 15168 22314 15300
rect 22384 15168 22394 15300
rect 22314 15162 22384 15168
rect 22442 15130 22496 15566
rect 22554 15300 22624 15306
rect 22544 15168 22554 15300
rect 22624 15168 22634 15300
rect 22554 15162 22624 15168
rect 22682 15158 22736 15310
rect 22794 15300 22864 15306
rect 22784 15168 22794 15300
rect 22864 15168 22874 15300
rect 22794 15162 22864 15168
rect 22922 15130 22976 15566
rect 23034 15300 23104 15306
rect 23024 15168 23034 15300
rect 23104 15168 23114 15300
rect 23034 15162 23104 15168
rect 23162 15158 23216 15310
rect 23274 15300 23344 15306
rect 23264 15168 23274 15300
rect 23344 15168 23354 15300
rect 23274 15162 23344 15168
rect 23402 15130 23456 15566
rect 23514 15300 23584 15306
rect 23504 15168 23514 15300
rect 23584 15168 23594 15300
rect 23514 15162 23584 15168
rect 23642 15158 23696 15310
rect 23754 15300 23824 15306
rect 23744 15168 23754 15300
rect 23824 15168 23834 15300
rect 23754 15162 23824 15168
rect 23882 15130 23936 15566
rect 23994 15300 24064 15306
rect 23984 15168 23994 15300
rect 24064 15168 24074 15300
rect 23994 15162 24064 15168
rect 24122 15158 24176 15310
rect 24234 15300 24304 15306
rect 24224 15168 24234 15300
rect 24304 15168 24314 15300
rect 24234 15162 24304 15168
rect 24362 15130 24416 15566
rect 24474 15300 24544 15306
rect 24464 15168 24474 15300
rect 24544 15168 24554 15300
rect 24474 15162 24544 15168
rect 24602 15158 24656 15310
rect 24714 15300 24784 15306
rect 24704 15168 24714 15300
rect 24784 15168 24794 15300
rect 24714 15162 24784 15168
rect 24842 15130 24896 15566
rect 24954 15300 25024 15306
rect 24944 15168 24954 15300
rect 25024 15168 25034 15300
rect 24954 15162 25024 15168
rect 25082 15158 25136 15310
rect 25194 15300 25264 15306
rect 25184 15168 25194 15300
rect 25264 15168 25274 15300
rect 25194 15162 25264 15168
rect 25322 15130 25376 15566
rect 25434 15300 25504 15306
rect 25424 15168 25434 15300
rect 25504 15168 25514 15300
rect 25434 15162 25504 15168
rect 25562 15158 25616 15310
rect 25674 15300 25744 15306
rect 25664 15168 25674 15300
rect 25744 15168 25754 15300
rect 25674 15162 25744 15168
rect 25802 15130 25856 15566
rect 25914 15300 25984 15306
rect 25904 15168 25914 15300
rect 25984 15168 25994 15300
rect 25914 15162 25984 15168
rect 26042 15158 26096 15310
rect 26154 15300 26224 15306
rect 26144 15168 26154 15300
rect 26224 15168 26234 15300
rect 26154 15162 26224 15168
rect 26282 15130 26336 15566
rect 26394 15300 26464 15306
rect 26384 15168 26394 15300
rect 26464 15168 26474 15300
rect 26394 15162 26464 15168
rect 26522 15158 26576 15310
rect 26634 15300 26704 15306
rect 26624 15168 26634 15300
rect 26704 15168 26714 15300
rect 26634 15162 26704 15168
rect 26762 15130 26816 15566
rect 26874 15300 26944 15306
rect 26864 15168 26874 15300
rect 26944 15168 26954 15300
rect 26874 15162 26944 15168
rect 27002 15158 27056 15310
rect 27114 15300 27184 15306
rect 27104 15168 27114 15300
rect 27184 15168 27194 15300
rect 27114 15162 27184 15168
rect 27242 15130 27296 15566
rect 27354 15300 27424 15306
rect 27344 15168 27354 15300
rect 27424 15168 27434 15300
rect 27354 15162 27424 15168
rect 27482 15158 27536 15310
rect 27594 15300 27664 15306
rect 27584 15168 27594 15300
rect 27664 15168 27674 15300
rect 27594 15162 27664 15168
rect 27722 15130 27776 15566
rect 27834 15300 27904 15306
rect 27824 15168 27834 15300
rect 27904 15168 27914 15300
rect 27834 15162 27904 15168
rect 27962 15158 28016 15310
rect 28074 15300 28144 15306
rect 28064 15168 28074 15300
rect 28144 15168 28154 15300
rect 28074 15162 28144 15168
rect 28202 15130 28256 15566
rect 28314 15300 28384 15306
rect 28304 15168 28314 15300
rect 28384 15168 28394 15300
rect 28314 15162 28384 15168
rect 28442 15158 28496 15310
rect 28554 15300 28624 15306
rect 28544 15168 28554 15300
rect 28624 15168 28634 15300
rect 28554 15162 28624 15168
rect 28682 15130 28736 15566
rect 28794 15300 28864 15306
rect 28784 15168 28794 15300
rect 28864 15168 28874 15300
rect 28794 15162 28864 15168
rect 28922 15158 28976 15310
rect 29034 15300 29104 15306
rect 29024 15168 29034 15300
rect 29104 15168 29114 15300
rect 29034 15162 29104 15168
rect 29162 15130 29216 15566
rect 29274 15300 29344 15306
rect 29264 15168 29274 15300
rect 29344 15168 29354 15300
rect 29274 15162 29344 15168
rect 19790 15118 19908 15130
rect 19790 14542 19868 15118
rect 19902 14542 19908 15118
rect 19790 14530 19908 14542
rect 19990 15118 20148 15130
rect 19990 14542 19996 15118
rect 20030 14542 20108 15118
rect 20142 14542 20148 15118
rect 19990 14530 20148 14542
rect 20230 15118 20388 15130
rect 20230 14542 20236 15118
rect 20270 14542 20348 15118
rect 20382 14542 20388 15118
rect 20230 14530 20388 14542
rect 20470 15118 20628 15130
rect 20470 14542 20476 15118
rect 20510 14542 20588 15118
rect 20622 14542 20628 15118
rect 20470 14530 20628 14542
rect 20710 15118 20868 15130
rect 20710 14542 20716 15118
rect 20750 14542 20828 15118
rect 20862 14542 20868 15118
rect 20710 14530 20868 14542
rect 20950 15118 21108 15130
rect 20950 14542 20956 15118
rect 20990 14542 21068 15118
rect 21102 14542 21108 15118
rect 20950 14530 21108 14542
rect 21190 15118 21348 15130
rect 21190 14542 21196 15118
rect 21230 14542 21308 15118
rect 21342 14542 21348 15118
rect 21190 14530 21348 14542
rect 21430 15118 21588 15130
rect 21430 14542 21436 15118
rect 21470 14542 21548 15118
rect 21582 14542 21588 15118
rect 21430 14530 21588 14542
rect 21670 15118 21828 15130
rect 21670 14542 21676 15118
rect 21710 14542 21788 15118
rect 21822 14542 21828 15118
rect 21670 14530 21828 14542
rect 21910 15118 22068 15130
rect 21910 14542 21916 15118
rect 21950 14542 22028 15118
rect 22062 14542 22068 15118
rect 21910 14530 22068 14542
rect 22150 15118 22308 15130
rect 22150 14542 22156 15118
rect 22190 14542 22268 15118
rect 22302 14542 22308 15118
rect 22150 14530 22308 14542
rect 22390 15118 22548 15130
rect 22390 14542 22396 15118
rect 22430 14542 22508 15118
rect 22542 14542 22548 15118
rect 22390 14530 22548 14542
rect 22630 15118 22788 15130
rect 22630 14542 22636 15118
rect 22670 14542 22748 15118
rect 22782 14542 22788 15118
rect 22630 14530 22788 14542
rect 22870 15118 23028 15130
rect 22870 14542 22876 15118
rect 22910 14542 22988 15118
rect 23022 14542 23028 15118
rect 22870 14530 23028 14542
rect 23110 15118 23268 15130
rect 23110 14542 23116 15118
rect 23150 14542 23228 15118
rect 23262 14542 23268 15118
rect 23110 14530 23268 14542
rect 23350 15118 23508 15130
rect 23350 14542 23356 15118
rect 23390 14542 23468 15118
rect 23502 14542 23508 15118
rect 23350 14530 23508 14542
rect 23590 15118 23748 15130
rect 23590 14542 23596 15118
rect 23630 14542 23708 15118
rect 23742 14542 23748 15118
rect 23590 14530 23748 14542
rect 23830 15118 23988 15130
rect 23830 14542 23836 15118
rect 23870 14542 23948 15118
rect 23982 14542 23988 15118
rect 23830 14530 23988 14542
rect 24070 15118 24228 15130
rect 24070 14542 24076 15118
rect 24110 14542 24188 15118
rect 24222 14542 24228 15118
rect 24070 14530 24228 14542
rect 24310 15118 24468 15130
rect 24310 14542 24316 15118
rect 24350 14542 24428 15118
rect 24462 14542 24468 15118
rect 24310 14530 24468 14542
rect 24550 15118 24708 15130
rect 24550 14542 24556 15118
rect 24590 14542 24668 15118
rect 24702 14542 24708 15118
rect 24550 14530 24708 14542
rect 24790 15118 24948 15130
rect 24790 14542 24796 15118
rect 24830 14542 24908 15118
rect 24942 14542 24948 15118
rect 24790 14530 24948 14542
rect 25030 15118 25188 15130
rect 25030 14542 25036 15118
rect 25070 14542 25148 15118
rect 25182 14542 25188 15118
rect 25030 14530 25188 14542
rect 25270 15118 25428 15130
rect 25270 14542 25276 15118
rect 25310 14542 25388 15118
rect 25422 14542 25428 15118
rect 25270 14530 25428 14542
rect 25510 15118 25668 15130
rect 25510 14542 25516 15118
rect 25550 14542 25628 15118
rect 25662 14542 25668 15118
rect 25510 14530 25668 14542
rect 25750 15118 25908 15130
rect 25750 14542 25756 15118
rect 25790 14542 25868 15118
rect 25902 14542 25908 15118
rect 25750 14530 25908 14542
rect 25990 15118 26148 15130
rect 25990 14542 25996 15118
rect 26030 14542 26108 15118
rect 26142 14542 26148 15118
rect 25990 14530 26148 14542
rect 26230 15118 26388 15130
rect 26230 14542 26236 15118
rect 26270 14542 26348 15118
rect 26382 14542 26388 15118
rect 26230 14530 26388 14542
rect 26470 15118 26628 15130
rect 26470 14542 26476 15118
rect 26510 14542 26588 15118
rect 26622 14542 26628 15118
rect 26470 14530 26628 14542
rect 26710 15118 26868 15130
rect 26710 14542 26716 15118
rect 26750 14542 26828 15118
rect 26862 14542 26868 15118
rect 26710 14530 26868 14542
rect 26950 15118 27108 15130
rect 26950 14542 26956 15118
rect 26990 14542 27068 15118
rect 27102 14542 27108 15118
rect 26950 14530 27108 14542
rect 27190 15118 27348 15130
rect 27190 14542 27196 15118
rect 27230 14542 27308 15118
rect 27342 14542 27348 15118
rect 27190 14530 27348 14542
rect 27430 15118 27588 15130
rect 27430 14542 27436 15118
rect 27470 14542 27548 15118
rect 27582 14542 27588 15118
rect 27430 14530 27588 14542
rect 27670 15118 27828 15130
rect 27670 14542 27676 15118
rect 27710 14542 27788 15118
rect 27822 14542 27828 15118
rect 27670 14530 27828 14542
rect 27910 15118 28068 15130
rect 27910 14542 27916 15118
rect 27950 14542 28028 15118
rect 28062 14542 28068 15118
rect 27910 14530 28068 14542
rect 28150 15118 28308 15130
rect 28150 14542 28156 15118
rect 28190 14542 28268 15118
rect 28302 14542 28308 15118
rect 28150 14530 28308 14542
rect 28390 15118 28548 15130
rect 28390 14542 28396 15118
rect 28430 14542 28508 15118
rect 28542 14542 28548 15118
rect 28390 14530 28548 14542
rect 28630 15118 28788 15130
rect 28630 14542 28636 15118
rect 28670 14542 28748 15118
rect 28782 14542 28788 15118
rect 28630 14530 28788 14542
rect 28870 15118 29028 15130
rect 28870 14542 28876 15118
rect 28910 14542 28988 15118
rect 29022 14542 29028 15118
rect 28870 14530 29028 14542
rect 29110 15118 29268 15130
rect 29110 14542 29116 15118
rect 29150 14542 29228 15118
rect 29262 14542 29268 15118
rect 29110 14530 29268 14542
rect 29350 15118 29468 15130
rect 29350 14542 29356 15118
rect 29390 14542 29468 15118
rect 29350 14530 29468 14542
rect 19790 14322 19868 14530
rect 19914 14492 19984 14498
rect 19904 14360 19914 14492
rect 19984 14360 19994 14492
rect 19914 14354 19984 14360
rect 20036 14322 20102 14530
rect 20154 14492 20224 14498
rect 20144 14360 20154 14492
rect 20224 14360 20234 14492
rect 20154 14354 20224 14360
rect 20276 14322 20342 14530
rect 20394 14492 20464 14498
rect 20384 14360 20394 14492
rect 20464 14360 20474 14492
rect 20394 14354 20464 14360
rect 20516 14322 20582 14530
rect 20634 14492 20704 14498
rect 20624 14360 20634 14492
rect 20704 14360 20714 14492
rect 20634 14354 20704 14360
rect 20750 14322 20828 14530
rect 20874 14492 20944 14498
rect 20864 14360 20874 14492
rect 20944 14360 20954 14492
rect 20874 14354 20944 14360
rect 20996 14322 21062 14530
rect 21114 14492 21184 14498
rect 21104 14360 21114 14492
rect 21184 14360 21194 14492
rect 21114 14354 21184 14360
rect 21236 14322 21302 14530
rect 21354 14492 21424 14498
rect 21344 14360 21354 14492
rect 21424 14360 21434 14492
rect 21354 14354 21424 14360
rect 21476 14322 21542 14530
rect 21594 14492 21664 14498
rect 21584 14360 21594 14492
rect 21664 14360 21674 14492
rect 21594 14354 21664 14360
rect 21710 14322 21788 14530
rect 21834 14492 21904 14498
rect 21824 14360 21834 14492
rect 21904 14360 21914 14492
rect 21834 14354 21904 14360
rect 21956 14322 22022 14530
rect 22074 14492 22144 14498
rect 22064 14360 22074 14492
rect 22144 14360 22154 14492
rect 22074 14354 22144 14360
rect 22196 14322 22262 14530
rect 22314 14492 22384 14498
rect 22304 14360 22314 14492
rect 22384 14360 22394 14492
rect 22314 14354 22384 14360
rect 22436 14322 22502 14530
rect 22554 14492 22624 14498
rect 22544 14360 22554 14492
rect 22624 14360 22634 14492
rect 22554 14354 22624 14360
rect 22670 14322 22748 14530
rect 22794 14492 22864 14498
rect 22784 14360 22794 14492
rect 22864 14360 22874 14492
rect 22794 14354 22864 14360
rect 22916 14322 22982 14530
rect 23034 14492 23104 14498
rect 23024 14360 23034 14492
rect 23104 14360 23114 14492
rect 23034 14354 23104 14360
rect 23156 14322 23222 14530
rect 23274 14492 23344 14498
rect 23264 14360 23274 14492
rect 23344 14360 23354 14492
rect 23274 14354 23344 14360
rect 23396 14322 23462 14530
rect 23514 14492 23584 14498
rect 23504 14360 23514 14492
rect 23584 14360 23594 14492
rect 23514 14354 23584 14360
rect 23630 14322 23708 14530
rect 23754 14492 23824 14498
rect 23744 14360 23754 14492
rect 23824 14360 23834 14492
rect 23754 14354 23824 14360
rect 23876 14322 23942 14530
rect 23994 14492 24064 14498
rect 23984 14360 23994 14492
rect 24064 14360 24074 14492
rect 23994 14354 24064 14360
rect 24116 14322 24182 14530
rect 24234 14492 24304 14498
rect 24224 14360 24234 14492
rect 24304 14360 24314 14492
rect 24234 14354 24304 14360
rect 24356 14322 24422 14530
rect 24474 14492 24544 14498
rect 24464 14360 24474 14492
rect 24544 14360 24554 14492
rect 24474 14354 24544 14360
rect 24590 14322 24668 14530
rect 24714 14492 24784 14498
rect 24704 14360 24714 14492
rect 24784 14360 24794 14492
rect 24714 14354 24784 14360
rect 24836 14322 24902 14530
rect 24954 14492 25024 14498
rect 24944 14360 24954 14492
rect 25024 14360 25034 14492
rect 24954 14354 25024 14360
rect 25076 14322 25142 14530
rect 25194 14492 25264 14498
rect 25184 14360 25194 14492
rect 25264 14360 25274 14492
rect 25194 14354 25264 14360
rect 25316 14322 25382 14530
rect 25434 14492 25504 14498
rect 25424 14360 25434 14492
rect 25504 14360 25514 14492
rect 25434 14354 25504 14360
rect 25550 14322 25628 14530
rect 25674 14492 25744 14498
rect 25664 14360 25674 14492
rect 25744 14360 25754 14492
rect 25674 14354 25744 14360
rect 25796 14322 25862 14530
rect 25914 14492 25984 14498
rect 25904 14360 25914 14492
rect 25984 14360 25994 14492
rect 25914 14354 25984 14360
rect 26036 14322 26102 14530
rect 26154 14492 26224 14498
rect 26144 14360 26154 14492
rect 26224 14360 26234 14492
rect 26154 14354 26224 14360
rect 26276 14322 26342 14530
rect 26394 14492 26464 14498
rect 26384 14360 26394 14492
rect 26464 14360 26474 14492
rect 26394 14354 26464 14360
rect 26510 14322 26588 14530
rect 26634 14492 26704 14498
rect 26624 14360 26634 14492
rect 26704 14360 26714 14492
rect 26634 14354 26704 14360
rect 26756 14322 26822 14530
rect 26874 14492 26944 14498
rect 26864 14360 26874 14492
rect 26944 14360 26954 14492
rect 26874 14354 26944 14360
rect 26996 14322 27062 14530
rect 27114 14492 27184 14498
rect 27104 14360 27114 14492
rect 27184 14360 27194 14492
rect 27114 14354 27184 14360
rect 27236 14322 27302 14530
rect 27354 14492 27424 14498
rect 27344 14360 27354 14492
rect 27424 14360 27434 14492
rect 27354 14354 27424 14360
rect 27470 14322 27548 14530
rect 27594 14492 27664 14498
rect 27584 14360 27594 14492
rect 27664 14360 27674 14492
rect 27594 14354 27664 14360
rect 27716 14322 27782 14530
rect 27834 14492 27904 14498
rect 27824 14360 27834 14492
rect 27904 14360 27914 14492
rect 27834 14354 27904 14360
rect 27956 14322 28022 14530
rect 28074 14492 28144 14498
rect 28064 14360 28074 14492
rect 28144 14360 28154 14492
rect 28074 14354 28144 14360
rect 28196 14322 28262 14530
rect 28314 14492 28384 14498
rect 28304 14360 28314 14492
rect 28384 14360 28394 14492
rect 28314 14354 28384 14360
rect 28430 14322 28508 14530
rect 28554 14492 28624 14498
rect 28544 14360 28554 14492
rect 28624 14360 28634 14492
rect 28554 14354 28624 14360
rect 28676 14322 28742 14530
rect 28794 14492 28864 14498
rect 28784 14360 28794 14492
rect 28864 14360 28874 14492
rect 28794 14354 28864 14360
rect 28916 14322 28982 14530
rect 29034 14492 29104 14498
rect 29024 14360 29034 14492
rect 29104 14360 29114 14492
rect 29034 14354 29104 14360
rect 29156 14322 29222 14530
rect 29274 14492 29344 14498
rect 29264 14360 29274 14492
rect 29344 14360 29354 14492
rect 29274 14354 29344 14360
rect 29390 14322 29468 14530
rect 19790 14310 19908 14322
rect 19790 13734 19868 14310
rect 19902 13734 19908 14310
rect 19790 13722 19908 13734
rect 19990 14310 20148 14322
rect 19990 13734 19996 14310
rect 20030 13734 20108 14310
rect 20142 13734 20148 14310
rect 19990 13722 20148 13734
rect 20230 14310 20388 14322
rect 20230 13734 20236 14310
rect 20270 13734 20348 14310
rect 20382 13734 20388 14310
rect 20230 13722 20388 13734
rect 20470 14310 20628 14322
rect 20470 13734 20476 14310
rect 20510 13734 20588 14310
rect 20622 13734 20628 14310
rect 20470 13722 20628 13734
rect 20710 14310 20868 14322
rect 20710 13734 20716 14310
rect 20750 13734 20828 14310
rect 20862 13734 20868 14310
rect 20710 13722 20868 13734
rect 20950 14310 21108 14322
rect 20950 13734 20956 14310
rect 20990 13734 21068 14310
rect 21102 13734 21108 14310
rect 20950 13722 21108 13734
rect 21190 14310 21348 14322
rect 21190 13734 21196 14310
rect 21230 13734 21308 14310
rect 21342 13734 21348 14310
rect 21190 13722 21348 13734
rect 21430 14310 21588 14322
rect 21430 13734 21436 14310
rect 21470 13734 21548 14310
rect 21582 13734 21588 14310
rect 21430 13722 21588 13734
rect 21670 14310 21828 14322
rect 21670 13734 21676 14310
rect 21710 13734 21788 14310
rect 21822 13734 21828 14310
rect 21670 13722 21828 13734
rect 21910 14310 22068 14322
rect 21910 13734 21916 14310
rect 21950 13734 22028 14310
rect 22062 13734 22068 14310
rect 21910 13722 22068 13734
rect 22150 14310 22308 14322
rect 22150 13734 22156 14310
rect 22190 13734 22268 14310
rect 22302 13734 22308 14310
rect 22150 13722 22308 13734
rect 22390 14310 22548 14322
rect 22390 13734 22396 14310
rect 22430 13734 22508 14310
rect 22542 13734 22548 14310
rect 22390 13722 22548 13734
rect 22630 14310 22788 14322
rect 22630 13734 22636 14310
rect 22670 13734 22748 14310
rect 22782 13734 22788 14310
rect 22630 13722 22788 13734
rect 22870 14310 23028 14322
rect 22870 13734 22876 14310
rect 22910 13734 22988 14310
rect 23022 13734 23028 14310
rect 22870 13722 23028 13734
rect 23110 14310 23268 14322
rect 23110 13734 23116 14310
rect 23150 13734 23228 14310
rect 23262 13734 23268 14310
rect 23110 13722 23268 13734
rect 23350 14310 23508 14322
rect 23350 13734 23356 14310
rect 23390 13734 23468 14310
rect 23502 13734 23508 14310
rect 23350 13722 23508 13734
rect 23590 14310 23748 14322
rect 23590 13734 23596 14310
rect 23630 13734 23708 14310
rect 23742 13734 23748 14310
rect 23590 13722 23748 13734
rect 23830 14310 23988 14322
rect 23830 13734 23836 14310
rect 23870 13734 23948 14310
rect 23982 13734 23988 14310
rect 23830 13722 23988 13734
rect 24070 14310 24228 14322
rect 24070 13734 24076 14310
rect 24110 13734 24188 14310
rect 24222 13734 24228 14310
rect 24070 13722 24228 13734
rect 24310 14310 24468 14322
rect 24310 13734 24316 14310
rect 24350 13734 24428 14310
rect 24462 13734 24468 14310
rect 24310 13722 24468 13734
rect 24550 14310 24708 14322
rect 24550 13734 24556 14310
rect 24590 13734 24668 14310
rect 24702 13734 24708 14310
rect 24550 13722 24708 13734
rect 24790 14310 24948 14322
rect 24790 13734 24796 14310
rect 24830 13734 24908 14310
rect 24942 13734 24948 14310
rect 24790 13722 24948 13734
rect 25030 14310 25188 14322
rect 25030 13734 25036 14310
rect 25070 13734 25148 14310
rect 25182 13734 25188 14310
rect 25030 13722 25188 13734
rect 25270 14310 25428 14322
rect 25270 13734 25276 14310
rect 25310 13734 25388 14310
rect 25422 13734 25428 14310
rect 25270 13722 25428 13734
rect 25510 14310 25668 14322
rect 25510 13734 25516 14310
rect 25550 13734 25628 14310
rect 25662 13734 25668 14310
rect 25510 13722 25668 13734
rect 25750 14310 25908 14322
rect 25750 13734 25756 14310
rect 25790 13734 25868 14310
rect 25902 13734 25908 14310
rect 25750 13722 25908 13734
rect 25990 14310 26148 14322
rect 25990 13734 25996 14310
rect 26030 13734 26108 14310
rect 26142 13734 26148 14310
rect 25990 13722 26148 13734
rect 26230 14310 26388 14322
rect 26230 13734 26236 14310
rect 26270 13734 26348 14310
rect 26382 13734 26388 14310
rect 26230 13722 26388 13734
rect 26470 14310 26628 14322
rect 26470 13734 26476 14310
rect 26510 13734 26588 14310
rect 26622 13734 26628 14310
rect 26470 13722 26628 13734
rect 26710 14310 26868 14322
rect 26710 13734 26716 14310
rect 26750 13734 26828 14310
rect 26862 13734 26868 14310
rect 26710 13722 26868 13734
rect 26950 14310 27108 14322
rect 26950 13734 26956 14310
rect 26990 13734 27068 14310
rect 27102 13734 27108 14310
rect 26950 13722 27108 13734
rect 27190 14310 27348 14322
rect 27190 13734 27196 14310
rect 27230 13734 27308 14310
rect 27342 13734 27348 14310
rect 27190 13722 27348 13734
rect 27430 14310 27588 14322
rect 27430 13734 27436 14310
rect 27470 13734 27548 14310
rect 27582 13734 27588 14310
rect 27430 13722 27588 13734
rect 27670 14310 27828 14322
rect 27670 13734 27676 14310
rect 27710 13734 27788 14310
rect 27822 13734 27828 14310
rect 27670 13722 27828 13734
rect 27910 14310 28068 14322
rect 27910 13734 27916 14310
rect 27950 13734 28028 14310
rect 28062 13734 28068 14310
rect 27910 13722 28068 13734
rect 28150 14310 28308 14322
rect 28150 13734 28156 14310
rect 28190 13734 28268 14310
rect 28302 13734 28308 14310
rect 28150 13722 28308 13734
rect 28390 14310 28548 14322
rect 28390 13734 28396 14310
rect 28430 13734 28508 14310
rect 28542 13734 28548 14310
rect 28390 13722 28548 13734
rect 28630 14310 28788 14322
rect 28630 13734 28636 14310
rect 28670 13734 28748 14310
rect 28782 13734 28788 14310
rect 28630 13722 28788 13734
rect 28870 14310 29028 14322
rect 28870 13734 28876 14310
rect 28910 13734 28988 14310
rect 29022 13734 29028 14310
rect 28870 13722 29028 13734
rect 29110 14310 29268 14322
rect 29110 13734 29116 14310
rect 29150 13734 29228 14310
rect 29262 13734 29268 14310
rect 29110 13722 29268 13734
rect 29350 14310 29468 14322
rect 29350 13734 29356 14310
rect 29390 13734 29468 14310
rect 29350 13722 29468 13734
rect 19790 12856 19856 13722
rect 19914 13684 19984 13690
rect 20154 13684 20224 13690
rect 19904 13552 19914 13684
rect 19984 13552 19994 13684
rect 20144 13552 20154 13684
rect 20224 13552 20234 13684
rect 19914 13546 19984 13552
rect 20154 13546 20224 13552
rect 20282 12856 20336 13722
rect 20394 13684 20464 13690
rect 20634 13684 20704 13690
rect 20384 13552 20394 13684
rect 20464 13552 20474 13684
rect 20624 13552 20634 13684
rect 20704 13552 20714 13684
rect 20394 13546 20464 13552
rect 20634 13546 20704 13552
rect 20762 12856 20816 13722
rect 20874 13684 20944 13690
rect 21114 13684 21184 13690
rect 20864 13552 20874 13684
rect 20944 13552 20954 13684
rect 21104 13552 21114 13684
rect 21184 13552 21194 13684
rect 20874 13546 20944 13552
rect 21114 13546 21184 13552
rect 21242 12856 21296 13722
rect 21354 13684 21424 13690
rect 21594 13684 21664 13690
rect 21344 13552 21354 13684
rect 21424 13552 21434 13684
rect 21584 13552 21594 13684
rect 21664 13552 21674 13684
rect 21354 13546 21424 13552
rect 21594 13546 21664 13552
rect 21722 12856 21776 13722
rect 21834 13684 21904 13690
rect 22074 13684 22144 13690
rect 21824 13552 21834 13684
rect 21904 13552 21914 13684
rect 22064 13552 22074 13684
rect 22144 13552 22154 13684
rect 21834 13546 21904 13552
rect 22074 13546 22144 13552
rect 22202 12856 22256 13722
rect 22314 13684 22384 13690
rect 22554 13684 22624 13690
rect 22304 13552 22314 13684
rect 22384 13552 22394 13684
rect 22544 13552 22554 13684
rect 22624 13552 22634 13684
rect 22314 13546 22384 13552
rect 22554 13546 22624 13552
rect 22682 12856 22736 13722
rect 22794 13684 22864 13690
rect 23034 13684 23104 13690
rect 22784 13552 22794 13684
rect 22864 13552 22874 13684
rect 23024 13552 23034 13684
rect 23104 13552 23114 13684
rect 22794 13546 22864 13552
rect 23034 13546 23104 13552
rect 23162 12856 23216 13722
rect 23274 13684 23344 13690
rect 23514 13684 23584 13690
rect 23264 13552 23274 13684
rect 23344 13552 23354 13684
rect 23504 13552 23514 13684
rect 23584 13552 23594 13684
rect 23274 13546 23344 13552
rect 23514 13546 23584 13552
rect 23642 12856 23696 13722
rect 23754 13684 23824 13690
rect 23994 13684 24064 13690
rect 23744 13552 23754 13684
rect 23824 13552 23834 13684
rect 23984 13552 23994 13684
rect 24064 13552 24074 13684
rect 23754 13546 23824 13552
rect 23994 13546 24064 13552
rect 24122 12856 24176 13722
rect 24234 13684 24304 13690
rect 24474 13684 24544 13690
rect 24224 13552 24234 13684
rect 24304 13552 24314 13684
rect 24464 13552 24474 13684
rect 24544 13552 24554 13684
rect 24234 13546 24304 13552
rect 24474 13546 24544 13552
rect 24602 12856 24656 13722
rect 24714 13684 24784 13690
rect 24954 13684 25024 13690
rect 24704 13552 24714 13684
rect 24784 13552 24794 13684
rect 24944 13552 24954 13684
rect 25024 13552 25034 13684
rect 24714 13546 24784 13552
rect 24954 13546 25024 13552
rect 25082 12856 25136 13722
rect 25194 13684 25264 13690
rect 25434 13684 25504 13690
rect 25184 13552 25194 13684
rect 25264 13552 25274 13684
rect 25424 13552 25434 13684
rect 25504 13552 25514 13684
rect 25194 13546 25264 13552
rect 25434 13546 25504 13552
rect 25562 12856 25616 13722
rect 25674 13684 25744 13690
rect 25914 13684 25984 13690
rect 25664 13552 25674 13684
rect 25744 13552 25754 13684
rect 25904 13552 25914 13684
rect 25984 13552 25994 13684
rect 25674 13546 25744 13552
rect 25914 13546 25984 13552
rect 26042 12856 26096 13722
rect 26154 13684 26224 13690
rect 26394 13684 26464 13690
rect 26144 13552 26154 13684
rect 26224 13552 26234 13684
rect 26384 13552 26394 13684
rect 26464 13552 26474 13684
rect 26154 13546 26224 13552
rect 26394 13546 26464 13552
rect 26522 12856 26576 13722
rect 26634 13684 26704 13690
rect 26874 13684 26944 13690
rect 26624 13552 26634 13684
rect 26704 13552 26714 13684
rect 26864 13552 26874 13684
rect 26944 13552 26954 13684
rect 26634 13546 26704 13552
rect 26874 13546 26944 13552
rect 27002 12856 27056 13722
rect 27114 13684 27184 13690
rect 27354 13684 27424 13690
rect 27104 13552 27114 13684
rect 27184 13552 27194 13684
rect 27344 13552 27354 13684
rect 27424 13552 27434 13684
rect 27114 13546 27184 13552
rect 27354 13546 27424 13552
rect 27482 12856 27536 13722
rect 27594 13684 27664 13690
rect 27834 13684 27904 13690
rect 27584 13552 27594 13684
rect 27664 13552 27674 13684
rect 27824 13552 27834 13684
rect 27904 13552 27914 13684
rect 27594 13546 27664 13552
rect 27834 13546 27904 13552
rect 27962 12856 28016 13722
rect 28074 13684 28144 13690
rect 28314 13684 28384 13690
rect 28064 13552 28074 13684
rect 28144 13552 28154 13684
rect 28304 13552 28314 13684
rect 28384 13552 28394 13684
rect 28074 13546 28144 13552
rect 28314 13546 28384 13552
rect 28442 12856 28496 13722
rect 28554 13684 28624 13690
rect 28794 13684 28864 13690
rect 28544 13552 28554 13684
rect 28624 13552 28634 13684
rect 28784 13552 28794 13684
rect 28864 13552 28874 13684
rect 28554 13546 28624 13552
rect 28794 13546 28864 13552
rect 28922 12856 28976 13722
rect 29034 13684 29104 13690
rect 29274 13684 29344 13690
rect 29024 13552 29034 13684
rect 29104 13552 29114 13684
rect 29264 13552 29274 13684
rect 29344 13552 29354 13684
rect 29034 13546 29104 13552
rect 29274 13546 29344 13552
rect 29402 12856 29468 13722
rect 10474 12658 38782 12856
rect 10474 12216 33856 12658
rect 34756 12216 38782 12658
rect 10474 12050 38782 12216
rect 10474 11112 10552 12050
rect 10614 11193 11006 11199
rect 10614 11159 10626 11193
rect 10994 11159 11006 11193
rect 10614 11153 11006 11159
rect 11202 11193 11594 11199
rect 11202 11159 11214 11193
rect 11582 11159 11594 11193
rect 11202 11153 11594 11159
rect 11656 11112 11728 12050
rect 11790 11193 12182 11199
rect 11790 11159 11802 11193
rect 12170 11159 12182 11193
rect 11790 11153 12182 11159
rect 12378 11193 12770 11199
rect 12378 11159 12390 11193
rect 12758 11159 12770 11193
rect 12378 11153 12770 11159
rect 12832 11112 12904 12050
rect 12966 11193 13358 11199
rect 12966 11159 12978 11193
rect 13346 11159 13358 11193
rect 12966 11153 13358 11159
rect 13554 11193 13946 11199
rect 13554 11159 13566 11193
rect 13934 11159 13946 11193
rect 13554 11153 13946 11159
rect 14008 11112 14080 12050
rect 14142 11193 14534 11199
rect 14142 11159 14154 11193
rect 14522 11159 14534 11193
rect 14142 11153 14534 11159
rect 14730 11193 15122 11199
rect 14730 11159 14742 11193
rect 15110 11159 15122 11193
rect 14730 11153 15122 11159
rect 15184 11112 15256 12050
rect 15318 11193 15710 11199
rect 15318 11159 15330 11193
rect 15698 11159 15710 11193
rect 15318 11153 15710 11159
rect 15906 11193 16298 11199
rect 15906 11159 15918 11193
rect 16286 11159 16298 11193
rect 15906 11153 16298 11159
rect 16360 11112 16432 12050
rect 16494 11193 16886 11199
rect 16494 11159 16506 11193
rect 16874 11159 16886 11193
rect 16494 11153 16886 11159
rect 17082 11193 17474 11199
rect 17082 11159 17094 11193
rect 17462 11159 17474 11193
rect 17082 11153 17474 11159
rect 17536 11112 17608 12050
rect 17670 11193 18062 11199
rect 17670 11159 17682 11193
rect 18050 11159 18062 11193
rect 17670 11153 18062 11159
rect 18258 11193 18650 11199
rect 18258 11159 18270 11193
rect 18638 11159 18650 11193
rect 18258 11153 18650 11159
rect 18712 11112 18784 12050
rect 18846 11193 19238 11199
rect 18846 11159 18858 11193
rect 19226 11159 19238 11193
rect 18846 11153 19238 11159
rect 19434 11193 19826 11199
rect 19434 11159 19446 11193
rect 19814 11159 19826 11193
rect 19434 11153 19826 11159
rect 19888 11112 19960 12050
rect 20022 11193 20414 11199
rect 20022 11159 20034 11193
rect 20402 11159 20414 11193
rect 20022 11153 20414 11159
rect 20610 11193 21002 11199
rect 20610 11159 20622 11193
rect 20990 11159 21002 11193
rect 20610 11153 21002 11159
rect 21064 11112 21136 12050
rect 21198 11193 21590 11199
rect 21198 11159 21210 11193
rect 21578 11159 21590 11193
rect 21198 11153 21590 11159
rect 21786 11193 22178 11199
rect 21786 11159 21798 11193
rect 22166 11159 22178 11193
rect 21786 11153 22178 11159
rect 22212 11112 22284 12050
rect 22374 11193 22766 11199
rect 22374 11159 22386 11193
rect 22754 11159 22766 11193
rect 22374 11153 22766 11159
rect 22962 11193 23354 11199
rect 22962 11159 22974 11193
rect 23342 11159 23354 11193
rect 22962 11153 23354 11159
rect 23550 11193 23942 11199
rect 23550 11159 23562 11193
rect 23930 11159 23942 11193
rect 23550 11153 23942 11159
rect 24138 11193 24530 11199
rect 24138 11159 24150 11193
rect 24518 11159 24530 11193
rect 24138 11153 24530 11159
rect 24726 11193 25118 11199
rect 24726 11159 24738 11193
rect 25106 11159 25118 11193
rect 24726 11153 25118 11159
rect 25314 11193 25706 11199
rect 25314 11159 25326 11193
rect 25694 11159 25706 11193
rect 25314 11153 25706 11159
rect 25902 11193 26294 11199
rect 25902 11159 25914 11193
rect 26282 11159 26294 11193
rect 25902 11153 26294 11159
rect 26490 11193 26882 11199
rect 26490 11159 26502 11193
rect 26870 11159 26882 11193
rect 26490 11153 26882 11159
rect 26972 11112 27044 12050
rect 27078 11193 27470 11199
rect 27078 11159 27090 11193
rect 27458 11159 27470 11193
rect 27078 11153 27470 11159
rect 27666 11193 28058 11199
rect 27666 11159 27678 11193
rect 28046 11159 28058 11193
rect 27666 11153 28058 11159
rect 28120 11112 28192 12050
rect 28254 11193 28646 11199
rect 28254 11159 28266 11193
rect 28634 11159 28646 11193
rect 28254 11153 28646 11159
rect 28842 11193 29234 11199
rect 28842 11159 28854 11193
rect 29222 11159 29234 11193
rect 28842 11153 29234 11159
rect 29296 11112 29368 12050
rect 29430 11193 29822 11199
rect 29430 11159 29442 11193
rect 29810 11159 29822 11193
rect 29430 11153 29822 11159
rect 30018 11193 30410 11199
rect 30018 11159 30030 11193
rect 30398 11159 30410 11193
rect 30018 11153 30410 11159
rect 30472 11112 30544 12050
rect 30606 11193 30998 11199
rect 30606 11159 30618 11193
rect 30986 11159 30998 11193
rect 30606 11153 30998 11159
rect 31194 11193 31586 11199
rect 31194 11159 31206 11193
rect 31574 11159 31586 11193
rect 31194 11153 31586 11159
rect 31648 11112 31720 12050
rect 31782 11193 32174 11199
rect 31782 11159 31794 11193
rect 32162 11159 32174 11193
rect 31782 11153 32174 11159
rect 32370 11193 32762 11199
rect 32370 11159 32382 11193
rect 32750 11159 32762 11193
rect 32370 11153 32762 11159
rect 32824 11112 32896 12050
rect 32958 11193 33350 11199
rect 32958 11159 32970 11193
rect 33338 11159 33350 11193
rect 32958 11153 33350 11159
rect 33546 11193 33938 11199
rect 33546 11159 33558 11193
rect 33926 11159 33938 11193
rect 33546 11153 33938 11159
rect 34000 11112 34072 12050
rect 34134 11193 34526 11199
rect 34134 11159 34146 11193
rect 34514 11159 34526 11193
rect 34134 11153 34526 11159
rect 34722 11193 35114 11199
rect 34722 11159 34734 11193
rect 35102 11159 35114 11193
rect 34722 11153 35114 11159
rect 35176 11112 35248 12050
rect 35310 11193 35702 11199
rect 35310 11159 35322 11193
rect 35690 11159 35702 11193
rect 35310 11153 35702 11159
rect 35898 11193 36290 11199
rect 35898 11159 35910 11193
rect 36278 11159 36290 11193
rect 35898 11153 36290 11159
rect 36352 11112 36424 12050
rect 36486 11193 36878 11199
rect 36486 11159 36498 11193
rect 36866 11159 36878 11193
rect 36486 11153 36878 11159
rect 37074 11193 37466 11199
rect 37074 11159 37086 11193
rect 37454 11159 37466 11193
rect 37074 11153 37466 11159
rect 37528 11112 37600 12050
rect 37662 11193 38054 11199
rect 37662 11159 37674 11193
rect 38042 11159 38054 11193
rect 37662 11153 38054 11159
rect 38250 11193 38642 11199
rect 38250 11159 38262 11193
rect 38630 11159 38642 11193
rect 38250 11153 38642 11159
rect 38704 11112 38782 12050
rect 10474 11100 10604 11112
rect 10474 10324 10564 11100
rect 10598 10324 10604 11100
rect 10474 10312 10604 10324
rect 11016 11100 11192 11112
rect 11016 10324 11022 11100
rect 11056 10324 11152 11100
rect 11186 10324 11192 11100
rect 11016 10312 11192 10324
rect 11604 11100 11780 11112
rect 11604 10324 11610 11100
rect 11644 10324 11740 11100
rect 11774 10324 11780 11100
rect 11604 10312 11780 10324
rect 12192 11100 12368 11112
rect 12192 10324 12198 11100
rect 12232 10324 12328 11100
rect 12362 10324 12368 11100
rect 12192 10312 12368 10324
rect 12780 11100 12956 11112
rect 12780 10324 12786 11100
rect 12820 10324 12916 11100
rect 12950 10324 12956 11100
rect 12780 10312 12956 10324
rect 13368 11100 13544 11112
rect 13368 10324 13374 11100
rect 13408 10324 13504 11100
rect 13538 10324 13544 11100
rect 13368 10312 13544 10324
rect 13956 11100 14132 11112
rect 13956 10324 13962 11100
rect 13996 10324 14092 11100
rect 14126 10324 14132 11100
rect 13956 10312 14132 10324
rect 14544 11100 14720 11112
rect 14544 10324 14550 11100
rect 14584 10324 14680 11100
rect 14714 10324 14720 11100
rect 14544 10312 14720 10324
rect 15132 11100 15308 11112
rect 15132 10324 15138 11100
rect 15172 10324 15268 11100
rect 15302 10324 15308 11100
rect 15132 10312 15308 10324
rect 15720 11100 15896 11112
rect 15720 10324 15726 11100
rect 15760 10324 15856 11100
rect 15890 10324 15896 11100
rect 15720 10312 15896 10324
rect 16308 11100 16484 11112
rect 16308 10324 16314 11100
rect 16348 10324 16444 11100
rect 16478 10324 16484 11100
rect 16308 10312 16484 10324
rect 16896 11100 17072 11112
rect 16896 10324 16902 11100
rect 16936 10324 17032 11100
rect 17066 10324 17072 11100
rect 16896 10312 17072 10324
rect 17484 11100 17660 11112
rect 17484 10324 17490 11100
rect 17524 10324 17620 11100
rect 17654 10324 17660 11100
rect 17484 10312 17660 10324
rect 18072 11100 18248 11112
rect 18072 10324 18078 11100
rect 18112 10324 18208 11100
rect 18242 10324 18248 11100
rect 18072 10312 18248 10324
rect 18660 11100 18836 11112
rect 18660 10324 18666 11100
rect 18700 10324 18796 11100
rect 18830 10324 18836 11100
rect 18660 10312 18836 10324
rect 19248 11100 19424 11112
rect 19248 10324 19254 11100
rect 19288 10324 19384 11100
rect 19418 10324 19424 11100
rect 19248 10312 19424 10324
rect 19836 11100 20012 11112
rect 19836 10324 19842 11100
rect 19876 10324 19972 11100
rect 20006 10324 20012 11100
rect 19836 10312 20012 10324
rect 20424 11100 20600 11112
rect 20424 10324 20430 11100
rect 20464 10324 20560 11100
rect 20594 10324 20600 11100
rect 20424 10312 20600 10324
rect 21012 11100 21188 11112
rect 21012 10324 21018 11100
rect 21052 10324 21148 11100
rect 21182 10324 21188 11100
rect 21012 10312 21188 10324
rect 21600 11100 21776 11112
rect 21600 10324 21606 11100
rect 21640 10324 21736 11100
rect 21770 10324 21776 11100
rect 21600 10312 21776 10324
rect 22188 11100 22284 11112
rect 22188 10324 22194 11100
rect 22228 10376 22284 11100
rect 22318 11100 22364 11112
rect 22228 10324 22286 10376
rect 22188 10312 22286 10324
rect 22318 10324 22324 11100
rect 22358 10324 22364 11100
rect 22318 10312 22364 10324
rect 22776 11100 22952 11112
rect 22776 10324 22782 11100
rect 22816 10324 22912 11100
rect 22946 10324 22952 11100
rect 22776 10312 22952 10324
rect 23364 11100 23540 11112
rect 23364 10324 23370 11100
rect 23404 10324 23500 11100
rect 23534 10324 23540 11100
rect 23364 10312 23540 10324
rect 23952 11100 24128 11112
rect 23952 10324 23958 11100
rect 23992 10324 24088 11100
rect 24122 10324 24128 11100
rect 23952 10312 24128 10324
rect 24540 11100 24586 11112
rect 24540 10324 24546 11100
rect 24580 10324 24586 11100
rect 24540 10312 24586 10324
rect 24670 11100 24716 11112
rect 24670 10324 24676 11100
rect 24710 10324 24716 11100
rect 24670 10312 24716 10324
rect 25128 11100 25304 11112
rect 25128 10324 25134 11100
rect 25168 10324 25264 11100
rect 25298 10324 25304 11100
rect 25128 10312 25304 10324
rect 25716 11100 25892 11112
rect 25716 10324 25722 11100
rect 25756 10324 25852 11100
rect 25886 10324 25892 11100
rect 25716 10312 25892 10324
rect 26304 11100 26480 11112
rect 26304 10324 26310 11100
rect 26344 10324 26440 11100
rect 26474 10324 26480 11100
rect 26304 10312 26480 10324
rect 26892 11100 26938 11112
rect 26892 10324 26898 11100
rect 26932 10324 26938 11100
rect 26892 10312 26938 10324
rect 26972 11100 27068 11112
rect 26972 10324 27028 11100
rect 27062 10324 27068 11100
rect 26972 10312 27068 10324
rect 27480 11100 27656 11112
rect 27480 10324 27486 11100
rect 27520 10324 27616 11100
rect 27650 10324 27656 11100
rect 27480 10312 27656 10324
rect 28068 11100 28244 11112
rect 28068 10324 28074 11100
rect 28108 10324 28204 11100
rect 28238 10324 28244 11100
rect 28068 10312 28244 10324
rect 28656 11100 28832 11112
rect 28656 10324 28662 11100
rect 28696 10324 28792 11100
rect 28826 10324 28832 11100
rect 28656 10312 28832 10324
rect 29244 11100 29420 11112
rect 29244 10324 29250 11100
rect 29284 10324 29380 11100
rect 29414 10324 29420 11100
rect 29244 10312 29420 10324
rect 29832 11100 30008 11112
rect 29832 10324 29838 11100
rect 29872 10324 29968 11100
rect 30002 10324 30008 11100
rect 29832 10312 30008 10324
rect 30420 11100 30596 11112
rect 30420 10324 30426 11100
rect 30460 10324 30556 11100
rect 30590 10324 30596 11100
rect 30420 10312 30596 10324
rect 31008 11100 31184 11112
rect 31008 10324 31014 11100
rect 31048 10324 31144 11100
rect 31178 10324 31184 11100
rect 31008 10312 31184 10324
rect 31596 11100 31772 11112
rect 31596 10324 31602 11100
rect 31636 10324 31732 11100
rect 31766 10324 31772 11100
rect 31596 10312 31772 10324
rect 32184 11100 32360 11112
rect 32184 10324 32190 11100
rect 32224 10324 32320 11100
rect 32354 10324 32360 11100
rect 32184 10312 32360 10324
rect 32772 11100 32948 11112
rect 32772 10324 32778 11100
rect 32812 10324 32908 11100
rect 32942 10324 32948 11100
rect 32772 10312 32948 10324
rect 33360 11100 33536 11112
rect 33360 10324 33366 11100
rect 33400 10324 33496 11100
rect 33530 10324 33536 11100
rect 33360 10312 33536 10324
rect 33948 11100 34124 11112
rect 33948 10324 33954 11100
rect 33988 10324 34084 11100
rect 34118 10324 34124 11100
rect 33948 10312 34124 10324
rect 34536 11100 34712 11112
rect 34536 10324 34542 11100
rect 34576 10324 34672 11100
rect 34706 10324 34712 11100
rect 34536 10312 34712 10324
rect 35124 11100 35300 11112
rect 35124 10324 35130 11100
rect 35164 10324 35260 11100
rect 35294 10324 35300 11100
rect 35124 10312 35300 10324
rect 35712 11100 35888 11112
rect 35712 10324 35718 11100
rect 35752 10324 35848 11100
rect 35882 10324 35888 11100
rect 35712 10312 35888 10324
rect 36300 11100 36476 11112
rect 36300 10324 36306 11100
rect 36340 10324 36436 11100
rect 36470 10324 36476 11100
rect 36300 10312 36476 10324
rect 36888 11100 37064 11112
rect 36888 10324 36894 11100
rect 36928 10324 37024 11100
rect 37058 10324 37064 11100
rect 36888 10312 37064 10324
rect 37476 11100 37652 11112
rect 37476 10324 37482 11100
rect 37516 10324 37612 11100
rect 37646 10324 37652 11100
rect 37476 10312 37652 10324
rect 38064 11100 38240 11112
rect 38064 10324 38070 11100
rect 38104 10324 38200 11100
rect 38234 10324 38240 11100
rect 38064 10312 38240 10324
rect 38652 11100 38782 11112
rect 38652 10324 38658 11100
rect 38692 10324 38782 11100
rect 38652 10312 38782 10324
rect 10474 10112 10558 10312
rect 10614 10265 11006 10271
rect 10614 10231 10626 10265
rect 10994 10231 11006 10265
rect 10614 10193 11006 10231
rect 10614 10159 10626 10193
rect 10994 10159 11006 10193
rect 10614 10153 11006 10159
rect 11062 10112 11146 10312
rect 11202 10265 11594 10271
rect 11202 10231 11214 10265
rect 11582 10231 11594 10265
rect 11202 10193 11594 10231
rect 11202 10159 11214 10193
rect 11582 10159 11594 10193
rect 11202 10153 11594 10159
rect 11650 10112 11734 10312
rect 11790 10265 12182 10271
rect 11790 10231 11802 10265
rect 12170 10231 12182 10265
rect 11790 10193 12182 10231
rect 11790 10159 11802 10193
rect 12170 10159 12182 10193
rect 11790 10153 12182 10159
rect 12238 10112 12322 10312
rect 12378 10265 12770 10271
rect 12378 10231 12390 10265
rect 12758 10231 12770 10265
rect 12378 10193 12770 10231
rect 12378 10159 12390 10193
rect 12758 10159 12770 10193
rect 12378 10153 12770 10159
rect 12826 10112 12910 10312
rect 12966 10265 13358 10271
rect 12966 10231 12978 10265
rect 13346 10231 13358 10265
rect 12966 10193 13358 10231
rect 12966 10159 12978 10193
rect 13346 10159 13358 10193
rect 12966 10153 13358 10159
rect 13414 10112 13498 10312
rect 13554 10265 13946 10271
rect 13554 10231 13566 10265
rect 13934 10231 13946 10265
rect 13554 10193 13946 10231
rect 13554 10159 13566 10193
rect 13934 10159 13946 10193
rect 13554 10153 13946 10159
rect 14002 10112 14086 10312
rect 14142 10265 14534 10271
rect 14142 10231 14154 10265
rect 14522 10231 14534 10265
rect 14142 10193 14534 10231
rect 14142 10159 14154 10193
rect 14522 10159 14534 10193
rect 14142 10153 14534 10159
rect 14590 10112 14674 10312
rect 14730 10265 15122 10271
rect 14730 10231 14742 10265
rect 15110 10231 15122 10265
rect 14730 10193 15122 10231
rect 14730 10159 14742 10193
rect 15110 10159 15122 10193
rect 14730 10153 15122 10159
rect 15178 10112 15262 10312
rect 15318 10265 15710 10271
rect 15318 10231 15330 10265
rect 15698 10231 15710 10265
rect 15318 10193 15710 10231
rect 15318 10159 15330 10193
rect 15698 10159 15710 10193
rect 15318 10153 15710 10159
rect 15766 10112 15850 10312
rect 15906 10265 16298 10271
rect 15906 10231 15918 10265
rect 16286 10231 16298 10265
rect 15906 10193 16298 10231
rect 15906 10159 15918 10193
rect 16286 10159 16298 10193
rect 15906 10153 16298 10159
rect 16354 10112 16438 10312
rect 16494 10265 16886 10271
rect 16494 10231 16506 10265
rect 16874 10231 16886 10265
rect 16494 10193 16886 10231
rect 16494 10159 16506 10193
rect 16874 10159 16886 10193
rect 16494 10153 16886 10159
rect 16942 10112 17026 10312
rect 17082 10265 17474 10271
rect 17082 10231 17094 10265
rect 17462 10231 17474 10265
rect 17082 10193 17474 10231
rect 17082 10159 17094 10193
rect 17462 10159 17474 10193
rect 17082 10153 17474 10159
rect 17530 10112 17614 10312
rect 17670 10265 18062 10271
rect 17670 10231 17682 10265
rect 18050 10231 18062 10265
rect 17670 10193 18062 10231
rect 17670 10159 17682 10193
rect 18050 10159 18062 10193
rect 17670 10153 18062 10159
rect 18118 10112 18202 10312
rect 18258 10265 18650 10271
rect 18258 10231 18270 10265
rect 18638 10231 18650 10265
rect 18258 10193 18650 10231
rect 18258 10159 18270 10193
rect 18638 10159 18650 10193
rect 18258 10153 18650 10159
rect 18706 10112 18790 10312
rect 18846 10265 19238 10271
rect 18846 10231 18858 10265
rect 19226 10231 19238 10265
rect 18846 10193 19238 10231
rect 18846 10159 18858 10193
rect 19226 10159 19238 10193
rect 18846 10153 19238 10159
rect 19294 10112 19378 10312
rect 19434 10265 19826 10271
rect 19434 10231 19446 10265
rect 19814 10231 19826 10265
rect 19434 10193 19826 10231
rect 19434 10159 19446 10193
rect 19814 10159 19826 10193
rect 19434 10153 19826 10159
rect 19882 10112 19966 10312
rect 20022 10265 20414 10271
rect 20022 10231 20034 10265
rect 20402 10231 20414 10265
rect 20022 10193 20414 10231
rect 20022 10159 20034 10193
rect 20402 10159 20414 10193
rect 20022 10153 20414 10159
rect 20470 10112 20554 10312
rect 20610 10265 21002 10271
rect 20610 10231 20622 10265
rect 20990 10231 21002 10265
rect 20610 10193 21002 10231
rect 20610 10159 20622 10193
rect 20990 10159 21002 10193
rect 20610 10153 21002 10159
rect 21058 10112 21142 10312
rect 21198 10265 21590 10271
rect 21198 10231 21210 10265
rect 21578 10231 21590 10265
rect 21198 10193 21590 10231
rect 21198 10159 21210 10193
rect 21578 10159 21590 10193
rect 21198 10153 21590 10159
rect 21646 10112 21730 10312
rect 21786 10265 22178 10271
rect 21786 10231 21798 10265
rect 22166 10231 22178 10265
rect 21786 10193 22178 10231
rect 21786 10159 21798 10193
rect 22166 10159 22178 10193
rect 21786 10153 22178 10159
rect 22228 10112 22286 10312
rect 22374 10265 22766 10271
rect 22374 10231 22386 10265
rect 22754 10231 22766 10265
rect 22374 10193 22766 10231
rect 22374 10159 22386 10193
rect 22754 10159 22766 10193
rect 22374 10153 22766 10159
rect 22822 10112 22906 10312
rect 22962 10265 23354 10271
rect 22962 10231 22974 10265
rect 23342 10231 23354 10265
rect 22962 10193 23354 10231
rect 22962 10159 22974 10193
rect 23342 10159 23354 10193
rect 22962 10153 23354 10159
rect 23410 10112 23494 10312
rect 23550 10265 23942 10271
rect 23550 10231 23562 10265
rect 23930 10231 23942 10265
rect 23550 10193 23942 10231
rect 23550 10159 23562 10193
rect 23930 10159 23942 10193
rect 23550 10153 23942 10159
rect 23998 10112 24082 10312
rect 24138 10265 24530 10271
rect 24138 10231 24150 10265
rect 24518 10231 24530 10265
rect 24138 10193 24530 10231
rect 24138 10159 24150 10193
rect 24518 10159 24530 10193
rect 24138 10153 24530 10159
rect 24726 10265 25118 10271
rect 24726 10231 24738 10265
rect 25106 10231 25118 10265
rect 24726 10193 25118 10231
rect 24726 10159 24738 10193
rect 25106 10159 25118 10193
rect 24726 10153 25118 10159
rect 25174 10112 25258 10312
rect 25314 10265 25706 10271
rect 25314 10231 25326 10265
rect 25694 10231 25706 10265
rect 25314 10193 25706 10231
rect 25314 10159 25326 10193
rect 25694 10159 25706 10193
rect 25314 10153 25706 10159
rect 25762 10112 25846 10312
rect 25902 10265 26294 10271
rect 25902 10231 25914 10265
rect 26282 10231 26294 10265
rect 25902 10193 26294 10231
rect 25902 10159 25914 10193
rect 26282 10159 26294 10193
rect 25902 10153 26294 10159
rect 26350 10112 26434 10312
rect 26490 10265 26882 10271
rect 26490 10231 26502 10265
rect 26870 10231 26882 10265
rect 26490 10193 26882 10231
rect 26490 10159 26502 10193
rect 26870 10159 26882 10193
rect 26490 10153 26882 10159
rect 26972 10112 27028 10312
rect 27078 10265 27470 10271
rect 27078 10231 27090 10265
rect 27458 10231 27470 10265
rect 27078 10193 27470 10231
rect 27078 10159 27090 10193
rect 27458 10159 27470 10193
rect 27078 10153 27470 10159
rect 27526 10112 27610 10312
rect 27666 10265 28058 10271
rect 27666 10231 27678 10265
rect 28046 10231 28058 10265
rect 27666 10193 28058 10231
rect 27666 10159 27678 10193
rect 28046 10159 28058 10193
rect 27666 10153 28058 10159
rect 28114 10112 28198 10312
rect 28254 10265 28646 10271
rect 28254 10231 28266 10265
rect 28634 10231 28646 10265
rect 28254 10193 28646 10231
rect 28254 10159 28266 10193
rect 28634 10159 28646 10193
rect 28254 10153 28646 10159
rect 28702 10112 28786 10312
rect 28842 10265 29234 10271
rect 28842 10231 28854 10265
rect 29222 10231 29234 10265
rect 28842 10193 29234 10231
rect 28842 10159 28854 10193
rect 29222 10159 29234 10193
rect 28842 10153 29234 10159
rect 29290 10112 29374 10312
rect 29430 10265 29822 10271
rect 29430 10231 29442 10265
rect 29810 10231 29822 10265
rect 29430 10193 29822 10231
rect 29430 10159 29442 10193
rect 29810 10159 29822 10193
rect 29430 10153 29822 10159
rect 29878 10112 29962 10312
rect 30018 10265 30410 10271
rect 30018 10231 30030 10265
rect 30398 10231 30410 10265
rect 30018 10193 30410 10231
rect 30018 10159 30030 10193
rect 30398 10159 30410 10193
rect 30018 10153 30410 10159
rect 30466 10112 30550 10312
rect 30606 10265 30998 10271
rect 30606 10231 30618 10265
rect 30986 10231 30998 10265
rect 30606 10193 30998 10231
rect 30606 10159 30618 10193
rect 30986 10159 30998 10193
rect 30606 10153 30998 10159
rect 31054 10112 31138 10312
rect 31194 10265 31586 10271
rect 31194 10231 31206 10265
rect 31574 10231 31586 10265
rect 31194 10193 31586 10231
rect 31194 10159 31206 10193
rect 31574 10159 31586 10193
rect 31194 10153 31586 10159
rect 31642 10112 31726 10312
rect 31782 10265 32174 10271
rect 31782 10231 31794 10265
rect 32162 10231 32174 10265
rect 31782 10193 32174 10231
rect 31782 10159 31794 10193
rect 32162 10159 32174 10193
rect 31782 10153 32174 10159
rect 32230 10112 32314 10312
rect 32370 10265 32762 10271
rect 32370 10231 32382 10265
rect 32750 10231 32762 10265
rect 32370 10193 32762 10231
rect 32370 10159 32382 10193
rect 32750 10159 32762 10193
rect 32370 10153 32762 10159
rect 32818 10112 32902 10312
rect 32958 10265 33350 10271
rect 32958 10231 32970 10265
rect 33338 10231 33350 10265
rect 32958 10193 33350 10231
rect 32958 10159 32970 10193
rect 33338 10159 33350 10193
rect 32958 10153 33350 10159
rect 33406 10112 33490 10312
rect 33546 10265 33938 10271
rect 33546 10231 33558 10265
rect 33926 10231 33938 10265
rect 33546 10193 33938 10231
rect 33546 10159 33558 10193
rect 33926 10159 33938 10193
rect 33546 10153 33938 10159
rect 33994 10112 34078 10312
rect 34134 10265 34526 10271
rect 34134 10231 34146 10265
rect 34514 10231 34526 10265
rect 34134 10193 34526 10231
rect 34134 10159 34146 10193
rect 34514 10159 34526 10193
rect 34134 10153 34526 10159
rect 34582 10112 34666 10312
rect 34722 10265 35114 10271
rect 34722 10231 34734 10265
rect 35102 10231 35114 10265
rect 34722 10193 35114 10231
rect 34722 10159 34734 10193
rect 35102 10159 35114 10193
rect 34722 10153 35114 10159
rect 35170 10112 35254 10312
rect 35310 10265 35702 10271
rect 35310 10231 35322 10265
rect 35690 10231 35702 10265
rect 35310 10193 35702 10231
rect 35310 10159 35322 10193
rect 35690 10159 35702 10193
rect 35310 10153 35702 10159
rect 35758 10112 35842 10312
rect 35898 10265 36290 10271
rect 35898 10231 35910 10265
rect 36278 10231 36290 10265
rect 35898 10193 36290 10231
rect 35898 10159 35910 10193
rect 36278 10159 36290 10193
rect 35898 10153 36290 10159
rect 36346 10112 36430 10312
rect 36486 10265 36878 10271
rect 36486 10231 36498 10265
rect 36866 10231 36878 10265
rect 36486 10193 36878 10231
rect 36486 10159 36498 10193
rect 36866 10159 36878 10193
rect 36486 10153 36878 10159
rect 36934 10112 37018 10312
rect 37074 10265 37466 10271
rect 37074 10231 37086 10265
rect 37454 10231 37466 10265
rect 37074 10193 37466 10231
rect 37074 10159 37086 10193
rect 37454 10159 37466 10193
rect 37074 10153 37466 10159
rect 37522 10112 37606 10312
rect 37662 10265 38054 10271
rect 37662 10231 37674 10265
rect 38042 10231 38054 10265
rect 37662 10193 38054 10231
rect 37662 10159 37674 10193
rect 38042 10159 38054 10193
rect 37662 10153 38054 10159
rect 38110 10112 38194 10312
rect 38250 10265 38642 10271
rect 38250 10231 38262 10265
rect 38630 10231 38642 10265
rect 38250 10193 38642 10231
rect 38250 10159 38262 10193
rect 38630 10159 38642 10193
rect 38250 10153 38642 10159
rect 38698 10112 38782 10312
rect 10474 10100 10604 10112
rect 10474 9324 10564 10100
rect 10598 9324 10604 10100
rect 10474 9312 10604 9324
rect 11016 10100 11192 10112
rect 11016 9324 11022 10100
rect 11056 9324 11152 10100
rect 11186 9324 11192 10100
rect 11016 9312 11192 9324
rect 11604 10100 11780 10112
rect 11604 9324 11610 10100
rect 11644 9324 11740 10100
rect 11774 9324 11780 10100
rect 11604 9312 11780 9324
rect 12192 10100 12368 10112
rect 12192 9324 12198 10100
rect 12232 9324 12328 10100
rect 12362 9324 12368 10100
rect 12192 9312 12368 9324
rect 12780 10100 12956 10112
rect 12780 9324 12786 10100
rect 12820 9324 12916 10100
rect 12950 9324 12956 10100
rect 12780 9312 12956 9324
rect 13368 10100 13544 10112
rect 13368 9324 13374 10100
rect 13408 9324 13504 10100
rect 13538 9324 13544 10100
rect 13368 9312 13544 9324
rect 13956 10100 14132 10112
rect 13956 9324 13962 10100
rect 13996 9324 14092 10100
rect 14126 9324 14132 10100
rect 13956 9312 14132 9324
rect 14544 10100 14720 10112
rect 14544 9324 14550 10100
rect 14584 9324 14680 10100
rect 14714 9324 14720 10100
rect 14544 9312 14720 9324
rect 15132 10100 15308 10112
rect 15132 9324 15138 10100
rect 15172 9324 15268 10100
rect 15302 9324 15308 10100
rect 15132 9312 15308 9324
rect 15720 10100 15896 10112
rect 15720 9324 15726 10100
rect 15760 9324 15856 10100
rect 15890 9324 15896 10100
rect 15720 9312 15896 9324
rect 16308 10100 16484 10112
rect 16308 9324 16314 10100
rect 16348 9324 16444 10100
rect 16478 9324 16484 10100
rect 16308 9312 16484 9324
rect 16896 10100 17072 10112
rect 16896 9324 16902 10100
rect 16936 9324 17032 10100
rect 17066 9324 17072 10100
rect 16896 9312 17072 9324
rect 17484 10100 17660 10112
rect 17484 9324 17490 10100
rect 17524 9324 17620 10100
rect 17654 9324 17660 10100
rect 17484 9312 17660 9324
rect 18072 10100 18248 10112
rect 18072 9324 18078 10100
rect 18112 9324 18208 10100
rect 18242 9324 18248 10100
rect 18072 9312 18248 9324
rect 18660 10100 18836 10112
rect 18660 9324 18666 10100
rect 18700 9324 18796 10100
rect 18830 9324 18836 10100
rect 18660 9312 18836 9324
rect 19248 10100 19424 10112
rect 19248 9324 19254 10100
rect 19288 9324 19384 10100
rect 19418 9324 19424 10100
rect 19248 9312 19424 9324
rect 19836 10100 20012 10112
rect 19836 9324 19842 10100
rect 19876 9324 19972 10100
rect 20006 9324 20012 10100
rect 19836 9312 20012 9324
rect 20424 10100 20600 10112
rect 20424 9324 20430 10100
rect 20464 9324 20560 10100
rect 20594 9324 20600 10100
rect 20424 9312 20600 9324
rect 21012 10100 21188 10112
rect 21012 9324 21018 10100
rect 21052 9324 21148 10100
rect 21182 9324 21188 10100
rect 21012 9312 21188 9324
rect 21600 10100 21776 10112
rect 21600 9324 21606 10100
rect 21640 9324 21736 10100
rect 21770 9324 21776 10100
rect 21600 9312 21776 9324
rect 22188 10100 22286 10112
rect 22188 9324 22194 10100
rect 22228 9324 22286 10100
rect 22188 9312 22286 9324
rect 22318 10100 22364 10112
rect 22318 9324 22324 10100
rect 22358 9324 22364 10100
rect 22318 9312 22364 9324
rect 22776 10100 22952 10112
rect 22776 9324 22782 10100
rect 22816 9324 22912 10100
rect 22946 9324 22952 10100
rect 22776 9312 22952 9324
rect 23364 10100 23540 10112
rect 23364 9324 23370 10100
rect 23404 9324 23500 10100
rect 23534 9324 23540 10100
rect 23364 9312 23540 9324
rect 23952 10100 24128 10112
rect 23952 9324 23958 10100
rect 23992 9324 24088 10100
rect 24122 9324 24128 10100
rect 23952 9312 24128 9324
rect 24540 10100 24586 10112
rect 24540 9324 24546 10100
rect 24580 9324 24586 10100
rect 24540 9312 24586 9324
rect 24670 10100 24716 10112
rect 24670 9324 24676 10100
rect 24710 9324 24716 10100
rect 24670 9312 24716 9324
rect 25128 10100 25304 10112
rect 25128 9324 25134 10100
rect 25168 9324 25264 10100
rect 25298 9324 25304 10100
rect 25128 9312 25304 9324
rect 25716 10100 25892 10112
rect 25716 9324 25722 10100
rect 25756 9324 25852 10100
rect 25886 9324 25892 10100
rect 25716 9312 25892 9324
rect 26304 10100 26480 10112
rect 26304 9324 26310 10100
rect 26344 9324 26440 10100
rect 26474 9324 26480 10100
rect 26304 9312 26480 9324
rect 26892 10100 26938 10112
rect 26892 9324 26898 10100
rect 26932 9324 26938 10100
rect 26892 9312 26938 9324
rect 26972 10100 27068 10112
rect 26972 9324 27028 10100
rect 27062 9324 27068 10100
rect 26972 9312 27068 9324
rect 27480 10100 27656 10112
rect 27480 9324 27486 10100
rect 27520 9324 27616 10100
rect 27650 9324 27656 10100
rect 27480 9312 27656 9324
rect 28068 10100 28244 10112
rect 28068 9324 28074 10100
rect 28108 9324 28204 10100
rect 28238 9324 28244 10100
rect 28068 9312 28244 9324
rect 28656 10100 28832 10112
rect 28656 9324 28662 10100
rect 28696 9324 28792 10100
rect 28826 9324 28832 10100
rect 28656 9312 28832 9324
rect 29244 10100 29420 10112
rect 29244 9324 29250 10100
rect 29284 9324 29380 10100
rect 29414 9324 29420 10100
rect 29244 9312 29420 9324
rect 29832 10100 30008 10112
rect 29832 9324 29838 10100
rect 29872 9324 29968 10100
rect 30002 9324 30008 10100
rect 29832 9312 30008 9324
rect 30420 10100 30596 10112
rect 30420 9324 30426 10100
rect 30460 9324 30556 10100
rect 30590 9324 30596 10100
rect 30420 9312 30596 9324
rect 31008 10100 31184 10112
rect 31008 9324 31014 10100
rect 31048 9324 31144 10100
rect 31178 9324 31184 10100
rect 31008 9312 31184 9324
rect 31596 10100 31772 10112
rect 31596 9324 31602 10100
rect 31636 9324 31732 10100
rect 31766 9324 31772 10100
rect 31596 9312 31772 9324
rect 32184 10100 32360 10112
rect 32184 9324 32190 10100
rect 32224 9324 32320 10100
rect 32354 9324 32360 10100
rect 32184 9312 32360 9324
rect 32772 10100 32948 10112
rect 32772 9324 32778 10100
rect 32812 9324 32908 10100
rect 32942 9324 32948 10100
rect 32772 9312 32948 9324
rect 33360 10100 33536 10112
rect 33360 9324 33366 10100
rect 33400 9324 33496 10100
rect 33530 9324 33536 10100
rect 33360 9312 33536 9324
rect 33948 10100 34124 10112
rect 33948 9324 33954 10100
rect 33988 9324 34084 10100
rect 34118 9324 34124 10100
rect 33948 9312 34124 9324
rect 34536 10100 34712 10112
rect 34536 9324 34542 10100
rect 34576 9324 34672 10100
rect 34706 9324 34712 10100
rect 34536 9312 34712 9324
rect 35124 10100 35300 10112
rect 35124 9324 35130 10100
rect 35164 9324 35260 10100
rect 35294 9324 35300 10100
rect 35124 9312 35300 9324
rect 35712 10100 35888 10112
rect 35712 9324 35718 10100
rect 35752 9324 35848 10100
rect 35882 9324 35888 10100
rect 35712 9312 35888 9324
rect 36300 10100 36476 10112
rect 36300 9324 36306 10100
rect 36340 9324 36436 10100
rect 36470 9324 36476 10100
rect 36300 9312 36476 9324
rect 36888 10100 37064 10112
rect 36888 9324 36894 10100
rect 36928 9324 37024 10100
rect 37058 9324 37064 10100
rect 36888 9312 37064 9324
rect 37476 10100 37652 10112
rect 37476 9324 37482 10100
rect 37516 9324 37612 10100
rect 37646 9324 37652 10100
rect 37476 9312 37652 9324
rect 38064 10100 38240 10112
rect 38064 9324 38070 10100
rect 38104 9324 38200 10100
rect 38234 9324 38240 10100
rect 38064 9312 38240 9324
rect 38652 10100 38782 10112
rect 38652 9324 38658 10100
rect 38692 9324 38782 10100
rect 38652 9312 38782 9324
rect 10474 9112 10558 9312
rect 10614 9265 11006 9271
rect 10614 9231 10626 9265
rect 10994 9231 11006 9265
rect 10614 9193 11006 9231
rect 10614 9159 10626 9193
rect 10994 9159 11006 9193
rect 10614 9153 11006 9159
rect 11062 9112 11146 9312
rect 11202 9265 11594 9271
rect 11202 9231 11214 9265
rect 11582 9231 11594 9265
rect 11202 9193 11594 9231
rect 11202 9159 11214 9193
rect 11582 9159 11594 9193
rect 11202 9153 11594 9159
rect 11650 9112 11734 9312
rect 11790 9265 12182 9271
rect 11790 9231 11802 9265
rect 12170 9231 12182 9265
rect 11790 9193 12182 9231
rect 11790 9159 11802 9193
rect 12170 9159 12182 9193
rect 11790 9153 12182 9159
rect 12238 9112 12322 9312
rect 12378 9265 12770 9271
rect 12378 9231 12390 9265
rect 12758 9231 12770 9265
rect 12378 9193 12770 9231
rect 12378 9159 12390 9193
rect 12758 9159 12770 9193
rect 12378 9153 12770 9159
rect 12826 9112 12910 9312
rect 12966 9265 13358 9271
rect 12966 9231 12978 9265
rect 13346 9231 13358 9265
rect 12966 9193 13358 9231
rect 12966 9159 12978 9193
rect 13346 9159 13358 9193
rect 12966 9153 13358 9159
rect 13414 9112 13498 9312
rect 13554 9265 13946 9271
rect 13554 9231 13566 9265
rect 13934 9231 13946 9265
rect 13554 9193 13946 9231
rect 13554 9159 13566 9193
rect 13934 9159 13946 9193
rect 13554 9153 13946 9159
rect 14002 9112 14086 9312
rect 14142 9265 14534 9271
rect 14142 9231 14154 9265
rect 14522 9231 14534 9265
rect 14142 9193 14534 9231
rect 14142 9159 14154 9193
rect 14522 9159 14534 9193
rect 14142 9153 14534 9159
rect 14590 9112 14674 9312
rect 14730 9265 15122 9271
rect 14730 9231 14742 9265
rect 15110 9231 15122 9265
rect 14730 9193 15122 9231
rect 14730 9159 14742 9193
rect 15110 9159 15122 9193
rect 14730 9153 15122 9159
rect 15178 9112 15262 9312
rect 15318 9265 15710 9271
rect 15318 9231 15330 9265
rect 15698 9231 15710 9265
rect 15318 9193 15710 9231
rect 15318 9159 15330 9193
rect 15698 9159 15710 9193
rect 15318 9153 15710 9159
rect 15766 9112 15850 9312
rect 15906 9265 16298 9271
rect 15906 9231 15918 9265
rect 16286 9231 16298 9265
rect 15906 9193 16298 9231
rect 15906 9159 15918 9193
rect 16286 9159 16298 9193
rect 15906 9153 16298 9159
rect 16354 9112 16438 9312
rect 16494 9265 16886 9271
rect 16494 9231 16506 9265
rect 16874 9231 16886 9265
rect 16494 9193 16886 9231
rect 16494 9159 16506 9193
rect 16874 9159 16886 9193
rect 16494 9153 16886 9159
rect 16942 9112 17026 9312
rect 17082 9265 17474 9271
rect 17082 9231 17094 9265
rect 17462 9231 17474 9265
rect 17082 9193 17474 9231
rect 17082 9159 17094 9193
rect 17462 9159 17474 9193
rect 17082 9153 17474 9159
rect 17530 9112 17614 9312
rect 17670 9265 18062 9271
rect 17670 9231 17682 9265
rect 18050 9231 18062 9265
rect 17670 9193 18062 9231
rect 17670 9159 17682 9193
rect 18050 9159 18062 9193
rect 17670 9153 18062 9159
rect 18118 9112 18202 9312
rect 18258 9265 18650 9271
rect 18258 9231 18270 9265
rect 18638 9231 18650 9265
rect 18258 9193 18650 9231
rect 18258 9159 18270 9193
rect 18638 9159 18650 9193
rect 18258 9153 18650 9159
rect 18706 9112 18790 9312
rect 18846 9265 19238 9271
rect 18846 9231 18858 9265
rect 19226 9231 19238 9265
rect 18846 9193 19238 9231
rect 18846 9159 18858 9193
rect 19226 9159 19238 9193
rect 18846 9153 19238 9159
rect 19294 9112 19378 9312
rect 19434 9265 19826 9271
rect 19434 9231 19446 9265
rect 19814 9231 19826 9265
rect 19434 9193 19826 9231
rect 19434 9159 19446 9193
rect 19814 9159 19826 9193
rect 19434 9153 19826 9159
rect 19882 9112 19966 9312
rect 20022 9265 20414 9271
rect 20022 9231 20034 9265
rect 20402 9231 20414 9265
rect 20022 9193 20414 9231
rect 20022 9159 20034 9193
rect 20402 9159 20414 9193
rect 20022 9153 20414 9159
rect 20470 9112 20554 9312
rect 20610 9265 21002 9271
rect 20610 9231 20622 9265
rect 20990 9231 21002 9265
rect 20610 9193 21002 9231
rect 20610 9159 20622 9193
rect 20990 9159 21002 9193
rect 20610 9153 21002 9159
rect 21058 9112 21142 9312
rect 21198 9265 21590 9271
rect 21198 9231 21210 9265
rect 21578 9231 21590 9265
rect 21198 9193 21590 9231
rect 21198 9159 21210 9193
rect 21578 9159 21590 9193
rect 21198 9153 21590 9159
rect 21646 9112 21730 9312
rect 21786 9265 22178 9271
rect 21786 9231 21798 9265
rect 22166 9231 22178 9265
rect 21786 9193 22178 9231
rect 21786 9159 21798 9193
rect 22166 9159 22178 9193
rect 21786 9153 22178 9159
rect 22228 9112 22286 9312
rect 22374 9265 22766 9271
rect 22374 9231 22386 9265
rect 22754 9231 22766 9265
rect 22374 9193 22766 9231
rect 22374 9159 22386 9193
rect 22754 9159 22766 9193
rect 22374 9153 22766 9159
rect 22822 9112 22906 9312
rect 22962 9265 23354 9271
rect 22962 9231 22974 9265
rect 23342 9231 23354 9265
rect 22962 9193 23354 9231
rect 22962 9159 22974 9193
rect 23342 9159 23354 9193
rect 22962 9153 23354 9159
rect 23410 9112 23494 9312
rect 23550 9265 23942 9271
rect 23550 9231 23562 9265
rect 23930 9231 23942 9265
rect 23550 9193 23942 9231
rect 23550 9159 23562 9193
rect 23930 9159 23942 9193
rect 23550 9153 23942 9159
rect 23998 9112 24082 9312
rect 24138 9265 24530 9271
rect 24138 9231 24150 9265
rect 24518 9231 24530 9265
rect 24138 9193 24530 9231
rect 24138 9159 24150 9193
rect 24518 9159 24530 9193
rect 24138 9153 24530 9159
rect 24726 9265 25118 9271
rect 24726 9231 24738 9265
rect 25106 9231 25118 9265
rect 24726 9193 25118 9231
rect 24726 9159 24738 9193
rect 25106 9159 25118 9193
rect 24726 9153 25118 9159
rect 25174 9112 25258 9312
rect 25314 9265 25706 9271
rect 25314 9231 25326 9265
rect 25694 9231 25706 9265
rect 25314 9193 25706 9231
rect 25314 9159 25326 9193
rect 25694 9159 25706 9193
rect 25314 9153 25706 9159
rect 25762 9112 25846 9312
rect 25902 9265 26294 9271
rect 25902 9231 25914 9265
rect 26282 9231 26294 9265
rect 25902 9193 26294 9231
rect 25902 9159 25914 9193
rect 26282 9159 26294 9193
rect 25902 9153 26294 9159
rect 26350 9112 26434 9312
rect 26490 9265 26882 9271
rect 26490 9231 26502 9265
rect 26870 9231 26882 9265
rect 26490 9193 26882 9231
rect 26490 9159 26502 9193
rect 26870 9159 26882 9193
rect 26490 9153 26882 9159
rect 26972 9112 27028 9312
rect 27078 9265 27470 9271
rect 27078 9231 27090 9265
rect 27458 9231 27470 9265
rect 27078 9193 27470 9231
rect 27078 9159 27090 9193
rect 27458 9159 27470 9193
rect 27078 9153 27470 9159
rect 27526 9112 27610 9312
rect 27666 9265 28058 9271
rect 27666 9231 27678 9265
rect 28046 9231 28058 9265
rect 27666 9193 28058 9231
rect 27666 9159 27678 9193
rect 28046 9159 28058 9193
rect 27666 9153 28058 9159
rect 28114 9112 28198 9312
rect 28254 9265 28646 9271
rect 28254 9231 28266 9265
rect 28634 9231 28646 9265
rect 28254 9193 28646 9231
rect 28254 9159 28266 9193
rect 28634 9159 28646 9193
rect 28254 9153 28646 9159
rect 28702 9112 28786 9312
rect 28842 9265 29234 9271
rect 28842 9231 28854 9265
rect 29222 9231 29234 9265
rect 28842 9193 29234 9231
rect 28842 9159 28854 9193
rect 29222 9159 29234 9193
rect 28842 9153 29234 9159
rect 29290 9112 29374 9312
rect 29430 9265 29822 9271
rect 29430 9231 29442 9265
rect 29810 9231 29822 9265
rect 29430 9193 29822 9231
rect 29430 9159 29442 9193
rect 29810 9159 29822 9193
rect 29430 9153 29822 9159
rect 29878 9112 29962 9312
rect 30018 9265 30410 9271
rect 30018 9231 30030 9265
rect 30398 9231 30410 9265
rect 30018 9193 30410 9231
rect 30018 9159 30030 9193
rect 30398 9159 30410 9193
rect 30018 9153 30410 9159
rect 30466 9112 30550 9312
rect 30606 9265 30998 9271
rect 30606 9231 30618 9265
rect 30986 9231 30998 9265
rect 30606 9193 30998 9231
rect 30606 9159 30618 9193
rect 30986 9159 30998 9193
rect 30606 9153 30998 9159
rect 31054 9112 31138 9312
rect 31194 9265 31586 9271
rect 31194 9231 31206 9265
rect 31574 9231 31586 9265
rect 31194 9193 31586 9231
rect 31194 9159 31206 9193
rect 31574 9159 31586 9193
rect 31194 9153 31586 9159
rect 31642 9112 31726 9312
rect 31782 9265 32174 9271
rect 31782 9231 31794 9265
rect 32162 9231 32174 9265
rect 31782 9193 32174 9231
rect 31782 9159 31794 9193
rect 32162 9159 32174 9193
rect 31782 9153 32174 9159
rect 32230 9112 32314 9312
rect 32370 9265 32762 9271
rect 32370 9231 32382 9265
rect 32750 9231 32762 9265
rect 32370 9193 32762 9231
rect 32370 9159 32382 9193
rect 32750 9159 32762 9193
rect 32370 9153 32762 9159
rect 32818 9112 32902 9312
rect 32958 9265 33350 9271
rect 32958 9231 32970 9265
rect 33338 9231 33350 9265
rect 32958 9193 33350 9231
rect 32958 9159 32970 9193
rect 33338 9159 33350 9193
rect 32958 9153 33350 9159
rect 33406 9112 33490 9312
rect 33546 9265 33938 9271
rect 33546 9231 33558 9265
rect 33926 9231 33938 9265
rect 33546 9193 33938 9231
rect 33546 9159 33558 9193
rect 33926 9159 33938 9193
rect 33546 9153 33938 9159
rect 33994 9112 34078 9312
rect 34134 9265 34526 9271
rect 34134 9231 34146 9265
rect 34514 9231 34526 9265
rect 34134 9193 34526 9231
rect 34134 9159 34146 9193
rect 34514 9159 34526 9193
rect 34134 9153 34526 9159
rect 34582 9112 34666 9312
rect 34722 9265 35114 9271
rect 34722 9231 34734 9265
rect 35102 9231 35114 9265
rect 34722 9193 35114 9231
rect 34722 9159 34734 9193
rect 35102 9159 35114 9193
rect 34722 9153 35114 9159
rect 35170 9112 35254 9312
rect 35310 9265 35702 9271
rect 35310 9231 35322 9265
rect 35690 9231 35702 9265
rect 35310 9193 35702 9231
rect 35310 9159 35322 9193
rect 35690 9159 35702 9193
rect 35310 9153 35702 9159
rect 35758 9112 35842 9312
rect 35898 9265 36290 9271
rect 35898 9231 35910 9265
rect 36278 9231 36290 9265
rect 35898 9193 36290 9231
rect 35898 9159 35910 9193
rect 36278 9159 36290 9193
rect 35898 9153 36290 9159
rect 36346 9112 36430 9312
rect 36486 9265 36878 9271
rect 36486 9231 36498 9265
rect 36866 9231 36878 9265
rect 36486 9193 36878 9231
rect 36486 9159 36498 9193
rect 36866 9159 36878 9193
rect 36486 9153 36878 9159
rect 36934 9112 37018 9312
rect 37074 9265 37466 9271
rect 37074 9231 37086 9265
rect 37454 9231 37466 9265
rect 37074 9193 37466 9231
rect 37074 9159 37086 9193
rect 37454 9159 37466 9193
rect 37074 9153 37466 9159
rect 37522 9112 37606 9312
rect 37662 9265 38054 9271
rect 37662 9231 37674 9265
rect 38042 9231 38054 9265
rect 37662 9193 38054 9231
rect 37662 9159 37674 9193
rect 38042 9159 38054 9193
rect 37662 9153 38054 9159
rect 38110 9112 38194 9312
rect 38250 9265 38642 9271
rect 38250 9231 38262 9265
rect 38630 9231 38642 9265
rect 38250 9193 38642 9231
rect 38250 9159 38262 9193
rect 38630 9159 38642 9193
rect 38250 9153 38642 9159
rect 38698 9112 38782 9312
rect 10474 9100 10604 9112
rect 10474 8324 10564 9100
rect 10598 8324 10604 9100
rect 10474 8312 10604 8324
rect 11016 9100 11192 9112
rect 11016 8324 11022 9100
rect 11056 8324 11152 9100
rect 11186 8324 11192 9100
rect 11016 8312 11192 8324
rect 11604 9100 11780 9112
rect 11604 8324 11610 9100
rect 11644 8324 11740 9100
rect 11774 8324 11780 9100
rect 11604 8312 11780 8324
rect 12192 9100 12368 9112
rect 12192 8324 12198 9100
rect 12232 8324 12328 9100
rect 12362 8324 12368 9100
rect 12192 8312 12368 8324
rect 12780 9100 12956 9112
rect 12780 8324 12786 9100
rect 12820 8324 12916 9100
rect 12950 8324 12956 9100
rect 12780 8312 12956 8324
rect 13368 9100 13544 9112
rect 13368 8324 13374 9100
rect 13408 8324 13504 9100
rect 13538 8324 13544 9100
rect 13368 8312 13544 8324
rect 13956 9100 14132 9112
rect 13956 8324 13962 9100
rect 13996 8324 14092 9100
rect 14126 8324 14132 9100
rect 13956 8312 14132 8324
rect 14544 9100 14720 9112
rect 14544 8324 14550 9100
rect 14584 8324 14680 9100
rect 14714 8324 14720 9100
rect 14544 8312 14720 8324
rect 15132 9100 15308 9112
rect 15132 8324 15138 9100
rect 15172 8324 15268 9100
rect 15302 8324 15308 9100
rect 15132 8312 15308 8324
rect 15720 9100 15896 9112
rect 15720 8324 15726 9100
rect 15760 8324 15856 9100
rect 15890 8324 15896 9100
rect 15720 8312 15896 8324
rect 16308 9100 16484 9112
rect 16308 8324 16314 9100
rect 16348 8324 16444 9100
rect 16478 8324 16484 9100
rect 16308 8312 16484 8324
rect 16896 9100 17072 9112
rect 16896 8324 16902 9100
rect 16936 8324 17032 9100
rect 17066 8324 17072 9100
rect 16896 8312 17072 8324
rect 17484 9100 17660 9112
rect 17484 8324 17490 9100
rect 17524 8324 17620 9100
rect 17654 8324 17660 9100
rect 17484 8312 17660 8324
rect 18072 9100 18248 9112
rect 18072 8324 18078 9100
rect 18112 8324 18208 9100
rect 18242 8324 18248 9100
rect 18072 8312 18248 8324
rect 18660 9100 18836 9112
rect 18660 8324 18666 9100
rect 18700 8324 18796 9100
rect 18830 8324 18836 9100
rect 18660 8312 18836 8324
rect 19248 9100 19424 9112
rect 19248 8324 19254 9100
rect 19288 8324 19384 9100
rect 19418 8324 19424 9100
rect 19248 8312 19424 8324
rect 19836 9100 20012 9112
rect 19836 8324 19842 9100
rect 19876 8324 19972 9100
rect 20006 8324 20012 9100
rect 19836 8312 20012 8324
rect 20424 9100 20600 9112
rect 20424 8324 20430 9100
rect 20464 8324 20560 9100
rect 20594 8324 20600 9100
rect 20424 8312 20600 8324
rect 21012 9100 21188 9112
rect 21012 8324 21018 9100
rect 21052 8324 21148 9100
rect 21182 8324 21188 9100
rect 21012 8312 21188 8324
rect 21600 9100 21776 9112
rect 21600 8324 21606 9100
rect 21640 8324 21736 9100
rect 21770 8324 21776 9100
rect 21600 8312 21776 8324
rect 22188 9100 22286 9112
rect 22188 8324 22194 9100
rect 22228 8324 22286 9100
rect 22188 8312 22286 8324
rect 22318 9100 22364 9112
rect 22318 8324 22324 9100
rect 22358 8324 22364 9100
rect 22318 8312 22364 8324
rect 22776 9100 22952 9112
rect 22776 8324 22782 9100
rect 22816 8324 22912 9100
rect 22946 8324 22952 9100
rect 22776 8312 22952 8324
rect 23364 9100 23540 9112
rect 23364 8324 23370 9100
rect 23404 8324 23500 9100
rect 23534 8324 23540 9100
rect 23364 8312 23540 8324
rect 23952 9100 24128 9112
rect 23952 8324 23958 9100
rect 23992 8324 24088 9100
rect 24122 8324 24128 9100
rect 23952 8312 24128 8324
rect 24540 9100 24586 9112
rect 24540 8324 24546 9100
rect 24580 8324 24586 9100
rect 24540 8312 24586 8324
rect 24670 9100 24716 9112
rect 24670 8324 24676 9100
rect 24710 8324 24716 9100
rect 24670 8312 24716 8324
rect 25128 9100 25304 9112
rect 25128 8324 25134 9100
rect 25168 8324 25264 9100
rect 25298 8324 25304 9100
rect 25128 8312 25304 8324
rect 25716 9100 25892 9112
rect 25716 8324 25722 9100
rect 25756 8324 25852 9100
rect 25886 8324 25892 9100
rect 25716 8312 25892 8324
rect 26304 9100 26480 9112
rect 26304 8324 26310 9100
rect 26344 8324 26440 9100
rect 26474 8324 26480 9100
rect 26304 8312 26480 8324
rect 26892 9100 26938 9112
rect 26892 8324 26898 9100
rect 26932 8324 26938 9100
rect 26892 8312 26938 8324
rect 26972 9100 27068 9112
rect 26972 8324 27028 9100
rect 27062 8324 27068 9100
rect 26972 8312 27068 8324
rect 27480 9100 27656 9112
rect 27480 8324 27486 9100
rect 27520 8324 27616 9100
rect 27650 8324 27656 9100
rect 27480 8312 27656 8324
rect 28068 9100 28244 9112
rect 28068 8324 28074 9100
rect 28108 8324 28204 9100
rect 28238 8324 28244 9100
rect 28068 8312 28244 8324
rect 28656 9100 28832 9112
rect 28656 8324 28662 9100
rect 28696 8324 28792 9100
rect 28826 8324 28832 9100
rect 28656 8312 28832 8324
rect 29244 9100 29420 9112
rect 29244 8324 29250 9100
rect 29284 8324 29380 9100
rect 29414 8324 29420 9100
rect 29244 8312 29420 8324
rect 29832 9100 30008 9112
rect 29832 8324 29838 9100
rect 29872 8324 29968 9100
rect 30002 8324 30008 9100
rect 29832 8312 30008 8324
rect 30420 9100 30596 9112
rect 30420 8324 30426 9100
rect 30460 8324 30556 9100
rect 30590 8324 30596 9100
rect 30420 8312 30596 8324
rect 31008 9100 31184 9112
rect 31008 8324 31014 9100
rect 31048 8324 31144 9100
rect 31178 8324 31184 9100
rect 31008 8312 31184 8324
rect 31596 9100 31772 9112
rect 31596 8324 31602 9100
rect 31636 8324 31732 9100
rect 31766 8324 31772 9100
rect 31596 8312 31772 8324
rect 32184 9100 32360 9112
rect 32184 8324 32190 9100
rect 32224 8324 32320 9100
rect 32354 8324 32360 9100
rect 32184 8312 32360 8324
rect 32772 9100 32948 9112
rect 32772 8324 32778 9100
rect 32812 8324 32908 9100
rect 32942 8324 32948 9100
rect 32772 8312 32948 8324
rect 33360 9100 33536 9112
rect 33360 8324 33366 9100
rect 33400 8324 33496 9100
rect 33530 8324 33536 9100
rect 33360 8312 33536 8324
rect 33948 9100 34124 9112
rect 33948 8324 33954 9100
rect 33988 8324 34084 9100
rect 34118 8324 34124 9100
rect 33948 8312 34124 8324
rect 34536 9100 34712 9112
rect 34536 8324 34542 9100
rect 34576 8324 34672 9100
rect 34706 8324 34712 9100
rect 34536 8312 34712 8324
rect 35124 9100 35300 9112
rect 35124 8324 35130 9100
rect 35164 8324 35260 9100
rect 35294 8324 35300 9100
rect 35124 8312 35300 8324
rect 35712 9100 35888 9112
rect 35712 8324 35718 9100
rect 35752 8324 35848 9100
rect 35882 8324 35888 9100
rect 35712 8312 35888 8324
rect 36300 9100 36476 9112
rect 36300 8324 36306 9100
rect 36340 8324 36436 9100
rect 36470 8324 36476 9100
rect 36300 8312 36476 8324
rect 36888 9100 37064 9112
rect 36888 8324 36894 9100
rect 36928 8324 37024 9100
rect 37058 8324 37064 9100
rect 36888 8312 37064 8324
rect 37476 9100 37652 9112
rect 37476 8324 37482 9100
rect 37516 8324 37612 9100
rect 37646 8324 37652 9100
rect 37476 8312 37652 8324
rect 38064 9100 38240 9112
rect 38064 8324 38070 9100
rect 38104 8324 38200 9100
rect 38234 8324 38240 9100
rect 38064 8312 38240 8324
rect 38652 9100 38782 9112
rect 38652 8324 38658 9100
rect 38692 8324 38782 9100
rect 38652 8312 38782 8324
rect 10614 8265 11006 8271
rect 10614 8231 10626 8265
rect 10994 8231 11006 8265
rect 10614 8225 11006 8231
rect 11068 7968 11140 8312
rect 11202 8265 11594 8271
rect 11202 8231 11214 8265
rect 11582 8231 11594 8265
rect 11202 8225 11594 8231
rect 11790 8265 12182 8271
rect 11790 8231 11802 8265
rect 12170 8231 12182 8265
rect 11790 8225 12182 8231
rect 12244 7968 12316 8312
rect 12378 8265 12770 8271
rect 12378 8231 12390 8265
rect 12758 8231 12770 8265
rect 12378 8225 12770 8231
rect 12966 8265 13358 8271
rect 12966 8231 12978 8265
rect 13346 8231 13358 8265
rect 12966 8225 13358 8231
rect 13420 7968 13492 8312
rect 13554 8265 13946 8271
rect 13554 8231 13566 8265
rect 13934 8231 13946 8265
rect 13554 8225 13946 8231
rect 14142 8265 14534 8271
rect 14142 8231 14154 8265
rect 14522 8231 14534 8265
rect 14142 8225 14534 8231
rect 14596 7968 14668 8312
rect 14730 8265 15122 8271
rect 14730 8231 14742 8265
rect 15110 8231 15122 8265
rect 14730 8225 15122 8231
rect 15318 8265 15710 8271
rect 15318 8231 15330 8265
rect 15698 8231 15710 8265
rect 15318 8225 15710 8231
rect 15772 7968 15844 8312
rect 15906 8265 16298 8271
rect 15906 8231 15918 8265
rect 16286 8231 16298 8265
rect 15906 8225 16298 8231
rect 16494 8265 16886 8271
rect 16494 8231 16506 8265
rect 16874 8231 16886 8265
rect 16494 8225 16886 8231
rect 16948 7968 17020 8312
rect 17082 8265 17474 8271
rect 17082 8231 17094 8265
rect 17462 8231 17474 8265
rect 17082 8225 17474 8231
rect 17670 8265 18062 8271
rect 17670 8231 17682 8265
rect 18050 8231 18062 8265
rect 17670 8225 18062 8231
rect 18124 7968 18196 8312
rect 18258 8265 18650 8271
rect 18258 8231 18270 8265
rect 18638 8231 18650 8265
rect 18258 8225 18650 8231
rect 18846 8265 19238 8271
rect 18846 8231 18858 8265
rect 19226 8231 19238 8265
rect 18846 8225 19238 8231
rect 19300 7968 19372 8312
rect 19434 8265 19826 8271
rect 19434 8231 19446 8265
rect 19814 8231 19826 8265
rect 19434 8225 19826 8231
rect 20022 8265 20414 8271
rect 20022 8231 20034 8265
rect 20402 8231 20414 8265
rect 20022 8225 20414 8231
rect 20476 7968 20548 8312
rect 20610 8265 21002 8271
rect 20610 8231 20622 8265
rect 20990 8231 21002 8265
rect 20610 8225 21002 8231
rect 21198 8265 21590 8271
rect 21198 8231 21210 8265
rect 21578 8231 21590 8265
rect 21198 8225 21590 8231
rect 21652 7968 21724 8312
rect 21786 8265 22178 8271
rect 21786 8231 21798 8265
rect 22166 8231 22178 8265
rect 21786 8225 22178 8231
rect 22374 8265 22766 8271
rect 22374 8231 22386 8265
rect 22754 8231 22766 8265
rect 22374 8225 22766 8231
rect 22828 7968 22900 8312
rect 22962 8265 23354 8271
rect 22962 8231 22974 8265
rect 23342 8231 23354 8265
rect 22962 8225 23354 8231
rect 10998 7962 11210 7968
rect 10998 7852 11010 7962
rect 11198 7852 11210 7962
rect 10998 7846 11210 7852
rect 12174 7962 12386 7968
rect 12174 7852 12186 7962
rect 12374 7852 12386 7962
rect 12174 7846 12386 7852
rect 13350 7962 13562 7968
rect 13350 7852 13362 7962
rect 13550 7852 13562 7962
rect 13350 7846 13562 7852
rect 14526 7962 14738 7968
rect 14526 7852 14538 7962
rect 14726 7852 14738 7962
rect 14526 7846 14738 7852
rect 15702 7962 15914 7968
rect 15702 7852 15714 7962
rect 15902 7852 15914 7962
rect 15702 7846 15914 7852
rect 16878 7962 17090 7968
rect 16878 7852 16890 7962
rect 17078 7852 17090 7962
rect 16878 7846 17090 7852
rect 18054 7962 18266 7968
rect 18054 7852 18066 7962
rect 18254 7852 18266 7962
rect 18054 7846 18266 7852
rect 19230 7962 19442 7968
rect 19230 7852 19242 7962
rect 19430 7852 19442 7962
rect 19230 7846 19442 7852
rect 20406 7962 20618 7968
rect 20406 7852 20418 7962
rect 20606 7852 20618 7962
rect 20406 7846 20618 7852
rect 21582 7962 21794 7968
rect 21582 7852 21594 7962
rect 21782 7852 21794 7962
rect 21582 7846 21794 7852
rect 22758 7962 22970 7968
rect 22758 7852 22770 7962
rect 22958 7852 22970 7962
rect 22758 7846 22970 7852
rect 23416 7460 23488 8312
rect 23550 8265 23942 8271
rect 23550 8231 23562 8265
rect 23930 8231 23942 8265
rect 23550 8225 23942 8231
rect 24004 7968 24076 8312
rect 24138 8265 24530 8271
rect 24138 8231 24150 8265
rect 24518 8231 24530 8265
rect 24138 8225 24530 8231
rect 24726 8265 25118 8271
rect 24726 8231 24738 8265
rect 25106 8231 25118 8265
rect 24726 8225 25118 8231
rect 25180 7968 25252 8312
rect 25314 8265 25706 8271
rect 25314 8231 25326 8265
rect 25694 8231 25706 8265
rect 25314 8225 25706 8231
rect 23934 7962 24146 7968
rect 23934 7852 23946 7962
rect 24134 7852 24146 7962
rect 23934 7846 24146 7852
rect 25110 7962 25322 7968
rect 25110 7852 25122 7962
rect 25310 7852 25322 7962
rect 25110 7846 25322 7852
rect 25768 7460 25840 8312
rect 25902 8265 26294 8271
rect 25902 8231 25914 8265
rect 26282 8231 26294 8265
rect 25902 8225 26294 8231
rect 26356 7968 26428 8312
rect 26490 8265 26882 8271
rect 26490 8231 26502 8265
rect 26870 8231 26882 8265
rect 26490 8225 26882 8231
rect 27078 8265 27470 8271
rect 27078 8231 27090 8265
rect 27458 8231 27470 8265
rect 27078 8225 27470 8231
rect 27532 7968 27604 8312
rect 27666 8265 28058 8271
rect 27666 8231 27678 8265
rect 28046 8231 28058 8265
rect 27666 8225 28058 8231
rect 28254 8265 28646 8271
rect 28254 8231 28266 8265
rect 28634 8231 28646 8265
rect 28254 8225 28646 8231
rect 28708 7968 28780 8312
rect 28842 8265 29234 8271
rect 28842 8231 28854 8265
rect 29222 8231 29234 8265
rect 28842 8225 29234 8231
rect 29430 8265 29822 8271
rect 29430 8231 29442 8265
rect 29810 8231 29822 8265
rect 29430 8225 29822 8231
rect 29884 7978 29956 8312
rect 30018 8265 30410 8271
rect 30018 8231 30030 8265
rect 30398 8231 30410 8265
rect 30018 8225 30410 8231
rect 30606 8265 30998 8271
rect 30606 8231 30618 8265
rect 30986 8231 30998 8265
rect 30606 8225 30998 8231
rect 29814 7972 30026 7978
rect 26286 7962 26498 7968
rect 26286 7852 26298 7962
rect 26486 7852 26498 7962
rect 26286 7846 26498 7852
rect 27462 7962 27674 7968
rect 27462 7852 27474 7962
rect 27662 7852 27674 7962
rect 27462 7846 27674 7852
rect 28638 7962 28850 7968
rect 28638 7852 28650 7962
rect 28838 7852 28850 7962
rect 29814 7862 29826 7972
rect 30014 7862 30026 7972
rect 31060 7968 31132 8312
rect 31194 8265 31586 8271
rect 31194 8231 31206 8265
rect 31574 8231 31586 8265
rect 31194 8225 31586 8231
rect 31782 8265 32174 8271
rect 31782 8231 31794 8265
rect 32162 8231 32174 8265
rect 31782 8225 32174 8231
rect 32236 7968 32308 8312
rect 32370 8265 32762 8271
rect 32370 8231 32382 8265
rect 32750 8231 32762 8265
rect 32370 8225 32762 8231
rect 32958 8265 33350 8271
rect 32958 8231 32970 8265
rect 33338 8231 33350 8265
rect 32958 8225 33350 8231
rect 33412 7968 33484 8312
rect 33546 8265 33938 8271
rect 33546 8231 33558 8265
rect 33926 8231 33938 8265
rect 33546 8225 33938 8231
rect 34134 8265 34526 8271
rect 34134 8231 34146 8265
rect 34514 8231 34526 8265
rect 34134 8225 34526 8231
rect 34588 7978 34660 8312
rect 34722 8265 35114 8271
rect 34722 8231 34734 8265
rect 35102 8231 35114 8265
rect 34722 8225 35114 8231
rect 35310 8265 35702 8271
rect 35310 8231 35322 8265
rect 35690 8231 35702 8265
rect 35310 8225 35702 8231
rect 34504 7972 34740 7978
rect 29814 7856 30026 7862
rect 30990 7962 31202 7968
rect 28638 7846 28850 7852
rect 30990 7852 31002 7962
rect 31190 7852 31202 7962
rect 30990 7846 31202 7852
rect 32166 7962 32378 7968
rect 32166 7852 32178 7962
rect 32366 7852 32378 7962
rect 32166 7846 32378 7852
rect 33342 7962 33554 7968
rect 33342 7852 33354 7962
rect 33542 7852 33554 7962
rect 33342 7846 33554 7852
rect 34504 7850 34516 7972
rect 34728 7850 34740 7972
rect 35764 7968 35836 8312
rect 35898 8265 36290 8271
rect 35898 8231 35910 8265
rect 36278 8231 36290 8265
rect 35898 8225 36290 8231
rect 36486 8265 36878 8271
rect 36486 8231 36498 8265
rect 36866 8231 36878 8265
rect 36486 8225 36878 8231
rect 36940 7968 37012 8312
rect 37074 8265 37466 8271
rect 37074 8231 37086 8265
rect 37454 8231 37466 8265
rect 37074 8225 37466 8231
rect 37662 8265 38054 8271
rect 37662 8231 37674 8265
rect 38042 8231 38054 8265
rect 37662 8225 38054 8231
rect 38116 7968 38188 8312
rect 38250 8265 38642 8271
rect 38250 8231 38262 8265
rect 38630 8231 38642 8265
rect 38250 8225 38642 8231
rect 34504 7844 34740 7850
rect 35694 7962 35906 7968
rect 35694 7852 35706 7962
rect 35894 7852 35906 7962
rect 35694 7846 35906 7852
rect 36870 7962 37082 7968
rect 36870 7852 36882 7962
rect 37070 7852 37082 7962
rect 36870 7846 37082 7852
rect 38046 7962 38258 7968
rect 38046 7852 38058 7962
rect 38246 7852 38258 7962
rect 38046 7846 38258 7852
rect 23416 7380 25840 7460
rect 23524 6666 23604 7380
rect 23660 6836 23734 6842
rect 23660 6704 23670 6836
rect 23724 6704 23734 6836
rect 23660 6698 23734 6704
rect 23926 6836 24000 6842
rect 23926 6704 23936 6836
rect 23990 6704 24000 6836
rect 23926 6698 24000 6704
rect 24056 6666 24136 7380
rect 24192 6836 24266 6842
rect 24192 6704 24202 6836
rect 24256 6704 24266 6836
rect 24192 6698 24266 6704
rect 24458 6836 24532 6842
rect 24458 6704 24468 6836
rect 24522 6704 24532 6836
rect 24458 6698 24532 6704
rect 24588 6666 24668 7380
rect 24724 6836 24798 6842
rect 24724 6704 24734 6836
rect 24788 6704 24798 6836
rect 24724 6698 24798 6704
rect 24990 6836 25064 6842
rect 24990 6704 25000 6836
rect 25054 6704 25064 6836
rect 24990 6698 25064 6704
rect 25120 6666 25200 7380
rect 25256 6836 25330 6842
rect 25256 6704 25266 6836
rect 25320 6704 25330 6836
rect 25256 6698 25330 6704
rect 25522 6836 25596 6842
rect 25522 6704 25532 6836
rect 25586 6704 25596 6836
rect 25522 6698 25596 6704
rect 25652 6666 25732 7380
rect 23524 6654 23656 6666
rect 23524 5878 23616 6654
rect 23650 5878 23656 6654
rect 23524 5866 23656 5878
rect 23738 6654 23922 6666
rect 23738 5878 23744 6654
rect 23778 5878 23882 6654
rect 23916 5878 23922 6654
rect 23738 5866 23922 5878
rect 24004 6654 24188 6666
rect 24004 5878 24010 6654
rect 24044 5878 24148 6654
rect 24182 5878 24188 6654
rect 24004 5866 24188 5878
rect 24270 6654 24454 6666
rect 24270 5878 24276 6654
rect 24310 5878 24414 6654
rect 24448 5878 24454 6654
rect 24270 5866 24454 5878
rect 24536 6654 24720 6666
rect 24536 5878 24542 6654
rect 24576 5878 24680 6654
rect 24714 5878 24720 6654
rect 24536 5866 24720 5878
rect 24802 6654 24986 6666
rect 24802 5878 24808 6654
rect 24842 5878 24946 6654
rect 24980 5878 24986 6654
rect 24802 5866 24986 5878
rect 25068 6654 25252 6666
rect 25068 5878 25074 6654
rect 25108 5878 25212 6654
rect 25246 5878 25252 6654
rect 25068 5866 25252 5878
rect 25334 6654 25518 6666
rect 25334 5878 25340 6654
rect 25374 5878 25478 6654
rect 25512 5878 25518 6654
rect 25334 5866 25518 5878
rect 25600 6654 25732 6666
rect 25600 5878 25606 6654
rect 25640 5878 25732 6654
rect 25600 5866 25732 5878
rect 23524 5656 23610 5866
rect 23660 5826 23734 5832
rect 23660 5694 23670 5826
rect 23724 5694 23734 5826
rect 23660 5688 23734 5694
rect 23784 5656 23876 5866
rect 23926 5826 24000 5832
rect 23926 5694 23936 5826
rect 23990 5694 24000 5826
rect 23926 5688 24000 5694
rect 24050 5656 24142 5866
rect 24192 5826 24266 5832
rect 24192 5694 24202 5826
rect 24256 5694 24266 5826
rect 24192 5688 24266 5694
rect 24316 5656 24408 5866
rect 24458 5826 24532 5832
rect 24458 5694 24468 5826
rect 24522 5694 24532 5826
rect 24458 5688 24532 5694
rect 24582 5656 24674 5866
rect 24724 5826 24798 5832
rect 24724 5694 24734 5826
rect 24788 5694 24798 5826
rect 24724 5688 24798 5694
rect 24848 5656 24940 5866
rect 24990 5826 25064 5832
rect 24990 5694 25000 5826
rect 25054 5694 25064 5826
rect 24990 5688 25064 5694
rect 25114 5656 25206 5866
rect 25256 5826 25330 5832
rect 25256 5694 25266 5826
rect 25320 5694 25330 5826
rect 25256 5688 25330 5694
rect 25380 5656 25472 5866
rect 25522 5826 25596 5832
rect 25522 5694 25532 5826
rect 25586 5694 25596 5826
rect 25522 5688 25596 5694
rect 25646 5656 25732 5866
rect 23524 5644 23656 5656
rect 23524 4868 23616 5644
rect 23650 4868 23656 5644
rect 23524 4856 23656 4868
rect 23738 5644 23922 5656
rect 23738 4868 23744 5644
rect 23778 4868 23882 5644
rect 23916 4868 23922 5644
rect 23738 4856 23922 4868
rect 24004 5644 24188 5656
rect 24004 4868 24010 5644
rect 24044 4868 24148 5644
rect 24182 4868 24188 5644
rect 24004 4856 24188 4868
rect 24270 5644 24454 5656
rect 24270 4868 24276 5644
rect 24310 4868 24414 5644
rect 24448 4868 24454 5644
rect 24270 4856 24454 4868
rect 24536 5644 24720 5656
rect 24536 4868 24542 5644
rect 24576 4868 24680 5644
rect 24714 4868 24720 5644
rect 24536 4856 24720 4868
rect 24802 5644 24986 5656
rect 24802 4868 24808 5644
rect 24842 4868 24946 5644
rect 24980 4868 24986 5644
rect 24802 4856 24986 4868
rect 25068 5644 25252 5656
rect 25068 4868 25074 5644
rect 25108 4868 25212 5644
rect 25246 4868 25252 5644
rect 25068 4856 25252 4868
rect 25334 5644 25518 5656
rect 25334 4868 25340 5644
rect 25374 4868 25478 5644
rect 25512 4868 25518 5644
rect 25334 4856 25518 4868
rect 25600 5644 25732 5656
rect 25600 4868 25606 5644
rect 25640 4868 25732 5644
rect 25600 4856 25732 4868
rect 23524 4646 23610 4856
rect 23660 4816 23734 4822
rect 23660 4684 23670 4816
rect 23724 4684 23734 4816
rect 23660 4678 23734 4684
rect 23784 4646 23876 4856
rect 23926 4816 24000 4822
rect 23926 4684 23936 4816
rect 23990 4684 24000 4816
rect 23926 4678 24000 4684
rect 24050 4646 24142 4856
rect 24192 4816 24266 4822
rect 24192 4684 24202 4816
rect 24256 4684 24266 4816
rect 24192 4678 24266 4684
rect 24316 4646 24408 4856
rect 24458 4816 24532 4822
rect 24458 4684 24468 4816
rect 24522 4684 24532 4816
rect 24458 4678 24532 4684
rect 24582 4646 24674 4856
rect 24724 4816 24798 4822
rect 24724 4684 24734 4816
rect 24788 4684 24798 4816
rect 24724 4678 24798 4684
rect 24848 4646 24940 4856
rect 24990 4816 25064 4822
rect 24990 4684 25000 4816
rect 25054 4684 25064 4816
rect 24990 4678 25064 4684
rect 25114 4646 25206 4856
rect 25256 4816 25330 4822
rect 25256 4684 25266 4816
rect 25320 4684 25330 4816
rect 25256 4678 25330 4684
rect 25380 4646 25472 4856
rect 25522 4816 25596 4822
rect 25522 4684 25532 4816
rect 25586 4684 25596 4816
rect 25522 4678 25596 4684
rect 25646 4646 25732 4856
rect 30570 4802 30580 5340
rect 31062 4802 31072 5340
rect 30791 4744 30797 4802
rect 30835 4744 30841 4802
rect 30791 4732 30841 4744
rect 23524 4634 23656 4646
rect 23524 3858 23616 4634
rect 23650 3858 23656 4634
rect 23524 3846 23656 3858
rect 23738 4634 23922 4646
rect 23738 3858 23744 4634
rect 23778 3858 23882 4634
rect 23916 3858 23922 4634
rect 23738 3846 23922 3858
rect 24004 4634 24188 4646
rect 24004 3858 24010 4634
rect 24044 3858 24148 4634
rect 24182 3858 24188 4634
rect 24004 3846 24188 3858
rect 24270 4634 24454 4646
rect 24270 3858 24276 4634
rect 24310 3858 24414 4634
rect 24448 3858 24454 4634
rect 24270 3846 24454 3858
rect 24536 4634 24720 4646
rect 24536 3858 24542 4634
rect 24576 3858 24680 4634
rect 24714 3858 24720 4634
rect 24536 3846 24720 3858
rect 24802 4634 24986 4646
rect 24802 3858 24808 4634
rect 24842 3858 24946 4634
rect 24980 3858 24986 4634
rect 24802 3846 24986 3858
rect 25068 4634 25252 4646
rect 25068 3858 25074 4634
rect 25108 3858 25212 4634
rect 25246 3858 25252 4634
rect 25068 3846 25252 3858
rect 25334 4634 25518 4646
rect 25334 3858 25340 4634
rect 25374 3858 25478 4634
rect 25512 3858 25518 4634
rect 25334 3846 25518 3858
rect 25600 4634 25732 4646
rect 25600 3858 25606 4634
rect 25640 3858 25732 4634
rect 31070 4534 31244 4554
rect 25600 3846 25732 3858
rect 30791 4150 30841 4162
rect 23660 3806 23734 3812
rect 23660 3674 23670 3806
rect 23724 3674 23734 3806
rect 23660 3668 23734 3674
rect 23790 2474 23870 3846
rect 23926 3806 24000 3812
rect 23926 3674 23936 3806
rect 23990 3674 24000 3806
rect 23926 3668 24000 3674
rect 24192 3806 24266 3812
rect 24192 3674 24202 3806
rect 24256 3674 24266 3806
rect 24192 3668 24266 3674
rect 24322 3290 24402 3846
rect 24458 3806 24532 3812
rect 24458 3674 24468 3806
rect 24522 3674 24532 3806
rect 24458 3668 24532 3674
rect 24724 3806 24798 3812
rect 24724 3674 24734 3806
rect 24788 3674 24798 3806
rect 24724 3668 24798 3674
rect 24854 3290 24934 3846
rect 24990 3806 25064 3812
rect 24990 3674 25000 3806
rect 25054 3674 25064 3806
rect 24990 3668 25064 3674
rect 25256 3806 25330 3812
rect 25256 3674 25266 3806
rect 25320 3674 25330 3806
rect 25256 3668 25330 3674
rect 24322 3258 24934 3290
rect 24322 3130 24368 3258
rect 24862 3130 24934 3258
rect 24322 3100 24934 3130
rect 24234 2638 24544 2644
rect 24234 2512 24250 2638
rect 24288 2512 24490 2638
rect 24528 2512 24544 2638
rect 24234 2506 24304 2512
rect 24474 2506 24544 2512
rect 24602 2474 24656 3100
rect 24714 2638 25024 2644
rect 24714 2512 24730 2638
rect 24768 2512 24970 2638
rect 25008 2512 25024 2638
rect 24714 2506 24784 2512
rect 24954 2506 25024 2512
rect 25386 2474 25466 3846
rect 25522 3806 25596 3812
rect 25522 3674 25532 3806
rect 25586 3674 25596 3806
rect 30791 3766 30797 4150
rect 25522 3668 25596 3674
rect 30780 3753 30797 3766
rect 30835 3766 30841 4150
rect 31070 4074 31086 4534
rect 31226 4074 31244 4534
rect 30835 3753 30852 3766
rect 30780 3348 30852 3753
rect 30566 2918 30576 3348
rect 30952 2918 30962 3348
rect 23790 2462 24228 2474
rect 23790 2404 24188 2462
rect 24138 1886 24188 2404
rect 24222 1886 24228 2462
rect 24138 1874 24228 1886
rect 24310 2462 24468 2474
rect 24310 1886 24316 2462
rect 24350 1886 24428 2462
rect 24462 1886 24468 2462
rect 24310 1874 24468 1886
rect 24550 2462 24708 2474
rect 24550 1886 24556 2462
rect 24590 1886 24668 2462
rect 24702 1886 24708 2462
rect 24550 1874 24708 1886
rect 24790 2462 24948 2474
rect 24790 1886 24796 2462
rect 24830 1886 24908 2462
rect 24942 1886 24948 2462
rect 24790 1874 24948 1886
rect 25030 2462 25466 2474
rect 25030 1886 25036 2462
rect 25070 2404 25466 2462
rect 25070 1886 25126 2404
rect 25030 1874 25126 1886
rect 24138 1666 24188 1874
rect 24234 1836 24304 1842
rect 24234 1704 24250 1836
rect 24288 1704 24304 1836
rect 24234 1698 24304 1704
rect 24356 1666 24422 1874
rect 24474 1836 24544 1842
rect 24474 1704 24490 1836
rect 24528 1704 24544 1836
rect 24474 1698 24544 1704
rect 24596 1666 24662 1874
rect 24714 1836 24784 1842
rect 24714 1704 24730 1836
rect 24768 1704 24784 1836
rect 24714 1698 24784 1704
rect 24836 1666 24902 1874
rect 24954 1836 25024 1842
rect 24954 1704 24970 1836
rect 25008 1704 25024 1836
rect 24954 1698 25024 1704
rect 25076 1666 25126 1874
rect 24138 1654 24228 1666
rect 24138 1078 24188 1654
rect 24222 1078 24228 1654
rect 24138 1066 24228 1078
rect 24310 1654 24468 1666
rect 24310 1078 24316 1654
rect 24350 1078 24428 1654
rect 24462 1078 24468 1654
rect 24310 1066 24468 1078
rect 24550 1654 24708 1666
rect 24550 1078 24556 1654
rect 24590 1078 24668 1654
rect 24702 1078 24708 1654
rect 24550 1066 24708 1078
rect 24790 1654 24948 1666
rect 24790 1078 24796 1654
rect 24830 1078 24908 1654
rect 24942 1078 24948 1654
rect 24790 1066 24948 1078
rect 25030 1654 25126 1666
rect 25030 1078 25036 1654
rect 25070 1078 25126 1654
rect 31070 1224 31244 4074
rect 25030 1066 25126 1078
rect 24234 1028 24304 1034
rect 24234 896 24250 1028
rect 24288 896 24304 1028
rect 24234 890 24304 896
rect 24362 650 24416 1066
rect 24474 1028 24544 1034
rect 24474 896 24490 1028
rect 24528 896 24544 1028
rect 24474 890 24544 896
rect 24714 1028 24784 1034
rect 24714 896 24730 1028
rect 24768 896 24784 1028
rect 24714 890 24784 896
rect 24842 650 24896 1066
rect 24954 1028 25024 1034
rect 24954 896 24970 1028
rect 25008 896 25024 1028
rect 24954 890 25024 896
rect 23928 644 25304 650
rect 23928 532 23940 644
rect 25292 532 25304 644
rect 30782 558 30792 1224
rect 31548 558 31558 1224
rect 23928 526 25304 532
<< via1 >>
rect 20014 15572 20124 15644
rect 20494 15572 20604 15644
rect 20974 15572 21084 15644
rect 21454 15572 21564 15644
rect 21934 15572 22044 15644
rect 22414 15572 22524 15644
rect 22894 15572 23004 15644
rect 23374 15572 23484 15644
rect 23854 15572 23964 15644
rect 24334 15572 24444 15644
rect 24814 15572 24924 15644
rect 25294 15572 25404 15644
rect 25774 15572 25884 15644
rect 26254 15572 26364 15644
rect 26734 15572 26844 15644
rect 27214 15572 27324 15644
rect 27694 15572 27804 15644
rect 28174 15572 28284 15644
rect 28654 15572 28764 15644
rect 29134 15572 29244 15644
rect 19914 15168 19930 15300
rect 19930 15168 19968 15300
rect 19968 15168 19984 15300
rect 20154 15168 20170 15300
rect 20170 15168 20208 15300
rect 20208 15168 20224 15300
rect 20394 15168 20410 15300
rect 20410 15168 20448 15300
rect 20448 15168 20464 15300
rect 20634 15168 20650 15300
rect 20650 15168 20688 15300
rect 20688 15168 20704 15300
rect 20874 15168 20890 15300
rect 20890 15168 20928 15300
rect 20928 15168 20944 15300
rect 21114 15168 21130 15300
rect 21130 15168 21168 15300
rect 21168 15168 21184 15300
rect 21354 15168 21370 15300
rect 21370 15168 21408 15300
rect 21408 15168 21424 15300
rect 21594 15168 21610 15300
rect 21610 15168 21648 15300
rect 21648 15168 21664 15300
rect 21834 15168 21850 15300
rect 21850 15168 21888 15300
rect 21888 15168 21904 15300
rect 22074 15168 22090 15300
rect 22090 15168 22128 15300
rect 22128 15168 22144 15300
rect 22314 15168 22330 15300
rect 22330 15168 22368 15300
rect 22368 15168 22384 15300
rect 22554 15168 22570 15300
rect 22570 15168 22608 15300
rect 22608 15168 22624 15300
rect 22794 15168 22810 15300
rect 22810 15168 22848 15300
rect 22848 15168 22864 15300
rect 23034 15168 23050 15300
rect 23050 15168 23088 15300
rect 23088 15168 23104 15300
rect 23274 15168 23290 15300
rect 23290 15168 23328 15300
rect 23328 15168 23344 15300
rect 23514 15168 23530 15300
rect 23530 15168 23568 15300
rect 23568 15168 23584 15300
rect 23754 15168 23770 15300
rect 23770 15168 23808 15300
rect 23808 15168 23824 15300
rect 23994 15168 24010 15300
rect 24010 15168 24048 15300
rect 24048 15168 24064 15300
rect 24234 15168 24250 15300
rect 24250 15168 24288 15300
rect 24288 15168 24304 15300
rect 24474 15168 24490 15300
rect 24490 15168 24528 15300
rect 24528 15168 24544 15300
rect 24714 15168 24730 15300
rect 24730 15168 24768 15300
rect 24768 15168 24784 15300
rect 24954 15168 24970 15300
rect 24970 15168 25008 15300
rect 25008 15168 25024 15300
rect 25194 15168 25210 15300
rect 25210 15168 25248 15300
rect 25248 15168 25264 15300
rect 25434 15168 25450 15300
rect 25450 15168 25488 15300
rect 25488 15168 25504 15300
rect 25674 15168 25690 15300
rect 25690 15168 25728 15300
rect 25728 15168 25744 15300
rect 25914 15168 25930 15300
rect 25930 15168 25968 15300
rect 25968 15168 25984 15300
rect 26154 15168 26170 15300
rect 26170 15168 26208 15300
rect 26208 15168 26224 15300
rect 26394 15168 26410 15300
rect 26410 15168 26448 15300
rect 26448 15168 26464 15300
rect 26634 15168 26650 15300
rect 26650 15168 26688 15300
rect 26688 15168 26704 15300
rect 26874 15168 26890 15300
rect 26890 15168 26928 15300
rect 26928 15168 26944 15300
rect 27114 15168 27130 15300
rect 27130 15168 27168 15300
rect 27168 15168 27184 15300
rect 27354 15168 27370 15300
rect 27370 15168 27408 15300
rect 27408 15168 27424 15300
rect 27594 15168 27610 15300
rect 27610 15168 27648 15300
rect 27648 15168 27664 15300
rect 27834 15168 27850 15300
rect 27850 15168 27888 15300
rect 27888 15168 27904 15300
rect 28074 15168 28090 15300
rect 28090 15168 28128 15300
rect 28128 15168 28144 15300
rect 28314 15168 28330 15300
rect 28330 15168 28368 15300
rect 28368 15168 28384 15300
rect 28554 15168 28570 15300
rect 28570 15168 28608 15300
rect 28608 15168 28624 15300
rect 28794 15168 28810 15300
rect 28810 15168 28848 15300
rect 28848 15168 28864 15300
rect 29034 15168 29050 15300
rect 29050 15168 29088 15300
rect 29088 15168 29104 15300
rect 29274 15168 29290 15300
rect 29290 15168 29328 15300
rect 29328 15168 29344 15300
rect 19914 14360 19930 14492
rect 19930 14360 19968 14492
rect 19968 14360 19984 14492
rect 20154 14360 20170 14492
rect 20170 14360 20208 14492
rect 20208 14360 20224 14492
rect 20394 14360 20410 14492
rect 20410 14360 20448 14492
rect 20448 14360 20464 14492
rect 20634 14360 20650 14492
rect 20650 14360 20688 14492
rect 20688 14360 20704 14492
rect 20874 14360 20890 14492
rect 20890 14360 20928 14492
rect 20928 14360 20944 14492
rect 21114 14360 21130 14492
rect 21130 14360 21168 14492
rect 21168 14360 21184 14492
rect 21354 14360 21370 14492
rect 21370 14360 21408 14492
rect 21408 14360 21424 14492
rect 21594 14360 21610 14492
rect 21610 14360 21648 14492
rect 21648 14360 21664 14492
rect 21834 14360 21850 14492
rect 21850 14360 21888 14492
rect 21888 14360 21904 14492
rect 22074 14360 22090 14492
rect 22090 14360 22128 14492
rect 22128 14360 22144 14492
rect 22314 14360 22330 14492
rect 22330 14360 22368 14492
rect 22368 14360 22384 14492
rect 22554 14360 22570 14492
rect 22570 14360 22608 14492
rect 22608 14360 22624 14492
rect 22794 14360 22810 14492
rect 22810 14360 22848 14492
rect 22848 14360 22864 14492
rect 23034 14360 23050 14492
rect 23050 14360 23088 14492
rect 23088 14360 23104 14492
rect 23274 14360 23290 14492
rect 23290 14360 23328 14492
rect 23328 14360 23344 14492
rect 23514 14360 23530 14492
rect 23530 14360 23568 14492
rect 23568 14360 23584 14492
rect 23754 14360 23770 14492
rect 23770 14360 23808 14492
rect 23808 14360 23824 14492
rect 23994 14360 24010 14492
rect 24010 14360 24048 14492
rect 24048 14360 24064 14492
rect 24234 14360 24250 14492
rect 24250 14360 24288 14492
rect 24288 14360 24304 14492
rect 24474 14360 24490 14492
rect 24490 14360 24528 14492
rect 24528 14360 24544 14492
rect 24714 14360 24730 14492
rect 24730 14360 24768 14492
rect 24768 14360 24784 14492
rect 24954 14360 24970 14492
rect 24970 14360 25008 14492
rect 25008 14360 25024 14492
rect 25194 14360 25210 14492
rect 25210 14360 25248 14492
rect 25248 14360 25264 14492
rect 25434 14360 25450 14492
rect 25450 14360 25488 14492
rect 25488 14360 25504 14492
rect 25674 14360 25690 14492
rect 25690 14360 25728 14492
rect 25728 14360 25744 14492
rect 25914 14360 25930 14492
rect 25930 14360 25968 14492
rect 25968 14360 25984 14492
rect 26154 14360 26170 14492
rect 26170 14360 26208 14492
rect 26208 14360 26224 14492
rect 26394 14360 26410 14492
rect 26410 14360 26448 14492
rect 26448 14360 26464 14492
rect 26634 14360 26650 14492
rect 26650 14360 26688 14492
rect 26688 14360 26704 14492
rect 26874 14360 26890 14492
rect 26890 14360 26928 14492
rect 26928 14360 26944 14492
rect 27114 14360 27130 14492
rect 27130 14360 27168 14492
rect 27168 14360 27184 14492
rect 27354 14360 27370 14492
rect 27370 14360 27408 14492
rect 27408 14360 27424 14492
rect 27594 14360 27610 14492
rect 27610 14360 27648 14492
rect 27648 14360 27664 14492
rect 27834 14360 27850 14492
rect 27850 14360 27888 14492
rect 27888 14360 27904 14492
rect 28074 14360 28090 14492
rect 28090 14360 28128 14492
rect 28128 14360 28144 14492
rect 28314 14360 28330 14492
rect 28330 14360 28368 14492
rect 28368 14360 28384 14492
rect 28554 14360 28570 14492
rect 28570 14360 28608 14492
rect 28608 14360 28624 14492
rect 28794 14360 28810 14492
rect 28810 14360 28848 14492
rect 28848 14360 28864 14492
rect 29034 14360 29050 14492
rect 29050 14360 29088 14492
rect 29088 14360 29104 14492
rect 29274 14360 29290 14492
rect 29290 14360 29328 14492
rect 29328 14360 29344 14492
rect 19914 13552 19930 13684
rect 19930 13552 19968 13684
rect 19968 13552 19984 13684
rect 20154 13552 20170 13684
rect 20170 13552 20208 13684
rect 20208 13552 20224 13684
rect 20394 13552 20410 13684
rect 20410 13552 20448 13684
rect 20448 13552 20464 13684
rect 20634 13552 20650 13684
rect 20650 13552 20688 13684
rect 20688 13552 20704 13684
rect 20874 13552 20890 13684
rect 20890 13552 20928 13684
rect 20928 13552 20944 13684
rect 21114 13552 21130 13684
rect 21130 13552 21168 13684
rect 21168 13552 21184 13684
rect 21354 13552 21370 13684
rect 21370 13552 21408 13684
rect 21408 13552 21424 13684
rect 21594 13552 21610 13684
rect 21610 13552 21648 13684
rect 21648 13552 21664 13684
rect 21834 13552 21850 13684
rect 21850 13552 21888 13684
rect 21888 13552 21904 13684
rect 22074 13552 22090 13684
rect 22090 13552 22128 13684
rect 22128 13552 22144 13684
rect 22314 13552 22330 13684
rect 22330 13552 22368 13684
rect 22368 13552 22384 13684
rect 22554 13552 22570 13684
rect 22570 13552 22608 13684
rect 22608 13552 22624 13684
rect 22794 13552 22810 13684
rect 22810 13552 22848 13684
rect 22848 13552 22864 13684
rect 23034 13552 23050 13684
rect 23050 13552 23088 13684
rect 23088 13552 23104 13684
rect 23274 13552 23290 13684
rect 23290 13552 23328 13684
rect 23328 13552 23344 13684
rect 23514 13552 23530 13684
rect 23530 13552 23568 13684
rect 23568 13552 23584 13684
rect 23754 13552 23770 13684
rect 23770 13552 23808 13684
rect 23808 13552 23824 13684
rect 23994 13552 24010 13684
rect 24010 13552 24048 13684
rect 24048 13552 24064 13684
rect 24234 13552 24250 13684
rect 24250 13552 24288 13684
rect 24288 13552 24304 13684
rect 24474 13552 24490 13684
rect 24490 13552 24528 13684
rect 24528 13552 24544 13684
rect 24714 13552 24730 13684
rect 24730 13552 24768 13684
rect 24768 13552 24784 13684
rect 24954 13552 24970 13684
rect 24970 13552 25008 13684
rect 25008 13552 25024 13684
rect 25194 13552 25210 13684
rect 25210 13552 25248 13684
rect 25248 13552 25264 13684
rect 25434 13552 25450 13684
rect 25450 13552 25488 13684
rect 25488 13552 25504 13684
rect 25674 13552 25690 13684
rect 25690 13552 25728 13684
rect 25728 13552 25744 13684
rect 25914 13552 25930 13684
rect 25930 13552 25968 13684
rect 25968 13552 25984 13684
rect 26154 13552 26170 13684
rect 26170 13552 26208 13684
rect 26208 13552 26224 13684
rect 26394 13552 26410 13684
rect 26410 13552 26448 13684
rect 26448 13552 26464 13684
rect 26634 13552 26650 13684
rect 26650 13552 26688 13684
rect 26688 13552 26704 13684
rect 26874 13552 26890 13684
rect 26890 13552 26928 13684
rect 26928 13552 26944 13684
rect 27114 13552 27130 13684
rect 27130 13552 27168 13684
rect 27168 13552 27184 13684
rect 27354 13552 27370 13684
rect 27370 13552 27408 13684
rect 27408 13552 27424 13684
rect 27594 13552 27610 13684
rect 27610 13552 27648 13684
rect 27648 13552 27664 13684
rect 27834 13552 27850 13684
rect 27850 13552 27888 13684
rect 27888 13552 27904 13684
rect 28074 13552 28090 13684
rect 28090 13552 28128 13684
rect 28128 13552 28144 13684
rect 28314 13552 28330 13684
rect 28330 13552 28368 13684
rect 28368 13552 28384 13684
rect 28554 13552 28570 13684
rect 28570 13552 28608 13684
rect 28608 13552 28624 13684
rect 28794 13552 28810 13684
rect 28810 13552 28848 13684
rect 28848 13552 28864 13684
rect 29034 13552 29050 13684
rect 29050 13552 29088 13684
rect 29088 13552 29104 13684
rect 29274 13552 29290 13684
rect 29290 13552 29328 13684
rect 29328 13552 29344 13684
rect 33856 12216 34756 12658
rect 11010 7852 11198 7962
rect 12186 7852 12374 7962
rect 13362 7852 13550 7962
rect 14538 7852 14726 7962
rect 15714 7852 15902 7962
rect 16890 7852 17078 7962
rect 18066 7852 18254 7962
rect 19242 7852 19430 7962
rect 20418 7852 20606 7962
rect 21594 7852 21782 7962
rect 22770 7852 22958 7962
rect 23946 7852 24134 7962
rect 25122 7852 25310 7962
rect 26298 7852 26486 7962
rect 27474 7852 27662 7962
rect 28650 7852 28838 7962
rect 31002 7852 31190 7962
rect 32178 7852 32366 7962
rect 33354 7852 33542 7962
rect 35706 7852 35894 7962
rect 36882 7852 37070 7962
rect 38058 7852 38246 7962
rect 23670 6704 23678 6836
rect 23678 6704 23716 6836
rect 23716 6704 23724 6836
rect 23936 6704 23944 6836
rect 23944 6704 23982 6836
rect 23982 6704 23990 6836
rect 24202 6704 24210 6836
rect 24210 6704 24248 6836
rect 24248 6704 24256 6836
rect 24468 6704 24476 6836
rect 24476 6704 24514 6836
rect 24514 6704 24522 6836
rect 24734 6704 24742 6836
rect 24742 6704 24780 6836
rect 24780 6704 24788 6836
rect 25000 6704 25008 6836
rect 25008 6704 25046 6836
rect 25046 6704 25054 6836
rect 25266 6704 25274 6836
rect 25274 6704 25312 6836
rect 25312 6704 25320 6836
rect 25532 6704 25540 6836
rect 25540 6704 25578 6836
rect 25578 6704 25586 6836
rect 23670 5694 23678 5826
rect 23678 5694 23716 5826
rect 23716 5694 23724 5826
rect 23936 5694 23944 5826
rect 23944 5694 23982 5826
rect 23982 5694 23990 5826
rect 24202 5694 24210 5826
rect 24210 5694 24248 5826
rect 24248 5694 24256 5826
rect 24468 5694 24476 5826
rect 24476 5694 24514 5826
rect 24514 5694 24522 5826
rect 24734 5694 24742 5826
rect 24742 5694 24780 5826
rect 24780 5694 24788 5826
rect 25000 5694 25008 5826
rect 25008 5694 25046 5826
rect 25046 5694 25054 5826
rect 25266 5694 25274 5826
rect 25274 5694 25312 5826
rect 25312 5694 25320 5826
rect 25532 5694 25540 5826
rect 25540 5694 25578 5826
rect 25578 5694 25586 5826
rect 23670 4684 23678 4816
rect 23678 4684 23716 4816
rect 23716 4684 23724 4816
rect 23936 4684 23944 4816
rect 23944 4684 23982 4816
rect 23982 4684 23990 4816
rect 24202 4684 24210 4816
rect 24210 4684 24248 4816
rect 24248 4684 24256 4816
rect 24468 4684 24476 4816
rect 24476 4684 24514 4816
rect 24514 4684 24522 4816
rect 24734 4684 24742 4816
rect 24742 4684 24780 4816
rect 24780 4684 24788 4816
rect 25000 4684 25008 4816
rect 25008 4684 25046 4816
rect 25046 4684 25054 4816
rect 25266 4684 25274 4816
rect 25274 4684 25312 4816
rect 25312 4684 25320 4816
rect 25532 4684 25540 4816
rect 25540 4684 25578 4816
rect 25578 4684 25586 4816
rect 30580 5141 31062 5340
rect 30580 4802 30797 5141
rect 30797 4802 30835 5141
rect 30835 4802 31062 5141
rect 23670 3674 23678 3806
rect 23678 3674 23716 3806
rect 23716 3674 23724 3806
rect 23936 3674 23944 3806
rect 23944 3674 23982 3806
rect 23982 3674 23990 3806
rect 24202 3674 24210 3806
rect 24210 3674 24248 3806
rect 24248 3674 24256 3806
rect 24468 3674 24476 3806
rect 24476 3674 24514 3806
rect 24514 3674 24522 3806
rect 24734 3674 24742 3806
rect 24742 3674 24780 3806
rect 24780 3674 24788 3806
rect 25000 3674 25008 3806
rect 25008 3674 25046 3806
rect 25046 3674 25054 3806
rect 25266 3674 25274 3806
rect 25274 3674 25312 3806
rect 25312 3674 25320 3806
rect 24368 3130 24862 3258
rect 25532 3674 25540 3806
rect 25540 3674 25578 3806
rect 25578 3674 25586 3806
rect 30576 2918 30952 3348
rect 23940 532 25292 644
rect 30792 558 31548 1224
<< metal2 >>
rect 20014 15644 20124 15654
rect 20014 15562 20124 15572
rect 20494 15644 20604 15654
rect 20494 15562 20604 15572
rect 20974 15644 21084 15654
rect 20974 15562 21084 15572
rect 21454 15644 21564 15654
rect 21454 15562 21564 15572
rect 21934 15644 22044 15654
rect 21934 15562 22044 15572
rect 22414 15644 22524 15654
rect 22414 15562 22524 15572
rect 22894 15644 23004 15654
rect 22894 15562 23004 15572
rect 23374 15644 23484 15654
rect 23374 15562 23484 15572
rect 23854 15644 23964 15654
rect 23854 15562 23964 15572
rect 24334 15644 24444 15654
rect 24334 15562 24444 15572
rect 24814 15644 24924 15654
rect 24814 15562 24924 15572
rect 25294 15644 25404 15654
rect 25294 15562 25404 15572
rect 25774 15644 25884 15654
rect 25774 15562 25884 15572
rect 26254 15644 26364 15654
rect 26254 15562 26364 15572
rect 26734 15644 26844 15654
rect 26734 15562 26844 15572
rect 27214 15644 27324 15654
rect 27214 15562 27324 15572
rect 27694 15644 27804 15654
rect 27694 15562 27804 15572
rect 28174 15644 28284 15654
rect 28174 15562 28284 15572
rect 28654 15644 28764 15654
rect 28654 15562 28764 15572
rect 29134 15644 29244 15654
rect 29134 15562 29244 15572
rect 29952 15458 30252 15468
rect 19904 15300 29952 15310
rect 19904 15168 19914 15300
rect 19984 15168 20154 15300
rect 20224 15168 20394 15300
rect 20464 15168 20634 15300
rect 20704 15168 20874 15300
rect 20944 15168 21114 15300
rect 21184 15168 21354 15300
rect 21424 15168 21594 15300
rect 21664 15168 21834 15300
rect 21904 15168 22074 15300
rect 22144 15168 22314 15300
rect 22384 15168 22554 15300
rect 22624 15168 22794 15300
rect 22864 15168 23034 15300
rect 23104 15168 23274 15300
rect 23344 15168 23514 15300
rect 23584 15168 23754 15300
rect 23824 15168 23994 15300
rect 24064 15168 24234 15300
rect 24304 15168 24474 15300
rect 24544 15168 24714 15300
rect 24784 15168 24954 15300
rect 25024 15168 25194 15300
rect 25264 15168 25434 15300
rect 25504 15168 25674 15300
rect 25744 15168 25914 15300
rect 25984 15168 26154 15300
rect 26224 15168 26394 15300
rect 26464 15168 26634 15300
rect 26704 15168 26874 15300
rect 26944 15168 27114 15300
rect 27184 15168 27354 15300
rect 27424 15168 27594 15300
rect 27664 15168 27834 15300
rect 27904 15168 28074 15300
rect 28144 15168 28314 15300
rect 28384 15168 28554 15300
rect 28624 15168 28794 15300
rect 28864 15168 29034 15300
rect 29104 15168 29274 15300
rect 29344 15168 29952 15300
rect 19904 15158 29952 15168
rect 29952 15148 30252 15158
rect 29952 14650 30252 14660
rect 19904 14492 29952 14502
rect 19904 14360 19914 14492
rect 19984 14360 20154 14492
rect 20224 14360 20394 14492
rect 20464 14360 20634 14492
rect 20704 14360 20874 14492
rect 20944 14360 21114 14492
rect 21184 14360 21354 14492
rect 21424 14360 21594 14492
rect 21664 14360 21834 14492
rect 21904 14360 22074 14492
rect 22144 14360 22314 14492
rect 22384 14360 22554 14492
rect 22624 14360 22794 14492
rect 22864 14360 23034 14492
rect 23104 14360 23274 14492
rect 23344 14360 23514 14492
rect 23584 14360 23754 14492
rect 23824 14360 23994 14492
rect 24064 14360 24234 14492
rect 24304 14360 24474 14492
rect 24544 14360 24714 14492
rect 24784 14360 24954 14492
rect 25024 14360 25194 14492
rect 25264 14360 25434 14492
rect 25504 14360 25674 14492
rect 25744 14360 25914 14492
rect 25984 14360 26154 14492
rect 26224 14360 26394 14492
rect 26464 14360 26634 14492
rect 26704 14360 26874 14492
rect 26944 14360 27114 14492
rect 27184 14360 27354 14492
rect 27424 14360 27594 14492
rect 27664 14360 27834 14492
rect 27904 14360 28074 14492
rect 28144 14360 28314 14492
rect 28384 14360 28554 14492
rect 28624 14360 28794 14492
rect 28864 14360 29034 14492
rect 29104 14360 29274 14492
rect 29344 14360 29952 14492
rect 19904 14350 29952 14360
rect 29952 14340 30252 14350
rect 29952 13842 30252 13852
rect 19904 13684 29952 13694
rect 19904 13552 19914 13684
rect 19984 13552 20154 13684
rect 20224 13552 20394 13684
rect 20464 13552 20634 13684
rect 20704 13552 20874 13684
rect 20944 13552 21114 13684
rect 21184 13552 21354 13684
rect 21424 13552 21594 13684
rect 21664 13552 21834 13684
rect 21904 13552 22074 13684
rect 22144 13552 22314 13684
rect 22384 13552 22554 13684
rect 22624 13552 22794 13684
rect 22864 13552 23034 13684
rect 23104 13552 23274 13684
rect 23344 13552 23514 13684
rect 23584 13552 23754 13684
rect 23824 13552 23994 13684
rect 24064 13552 24234 13684
rect 24304 13552 24474 13684
rect 24544 13552 24714 13684
rect 24784 13552 24954 13684
rect 25024 13552 25194 13684
rect 25264 13552 25434 13684
rect 25504 13552 25674 13684
rect 25744 13552 25914 13684
rect 25984 13552 26154 13684
rect 26224 13552 26394 13684
rect 26464 13552 26634 13684
rect 26704 13552 26874 13684
rect 26944 13552 27114 13684
rect 27184 13552 27354 13684
rect 27424 13552 27594 13684
rect 27664 13552 27834 13684
rect 27904 13552 28074 13684
rect 28144 13552 28314 13684
rect 28384 13552 28554 13684
rect 28624 13552 28794 13684
rect 28864 13552 29034 13684
rect 29104 13552 29274 13684
rect 29344 13552 29952 13684
rect 19904 13542 29952 13552
rect 29952 13532 30252 13542
rect 33856 12658 34756 12668
rect 33856 12206 34756 12216
rect 11010 7962 11198 7972
rect 11010 7842 11198 7852
rect 12186 7962 12374 7972
rect 12186 7842 12374 7852
rect 13362 7962 13550 7972
rect 13362 7842 13550 7852
rect 14538 7962 14726 7972
rect 14538 7842 14726 7852
rect 15714 7962 15902 7972
rect 15714 7842 15902 7852
rect 16890 7962 17078 7972
rect 16890 7842 17078 7852
rect 18066 7962 18254 7972
rect 18066 7842 18254 7852
rect 19242 7962 19430 7972
rect 19242 7842 19430 7852
rect 20418 7962 20606 7972
rect 20418 7842 20606 7852
rect 21594 7962 21782 7972
rect 21594 7842 21782 7852
rect 22770 7962 22958 7972
rect 22770 7842 22958 7852
rect 23946 7962 24134 7972
rect 23946 7842 24134 7852
rect 25122 7962 25310 7972
rect 25122 7842 25310 7852
rect 26298 7962 26486 7972
rect 26298 7842 26486 7852
rect 27474 7962 27662 7972
rect 27474 7842 27662 7852
rect 28650 7962 28838 7972
rect 28650 7842 28838 7852
rect 31002 7962 31190 7972
rect 31002 7842 31190 7852
rect 32178 7962 32366 7972
rect 32178 7842 32366 7852
rect 33354 7962 33542 7972
rect 33354 7842 33542 7852
rect 35706 7962 35894 7972
rect 35706 7842 35894 7852
rect 36882 7962 37070 7972
rect 36882 7842 37070 7852
rect 38058 7962 38246 7972
rect 38058 7842 38246 7852
rect 24202 6960 26348 7086
rect 24202 6846 24522 6960
rect 23670 6836 23990 6846
rect 23724 6704 23936 6836
rect 23670 6580 23990 6704
rect 24202 6836 24256 6846
rect 24202 6694 24256 6704
rect 24468 6836 24522 6846
rect 24468 6694 24522 6704
rect 24734 6836 25054 6960
rect 24788 6704 25000 6836
rect 24734 6698 25054 6704
rect 25266 6836 25320 6846
rect 25266 6698 25320 6704
rect 25532 6836 25586 6846
rect 25532 6698 25586 6704
rect 25266 6580 25586 6698
rect 22908 6454 25586 6580
rect 22908 5570 23124 6454
rect 26132 6076 26348 6960
rect 24202 5950 26348 6076
rect 24202 5836 24522 5950
rect 24742 5836 25062 5950
rect 23670 5826 23724 5836
rect 23670 5684 23724 5694
rect 23936 5826 23990 5836
rect 23936 5684 23990 5694
rect 24202 5826 24256 5836
rect 24202 5684 24256 5694
rect 24468 5826 24522 5836
rect 24468 5684 24522 5694
rect 24734 5826 24788 5836
rect 24734 5684 24788 5694
rect 25000 5826 25054 5836
rect 25000 5684 25054 5694
rect 25266 5826 25320 5836
rect 25266 5684 25320 5694
rect 25532 5826 25586 5836
rect 25532 5684 25586 5694
rect 23670 5570 23990 5684
rect 25266 5570 25586 5684
rect 22908 5444 25586 5570
rect 22908 4560 23124 5444
rect 26132 5066 26348 5950
rect 24202 4940 26348 5066
rect 24202 4826 24522 4940
rect 23670 4816 23724 4826
rect 23670 4674 23724 4684
rect 23936 4816 23990 4826
rect 23936 4674 23990 4684
rect 24202 4816 24256 4826
rect 24202 4674 24256 4684
rect 24468 4816 24522 4826
rect 24468 4674 24522 4684
rect 24734 4822 25054 4940
rect 24734 4816 24788 4822
rect 24734 4674 24788 4684
rect 25000 4816 25054 4822
rect 25000 4674 25054 4684
rect 25266 4816 25320 4826
rect 25266 4674 25320 4684
rect 25532 4816 25586 4826
rect 25532 4674 25586 4684
rect 23670 4560 23990 4674
rect 25266 4560 25586 4674
rect 22908 4434 25586 4560
rect 22908 3550 23124 4434
rect 26132 4056 26348 4940
rect 30580 5340 31062 5350
rect 31886 5304 32474 5314
rect 31062 4984 31886 5150
rect 30580 4792 31062 4802
rect 31886 4746 32474 4756
rect 24202 3930 26348 4056
rect 24202 3816 24522 3930
rect 23670 3806 23724 3816
rect 23670 3664 23724 3674
rect 23936 3806 23990 3816
rect 23936 3664 23990 3674
rect 24202 3806 24256 3816
rect 24202 3664 24256 3674
rect 24468 3806 24522 3816
rect 24468 3664 24522 3674
rect 24734 3816 25054 3930
rect 24734 3806 24788 3816
rect 24734 3664 24788 3674
rect 25000 3806 25054 3816
rect 25000 3664 25054 3674
rect 25266 3806 25320 3816
rect 25266 3664 25320 3674
rect 25532 3806 25586 3816
rect 25532 3664 25586 3674
rect 23670 3550 23990 3664
rect 25266 3550 25586 3664
rect 22908 3424 25586 3550
rect 29724 3712 30504 3722
rect 24368 3258 29724 3268
rect 24862 3130 29724 3258
rect 24368 3120 29724 3130
rect 30576 3348 30952 3358
rect 30504 3120 30576 3268
rect 30576 2908 30952 2918
rect 29724 2892 30504 2902
rect 30792 1224 31548 1234
rect 23940 644 25292 654
rect 30792 548 31548 558
rect 23940 522 25292 532
<< via2 >>
rect 20014 15572 20124 15644
rect 20494 15572 20604 15644
rect 20974 15572 21084 15644
rect 21454 15572 21564 15644
rect 21934 15572 22044 15644
rect 22414 15572 22524 15644
rect 22894 15572 23004 15644
rect 23374 15572 23484 15644
rect 23854 15572 23964 15644
rect 24334 15572 24444 15644
rect 24814 15572 24924 15644
rect 25294 15572 25404 15644
rect 25774 15572 25884 15644
rect 26254 15572 26364 15644
rect 26734 15572 26844 15644
rect 27214 15572 27324 15644
rect 27694 15572 27804 15644
rect 28174 15572 28284 15644
rect 28654 15572 28764 15644
rect 29134 15572 29244 15644
rect 29952 15158 30252 15458
rect 29952 14350 30252 14650
rect 29952 13542 30252 13842
rect 33856 12216 34756 12658
rect 11010 7852 11198 7962
rect 12186 7852 12374 7962
rect 13362 7852 13550 7962
rect 14538 7852 14726 7962
rect 15714 7852 15902 7962
rect 16890 7852 17078 7962
rect 18066 7852 18254 7962
rect 19242 7852 19430 7962
rect 20418 7852 20606 7962
rect 21594 7852 21782 7962
rect 22770 7852 22958 7962
rect 23946 7852 24134 7962
rect 25122 7852 25310 7962
rect 26298 7852 26486 7962
rect 27474 7852 27662 7962
rect 28650 7852 28838 7962
rect 31002 7852 31190 7962
rect 32178 7852 32366 7962
rect 33354 7852 33542 7962
rect 35706 7852 35894 7962
rect 36882 7852 37070 7962
rect 38058 7852 38246 7962
rect 31886 4756 32474 5304
rect 29724 2902 30504 3712
rect 23940 532 25292 644
rect 30792 558 31548 1224
<< metal3 >>
rect 20004 15644 20134 15649
rect 20004 15572 20014 15644
rect 20124 15572 20134 15644
rect 20004 15567 20134 15572
rect 20484 15644 20614 15649
rect 20484 15572 20494 15644
rect 20604 15572 20614 15644
rect 20484 15567 20614 15572
rect 20964 15644 21094 15649
rect 20964 15572 20974 15644
rect 21084 15572 21094 15644
rect 20964 15567 21094 15572
rect 21444 15644 21574 15649
rect 21444 15572 21454 15644
rect 21564 15572 21574 15644
rect 21444 15567 21574 15572
rect 21924 15644 22054 15649
rect 21924 15572 21934 15644
rect 22044 15572 22054 15644
rect 21924 15567 22054 15572
rect 22404 15644 22534 15649
rect 22404 15572 22414 15644
rect 22524 15572 22534 15644
rect 22404 15567 22534 15572
rect 22884 15644 23014 15649
rect 22884 15572 22894 15644
rect 23004 15572 23014 15644
rect 22884 15567 23014 15572
rect 23364 15644 23494 15649
rect 23364 15572 23374 15644
rect 23484 15572 23494 15644
rect 23364 15567 23494 15572
rect 23844 15644 23974 15649
rect 23844 15572 23854 15644
rect 23964 15572 23974 15644
rect 23844 15567 23974 15572
rect 24324 15644 24454 15649
rect 24324 15572 24334 15644
rect 24444 15572 24454 15644
rect 24324 15567 24454 15572
rect 24804 15644 24934 15649
rect 24804 15572 24814 15644
rect 24924 15572 24934 15644
rect 24804 15567 24934 15572
rect 25284 15644 25414 15649
rect 25284 15572 25294 15644
rect 25404 15572 25414 15644
rect 25284 15567 25414 15572
rect 25764 15644 25894 15649
rect 25764 15572 25774 15644
rect 25884 15572 25894 15644
rect 25764 15567 25894 15572
rect 26244 15644 26374 15649
rect 26244 15572 26254 15644
rect 26364 15572 26374 15644
rect 26244 15567 26374 15572
rect 26724 15644 26854 15649
rect 26724 15572 26734 15644
rect 26844 15572 26854 15644
rect 26724 15567 26854 15572
rect 27204 15644 27334 15649
rect 27204 15572 27214 15644
rect 27324 15572 27334 15644
rect 27204 15567 27334 15572
rect 27684 15644 27814 15649
rect 27684 15572 27694 15644
rect 27804 15572 27814 15644
rect 27684 15567 27814 15572
rect 28164 15644 28294 15649
rect 28164 15572 28174 15644
rect 28284 15572 28294 15644
rect 28164 15567 28294 15572
rect 28644 15644 28774 15649
rect 28644 15572 28654 15644
rect 28764 15572 28774 15644
rect 28644 15567 28774 15572
rect 29124 15644 29254 15649
rect 29124 15572 29134 15644
rect 29244 15572 29254 15644
rect 29124 15567 29254 15572
rect 29942 15462 30262 15463
rect 29942 15458 30272 15462
rect 29942 15158 29952 15458
rect 30252 15158 30272 15458
rect 29942 15153 30272 15158
rect 29952 14655 30272 15153
rect 29942 14650 30272 14655
rect 29942 14350 29952 14650
rect 30252 14350 30272 14650
rect 29942 14345 30272 14350
rect 29952 13847 30272 14345
rect 29942 13842 30272 13847
rect 29942 13542 29952 13842
rect 30252 13542 30272 13842
rect 29942 13537 30272 13542
rect 11000 7962 11208 7967
rect 11000 7852 11010 7962
rect 11198 7852 11208 7962
rect 11000 7847 11208 7852
rect 12176 7962 12384 7967
rect 12176 7852 12186 7962
rect 12374 7852 12384 7962
rect 12176 7847 12384 7852
rect 13352 7962 13560 7967
rect 13352 7852 13362 7962
rect 13550 7852 13560 7962
rect 13352 7847 13560 7852
rect 14528 7962 14736 7967
rect 14528 7852 14538 7962
rect 14726 7852 14736 7962
rect 14528 7847 14736 7852
rect 15704 7962 15912 7967
rect 15704 7852 15714 7962
rect 15902 7852 15912 7962
rect 15704 7847 15912 7852
rect 16880 7962 17088 7967
rect 16880 7852 16890 7962
rect 17078 7852 17088 7962
rect 16880 7847 17088 7852
rect 18056 7962 18264 7967
rect 18056 7852 18066 7962
rect 18254 7852 18264 7962
rect 18056 7847 18264 7852
rect 19232 7962 19440 7967
rect 19232 7852 19242 7962
rect 19430 7852 19440 7962
rect 19232 7847 19440 7852
rect 20408 7962 20616 7967
rect 20408 7852 20418 7962
rect 20606 7852 20616 7962
rect 20408 7847 20616 7852
rect 21584 7962 21792 7967
rect 21584 7852 21594 7962
rect 21782 7852 21792 7962
rect 21584 7847 21792 7852
rect 22760 7962 22968 7967
rect 22760 7852 22770 7962
rect 22958 7852 22968 7962
rect 22760 7847 22968 7852
rect 23936 7962 24144 7967
rect 23936 7852 23946 7962
rect 24134 7852 24144 7962
rect 23936 7847 24144 7852
rect 25112 7962 25320 7967
rect 25112 7852 25122 7962
rect 25310 7852 25320 7962
rect 25112 7847 25320 7852
rect 26288 7962 26496 7967
rect 26288 7852 26298 7962
rect 26486 7852 26496 7962
rect 26288 7847 26496 7852
rect 27464 7962 27672 7967
rect 27464 7852 27474 7962
rect 27662 7852 27672 7962
rect 27464 7847 27672 7852
rect 28640 7962 28848 7967
rect 28640 7852 28650 7962
rect 28838 7852 28848 7962
rect 28640 7847 28848 7852
rect 29952 3717 30272 13537
rect 33846 12658 34766 12663
rect 33846 12216 33856 12658
rect 34756 12216 34766 12658
rect 33846 12211 34766 12216
rect 30992 7962 31200 7967
rect 30992 7852 31002 7962
rect 31190 7852 31200 7962
rect 30992 7847 31200 7852
rect 32168 7962 32376 7967
rect 32168 7852 32178 7962
rect 32366 7852 32376 7962
rect 32168 7847 32376 7852
rect 33344 7962 33552 7967
rect 33344 7852 33354 7962
rect 33542 7852 33552 7962
rect 33344 7847 33552 7852
rect 33900 7092 34738 12211
rect 35696 7962 35904 7967
rect 35696 7852 35706 7962
rect 35894 7852 35904 7962
rect 35696 7847 35904 7852
rect 36872 7962 37080 7967
rect 36872 7852 36882 7962
rect 37070 7852 37080 7962
rect 36872 7847 37080 7852
rect 38048 7962 38256 7967
rect 38048 7852 38058 7962
rect 38246 7852 38256 7962
rect 38048 7847 38256 7852
rect 33862 6192 33872 7092
rect 34772 6192 34782 7092
rect 31876 5304 32484 5309
rect 31876 4756 31886 5304
rect 32474 5148 32484 5304
rect 33046 5148 36230 5294
rect 32474 4836 36230 5148
rect 32474 4756 32484 4836
rect 31876 4751 32484 4756
rect 29714 3712 30514 3717
rect 29714 2902 29724 3712
rect 30504 2902 30514 3712
rect 29714 2897 30514 2902
rect 33046 2094 36230 4836
rect 30782 1224 31558 1229
rect 23930 644 25302 649
rect 23930 532 23940 644
rect 25292 532 25302 644
rect 30782 558 30792 1224
rect 31548 558 31558 1224
rect 30782 553 31558 558
rect 23930 527 25302 532
<< via3 >>
rect 20014 15572 20124 15644
rect 20494 15572 20604 15644
rect 20974 15572 21084 15644
rect 21454 15572 21564 15644
rect 21934 15572 22044 15644
rect 22414 15572 22524 15644
rect 22894 15572 23004 15644
rect 23374 15572 23484 15644
rect 23854 15572 23964 15644
rect 24334 15572 24444 15644
rect 24814 15572 24924 15644
rect 25294 15572 25404 15644
rect 25774 15572 25884 15644
rect 26254 15572 26364 15644
rect 26734 15572 26844 15644
rect 27214 15572 27324 15644
rect 27694 15572 27804 15644
rect 28174 15572 28284 15644
rect 28654 15572 28764 15644
rect 29134 15572 29244 15644
rect 11010 7852 11198 7962
rect 12186 7852 12374 7962
rect 13362 7852 13550 7962
rect 14538 7852 14726 7962
rect 15714 7852 15902 7962
rect 16890 7852 17078 7962
rect 18066 7852 18254 7962
rect 19242 7852 19430 7962
rect 20418 7852 20606 7962
rect 21594 7852 21782 7962
rect 22770 7852 22958 7962
rect 23946 7852 24134 7962
rect 25122 7852 25310 7962
rect 26298 7852 26486 7962
rect 27474 7852 27662 7962
rect 28650 7852 28838 7962
rect 31002 7852 31190 7962
rect 32178 7852 32366 7962
rect 33354 7852 33542 7962
rect 35706 7852 35894 7962
rect 36882 7852 37070 7962
rect 38058 7852 38246 7962
rect 33872 6192 34772 7092
rect 23940 532 25292 644
rect 30792 558 31548 1224
<< mimcap >>
rect 33146 5154 36146 5194
rect 33146 2234 33186 5154
rect 36106 2234 36146 5154
rect 33146 2194 36146 2234
<< mimcapcontact >>
rect 33186 2234 36106 5154
<< metal4 >>
rect 7082 15644 35696 16350
rect 7082 15572 20014 15644
rect 20124 15572 20494 15644
rect 20604 15572 20974 15644
rect 21084 15572 21454 15644
rect 21564 15572 21934 15644
rect 22044 15572 22414 15644
rect 22524 15572 22894 15644
rect 23004 15572 23374 15644
rect 23484 15572 23854 15644
rect 23964 15572 24334 15644
rect 24444 15572 24814 15644
rect 24924 15572 25294 15644
rect 25404 15572 25774 15644
rect 25884 15572 26254 15644
rect 26364 15572 26734 15644
rect 26844 15572 27214 15644
rect 27324 15572 27694 15644
rect 27804 15572 28174 15644
rect 28284 15572 28654 15644
rect 28764 15572 29134 15644
rect 29244 15572 35696 15644
rect 7082 15086 35696 15572
rect 7082 15084 13862 15086
rect 7082 1538 8398 15084
rect 8986 7962 39470 8826
rect 8986 7852 11010 7962
rect 11198 7852 12186 7962
rect 12374 7852 13362 7962
rect 13550 7852 14538 7962
rect 14726 7852 15714 7962
rect 15902 7852 16890 7962
rect 17078 7852 18066 7962
rect 18254 7852 19242 7962
rect 19430 7852 20418 7962
rect 20606 7852 21594 7962
rect 21782 7852 22770 7962
rect 22958 7852 23946 7962
rect 24134 7852 25122 7962
rect 25310 7852 26298 7962
rect 26486 7852 27474 7962
rect 27662 7852 28650 7962
rect 28838 7852 31002 7962
rect 31190 7852 32178 7962
rect 32366 7852 33354 7962
rect 33542 7852 35706 7962
rect 35894 7852 36882 7962
rect 37070 7852 38058 7962
rect 38246 7852 39470 7962
rect 8986 7294 39470 7852
rect 33871 7092 34773 7093
rect 33871 6192 33872 7092
rect 34772 6192 34773 7092
rect 33871 6191 34773 6192
rect 33928 5155 34730 6191
rect 33185 5154 36107 5155
rect 33185 2234 33186 5154
rect 36106 2234 36107 5154
rect 33185 2233 36107 2234
rect 7082 1224 31958 1538
rect 7082 644 30792 1224
rect 7082 532 23940 644
rect 25292 558 30792 644
rect 31548 558 31958 1224
rect 25292 532 31958 558
rect 7082 6 31958 532
<< labels >>
flabel metal4 9160 8150 9160 8150 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal4 9644 400 9644 400 0 FreeSans 1600 0 0 0 vss
port 4 nsew
flabel metal1 37260 12404 37260 12404 0 FreeSans 1600 0 0 0 vout
port 5 nsew
flabel metal1 10784 9208 10784 9208 0 FreeSans 1600 0 0 0 vbias
port 3 nsew
flabel metal2 23010 5540 23010 5540 0 FreeSans 1600 0 0 0 vn
port 2 nsew
flabel metal2 26244 5942 26244 5942 0 FreeSans 1600 0 0 0 vp
port 1 nsew
<< end >>
