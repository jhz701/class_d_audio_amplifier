magic
tech sky130A
magscale 1 2
timestamp 1627371027
<< nwell >>
rect 42914 9266 71934 13130
rect 55926 4726 58922 8756
<< pwell >>
rect 52218 14650 62632 17286
rect 56538 1948 58312 4564
<< pmoslvt >>
rect 43406 11798 43806 12598
rect 43994 11798 44394 12598
rect 44582 11798 44982 12598
rect 45170 11798 45570 12598
rect 45758 11798 46158 12598
rect 46346 11798 46746 12598
rect 46934 11798 47334 12598
rect 47522 11798 47922 12598
rect 48110 11798 48510 12598
rect 48698 11798 49098 12598
rect 49286 11798 49686 12598
rect 49874 11798 50274 12598
rect 50462 11798 50862 12598
rect 51050 11798 51450 12598
rect 51638 11798 52038 12598
rect 52226 11798 52626 12598
rect 52814 11798 53214 12598
rect 53402 11798 53802 12598
rect 53990 11798 54390 12598
rect 54578 11798 54978 12598
rect 55166 11798 55566 12598
rect 55754 11798 56154 12598
rect 56342 11798 56742 12598
rect 56930 11798 57330 12598
rect 57518 11798 57918 12598
rect 58106 11798 58506 12598
rect 58694 11798 59094 12598
rect 59282 11798 59682 12598
rect 59870 11798 60270 12598
rect 60458 11798 60858 12598
rect 61046 11798 61446 12598
rect 61634 11798 62034 12598
rect 62222 11798 62622 12598
rect 62810 11798 63210 12598
rect 63398 11798 63798 12598
rect 63986 11798 64386 12598
rect 64574 11798 64974 12598
rect 65162 11798 65562 12598
rect 65750 11798 66150 12598
rect 66338 11798 66738 12598
rect 66926 11798 67326 12598
rect 67514 11798 67914 12598
rect 68102 11798 68502 12598
rect 68690 11798 69090 12598
rect 69278 11798 69678 12598
rect 69866 11798 70266 12598
rect 70454 11798 70854 12598
rect 71042 11798 71442 12598
rect 43406 10798 43806 11598
rect 43994 10798 44394 11598
rect 44582 10798 44982 11598
rect 45170 10798 45570 11598
rect 45758 10798 46158 11598
rect 46346 10798 46746 11598
rect 46934 10798 47334 11598
rect 47522 10798 47922 11598
rect 48110 10798 48510 11598
rect 48698 10798 49098 11598
rect 49286 10798 49686 11598
rect 49874 10798 50274 11598
rect 50462 10798 50862 11598
rect 51050 10798 51450 11598
rect 51638 10798 52038 11598
rect 52226 10798 52626 11598
rect 52814 10798 53214 11598
rect 53402 10798 53802 11598
rect 53990 10798 54390 11598
rect 54578 10798 54978 11598
rect 55166 10798 55566 11598
rect 55754 10798 56154 11598
rect 56342 10798 56742 11598
rect 56930 10798 57330 11598
rect 57518 10798 57918 11598
rect 58106 10798 58506 11598
rect 58694 10798 59094 11598
rect 59282 10798 59682 11598
rect 59870 10798 60270 11598
rect 60458 10798 60858 11598
rect 61046 10798 61446 11598
rect 61634 10798 62034 11598
rect 62222 10798 62622 11598
rect 62810 10798 63210 11598
rect 63398 10798 63798 11598
rect 63986 10798 64386 11598
rect 64574 10798 64974 11598
rect 65162 10798 65562 11598
rect 65750 10798 66150 11598
rect 66338 10798 66738 11598
rect 66926 10798 67326 11598
rect 67514 10798 67914 11598
rect 68102 10798 68502 11598
rect 68690 10798 69090 11598
rect 69278 10798 69678 11598
rect 69866 10798 70266 11598
rect 70454 10798 70854 11598
rect 71042 10798 71442 11598
rect 43406 9798 43806 10598
rect 43994 9798 44394 10598
rect 44582 9798 44982 10598
rect 45170 9798 45570 10598
rect 45758 9798 46158 10598
rect 46346 9798 46746 10598
rect 46934 9798 47334 10598
rect 47522 9798 47922 10598
rect 48110 9798 48510 10598
rect 48698 9798 49098 10598
rect 49286 9798 49686 10598
rect 49874 9798 50274 10598
rect 50462 9798 50862 10598
rect 51050 9798 51450 10598
rect 51638 9798 52038 10598
rect 52226 9798 52626 10598
rect 52814 9798 53214 10598
rect 53402 9798 53802 10598
rect 53990 9798 54390 10598
rect 54578 9798 54978 10598
rect 55166 9798 55566 10598
rect 55754 9798 56154 10598
rect 56342 9798 56742 10598
rect 56930 9798 57330 10598
rect 57518 9798 57918 10598
rect 58106 9798 58506 10598
rect 58694 9798 59094 10598
rect 59282 9798 59682 10598
rect 59870 9798 60270 10598
rect 60458 9798 60858 10598
rect 61046 9798 61446 10598
rect 61634 9798 62034 10598
rect 62222 9798 62622 10598
rect 62810 9798 63210 10598
rect 63398 9798 63798 10598
rect 63986 9798 64386 10598
rect 64574 9798 64974 10598
rect 65162 9798 65562 10598
rect 65750 9798 66150 10598
rect 66338 9798 66738 10598
rect 66926 9798 67326 10598
rect 67514 9798 67914 10598
rect 68102 9798 68502 10598
rect 68690 9798 69090 10598
rect 69278 9798 69678 10598
rect 69866 9798 70266 10598
rect 70454 9798 70854 10598
rect 71042 9798 71442 10598
rect 56458 7352 56528 8152
rect 56724 7352 56794 8152
rect 56990 7352 57060 8152
rect 57256 7352 57326 8152
rect 57522 7352 57592 8152
rect 57788 7352 57858 8152
rect 58054 7352 58124 8152
rect 58320 7352 58390 8152
rect 56458 6342 56528 7142
rect 56724 6342 56794 7142
rect 56990 6342 57060 7142
rect 57256 6342 57326 7142
rect 57522 6342 57592 7142
rect 57788 6342 57858 7142
rect 58054 6342 58124 7142
rect 58320 6342 58390 7142
rect 56458 5332 56528 6132
rect 56724 5332 56794 6132
rect 56990 5332 57060 6132
rect 57256 5332 57326 6132
rect 57522 5332 57592 6132
rect 57788 5332 57858 6132
rect 58054 5332 58124 6132
rect 58320 5332 58390 6132
<< nmoslvt >>
rect 52710 16072 52780 16672
rect 52950 16072 53020 16672
rect 53190 16072 53260 16672
rect 53430 16072 53500 16672
rect 53670 16072 53740 16672
rect 53910 16072 53980 16672
rect 54150 16072 54220 16672
rect 54390 16072 54460 16672
rect 54630 16072 54700 16672
rect 54870 16072 54940 16672
rect 55110 16072 55180 16672
rect 55350 16072 55420 16672
rect 55590 16072 55660 16672
rect 55830 16072 55900 16672
rect 56070 16072 56140 16672
rect 56310 16072 56380 16672
rect 56550 16072 56620 16672
rect 56790 16072 56860 16672
rect 57030 16072 57100 16672
rect 57270 16072 57340 16672
rect 57510 16072 57580 16672
rect 57750 16072 57820 16672
rect 57990 16072 58060 16672
rect 58230 16072 58300 16672
rect 58470 16072 58540 16672
rect 58710 16072 58780 16672
rect 58950 16072 59020 16672
rect 59190 16072 59260 16672
rect 59430 16072 59500 16672
rect 59670 16072 59740 16672
rect 59910 16072 59980 16672
rect 60150 16072 60220 16672
rect 60390 16072 60460 16672
rect 60630 16072 60700 16672
rect 60870 16072 60940 16672
rect 61110 16072 61180 16672
rect 61350 16072 61420 16672
rect 61590 16072 61660 16672
rect 61830 16072 61900 16672
rect 62070 16072 62140 16672
rect 52710 15264 52780 15864
rect 52950 15264 53020 15864
rect 53190 15264 53260 15864
rect 53430 15264 53500 15864
rect 53670 15264 53740 15864
rect 53910 15264 53980 15864
rect 54150 15264 54220 15864
rect 54390 15264 54460 15864
rect 54630 15264 54700 15864
rect 54870 15264 54940 15864
rect 55110 15264 55180 15864
rect 55350 15264 55420 15864
rect 55590 15264 55660 15864
rect 55830 15264 55900 15864
rect 56070 15264 56140 15864
rect 56310 15264 56380 15864
rect 56550 15264 56620 15864
rect 56790 15264 56860 15864
rect 57030 15264 57100 15864
rect 57270 15264 57340 15864
rect 57510 15264 57580 15864
rect 57750 15264 57820 15864
rect 57990 15264 58060 15864
rect 58230 15264 58300 15864
rect 58470 15264 58540 15864
rect 58710 15264 58780 15864
rect 58950 15264 59020 15864
rect 59190 15264 59260 15864
rect 59430 15264 59500 15864
rect 59670 15264 59740 15864
rect 59910 15264 59980 15864
rect 60150 15264 60220 15864
rect 60390 15264 60460 15864
rect 60630 15264 60700 15864
rect 60870 15264 60940 15864
rect 61110 15264 61180 15864
rect 61350 15264 61420 15864
rect 61590 15264 61660 15864
rect 61830 15264 61900 15864
rect 62070 15264 62140 15864
rect 57030 3360 57100 3960
rect 57270 3360 57340 3960
rect 57510 3360 57580 3960
rect 57750 3360 57820 3960
rect 57030 2552 57100 3152
rect 57270 2552 57340 3152
rect 57510 2552 57580 3152
rect 57750 2552 57820 3152
<< ndiff >>
rect 52652 16660 52710 16672
rect 52652 16084 52664 16660
rect 52698 16084 52710 16660
rect 52652 16072 52710 16084
rect 52780 16660 52838 16672
rect 52780 16084 52792 16660
rect 52826 16084 52838 16660
rect 52780 16072 52838 16084
rect 52892 16660 52950 16672
rect 52892 16084 52904 16660
rect 52938 16084 52950 16660
rect 52892 16072 52950 16084
rect 53020 16660 53078 16672
rect 53020 16084 53032 16660
rect 53066 16084 53078 16660
rect 53020 16072 53078 16084
rect 53132 16660 53190 16672
rect 53132 16084 53144 16660
rect 53178 16084 53190 16660
rect 53132 16072 53190 16084
rect 53260 16660 53318 16672
rect 53260 16084 53272 16660
rect 53306 16084 53318 16660
rect 53260 16072 53318 16084
rect 53372 16660 53430 16672
rect 53372 16084 53384 16660
rect 53418 16084 53430 16660
rect 53372 16072 53430 16084
rect 53500 16660 53558 16672
rect 53500 16084 53512 16660
rect 53546 16084 53558 16660
rect 53500 16072 53558 16084
rect 53612 16660 53670 16672
rect 53612 16084 53624 16660
rect 53658 16084 53670 16660
rect 53612 16072 53670 16084
rect 53740 16660 53798 16672
rect 53740 16084 53752 16660
rect 53786 16084 53798 16660
rect 53740 16072 53798 16084
rect 53852 16660 53910 16672
rect 53852 16084 53864 16660
rect 53898 16084 53910 16660
rect 53852 16072 53910 16084
rect 53980 16660 54038 16672
rect 53980 16084 53992 16660
rect 54026 16084 54038 16660
rect 53980 16072 54038 16084
rect 54092 16660 54150 16672
rect 54092 16084 54104 16660
rect 54138 16084 54150 16660
rect 54092 16072 54150 16084
rect 54220 16660 54278 16672
rect 54220 16084 54232 16660
rect 54266 16084 54278 16660
rect 54220 16072 54278 16084
rect 54332 16660 54390 16672
rect 54332 16084 54344 16660
rect 54378 16084 54390 16660
rect 54332 16072 54390 16084
rect 54460 16660 54518 16672
rect 54460 16084 54472 16660
rect 54506 16084 54518 16660
rect 54460 16072 54518 16084
rect 54572 16660 54630 16672
rect 54572 16084 54584 16660
rect 54618 16084 54630 16660
rect 54572 16072 54630 16084
rect 54700 16660 54758 16672
rect 54700 16084 54712 16660
rect 54746 16084 54758 16660
rect 54700 16072 54758 16084
rect 54812 16660 54870 16672
rect 54812 16084 54824 16660
rect 54858 16084 54870 16660
rect 54812 16072 54870 16084
rect 54940 16660 54998 16672
rect 54940 16084 54952 16660
rect 54986 16084 54998 16660
rect 54940 16072 54998 16084
rect 55052 16660 55110 16672
rect 55052 16084 55064 16660
rect 55098 16084 55110 16660
rect 55052 16072 55110 16084
rect 55180 16660 55238 16672
rect 55180 16084 55192 16660
rect 55226 16084 55238 16660
rect 55180 16072 55238 16084
rect 55292 16660 55350 16672
rect 55292 16084 55304 16660
rect 55338 16084 55350 16660
rect 55292 16072 55350 16084
rect 55420 16660 55478 16672
rect 55420 16084 55432 16660
rect 55466 16084 55478 16660
rect 55420 16072 55478 16084
rect 55532 16660 55590 16672
rect 55532 16084 55544 16660
rect 55578 16084 55590 16660
rect 55532 16072 55590 16084
rect 55660 16660 55718 16672
rect 55660 16084 55672 16660
rect 55706 16084 55718 16660
rect 55660 16072 55718 16084
rect 55772 16660 55830 16672
rect 55772 16084 55784 16660
rect 55818 16084 55830 16660
rect 55772 16072 55830 16084
rect 55900 16660 55958 16672
rect 55900 16084 55912 16660
rect 55946 16084 55958 16660
rect 55900 16072 55958 16084
rect 56012 16660 56070 16672
rect 56012 16084 56024 16660
rect 56058 16084 56070 16660
rect 56012 16072 56070 16084
rect 56140 16660 56198 16672
rect 56140 16084 56152 16660
rect 56186 16084 56198 16660
rect 56140 16072 56198 16084
rect 56252 16660 56310 16672
rect 56252 16084 56264 16660
rect 56298 16084 56310 16660
rect 56252 16072 56310 16084
rect 56380 16660 56438 16672
rect 56380 16084 56392 16660
rect 56426 16084 56438 16660
rect 56380 16072 56438 16084
rect 56492 16660 56550 16672
rect 56492 16084 56504 16660
rect 56538 16084 56550 16660
rect 56492 16072 56550 16084
rect 56620 16660 56678 16672
rect 56620 16084 56632 16660
rect 56666 16084 56678 16660
rect 56620 16072 56678 16084
rect 56732 16660 56790 16672
rect 56732 16084 56744 16660
rect 56778 16084 56790 16660
rect 56732 16072 56790 16084
rect 56860 16660 56918 16672
rect 56860 16084 56872 16660
rect 56906 16084 56918 16660
rect 56860 16072 56918 16084
rect 56972 16660 57030 16672
rect 56972 16084 56984 16660
rect 57018 16084 57030 16660
rect 56972 16072 57030 16084
rect 57100 16660 57158 16672
rect 57100 16084 57112 16660
rect 57146 16084 57158 16660
rect 57100 16072 57158 16084
rect 57212 16660 57270 16672
rect 57212 16084 57224 16660
rect 57258 16084 57270 16660
rect 57212 16072 57270 16084
rect 57340 16660 57398 16672
rect 57340 16084 57352 16660
rect 57386 16084 57398 16660
rect 57340 16072 57398 16084
rect 57452 16660 57510 16672
rect 57452 16084 57464 16660
rect 57498 16084 57510 16660
rect 57452 16072 57510 16084
rect 57580 16660 57638 16672
rect 57580 16084 57592 16660
rect 57626 16084 57638 16660
rect 57580 16072 57638 16084
rect 57692 16660 57750 16672
rect 57692 16084 57704 16660
rect 57738 16084 57750 16660
rect 57692 16072 57750 16084
rect 57820 16660 57878 16672
rect 57820 16084 57832 16660
rect 57866 16084 57878 16660
rect 57820 16072 57878 16084
rect 57932 16660 57990 16672
rect 57932 16084 57944 16660
rect 57978 16084 57990 16660
rect 57932 16072 57990 16084
rect 58060 16660 58118 16672
rect 58060 16084 58072 16660
rect 58106 16084 58118 16660
rect 58060 16072 58118 16084
rect 58172 16660 58230 16672
rect 58172 16084 58184 16660
rect 58218 16084 58230 16660
rect 58172 16072 58230 16084
rect 58300 16660 58358 16672
rect 58300 16084 58312 16660
rect 58346 16084 58358 16660
rect 58300 16072 58358 16084
rect 58412 16660 58470 16672
rect 58412 16084 58424 16660
rect 58458 16084 58470 16660
rect 58412 16072 58470 16084
rect 58540 16660 58598 16672
rect 58540 16084 58552 16660
rect 58586 16084 58598 16660
rect 58540 16072 58598 16084
rect 58652 16660 58710 16672
rect 58652 16084 58664 16660
rect 58698 16084 58710 16660
rect 58652 16072 58710 16084
rect 58780 16660 58838 16672
rect 58780 16084 58792 16660
rect 58826 16084 58838 16660
rect 58780 16072 58838 16084
rect 58892 16660 58950 16672
rect 58892 16084 58904 16660
rect 58938 16084 58950 16660
rect 58892 16072 58950 16084
rect 59020 16660 59078 16672
rect 59020 16084 59032 16660
rect 59066 16084 59078 16660
rect 59020 16072 59078 16084
rect 59132 16660 59190 16672
rect 59132 16084 59144 16660
rect 59178 16084 59190 16660
rect 59132 16072 59190 16084
rect 59260 16660 59318 16672
rect 59260 16084 59272 16660
rect 59306 16084 59318 16660
rect 59260 16072 59318 16084
rect 59372 16660 59430 16672
rect 59372 16084 59384 16660
rect 59418 16084 59430 16660
rect 59372 16072 59430 16084
rect 59500 16660 59558 16672
rect 59500 16084 59512 16660
rect 59546 16084 59558 16660
rect 59500 16072 59558 16084
rect 59612 16660 59670 16672
rect 59612 16084 59624 16660
rect 59658 16084 59670 16660
rect 59612 16072 59670 16084
rect 59740 16660 59798 16672
rect 59740 16084 59752 16660
rect 59786 16084 59798 16660
rect 59740 16072 59798 16084
rect 59852 16660 59910 16672
rect 59852 16084 59864 16660
rect 59898 16084 59910 16660
rect 59852 16072 59910 16084
rect 59980 16660 60038 16672
rect 59980 16084 59992 16660
rect 60026 16084 60038 16660
rect 59980 16072 60038 16084
rect 60092 16660 60150 16672
rect 60092 16084 60104 16660
rect 60138 16084 60150 16660
rect 60092 16072 60150 16084
rect 60220 16660 60278 16672
rect 60220 16084 60232 16660
rect 60266 16084 60278 16660
rect 60220 16072 60278 16084
rect 60332 16660 60390 16672
rect 60332 16084 60344 16660
rect 60378 16084 60390 16660
rect 60332 16072 60390 16084
rect 60460 16660 60518 16672
rect 60460 16084 60472 16660
rect 60506 16084 60518 16660
rect 60460 16072 60518 16084
rect 60572 16660 60630 16672
rect 60572 16084 60584 16660
rect 60618 16084 60630 16660
rect 60572 16072 60630 16084
rect 60700 16660 60758 16672
rect 60700 16084 60712 16660
rect 60746 16084 60758 16660
rect 60700 16072 60758 16084
rect 60812 16660 60870 16672
rect 60812 16084 60824 16660
rect 60858 16084 60870 16660
rect 60812 16072 60870 16084
rect 60940 16660 60998 16672
rect 60940 16084 60952 16660
rect 60986 16084 60998 16660
rect 60940 16072 60998 16084
rect 61052 16660 61110 16672
rect 61052 16084 61064 16660
rect 61098 16084 61110 16660
rect 61052 16072 61110 16084
rect 61180 16660 61238 16672
rect 61180 16084 61192 16660
rect 61226 16084 61238 16660
rect 61180 16072 61238 16084
rect 61292 16660 61350 16672
rect 61292 16084 61304 16660
rect 61338 16084 61350 16660
rect 61292 16072 61350 16084
rect 61420 16660 61478 16672
rect 61420 16084 61432 16660
rect 61466 16084 61478 16660
rect 61420 16072 61478 16084
rect 61532 16660 61590 16672
rect 61532 16084 61544 16660
rect 61578 16084 61590 16660
rect 61532 16072 61590 16084
rect 61660 16660 61718 16672
rect 61660 16084 61672 16660
rect 61706 16084 61718 16660
rect 61660 16072 61718 16084
rect 61772 16660 61830 16672
rect 61772 16084 61784 16660
rect 61818 16084 61830 16660
rect 61772 16072 61830 16084
rect 61900 16660 61958 16672
rect 61900 16084 61912 16660
rect 61946 16084 61958 16660
rect 61900 16072 61958 16084
rect 62012 16660 62070 16672
rect 62012 16084 62024 16660
rect 62058 16084 62070 16660
rect 62012 16072 62070 16084
rect 62140 16660 62198 16672
rect 62140 16084 62152 16660
rect 62186 16084 62198 16660
rect 62140 16072 62198 16084
rect 52652 15852 52710 15864
rect 52652 15276 52664 15852
rect 52698 15276 52710 15852
rect 52652 15264 52710 15276
rect 52780 15852 52838 15864
rect 52780 15276 52792 15852
rect 52826 15276 52838 15852
rect 52780 15264 52838 15276
rect 52892 15852 52950 15864
rect 52892 15276 52904 15852
rect 52938 15276 52950 15852
rect 52892 15264 52950 15276
rect 53020 15852 53078 15864
rect 53020 15276 53032 15852
rect 53066 15276 53078 15852
rect 53020 15264 53078 15276
rect 53132 15852 53190 15864
rect 53132 15276 53144 15852
rect 53178 15276 53190 15852
rect 53132 15264 53190 15276
rect 53260 15852 53318 15864
rect 53260 15276 53272 15852
rect 53306 15276 53318 15852
rect 53260 15264 53318 15276
rect 53372 15852 53430 15864
rect 53372 15276 53384 15852
rect 53418 15276 53430 15852
rect 53372 15264 53430 15276
rect 53500 15852 53558 15864
rect 53500 15276 53512 15852
rect 53546 15276 53558 15852
rect 53500 15264 53558 15276
rect 53612 15852 53670 15864
rect 53612 15276 53624 15852
rect 53658 15276 53670 15852
rect 53612 15264 53670 15276
rect 53740 15852 53798 15864
rect 53740 15276 53752 15852
rect 53786 15276 53798 15852
rect 53740 15264 53798 15276
rect 53852 15852 53910 15864
rect 53852 15276 53864 15852
rect 53898 15276 53910 15852
rect 53852 15264 53910 15276
rect 53980 15852 54038 15864
rect 53980 15276 53992 15852
rect 54026 15276 54038 15852
rect 53980 15264 54038 15276
rect 54092 15852 54150 15864
rect 54092 15276 54104 15852
rect 54138 15276 54150 15852
rect 54092 15264 54150 15276
rect 54220 15852 54278 15864
rect 54220 15276 54232 15852
rect 54266 15276 54278 15852
rect 54220 15264 54278 15276
rect 54332 15852 54390 15864
rect 54332 15276 54344 15852
rect 54378 15276 54390 15852
rect 54332 15264 54390 15276
rect 54460 15852 54518 15864
rect 54460 15276 54472 15852
rect 54506 15276 54518 15852
rect 54460 15264 54518 15276
rect 54572 15852 54630 15864
rect 54572 15276 54584 15852
rect 54618 15276 54630 15852
rect 54572 15264 54630 15276
rect 54700 15852 54758 15864
rect 54700 15276 54712 15852
rect 54746 15276 54758 15852
rect 54700 15264 54758 15276
rect 54812 15852 54870 15864
rect 54812 15276 54824 15852
rect 54858 15276 54870 15852
rect 54812 15264 54870 15276
rect 54940 15852 54998 15864
rect 54940 15276 54952 15852
rect 54986 15276 54998 15852
rect 54940 15264 54998 15276
rect 55052 15852 55110 15864
rect 55052 15276 55064 15852
rect 55098 15276 55110 15852
rect 55052 15264 55110 15276
rect 55180 15852 55238 15864
rect 55180 15276 55192 15852
rect 55226 15276 55238 15852
rect 55180 15264 55238 15276
rect 55292 15852 55350 15864
rect 55292 15276 55304 15852
rect 55338 15276 55350 15852
rect 55292 15264 55350 15276
rect 55420 15852 55478 15864
rect 55420 15276 55432 15852
rect 55466 15276 55478 15852
rect 55420 15264 55478 15276
rect 55532 15852 55590 15864
rect 55532 15276 55544 15852
rect 55578 15276 55590 15852
rect 55532 15264 55590 15276
rect 55660 15852 55718 15864
rect 55660 15276 55672 15852
rect 55706 15276 55718 15852
rect 55660 15264 55718 15276
rect 55772 15852 55830 15864
rect 55772 15276 55784 15852
rect 55818 15276 55830 15852
rect 55772 15264 55830 15276
rect 55900 15852 55958 15864
rect 55900 15276 55912 15852
rect 55946 15276 55958 15852
rect 55900 15264 55958 15276
rect 56012 15852 56070 15864
rect 56012 15276 56024 15852
rect 56058 15276 56070 15852
rect 56012 15264 56070 15276
rect 56140 15852 56198 15864
rect 56140 15276 56152 15852
rect 56186 15276 56198 15852
rect 56140 15264 56198 15276
rect 56252 15852 56310 15864
rect 56252 15276 56264 15852
rect 56298 15276 56310 15852
rect 56252 15264 56310 15276
rect 56380 15852 56438 15864
rect 56380 15276 56392 15852
rect 56426 15276 56438 15852
rect 56380 15264 56438 15276
rect 56492 15852 56550 15864
rect 56492 15276 56504 15852
rect 56538 15276 56550 15852
rect 56492 15264 56550 15276
rect 56620 15852 56678 15864
rect 56620 15276 56632 15852
rect 56666 15276 56678 15852
rect 56620 15264 56678 15276
rect 56732 15852 56790 15864
rect 56732 15276 56744 15852
rect 56778 15276 56790 15852
rect 56732 15264 56790 15276
rect 56860 15852 56918 15864
rect 56860 15276 56872 15852
rect 56906 15276 56918 15852
rect 56860 15264 56918 15276
rect 56972 15852 57030 15864
rect 56972 15276 56984 15852
rect 57018 15276 57030 15852
rect 56972 15264 57030 15276
rect 57100 15852 57158 15864
rect 57100 15276 57112 15852
rect 57146 15276 57158 15852
rect 57100 15264 57158 15276
rect 57212 15852 57270 15864
rect 57212 15276 57224 15852
rect 57258 15276 57270 15852
rect 57212 15264 57270 15276
rect 57340 15852 57398 15864
rect 57340 15276 57352 15852
rect 57386 15276 57398 15852
rect 57340 15264 57398 15276
rect 57452 15852 57510 15864
rect 57452 15276 57464 15852
rect 57498 15276 57510 15852
rect 57452 15264 57510 15276
rect 57580 15852 57638 15864
rect 57580 15276 57592 15852
rect 57626 15276 57638 15852
rect 57580 15264 57638 15276
rect 57692 15852 57750 15864
rect 57692 15276 57704 15852
rect 57738 15276 57750 15852
rect 57692 15264 57750 15276
rect 57820 15852 57878 15864
rect 57820 15276 57832 15852
rect 57866 15276 57878 15852
rect 57820 15264 57878 15276
rect 57932 15852 57990 15864
rect 57932 15276 57944 15852
rect 57978 15276 57990 15852
rect 57932 15264 57990 15276
rect 58060 15852 58118 15864
rect 58060 15276 58072 15852
rect 58106 15276 58118 15852
rect 58060 15264 58118 15276
rect 58172 15852 58230 15864
rect 58172 15276 58184 15852
rect 58218 15276 58230 15852
rect 58172 15264 58230 15276
rect 58300 15852 58358 15864
rect 58300 15276 58312 15852
rect 58346 15276 58358 15852
rect 58300 15264 58358 15276
rect 58412 15852 58470 15864
rect 58412 15276 58424 15852
rect 58458 15276 58470 15852
rect 58412 15264 58470 15276
rect 58540 15852 58598 15864
rect 58540 15276 58552 15852
rect 58586 15276 58598 15852
rect 58540 15264 58598 15276
rect 58652 15852 58710 15864
rect 58652 15276 58664 15852
rect 58698 15276 58710 15852
rect 58652 15264 58710 15276
rect 58780 15852 58838 15864
rect 58780 15276 58792 15852
rect 58826 15276 58838 15852
rect 58780 15264 58838 15276
rect 58892 15852 58950 15864
rect 58892 15276 58904 15852
rect 58938 15276 58950 15852
rect 58892 15264 58950 15276
rect 59020 15852 59078 15864
rect 59020 15276 59032 15852
rect 59066 15276 59078 15852
rect 59020 15264 59078 15276
rect 59132 15852 59190 15864
rect 59132 15276 59144 15852
rect 59178 15276 59190 15852
rect 59132 15264 59190 15276
rect 59260 15852 59318 15864
rect 59260 15276 59272 15852
rect 59306 15276 59318 15852
rect 59260 15264 59318 15276
rect 59372 15852 59430 15864
rect 59372 15276 59384 15852
rect 59418 15276 59430 15852
rect 59372 15264 59430 15276
rect 59500 15852 59558 15864
rect 59500 15276 59512 15852
rect 59546 15276 59558 15852
rect 59500 15264 59558 15276
rect 59612 15852 59670 15864
rect 59612 15276 59624 15852
rect 59658 15276 59670 15852
rect 59612 15264 59670 15276
rect 59740 15852 59798 15864
rect 59740 15276 59752 15852
rect 59786 15276 59798 15852
rect 59740 15264 59798 15276
rect 59852 15852 59910 15864
rect 59852 15276 59864 15852
rect 59898 15276 59910 15852
rect 59852 15264 59910 15276
rect 59980 15852 60038 15864
rect 59980 15276 59992 15852
rect 60026 15276 60038 15852
rect 59980 15264 60038 15276
rect 60092 15852 60150 15864
rect 60092 15276 60104 15852
rect 60138 15276 60150 15852
rect 60092 15264 60150 15276
rect 60220 15852 60278 15864
rect 60220 15276 60232 15852
rect 60266 15276 60278 15852
rect 60220 15264 60278 15276
rect 60332 15852 60390 15864
rect 60332 15276 60344 15852
rect 60378 15276 60390 15852
rect 60332 15264 60390 15276
rect 60460 15852 60518 15864
rect 60460 15276 60472 15852
rect 60506 15276 60518 15852
rect 60460 15264 60518 15276
rect 60572 15852 60630 15864
rect 60572 15276 60584 15852
rect 60618 15276 60630 15852
rect 60572 15264 60630 15276
rect 60700 15852 60758 15864
rect 60700 15276 60712 15852
rect 60746 15276 60758 15852
rect 60700 15264 60758 15276
rect 60812 15852 60870 15864
rect 60812 15276 60824 15852
rect 60858 15276 60870 15852
rect 60812 15264 60870 15276
rect 60940 15852 60998 15864
rect 60940 15276 60952 15852
rect 60986 15276 60998 15852
rect 60940 15264 60998 15276
rect 61052 15852 61110 15864
rect 61052 15276 61064 15852
rect 61098 15276 61110 15852
rect 61052 15264 61110 15276
rect 61180 15852 61238 15864
rect 61180 15276 61192 15852
rect 61226 15276 61238 15852
rect 61180 15264 61238 15276
rect 61292 15852 61350 15864
rect 61292 15276 61304 15852
rect 61338 15276 61350 15852
rect 61292 15264 61350 15276
rect 61420 15852 61478 15864
rect 61420 15276 61432 15852
rect 61466 15276 61478 15852
rect 61420 15264 61478 15276
rect 61532 15852 61590 15864
rect 61532 15276 61544 15852
rect 61578 15276 61590 15852
rect 61532 15264 61590 15276
rect 61660 15852 61718 15864
rect 61660 15276 61672 15852
rect 61706 15276 61718 15852
rect 61660 15264 61718 15276
rect 61772 15852 61830 15864
rect 61772 15276 61784 15852
rect 61818 15276 61830 15852
rect 61772 15264 61830 15276
rect 61900 15852 61958 15864
rect 61900 15276 61912 15852
rect 61946 15276 61958 15852
rect 61900 15264 61958 15276
rect 62012 15852 62070 15864
rect 62012 15276 62024 15852
rect 62058 15276 62070 15852
rect 62012 15264 62070 15276
rect 62140 15852 62198 15864
rect 62140 15276 62152 15852
rect 62186 15276 62198 15852
rect 62140 15264 62198 15276
rect 56972 3948 57030 3960
rect 56972 3372 56984 3948
rect 57018 3372 57030 3948
rect 56972 3360 57030 3372
rect 57100 3948 57158 3960
rect 57100 3372 57112 3948
rect 57146 3372 57158 3948
rect 57100 3360 57158 3372
rect 57212 3948 57270 3960
rect 57212 3372 57224 3948
rect 57258 3372 57270 3948
rect 57212 3360 57270 3372
rect 57340 3948 57398 3960
rect 57340 3372 57352 3948
rect 57386 3372 57398 3948
rect 57340 3360 57398 3372
rect 57452 3948 57510 3960
rect 57452 3372 57464 3948
rect 57498 3372 57510 3948
rect 57452 3360 57510 3372
rect 57580 3948 57638 3960
rect 57580 3372 57592 3948
rect 57626 3372 57638 3948
rect 57580 3360 57638 3372
rect 57692 3948 57750 3960
rect 57692 3372 57704 3948
rect 57738 3372 57750 3948
rect 57692 3360 57750 3372
rect 57820 3948 57878 3960
rect 57820 3372 57832 3948
rect 57866 3372 57878 3948
rect 57820 3360 57878 3372
rect 56972 3140 57030 3152
rect 56972 2564 56984 3140
rect 57018 2564 57030 3140
rect 56972 2552 57030 2564
rect 57100 3140 57158 3152
rect 57100 2564 57112 3140
rect 57146 2564 57158 3140
rect 57100 2552 57158 2564
rect 57212 3140 57270 3152
rect 57212 2564 57224 3140
rect 57258 2564 57270 3140
rect 57212 2552 57270 2564
rect 57340 3140 57398 3152
rect 57340 2564 57352 3140
rect 57386 2564 57398 3140
rect 57340 2552 57398 2564
rect 57452 3140 57510 3152
rect 57452 2564 57464 3140
rect 57498 2564 57510 3140
rect 57452 2552 57510 2564
rect 57580 3140 57638 3152
rect 57580 2564 57592 3140
rect 57626 2564 57638 3140
rect 57580 2552 57638 2564
rect 57692 3140 57750 3152
rect 57692 2564 57704 3140
rect 57738 2564 57750 3140
rect 57692 2552 57750 2564
rect 57820 3140 57878 3152
rect 57820 2564 57832 3140
rect 57866 2564 57878 3140
rect 57820 2552 57878 2564
<< pdiff >>
rect 43348 12586 43406 12598
rect 43348 11810 43360 12586
rect 43394 11810 43406 12586
rect 43348 11798 43406 11810
rect 43806 12586 43864 12598
rect 43806 11810 43818 12586
rect 43852 11810 43864 12586
rect 43806 11798 43864 11810
rect 43936 12586 43994 12598
rect 43936 11810 43948 12586
rect 43982 11810 43994 12586
rect 43936 11798 43994 11810
rect 44394 12586 44452 12598
rect 44394 11810 44406 12586
rect 44440 11810 44452 12586
rect 44394 11798 44452 11810
rect 44524 12586 44582 12598
rect 44524 11810 44536 12586
rect 44570 11810 44582 12586
rect 44524 11798 44582 11810
rect 44982 12586 45040 12598
rect 44982 11810 44994 12586
rect 45028 11810 45040 12586
rect 44982 11798 45040 11810
rect 45112 12586 45170 12598
rect 45112 11810 45124 12586
rect 45158 11810 45170 12586
rect 45112 11798 45170 11810
rect 45570 12586 45628 12598
rect 45570 11810 45582 12586
rect 45616 11810 45628 12586
rect 45570 11798 45628 11810
rect 45700 12586 45758 12598
rect 45700 11810 45712 12586
rect 45746 11810 45758 12586
rect 45700 11798 45758 11810
rect 46158 12586 46216 12598
rect 46158 11810 46170 12586
rect 46204 11810 46216 12586
rect 46158 11798 46216 11810
rect 46288 12586 46346 12598
rect 46288 11810 46300 12586
rect 46334 11810 46346 12586
rect 46288 11798 46346 11810
rect 46746 12586 46804 12598
rect 46746 11810 46758 12586
rect 46792 11810 46804 12586
rect 46746 11798 46804 11810
rect 46876 12586 46934 12598
rect 46876 11810 46888 12586
rect 46922 11810 46934 12586
rect 46876 11798 46934 11810
rect 47334 12586 47392 12598
rect 47334 11810 47346 12586
rect 47380 11810 47392 12586
rect 47334 11798 47392 11810
rect 47464 12586 47522 12598
rect 47464 11810 47476 12586
rect 47510 11810 47522 12586
rect 47464 11798 47522 11810
rect 47922 12586 47980 12598
rect 47922 11810 47934 12586
rect 47968 11810 47980 12586
rect 47922 11798 47980 11810
rect 48052 12586 48110 12598
rect 48052 11810 48064 12586
rect 48098 11810 48110 12586
rect 48052 11798 48110 11810
rect 48510 12586 48568 12598
rect 48510 11810 48522 12586
rect 48556 11810 48568 12586
rect 48510 11798 48568 11810
rect 48640 12586 48698 12598
rect 48640 11810 48652 12586
rect 48686 11810 48698 12586
rect 48640 11798 48698 11810
rect 49098 12586 49156 12598
rect 49098 11810 49110 12586
rect 49144 11810 49156 12586
rect 49098 11798 49156 11810
rect 49228 12586 49286 12598
rect 49228 11810 49240 12586
rect 49274 11810 49286 12586
rect 49228 11798 49286 11810
rect 49686 12586 49744 12598
rect 49686 11810 49698 12586
rect 49732 11810 49744 12586
rect 49686 11798 49744 11810
rect 49816 12586 49874 12598
rect 49816 11810 49828 12586
rect 49862 11810 49874 12586
rect 49816 11798 49874 11810
rect 50274 12586 50332 12598
rect 50274 11810 50286 12586
rect 50320 11810 50332 12586
rect 50274 11798 50332 11810
rect 50404 12586 50462 12598
rect 50404 11810 50416 12586
rect 50450 11810 50462 12586
rect 50404 11798 50462 11810
rect 50862 12586 50920 12598
rect 50862 11810 50874 12586
rect 50908 11810 50920 12586
rect 50862 11798 50920 11810
rect 50992 12586 51050 12598
rect 50992 11810 51004 12586
rect 51038 11810 51050 12586
rect 50992 11798 51050 11810
rect 51450 12586 51508 12598
rect 51450 11810 51462 12586
rect 51496 11810 51508 12586
rect 51450 11798 51508 11810
rect 51580 12586 51638 12598
rect 51580 11810 51592 12586
rect 51626 11810 51638 12586
rect 51580 11798 51638 11810
rect 52038 12586 52096 12598
rect 52038 11810 52050 12586
rect 52084 11810 52096 12586
rect 52038 11798 52096 11810
rect 52168 12586 52226 12598
rect 52168 11810 52180 12586
rect 52214 11810 52226 12586
rect 52168 11798 52226 11810
rect 52626 12586 52684 12598
rect 52626 11810 52638 12586
rect 52672 11810 52684 12586
rect 52626 11798 52684 11810
rect 52756 12586 52814 12598
rect 52756 11810 52768 12586
rect 52802 11810 52814 12586
rect 52756 11798 52814 11810
rect 53214 12586 53272 12598
rect 53214 11810 53226 12586
rect 53260 11810 53272 12586
rect 53214 11798 53272 11810
rect 53344 12586 53402 12598
rect 53344 11810 53356 12586
rect 53390 11810 53402 12586
rect 53344 11798 53402 11810
rect 53802 12586 53860 12598
rect 53802 11810 53814 12586
rect 53848 11810 53860 12586
rect 53802 11798 53860 11810
rect 53932 12586 53990 12598
rect 53932 11810 53944 12586
rect 53978 11810 53990 12586
rect 53932 11798 53990 11810
rect 54390 12586 54448 12598
rect 54390 11810 54402 12586
rect 54436 11810 54448 12586
rect 54390 11798 54448 11810
rect 54520 12586 54578 12598
rect 54520 11810 54532 12586
rect 54566 11810 54578 12586
rect 54520 11798 54578 11810
rect 54978 12586 55036 12598
rect 54978 11810 54990 12586
rect 55024 11810 55036 12586
rect 54978 11798 55036 11810
rect 55108 12586 55166 12598
rect 55108 11810 55120 12586
rect 55154 11810 55166 12586
rect 55108 11798 55166 11810
rect 55566 12586 55624 12598
rect 55566 11810 55578 12586
rect 55612 11810 55624 12586
rect 55566 11798 55624 11810
rect 55696 12586 55754 12598
rect 55696 11810 55708 12586
rect 55742 11810 55754 12586
rect 55696 11798 55754 11810
rect 56154 12586 56212 12598
rect 56154 11810 56166 12586
rect 56200 11810 56212 12586
rect 56154 11798 56212 11810
rect 56284 12586 56342 12598
rect 56284 11810 56296 12586
rect 56330 11810 56342 12586
rect 56284 11798 56342 11810
rect 56742 12586 56800 12598
rect 56742 11810 56754 12586
rect 56788 11810 56800 12586
rect 56742 11798 56800 11810
rect 56872 12586 56930 12598
rect 56872 11810 56884 12586
rect 56918 11810 56930 12586
rect 56872 11798 56930 11810
rect 57330 12586 57388 12598
rect 57330 11810 57342 12586
rect 57376 11810 57388 12586
rect 57330 11798 57388 11810
rect 57460 12586 57518 12598
rect 57460 11810 57472 12586
rect 57506 11810 57518 12586
rect 57460 11798 57518 11810
rect 57918 12586 57976 12598
rect 57918 11810 57930 12586
rect 57964 11810 57976 12586
rect 57918 11798 57976 11810
rect 58048 12586 58106 12598
rect 58048 11810 58060 12586
rect 58094 11810 58106 12586
rect 58048 11798 58106 11810
rect 58506 12586 58564 12598
rect 58506 11810 58518 12586
rect 58552 11810 58564 12586
rect 58506 11798 58564 11810
rect 58636 12586 58694 12598
rect 58636 11810 58648 12586
rect 58682 11810 58694 12586
rect 58636 11798 58694 11810
rect 59094 12586 59152 12598
rect 59094 11810 59106 12586
rect 59140 11810 59152 12586
rect 59094 11798 59152 11810
rect 59224 12586 59282 12598
rect 59224 11810 59236 12586
rect 59270 11810 59282 12586
rect 59224 11798 59282 11810
rect 59682 12586 59740 12598
rect 59682 11810 59694 12586
rect 59728 11810 59740 12586
rect 59682 11798 59740 11810
rect 59812 12586 59870 12598
rect 59812 11810 59824 12586
rect 59858 11810 59870 12586
rect 59812 11798 59870 11810
rect 60270 12586 60328 12598
rect 60270 11810 60282 12586
rect 60316 11810 60328 12586
rect 60270 11798 60328 11810
rect 60400 12586 60458 12598
rect 60400 11810 60412 12586
rect 60446 11810 60458 12586
rect 60400 11798 60458 11810
rect 60858 12586 60916 12598
rect 60858 11810 60870 12586
rect 60904 11810 60916 12586
rect 60858 11798 60916 11810
rect 60988 12586 61046 12598
rect 60988 11810 61000 12586
rect 61034 11810 61046 12586
rect 60988 11798 61046 11810
rect 61446 12586 61504 12598
rect 61446 11810 61458 12586
rect 61492 11810 61504 12586
rect 61446 11798 61504 11810
rect 61576 12586 61634 12598
rect 61576 11810 61588 12586
rect 61622 11810 61634 12586
rect 61576 11798 61634 11810
rect 62034 12586 62092 12598
rect 62034 11810 62046 12586
rect 62080 11810 62092 12586
rect 62034 11798 62092 11810
rect 62164 12586 62222 12598
rect 62164 11810 62176 12586
rect 62210 11810 62222 12586
rect 62164 11798 62222 11810
rect 62622 12586 62680 12598
rect 62622 11810 62634 12586
rect 62668 11810 62680 12586
rect 62622 11798 62680 11810
rect 62752 12586 62810 12598
rect 62752 11810 62764 12586
rect 62798 11810 62810 12586
rect 62752 11798 62810 11810
rect 63210 12586 63268 12598
rect 63210 11810 63222 12586
rect 63256 11810 63268 12586
rect 63210 11798 63268 11810
rect 63340 12586 63398 12598
rect 63340 11810 63352 12586
rect 63386 11810 63398 12586
rect 63340 11798 63398 11810
rect 63798 12586 63856 12598
rect 63798 11810 63810 12586
rect 63844 11810 63856 12586
rect 63798 11798 63856 11810
rect 63928 12586 63986 12598
rect 63928 11810 63940 12586
rect 63974 11810 63986 12586
rect 63928 11798 63986 11810
rect 64386 12586 64444 12598
rect 64386 11810 64398 12586
rect 64432 11810 64444 12586
rect 64386 11798 64444 11810
rect 64516 12586 64574 12598
rect 64516 11810 64528 12586
rect 64562 11810 64574 12586
rect 64516 11798 64574 11810
rect 64974 12586 65032 12598
rect 64974 11810 64986 12586
rect 65020 11810 65032 12586
rect 64974 11798 65032 11810
rect 65104 12586 65162 12598
rect 65104 11810 65116 12586
rect 65150 11810 65162 12586
rect 65104 11798 65162 11810
rect 65562 12586 65620 12598
rect 65562 11810 65574 12586
rect 65608 11810 65620 12586
rect 65562 11798 65620 11810
rect 65692 12586 65750 12598
rect 65692 11810 65704 12586
rect 65738 11810 65750 12586
rect 65692 11798 65750 11810
rect 66150 12586 66208 12598
rect 66150 11810 66162 12586
rect 66196 11810 66208 12586
rect 66150 11798 66208 11810
rect 66280 12586 66338 12598
rect 66280 11810 66292 12586
rect 66326 11810 66338 12586
rect 66280 11798 66338 11810
rect 66738 12586 66796 12598
rect 66738 11810 66750 12586
rect 66784 11810 66796 12586
rect 66738 11798 66796 11810
rect 66868 12586 66926 12598
rect 66868 11810 66880 12586
rect 66914 11810 66926 12586
rect 66868 11798 66926 11810
rect 67326 12586 67384 12598
rect 67326 11810 67338 12586
rect 67372 11810 67384 12586
rect 67326 11798 67384 11810
rect 67456 12586 67514 12598
rect 67456 11810 67468 12586
rect 67502 11810 67514 12586
rect 67456 11798 67514 11810
rect 67914 12586 67972 12598
rect 67914 11810 67926 12586
rect 67960 11810 67972 12586
rect 67914 11798 67972 11810
rect 68044 12586 68102 12598
rect 68044 11810 68056 12586
rect 68090 11810 68102 12586
rect 68044 11798 68102 11810
rect 68502 12586 68560 12598
rect 68502 11810 68514 12586
rect 68548 11810 68560 12586
rect 68502 11798 68560 11810
rect 68632 12586 68690 12598
rect 68632 11810 68644 12586
rect 68678 11810 68690 12586
rect 68632 11798 68690 11810
rect 69090 12586 69148 12598
rect 69090 11810 69102 12586
rect 69136 11810 69148 12586
rect 69090 11798 69148 11810
rect 69220 12586 69278 12598
rect 69220 11810 69232 12586
rect 69266 11810 69278 12586
rect 69220 11798 69278 11810
rect 69678 12586 69736 12598
rect 69678 11810 69690 12586
rect 69724 11810 69736 12586
rect 69678 11798 69736 11810
rect 69808 12586 69866 12598
rect 69808 11810 69820 12586
rect 69854 11810 69866 12586
rect 69808 11798 69866 11810
rect 70266 12586 70324 12598
rect 70266 11810 70278 12586
rect 70312 11810 70324 12586
rect 70266 11798 70324 11810
rect 70396 12586 70454 12598
rect 70396 11810 70408 12586
rect 70442 11810 70454 12586
rect 70396 11798 70454 11810
rect 70854 12586 70912 12598
rect 70854 11810 70866 12586
rect 70900 11810 70912 12586
rect 70854 11798 70912 11810
rect 70984 12586 71042 12598
rect 70984 11810 70996 12586
rect 71030 11810 71042 12586
rect 70984 11798 71042 11810
rect 71442 12586 71500 12598
rect 71442 11810 71454 12586
rect 71488 11810 71500 12586
rect 71442 11798 71500 11810
rect 43348 11586 43406 11598
rect 43348 10810 43360 11586
rect 43394 10810 43406 11586
rect 43348 10798 43406 10810
rect 43806 11586 43864 11598
rect 43806 10810 43818 11586
rect 43852 10810 43864 11586
rect 43806 10798 43864 10810
rect 43936 11586 43994 11598
rect 43936 10810 43948 11586
rect 43982 10810 43994 11586
rect 43936 10798 43994 10810
rect 44394 11586 44452 11598
rect 44394 10810 44406 11586
rect 44440 10810 44452 11586
rect 44394 10798 44452 10810
rect 44524 11586 44582 11598
rect 44524 10810 44536 11586
rect 44570 10810 44582 11586
rect 44524 10798 44582 10810
rect 44982 11586 45040 11598
rect 44982 10810 44994 11586
rect 45028 10810 45040 11586
rect 44982 10798 45040 10810
rect 45112 11586 45170 11598
rect 45112 10810 45124 11586
rect 45158 10810 45170 11586
rect 45112 10798 45170 10810
rect 45570 11586 45628 11598
rect 45570 10810 45582 11586
rect 45616 10810 45628 11586
rect 45570 10798 45628 10810
rect 45700 11586 45758 11598
rect 45700 10810 45712 11586
rect 45746 10810 45758 11586
rect 45700 10798 45758 10810
rect 46158 11586 46216 11598
rect 46158 10810 46170 11586
rect 46204 10810 46216 11586
rect 46158 10798 46216 10810
rect 46288 11586 46346 11598
rect 46288 10810 46300 11586
rect 46334 10810 46346 11586
rect 46288 10798 46346 10810
rect 46746 11586 46804 11598
rect 46746 10810 46758 11586
rect 46792 10810 46804 11586
rect 46746 10798 46804 10810
rect 46876 11586 46934 11598
rect 46876 10810 46888 11586
rect 46922 10810 46934 11586
rect 46876 10798 46934 10810
rect 47334 11586 47392 11598
rect 47334 10810 47346 11586
rect 47380 10810 47392 11586
rect 47334 10798 47392 10810
rect 47464 11586 47522 11598
rect 47464 10810 47476 11586
rect 47510 10810 47522 11586
rect 47464 10798 47522 10810
rect 47922 11586 47980 11598
rect 47922 10810 47934 11586
rect 47968 10810 47980 11586
rect 47922 10798 47980 10810
rect 48052 11586 48110 11598
rect 48052 10810 48064 11586
rect 48098 10810 48110 11586
rect 48052 10798 48110 10810
rect 48510 11586 48568 11598
rect 48510 10810 48522 11586
rect 48556 10810 48568 11586
rect 48510 10798 48568 10810
rect 48640 11586 48698 11598
rect 48640 10810 48652 11586
rect 48686 10810 48698 11586
rect 48640 10798 48698 10810
rect 49098 11586 49156 11598
rect 49098 10810 49110 11586
rect 49144 10810 49156 11586
rect 49098 10798 49156 10810
rect 49228 11586 49286 11598
rect 49228 10810 49240 11586
rect 49274 10810 49286 11586
rect 49228 10798 49286 10810
rect 49686 11586 49744 11598
rect 49686 10810 49698 11586
rect 49732 10810 49744 11586
rect 49686 10798 49744 10810
rect 49816 11586 49874 11598
rect 49816 10810 49828 11586
rect 49862 10810 49874 11586
rect 49816 10798 49874 10810
rect 50274 11586 50332 11598
rect 50274 10810 50286 11586
rect 50320 10810 50332 11586
rect 50274 10798 50332 10810
rect 50404 11586 50462 11598
rect 50404 10810 50416 11586
rect 50450 10810 50462 11586
rect 50404 10798 50462 10810
rect 50862 11586 50920 11598
rect 50862 10810 50874 11586
rect 50908 10810 50920 11586
rect 50862 10798 50920 10810
rect 50992 11586 51050 11598
rect 50992 10810 51004 11586
rect 51038 10810 51050 11586
rect 50992 10798 51050 10810
rect 51450 11586 51508 11598
rect 51450 10810 51462 11586
rect 51496 10810 51508 11586
rect 51450 10798 51508 10810
rect 51580 11586 51638 11598
rect 51580 10810 51592 11586
rect 51626 10810 51638 11586
rect 51580 10798 51638 10810
rect 52038 11586 52096 11598
rect 52038 10810 52050 11586
rect 52084 10810 52096 11586
rect 52038 10798 52096 10810
rect 52168 11586 52226 11598
rect 52168 10810 52180 11586
rect 52214 10810 52226 11586
rect 52168 10798 52226 10810
rect 52626 11586 52684 11598
rect 52626 10810 52638 11586
rect 52672 10810 52684 11586
rect 52626 10798 52684 10810
rect 52756 11586 52814 11598
rect 52756 10810 52768 11586
rect 52802 10810 52814 11586
rect 52756 10798 52814 10810
rect 53214 11586 53272 11598
rect 53214 10810 53226 11586
rect 53260 10810 53272 11586
rect 53214 10798 53272 10810
rect 53344 11586 53402 11598
rect 53344 10810 53356 11586
rect 53390 10810 53402 11586
rect 53344 10798 53402 10810
rect 53802 11586 53860 11598
rect 53802 10810 53814 11586
rect 53848 10810 53860 11586
rect 53802 10798 53860 10810
rect 53932 11586 53990 11598
rect 53932 10810 53944 11586
rect 53978 10810 53990 11586
rect 53932 10798 53990 10810
rect 54390 11586 54448 11598
rect 54390 10810 54402 11586
rect 54436 10810 54448 11586
rect 54390 10798 54448 10810
rect 54520 11586 54578 11598
rect 54520 10810 54532 11586
rect 54566 10810 54578 11586
rect 54520 10798 54578 10810
rect 54978 11586 55036 11598
rect 54978 10810 54990 11586
rect 55024 10810 55036 11586
rect 54978 10798 55036 10810
rect 55108 11586 55166 11598
rect 55108 10810 55120 11586
rect 55154 10810 55166 11586
rect 55108 10798 55166 10810
rect 55566 11586 55624 11598
rect 55566 10810 55578 11586
rect 55612 10810 55624 11586
rect 55566 10798 55624 10810
rect 55696 11586 55754 11598
rect 55696 10810 55708 11586
rect 55742 10810 55754 11586
rect 55696 10798 55754 10810
rect 56154 11586 56212 11598
rect 56154 10810 56166 11586
rect 56200 10810 56212 11586
rect 56154 10798 56212 10810
rect 56284 11586 56342 11598
rect 56284 10810 56296 11586
rect 56330 10810 56342 11586
rect 56284 10798 56342 10810
rect 56742 11586 56800 11598
rect 56742 10810 56754 11586
rect 56788 10810 56800 11586
rect 56742 10798 56800 10810
rect 56872 11586 56930 11598
rect 56872 10810 56884 11586
rect 56918 10810 56930 11586
rect 56872 10798 56930 10810
rect 57330 11586 57388 11598
rect 57330 10810 57342 11586
rect 57376 10810 57388 11586
rect 57330 10798 57388 10810
rect 57460 11586 57518 11598
rect 57460 10810 57472 11586
rect 57506 10810 57518 11586
rect 57460 10798 57518 10810
rect 57918 11586 57976 11598
rect 57918 10810 57930 11586
rect 57964 10810 57976 11586
rect 57918 10798 57976 10810
rect 58048 11586 58106 11598
rect 58048 10810 58060 11586
rect 58094 10810 58106 11586
rect 58048 10798 58106 10810
rect 58506 11586 58564 11598
rect 58506 10810 58518 11586
rect 58552 10810 58564 11586
rect 58506 10798 58564 10810
rect 58636 11586 58694 11598
rect 58636 10810 58648 11586
rect 58682 10810 58694 11586
rect 58636 10798 58694 10810
rect 59094 11586 59152 11598
rect 59094 10810 59106 11586
rect 59140 10810 59152 11586
rect 59094 10798 59152 10810
rect 59224 11586 59282 11598
rect 59224 10810 59236 11586
rect 59270 10810 59282 11586
rect 59224 10798 59282 10810
rect 59682 11586 59740 11598
rect 59682 10810 59694 11586
rect 59728 10810 59740 11586
rect 59682 10798 59740 10810
rect 59812 11586 59870 11598
rect 59812 10810 59824 11586
rect 59858 10810 59870 11586
rect 59812 10798 59870 10810
rect 60270 11586 60328 11598
rect 60270 10810 60282 11586
rect 60316 10810 60328 11586
rect 60270 10798 60328 10810
rect 60400 11586 60458 11598
rect 60400 10810 60412 11586
rect 60446 10810 60458 11586
rect 60400 10798 60458 10810
rect 60858 11586 60916 11598
rect 60858 10810 60870 11586
rect 60904 10810 60916 11586
rect 60858 10798 60916 10810
rect 60988 11586 61046 11598
rect 60988 10810 61000 11586
rect 61034 10810 61046 11586
rect 60988 10798 61046 10810
rect 61446 11586 61504 11598
rect 61446 10810 61458 11586
rect 61492 10810 61504 11586
rect 61446 10798 61504 10810
rect 61576 11586 61634 11598
rect 61576 10810 61588 11586
rect 61622 10810 61634 11586
rect 61576 10798 61634 10810
rect 62034 11586 62092 11598
rect 62034 10810 62046 11586
rect 62080 10810 62092 11586
rect 62034 10798 62092 10810
rect 62164 11586 62222 11598
rect 62164 10810 62176 11586
rect 62210 10810 62222 11586
rect 62164 10798 62222 10810
rect 62622 11586 62680 11598
rect 62622 10810 62634 11586
rect 62668 10810 62680 11586
rect 62622 10798 62680 10810
rect 62752 11586 62810 11598
rect 62752 10810 62764 11586
rect 62798 10810 62810 11586
rect 62752 10798 62810 10810
rect 63210 11586 63268 11598
rect 63210 10810 63222 11586
rect 63256 10810 63268 11586
rect 63210 10798 63268 10810
rect 63340 11586 63398 11598
rect 63340 10810 63352 11586
rect 63386 10810 63398 11586
rect 63340 10798 63398 10810
rect 63798 11586 63856 11598
rect 63798 10810 63810 11586
rect 63844 10810 63856 11586
rect 63798 10798 63856 10810
rect 63928 11586 63986 11598
rect 63928 10810 63940 11586
rect 63974 10810 63986 11586
rect 63928 10798 63986 10810
rect 64386 11586 64444 11598
rect 64386 10810 64398 11586
rect 64432 10810 64444 11586
rect 64386 10798 64444 10810
rect 64516 11586 64574 11598
rect 64516 10810 64528 11586
rect 64562 10810 64574 11586
rect 64516 10798 64574 10810
rect 64974 11586 65032 11598
rect 64974 10810 64986 11586
rect 65020 10810 65032 11586
rect 64974 10798 65032 10810
rect 65104 11586 65162 11598
rect 65104 10810 65116 11586
rect 65150 10810 65162 11586
rect 65104 10798 65162 10810
rect 65562 11586 65620 11598
rect 65562 10810 65574 11586
rect 65608 10810 65620 11586
rect 65562 10798 65620 10810
rect 65692 11586 65750 11598
rect 65692 10810 65704 11586
rect 65738 10810 65750 11586
rect 65692 10798 65750 10810
rect 66150 11586 66208 11598
rect 66150 10810 66162 11586
rect 66196 10810 66208 11586
rect 66150 10798 66208 10810
rect 66280 11586 66338 11598
rect 66280 10810 66292 11586
rect 66326 10810 66338 11586
rect 66280 10798 66338 10810
rect 66738 11586 66796 11598
rect 66738 10810 66750 11586
rect 66784 10810 66796 11586
rect 66738 10798 66796 10810
rect 66868 11586 66926 11598
rect 66868 10810 66880 11586
rect 66914 10810 66926 11586
rect 66868 10798 66926 10810
rect 67326 11586 67384 11598
rect 67326 10810 67338 11586
rect 67372 10810 67384 11586
rect 67326 10798 67384 10810
rect 67456 11586 67514 11598
rect 67456 10810 67468 11586
rect 67502 10810 67514 11586
rect 67456 10798 67514 10810
rect 67914 11586 67972 11598
rect 67914 10810 67926 11586
rect 67960 10810 67972 11586
rect 67914 10798 67972 10810
rect 68044 11586 68102 11598
rect 68044 10810 68056 11586
rect 68090 10810 68102 11586
rect 68044 10798 68102 10810
rect 68502 11586 68560 11598
rect 68502 10810 68514 11586
rect 68548 10810 68560 11586
rect 68502 10798 68560 10810
rect 68632 11586 68690 11598
rect 68632 10810 68644 11586
rect 68678 10810 68690 11586
rect 68632 10798 68690 10810
rect 69090 11586 69148 11598
rect 69090 10810 69102 11586
rect 69136 10810 69148 11586
rect 69090 10798 69148 10810
rect 69220 11586 69278 11598
rect 69220 10810 69232 11586
rect 69266 10810 69278 11586
rect 69220 10798 69278 10810
rect 69678 11586 69736 11598
rect 69678 10810 69690 11586
rect 69724 10810 69736 11586
rect 69678 10798 69736 10810
rect 69808 11586 69866 11598
rect 69808 10810 69820 11586
rect 69854 10810 69866 11586
rect 69808 10798 69866 10810
rect 70266 11586 70324 11598
rect 70266 10810 70278 11586
rect 70312 10810 70324 11586
rect 70266 10798 70324 10810
rect 70396 11586 70454 11598
rect 70396 10810 70408 11586
rect 70442 10810 70454 11586
rect 70396 10798 70454 10810
rect 70854 11586 70912 11598
rect 70854 10810 70866 11586
rect 70900 10810 70912 11586
rect 70854 10798 70912 10810
rect 70984 11586 71042 11598
rect 70984 10810 70996 11586
rect 71030 10810 71042 11586
rect 70984 10798 71042 10810
rect 71442 11586 71500 11598
rect 71442 10810 71454 11586
rect 71488 10810 71500 11586
rect 71442 10798 71500 10810
rect 43348 10586 43406 10598
rect 43348 9810 43360 10586
rect 43394 9810 43406 10586
rect 43348 9798 43406 9810
rect 43806 10586 43864 10598
rect 43806 9810 43818 10586
rect 43852 9810 43864 10586
rect 43806 9798 43864 9810
rect 43936 10586 43994 10598
rect 43936 9810 43948 10586
rect 43982 9810 43994 10586
rect 43936 9798 43994 9810
rect 44394 10586 44452 10598
rect 44394 9810 44406 10586
rect 44440 9810 44452 10586
rect 44394 9798 44452 9810
rect 44524 10586 44582 10598
rect 44524 9810 44536 10586
rect 44570 9810 44582 10586
rect 44524 9798 44582 9810
rect 44982 10586 45040 10598
rect 44982 9810 44994 10586
rect 45028 9810 45040 10586
rect 44982 9798 45040 9810
rect 45112 10586 45170 10598
rect 45112 9810 45124 10586
rect 45158 9810 45170 10586
rect 45112 9798 45170 9810
rect 45570 10586 45628 10598
rect 45570 9810 45582 10586
rect 45616 9810 45628 10586
rect 45570 9798 45628 9810
rect 45700 10586 45758 10598
rect 45700 9810 45712 10586
rect 45746 9810 45758 10586
rect 45700 9798 45758 9810
rect 46158 10586 46216 10598
rect 46158 9810 46170 10586
rect 46204 9810 46216 10586
rect 46158 9798 46216 9810
rect 46288 10586 46346 10598
rect 46288 9810 46300 10586
rect 46334 9810 46346 10586
rect 46288 9798 46346 9810
rect 46746 10586 46804 10598
rect 46746 9810 46758 10586
rect 46792 9810 46804 10586
rect 46746 9798 46804 9810
rect 46876 10586 46934 10598
rect 46876 9810 46888 10586
rect 46922 9810 46934 10586
rect 46876 9798 46934 9810
rect 47334 10586 47392 10598
rect 47334 9810 47346 10586
rect 47380 9810 47392 10586
rect 47334 9798 47392 9810
rect 47464 10586 47522 10598
rect 47464 9810 47476 10586
rect 47510 9810 47522 10586
rect 47464 9798 47522 9810
rect 47922 10586 47980 10598
rect 47922 9810 47934 10586
rect 47968 9810 47980 10586
rect 47922 9798 47980 9810
rect 48052 10586 48110 10598
rect 48052 9810 48064 10586
rect 48098 9810 48110 10586
rect 48052 9798 48110 9810
rect 48510 10586 48568 10598
rect 48510 9810 48522 10586
rect 48556 9810 48568 10586
rect 48510 9798 48568 9810
rect 48640 10586 48698 10598
rect 48640 9810 48652 10586
rect 48686 9810 48698 10586
rect 48640 9798 48698 9810
rect 49098 10586 49156 10598
rect 49098 9810 49110 10586
rect 49144 9810 49156 10586
rect 49098 9798 49156 9810
rect 49228 10586 49286 10598
rect 49228 9810 49240 10586
rect 49274 9810 49286 10586
rect 49228 9798 49286 9810
rect 49686 10586 49744 10598
rect 49686 9810 49698 10586
rect 49732 9810 49744 10586
rect 49686 9798 49744 9810
rect 49816 10586 49874 10598
rect 49816 9810 49828 10586
rect 49862 9810 49874 10586
rect 49816 9798 49874 9810
rect 50274 10586 50332 10598
rect 50274 9810 50286 10586
rect 50320 9810 50332 10586
rect 50274 9798 50332 9810
rect 50404 10586 50462 10598
rect 50404 9810 50416 10586
rect 50450 9810 50462 10586
rect 50404 9798 50462 9810
rect 50862 10586 50920 10598
rect 50862 9810 50874 10586
rect 50908 9810 50920 10586
rect 50862 9798 50920 9810
rect 50992 10586 51050 10598
rect 50992 9810 51004 10586
rect 51038 9810 51050 10586
rect 50992 9798 51050 9810
rect 51450 10586 51508 10598
rect 51450 9810 51462 10586
rect 51496 9810 51508 10586
rect 51450 9798 51508 9810
rect 51580 10586 51638 10598
rect 51580 9810 51592 10586
rect 51626 9810 51638 10586
rect 51580 9798 51638 9810
rect 52038 10586 52096 10598
rect 52038 9810 52050 10586
rect 52084 9810 52096 10586
rect 52038 9798 52096 9810
rect 52168 10586 52226 10598
rect 52168 9810 52180 10586
rect 52214 9810 52226 10586
rect 52168 9798 52226 9810
rect 52626 10586 52684 10598
rect 52626 9810 52638 10586
rect 52672 9810 52684 10586
rect 52626 9798 52684 9810
rect 52756 10586 52814 10598
rect 52756 9810 52768 10586
rect 52802 9810 52814 10586
rect 52756 9798 52814 9810
rect 53214 10586 53272 10598
rect 53214 9810 53226 10586
rect 53260 9810 53272 10586
rect 53214 9798 53272 9810
rect 53344 10586 53402 10598
rect 53344 9810 53356 10586
rect 53390 9810 53402 10586
rect 53344 9798 53402 9810
rect 53802 10586 53860 10598
rect 53802 9810 53814 10586
rect 53848 9810 53860 10586
rect 53802 9798 53860 9810
rect 53932 10586 53990 10598
rect 53932 9810 53944 10586
rect 53978 9810 53990 10586
rect 53932 9798 53990 9810
rect 54390 10586 54448 10598
rect 54390 9810 54402 10586
rect 54436 9810 54448 10586
rect 54390 9798 54448 9810
rect 54520 10586 54578 10598
rect 54520 9810 54532 10586
rect 54566 9810 54578 10586
rect 54520 9798 54578 9810
rect 54978 10586 55036 10598
rect 54978 9810 54990 10586
rect 55024 9810 55036 10586
rect 54978 9798 55036 9810
rect 55108 10586 55166 10598
rect 55108 9810 55120 10586
rect 55154 9810 55166 10586
rect 55108 9798 55166 9810
rect 55566 10586 55624 10598
rect 55566 9810 55578 10586
rect 55612 9810 55624 10586
rect 55566 9798 55624 9810
rect 55696 10586 55754 10598
rect 55696 9810 55708 10586
rect 55742 9810 55754 10586
rect 55696 9798 55754 9810
rect 56154 10586 56212 10598
rect 56154 9810 56166 10586
rect 56200 9810 56212 10586
rect 56154 9798 56212 9810
rect 56284 10586 56342 10598
rect 56284 9810 56296 10586
rect 56330 9810 56342 10586
rect 56284 9798 56342 9810
rect 56742 10586 56800 10598
rect 56742 9810 56754 10586
rect 56788 9810 56800 10586
rect 56742 9798 56800 9810
rect 56872 10586 56930 10598
rect 56872 9810 56884 10586
rect 56918 9810 56930 10586
rect 56872 9798 56930 9810
rect 57330 10586 57388 10598
rect 57330 9810 57342 10586
rect 57376 9810 57388 10586
rect 57330 9798 57388 9810
rect 57460 10586 57518 10598
rect 57460 9810 57472 10586
rect 57506 9810 57518 10586
rect 57460 9798 57518 9810
rect 57918 10586 57976 10598
rect 57918 9810 57930 10586
rect 57964 9810 57976 10586
rect 57918 9798 57976 9810
rect 58048 10586 58106 10598
rect 58048 9810 58060 10586
rect 58094 9810 58106 10586
rect 58048 9798 58106 9810
rect 58506 10586 58564 10598
rect 58506 9810 58518 10586
rect 58552 9810 58564 10586
rect 58506 9798 58564 9810
rect 58636 10586 58694 10598
rect 58636 9810 58648 10586
rect 58682 9810 58694 10586
rect 58636 9798 58694 9810
rect 59094 10586 59152 10598
rect 59094 9810 59106 10586
rect 59140 9810 59152 10586
rect 59094 9798 59152 9810
rect 59224 10586 59282 10598
rect 59224 9810 59236 10586
rect 59270 9810 59282 10586
rect 59224 9798 59282 9810
rect 59682 10586 59740 10598
rect 59682 9810 59694 10586
rect 59728 9810 59740 10586
rect 59682 9798 59740 9810
rect 59812 10586 59870 10598
rect 59812 9810 59824 10586
rect 59858 9810 59870 10586
rect 59812 9798 59870 9810
rect 60270 10586 60328 10598
rect 60270 9810 60282 10586
rect 60316 9810 60328 10586
rect 60270 9798 60328 9810
rect 60400 10586 60458 10598
rect 60400 9810 60412 10586
rect 60446 9810 60458 10586
rect 60400 9798 60458 9810
rect 60858 10586 60916 10598
rect 60858 9810 60870 10586
rect 60904 9810 60916 10586
rect 60858 9798 60916 9810
rect 60988 10586 61046 10598
rect 60988 9810 61000 10586
rect 61034 9810 61046 10586
rect 60988 9798 61046 9810
rect 61446 10586 61504 10598
rect 61446 9810 61458 10586
rect 61492 9810 61504 10586
rect 61446 9798 61504 9810
rect 61576 10586 61634 10598
rect 61576 9810 61588 10586
rect 61622 9810 61634 10586
rect 61576 9798 61634 9810
rect 62034 10586 62092 10598
rect 62034 9810 62046 10586
rect 62080 9810 62092 10586
rect 62034 9798 62092 9810
rect 62164 10586 62222 10598
rect 62164 9810 62176 10586
rect 62210 9810 62222 10586
rect 62164 9798 62222 9810
rect 62622 10586 62680 10598
rect 62622 9810 62634 10586
rect 62668 9810 62680 10586
rect 62622 9798 62680 9810
rect 62752 10586 62810 10598
rect 62752 9810 62764 10586
rect 62798 9810 62810 10586
rect 62752 9798 62810 9810
rect 63210 10586 63268 10598
rect 63210 9810 63222 10586
rect 63256 9810 63268 10586
rect 63210 9798 63268 9810
rect 63340 10586 63398 10598
rect 63340 9810 63352 10586
rect 63386 9810 63398 10586
rect 63340 9798 63398 9810
rect 63798 10586 63856 10598
rect 63798 9810 63810 10586
rect 63844 9810 63856 10586
rect 63798 9798 63856 9810
rect 63928 10586 63986 10598
rect 63928 9810 63940 10586
rect 63974 9810 63986 10586
rect 63928 9798 63986 9810
rect 64386 10586 64444 10598
rect 64386 9810 64398 10586
rect 64432 9810 64444 10586
rect 64386 9798 64444 9810
rect 64516 10586 64574 10598
rect 64516 9810 64528 10586
rect 64562 9810 64574 10586
rect 64516 9798 64574 9810
rect 64974 10586 65032 10598
rect 64974 9810 64986 10586
rect 65020 9810 65032 10586
rect 64974 9798 65032 9810
rect 65104 10586 65162 10598
rect 65104 9810 65116 10586
rect 65150 9810 65162 10586
rect 65104 9798 65162 9810
rect 65562 10586 65620 10598
rect 65562 9810 65574 10586
rect 65608 9810 65620 10586
rect 65562 9798 65620 9810
rect 65692 10586 65750 10598
rect 65692 9810 65704 10586
rect 65738 9810 65750 10586
rect 65692 9798 65750 9810
rect 66150 10586 66208 10598
rect 66150 9810 66162 10586
rect 66196 9810 66208 10586
rect 66150 9798 66208 9810
rect 66280 10586 66338 10598
rect 66280 9810 66292 10586
rect 66326 9810 66338 10586
rect 66280 9798 66338 9810
rect 66738 10586 66796 10598
rect 66738 9810 66750 10586
rect 66784 9810 66796 10586
rect 66738 9798 66796 9810
rect 66868 10586 66926 10598
rect 66868 9810 66880 10586
rect 66914 9810 66926 10586
rect 66868 9798 66926 9810
rect 67326 10586 67384 10598
rect 67326 9810 67338 10586
rect 67372 9810 67384 10586
rect 67326 9798 67384 9810
rect 67456 10586 67514 10598
rect 67456 9810 67468 10586
rect 67502 9810 67514 10586
rect 67456 9798 67514 9810
rect 67914 10586 67972 10598
rect 67914 9810 67926 10586
rect 67960 9810 67972 10586
rect 67914 9798 67972 9810
rect 68044 10586 68102 10598
rect 68044 9810 68056 10586
rect 68090 9810 68102 10586
rect 68044 9798 68102 9810
rect 68502 10586 68560 10598
rect 68502 9810 68514 10586
rect 68548 9810 68560 10586
rect 68502 9798 68560 9810
rect 68632 10586 68690 10598
rect 68632 9810 68644 10586
rect 68678 9810 68690 10586
rect 68632 9798 68690 9810
rect 69090 10586 69148 10598
rect 69090 9810 69102 10586
rect 69136 9810 69148 10586
rect 69090 9798 69148 9810
rect 69220 10586 69278 10598
rect 69220 9810 69232 10586
rect 69266 9810 69278 10586
rect 69220 9798 69278 9810
rect 69678 10586 69736 10598
rect 69678 9810 69690 10586
rect 69724 9810 69736 10586
rect 69678 9798 69736 9810
rect 69808 10586 69866 10598
rect 69808 9810 69820 10586
rect 69854 9810 69866 10586
rect 69808 9798 69866 9810
rect 70266 10586 70324 10598
rect 70266 9810 70278 10586
rect 70312 9810 70324 10586
rect 70266 9798 70324 9810
rect 70396 10586 70454 10598
rect 70396 9810 70408 10586
rect 70442 9810 70454 10586
rect 70396 9798 70454 9810
rect 70854 10586 70912 10598
rect 70854 9810 70866 10586
rect 70900 9810 70912 10586
rect 70854 9798 70912 9810
rect 70984 10586 71042 10598
rect 70984 9810 70996 10586
rect 71030 9810 71042 10586
rect 70984 9798 71042 9810
rect 71442 10586 71500 10598
rect 71442 9810 71454 10586
rect 71488 9810 71500 10586
rect 71442 9798 71500 9810
rect 56400 8140 56458 8152
rect 56400 7364 56412 8140
rect 56446 7364 56458 8140
rect 56400 7352 56458 7364
rect 56528 8140 56586 8152
rect 56528 7364 56540 8140
rect 56574 7364 56586 8140
rect 56528 7352 56586 7364
rect 56666 8140 56724 8152
rect 56666 7364 56678 8140
rect 56712 7364 56724 8140
rect 56666 7352 56724 7364
rect 56794 8140 56852 8152
rect 56794 7364 56806 8140
rect 56840 7364 56852 8140
rect 56794 7352 56852 7364
rect 56932 8140 56990 8152
rect 56932 7364 56944 8140
rect 56978 7364 56990 8140
rect 56932 7352 56990 7364
rect 57060 8140 57118 8152
rect 57060 7364 57072 8140
rect 57106 7364 57118 8140
rect 57060 7352 57118 7364
rect 57198 8140 57256 8152
rect 57198 7364 57210 8140
rect 57244 7364 57256 8140
rect 57198 7352 57256 7364
rect 57326 8140 57384 8152
rect 57326 7364 57338 8140
rect 57372 7364 57384 8140
rect 57326 7352 57384 7364
rect 57464 8140 57522 8152
rect 57464 7364 57476 8140
rect 57510 7364 57522 8140
rect 57464 7352 57522 7364
rect 57592 8140 57650 8152
rect 57592 7364 57604 8140
rect 57638 7364 57650 8140
rect 57592 7352 57650 7364
rect 57730 8140 57788 8152
rect 57730 7364 57742 8140
rect 57776 7364 57788 8140
rect 57730 7352 57788 7364
rect 57858 8140 57916 8152
rect 57858 7364 57870 8140
rect 57904 7364 57916 8140
rect 57858 7352 57916 7364
rect 57996 8140 58054 8152
rect 57996 7364 58008 8140
rect 58042 7364 58054 8140
rect 57996 7352 58054 7364
rect 58124 8140 58182 8152
rect 58124 7364 58136 8140
rect 58170 7364 58182 8140
rect 58124 7352 58182 7364
rect 58262 8140 58320 8152
rect 58262 7364 58274 8140
rect 58308 7364 58320 8140
rect 58262 7352 58320 7364
rect 58390 8140 58448 8152
rect 58390 7364 58402 8140
rect 58436 7364 58448 8140
rect 58390 7352 58448 7364
rect 56400 7130 56458 7142
rect 56400 6354 56412 7130
rect 56446 6354 56458 7130
rect 56400 6342 56458 6354
rect 56528 7130 56586 7142
rect 56528 6354 56540 7130
rect 56574 6354 56586 7130
rect 56528 6342 56586 6354
rect 56666 7130 56724 7142
rect 56666 6354 56678 7130
rect 56712 6354 56724 7130
rect 56666 6342 56724 6354
rect 56794 7130 56852 7142
rect 56794 6354 56806 7130
rect 56840 6354 56852 7130
rect 56794 6342 56852 6354
rect 56932 7130 56990 7142
rect 56932 6354 56944 7130
rect 56978 6354 56990 7130
rect 56932 6342 56990 6354
rect 57060 7130 57118 7142
rect 57060 6354 57072 7130
rect 57106 6354 57118 7130
rect 57060 6342 57118 6354
rect 57198 7130 57256 7142
rect 57198 6354 57210 7130
rect 57244 6354 57256 7130
rect 57198 6342 57256 6354
rect 57326 7130 57384 7142
rect 57326 6354 57338 7130
rect 57372 6354 57384 7130
rect 57326 6342 57384 6354
rect 57464 7130 57522 7142
rect 57464 6354 57476 7130
rect 57510 6354 57522 7130
rect 57464 6342 57522 6354
rect 57592 7130 57650 7142
rect 57592 6354 57604 7130
rect 57638 6354 57650 7130
rect 57592 6342 57650 6354
rect 57730 7130 57788 7142
rect 57730 6354 57742 7130
rect 57776 6354 57788 7130
rect 57730 6342 57788 6354
rect 57858 7130 57916 7142
rect 57858 6354 57870 7130
rect 57904 6354 57916 7130
rect 57858 6342 57916 6354
rect 57996 7130 58054 7142
rect 57996 6354 58008 7130
rect 58042 6354 58054 7130
rect 57996 6342 58054 6354
rect 58124 7130 58182 7142
rect 58124 6354 58136 7130
rect 58170 6354 58182 7130
rect 58124 6342 58182 6354
rect 58262 7130 58320 7142
rect 58262 6354 58274 7130
rect 58308 6354 58320 7130
rect 58262 6342 58320 6354
rect 58390 7130 58448 7142
rect 58390 6354 58402 7130
rect 58436 6354 58448 7130
rect 58390 6342 58448 6354
rect 56400 6120 56458 6132
rect 56400 5344 56412 6120
rect 56446 5344 56458 6120
rect 56400 5332 56458 5344
rect 56528 6120 56586 6132
rect 56528 5344 56540 6120
rect 56574 5344 56586 6120
rect 56528 5332 56586 5344
rect 56666 6120 56724 6132
rect 56666 5344 56678 6120
rect 56712 5344 56724 6120
rect 56666 5332 56724 5344
rect 56794 6120 56852 6132
rect 56794 5344 56806 6120
rect 56840 5344 56852 6120
rect 56794 5332 56852 5344
rect 56932 6120 56990 6132
rect 56932 5344 56944 6120
rect 56978 5344 56990 6120
rect 56932 5332 56990 5344
rect 57060 6120 57118 6132
rect 57060 5344 57072 6120
rect 57106 5344 57118 6120
rect 57060 5332 57118 5344
rect 57198 6120 57256 6132
rect 57198 5344 57210 6120
rect 57244 5344 57256 6120
rect 57198 5332 57256 5344
rect 57326 6120 57384 6132
rect 57326 5344 57338 6120
rect 57372 5344 57384 6120
rect 57326 5332 57384 5344
rect 57464 6120 57522 6132
rect 57464 5344 57476 6120
rect 57510 5344 57522 6120
rect 57464 5332 57522 5344
rect 57592 6120 57650 6132
rect 57592 5344 57604 6120
rect 57638 5344 57650 6120
rect 57592 5332 57650 5344
rect 57730 6120 57788 6132
rect 57730 5344 57742 6120
rect 57776 5344 57788 6120
rect 57730 5332 57788 5344
rect 57858 6120 57916 6132
rect 57858 5344 57870 6120
rect 57904 5344 57916 6120
rect 57858 5332 57916 5344
rect 57996 6120 58054 6132
rect 57996 5344 58008 6120
rect 58042 5344 58054 6120
rect 57996 5332 58054 5344
rect 58124 6120 58182 6132
rect 58124 5344 58136 6120
rect 58170 5344 58182 6120
rect 58124 5332 58182 5344
rect 58262 6120 58320 6132
rect 58262 5344 58274 6120
rect 58308 5344 58320 6120
rect 58262 5332 58320 5344
rect 58390 6120 58448 6132
rect 58390 5344 58402 6120
rect 58436 5344 58448 6120
rect 58390 5332 58448 5344
<< ndiffc >>
rect 52664 16084 52698 16660
rect 52792 16084 52826 16660
rect 52904 16084 52938 16660
rect 53032 16084 53066 16660
rect 53144 16084 53178 16660
rect 53272 16084 53306 16660
rect 53384 16084 53418 16660
rect 53512 16084 53546 16660
rect 53624 16084 53658 16660
rect 53752 16084 53786 16660
rect 53864 16084 53898 16660
rect 53992 16084 54026 16660
rect 54104 16084 54138 16660
rect 54232 16084 54266 16660
rect 54344 16084 54378 16660
rect 54472 16084 54506 16660
rect 54584 16084 54618 16660
rect 54712 16084 54746 16660
rect 54824 16084 54858 16660
rect 54952 16084 54986 16660
rect 55064 16084 55098 16660
rect 55192 16084 55226 16660
rect 55304 16084 55338 16660
rect 55432 16084 55466 16660
rect 55544 16084 55578 16660
rect 55672 16084 55706 16660
rect 55784 16084 55818 16660
rect 55912 16084 55946 16660
rect 56024 16084 56058 16660
rect 56152 16084 56186 16660
rect 56264 16084 56298 16660
rect 56392 16084 56426 16660
rect 56504 16084 56538 16660
rect 56632 16084 56666 16660
rect 56744 16084 56778 16660
rect 56872 16084 56906 16660
rect 56984 16084 57018 16660
rect 57112 16084 57146 16660
rect 57224 16084 57258 16660
rect 57352 16084 57386 16660
rect 57464 16084 57498 16660
rect 57592 16084 57626 16660
rect 57704 16084 57738 16660
rect 57832 16084 57866 16660
rect 57944 16084 57978 16660
rect 58072 16084 58106 16660
rect 58184 16084 58218 16660
rect 58312 16084 58346 16660
rect 58424 16084 58458 16660
rect 58552 16084 58586 16660
rect 58664 16084 58698 16660
rect 58792 16084 58826 16660
rect 58904 16084 58938 16660
rect 59032 16084 59066 16660
rect 59144 16084 59178 16660
rect 59272 16084 59306 16660
rect 59384 16084 59418 16660
rect 59512 16084 59546 16660
rect 59624 16084 59658 16660
rect 59752 16084 59786 16660
rect 59864 16084 59898 16660
rect 59992 16084 60026 16660
rect 60104 16084 60138 16660
rect 60232 16084 60266 16660
rect 60344 16084 60378 16660
rect 60472 16084 60506 16660
rect 60584 16084 60618 16660
rect 60712 16084 60746 16660
rect 60824 16084 60858 16660
rect 60952 16084 60986 16660
rect 61064 16084 61098 16660
rect 61192 16084 61226 16660
rect 61304 16084 61338 16660
rect 61432 16084 61466 16660
rect 61544 16084 61578 16660
rect 61672 16084 61706 16660
rect 61784 16084 61818 16660
rect 61912 16084 61946 16660
rect 62024 16084 62058 16660
rect 62152 16084 62186 16660
rect 52664 15276 52698 15852
rect 52792 15276 52826 15852
rect 52904 15276 52938 15852
rect 53032 15276 53066 15852
rect 53144 15276 53178 15852
rect 53272 15276 53306 15852
rect 53384 15276 53418 15852
rect 53512 15276 53546 15852
rect 53624 15276 53658 15852
rect 53752 15276 53786 15852
rect 53864 15276 53898 15852
rect 53992 15276 54026 15852
rect 54104 15276 54138 15852
rect 54232 15276 54266 15852
rect 54344 15276 54378 15852
rect 54472 15276 54506 15852
rect 54584 15276 54618 15852
rect 54712 15276 54746 15852
rect 54824 15276 54858 15852
rect 54952 15276 54986 15852
rect 55064 15276 55098 15852
rect 55192 15276 55226 15852
rect 55304 15276 55338 15852
rect 55432 15276 55466 15852
rect 55544 15276 55578 15852
rect 55672 15276 55706 15852
rect 55784 15276 55818 15852
rect 55912 15276 55946 15852
rect 56024 15276 56058 15852
rect 56152 15276 56186 15852
rect 56264 15276 56298 15852
rect 56392 15276 56426 15852
rect 56504 15276 56538 15852
rect 56632 15276 56666 15852
rect 56744 15276 56778 15852
rect 56872 15276 56906 15852
rect 56984 15276 57018 15852
rect 57112 15276 57146 15852
rect 57224 15276 57258 15852
rect 57352 15276 57386 15852
rect 57464 15276 57498 15852
rect 57592 15276 57626 15852
rect 57704 15276 57738 15852
rect 57832 15276 57866 15852
rect 57944 15276 57978 15852
rect 58072 15276 58106 15852
rect 58184 15276 58218 15852
rect 58312 15276 58346 15852
rect 58424 15276 58458 15852
rect 58552 15276 58586 15852
rect 58664 15276 58698 15852
rect 58792 15276 58826 15852
rect 58904 15276 58938 15852
rect 59032 15276 59066 15852
rect 59144 15276 59178 15852
rect 59272 15276 59306 15852
rect 59384 15276 59418 15852
rect 59512 15276 59546 15852
rect 59624 15276 59658 15852
rect 59752 15276 59786 15852
rect 59864 15276 59898 15852
rect 59992 15276 60026 15852
rect 60104 15276 60138 15852
rect 60232 15276 60266 15852
rect 60344 15276 60378 15852
rect 60472 15276 60506 15852
rect 60584 15276 60618 15852
rect 60712 15276 60746 15852
rect 60824 15276 60858 15852
rect 60952 15276 60986 15852
rect 61064 15276 61098 15852
rect 61192 15276 61226 15852
rect 61304 15276 61338 15852
rect 61432 15276 61466 15852
rect 61544 15276 61578 15852
rect 61672 15276 61706 15852
rect 61784 15276 61818 15852
rect 61912 15276 61946 15852
rect 62024 15276 62058 15852
rect 62152 15276 62186 15852
rect 56984 3372 57018 3948
rect 57112 3372 57146 3948
rect 57224 3372 57258 3948
rect 57352 3372 57386 3948
rect 57464 3372 57498 3948
rect 57592 3372 57626 3948
rect 57704 3372 57738 3948
rect 57832 3372 57866 3948
rect 56984 2564 57018 3140
rect 57112 2564 57146 3140
rect 57224 2564 57258 3140
rect 57352 2564 57386 3140
rect 57464 2564 57498 3140
rect 57592 2564 57626 3140
rect 57704 2564 57738 3140
rect 57832 2564 57866 3140
<< pdiffc >>
rect 43360 11810 43394 12586
rect 43818 11810 43852 12586
rect 43948 11810 43982 12586
rect 44406 11810 44440 12586
rect 44536 11810 44570 12586
rect 44994 11810 45028 12586
rect 45124 11810 45158 12586
rect 45582 11810 45616 12586
rect 45712 11810 45746 12586
rect 46170 11810 46204 12586
rect 46300 11810 46334 12586
rect 46758 11810 46792 12586
rect 46888 11810 46922 12586
rect 47346 11810 47380 12586
rect 47476 11810 47510 12586
rect 47934 11810 47968 12586
rect 48064 11810 48098 12586
rect 48522 11810 48556 12586
rect 48652 11810 48686 12586
rect 49110 11810 49144 12586
rect 49240 11810 49274 12586
rect 49698 11810 49732 12586
rect 49828 11810 49862 12586
rect 50286 11810 50320 12586
rect 50416 11810 50450 12586
rect 50874 11810 50908 12586
rect 51004 11810 51038 12586
rect 51462 11810 51496 12586
rect 51592 11810 51626 12586
rect 52050 11810 52084 12586
rect 52180 11810 52214 12586
rect 52638 11810 52672 12586
rect 52768 11810 52802 12586
rect 53226 11810 53260 12586
rect 53356 11810 53390 12586
rect 53814 11810 53848 12586
rect 53944 11810 53978 12586
rect 54402 11810 54436 12586
rect 54532 11810 54566 12586
rect 54990 11810 55024 12586
rect 55120 11810 55154 12586
rect 55578 11810 55612 12586
rect 55708 11810 55742 12586
rect 56166 11810 56200 12586
rect 56296 11810 56330 12586
rect 56754 11810 56788 12586
rect 56884 11810 56918 12586
rect 57342 11810 57376 12586
rect 57472 11810 57506 12586
rect 57930 11810 57964 12586
rect 58060 11810 58094 12586
rect 58518 11810 58552 12586
rect 58648 11810 58682 12586
rect 59106 11810 59140 12586
rect 59236 11810 59270 12586
rect 59694 11810 59728 12586
rect 59824 11810 59858 12586
rect 60282 11810 60316 12586
rect 60412 11810 60446 12586
rect 60870 11810 60904 12586
rect 61000 11810 61034 12586
rect 61458 11810 61492 12586
rect 61588 11810 61622 12586
rect 62046 11810 62080 12586
rect 62176 11810 62210 12586
rect 62634 11810 62668 12586
rect 62764 11810 62798 12586
rect 63222 11810 63256 12586
rect 63352 11810 63386 12586
rect 63810 11810 63844 12586
rect 63940 11810 63974 12586
rect 64398 11810 64432 12586
rect 64528 11810 64562 12586
rect 64986 11810 65020 12586
rect 65116 11810 65150 12586
rect 65574 11810 65608 12586
rect 65704 11810 65738 12586
rect 66162 11810 66196 12586
rect 66292 11810 66326 12586
rect 66750 11810 66784 12586
rect 66880 11810 66914 12586
rect 67338 11810 67372 12586
rect 67468 11810 67502 12586
rect 67926 11810 67960 12586
rect 68056 11810 68090 12586
rect 68514 11810 68548 12586
rect 68644 11810 68678 12586
rect 69102 11810 69136 12586
rect 69232 11810 69266 12586
rect 69690 11810 69724 12586
rect 69820 11810 69854 12586
rect 70278 11810 70312 12586
rect 70408 11810 70442 12586
rect 70866 11810 70900 12586
rect 70996 11810 71030 12586
rect 71454 11810 71488 12586
rect 43360 10810 43394 11586
rect 43818 10810 43852 11586
rect 43948 10810 43982 11586
rect 44406 10810 44440 11586
rect 44536 10810 44570 11586
rect 44994 10810 45028 11586
rect 45124 10810 45158 11586
rect 45582 10810 45616 11586
rect 45712 10810 45746 11586
rect 46170 10810 46204 11586
rect 46300 10810 46334 11586
rect 46758 10810 46792 11586
rect 46888 10810 46922 11586
rect 47346 10810 47380 11586
rect 47476 10810 47510 11586
rect 47934 10810 47968 11586
rect 48064 10810 48098 11586
rect 48522 10810 48556 11586
rect 48652 10810 48686 11586
rect 49110 10810 49144 11586
rect 49240 10810 49274 11586
rect 49698 10810 49732 11586
rect 49828 10810 49862 11586
rect 50286 10810 50320 11586
rect 50416 10810 50450 11586
rect 50874 10810 50908 11586
rect 51004 10810 51038 11586
rect 51462 10810 51496 11586
rect 51592 10810 51626 11586
rect 52050 10810 52084 11586
rect 52180 10810 52214 11586
rect 52638 10810 52672 11586
rect 52768 10810 52802 11586
rect 53226 10810 53260 11586
rect 53356 10810 53390 11586
rect 53814 10810 53848 11586
rect 53944 10810 53978 11586
rect 54402 10810 54436 11586
rect 54532 10810 54566 11586
rect 54990 10810 55024 11586
rect 55120 10810 55154 11586
rect 55578 10810 55612 11586
rect 55708 10810 55742 11586
rect 56166 10810 56200 11586
rect 56296 10810 56330 11586
rect 56754 10810 56788 11586
rect 56884 10810 56918 11586
rect 57342 10810 57376 11586
rect 57472 10810 57506 11586
rect 57930 10810 57964 11586
rect 58060 10810 58094 11586
rect 58518 10810 58552 11586
rect 58648 10810 58682 11586
rect 59106 10810 59140 11586
rect 59236 10810 59270 11586
rect 59694 10810 59728 11586
rect 59824 10810 59858 11586
rect 60282 10810 60316 11586
rect 60412 10810 60446 11586
rect 60870 10810 60904 11586
rect 61000 10810 61034 11586
rect 61458 10810 61492 11586
rect 61588 10810 61622 11586
rect 62046 10810 62080 11586
rect 62176 10810 62210 11586
rect 62634 10810 62668 11586
rect 62764 10810 62798 11586
rect 63222 10810 63256 11586
rect 63352 10810 63386 11586
rect 63810 10810 63844 11586
rect 63940 10810 63974 11586
rect 64398 10810 64432 11586
rect 64528 10810 64562 11586
rect 64986 10810 65020 11586
rect 65116 10810 65150 11586
rect 65574 10810 65608 11586
rect 65704 10810 65738 11586
rect 66162 10810 66196 11586
rect 66292 10810 66326 11586
rect 66750 10810 66784 11586
rect 66880 10810 66914 11586
rect 67338 10810 67372 11586
rect 67468 10810 67502 11586
rect 67926 10810 67960 11586
rect 68056 10810 68090 11586
rect 68514 10810 68548 11586
rect 68644 10810 68678 11586
rect 69102 10810 69136 11586
rect 69232 10810 69266 11586
rect 69690 10810 69724 11586
rect 69820 10810 69854 11586
rect 70278 10810 70312 11586
rect 70408 10810 70442 11586
rect 70866 10810 70900 11586
rect 70996 10810 71030 11586
rect 71454 10810 71488 11586
rect 43360 9810 43394 10586
rect 43818 9810 43852 10586
rect 43948 9810 43982 10586
rect 44406 9810 44440 10586
rect 44536 9810 44570 10586
rect 44994 9810 45028 10586
rect 45124 9810 45158 10586
rect 45582 9810 45616 10586
rect 45712 9810 45746 10586
rect 46170 9810 46204 10586
rect 46300 9810 46334 10586
rect 46758 9810 46792 10586
rect 46888 9810 46922 10586
rect 47346 9810 47380 10586
rect 47476 9810 47510 10586
rect 47934 9810 47968 10586
rect 48064 9810 48098 10586
rect 48522 9810 48556 10586
rect 48652 9810 48686 10586
rect 49110 9810 49144 10586
rect 49240 9810 49274 10586
rect 49698 9810 49732 10586
rect 49828 9810 49862 10586
rect 50286 9810 50320 10586
rect 50416 9810 50450 10586
rect 50874 9810 50908 10586
rect 51004 9810 51038 10586
rect 51462 9810 51496 10586
rect 51592 9810 51626 10586
rect 52050 9810 52084 10586
rect 52180 9810 52214 10586
rect 52638 9810 52672 10586
rect 52768 9810 52802 10586
rect 53226 9810 53260 10586
rect 53356 9810 53390 10586
rect 53814 9810 53848 10586
rect 53944 9810 53978 10586
rect 54402 9810 54436 10586
rect 54532 9810 54566 10586
rect 54990 9810 55024 10586
rect 55120 9810 55154 10586
rect 55578 9810 55612 10586
rect 55708 9810 55742 10586
rect 56166 9810 56200 10586
rect 56296 9810 56330 10586
rect 56754 9810 56788 10586
rect 56884 9810 56918 10586
rect 57342 9810 57376 10586
rect 57472 9810 57506 10586
rect 57930 9810 57964 10586
rect 58060 9810 58094 10586
rect 58518 9810 58552 10586
rect 58648 9810 58682 10586
rect 59106 9810 59140 10586
rect 59236 9810 59270 10586
rect 59694 9810 59728 10586
rect 59824 9810 59858 10586
rect 60282 9810 60316 10586
rect 60412 9810 60446 10586
rect 60870 9810 60904 10586
rect 61000 9810 61034 10586
rect 61458 9810 61492 10586
rect 61588 9810 61622 10586
rect 62046 9810 62080 10586
rect 62176 9810 62210 10586
rect 62634 9810 62668 10586
rect 62764 9810 62798 10586
rect 63222 9810 63256 10586
rect 63352 9810 63386 10586
rect 63810 9810 63844 10586
rect 63940 9810 63974 10586
rect 64398 9810 64432 10586
rect 64528 9810 64562 10586
rect 64986 9810 65020 10586
rect 65116 9810 65150 10586
rect 65574 9810 65608 10586
rect 65704 9810 65738 10586
rect 66162 9810 66196 10586
rect 66292 9810 66326 10586
rect 66750 9810 66784 10586
rect 66880 9810 66914 10586
rect 67338 9810 67372 10586
rect 67468 9810 67502 10586
rect 67926 9810 67960 10586
rect 68056 9810 68090 10586
rect 68514 9810 68548 10586
rect 68644 9810 68678 10586
rect 69102 9810 69136 10586
rect 69232 9810 69266 10586
rect 69690 9810 69724 10586
rect 69820 9810 69854 10586
rect 70278 9810 70312 10586
rect 70408 9810 70442 10586
rect 70866 9810 70900 10586
rect 70996 9810 71030 10586
rect 71454 9810 71488 10586
rect 56412 7364 56446 8140
rect 56540 7364 56574 8140
rect 56678 7364 56712 8140
rect 56806 7364 56840 8140
rect 56944 7364 56978 8140
rect 57072 7364 57106 8140
rect 57210 7364 57244 8140
rect 57338 7364 57372 8140
rect 57476 7364 57510 8140
rect 57604 7364 57638 8140
rect 57742 7364 57776 8140
rect 57870 7364 57904 8140
rect 58008 7364 58042 8140
rect 58136 7364 58170 8140
rect 58274 7364 58308 8140
rect 58402 7364 58436 8140
rect 56412 6354 56446 7130
rect 56540 6354 56574 7130
rect 56678 6354 56712 7130
rect 56806 6354 56840 7130
rect 56944 6354 56978 7130
rect 57072 6354 57106 7130
rect 57210 6354 57244 7130
rect 57338 6354 57372 7130
rect 57476 6354 57510 7130
rect 57604 6354 57638 7130
rect 57742 6354 57776 7130
rect 57870 6354 57904 7130
rect 58008 6354 58042 7130
rect 58136 6354 58170 7130
rect 58274 6354 58308 7130
rect 58402 6354 58436 7130
rect 56412 5344 56446 6120
rect 56540 5344 56574 6120
rect 56678 5344 56712 6120
rect 56806 5344 56840 6120
rect 56944 5344 56978 6120
rect 57072 5344 57106 6120
rect 57210 5344 57244 6120
rect 57338 5344 57372 6120
rect 57476 5344 57510 6120
rect 57604 5344 57638 6120
rect 57742 5344 57776 6120
rect 57870 5344 57904 6120
rect 58008 5344 58042 6120
rect 58136 5344 58170 6120
rect 58274 5344 58308 6120
rect 58402 5344 58436 6120
<< nsubdiff >>
rect 56026 8622 56060 8656
rect 58788 8622 58822 8656
rect 56026 4826 56060 4860
rect 58788 4826 58822 4860
<< psubdiffcont >>
rect 52406 17152 62444 17186
rect 52318 14838 52352 17118
rect 62498 14838 62532 17120
rect 52352 14750 62498 14784
rect 56784 4430 57994 4464
rect 56638 2082 56672 4430
rect 58178 2082 58212 4430
rect 56796 2048 58006 2082
<< nsubdiffcont >>
rect 43174 12996 71696 13030
rect 43014 9420 43048 12968
rect 71800 9454 71834 13002
rect 43132 9366 71746 9400
rect 56060 8622 58788 8656
rect 56026 4860 56060 8622
rect 58788 4860 58822 8622
rect 56060 4826 58788 4860
<< poly >>
rect 52710 16842 52780 16852
rect 52710 16710 52726 16842
rect 52764 16710 52780 16842
rect 52710 16672 52780 16710
rect 52950 16842 53020 16852
rect 52950 16710 52966 16842
rect 53004 16710 53020 16842
rect 52950 16672 53020 16710
rect 53190 16842 53260 16852
rect 53190 16710 53206 16842
rect 53244 16710 53260 16842
rect 53190 16672 53260 16710
rect 53430 16842 53500 16852
rect 53430 16710 53446 16842
rect 53484 16710 53500 16842
rect 53430 16672 53500 16710
rect 53670 16842 53740 16852
rect 53670 16710 53686 16842
rect 53724 16710 53740 16842
rect 53670 16672 53740 16710
rect 53910 16842 53980 16852
rect 53910 16710 53926 16842
rect 53964 16710 53980 16842
rect 53910 16672 53980 16710
rect 54150 16842 54220 16852
rect 54150 16710 54166 16842
rect 54204 16710 54220 16842
rect 54150 16672 54220 16710
rect 54390 16842 54460 16852
rect 54390 16710 54406 16842
rect 54444 16710 54460 16842
rect 54390 16672 54460 16710
rect 54630 16842 54700 16852
rect 54630 16710 54646 16842
rect 54684 16710 54700 16842
rect 54630 16672 54700 16710
rect 54870 16842 54940 16852
rect 54870 16710 54886 16842
rect 54924 16710 54940 16842
rect 54870 16672 54940 16710
rect 55110 16842 55180 16852
rect 55110 16710 55126 16842
rect 55164 16710 55180 16842
rect 55110 16672 55180 16710
rect 55350 16842 55420 16852
rect 55350 16710 55366 16842
rect 55404 16710 55420 16842
rect 55350 16672 55420 16710
rect 55590 16842 55660 16852
rect 55590 16710 55606 16842
rect 55644 16710 55660 16842
rect 55590 16672 55660 16710
rect 55830 16842 55900 16852
rect 55830 16710 55846 16842
rect 55884 16710 55900 16842
rect 55830 16672 55900 16710
rect 56070 16842 56140 16852
rect 56070 16710 56086 16842
rect 56124 16710 56140 16842
rect 56070 16672 56140 16710
rect 56310 16842 56380 16852
rect 56310 16710 56326 16842
rect 56364 16710 56380 16842
rect 56310 16672 56380 16710
rect 56550 16842 56620 16852
rect 56550 16710 56566 16842
rect 56604 16710 56620 16842
rect 56550 16672 56620 16710
rect 56790 16842 56860 16852
rect 56790 16710 56806 16842
rect 56844 16710 56860 16842
rect 56790 16672 56860 16710
rect 57030 16842 57100 16852
rect 57030 16710 57046 16842
rect 57084 16710 57100 16842
rect 57030 16672 57100 16710
rect 57270 16842 57340 16852
rect 57270 16710 57286 16842
rect 57324 16710 57340 16842
rect 57270 16672 57340 16710
rect 57510 16842 57580 16852
rect 57510 16710 57526 16842
rect 57564 16710 57580 16842
rect 57510 16672 57580 16710
rect 57750 16842 57820 16852
rect 57750 16710 57766 16842
rect 57804 16710 57820 16842
rect 57750 16672 57820 16710
rect 57990 16842 58060 16852
rect 57990 16710 58006 16842
rect 58044 16710 58060 16842
rect 57990 16672 58060 16710
rect 58230 16842 58300 16852
rect 58230 16710 58246 16842
rect 58284 16710 58300 16842
rect 58230 16672 58300 16710
rect 58470 16842 58540 16852
rect 58470 16710 58486 16842
rect 58524 16710 58540 16842
rect 58470 16672 58540 16710
rect 58710 16842 58780 16852
rect 58710 16710 58726 16842
rect 58764 16710 58780 16842
rect 58710 16672 58780 16710
rect 58950 16842 59020 16852
rect 58950 16710 58966 16842
rect 59004 16710 59020 16842
rect 58950 16672 59020 16710
rect 59190 16842 59260 16852
rect 59190 16710 59206 16842
rect 59244 16710 59260 16842
rect 59190 16672 59260 16710
rect 59430 16842 59500 16852
rect 59430 16710 59446 16842
rect 59484 16710 59500 16842
rect 59430 16672 59500 16710
rect 59670 16842 59740 16852
rect 59670 16710 59686 16842
rect 59724 16710 59740 16842
rect 59670 16672 59740 16710
rect 59910 16842 59980 16852
rect 59910 16710 59926 16842
rect 59964 16710 59980 16842
rect 59910 16672 59980 16710
rect 60150 16842 60220 16852
rect 60150 16710 60166 16842
rect 60204 16710 60220 16842
rect 60150 16672 60220 16710
rect 60390 16842 60460 16852
rect 60390 16710 60406 16842
rect 60444 16710 60460 16842
rect 60390 16672 60460 16710
rect 60630 16842 60700 16852
rect 60630 16710 60646 16842
rect 60684 16710 60700 16842
rect 60630 16672 60700 16710
rect 60870 16842 60940 16852
rect 60870 16710 60886 16842
rect 60924 16710 60940 16842
rect 60870 16672 60940 16710
rect 61110 16842 61180 16852
rect 61110 16710 61126 16842
rect 61164 16710 61180 16842
rect 61110 16672 61180 16710
rect 61350 16842 61420 16852
rect 61350 16710 61366 16842
rect 61404 16710 61420 16842
rect 61350 16672 61420 16710
rect 61590 16842 61660 16852
rect 61590 16710 61606 16842
rect 61644 16710 61660 16842
rect 61590 16672 61660 16710
rect 61830 16842 61900 16852
rect 61830 16710 61846 16842
rect 61884 16710 61900 16842
rect 61830 16672 61900 16710
rect 62070 16842 62140 16852
rect 62070 16710 62086 16842
rect 62124 16710 62140 16842
rect 62070 16672 62140 16710
rect 52710 16034 52780 16072
rect 52710 15902 52726 16034
rect 52764 15902 52780 16034
rect 52710 15864 52780 15902
rect 52950 16034 53020 16072
rect 52950 15902 52966 16034
rect 53004 15902 53020 16034
rect 52950 15864 53020 15902
rect 53190 16034 53260 16072
rect 53190 15902 53206 16034
rect 53244 15902 53260 16034
rect 53190 15864 53260 15902
rect 53430 16034 53500 16072
rect 53430 15902 53446 16034
rect 53484 15902 53500 16034
rect 53430 15864 53500 15902
rect 53670 16034 53740 16072
rect 53670 15902 53686 16034
rect 53724 15902 53740 16034
rect 53670 15864 53740 15902
rect 53910 16034 53980 16072
rect 53910 15902 53926 16034
rect 53964 15902 53980 16034
rect 53910 15864 53980 15902
rect 54150 16034 54220 16072
rect 54150 15902 54166 16034
rect 54204 15902 54220 16034
rect 54150 15864 54220 15902
rect 54390 16034 54460 16072
rect 54390 15902 54406 16034
rect 54444 15902 54460 16034
rect 54390 15864 54460 15902
rect 54630 16034 54700 16072
rect 54630 15902 54646 16034
rect 54684 15902 54700 16034
rect 54630 15864 54700 15902
rect 54870 16034 54940 16072
rect 54870 15902 54886 16034
rect 54924 15902 54940 16034
rect 54870 15864 54940 15902
rect 55110 16034 55180 16072
rect 55110 15902 55126 16034
rect 55164 15902 55180 16034
rect 55110 15864 55180 15902
rect 55350 16034 55420 16072
rect 55350 15902 55366 16034
rect 55404 15902 55420 16034
rect 55350 15864 55420 15902
rect 55590 16034 55660 16072
rect 55590 15902 55606 16034
rect 55644 15902 55660 16034
rect 55590 15864 55660 15902
rect 55830 16034 55900 16072
rect 55830 15902 55846 16034
rect 55884 15902 55900 16034
rect 55830 15864 55900 15902
rect 56070 16034 56140 16072
rect 56070 15902 56086 16034
rect 56124 15902 56140 16034
rect 56070 15864 56140 15902
rect 56310 16034 56380 16072
rect 56310 15902 56326 16034
rect 56364 15902 56380 16034
rect 56310 15864 56380 15902
rect 56550 16034 56620 16072
rect 56550 15902 56566 16034
rect 56604 15902 56620 16034
rect 56550 15864 56620 15902
rect 56790 16034 56860 16072
rect 56790 15902 56806 16034
rect 56844 15902 56860 16034
rect 56790 15864 56860 15902
rect 57030 16034 57100 16072
rect 57030 15902 57046 16034
rect 57084 15902 57100 16034
rect 57030 15864 57100 15902
rect 57270 16034 57340 16072
rect 57270 15902 57286 16034
rect 57324 15902 57340 16034
rect 57270 15864 57340 15902
rect 57510 16034 57580 16072
rect 57510 15902 57526 16034
rect 57564 15902 57580 16034
rect 57510 15864 57580 15902
rect 57750 16034 57820 16072
rect 57750 15902 57766 16034
rect 57804 15902 57820 16034
rect 57750 15864 57820 15902
rect 57990 16034 58060 16072
rect 57990 15902 58006 16034
rect 58044 15902 58060 16034
rect 57990 15864 58060 15902
rect 58230 16034 58300 16072
rect 58230 15902 58246 16034
rect 58284 15902 58300 16034
rect 58230 15864 58300 15902
rect 58470 16034 58540 16072
rect 58470 15902 58486 16034
rect 58524 15902 58540 16034
rect 58470 15864 58540 15902
rect 58710 16034 58780 16072
rect 58710 15902 58726 16034
rect 58764 15902 58780 16034
rect 58710 15864 58780 15902
rect 58950 16034 59020 16072
rect 58950 15902 58966 16034
rect 59004 15902 59020 16034
rect 58950 15864 59020 15902
rect 59190 16034 59260 16072
rect 59190 15902 59206 16034
rect 59244 15902 59260 16034
rect 59190 15864 59260 15902
rect 59430 16034 59500 16072
rect 59430 15902 59446 16034
rect 59484 15902 59500 16034
rect 59430 15864 59500 15902
rect 59670 16034 59740 16072
rect 59670 15902 59686 16034
rect 59724 15902 59740 16034
rect 59670 15864 59740 15902
rect 59910 16034 59980 16072
rect 59910 15902 59926 16034
rect 59964 15902 59980 16034
rect 59910 15864 59980 15902
rect 60150 16034 60220 16072
rect 60150 15902 60166 16034
rect 60204 15902 60220 16034
rect 60150 15864 60220 15902
rect 60390 16034 60460 16072
rect 60390 15902 60406 16034
rect 60444 15902 60460 16034
rect 60390 15864 60460 15902
rect 60630 16034 60700 16072
rect 60630 15902 60646 16034
rect 60684 15902 60700 16034
rect 60630 15864 60700 15902
rect 60870 16034 60940 16072
rect 60870 15902 60886 16034
rect 60924 15902 60940 16034
rect 60870 15864 60940 15902
rect 61110 16034 61180 16072
rect 61110 15902 61126 16034
rect 61164 15902 61180 16034
rect 61110 15864 61180 15902
rect 61350 16034 61420 16072
rect 61350 15902 61366 16034
rect 61404 15902 61420 16034
rect 61350 15864 61420 15902
rect 61590 16034 61660 16072
rect 61590 15902 61606 16034
rect 61644 15902 61660 16034
rect 61590 15864 61660 15902
rect 61830 16034 61900 16072
rect 61830 15902 61846 16034
rect 61884 15902 61900 16034
rect 61830 15864 61900 15902
rect 62070 16034 62140 16072
rect 62070 15902 62086 16034
rect 62124 15902 62140 16034
rect 62070 15864 62140 15902
rect 52710 15226 52780 15264
rect 52710 15094 52726 15226
rect 52764 15094 52780 15226
rect 52710 15084 52780 15094
rect 52950 15226 53020 15264
rect 52950 15094 52966 15226
rect 53004 15094 53020 15226
rect 52950 15084 53020 15094
rect 53190 15226 53260 15264
rect 53190 15094 53206 15226
rect 53244 15094 53260 15226
rect 53190 15084 53260 15094
rect 53430 15226 53500 15264
rect 53430 15094 53446 15226
rect 53484 15094 53500 15226
rect 53430 15084 53500 15094
rect 53670 15226 53740 15264
rect 53670 15094 53686 15226
rect 53724 15094 53740 15226
rect 53670 15084 53740 15094
rect 53910 15226 53980 15264
rect 53910 15094 53926 15226
rect 53964 15094 53980 15226
rect 53910 15084 53980 15094
rect 54150 15226 54220 15264
rect 54150 15094 54166 15226
rect 54204 15094 54220 15226
rect 54150 15084 54220 15094
rect 54390 15226 54460 15264
rect 54390 15094 54406 15226
rect 54444 15094 54460 15226
rect 54390 15084 54460 15094
rect 54630 15226 54700 15264
rect 54630 15094 54646 15226
rect 54684 15094 54700 15226
rect 54630 15084 54700 15094
rect 54870 15226 54940 15264
rect 54870 15094 54886 15226
rect 54924 15094 54940 15226
rect 54870 15084 54940 15094
rect 55110 15226 55180 15264
rect 55110 15094 55126 15226
rect 55164 15094 55180 15226
rect 55110 15084 55180 15094
rect 55350 15226 55420 15264
rect 55350 15094 55366 15226
rect 55404 15094 55420 15226
rect 55350 15084 55420 15094
rect 55590 15226 55660 15264
rect 55590 15094 55606 15226
rect 55644 15094 55660 15226
rect 55590 15084 55660 15094
rect 55830 15226 55900 15264
rect 55830 15094 55846 15226
rect 55884 15094 55900 15226
rect 55830 15084 55900 15094
rect 56070 15226 56140 15264
rect 56070 15094 56086 15226
rect 56124 15094 56140 15226
rect 56070 15084 56140 15094
rect 56310 15226 56380 15264
rect 56310 15094 56326 15226
rect 56364 15094 56380 15226
rect 56310 15084 56380 15094
rect 56550 15226 56620 15264
rect 56550 15094 56566 15226
rect 56604 15094 56620 15226
rect 56550 15084 56620 15094
rect 56790 15226 56860 15264
rect 56790 15094 56806 15226
rect 56844 15094 56860 15226
rect 56790 15084 56860 15094
rect 57030 15226 57100 15264
rect 57030 15094 57046 15226
rect 57084 15094 57100 15226
rect 57030 15084 57100 15094
rect 57270 15226 57340 15264
rect 57270 15094 57286 15226
rect 57324 15094 57340 15226
rect 57270 15084 57340 15094
rect 57510 15226 57580 15264
rect 57510 15094 57526 15226
rect 57564 15094 57580 15226
rect 57510 15084 57580 15094
rect 57750 15226 57820 15264
rect 57750 15094 57766 15226
rect 57804 15094 57820 15226
rect 57750 15084 57820 15094
rect 57990 15226 58060 15264
rect 57990 15094 58006 15226
rect 58044 15094 58060 15226
rect 57990 15084 58060 15094
rect 58230 15226 58300 15264
rect 58230 15094 58246 15226
rect 58284 15094 58300 15226
rect 58230 15084 58300 15094
rect 58470 15226 58540 15264
rect 58470 15094 58486 15226
rect 58524 15094 58540 15226
rect 58470 15084 58540 15094
rect 58710 15226 58780 15264
rect 58710 15094 58726 15226
rect 58764 15094 58780 15226
rect 58710 15084 58780 15094
rect 58950 15226 59020 15264
rect 58950 15094 58966 15226
rect 59004 15094 59020 15226
rect 58950 15084 59020 15094
rect 59190 15226 59260 15264
rect 59190 15094 59206 15226
rect 59244 15094 59260 15226
rect 59190 15084 59260 15094
rect 59430 15226 59500 15264
rect 59430 15094 59446 15226
rect 59484 15094 59500 15226
rect 59430 15084 59500 15094
rect 59670 15226 59740 15264
rect 59670 15094 59686 15226
rect 59724 15094 59740 15226
rect 59670 15084 59740 15094
rect 59910 15226 59980 15264
rect 59910 15094 59926 15226
rect 59964 15094 59980 15226
rect 59910 15084 59980 15094
rect 60150 15226 60220 15264
rect 60150 15094 60166 15226
rect 60204 15094 60220 15226
rect 60150 15084 60220 15094
rect 60390 15226 60460 15264
rect 60390 15094 60406 15226
rect 60444 15094 60460 15226
rect 60390 15084 60460 15094
rect 60630 15226 60700 15264
rect 60630 15094 60646 15226
rect 60684 15094 60700 15226
rect 60630 15084 60700 15094
rect 60870 15226 60940 15264
rect 60870 15094 60886 15226
rect 60924 15094 60940 15226
rect 60870 15084 60940 15094
rect 61110 15226 61180 15264
rect 61110 15094 61126 15226
rect 61164 15094 61180 15226
rect 61110 15084 61180 15094
rect 61350 15226 61420 15264
rect 61350 15094 61366 15226
rect 61404 15094 61420 15226
rect 61350 15084 61420 15094
rect 61590 15226 61660 15264
rect 61590 15094 61606 15226
rect 61644 15094 61660 15226
rect 61590 15084 61660 15094
rect 61830 15226 61900 15264
rect 61830 15094 61846 15226
rect 61884 15094 61900 15226
rect 61830 15084 61900 15094
rect 62070 15226 62140 15264
rect 62070 15094 62086 15226
rect 62124 15094 62140 15226
rect 62070 15084 62140 15094
rect 43406 12679 43806 12695
rect 43406 12645 43422 12679
rect 43790 12645 43806 12679
rect 43406 12598 43806 12645
rect 43994 12679 44394 12695
rect 43994 12645 44010 12679
rect 44378 12645 44394 12679
rect 43994 12598 44394 12645
rect 44582 12679 44982 12695
rect 44582 12645 44598 12679
rect 44966 12645 44982 12679
rect 44582 12598 44982 12645
rect 45170 12679 45570 12695
rect 45170 12645 45186 12679
rect 45554 12645 45570 12679
rect 45170 12598 45570 12645
rect 45758 12679 46158 12695
rect 45758 12645 45774 12679
rect 46142 12645 46158 12679
rect 45758 12598 46158 12645
rect 46346 12679 46746 12695
rect 46346 12645 46362 12679
rect 46730 12645 46746 12679
rect 46346 12598 46746 12645
rect 46934 12679 47334 12695
rect 46934 12645 46950 12679
rect 47318 12645 47334 12679
rect 46934 12598 47334 12645
rect 47522 12679 47922 12695
rect 47522 12645 47538 12679
rect 47906 12645 47922 12679
rect 47522 12598 47922 12645
rect 48110 12679 48510 12695
rect 48110 12645 48126 12679
rect 48494 12645 48510 12679
rect 48110 12598 48510 12645
rect 48698 12679 49098 12695
rect 48698 12645 48714 12679
rect 49082 12645 49098 12679
rect 48698 12598 49098 12645
rect 49286 12679 49686 12695
rect 49286 12645 49302 12679
rect 49670 12645 49686 12679
rect 49286 12598 49686 12645
rect 49874 12679 50274 12695
rect 49874 12645 49890 12679
rect 50258 12645 50274 12679
rect 49874 12598 50274 12645
rect 50462 12679 50862 12695
rect 50462 12645 50478 12679
rect 50846 12645 50862 12679
rect 50462 12598 50862 12645
rect 51050 12679 51450 12695
rect 51050 12645 51066 12679
rect 51434 12645 51450 12679
rect 51050 12598 51450 12645
rect 51638 12679 52038 12695
rect 51638 12645 51654 12679
rect 52022 12645 52038 12679
rect 51638 12598 52038 12645
rect 52226 12679 52626 12695
rect 52226 12645 52242 12679
rect 52610 12645 52626 12679
rect 52226 12598 52626 12645
rect 52814 12679 53214 12695
rect 52814 12645 52830 12679
rect 53198 12645 53214 12679
rect 52814 12598 53214 12645
rect 53402 12679 53802 12695
rect 53402 12645 53418 12679
rect 53786 12645 53802 12679
rect 53402 12598 53802 12645
rect 53990 12679 54390 12695
rect 53990 12645 54006 12679
rect 54374 12645 54390 12679
rect 53990 12598 54390 12645
rect 54578 12679 54978 12695
rect 54578 12645 54594 12679
rect 54962 12645 54978 12679
rect 54578 12598 54978 12645
rect 55166 12679 55566 12695
rect 55166 12645 55182 12679
rect 55550 12645 55566 12679
rect 55166 12598 55566 12645
rect 55754 12679 56154 12695
rect 55754 12645 55770 12679
rect 56138 12645 56154 12679
rect 55754 12598 56154 12645
rect 56342 12679 56742 12695
rect 56342 12645 56358 12679
rect 56726 12645 56742 12679
rect 56342 12598 56742 12645
rect 56930 12679 57330 12695
rect 56930 12645 56946 12679
rect 57314 12645 57330 12679
rect 56930 12598 57330 12645
rect 57518 12679 57918 12695
rect 57518 12645 57534 12679
rect 57902 12645 57918 12679
rect 57518 12598 57918 12645
rect 58106 12679 58506 12695
rect 58106 12645 58122 12679
rect 58490 12645 58506 12679
rect 58106 12598 58506 12645
rect 58694 12679 59094 12695
rect 58694 12645 58710 12679
rect 59078 12645 59094 12679
rect 58694 12598 59094 12645
rect 59282 12679 59682 12695
rect 59282 12645 59298 12679
rect 59666 12645 59682 12679
rect 59282 12598 59682 12645
rect 59870 12679 60270 12695
rect 59870 12645 59886 12679
rect 60254 12645 60270 12679
rect 59870 12598 60270 12645
rect 60458 12679 60858 12695
rect 60458 12645 60474 12679
rect 60842 12645 60858 12679
rect 60458 12598 60858 12645
rect 61046 12679 61446 12695
rect 61046 12645 61062 12679
rect 61430 12645 61446 12679
rect 61046 12598 61446 12645
rect 61634 12679 62034 12695
rect 61634 12645 61650 12679
rect 62018 12645 62034 12679
rect 61634 12598 62034 12645
rect 62222 12679 62622 12695
rect 62222 12645 62238 12679
rect 62606 12645 62622 12679
rect 62222 12598 62622 12645
rect 62810 12679 63210 12695
rect 62810 12645 62826 12679
rect 63194 12645 63210 12679
rect 62810 12598 63210 12645
rect 63398 12679 63798 12695
rect 63398 12645 63414 12679
rect 63782 12645 63798 12679
rect 63398 12598 63798 12645
rect 63986 12679 64386 12695
rect 63986 12645 64002 12679
rect 64370 12645 64386 12679
rect 63986 12598 64386 12645
rect 64574 12679 64974 12695
rect 64574 12645 64590 12679
rect 64958 12645 64974 12679
rect 64574 12598 64974 12645
rect 65162 12679 65562 12695
rect 65162 12645 65178 12679
rect 65546 12645 65562 12679
rect 65162 12598 65562 12645
rect 65750 12679 66150 12695
rect 65750 12645 65766 12679
rect 66134 12645 66150 12679
rect 65750 12598 66150 12645
rect 66338 12679 66738 12695
rect 66338 12645 66354 12679
rect 66722 12645 66738 12679
rect 66338 12598 66738 12645
rect 66926 12679 67326 12695
rect 66926 12645 66942 12679
rect 67310 12645 67326 12679
rect 66926 12598 67326 12645
rect 67514 12679 67914 12695
rect 67514 12645 67530 12679
rect 67898 12645 67914 12679
rect 67514 12598 67914 12645
rect 68102 12679 68502 12695
rect 68102 12645 68118 12679
rect 68486 12645 68502 12679
rect 68102 12598 68502 12645
rect 68690 12679 69090 12695
rect 68690 12645 68706 12679
rect 69074 12645 69090 12679
rect 68690 12598 69090 12645
rect 69278 12679 69678 12695
rect 69278 12645 69294 12679
rect 69662 12645 69678 12679
rect 69278 12598 69678 12645
rect 69866 12679 70266 12695
rect 69866 12645 69882 12679
rect 70250 12645 70266 12679
rect 69866 12598 70266 12645
rect 70454 12679 70854 12695
rect 70454 12645 70470 12679
rect 70838 12645 70854 12679
rect 70454 12598 70854 12645
rect 71042 12679 71442 12695
rect 71042 12645 71058 12679
rect 71426 12645 71442 12679
rect 71042 12598 71442 12645
rect 43406 11751 43806 11798
rect 43406 11717 43422 11751
rect 43790 11717 43806 11751
rect 43406 11679 43806 11717
rect 43406 11645 43422 11679
rect 43790 11645 43806 11679
rect 43406 11598 43806 11645
rect 43994 11751 44394 11798
rect 43994 11717 44010 11751
rect 44378 11717 44394 11751
rect 43994 11679 44394 11717
rect 43994 11645 44010 11679
rect 44378 11645 44394 11679
rect 43994 11598 44394 11645
rect 44582 11751 44982 11798
rect 44582 11717 44598 11751
rect 44966 11717 44982 11751
rect 44582 11679 44982 11717
rect 44582 11645 44598 11679
rect 44966 11645 44982 11679
rect 44582 11598 44982 11645
rect 45170 11751 45570 11798
rect 45170 11717 45186 11751
rect 45554 11717 45570 11751
rect 45170 11679 45570 11717
rect 45170 11645 45186 11679
rect 45554 11645 45570 11679
rect 45170 11598 45570 11645
rect 45758 11751 46158 11798
rect 45758 11717 45774 11751
rect 46142 11717 46158 11751
rect 45758 11679 46158 11717
rect 45758 11645 45774 11679
rect 46142 11645 46158 11679
rect 45758 11598 46158 11645
rect 46346 11751 46746 11798
rect 46346 11717 46362 11751
rect 46730 11717 46746 11751
rect 46346 11679 46746 11717
rect 46346 11645 46362 11679
rect 46730 11645 46746 11679
rect 46346 11598 46746 11645
rect 46934 11751 47334 11798
rect 46934 11717 46950 11751
rect 47318 11717 47334 11751
rect 46934 11679 47334 11717
rect 46934 11645 46950 11679
rect 47318 11645 47334 11679
rect 46934 11598 47334 11645
rect 47522 11751 47922 11798
rect 47522 11717 47538 11751
rect 47906 11717 47922 11751
rect 47522 11679 47922 11717
rect 47522 11645 47538 11679
rect 47906 11645 47922 11679
rect 47522 11598 47922 11645
rect 48110 11751 48510 11798
rect 48110 11717 48126 11751
rect 48494 11717 48510 11751
rect 48110 11679 48510 11717
rect 48110 11645 48126 11679
rect 48494 11645 48510 11679
rect 48110 11598 48510 11645
rect 48698 11751 49098 11798
rect 48698 11717 48714 11751
rect 49082 11717 49098 11751
rect 48698 11679 49098 11717
rect 48698 11645 48714 11679
rect 49082 11645 49098 11679
rect 48698 11598 49098 11645
rect 49286 11751 49686 11798
rect 49286 11717 49302 11751
rect 49670 11717 49686 11751
rect 49286 11679 49686 11717
rect 49286 11645 49302 11679
rect 49670 11645 49686 11679
rect 49286 11598 49686 11645
rect 49874 11751 50274 11798
rect 49874 11717 49890 11751
rect 50258 11717 50274 11751
rect 49874 11679 50274 11717
rect 49874 11645 49890 11679
rect 50258 11645 50274 11679
rect 49874 11598 50274 11645
rect 50462 11751 50862 11798
rect 50462 11717 50478 11751
rect 50846 11717 50862 11751
rect 50462 11679 50862 11717
rect 50462 11645 50478 11679
rect 50846 11645 50862 11679
rect 50462 11598 50862 11645
rect 51050 11751 51450 11798
rect 51050 11717 51066 11751
rect 51434 11717 51450 11751
rect 51050 11679 51450 11717
rect 51050 11645 51066 11679
rect 51434 11645 51450 11679
rect 51050 11598 51450 11645
rect 51638 11751 52038 11798
rect 51638 11717 51654 11751
rect 52022 11717 52038 11751
rect 51638 11679 52038 11717
rect 51638 11645 51654 11679
rect 52022 11645 52038 11679
rect 51638 11598 52038 11645
rect 52226 11751 52626 11798
rect 52226 11717 52242 11751
rect 52610 11717 52626 11751
rect 52226 11679 52626 11717
rect 52226 11645 52242 11679
rect 52610 11645 52626 11679
rect 52226 11598 52626 11645
rect 52814 11751 53214 11798
rect 52814 11717 52830 11751
rect 53198 11717 53214 11751
rect 52814 11679 53214 11717
rect 52814 11645 52830 11679
rect 53198 11645 53214 11679
rect 52814 11598 53214 11645
rect 53402 11751 53802 11798
rect 53402 11717 53418 11751
rect 53786 11717 53802 11751
rect 53402 11679 53802 11717
rect 53402 11645 53418 11679
rect 53786 11645 53802 11679
rect 53402 11598 53802 11645
rect 53990 11751 54390 11798
rect 53990 11717 54006 11751
rect 54374 11717 54390 11751
rect 53990 11679 54390 11717
rect 53990 11645 54006 11679
rect 54374 11645 54390 11679
rect 53990 11598 54390 11645
rect 54578 11751 54978 11798
rect 54578 11717 54594 11751
rect 54962 11717 54978 11751
rect 54578 11679 54978 11717
rect 54578 11645 54594 11679
rect 54962 11645 54978 11679
rect 54578 11598 54978 11645
rect 55166 11751 55566 11798
rect 55166 11717 55182 11751
rect 55550 11717 55566 11751
rect 55166 11679 55566 11717
rect 55166 11645 55182 11679
rect 55550 11645 55566 11679
rect 55166 11598 55566 11645
rect 55754 11751 56154 11798
rect 55754 11717 55770 11751
rect 56138 11717 56154 11751
rect 55754 11679 56154 11717
rect 55754 11645 55770 11679
rect 56138 11645 56154 11679
rect 55754 11598 56154 11645
rect 56342 11751 56742 11798
rect 56342 11717 56358 11751
rect 56726 11717 56742 11751
rect 56342 11679 56742 11717
rect 56342 11645 56358 11679
rect 56726 11645 56742 11679
rect 56342 11598 56742 11645
rect 56930 11751 57330 11798
rect 56930 11717 56946 11751
rect 57314 11717 57330 11751
rect 56930 11679 57330 11717
rect 56930 11645 56946 11679
rect 57314 11645 57330 11679
rect 56930 11598 57330 11645
rect 57518 11751 57918 11798
rect 57518 11717 57534 11751
rect 57902 11717 57918 11751
rect 57518 11679 57918 11717
rect 57518 11645 57534 11679
rect 57902 11645 57918 11679
rect 57518 11598 57918 11645
rect 58106 11751 58506 11798
rect 58106 11717 58122 11751
rect 58490 11717 58506 11751
rect 58106 11679 58506 11717
rect 58106 11645 58122 11679
rect 58490 11645 58506 11679
rect 58106 11598 58506 11645
rect 58694 11751 59094 11798
rect 58694 11717 58710 11751
rect 59078 11717 59094 11751
rect 58694 11679 59094 11717
rect 58694 11645 58710 11679
rect 59078 11645 59094 11679
rect 58694 11598 59094 11645
rect 59282 11751 59682 11798
rect 59282 11717 59298 11751
rect 59666 11717 59682 11751
rect 59282 11679 59682 11717
rect 59282 11645 59298 11679
rect 59666 11645 59682 11679
rect 59282 11598 59682 11645
rect 59870 11751 60270 11798
rect 59870 11717 59886 11751
rect 60254 11717 60270 11751
rect 59870 11679 60270 11717
rect 59870 11645 59886 11679
rect 60254 11645 60270 11679
rect 59870 11598 60270 11645
rect 60458 11751 60858 11798
rect 60458 11717 60474 11751
rect 60842 11717 60858 11751
rect 60458 11679 60858 11717
rect 60458 11645 60474 11679
rect 60842 11645 60858 11679
rect 60458 11598 60858 11645
rect 61046 11751 61446 11798
rect 61046 11717 61062 11751
rect 61430 11717 61446 11751
rect 61046 11679 61446 11717
rect 61046 11645 61062 11679
rect 61430 11645 61446 11679
rect 61046 11598 61446 11645
rect 61634 11751 62034 11798
rect 61634 11717 61650 11751
rect 62018 11717 62034 11751
rect 61634 11679 62034 11717
rect 61634 11645 61650 11679
rect 62018 11645 62034 11679
rect 61634 11598 62034 11645
rect 62222 11751 62622 11798
rect 62222 11717 62238 11751
rect 62606 11717 62622 11751
rect 62222 11679 62622 11717
rect 62222 11645 62238 11679
rect 62606 11645 62622 11679
rect 62222 11598 62622 11645
rect 62810 11751 63210 11798
rect 62810 11717 62826 11751
rect 63194 11717 63210 11751
rect 62810 11679 63210 11717
rect 62810 11645 62826 11679
rect 63194 11645 63210 11679
rect 62810 11598 63210 11645
rect 63398 11751 63798 11798
rect 63398 11717 63414 11751
rect 63782 11717 63798 11751
rect 63398 11679 63798 11717
rect 63398 11645 63414 11679
rect 63782 11645 63798 11679
rect 63398 11598 63798 11645
rect 63986 11751 64386 11798
rect 63986 11717 64002 11751
rect 64370 11717 64386 11751
rect 63986 11679 64386 11717
rect 63986 11645 64002 11679
rect 64370 11645 64386 11679
rect 63986 11598 64386 11645
rect 64574 11751 64974 11798
rect 64574 11717 64590 11751
rect 64958 11717 64974 11751
rect 64574 11679 64974 11717
rect 64574 11645 64590 11679
rect 64958 11645 64974 11679
rect 64574 11598 64974 11645
rect 65162 11751 65562 11798
rect 65162 11717 65178 11751
rect 65546 11717 65562 11751
rect 65162 11679 65562 11717
rect 65162 11645 65178 11679
rect 65546 11645 65562 11679
rect 65162 11598 65562 11645
rect 65750 11751 66150 11798
rect 65750 11717 65766 11751
rect 66134 11717 66150 11751
rect 65750 11679 66150 11717
rect 65750 11645 65766 11679
rect 66134 11645 66150 11679
rect 65750 11598 66150 11645
rect 66338 11751 66738 11798
rect 66338 11717 66354 11751
rect 66722 11717 66738 11751
rect 66338 11679 66738 11717
rect 66338 11645 66354 11679
rect 66722 11645 66738 11679
rect 66338 11598 66738 11645
rect 66926 11751 67326 11798
rect 66926 11717 66942 11751
rect 67310 11717 67326 11751
rect 66926 11679 67326 11717
rect 66926 11645 66942 11679
rect 67310 11645 67326 11679
rect 66926 11598 67326 11645
rect 67514 11751 67914 11798
rect 67514 11717 67530 11751
rect 67898 11717 67914 11751
rect 67514 11679 67914 11717
rect 67514 11645 67530 11679
rect 67898 11645 67914 11679
rect 67514 11598 67914 11645
rect 68102 11751 68502 11798
rect 68102 11717 68118 11751
rect 68486 11717 68502 11751
rect 68102 11679 68502 11717
rect 68102 11645 68118 11679
rect 68486 11645 68502 11679
rect 68102 11598 68502 11645
rect 68690 11751 69090 11798
rect 68690 11717 68706 11751
rect 69074 11717 69090 11751
rect 68690 11679 69090 11717
rect 68690 11645 68706 11679
rect 69074 11645 69090 11679
rect 68690 11598 69090 11645
rect 69278 11751 69678 11798
rect 69278 11717 69294 11751
rect 69662 11717 69678 11751
rect 69278 11679 69678 11717
rect 69278 11645 69294 11679
rect 69662 11645 69678 11679
rect 69278 11598 69678 11645
rect 69866 11751 70266 11798
rect 69866 11717 69882 11751
rect 70250 11717 70266 11751
rect 69866 11679 70266 11717
rect 69866 11645 69882 11679
rect 70250 11645 70266 11679
rect 69866 11598 70266 11645
rect 70454 11751 70854 11798
rect 70454 11717 70470 11751
rect 70838 11717 70854 11751
rect 70454 11679 70854 11717
rect 70454 11645 70470 11679
rect 70838 11645 70854 11679
rect 70454 11598 70854 11645
rect 71042 11751 71442 11798
rect 71042 11717 71058 11751
rect 71426 11717 71442 11751
rect 71042 11679 71442 11717
rect 71042 11645 71058 11679
rect 71426 11645 71442 11679
rect 71042 11598 71442 11645
rect 43406 10751 43806 10798
rect 43406 10717 43422 10751
rect 43790 10717 43806 10751
rect 43406 10679 43806 10717
rect 43406 10645 43422 10679
rect 43790 10645 43806 10679
rect 43406 10598 43806 10645
rect 43994 10751 44394 10798
rect 43994 10717 44010 10751
rect 44378 10717 44394 10751
rect 43994 10679 44394 10717
rect 43994 10645 44010 10679
rect 44378 10645 44394 10679
rect 43994 10598 44394 10645
rect 44582 10751 44982 10798
rect 44582 10717 44598 10751
rect 44966 10717 44982 10751
rect 44582 10679 44982 10717
rect 44582 10645 44598 10679
rect 44966 10645 44982 10679
rect 44582 10598 44982 10645
rect 45170 10751 45570 10798
rect 45170 10717 45186 10751
rect 45554 10717 45570 10751
rect 45170 10679 45570 10717
rect 45170 10645 45186 10679
rect 45554 10645 45570 10679
rect 45170 10598 45570 10645
rect 45758 10751 46158 10798
rect 45758 10717 45774 10751
rect 46142 10717 46158 10751
rect 45758 10679 46158 10717
rect 45758 10645 45774 10679
rect 46142 10645 46158 10679
rect 45758 10598 46158 10645
rect 46346 10751 46746 10798
rect 46346 10717 46362 10751
rect 46730 10717 46746 10751
rect 46346 10679 46746 10717
rect 46346 10645 46362 10679
rect 46730 10645 46746 10679
rect 46346 10598 46746 10645
rect 46934 10751 47334 10798
rect 46934 10717 46950 10751
rect 47318 10717 47334 10751
rect 46934 10679 47334 10717
rect 46934 10645 46950 10679
rect 47318 10645 47334 10679
rect 46934 10598 47334 10645
rect 47522 10751 47922 10798
rect 47522 10717 47538 10751
rect 47906 10717 47922 10751
rect 47522 10679 47922 10717
rect 47522 10645 47538 10679
rect 47906 10645 47922 10679
rect 47522 10598 47922 10645
rect 48110 10751 48510 10798
rect 48110 10717 48126 10751
rect 48494 10717 48510 10751
rect 48110 10679 48510 10717
rect 48110 10645 48126 10679
rect 48494 10645 48510 10679
rect 48110 10598 48510 10645
rect 48698 10751 49098 10798
rect 48698 10717 48714 10751
rect 49082 10717 49098 10751
rect 48698 10679 49098 10717
rect 48698 10645 48714 10679
rect 49082 10645 49098 10679
rect 48698 10598 49098 10645
rect 49286 10751 49686 10798
rect 49286 10717 49302 10751
rect 49670 10717 49686 10751
rect 49286 10679 49686 10717
rect 49286 10645 49302 10679
rect 49670 10645 49686 10679
rect 49286 10598 49686 10645
rect 49874 10751 50274 10798
rect 49874 10717 49890 10751
rect 50258 10717 50274 10751
rect 49874 10679 50274 10717
rect 49874 10645 49890 10679
rect 50258 10645 50274 10679
rect 49874 10598 50274 10645
rect 50462 10751 50862 10798
rect 50462 10717 50478 10751
rect 50846 10717 50862 10751
rect 50462 10679 50862 10717
rect 50462 10645 50478 10679
rect 50846 10645 50862 10679
rect 50462 10598 50862 10645
rect 51050 10751 51450 10798
rect 51050 10717 51066 10751
rect 51434 10717 51450 10751
rect 51050 10679 51450 10717
rect 51050 10645 51066 10679
rect 51434 10645 51450 10679
rect 51050 10598 51450 10645
rect 51638 10751 52038 10798
rect 51638 10717 51654 10751
rect 52022 10717 52038 10751
rect 51638 10679 52038 10717
rect 51638 10645 51654 10679
rect 52022 10645 52038 10679
rect 51638 10598 52038 10645
rect 52226 10751 52626 10798
rect 52226 10717 52242 10751
rect 52610 10717 52626 10751
rect 52226 10679 52626 10717
rect 52226 10645 52242 10679
rect 52610 10645 52626 10679
rect 52226 10598 52626 10645
rect 52814 10751 53214 10798
rect 52814 10717 52830 10751
rect 53198 10717 53214 10751
rect 52814 10679 53214 10717
rect 52814 10645 52830 10679
rect 53198 10645 53214 10679
rect 52814 10598 53214 10645
rect 53402 10751 53802 10798
rect 53402 10717 53418 10751
rect 53786 10717 53802 10751
rect 53402 10679 53802 10717
rect 53402 10645 53418 10679
rect 53786 10645 53802 10679
rect 53402 10598 53802 10645
rect 53990 10751 54390 10798
rect 53990 10717 54006 10751
rect 54374 10717 54390 10751
rect 53990 10679 54390 10717
rect 53990 10645 54006 10679
rect 54374 10645 54390 10679
rect 53990 10598 54390 10645
rect 54578 10751 54978 10798
rect 54578 10717 54594 10751
rect 54962 10717 54978 10751
rect 54578 10679 54978 10717
rect 54578 10645 54594 10679
rect 54962 10645 54978 10679
rect 54578 10598 54978 10645
rect 55166 10751 55566 10798
rect 55166 10717 55182 10751
rect 55550 10717 55566 10751
rect 55166 10679 55566 10717
rect 55166 10645 55182 10679
rect 55550 10645 55566 10679
rect 55166 10598 55566 10645
rect 55754 10751 56154 10798
rect 55754 10717 55770 10751
rect 56138 10717 56154 10751
rect 55754 10679 56154 10717
rect 55754 10645 55770 10679
rect 56138 10645 56154 10679
rect 55754 10598 56154 10645
rect 56342 10751 56742 10798
rect 56342 10717 56358 10751
rect 56726 10717 56742 10751
rect 56342 10679 56742 10717
rect 56342 10645 56358 10679
rect 56726 10645 56742 10679
rect 56342 10598 56742 10645
rect 56930 10751 57330 10798
rect 56930 10717 56946 10751
rect 57314 10717 57330 10751
rect 56930 10679 57330 10717
rect 56930 10645 56946 10679
rect 57314 10645 57330 10679
rect 56930 10598 57330 10645
rect 57518 10751 57918 10798
rect 57518 10717 57534 10751
rect 57902 10717 57918 10751
rect 57518 10679 57918 10717
rect 57518 10645 57534 10679
rect 57902 10645 57918 10679
rect 57518 10598 57918 10645
rect 58106 10751 58506 10798
rect 58106 10717 58122 10751
rect 58490 10717 58506 10751
rect 58106 10679 58506 10717
rect 58106 10645 58122 10679
rect 58490 10645 58506 10679
rect 58106 10598 58506 10645
rect 58694 10751 59094 10798
rect 58694 10717 58710 10751
rect 59078 10717 59094 10751
rect 58694 10679 59094 10717
rect 58694 10645 58710 10679
rect 59078 10645 59094 10679
rect 58694 10598 59094 10645
rect 59282 10751 59682 10798
rect 59282 10717 59298 10751
rect 59666 10717 59682 10751
rect 59282 10679 59682 10717
rect 59282 10645 59298 10679
rect 59666 10645 59682 10679
rect 59282 10598 59682 10645
rect 59870 10751 60270 10798
rect 59870 10717 59886 10751
rect 60254 10717 60270 10751
rect 59870 10679 60270 10717
rect 59870 10645 59886 10679
rect 60254 10645 60270 10679
rect 59870 10598 60270 10645
rect 60458 10751 60858 10798
rect 60458 10717 60474 10751
rect 60842 10717 60858 10751
rect 60458 10679 60858 10717
rect 60458 10645 60474 10679
rect 60842 10645 60858 10679
rect 60458 10598 60858 10645
rect 61046 10751 61446 10798
rect 61046 10717 61062 10751
rect 61430 10717 61446 10751
rect 61046 10679 61446 10717
rect 61046 10645 61062 10679
rect 61430 10645 61446 10679
rect 61046 10598 61446 10645
rect 61634 10751 62034 10798
rect 61634 10717 61650 10751
rect 62018 10717 62034 10751
rect 61634 10679 62034 10717
rect 61634 10645 61650 10679
rect 62018 10645 62034 10679
rect 61634 10598 62034 10645
rect 62222 10751 62622 10798
rect 62222 10717 62238 10751
rect 62606 10717 62622 10751
rect 62222 10679 62622 10717
rect 62222 10645 62238 10679
rect 62606 10645 62622 10679
rect 62222 10598 62622 10645
rect 62810 10751 63210 10798
rect 62810 10717 62826 10751
rect 63194 10717 63210 10751
rect 62810 10679 63210 10717
rect 62810 10645 62826 10679
rect 63194 10645 63210 10679
rect 62810 10598 63210 10645
rect 63398 10751 63798 10798
rect 63398 10717 63414 10751
rect 63782 10717 63798 10751
rect 63398 10679 63798 10717
rect 63398 10645 63414 10679
rect 63782 10645 63798 10679
rect 63398 10598 63798 10645
rect 63986 10751 64386 10798
rect 63986 10717 64002 10751
rect 64370 10717 64386 10751
rect 63986 10679 64386 10717
rect 63986 10645 64002 10679
rect 64370 10645 64386 10679
rect 63986 10598 64386 10645
rect 64574 10751 64974 10798
rect 64574 10717 64590 10751
rect 64958 10717 64974 10751
rect 64574 10679 64974 10717
rect 64574 10645 64590 10679
rect 64958 10645 64974 10679
rect 64574 10598 64974 10645
rect 65162 10751 65562 10798
rect 65162 10717 65178 10751
rect 65546 10717 65562 10751
rect 65162 10679 65562 10717
rect 65162 10645 65178 10679
rect 65546 10645 65562 10679
rect 65162 10598 65562 10645
rect 65750 10751 66150 10798
rect 65750 10717 65766 10751
rect 66134 10717 66150 10751
rect 65750 10679 66150 10717
rect 65750 10645 65766 10679
rect 66134 10645 66150 10679
rect 65750 10598 66150 10645
rect 66338 10751 66738 10798
rect 66338 10717 66354 10751
rect 66722 10717 66738 10751
rect 66338 10679 66738 10717
rect 66338 10645 66354 10679
rect 66722 10645 66738 10679
rect 66338 10598 66738 10645
rect 66926 10751 67326 10798
rect 66926 10717 66942 10751
rect 67310 10717 67326 10751
rect 66926 10679 67326 10717
rect 66926 10645 66942 10679
rect 67310 10645 67326 10679
rect 66926 10598 67326 10645
rect 67514 10751 67914 10798
rect 67514 10717 67530 10751
rect 67898 10717 67914 10751
rect 67514 10679 67914 10717
rect 67514 10645 67530 10679
rect 67898 10645 67914 10679
rect 67514 10598 67914 10645
rect 68102 10751 68502 10798
rect 68102 10717 68118 10751
rect 68486 10717 68502 10751
rect 68102 10679 68502 10717
rect 68102 10645 68118 10679
rect 68486 10645 68502 10679
rect 68102 10598 68502 10645
rect 68690 10751 69090 10798
rect 68690 10717 68706 10751
rect 69074 10717 69090 10751
rect 68690 10679 69090 10717
rect 68690 10645 68706 10679
rect 69074 10645 69090 10679
rect 68690 10598 69090 10645
rect 69278 10751 69678 10798
rect 69278 10717 69294 10751
rect 69662 10717 69678 10751
rect 69278 10679 69678 10717
rect 69278 10645 69294 10679
rect 69662 10645 69678 10679
rect 69278 10598 69678 10645
rect 69866 10751 70266 10798
rect 69866 10717 69882 10751
rect 70250 10717 70266 10751
rect 69866 10679 70266 10717
rect 69866 10645 69882 10679
rect 70250 10645 70266 10679
rect 69866 10598 70266 10645
rect 70454 10751 70854 10798
rect 70454 10717 70470 10751
rect 70838 10717 70854 10751
rect 70454 10679 70854 10717
rect 70454 10645 70470 10679
rect 70838 10645 70854 10679
rect 70454 10598 70854 10645
rect 71042 10751 71442 10798
rect 71042 10717 71058 10751
rect 71426 10717 71442 10751
rect 71042 10679 71442 10717
rect 71042 10645 71058 10679
rect 71426 10645 71442 10679
rect 71042 10598 71442 10645
rect 43406 9751 43806 9798
rect 43406 9717 43422 9751
rect 43790 9717 43806 9751
rect 43406 9701 43806 9717
rect 43994 9751 44394 9798
rect 43994 9717 44010 9751
rect 44378 9717 44394 9751
rect 43994 9701 44394 9717
rect 44582 9751 44982 9798
rect 44582 9717 44598 9751
rect 44966 9717 44982 9751
rect 44582 9701 44982 9717
rect 45170 9751 45570 9798
rect 45170 9717 45186 9751
rect 45554 9717 45570 9751
rect 45170 9701 45570 9717
rect 45758 9751 46158 9798
rect 45758 9717 45774 9751
rect 46142 9717 46158 9751
rect 45758 9701 46158 9717
rect 46346 9751 46746 9798
rect 46346 9717 46362 9751
rect 46730 9717 46746 9751
rect 46346 9701 46746 9717
rect 46934 9751 47334 9798
rect 46934 9717 46950 9751
rect 47318 9717 47334 9751
rect 46934 9701 47334 9717
rect 47522 9751 47922 9798
rect 47522 9717 47538 9751
rect 47906 9717 47922 9751
rect 47522 9701 47922 9717
rect 48110 9751 48510 9798
rect 48110 9717 48126 9751
rect 48494 9717 48510 9751
rect 48110 9701 48510 9717
rect 48698 9751 49098 9798
rect 48698 9717 48714 9751
rect 49082 9717 49098 9751
rect 48698 9701 49098 9717
rect 49286 9751 49686 9798
rect 49286 9717 49302 9751
rect 49670 9717 49686 9751
rect 49286 9701 49686 9717
rect 49874 9751 50274 9798
rect 49874 9717 49890 9751
rect 50258 9717 50274 9751
rect 49874 9701 50274 9717
rect 50462 9751 50862 9798
rect 50462 9717 50478 9751
rect 50846 9717 50862 9751
rect 50462 9701 50862 9717
rect 51050 9751 51450 9798
rect 51050 9717 51066 9751
rect 51434 9717 51450 9751
rect 51050 9701 51450 9717
rect 51638 9751 52038 9798
rect 51638 9717 51654 9751
rect 52022 9717 52038 9751
rect 51638 9701 52038 9717
rect 52226 9751 52626 9798
rect 52226 9717 52242 9751
rect 52610 9717 52626 9751
rect 52226 9701 52626 9717
rect 52814 9751 53214 9798
rect 52814 9717 52830 9751
rect 53198 9717 53214 9751
rect 52814 9701 53214 9717
rect 53402 9751 53802 9798
rect 53402 9717 53418 9751
rect 53786 9717 53802 9751
rect 53402 9701 53802 9717
rect 53990 9751 54390 9798
rect 53990 9717 54006 9751
rect 54374 9717 54390 9751
rect 53990 9701 54390 9717
rect 54578 9751 54978 9798
rect 54578 9717 54594 9751
rect 54962 9717 54978 9751
rect 54578 9701 54978 9717
rect 55166 9751 55566 9798
rect 55166 9717 55182 9751
rect 55550 9717 55566 9751
rect 55166 9701 55566 9717
rect 55754 9751 56154 9798
rect 55754 9717 55770 9751
rect 56138 9717 56154 9751
rect 55754 9701 56154 9717
rect 56342 9751 56742 9798
rect 56342 9717 56358 9751
rect 56726 9717 56742 9751
rect 56342 9701 56742 9717
rect 56930 9751 57330 9798
rect 56930 9717 56946 9751
rect 57314 9717 57330 9751
rect 56930 9701 57330 9717
rect 57518 9751 57918 9798
rect 57518 9717 57534 9751
rect 57902 9717 57918 9751
rect 57518 9701 57918 9717
rect 58106 9751 58506 9798
rect 58106 9717 58122 9751
rect 58490 9717 58506 9751
rect 58106 9701 58506 9717
rect 58694 9751 59094 9798
rect 58694 9717 58710 9751
rect 59078 9717 59094 9751
rect 58694 9701 59094 9717
rect 59282 9751 59682 9798
rect 59282 9717 59298 9751
rect 59666 9717 59682 9751
rect 59282 9701 59682 9717
rect 59870 9751 60270 9798
rect 59870 9717 59886 9751
rect 60254 9717 60270 9751
rect 59870 9701 60270 9717
rect 60458 9751 60858 9798
rect 60458 9717 60474 9751
rect 60842 9717 60858 9751
rect 60458 9701 60858 9717
rect 61046 9751 61446 9798
rect 61046 9717 61062 9751
rect 61430 9717 61446 9751
rect 61046 9701 61446 9717
rect 61634 9751 62034 9798
rect 61634 9717 61650 9751
rect 62018 9717 62034 9751
rect 61634 9701 62034 9717
rect 62222 9751 62622 9798
rect 62222 9717 62238 9751
rect 62606 9717 62622 9751
rect 62222 9701 62622 9717
rect 62810 9751 63210 9798
rect 62810 9717 62826 9751
rect 63194 9717 63210 9751
rect 62810 9701 63210 9717
rect 63398 9751 63798 9798
rect 63398 9717 63414 9751
rect 63782 9717 63798 9751
rect 63398 9701 63798 9717
rect 63986 9751 64386 9798
rect 63986 9717 64002 9751
rect 64370 9717 64386 9751
rect 63986 9701 64386 9717
rect 64574 9751 64974 9798
rect 64574 9717 64590 9751
rect 64958 9717 64974 9751
rect 64574 9701 64974 9717
rect 65162 9751 65562 9798
rect 65162 9717 65178 9751
rect 65546 9717 65562 9751
rect 65162 9701 65562 9717
rect 65750 9751 66150 9798
rect 65750 9717 65766 9751
rect 66134 9717 66150 9751
rect 65750 9701 66150 9717
rect 66338 9751 66738 9798
rect 66338 9717 66354 9751
rect 66722 9717 66738 9751
rect 66338 9701 66738 9717
rect 66926 9751 67326 9798
rect 66926 9717 66942 9751
rect 67310 9717 67326 9751
rect 66926 9701 67326 9717
rect 67514 9751 67914 9798
rect 67514 9717 67530 9751
rect 67898 9717 67914 9751
rect 67514 9701 67914 9717
rect 68102 9751 68502 9798
rect 68102 9717 68118 9751
rect 68486 9717 68502 9751
rect 68102 9701 68502 9717
rect 68690 9751 69090 9798
rect 68690 9717 68706 9751
rect 69074 9717 69090 9751
rect 68690 9701 69090 9717
rect 69278 9751 69678 9798
rect 69278 9717 69294 9751
rect 69662 9717 69678 9751
rect 69278 9701 69678 9717
rect 69866 9751 70266 9798
rect 69866 9717 69882 9751
rect 70250 9717 70266 9751
rect 69866 9701 70266 9717
rect 70454 9751 70854 9798
rect 70454 9717 70470 9751
rect 70838 9717 70854 9751
rect 70454 9701 70854 9717
rect 71042 9751 71442 9798
rect 71042 9717 71058 9751
rect 71426 9717 71442 9751
rect 71042 9701 71442 9717
rect 56458 8322 56528 8328
rect 56458 8190 56474 8322
rect 56512 8190 56528 8322
rect 56458 8152 56528 8190
rect 56724 8322 56794 8328
rect 56724 8190 56740 8322
rect 56778 8190 56794 8322
rect 56724 8152 56794 8190
rect 56990 8322 57060 8328
rect 56990 8190 57006 8322
rect 57044 8190 57060 8322
rect 56990 8152 57060 8190
rect 57256 8322 57326 8328
rect 57256 8190 57272 8322
rect 57310 8190 57326 8322
rect 57256 8152 57326 8190
rect 57522 8322 57592 8328
rect 57522 8190 57538 8322
rect 57576 8190 57592 8322
rect 57522 8152 57592 8190
rect 57788 8322 57858 8328
rect 57788 8190 57804 8322
rect 57842 8190 57858 8322
rect 57788 8152 57858 8190
rect 58054 8322 58124 8328
rect 58054 8190 58070 8322
rect 58108 8190 58124 8322
rect 58054 8152 58124 8190
rect 58320 8322 58390 8328
rect 58320 8190 58336 8322
rect 58374 8190 58390 8322
rect 58320 8152 58390 8190
rect 56458 7312 56528 7352
rect 56458 7180 56474 7312
rect 56512 7180 56528 7312
rect 56458 7142 56528 7180
rect 56724 7312 56794 7352
rect 56724 7180 56740 7312
rect 56778 7180 56794 7312
rect 56724 7142 56794 7180
rect 56990 7312 57060 7352
rect 56990 7180 57006 7312
rect 57044 7180 57060 7312
rect 56990 7142 57060 7180
rect 57256 7312 57326 7352
rect 57256 7180 57272 7312
rect 57310 7180 57326 7312
rect 57256 7142 57326 7180
rect 57522 7312 57592 7352
rect 57522 7180 57538 7312
rect 57576 7180 57592 7312
rect 57522 7142 57592 7180
rect 57788 7312 57858 7352
rect 57788 7180 57804 7312
rect 57842 7180 57858 7312
rect 57788 7142 57858 7180
rect 58054 7312 58124 7352
rect 58054 7180 58070 7312
rect 58108 7180 58124 7312
rect 58054 7142 58124 7180
rect 58320 7312 58390 7352
rect 58320 7180 58336 7312
rect 58374 7180 58390 7312
rect 58320 7142 58390 7180
rect 56458 6302 56528 6342
rect 56458 6170 56474 6302
rect 56512 6170 56528 6302
rect 56458 6132 56528 6170
rect 56724 6302 56794 6342
rect 56724 6170 56740 6302
rect 56778 6170 56794 6302
rect 56724 6132 56794 6170
rect 56990 6302 57060 6342
rect 56990 6170 57006 6302
rect 57044 6170 57060 6302
rect 56990 6132 57060 6170
rect 57256 6302 57326 6342
rect 57256 6170 57272 6302
rect 57310 6170 57326 6302
rect 57256 6132 57326 6170
rect 57522 6302 57592 6342
rect 57522 6170 57538 6302
rect 57576 6170 57592 6302
rect 57522 6132 57592 6170
rect 57788 6302 57858 6342
rect 57788 6170 57804 6302
rect 57842 6170 57858 6302
rect 57788 6132 57858 6170
rect 58054 6302 58124 6342
rect 58054 6170 58070 6302
rect 58108 6170 58124 6302
rect 58054 6132 58124 6170
rect 58320 6302 58390 6342
rect 58320 6170 58336 6302
rect 58374 6170 58390 6302
rect 58320 6132 58390 6170
rect 56458 5292 56528 5332
rect 56458 5160 56474 5292
rect 56512 5160 56528 5292
rect 56458 5150 56528 5160
rect 56724 5292 56794 5332
rect 56724 5160 56740 5292
rect 56778 5160 56794 5292
rect 56724 5150 56794 5160
rect 56990 5292 57060 5332
rect 56990 5160 57006 5292
rect 57044 5160 57060 5292
rect 56990 5150 57060 5160
rect 57256 5292 57326 5332
rect 57256 5160 57272 5292
rect 57310 5160 57326 5292
rect 57256 5150 57326 5160
rect 57522 5292 57592 5332
rect 57522 5160 57538 5292
rect 57576 5160 57592 5292
rect 57522 5150 57592 5160
rect 57788 5292 57858 5332
rect 57788 5160 57804 5292
rect 57842 5160 57858 5292
rect 57788 5150 57858 5160
rect 58054 5292 58124 5332
rect 58054 5160 58070 5292
rect 58108 5160 58124 5292
rect 58054 5150 58124 5160
rect 58320 5292 58390 5332
rect 58320 5160 58336 5292
rect 58374 5160 58390 5292
rect 58320 5150 58390 5160
rect 57030 4124 57100 4130
rect 57030 3998 57046 4124
rect 57084 3998 57100 4124
rect 57030 3960 57100 3998
rect 57270 4124 57340 4130
rect 57270 3998 57286 4124
rect 57324 3998 57340 4124
rect 57270 3960 57340 3998
rect 57510 4124 57580 4130
rect 57510 3998 57526 4124
rect 57564 3998 57580 4124
rect 57510 3960 57580 3998
rect 57750 4124 57820 4130
rect 57750 3998 57766 4124
rect 57804 3998 57820 4124
rect 57750 3960 57820 3998
rect 57030 3322 57100 3360
rect 57030 3190 57046 3322
rect 57084 3190 57100 3322
rect 57030 3152 57100 3190
rect 57270 3322 57340 3360
rect 57270 3190 57286 3322
rect 57324 3190 57340 3322
rect 57270 3152 57340 3190
rect 57510 3322 57580 3360
rect 57510 3190 57526 3322
rect 57564 3190 57580 3322
rect 57510 3152 57580 3190
rect 57750 3322 57820 3360
rect 57750 3190 57766 3322
rect 57804 3190 57820 3322
rect 57750 3152 57820 3190
rect 57030 2514 57100 2552
rect 57030 2382 57046 2514
rect 57084 2382 57100 2514
rect 57270 2514 57340 2552
rect 57270 2382 57286 2514
rect 57324 2382 57340 2514
rect 57510 2514 57580 2552
rect 57510 2382 57526 2514
rect 57564 2382 57580 2514
rect 57750 2514 57820 2552
rect 57750 2382 57766 2514
rect 57804 2382 57820 2514
<< polycont >>
rect 52726 16710 52764 16842
rect 52966 16710 53004 16842
rect 53206 16710 53244 16842
rect 53446 16710 53484 16842
rect 53686 16710 53724 16842
rect 53926 16710 53964 16842
rect 54166 16710 54204 16842
rect 54406 16710 54444 16842
rect 54646 16710 54684 16842
rect 54886 16710 54924 16842
rect 55126 16710 55164 16842
rect 55366 16710 55404 16842
rect 55606 16710 55644 16842
rect 55846 16710 55884 16842
rect 56086 16710 56124 16842
rect 56326 16710 56364 16842
rect 56566 16710 56604 16842
rect 56806 16710 56844 16842
rect 57046 16710 57084 16842
rect 57286 16710 57324 16842
rect 57526 16710 57564 16842
rect 57766 16710 57804 16842
rect 58006 16710 58044 16842
rect 58246 16710 58284 16842
rect 58486 16710 58524 16842
rect 58726 16710 58764 16842
rect 58966 16710 59004 16842
rect 59206 16710 59244 16842
rect 59446 16710 59484 16842
rect 59686 16710 59724 16842
rect 59926 16710 59964 16842
rect 60166 16710 60204 16842
rect 60406 16710 60444 16842
rect 60646 16710 60684 16842
rect 60886 16710 60924 16842
rect 61126 16710 61164 16842
rect 61366 16710 61404 16842
rect 61606 16710 61644 16842
rect 61846 16710 61884 16842
rect 62086 16710 62124 16842
rect 52726 15902 52764 16034
rect 52966 15902 53004 16034
rect 53206 15902 53244 16034
rect 53446 15902 53484 16034
rect 53686 15902 53724 16034
rect 53926 15902 53964 16034
rect 54166 15902 54204 16034
rect 54406 15902 54444 16034
rect 54646 15902 54684 16034
rect 54886 15902 54924 16034
rect 55126 15902 55164 16034
rect 55366 15902 55404 16034
rect 55606 15902 55644 16034
rect 55846 15902 55884 16034
rect 56086 15902 56124 16034
rect 56326 15902 56364 16034
rect 56566 15902 56604 16034
rect 56806 15902 56844 16034
rect 57046 15902 57084 16034
rect 57286 15902 57324 16034
rect 57526 15902 57564 16034
rect 57766 15902 57804 16034
rect 58006 15902 58044 16034
rect 58246 15902 58284 16034
rect 58486 15902 58524 16034
rect 58726 15902 58764 16034
rect 58966 15902 59004 16034
rect 59206 15902 59244 16034
rect 59446 15902 59484 16034
rect 59686 15902 59724 16034
rect 59926 15902 59964 16034
rect 60166 15902 60204 16034
rect 60406 15902 60444 16034
rect 60646 15902 60684 16034
rect 60886 15902 60924 16034
rect 61126 15902 61164 16034
rect 61366 15902 61404 16034
rect 61606 15902 61644 16034
rect 61846 15902 61884 16034
rect 62086 15902 62124 16034
rect 52726 15094 52764 15226
rect 52966 15094 53004 15226
rect 53206 15094 53244 15226
rect 53446 15094 53484 15226
rect 53686 15094 53724 15226
rect 53926 15094 53964 15226
rect 54166 15094 54204 15226
rect 54406 15094 54444 15226
rect 54646 15094 54684 15226
rect 54886 15094 54924 15226
rect 55126 15094 55164 15226
rect 55366 15094 55404 15226
rect 55606 15094 55644 15226
rect 55846 15094 55884 15226
rect 56086 15094 56124 15226
rect 56326 15094 56364 15226
rect 56566 15094 56604 15226
rect 56806 15094 56844 15226
rect 57046 15094 57084 15226
rect 57286 15094 57324 15226
rect 57526 15094 57564 15226
rect 57766 15094 57804 15226
rect 58006 15094 58044 15226
rect 58246 15094 58284 15226
rect 58486 15094 58524 15226
rect 58726 15094 58764 15226
rect 58966 15094 59004 15226
rect 59206 15094 59244 15226
rect 59446 15094 59484 15226
rect 59686 15094 59724 15226
rect 59926 15094 59964 15226
rect 60166 15094 60204 15226
rect 60406 15094 60444 15226
rect 60646 15094 60684 15226
rect 60886 15094 60924 15226
rect 61126 15094 61164 15226
rect 61366 15094 61404 15226
rect 61606 15094 61644 15226
rect 61846 15094 61884 15226
rect 62086 15094 62124 15226
rect 43422 12645 43790 12679
rect 44010 12645 44378 12679
rect 44598 12645 44966 12679
rect 45186 12645 45554 12679
rect 45774 12645 46142 12679
rect 46362 12645 46730 12679
rect 46950 12645 47318 12679
rect 47538 12645 47906 12679
rect 48126 12645 48494 12679
rect 48714 12645 49082 12679
rect 49302 12645 49670 12679
rect 49890 12645 50258 12679
rect 50478 12645 50846 12679
rect 51066 12645 51434 12679
rect 51654 12645 52022 12679
rect 52242 12645 52610 12679
rect 52830 12645 53198 12679
rect 53418 12645 53786 12679
rect 54006 12645 54374 12679
rect 54594 12645 54962 12679
rect 55182 12645 55550 12679
rect 55770 12645 56138 12679
rect 56358 12645 56726 12679
rect 56946 12645 57314 12679
rect 57534 12645 57902 12679
rect 58122 12645 58490 12679
rect 58710 12645 59078 12679
rect 59298 12645 59666 12679
rect 59886 12645 60254 12679
rect 60474 12645 60842 12679
rect 61062 12645 61430 12679
rect 61650 12645 62018 12679
rect 62238 12645 62606 12679
rect 62826 12645 63194 12679
rect 63414 12645 63782 12679
rect 64002 12645 64370 12679
rect 64590 12645 64958 12679
rect 65178 12645 65546 12679
rect 65766 12645 66134 12679
rect 66354 12645 66722 12679
rect 66942 12645 67310 12679
rect 67530 12645 67898 12679
rect 68118 12645 68486 12679
rect 68706 12645 69074 12679
rect 69294 12645 69662 12679
rect 69882 12645 70250 12679
rect 70470 12645 70838 12679
rect 71058 12645 71426 12679
rect 43422 11717 43790 11751
rect 43422 11645 43790 11679
rect 44010 11717 44378 11751
rect 44010 11645 44378 11679
rect 44598 11717 44966 11751
rect 44598 11645 44966 11679
rect 45186 11717 45554 11751
rect 45186 11645 45554 11679
rect 45774 11717 46142 11751
rect 45774 11645 46142 11679
rect 46362 11717 46730 11751
rect 46362 11645 46730 11679
rect 46950 11717 47318 11751
rect 46950 11645 47318 11679
rect 47538 11717 47906 11751
rect 47538 11645 47906 11679
rect 48126 11717 48494 11751
rect 48126 11645 48494 11679
rect 48714 11717 49082 11751
rect 48714 11645 49082 11679
rect 49302 11717 49670 11751
rect 49302 11645 49670 11679
rect 49890 11717 50258 11751
rect 49890 11645 50258 11679
rect 50478 11717 50846 11751
rect 50478 11645 50846 11679
rect 51066 11717 51434 11751
rect 51066 11645 51434 11679
rect 51654 11717 52022 11751
rect 51654 11645 52022 11679
rect 52242 11717 52610 11751
rect 52242 11645 52610 11679
rect 52830 11717 53198 11751
rect 52830 11645 53198 11679
rect 53418 11717 53786 11751
rect 53418 11645 53786 11679
rect 54006 11717 54374 11751
rect 54006 11645 54374 11679
rect 54594 11717 54962 11751
rect 54594 11645 54962 11679
rect 55182 11717 55550 11751
rect 55182 11645 55550 11679
rect 55770 11717 56138 11751
rect 55770 11645 56138 11679
rect 56358 11717 56726 11751
rect 56358 11645 56726 11679
rect 56946 11717 57314 11751
rect 56946 11645 57314 11679
rect 57534 11717 57902 11751
rect 57534 11645 57902 11679
rect 58122 11717 58490 11751
rect 58122 11645 58490 11679
rect 58710 11717 59078 11751
rect 58710 11645 59078 11679
rect 59298 11717 59666 11751
rect 59298 11645 59666 11679
rect 59886 11717 60254 11751
rect 59886 11645 60254 11679
rect 60474 11717 60842 11751
rect 60474 11645 60842 11679
rect 61062 11717 61430 11751
rect 61062 11645 61430 11679
rect 61650 11717 62018 11751
rect 61650 11645 62018 11679
rect 62238 11717 62606 11751
rect 62238 11645 62606 11679
rect 62826 11717 63194 11751
rect 62826 11645 63194 11679
rect 63414 11717 63782 11751
rect 63414 11645 63782 11679
rect 64002 11717 64370 11751
rect 64002 11645 64370 11679
rect 64590 11717 64958 11751
rect 64590 11645 64958 11679
rect 65178 11717 65546 11751
rect 65178 11645 65546 11679
rect 65766 11717 66134 11751
rect 65766 11645 66134 11679
rect 66354 11717 66722 11751
rect 66354 11645 66722 11679
rect 66942 11717 67310 11751
rect 66942 11645 67310 11679
rect 67530 11717 67898 11751
rect 67530 11645 67898 11679
rect 68118 11717 68486 11751
rect 68118 11645 68486 11679
rect 68706 11717 69074 11751
rect 68706 11645 69074 11679
rect 69294 11717 69662 11751
rect 69294 11645 69662 11679
rect 69882 11717 70250 11751
rect 69882 11645 70250 11679
rect 70470 11717 70838 11751
rect 70470 11645 70838 11679
rect 71058 11717 71426 11751
rect 71058 11645 71426 11679
rect 43422 10717 43790 10751
rect 43422 10645 43790 10679
rect 44010 10717 44378 10751
rect 44010 10645 44378 10679
rect 44598 10717 44966 10751
rect 44598 10645 44966 10679
rect 45186 10717 45554 10751
rect 45186 10645 45554 10679
rect 45774 10717 46142 10751
rect 45774 10645 46142 10679
rect 46362 10717 46730 10751
rect 46362 10645 46730 10679
rect 46950 10717 47318 10751
rect 46950 10645 47318 10679
rect 47538 10717 47906 10751
rect 47538 10645 47906 10679
rect 48126 10717 48494 10751
rect 48126 10645 48494 10679
rect 48714 10717 49082 10751
rect 48714 10645 49082 10679
rect 49302 10717 49670 10751
rect 49302 10645 49670 10679
rect 49890 10717 50258 10751
rect 49890 10645 50258 10679
rect 50478 10717 50846 10751
rect 50478 10645 50846 10679
rect 51066 10717 51434 10751
rect 51066 10645 51434 10679
rect 51654 10717 52022 10751
rect 51654 10645 52022 10679
rect 52242 10717 52610 10751
rect 52242 10645 52610 10679
rect 52830 10717 53198 10751
rect 52830 10645 53198 10679
rect 53418 10717 53786 10751
rect 53418 10645 53786 10679
rect 54006 10717 54374 10751
rect 54006 10645 54374 10679
rect 54594 10717 54962 10751
rect 54594 10645 54962 10679
rect 55182 10717 55550 10751
rect 55182 10645 55550 10679
rect 55770 10717 56138 10751
rect 55770 10645 56138 10679
rect 56358 10717 56726 10751
rect 56358 10645 56726 10679
rect 56946 10717 57314 10751
rect 56946 10645 57314 10679
rect 57534 10717 57902 10751
rect 57534 10645 57902 10679
rect 58122 10717 58490 10751
rect 58122 10645 58490 10679
rect 58710 10717 59078 10751
rect 58710 10645 59078 10679
rect 59298 10717 59666 10751
rect 59298 10645 59666 10679
rect 59886 10717 60254 10751
rect 59886 10645 60254 10679
rect 60474 10717 60842 10751
rect 60474 10645 60842 10679
rect 61062 10717 61430 10751
rect 61062 10645 61430 10679
rect 61650 10717 62018 10751
rect 61650 10645 62018 10679
rect 62238 10717 62606 10751
rect 62238 10645 62606 10679
rect 62826 10717 63194 10751
rect 62826 10645 63194 10679
rect 63414 10717 63782 10751
rect 63414 10645 63782 10679
rect 64002 10717 64370 10751
rect 64002 10645 64370 10679
rect 64590 10717 64958 10751
rect 64590 10645 64958 10679
rect 65178 10717 65546 10751
rect 65178 10645 65546 10679
rect 65766 10717 66134 10751
rect 65766 10645 66134 10679
rect 66354 10717 66722 10751
rect 66354 10645 66722 10679
rect 66942 10717 67310 10751
rect 66942 10645 67310 10679
rect 67530 10717 67898 10751
rect 67530 10645 67898 10679
rect 68118 10717 68486 10751
rect 68118 10645 68486 10679
rect 68706 10717 69074 10751
rect 68706 10645 69074 10679
rect 69294 10717 69662 10751
rect 69294 10645 69662 10679
rect 69882 10717 70250 10751
rect 69882 10645 70250 10679
rect 70470 10717 70838 10751
rect 70470 10645 70838 10679
rect 71058 10717 71426 10751
rect 71058 10645 71426 10679
rect 43422 9717 43790 9751
rect 44010 9717 44378 9751
rect 44598 9717 44966 9751
rect 45186 9717 45554 9751
rect 45774 9717 46142 9751
rect 46362 9717 46730 9751
rect 46950 9717 47318 9751
rect 47538 9717 47906 9751
rect 48126 9717 48494 9751
rect 48714 9717 49082 9751
rect 49302 9717 49670 9751
rect 49890 9717 50258 9751
rect 50478 9717 50846 9751
rect 51066 9717 51434 9751
rect 51654 9717 52022 9751
rect 52242 9717 52610 9751
rect 52830 9717 53198 9751
rect 53418 9717 53786 9751
rect 54006 9717 54374 9751
rect 54594 9717 54962 9751
rect 55182 9717 55550 9751
rect 55770 9717 56138 9751
rect 56358 9717 56726 9751
rect 56946 9717 57314 9751
rect 57534 9717 57902 9751
rect 58122 9717 58490 9751
rect 58710 9717 59078 9751
rect 59298 9717 59666 9751
rect 59886 9717 60254 9751
rect 60474 9717 60842 9751
rect 61062 9717 61430 9751
rect 61650 9717 62018 9751
rect 62238 9717 62606 9751
rect 62826 9717 63194 9751
rect 63414 9717 63782 9751
rect 64002 9717 64370 9751
rect 64590 9717 64958 9751
rect 65178 9717 65546 9751
rect 65766 9717 66134 9751
rect 66354 9717 66722 9751
rect 66942 9717 67310 9751
rect 67530 9717 67898 9751
rect 68118 9717 68486 9751
rect 68706 9717 69074 9751
rect 69294 9717 69662 9751
rect 69882 9717 70250 9751
rect 70470 9717 70838 9751
rect 71058 9717 71426 9751
rect 56474 8190 56512 8322
rect 56740 8190 56778 8322
rect 57006 8190 57044 8322
rect 57272 8190 57310 8322
rect 57538 8190 57576 8322
rect 57804 8190 57842 8322
rect 58070 8190 58108 8322
rect 58336 8190 58374 8322
rect 56474 7180 56512 7312
rect 56740 7180 56778 7312
rect 57006 7180 57044 7312
rect 57272 7180 57310 7312
rect 57538 7180 57576 7312
rect 57804 7180 57842 7312
rect 58070 7180 58108 7312
rect 58336 7180 58374 7312
rect 56474 6170 56512 6302
rect 56740 6170 56778 6302
rect 57006 6170 57044 6302
rect 57272 6170 57310 6302
rect 57538 6170 57576 6302
rect 57804 6170 57842 6302
rect 58070 6170 58108 6302
rect 58336 6170 58374 6302
rect 56474 5160 56512 5292
rect 56740 5160 56778 5292
rect 57006 5160 57044 5292
rect 57272 5160 57310 5292
rect 57538 5160 57576 5292
rect 57804 5160 57842 5292
rect 58070 5160 58108 5292
rect 58336 5160 58374 5292
rect 57046 3998 57084 4124
rect 57286 3998 57324 4124
rect 57526 3998 57564 4124
rect 57766 3998 57804 4124
rect 57046 3190 57084 3322
rect 57286 3190 57324 3322
rect 57526 3190 57564 3322
rect 57766 3190 57804 3322
rect 57046 2382 57084 2514
rect 57286 2382 57324 2514
rect 57526 2382 57564 2514
rect 57766 2382 57804 2514
<< locali >>
rect 52318 17152 52406 17186
rect 62444 17152 62532 17186
rect 52318 17118 52352 17152
rect 62498 17120 62532 17152
rect 52710 16710 52726 16842
rect 52764 16710 52966 16842
rect 53004 16710 53206 16842
rect 53244 16710 53446 16842
rect 53484 16710 53686 16842
rect 53724 16710 53926 16842
rect 53964 16710 54166 16842
rect 54204 16710 54406 16842
rect 54444 16710 54646 16842
rect 54684 16710 54886 16842
rect 54924 16710 55126 16842
rect 55164 16710 55366 16842
rect 55404 16710 55606 16842
rect 55644 16710 55846 16842
rect 55884 16710 56086 16842
rect 56124 16710 56326 16842
rect 56364 16710 56566 16842
rect 56604 16710 56806 16842
rect 56844 16710 57046 16842
rect 57084 16710 57286 16842
rect 57324 16710 57526 16842
rect 57564 16710 57766 16842
rect 57804 16710 58006 16842
rect 58044 16710 58246 16842
rect 58284 16710 58486 16842
rect 58524 16710 58726 16842
rect 58764 16710 58966 16842
rect 59004 16710 59206 16842
rect 59244 16710 59446 16842
rect 59484 16710 59686 16842
rect 59724 16710 59926 16842
rect 59964 16710 60166 16842
rect 60204 16710 60406 16842
rect 60444 16710 60646 16842
rect 60684 16710 60886 16842
rect 60924 16710 61126 16842
rect 61164 16710 61366 16842
rect 61404 16710 61606 16842
rect 61644 16710 61846 16842
rect 61884 16710 62086 16842
rect 62124 16710 62150 16842
rect 52664 16660 52698 16676
rect 52664 16068 52698 16084
rect 52792 16660 52826 16676
rect 52792 16068 52826 16084
rect 52904 16660 52938 16676
rect 52904 16068 52938 16084
rect 53032 16660 53066 16676
rect 53032 16068 53066 16084
rect 53144 16660 53178 16676
rect 53144 16068 53178 16084
rect 53272 16660 53306 16676
rect 53272 16068 53306 16084
rect 53384 16660 53418 16676
rect 53384 16068 53418 16084
rect 53512 16660 53546 16676
rect 53512 16068 53546 16084
rect 53624 16660 53658 16676
rect 53624 16068 53658 16084
rect 53752 16660 53786 16676
rect 53752 16068 53786 16084
rect 53864 16660 53898 16676
rect 53864 16068 53898 16084
rect 53992 16660 54026 16676
rect 53992 16068 54026 16084
rect 54104 16660 54138 16676
rect 54104 16068 54138 16084
rect 54232 16660 54266 16676
rect 54232 16068 54266 16084
rect 54344 16660 54378 16676
rect 54344 16068 54378 16084
rect 54472 16660 54506 16676
rect 54472 16068 54506 16084
rect 54584 16660 54618 16676
rect 54584 16068 54618 16084
rect 54712 16660 54746 16676
rect 54712 16068 54746 16084
rect 54824 16660 54858 16676
rect 54824 16068 54858 16084
rect 54952 16660 54986 16676
rect 54952 16068 54986 16084
rect 55064 16660 55098 16676
rect 55064 16068 55098 16084
rect 55192 16660 55226 16676
rect 55192 16068 55226 16084
rect 55304 16660 55338 16676
rect 55304 16068 55338 16084
rect 55432 16660 55466 16676
rect 55432 16068 55466 16084
rect 55544 16660 55578 16676
rect 55544 16068 55578 16084
rect 55672 16660 55706 16676
rect 55672 16068 55706 16084
rect 55784 16660 55818 16676
rect 55784 16068 55818 16084
rect 55912 16660 55946 16676
rect 55912 16068 55946 16084
rect 56024 16660 56058 16676
rect 56024 16068 56058 16084
rect 56152 16660 56186 16676
rect 56152 16068 56186 16084
rect 56264 16660 56298 16676
rect 56264 16068 56298 16084
rect 56392 16660 56426 16676
rect 56392 16068 56426 16084
rect 56504 16660 56538 16676
rect 56504 16068 56538 16084
rect 56632 16660 56666 16676
rect 56632 16068 56666 16084
rect 56744 16660 56778 16676
rect 56744 16068 56778 16084
rect 56872 16660 56906 16676
rect 56872 16068 56906 16084
rect 56984 16660 57018 16676
rect 56984 16068 57018 16084
rect 57112 16660 57146 16676
rect 57112 16068 57146 16084
rect 57224 16660 57258 16676
rect 57224 16068 57258 16084
rect 57352 16660 57386 16676
rect 57352 16068 57386 16084
rect 57464 16660 57498 16676
rect 57464 16068 57498 16084
rect 57592 16660 57626 16676
rect 57592 16068 57626 16084
rect 57704 16660 57738 16676
rect 57704 16068 57738 16084
rect 57832 16660 57866 16676
rect 57832 16068 57866 16084
rect 57944 16660 57978 16676
rect 57944 16068 57978 16084
rect 58072 16660 58106 16676
rect 58072 16068 58106 16084
rect 58184 16660 58218 16676
rect 58184 16068 58218 16084
rect 58312 16660 58346 16676
rect 58312 16068 58346 16084
rect 58424 16660 58458 16676
rect 58424 16068 58458 16084
rect 58552 16660 58586 16676
rect 58552 16068 58586 16084
rect 58664 16660 58698 16676
rect 58664 16068 58698 16084
rect 58792 16660 58826 16676
rect 58792 16068 58826 16084
rect 58904 16660 58938 16676
rect 58904 16068 58938 16084
rect 59032 16660 59066 16676
rect 59032 16068 59066 16084
rect 59144 16660 59178 16676
rect 59144 16068 59178 16084
rect 59272 16660 59306 16676
rect 59272 16068 59306 16084
rect 59384 16660 59418 16676
rect 59384 16068 59418 16084
rect 59512 16660 59546 16676
rect 59512 16068 59546 16084
rect 59624 16660 59658 16676
rect 59624 16068 59658 16084
rect 59752 16660 59786 16676
rect 59752 16068 59786 16084
rect 59864 16660 59898 16676
rect 59864 16068 59898 16084
rect 59992 16660 60026 16676
rect 59992 16068 60026 16084
rect 60104 16660 60138 16676
rect 60104 16068 60138 16084
rect 60232 16660 60266 16676
rect 60232 16068 60266 16084
rect 60344 16660 60378 16676
rect 60344 16068 60378 16084
rect 60472 16660 60506 16676
rect 60472 16068 60506 16084
rect 60584 16660 60618 16676
rect 60584 16068 60618 16084
rect 60712 16660 60746 16676
rect 60712 16068 60746 16084
rect 60824 16660 60858 16676
rect 60824 16068 60858 16084
rect 60952 16660 60986 16676
rect 60952 16068 60986 16084
rect 61064 16660 61098 16676
rect 61064 16068 61098 16084
rect 61192 16660 61226 16676
rect 61192 16068 61226 16084
rect 61304 16660 61338 16676
rect 61304 16068 61338 16084
rect 61432 16660 61466 16676
rect 61432 16068 61466 16084
rect 61544 16660 61578 16676
rect 61544 16068 61578 16084
rect 61672 16660 61706 16676
rect 61672 16068 61706 16084
rect 61784 16660 61818 16676
rect 61784 16068 61818 16084
rect 61912 16660 61946 16676
rect 61912 16068 61946 16084
rect 62024 16660 62058 16676
rect 62024 16068 62058 16084
rect 62152 16660 62186 16676
rect 62152 16068 62186 16084
rect 52710 15902 52726 16034
rect 52764 15902 52966 16034
rect 53004 15902 53206 16034
rect 53244 15902 53446 16034
rect 53484 15902 53686 16034
rect 53724 15902 53926 16034
rect 53964 15902 54166 16034
rect 54204 15902 54406 16034
rect 54444 15902 54646 16034
rect 54684 15902 54886 16034
rect 54924 15902 55126 16034
rect 55164 15902 55366 16034
rect 55404 15902 55606 16034
rect 55644 15902 55846 16034
rect 55884 15902 56086 16034
rect 56124 15902 56326 16034
rect 56364 15902 56566 16034
rect 56604 15902 56806 16034
rect 56844 15902 57046 16034
rect 57084 15902 57286 16034
rect 57324 15902 57526 16034
rect 57564 15902 57766 16034
rect 57804 15902 58006 16034
rect 58044 15902 58246 16034
rect 58284 15902 58486 16034
rect 58524 15902 58726 16034
rect 58764 15902 58966 16034
rect 59004 15902 59206 16034
rect 59244 15902 59446 16034
rect 59484 15902 59686 16034
rect 59724 15902 59926 16034
rect 59964 15902 60166 16034
rect 60204 15902 60406 16034
rect 60444 15902 60646 16034
rect 60684 15902 60886 16034
rect 60924 15902 61126 16034
rect 61164 15902 61366 16034
rect 61404 15902 61606 16034
rect 61644 15902 61846 16034
rect 61884 15902 62086 16034
rect 62124 15902 62150 16034
rect 52664 15852 52698 15868
rect 52664 15260 52698 15276
rect 52792 15852 52826 15868
rect 52792 15260 52826 15276
rect 52904 15852 52938 15868
rect 52904 15260 52938 15276
rect 53032 15852 53066 15868
rect 53032 15260 53066 15276
rect 53144 15852 53178 15868
rect 53144 15260 53178 15276
rect 53272 15852 53306 15868
rect 53272 15260 53306 15276
rect 53384 15852 53418 15868
rect 53384 15260 53418 15276
rect 53512 15852 53546 15868
rect 53512 15260 53546 15276
rect 53624 15852 53658 15868
rect 53624 15260 53658 15276
rect 53752 15852 53786 15868
rect 53752 15260 53786 15276
rect 53864 15852 53898 15868
rect 53864 15260 53898 15276
rect 53992 15852 54026 15868
rect 53992 15260 54026 15276
rect 54104 15852 54138 15868
rect 54104 15260 54138 15276
rect 54232 15852 54266 15868
rect 54232 15260 54266 15276
rect 54344 15852 54378 15868
rect 54344 15260 54378 15276
rect 54472 15852 54506 15868
rect 54472 15260 54506 15276
rect 54584 15852 54618 15868
rect 54584 15260 54618 15276
rect 54712 15852 54746 15868
rect 54712 15260 54746 15276
rect 54824 15852 54858 15868
rect 54824 15260 54858 15276
rect 54952 15852 54986 15868
rect 54952 15260 54986 15276
rect 55064 15852 55098 15868
rect 55064 15260 55098 15276
rect 55192 15852 55226 15868
rect 55192 15260 55226 15276
rect 55304 15852 55338 15868
rect 55304 15260 55338 15276
rect 55432 15852 55466 15868
rect 55432 15260 55466 15276
rect 55544 15852 55578 15868
rect 55544 15260 55578 15276
rect 55672 15852 55706 15868
rect 55672 15260 55706 15276
rect 55784 15852 55818 15868
rect 55784 15260 55818 15276
rect 55912 15852 55946 15868
rect 55912 15260 55946 15276
rect 56024 15852 56058 15868
rect 56024 15260 56058 15276
rect 56152 15852 56186 15868
rect 56152 15260 56186 15276
rect 56264 15852 56298 15868
rect 56264 15260 56298 15276
rect 56392 15852 56426 15868
rect 56392 15260 56426 15276
rect 56504 15852 56538 15868
rect 56504 15260 56538 15276
rect 56632 15852 56666 15868
rect 56632 15260 56666 15276
rect 56744 15852 56778 15868
rect 56744 15260 56778 15276
rect 56872 15852 56906 15868
rect 56872 15260 56906 15276
rect 56984 15852 57018 15868
rect 56984 15260 57018 15276
rect 57112 15852 57146 15868
rect 57112 15260 57146 15276
rect 57224 15852 57258 15868
rect 57224 15260 57258 15276
rect 57352 15852 57386 15868
rect 57352 15260 57386 15276
rect 57464 15852 57498 15868
rect 57464 15260 57498 15276
rect 57592 15852 57626 15868
rect 57592 15260 57626 15276
rect 57704 15852 57738 15868
rect 57704 15260 57738 15276
rect 57832 15852 57866 15868
rect 57832 15260 57866 15276
rect 57944 15852 57978 15868
rect 57944 15260 57978 15276
rect 58072 15852 58106 15868
rect 58072 15260 58106 15276
rect 58184 15852 58218 15868
rect 58184 15260 58218 15276
rect 58312 15852 58346 15868
rect 58312 15260 58346 15276
rect 58424 15852 58458 15868
rect 58424 15260 58458 15276
rect 58552 15852 58586 15868
rect 58552 15260 58586 15276
rect 58664 15852 58698 15868
rect 58664 15260 58698 15276
rect 58792 15852 58826 15868
rect 58792 15260 58826 15276
rect 58904 15852 58938 15868
rect 58904 15260 58938 15276
rect 59032 15852 59066 15868
rect 59032 15260 59066 15276
rect 59144 15852 59178 15868
rect 59144 15260 59178 15276
rect 59272 15852 59306 15868
rect 59272 15260 59306 15276
rect 59384 15852 59418 15868
rect 59384 15260 59418 15276
rect 59512 15852 59546 15868
rect 59512 15260 59546 15276
rect 59624 15852 59658 15868
rect 59624 15260 59658 15276
rect 59752 15852 59786 15868
rect 59752 15260 59786 15276
rect 59864 15852 59898 15868
rect 59864 15260 59898 15276
rect 59992 15852 60026 15868
rect 59992 15260 60026 15276
rect 60104 15852 60138 15868
rect 60104 15260 60138 15276
rect 60232 15852 60266 15868
rect 60232 15260 60266 15276
rect 60344 15852 60378 15868
rect 60344 15260 60378 15276
rect 60472 15852 60506 15868
rect 60472 15260 60506 15276
rect 60584 15852 60618 15868
rect 60584 15260 60618 15276
rect 60712 15852 60746 15868
rect 60712 15260 60746 15276
rect 60824 15852 60858 15868
rect 60824 15260 60858 15276
rect 60952 15852 60986 15868
rect 60952 15260 60986 15276
rect 61064 15852 61098 15868
rect 61064 15260 61098 15276
rect 61192 15852 61226 15868
rect 61192 15260 61226 15276
rect 61304 15852 61338 15868
rect 61304 15260 61338 15276
rect 61432 15852 61466 15868
rect 61432 15260 61466 15276
rect 61544 15852 61578 15868
rect 61544 15260 61578 15276
rect 61672 15852 61706 15868
rect 61672 15260 61706 15276
rect 61784 15852 61818 15868
rect 61784 15260 61818 15276
rect 61912 15852 61946 15868
rect 61912 15260 61946 15276
rect 62024 15852 62058 15868
rect 62024 15260 62058 15276
rect 62152 15852 62186 15868
rect 62152 15260 62186 15276
rect 52710 15094 52726 15226
rect 52764 15094 52966 15226
rect 53004 15094 53206 15226
rect 53244 15094 53446 15226
rect 53484 15094 53686 15226
rect 53724 15094 53926 15226
rect 53964 15094 54166 15226
rect 54204 15094 54406 15226
rect 54444 15094 54646 15226
rect 54684 15094 54886 15226
rect 54924 15094 55126 15226
rect 55164 15094 55366 15226
rect 55404 15094 55606 15226
rect 55644 15094 55846 15226
rect 55884 15094 56086 15226
rect 56124 15094 56326 15226
rect 56364 15094 56566 15226
rect 56604 15094 56806 15226
rect 56844 15094 57046 15226
rect 57084 15094 57286 15226
rect 57324 15094 57526 15226
rect 57564 15094 57766 15226
rect 57804 15094 58006 15226
rect 58044 15094 58246 15226
rect 58284 15094 58486 15226
rect 58524 15094 58726 15226
rect 58764 15094 58966 15226
rect 59004 15094 59206 15226
rect 59244 15094 59446 15226
rect 59484 15094 59686 15226
rect 59724 15094 59926 15226
rect 59964 15094 60166 15226
rect 60204 15094 60406 15226
rect 60444 15094 60646 15226
rect 60684 15094 60886 15226
rect 60924 15094 61126 15226
rect 61164 15094 61366 15226
rect 61404 15094 61606 15226
rect 61644 15094 61846 15226
rect 61884 15094 62086 15226
rect 62124 15094 62150 15226
rect 52318 14750 52352 14838
rect 62498 14750 62532 14838
rect 43014 12996 43174 13030
rect 71696 13002 71834 13030
rect 71696 12996 71800 13002
rect 43014 12968 43048 12996
rect 43406 12679 55166 12680
rect 55566 12679 55754 12680
rect 56154 12679 56342 12680
rect 56742 12679 56930 12680
rect 57330 12679 57518 12680
rect 57918 12679 58106 12680
rect 58506 12679 58694 12680
rect 59094 12679 59282 12680
rect 59682 12679 71442 12680
rect 43406 12645 43422 12679
rect 43790 12645 44010 12679
rect 44378 12645 44598 12679
rect 44966 12645 45186 12679
rect 45554 12645 45774 12679
rect 46142 12645 46362 12679
rect 46730 12645 46950 12679
rect 47318 12645 47538 12679
rect 47906 12645 48126 12679
rect 48494 12645 48714 12679
rect 49082 12645 49302 12679
rect 49670 12645 49890 12679
rect 50258 12645 50478 12679
rect 50846 12645 51066 12679
rect 51434 12645 51654 12679
rect 52022 12645 52242 12679
rect 52610 12645 52830 12679
rect 53198 12645 53418 12679
rect 53786 12645 54006 12679
rect 54374 12645 54594 12679
rect 54962 12645 55182 12679
rect 55550 12645 55770 12679
rect 56138 12645 56358 12679
rect 56726 12645 56946 12679
rect 57314 12645 57534 12679
rect 57902 12645 58122 12679
rect 58490 12645 58710 12679
rect 59078 12645 59298 12679
rect 59666 12645 59886 12679
rect 60254 12645 60474 12679
rect 60842 12645 61062 12679
rect 61430 12645 61650 12679
rect 62018 12645 62238 12679
rect 62606 12645 62826 12679
rect 63194 12645 63414 12679
rect 63782 12645 64002 12679
rect 64370 12645 64590 12679
rect 64958 12645 65178 12679
rect 65546 12645 65766 12679
rect 66134 12645 66354 12679
rect 66722 12645 66942 12679
rect 67310 12645 67530 12679
rect 67898 12645 68118 12679
rect 68486 12645 68706 12679
rect 69074 12645 69294 12679
rect 69662 12645 69882 12679
rect 70250 12645 70470 12679
rect 70838 12645 71058 12679
rect 71426 12645 71442 12679
rect 43406 12644 55166 12645
rect 55566 12644 55754 12645
rect 56154 12644 56342 12645
rect 56742 12644 56930 12645
rect 55120 12602 55166 12644
rect 57330 12602 57518 12645
rect 57918 12644 58106 12645
rect 58506 12644 58694 12645
rect 59094 12644 59282 12645
rect 59682 12644 71442 12645
rect 59682 12602 59728 12644
rect 43360 12586 43394 12602
rect 43360 11794 43394 11810
rect 43818 12586 43852 12602
rect 43818 11794 43852 11810
rect 43948 12586 43982 12602
rect 43948 11794 43982 11810
rect 44406 12586 44440 12602
rect 44406 11794 44440 11810
rect 44536 12586 44570 12602
rect 44536 11794 44570 11810
rect 44994 12586 45028 12602
rect 44994 11794 45028 11810
rect 45124 12586 45158 12602
rect 45124 11794 45158 11810
rect 45582 12586 45616 12602
rect 45582 11794 45616 11810
rect 45712 12586 45746 12602
rect 45712 11794 45746 11810
rect 46170 12586 46204 12602
rect 46170 11794 46204 11810
rect 46300 12586 46334 12602
rect 46300 11794 46334 11810
rect 46758 12586 46792 12602
rect 46758 11794 46792 11810
rect 46888 12586 46922 12602
rect 46888 11794 46922 11810
rect 47346 12586 47380 12602
rect 47346 11794 47380 11810
rect 47476 12586 47510 12602
rect 47476 11794 47510 11810
rect 47934 12586 47968 12602
rect 47934 11794 47968 11810
rect 48064 12586 48098 12602
rect 48064 11794 48098 11810
rect 48522 12586 48556 12602
rect 48522 11794 48556 11810
rect 48652 12586 48686 12602
rect 48652 11794 48686 11810
rect 49110 12586 49144 12602
rect 49110 11794 49144 11810
rect 49240 12586 49274 12602
rect 49240 11794 49274 11810
rect 49698 12586 49732 12602
rect 49698 11794 49732 11810
rect 49828 12586 49862 12602
rect 49828 11794 49862 11810
rect 50286 12586 50320 12602
rect 50286 11794 50320 11810
rect 50416 12586 50450 12602
rect 50416 11794 50450 11810
rect 50874 12586 50908 12602
rect 50874 11794 50908 11810
rect 51004 12586 51038 12602
rect 51004 11794 51038 11810
rect 51462 12586 51496 12602
rect 51462 11794 51496 11810
rect 51592 12586 51626 12602
rect 51592 11794 51626 11810
rect 52050 12586 52084 12602
rect 52050 11794 52084 11810
rect 52180 12586 52214 12602
rect 52180 11794 52214 11810
rect 52638 12586 52672 12602
rect 52638 11794 52672 11810
rect 52768 12586 52802 12602
rect 52768 11794 52802 11810
rect 53226 12586 53260 12602
rect 53226 11794 53260 11810
rect 53356 12586 53390 12602
rect 53356 11794 53390 11810
rect 53814 12586 53848 12602
rect 53814 11794 53848 11810
rect 53944 12586 53978 12602
rect 53944 11794 53978 11810
rect 54402 12586 54436 12602
rect 54402 11794 54436 11810
rect 54532 12586 54566 12602
rect 54532 11794 54566 11810
rect 54990 12586 55024 12602
rect 54990 11794 55024 11810
rect 55120 12586 55154 12602
rect 55120 11752 55154 11810
rect 55578 12586 55612 12602
rect 55578 11794 55612 11810
rect 55708 12586 55742 12602
rect 55708 11794 55742 11810
rect 56166 12586 56200 12602
rect 56166 11794 56200 11810
rect 56296 12586 56330 12602
rect 56296 11794 56330 11810
rect 56754 12586 56788 12602
rect 56754 11794 56788 11810
rect 56884 12586 56918 12602
rect 56884 11794 56918 11810
rect 57342 12586 57506 12602
rect 57376 11810 57472 12586
rect 57342 11752 57506 11810
rect 57930 12586 57964 12602
rect 57930 11794 57964 11810
rect 58060 12586 58094 12602
rect 58060 11794 58094 11810
rect 58518 12586 58552 12602
rect 58518 11794 58552 11810
rect 58648 12586 58682 12602
rect 58648 11794 58682 11810
rect 59106 12586 59140 12602
rect 59106 11794 59140 11810
rect 59236 12586 59270 12602
rect 59236 11794 59270 11810
rect 59694 12586 59728 12602
rect 59694 11752 59728 11810
rect 59824 12586 59858 12602
rect 59824 11794 59858 11810
rect 60282 12586 60316 12602
rect 60282 11794 60316 11810
rect 60412 12586 60446 12602
rect 60412 11794 60446 11810
rect 60870 12586 60904 12602
rect 60870 11794 60904 11810
rect 61000 12586 61034 12602
rect 61000 11794 61034 11810
rect 61458 12586 61492 12602
rect 61458 11794 61492 11810
rect 61588 12586 61622 12602
rect 61588 11794 61622 11810
rect 62046 12586 62080 12602
rect 62046 11794 62080 11810
rect 62176 12586 62210 12602
rect 62176 11794 62210 11810
rect 62634 12586 62668 12602
rect 62634 11794 62668 11810
rect 62764 12586 62798 12602
rect 62764 11794 62798 11810
rect 63222 12586 63256 12602
rect 63222 11794 63256 11810
rect 63352 12586 63386 12602
rect 63352 11794 63386 11810
rect 63810 12586 63844 12602
rect 63810 11794 63844 11810
rect 63940 12586 63974 12602
rect 63940 11794 63974 11810
rect 64398 12586 64432 12602
rect 64398 11794 64432 11810
rect 64528 12586 64562 12602
rect 64528 11794 64562 11810
rect 64986 12586 65020 12602
rect 64986 11794 65020 11810
rect 65116 12586 65150 12602
rect 65116 11794 65150 11810
rect 65574 12586 65608 12602
rect 65574 11794 65608 11810
rect 65704 12586 65738 12602
rect 65704 11794 65738 11810
rect 66162 12586 66196 12602
rect 66162 11794 66196 11810
rect 66292 12586 66326 12602
rect 66292 11794 66326 11810
rect 66750 12586 66784 12602
rect 66750 11794 66784 11810
rect 66880 12586 66914 12602
rect 66880 11794 66914 11810
rect 67338 12586 67372 12602
rect 67338 11794 67372 11810
rect 67468 12586 67502 12602
rect 67468 11794 67502 11810
rect 67926 12586 67960 12602
rect 67926 11794 67960 11810
rect 68056 12586 68090 12602
rect 68056 11794 68090 11810
rect 68514 12586 68548 12602
rect 68514 11794 68548 11810
rect 68644 12586 68678 12602
rect 68644 11794 68678 11810
rect 69102 12586 69136 12602
rect 69102 11794 69136 11810
rect 69232 12586 69266 12602
rect 69232 11794 69266 11810
rect 69690 12586 69724 12602
rect 69690 11794 69724 11810
rect 69820 12586 69854 12602
rect 69820 11794 69854 11810
rect 70278 12586 70312 12602
rect 70278 11794 70312 11810
rect 70408 12586 70442 12602
rect 70408 11794 70442 11810
rect 70866 12586 70900 12602
rect 70866 11794 70900 11810
rect 70996 12586 71030 12602
rect 70996 11794 71030 11810
rect 71454 12586 71488 12602
rect 71454 11794 71488 11810
rect 43406 11751 55166 11752
rect 55566 11751 55754 11752
rect 56154 11751 56342 11752
rect 56742 11751 56930 11752
rect 57330 11751 57518 11752
rect 57918 11751 58106 11752
rect 58506 11751 58694 11752
rect 59094 11751 59282 11752
rect 59682 11751 71442 11752
rect 43406 11717 43422 11751
rect 43790 11717 44010 11751
rect 44378 11717 44598 11751
rect 44966 11717 45186 11751
rect 45554 11717 45774 11751
rect 46142 11717 46362 11751
rect 46730 11717 46950 11751
rect 47318 11717 47538 11751
rect 47906 11717 48126 11751
rect 48494 11717 48714 11751
rect 49082 11717 49302 11751
rect 49670 11717 49890 11751
rect 50258 11717 50478 11751
rect 50846 11717 51066 11751
rect 51434 11717 51654 11751
rect 52022 11717 52242 11751
rect 52610 11717 52830 11751
rect 53198 11717 53418 11751
rect 53786 11717 54006 11751
rect 54374 11717 54594 11751
rect 54962 11717 55182 11751
rect 55550 11717 55770 11751
rect 56138 11717 56358 11751
rect 56726 11717 56946 11751
rect 57314 11717 57534 11751
rect 57902 11717 58122 11751
rect 58490 11717 58710 11751
rect 59078 11717 59298 11751
rect 59666 11717 59886 11751
rect 60254 11717 60474 11751
rect 60842 11717 61062 11751
rect 61430 11717 61650 11751
rect 62018 11717 62238 11751
rect 62606 11717 62826 11751
rect 63194 11717 63414 11751
rect 63782 11717 64002 11751
rect 64370 11717 64590 11751
rect 64958 11717 65178 11751
rect 65546 11717 65766 11751
rect 66134 11717 66354 11751
rect 66722 11717 66942 11751
rect 67310 11717 67530 11751
rect 67898 11717 68118 11751
rect 68486 11717 68706 11751
rect 69074 11717 69294 11751
rect 69662 11717 69882 11751
rect 70250 11717 70470 11751
rect 70838 11717 71058 11751
rect 71426 11717 71442 11751
rect 43406 11679 55166 11717
rect 55566 11679 55754 11717
rect 56154 11716 56342 11717
rect 56154 11679 56342 11680
rect 56742 11679 56930 11717
rect 57330 11679 57518 11717
rect 57918 11679 58106 11717
rect 58506 11716 58694 11717
rect 58506 11679 58694 11680
rect 59094 11679 59282 11717
rect 59682 11679 71442 11717
rect 43406 11645 43422 11679
rect 43790 11645 44010 11679
rect 44378 11645 44598 11679
rect 44966 11645 45186 11679
rect 45554 11645 45774 11679
rect 46142 11645 46362 11679
rect 46730 11645 46950 11679
rect 47318 11645 47538 11679
rect 47906 11645 48126 11679
rect 48494 11645 48714 11679
rect 49082 11645 49302 11679
rect 49670 11645 49890 11679
rect 50258 11645 50478 11679
rect 50846 11645 51066 11679
rect 51434 11645 51654 11679
rect 52022 11645 52242 11679
rect 52610 11645 52830 11679
rect 53198 11645 53418 11679
rect 53786 11645 54006 11679
rect 54374 11645 54594 11679
rect 54962 11645 55182 11679
rect 55550 11645 55770 11679
rect 56138 11645 56358 11679
rect 56726 11645 56946 11679
rect 57314 11645 57534 11679
rect 57902 11645 58122 11679
rect 58490 11645 58710 11679
rect 59078 11645 59298 11679
rect 59666 11645 59886 11679
rect 60254 11645 60474 11679
rect 60842 11645 61062 11679
rect 61430 11645 61650 11679
rect 62018 11645 62238 11679
rect 62606 11645 62826 11679
rect 63194 11645 63414 11679
rect 63782 11645 64002 11679
rect 64370 11645 64590 11679
rect 64958 11645 65178 11679
rect 65546 11645 65766 11679
rect 66134 11645 66354 11679
rect 66722 11645 66942 11679
rect 67310 11645 67530 11679
rect 67898 11645 68118 11679
rect 68486 11645 68706 11679
rect 69074 11645 69294 11679
rect 69662 11645 69882 11679
rect 70250 11645 70470 11679
rect 70838 11645 71058 11679
rect 71426 11645 71442 11679
rect 43406 11644 55166 11645
rect 55566 11644 55754 11645
rect 56154 11644 56342 11645
rect 56742 11644 56930 11645
rect 57330 11644 57518 11645
rect 57918 11644 58106 11645
rect 58506 11644 58694 11645
rect 59094 11644 59282 11645
rect 59682 11644 71442 11645
rect 43360 11586 43394 11602
rect 43360 10794 43394 10810
rect 43818 11586 43852 11602
rect 43818 10794 43852 10810
rect 43948 11586 43982 11602
rect 43948 10794 43982 10810
rect 44406 11586 44440 11602
rect 44406 10794 44440 10810
rect 44536 11586 44570 11602
rect 44536 10794 44570 10810
rect 44994 11586 45028 11602
rect 44994 10794 45028 10810
rect 45124 11586 45158 11602
rect 45124 10794 45158 10810
rect 45582 11586 45616 11602
rect 45582 10794 45616 10810
rect 45712 11586 45746 11602
rect 45712 10794 45746 10810
rect 46170 11586 46204 11602
rect 46170 10794 46204 10810
rect 46300 11586 46334 11602
rect 46300 10794 46334 10810
rect 46758 11586 46792 11602
rect 46758 10794 46792 10810
rect 46888 11586 46922 11602
rect 46888 10794 46922 10810
rect 47346 11586 47380 11602
rect 47346 10794 47380 10810
rect 47476 11586 47510 11602
rect 47476 10794 47510 10810
rect 47934 11586 47968 11602
rect 47934 10794 47968 10810
rect 48064 11586 48098 11602
rect 48064 10794 48098 10810
rect 48522 11586 48556 11602
rect 48522 10794 48556 10810
rect 48652 11586 48686 11602
rect 48652 10794 48686 10810
rect 49110 11586 49144 11602
rect 49110 10794 49144 10810
rect 49240 11586 49274 11602
rect 49240 10794 49274 10810
rect 49698 11586 49732 11602
rect 49698 10794 49732 10810
rect 49828 11586 49862 11602
rect 49828 10794 49862 10810
rect 50286 11586 50320 11602
rect 50286 10794 50320 10810
rect 50416 11586 50450 11602
rect 50416 10794 50450 10810
rect 50874 11586 50908 11602
rect 50874 10794 50908 10810
rect 51004 11586 51038 11602
rect 51004 10794 51038 10810
rect 51462 11586 51496 11602
rect 51462 10794 51496 10810
rect 51592 11586 51626 11602
rect 51592 10794 51626 10810
rect 52050 11586 52084 11602
rect 52050 10794 52084 10810
rect 52180 11586 52214 11602
rect 52180 10794 52214 10810
rect 52638 11586 52672 11602
rect 52638 10794 52672 10810
rect 52768 11586 52802 11602
rect 52768 10794 52802 10810
rect 53226 11586 53260 11602
rect 53226 10794 53260 10810
rect 53356 11586 53390 11602
rect 53356 10794 53390 10810
rect 53814 11586 53848 11602
rect 53814 10794 53848 10810
rect 53944 11586 53978 11602
rect 53944 10794 53978 10810
rect 54402 11586 54436 11602
rect 54402 10794 54436 10810
rect 54532 11586 54566 11602
rect 54532 10794 54566 10810
rect 54990 11586 55024 11602
rect 54990 10794 55024 10810
rect 55120 11586 55154 11644
rect 55120 10752 55154 10810
rect 55578 11586 55612 11602
rect 55578 10794 55612 10810
rect 55708 11586 55742 11602
rect 55708 10794 55742 10810
rect 56166 11586 56200 11602
rect 56166 10794 56200 10810
rect 56296 11586 56330 11602
rect 56296 10794 56330 10810
rect 56754 11586 56788 11602
rect 56754 10794 56788 10810
rect 56884 11586 56918 11602
rect 56884 10794 56918 10810
rect 57342 11586 57506 11644
rect 57376 10810 57472 11586
rect 57342 10752 57506 10810
rect 57930 11586 57964 11602
rect 57930 10794 57964 10810
rect 58060 11586 58094 11602
rect 58060 10794 58094 10810
rect 58518 11586 58552 11602
rect 58518 10794 58552 10810
rect 58648 11586 58682 11602
rect 58648 10794 58682 10810
rect 59106 11586 59140 11602
rect 59106 10794 59140 10810
rect 59236 11586 59270 11602
rect 59236 10794 59270 10810
rect 59694 11586 59728 11644
rect 59694 10752 59728 10810
rect 59824 11586 59858 11602
rect 59824 10794 59858 10810
rect 60282 11586 60316 11602
rect 60282 10794 60316 10810
rect 60412 11586 60446 11602
rect 60412 10794 60446 10810
rect 60870 11586 60904 11602
rect 60870 10794 60904 10810
rect 61000 11586 61034 11602
rect 61000 10794 61034 10810
rect 61458 11586 61492 11602
rect 61458 10794 61492 10810
rect 61588 11586 61622 11602
rect 61588 10794 61622 10810
rect 62046 11586 62080 11602
rect 62046 10794 62080 10810
rect 62176 11586 62210 11602
rect 62176 10794 62210 10810
rect 62634 11586 62668 11602
rect 62634 10794 62668 10810
rect 62764 11586 62798 11602
rect 62764 10794 62798 10810
rect 63222 11586 63256 11602
rect 63222 10794 63256 10810
rect 63352 11586 63386 11602
rect 63352 10794 63386 10810
rect 63810 11586 63844 11602
rect 63810 10794 63844 10810
rect 63940 11586 63974 11602
rect 63940 10794 63974 10810
rect 64398 11586 64432 11602
rect 64398 10794 64432 10810
rect 64528 11586 64562 11602
rect 64528 10794 64562 10810
rect 64986 11586 65020 11602
rect 64986 10794 65020 10810
rect 65116 11586 65150 11602
rect 65116 10794 65150 10810
rect 65574 11586 65608 11602
rect 65574 10794 65608 10810
rect 65704 11586 65738 11602
rect 65704 10794 65738 10810
rect 66162 11586 66196 11602
rect 66162 10794 66196 10810
rect 66292 11586 66326 11602
rect 66292 10794 66326 10810
rect 66750 11586 66784 11602
rect 66750 10794 66784 10810
rect 66880 11586 66914 11602
rect 66880 10794 66914 10810
rect 67338 11586 67372 11602
rect 67338 10794 67372 10810
rect 67468 11586 67502 11602
rect 67468 10794 67502 10810
rect 67926 11586 67960 11602
rect 67926 10794 67960 10810
rect 68056 11586 68090 11602
rect 68056 10794 68090 10810
rect 68514 11586 68548 11602
rect 68514 10794 68548 10810
rect 68644 11586 68678 11602
rect 68644 10794 68678 10810
rect 69102 11586 69136 11602
rect 69102 10794 69136 10810
rect 69232 11586 69266 11602
rect 69232 10794 69266 10810
rect 69690 11586 69724 11602
rect 69690 10794 69724 10810
rect 69820 11586 69854 11602
rect 69820 10794 69854 10810
rect 70278 11586 70312 11602
rect 70278 10794 70312 10810
rect 70408 11586 70442 11602
rect 70408 10794 70442 10810
rect 70866 11586 70900 11602
rect 70866 10794 70900 10810
rect 70996 11586 71030 11602
rect 70996 10794 71030 10810
rect 71454 11586 71488 11602
rect 71454 10794 71488 10810
rect 43406 10751 55166 10752
rect 55566 10751 55754 10752
rect 56154 10751 56342 10752
rect 56742 10751 56930 10752
rect 57330 10751 57518 10752
rect 57918 10751 58106 10752
rect 58506 10751 58694 10752
rect 59094 10751 59282 10752
rect 59682 10751 71442 10752
rect 43406 10717 43422 10751
rect 43790 10717 44010 10751
rect 44378 10717 44598 10751
rect 44966 10717 45186 10751
rect 45554 10717 45774 10751
rect 46142 10717 46362 10751
rect 46730 10717 46950 10751
rect 47318 10717 47538 10751
rect 47906 10717 48126 10751
rect 48494 10717 48714 10751
rect 49082 10717 49302 10751
rect 49670 10717 49890 10751
rect 50258 10717 50478 10751
rect 50846 10717 51066 10751
rect 51434 10717 51654 10751
rect 52022 10717 52242 10751
rect 52610 10717 52830 10751
rect 53198 10717 53418 10751
rect 53786 10717 54006 10751
rect 54374 10717 54594 10751
rect 54962 10717 55182 10751
rect 55550 10717 55770 10751
rect 56138 10717 56358 10751
rect 56726 10717 56946 10751
rect 57314 10717 57534 10751
rect 57902 10717 58122 10751
rect 58490 10717 58710 10751
rect 59078 10717 59298 10751
rect 59666 10717 59886 10751
rect 60254 10717 60474 10751
rect 60842 10717 61062 10751
rect 61430 10717 61650 10751
rect 62018 10717 62238 10751
rect 62606 10717 62826 10751
rect 63194 10717 63414 10751
rect 63782 10717 64002 10751
rect 64370 10717 64590 10751
rect 64958 10717 65178 10751
rect 65546 10717 65766 10751
rect 66134 10717 66354 10751
rect 66722 10717 66942 10751
rect 67310 10717 67530 10751
rect 67898 10717 68118 10751
rect 68486 10717 68706 10751
rect 69074 10717 69294 10751
rect 69662 10717 69882 10751
rect 70250 10717 70470 10751
rect 70838 10717 71058 10751
rect 71426 10717 71442 10751
rect 43406 10679 55166 10717
rect 55566 10679 55754 10717
rect 56154 10716 56342 10717
rect 56154 10679 56342 10680
rect 56742 10679 56930 10717
rect 57330 10679 57518 10717
rect 57918 10679 58106 10717
rect 58506 10716 58694 10717
rect 58506 10679 58694 10680
rect 59094 10679 59282 10717
rect 59682 10679 71442 10717
rect 43406 10645 43422 10679
rect 43790 10645 44010 10679
rect 44378 10645 44598 10679
rect 44966 10645 45186 10679
rect 45554 10645 45774 10679
rect 46142 10645 46362 10679
rect 46730 10645 46950 10679
rect 47318 10645 47538 10679
rect 47906 10645 48126 10679
rect 48494 10645 48714 10679
rect 49082 10645 49302 10679
rect 49670 10645 49890 10679
rect 50258 10645 50478 10679
rect 50846 10645 51066 10679
rect 51434 10645 51654 10679
rect 52022 10645 52242 10679
rect 52610 10645 52830 10679
rect 53198 10645 53418 10679
rect 53786 10645 54006 10679
rect 54374 10645 54594 10679
rect 54962 10645 55182 10679
rect 55550 10645 55770 10679
rect 56138 10645 56358 10679
rect 56726 10645 56946 10679
rect 57314 10645 57534 10679
rect 57902 10645 58122 10679
rect 58490 10645 58710 10679
rect 59078 10645 59298 10679
rect 59666 10645 59886 10679
rect 60254 10645 60474 10679
rect 60842 10645 61062 10679
rect 61430 10645 61650 10679
rect 62018 10645 62238 10679
rect 62606 10645 62826 10679
rect 63194 10645 63414 10679
rect 63782 10645 64002 10679
rect 64370 10645 64590 10679
rect 64958 10645 65178 10679
rect 65546 10645 65766 10679
rect 66134 10645 66354 10679
rect 66722 10645 66942 10679
rect 67310 10645 67530 10679
rect 67898 10645 68118 10679
rect 68486 10645 68706 10679
rect 69074 10645 69294 10679
rect 69662 10645 69882 10679
rect 70250 10645 70470 10679
rect 70838 10645 71058 10679
rect 71426 10645 71442 10679
rect 43406 10644 55166 10645
rect 55566 10644 55754 10645
rect 56154 10644 56342 10645
rect 56742 10644 56930 10645
rect 57330 10644 57518 10645
rect 57918 10644 58106 10645
rect 58506 10644 58694 10645
rect 59094 10644 59282 10645
rect 59682 10644 71442 10645
rect 43360 10586 43394 10602
rect 43360 9794 43394 9810
rect 43818 10586 43852 10602
rect 43818 9794 43852 9810
rect 43948 10586 43982 10602
rect 43948 9794 43982 9810
rect 44406 10586 44440 10602
rect 44406 9794 44440 9810
rect 44536 10586 44570 10602
rect 44536 9794 44570 9810
rect 44994 10586 45028 10602
rect 44994 9794 45028 9810
rect 45124 10586 45158 10602
rect 45124 9794 45158 9810
rect 45582 10586 45616 10602
rect 45582 9794 45616 9810
rect 45712 10586 45746 10602
rect 45712 9794 45746 9810
rect 46170 10586 46204 10602
rect 46170 9794 46204 9810
rect 46300 10586 46334 10602
rect 46300 9794 46334 9810
rect 46758 10586 46792 10602
rect 46758 9794 46792 9810
rect 46888 10586 46922 10602
rect 46888 9794 46922 9810
rect 47346 10586 47380 10602
rect 47346 9794 47380 9810
rect 47476 10586 47510 10602
rect 47476 9794 47510 9810
rect 47934 10586 47968 10602
rect 47934 9794 47968 9810
rect 48064 10586 48098 10602
rect 48064 9794 48098 9810
rect 48522 10586 48556 10602
rect 48522 9794 48556 9810
rect 48652 10586 48686 10602
rect 48652 9794 48686 9810
rect 49110 10586 49144 10602
rect 49110 9794 49144 9810
rect 49240 10586 49274 10602
rect 49240 9794 49274 9810
rect 49698 10586 49732 10602
rect 49698 9794 49732 9810
rect 49828 10586 49862 10602
rect 49828 9794 49862 9810
rect 50286 10586 50320 10602
rect 50286 9794 50320 9810
rect 50416 10586 50450 10602
rect 50416 9794 50450 9810
rect 50874 10586 50908 10602
rect 50874 9794 50908 9810
rect 51004 10586 51038 10602
rect 51004 9794 51038 9810
rect 51462 10586 51496 10602
rect 51462 9794 51496 9810
rect 51592 10586 51626 10602
rect 51592 9794 51626 9810
rect 52050 10586 52084 10602
rect 52050 9794 52084 9810
rect 52180 10586 52214 10602
rect 52180 9794 52214 9810
rect 52638 10586 52672 10602
rect 52638 9794 52672 9810
rect 52768 10586 52802 10602
rect 52768 9794 52802 9810
rect 53226 10586 53260 10602
rect 53226 9794 53260 9810
rect 53356 10586 53390 10602
rect 53356 9794 53390 9810
rect 53814 10586 53848 10602
rect 53814 9794 53848 9810
rect 53944 10586 53978 10602
rect 53944 9794 53978 9810
rect 54402 10586 54436 10602
rect 54402 9794 54436 9810
rect 54532 10586 54566 10602
rect 54532 9794 54566 9810
rect 54990 10586 55024 10602
rect 54990 9794 55024 9810
rect 55120 10586 55154 10644
rect 55120 9794 55154 9810
rect 55578 10586 55612 10602
rect 55578 9794 55612 9810
rect 55708 10586 55742 10602
rect 55708 9794 55742 9810
rect 56166 10586 56200 10602
rect 56166 9794 56200 9810
rect 56296 10586 56330 10602
rect 56296 9794 56330 9810
rect 56754 10586 56788 10602
rect 56754 9794 56788 9810
rect 56884 10586 56918 10602
rect 56884 9794 56918 9810
rect 57342 10586 57506 10644
rect 57376 9810 57472 10586
rect 57342 9794 57506 9810
rect 57930 10586 57964 10602
rect 57930 9794 57964 9810
rect 58060 10586 58094 10602
rect 58060 9794 58094 9810
rect 58518 10586 58552 10602
rect 58518 9794 58552 9810
rect 58648 10586 58682 10602
rect 58648 9794 58682 9810
rect 59106 10586 59140 10602
rect 59106 9794 59140 9810
rect 59236 10586 59270 10602
rect 59236 9794 59270 9810
rect 59694 10586 59728 10644
rect 59694 9794 59728 9810
rect 59824 10586 59858 10602
rect 59824 9794 59858 9810
rect 60282 10586 60316 10602
rect 60282 9794 60316 9810
rect 60412 10586 60446 10602
rect 60412 9794 60446 9810
rect 60870 10586 60904 10602
rect 60870 9794 60904 9810
rect 61000 10586 61034 10602
rect 61000 9794 61034 9810
rect 61458 10586 61492 10602
rect 61458 9794 61492 9810
rect 61588 10586 61622 10602
rect 61588 9794 61622 9810
rect 62046 10586 62080 10602
rect 62046 9794 62080 9810
rect 62176 10586 62210 10602
rect 62176 9794 62210 9810
rect 62634 10586 62668 10602
rect 62634 9794 62668 9810
rect 62764 10586 62798 10602
rect 62764 9794 62798 9810
rect 63222 10586 63256 10602
rect 63222 9794 63256 9810
rect 63352 10586 63386 10602
rect 63352 9794 63386 9810
rect 63810 10586 63844 10602
rect 63810 9794 63844 9810
rect 63940 10586 63974 10602
rect 63940 9794 63974 9810
rect 64398 10586 64432 10602
rect 64398 9794 64432 9810
rect 64528 10586 64562 10602
rect 64528 9794 64562 9810
rect 64986 10586 65020 10602
rect 64986 9794 65020 9810
rect 65116 10586 65150 10602
rect 65116 9794 65150 9810
rect 65574 10586 65608 10602
rect 65574 9794 65608 9810
rect 65704 10586 65738 10602
rect 65704 9794 65738 9810
rect 66162 10586 66196 10602
rect 66162 9794 66196 9810
rect 66292 10586 66326 10602
rect 66292 9794 66326 9810
rect 66750 10586 66784 10602
rect 66750 9794 66784 9810
rect 66880 10586 66914 10602
rect 66880 9794 66914 9810
rect 67338 10586 67372 10602
rect 67338 9794 67372 9810
rect 67468 10586 67502 10602
rect 67468 9794 67502 9810
rect 67926 10586 67960 10602
rect 67926 9794 67960 9810
rect 68056 10586 68090 10602
rect 68056 9794 68090 9810
rect 68514 10586 68548 10602
rect 68514 9794 68548 9810
rect 68644 10586 68678 10602
rect 68644 9794 68678 9810
rect 69102 10586 69136 10602
rect 69102 9794 69136 9810
rect 69232 10586 69266 10602
rect 69232 9794 69266 9810
rect 69690 10586 69724 10602
rect 69690 9794 69724 9810
rect 69820 10586 69854 10602
rect 69820 9794 69854 9810
rect 70278 10586 70312 10602
rect 70278 9794 70312 9810
rect 70408 10586 70442 10602
rect 70408 9794 70442 9810
rect 70866 10586 70900 10602
rect 70866 9794 70900 9810
rect 70996 10586 71030 10602
rect 70996 9794 71030 9810
rect 71454 10586 71488 10602
rect 71454 9794 71488 9810
rect 55120 9752 55166 9794
rect 43406 9751 55166 9752
rect 55566 9751 55754 9752
rect 56154 9751 56342 9752
rect 56742 9751 56930 9752
rect 57330 9751 57518 9794
rect 59682 9752 59728 9794
rect 57918 9751 58106 9752
rect 58506 9751 58694 9752
rect 59094 9751 59282 9752
rect 59682 9751 71442 9752
rect 43406 9717 43422 9751
rect 43790 9717 44010 9751
rect 44378 9717 44598 9751
rect 44966 9717 45186 9751
rect 45554 9717 45774 9751
rect 46142 9717 46362 9751
rect 46730 9717 46950 9751
rect 47318 9717 47538 9751
rect 47906 9717 48126 9751
rect 48494 9717 48714 9751
rect 49082 9717 49302 9751
rect 49670 9717 49890 9751
rect 50258 9717 50478 9751
rect 50846 9717 51066 9751
rect 51434 9717 51654 9751
rect 52022 9717 52242 9751
rect 52610 9717 52830 9751
rect 53198 9717 53418 9751
rect 53786 9717 54006 9751
rect 54374 9717 54594 9751
rect 54962 9717 55182 9751
rect 55550 9717 55770 9751
rect 56138 9717 56358 9751
rect 56726 9717 56946 9751
rect 57314 9717 57534 9751
rect 57902 9717 58122 9751
rect 58490 9717 58710 9751
rect 59078 9717 59298 9751
rect 59666 9717 59886 9751
rect 60254 9717 60474 9751
rect 60842 9717 61062 9751
rect 61430 9717 61650 9751
rect 62018 9717 62238 9751
rect 62606 9717 62826 9751
rect 63194 9717 63414 9751
rect 63782 9717 64002 9751
rect 64370 9717 64590 9751
rect 64958 9717 65178 9751
rect 65546 9717 65766 9751
rect 66134 9717 66354 9751
rect 66722 9717 66942 9751
rect 67310 9717 67530 9751
rect 67898 9717 68118 9751
rect 68486 9717 68706 9751
rect 69074 9717 69294 9751
rect 69662 9717 69882 9751
rect 70250 9717 70470 9751
rect 70838 9717 71058 9751
rect 71426 9717 71442 9751
rect 43406 9716 55166 9717
rect 55566 9716 55754 9717
rect 56154 9716 56342 9717
rect 56742 9716 56930 9717
rect 57330 9716 57518 9717
rect 57918 9716 58106 9717
rect 58506 9716 58694 9717
rect 59094 9716 59282 9717
rect 59682 9716 71442 9717
rect 43014 9400 43048 9420
rect 71800 9400 71834 9454
rect 43014 9366 43132 9400
rect 71746 9366 71834 9400
rect 56716 9338 56742 9366
rect 56930 9338 56960 9366
rect 56716 8656 56960 9338
rect 57890 9338 57918 9366
rect 58106 9338 58134 9366
rect 57890 8656 58134 9338
rect 56026 8622 56060 8656
rect 58788 8622 58822 8656
rect 56458 8190 56474 8322
rect 56512 8190 56740 8322
rect 56778 8190 56796 8322
rect 56990 8190 57006 8322
rect 57044 8190 57272 8322
rect 57310 8190 57328 8322
rect 57522 8190 57538 8322
rect 57576 8190 57804 8322
rect 57842 8190 57860 8322
rect 58054 8190 58070 8322
rect 58108 8190 58336 8322
rect 58374 8190 58392 8322
rect 56412 8140 56446 8156
rect 56412 7348 56446 7364
rect 56540 8140 56574 8156
rect 56540 7348 56574 7364
rect 56678 8140 56712 8156
rect 56678 7348 56712 7364
rect 56806 8140 56840 8156
rect 56806 7348 56840 7364
rect 56944 8140 56978 8156
rect 56944 7348 56978 7364
rect 57072 8140 57106 8156
rect 57072 7348 57106 7364
rect 57210 8140 57244 8156
rect 57210 7348 57244 7364
rect 57338 8140 57372 8156
rect 57338 7348 57372 7364
rect 57476 8140 57510 8156
rect 57476 7348 57510 7364
rect 57604 8140 57638 8156
rect 57604 7348 57638 7364
rect 57742 8140 57776 8156
rect 57742 7348 57776 7364
rect 57870 8140 57904 8156
rect 57870 7348 57904 7364
rect 58008 8140 58042 8156
rect 58008 7348 58042 7364
rect 58136 8140 58170 8156
rect 58136 7348 58170 7364
rect 58274 8140 58308 8156
rect 58274 7348 58308 7364
rect 58402 8140 58436 8156
rect 58402 7348 58436 7364
rect 56458 7180 56474 7312
rect 56512 7180 56740 7312
rect 56778 7180 56796 7312
rect 56990 7180 57006 7312
rect 57044 7180 57272 7312
rect 57310 7180 57328 7312
rect 57522 7180 57538 7312
rect 57576 7180 57804 7312
rect 57842 7180 57860 7312
rect 58054 7180 58070 7312
rect 58108 7180 58336 7312
rect 58374 7180 58392 7312
rect 56412 7130 56446 7146
rect 56412 6338 56446 6354
rect 56540 7130 56574 7146
rect 56540 6338 56574 6354
rect 56678 7130 56712 7146
rect 56678 6338 56712 6354
rect 56806 7130 56840 7146
rect 56806 6338 56840 6354
rect 56944 7130 56978 7146
rect 56944 6338 56978 6354
rect 57072 7130 57106 7146
rect 57072 6338 57106 6354
rect 57210 7130 57244 7146
rect 57210 6338 57244 6354
rect 57338 7130 57372 7146
rect 57338 6338 57372 6354
rect 57476 7130 57510 7146
rect 57476 6338 57510 6354
rect 57604 7130 57638 7146
rect 57604 6338 57638 6354
rect 57742 7130 57776 7146
rect 57742 6338 57776 6354
rect 57870 7130 57904 7146
rect 57870 6338 57904 6354
rect 58008 7130 58042 7146
rect 58008 6338 58042 6354
rect 58136 7130 58170 7146
rect 58136 6338 58170 6354
rect 58274 7130 58308 7146
rect 58274 6338 58308 6354
rect 58402 7130 58436 7146
rect 58402 6338 58436 6354
rect 56458 6170 56474 6302
rect 56512 6170 56740 6302
rect 56778 6170 56796 6302
rect 56990 6170 57006 6302
rect 57044 6170 57272 6302
rect 57310 6170 57328 6302
rect 57522 6170 57538 6302
rect 57576 6170 57804 6302
rect 57842 6170 57860 6302
rect 58054 6170 58070 6302
rect 58108 6170 58336 6302
rect 58374 6170 58392 6302
rect 56412 6120 56446 6136
rect 56412 5328 56446 5344
rect 56540 6120 56574 6136
rect 56540 5328 56574 5344
rect 56678 6120 56712 6136
rect 56678 5328 56712 5344
rect 56806 6120 56840 6136
rect 56806 5328 56840 5344
rect 56944 6120 56978 6136
rect 56944 5328 56978 5344
rect 57072 6120 57106 6136
rect 57072 5328 57106 5344
rect 57210 6120 57244 6136
rect 57210 5328 57244 5344
rect 57338 6120 57372 6136
rect 57338 5328 57372 5344
rect 57476 6120 57510 6136
rect 57476 5328 57510 5344
rect 57604 6120 57638 6136
rect 57604 5328 57638 5344
rect 57742 6120 57776 6136
rect 57742 5328 57776 5344
rect 57870 6120 57904 6136
rect 57870 5328 57904 5344
rect 58008 6120 58042 6136
rect 58008 5328 58042 5344
rect 58136 6120 58170 6136
rect 58136 5328 58170 5344
rect 58274 6120 58308 6136
rect 58274 5328 58308 5344
rect 58402 6120 58436 6136
rect 58402 5328 58436 5344
rect 56458 5160 56474 5292
rect 56512 5160 56740 5292
rect 56778 5160 56796 5292
rect 56990 5160 57006 5292
rect 57044 5160 57272 5292
rect 57310 5160 57328 5292
rect 57522 5160 57538 5292
rect 57576 5160 57804 5292
rect 57842 5160 57860 5292
rect 58054 5160 58070 5292
rect 58108 5160 58336 5292
rect 58374 5160 58392 5292
rect 56026 4826 56060 4860
rect 58788 4826 58822 4860
rect 56638 4430 56784 4464
rect 57994 4430 58212 4464
rect 56984 4124 57866 4130
rect 56984 3998 57046 4124
rect 57084 3998 57286 4124
rect 57324 3998 57526 4124
rect 57564 3998 57766 4124
rect 57804 3998 57866 4124
rect 56984 3948 57018 3998
rect 56984 3322 57018 3372
rect 57112 3948 57146 3964
rect 57112 3356 57146 3372
rect 57224 3948 57258 3964
rect 57224 3356 57258 3372
rect 57352 3948 57386 3964
rect 57352 3356 57386 3372
rect 57464 3948 57498 3964
rect 57464 3356 57498 3372
rect 57592 3948 57626 3964
rect 57592 3356 57626 3372
rect 57704 3948 57738 3964
rect 57704 3356 57738 3372
rect 57832 3948 57866 3998
rect 57832 3322 57866 3372
rect 56984 3190 57046 3322
rect 57084 3190 57286 3322
rect 57324 3190 57526 3322
rect 57564 3190 57766 3322
rect 57804 3190 57866 3322
rect 56984 3140 57018 3190
rect 56984 2514 57018 2564
rect 57112 3140 57146 3156
rect 57112 2548 57146 2564
rect 57224 3140 57258 3156
rect 57224 2548 57258 2564
rect 57352 3140 57386 3156
rect 57352 2548 57386 2564
rect 57464 3140 57498 3156
rect 57464 2548 57498 2564
rect 57592 3140 57626 3156
rect 57592 2548 57626 2564
rect 57704 3140 57738 3156
rect 57704 2548 57738 2564
rect 57832 3140 57866 3190
rect 57832 2514 57866 2564
rect 56984 2382 57046 2514
rect 57084 2382 57286 2514
rect 57324 2382 57526 2514
rect 57564 2382 57766 2514
rect 57804 2382 57866 2514
rect 56638 2048 56736 2082
rect 58088 2048 58212 2082
<< viali >>
rect 52810 17152 52920 17186
rect 53290 17152 53400 17186
rect 53770 17152 53880 17186
rect 54250 17152 54360 17186
rect 54730 17152 54840 17186
rect 55210 17152 55320 17186
rect 55690 17152 55800 17186
rect 56170 17152 56280 17186
rect 56650 17152 56760 17186
rect 57130 17152 57240 17186
rect 57610 17152 57720 17186
rect 58090 17152 58200 17186
rect 58570 17152 58680 17186
rect 59050 17152 59160 17186
rect 59530 17152 59640 17186
rect 60010 17152 60120 17186
rect 60490 17152 60600 17186
rect 60970 17152 61080 17186
rect 61450 17152 61560 17186
rect 61930 17152 62040 17186
rect 52810 17114 52920 17152
rect 53290 17114 53400 17152
rect 53770 17114 53880 17152
rect 54250 17114 54360 17152
rect 54730 17114 54840 17152
rect 55210 17114 55320 17152
rect 55690 17114 55800 17152
rect 56170 17114 56280 17152
rect 56650 17114 56760 17152
rect 57130 17114 57240 17152
rect 57610 17114 57720 17152
rect 58090 17114 58200 17152
rect 58570 17114 58680 17152
rect 59050 17114 59160 17152
rect 59530 17114 59640 17152
rect 60010 17114 60120 17152
rect 60490 17114 60600 17152
rect 60970 17114 61080 17152
rect 61450 17114 61560 17152
rect 61930 17114 62040 17152
rect 52726 16710 52764 16842
rect 52966 16710 53004 16842
rect 53206 16710 53244 16842
rect 53446 16710 53484 16842
rect 53686 16710 53724 16842
rect 53926 16710 53964 16842
rect 54166 16710 54204 16842
rect 54406 16710 54444 16842
rect 54646 16710 54684 16842
rect 54886 16710 54924 16842
rect 55126 16710 55164 16842
rect 55366 16710 55404 16842
rect 55606 16710 55644 16842
rect 55846 16710 55884 16842
rect 56086 16710 56124 16842
rect 56326 16710 56364 16842
rect 56566 16710 56604 16842
rect 56806 16710 56844 16842
rect 57046 16710 57084 16842
rect 57286 16710 57324 16842
rect 57526 16710 57564 16842
rect 57766 16710 57804 16842
rect 58006 16710 58044 16842
rect 58246 16710 58284 16842
rect 58486 16710 58524 16842
rect 58726 16710 58764 16842
rect 58966 16710 59004 16842
rect 59206 16710 59244 16842
rect 59446 16710 59484 16842
rect 59686 16710 59724 16842
rect 59926 16710 59964 16842
rect 60166 16710 60204 16842
rect 60406 16710 60444 16842
rect 60646 16710 60684 16842
rect 60886 16710 60924 16842
rect 61126 16710 61164 16842
rect 61366 16710 61404 16842
rect 61606 16710 61644 16842
rect 61846 16710 61884 16842
rect 62086 16710 62124 16842
rect 52664 16084 52698 16660
rect 52792 16084 52826 16660
rect 52904 16084 52938 16660
rect 53032 16084 53066 16660
rect 53144 16084 53178 16660
rect 53272 16084 53306 16660
rect 53384 16084 53418 16660
rect 53512 16084 53546 16660
rect 53624 16084 53658 16660
rect 53752 16084 53786 16660
rect 53864 16084 53898 16660
rect 53992 16084 54026 16660
rect 54104 16084 54138 16660
rect 54232 16084 54266 16660
rect 54344 16084 54378 16660
rect 54472 16084 54506 16660
rect 54584 16084 54618 16660
rect 54712 16084 54746 16660
rect 54824 16084 54858 16660
rect 54952 16084 54986 16660
rect 55064 16084 55098 16660
rect 55192 16084 55226 16660
rect 55304 16084 55338 16660
rect 55432 16084 55466 16660
rect 55544 16084 55578 16660
rect 55672 16084 55706 16660
rect 55784 16084 55818 16660
rect 55912 16084 55946 16660
rect 56024 16084 56058 16660
rect 56152 16084 56186 16660
rect 56264 16084 56298 16660
rect 56392 16084 56426 16660
rect 56504 16084 56538 16660
rect 56632 16084 56666 16660
rect 56744 16084 56778 16660
rect 56872 16084 56906 16660
rect 56984 16084 57018 16660
rect 57112 16084 57146 16660
rect 57224 16084 57258 16660
rect 57352 16084 57386 16660
rect 57464 16084 57498 16660
rect 57592 16084 57626 16660
rect 57704 16084 57738 16660
rect 57832 16084 57866 16660
rect 57944 16084 57978 16660
rect 58072 16084 58106 16660
rect 58184 16084 58218 16660
rect 58312 16084 58346 16660
rect 58424 16084 58458 16660
rect 58552 16084 58586 16660
rect 58664 16084 58698 16660
rect 58792 16084 58826 16660
rect 58904 16084 58938 16660
rect 59032 16084 59066 16660
rect 59144 16084 59178 16660
rect 59272 16084 59306 16660
rect 59384 16084 59418 16660
rect 59512 16084 59546 16660
rect 59624 16084 59658 16660
rect 59752 16084 59786 16660
rect 59864 16084 59898 16660
rect 59992 16084 60026 16660
rect 60104 16084 60138 16660
rect 60232 16084 60266 16660
rect 60344 16084 60378 16660
rect 60472 16084 60506 16660
rect 60584 16084 60618 16660
rect 60712 16084 60746 16660
rect 60824 16084 60858 16660
rect 60952 16084 60986 16660
rect 61064 16084 61098 16660
rect 61192 16084 61226 16660
rect 61304 16084 61338 16660
rect 61432 16084 61466 16660
rect 61544 16084 61578 16660
rect 61672 16084 61706 16660
rect 61784 16084 61818 16660
rect 61912 16084 61946 16660
rect 62024 16084 62058 16660
rect 62152 16084 62186 16660
rect 52726 15902 52764 16034
rect 52966 15902 53004 16034
rect 53206 15902 53244 16034
rect 53446 15902 53484 16034
rect 53686 15902 53724 16034
rect 53926 15902 53964 16034
rect 54166 15902 54204 16034
rect 54406 15902 54444 16034
rect 54646 15902 54684 16034
rect 54886 15902 54924 16034
rect 55126 15902 55164 16034
rect 55366 15902 55404 16034
rect 55606 15902 55644 16034
rect 55846 15902 55884 16034
rect 56086 15902 56124 16034
rect 56326 15902 56364 16034
rect 56566 15902 56604 16034
rect 56806 15902 56844 16034
rect 57046 15902 57084 16034
rect 57286 15902 57324 16034
rect 57526 15902 57564 16034
rect 57766 15902 57804 16034
rect 58006 15902 58044 16034
rect 58246 15902 58284 16034
rect 58486 15902 58524 16034
rect 58726 15902 58764 16034
rect 58966 15902 59004 16034
rect 59206 15902 59244 16034
rect 59446 15902 59484 16034
rect 59686 15902 59724 16034
rect 59926 15902 59964 16034
rect 60166 15902 60204 16034
rect 60406 15902 60444 16034
rect 60646 15902 60684 16034
rect 60886 15902 60924 16034
rect 61126 15902 61164 16034
rect 61366 15902 61404 16034
rect 61606 15902 61644 16034
rect 61846 15902 61884 16034
rect 62086 15902 62124 16034
rect 52664 15276 52698 15852
rect 52792 15276 52826 15852
rect 52904 15276 52938 15852
rect 53032 15276 53066 15852
rect 53144 15276 53178 15852
rect 53272 15276 53306 15852
rect 53384 15276 53418 15852
rect 53512 15276 53546 15852
rect 53624 15276 53658 15852
rect 53752 15276 53786 15852
rect 53864 15276 53898 15852
rect 53992 15276 54026 15852
rect 54104 15276 54138 15852
rect 54232 15276 54266 15852
rect 54344 15276 54378 15852
rect 54472 15276 54506 15852
rect 54584 15276 54618 15852
rect 54712 15276 54746 15852
rect 54824 15276 54858 15852
rect 54952 15276 54986 15852
rect 55064 15276 55098 15852
rect 55192 15276 55226 15852
rect 55304 15276 55338 15852
rect 55432 15276 55466 15852
rect 55544 15276 55578 15852
rect 55672 15276 55706 15852
rect 55784 15276 55818 15852
rect 55912 15276 55946 15852
rect 56024 15276 56058 15852
rect 56152 15276 56186 15852
rect 56264 15276 56298 15852
rect 56392 15276 56426 15852
rect 56504 15276 56538 15852
rect 56632 15276 56666 15852
rect 56744 15276 56778 15852
rect 56872 15276 56906 15852
rect 56984 15276 57018 15852
rect 57112 15276 57146 15852
rect 57224 15276 57258 15852
rect 57352 15276 57386 15852
rect 57464 15276 57498 15852
rect 57592 15276 57626 15852
rect 57704 15276 57738 15852
rect 57832 15276 57866 15852
rect 57944 15276 57978 15852
rect 58072 15276 58106 15852
rect 58184 15276 58218 15852
rect 58312 15276 58346 15852
rect 58424 15276 58458 15852
rect 58552 15276 58586 15852
rect 58664 15276 58698 15852
rect 58792 15276 58826 15852
rect 58904 15276 58938 15852
rect 59032 15276 59066 15852
rect 59144 15276 59178 15852
rect 59272 15276 59306 15852
rect 59384 15276 59418 15852
rect 59512 15276 59546 15852
rect 59624 15276 59658 15852
rect 59752 15276 59786 15852
rect 59864 15276 59898 15852
rect 59992 15276 60026 15852
rect 60104 15276 60138 15852
rect 60232 15276 60266 15852
rect 60344 15276 60378 15852
rect 60472 15276 60506 15852
rect 60584 15276 60618 15852
rect 60712 15276 60746 15852
rect 60824 15276 60858 15852
rect 60952 15276 60986 15852
rect 61064 15276 61098 15852
rect 61192 15276 61226 15852
rect 61304 15276 61338 15852
rect 61432 15276 61466 15852
rect 61544 15276 61578 15852
rect 61672 15276 61706 15852
rect 61784 15276 61818 15852
rect 61912 15276 61946 15852
rect 62024 15276 62058 15852
rect 62152 15276 62186 15852
rect 52726 15094 52764 15226
rect 52966 15094 53004 15226
rect 53206 15094 53244 15226
rect 53446 15094 53484 15226
rect 53686 15094 53724 15226
rect 53926 15094 53964 15226
rect 54166 15094 54204 15226
rect 54406 15094 54444 15226
rect 54646 15094 54684 15226
rect 54886 15094 54924 15226
rect 55126 15094 55164 15226
rect 55366 15094 55404 15226
rect 55606 15094 55644 15226
rect 55846 15094 55884 15226
rect 56086 15094 56124 15226
rect 56326 15094 56364 15226
rect 56566 15094 56604 15226
rect 56806 15094 56844 15226
rect 57046 15094 57084 15226
rect 57286 15094 57324 15226
rect 57526 15094 57564 15226
rect 57766 15094 57804 15226
rect 58006 15094 58044 15226
rect 58246 15094 58284 15226
rect 58486 15094 58524 15226
rect 58726 15094 58764 15226
rect 58966 15094 59004 15226
rect 59206 15094 59244 15226
rect 59446 15094 59484 15226
rect 59686 15094 59724 15226
rect 59926 15094 59964 15226
rect 60166 15094 60204 15226
rect 60406 15094 60444 15226
rect 60646 15094 60684 15226
rect 60886 15094 60924 15226
rect 61126 15094 61164 15226
rect 61366 15094 61404 15226
rect 61606 15094 61644 15226
rect 61846 15094 61884 15226
rect 62086 15094 62124 15226
rect 43422 12645 43790 12679
rect 44010 12645 44378 12679
rect 44598 12645 44966 12679
rect 45186 12645 45554 12679
rect 45774 12645 46142 12679
rect 46362 12645 46730 12679
rect 46950 12645 47318 12679
rect 47538 12645 47906 12679
rect 48126 12645 48494 12679
rect 48714 12645 49082 12679
rect 49302 12645 49670 12679
rect 49890 12645 50258 12679
rect 50478 12645 50846 12679
rect 51066 12645 51434 12679
rect 51654 12645 52022 12679
rect 52242 12645 52610 12679
rect 52830 12645 53198 12679
rect 53418 12645 53786 12679
rect 54006 12645 54374 12679
rect 54594 12645 54962 12679
rect 55182 12645 55550 12679
rect 55770 12645 56138 12679
rect 56358 12645 56726 12679
rect 56946 12645 57314 12679
rect 57534 12645 57902 12679
rect 58122 12645 58490 12679
rect 58710 12645 59078 12679
rect 59298 12645 59666 12679
rect 59886 12645 60254 12679
rect 60474 12645 60842 12679
rect 61062 12645 61430 12679
rect 61650 12645 62018 12679
rect 62238 12645 62606 12679
rect 62826 12645 63194 12679
rect 63414 12645 63782 12679
rect 64002 12645 64370 12679
rect 64590 12645 64958 12679
rect 65178 12645 65546 12679
rect 65766 12645 66134 12679
rect 66354 12645 66722 12679
rect 66942 12645 67310 12679
rect 67530 12645 67898 12679
rect 68118 12645 68486 12679
rect 68706 12645 69074 12679
rect 69294 12645 69662 12679
rect 69882 12645 70250 12679
rect 70470 12645 70838 12679
rect 71058 12645 71426 12679
rect 43360 11810 43394 12586
rect 43818 11810 43852 12586
rect 43948 11810 43982 12586
rect 44406 11810 44440 12586
rect 44536 11810 44570 12586
rect 44994 11810 45028 12586
rect 45124 11810 45158 12586
rect 45582 11810 45616 12586
rect 45712 11810 45746 12586
rect 46170 11810 46204 12586
rect 46300 11810 46334 12586
rect 46758 11810 46792 12586
rect 46888 11810 46922 12586
rect 47346 11810 47380 12586
rect 47476 11810 47510 12586
rect 47934 11810 47968 12586
rect 48064 11810 48098 12586
rect 48522 11810 48556 12586
rect 48652 11810 48686 12586
rect 49110 11810 49144 12586
rect 49240 11810 49274 12586
rect 49698 11810 49732 12586
rect 49828 11810 49862 12586
rect 50286 11810 50320 12586
rect 50416 11810 50450 12586
rect 50874 11810 50908 12586
rect 51004 11810 51038 12586
rect 51462 11810 51496 12586
rect 51592 11810 51626 12586
rect 52050 11810 52084 12586
rect 52180 11810 52214 12586
rect 52638 11810 52672 12586
rect 52768 11810 52802 12586
rect 53226 11810 53260 12586
rect 53356 11810 53390 12586
rect 53814 11810 53848 12586
rect 53944 11810 53978 12586
rect 54402 11810 54436 12586
rect 54532 11810 54566 12586
rect 54990 11810 55024 12586
rect 55120 11810 55154 12586
rect 55578 11810 55612 12586
rect 55708 11810 55742 12586
rect 56166 11810 56200 12586
rect 56296 11810 56330 12586
rect 56754 11810 56788 12586
rect 56884 11810 56918 12586
rect 57342 11810 57376 12586
rect 57472 11810 57506 12586
rect 57930 11810 57964 12586
rect 58060 11810 58094 12586
rect 58518 11810 58552 12586
rect 58648 11810 58682 12586
rect 59106 11810 59140 12586
rect 59236 11810 59270 12586
rect 59694 11810 59728 12586
rect 59824 11810 59858 12586
rect 60282 11810 60316 12586
rect 60412 11810 60446 12586
rect 60870 11810 60904 12586
rect 61000 11810 61034 12586
rect 61458 11810 61492 12586
rect 61588 11810 61622 12586
rect 62046 11810 62080 12586
rect 62176 11810 62210 12586
rect 62634 11810 62668 12586
rect 62764 11810 62798 12586
rect 63222 11810 63256 12586
rect 63352 11810 63386 12586
rect 63810 11810 63844 12586
rect 63940 11810 63974 12586
rect 64398 11810 64432 12586
rect 64528 11810 64562 12586
rect 64986 11810 65020 12586
rect 65116 11810 65150 12586
rect 65574 11810 65608 12586
rect 65704 11810 65738 12586
rect 66162 11810 66196 12586
rect 66292 11810 66326 12586
rect 66750 11810 66784 12586
rect 66880 11810 66914 12586
rect 67338 11810 67372 12586
rect 67468 11810 67502 12586
rect 67926 11810 67960 12586
rect 68056 11810 68090 12586
rect 68514 11810 68548 12586
rect 68644 11810 68678 12586
rect 69102 11810 69136 12586
rect 69232 11810 69266 12586
rect 69690 11810 69724 12586
rect 69820 11810 69854 12586
rect 70278 11810 70312 12586
rect 70408 11810 70442 12586
rect 70866 11810 70900 12586
rect 70996 11810 71030 12586
rect 71454 11810 71488 12586
rect 43422 11717 43790 11751
rect 44010 11717 44378 11751
rect 44598 11717 44966 11751
rect 45186 11717 45554 11751
rect 45774 11717 46142 11751
rect 46362 11717 46730 11751
rect 46950 11717 47318 11751
rect 47538 11717 47906 11751
rect 48126 11717 48494 11751
rect 48714 11717 49082 11751
rect 49302 11717 49670 11751
rect 49890 11717 50258 11751
rect 50478 11717 50846 11751
rect 51066 11717 51434 11751
rect 51654 11717 52022 11751
rect 52242 11717 52610 11751
rect 52830 11717 53198 11751
rect 53418 11717 53786 11751
rect 54006 11717 54374 11751
rect 54594 11717 54962 11751
rect 55182 11717 55550 11751
rect 55770 11717 56138 11751
rect 56358 11717 56726 11751
rect 56946 11717 57314 11751
rect 57534 11717 57902 11751
rect 58122 11717 58490 11751
rect 58710 11717 59078 11751
rect 59298 11717 59666 11751
rect 59886 11717 60254 11751
rect 60474 11717 60842 11751
rect 61062 11717 61430 11751
rect 61650 11717 62018 11751
rect 62238 11717 62606 11751
rect 62826 11717 63194 11751
rect 63414 11717 63782 11751
rect 64002 11717 64370 11751
rect 64590 11717 64958 11751
rect 65178 11717 65546 11751
rect 65766 11717 66134 11751
rect 66354 11717 66722 11751
rect 66942 11717 67310 11751
rect 67530 11717 67898 11751
rect 68118 11717 68486 11751
rect 68706 11717 69074 11751
rect 69294 11717 69662 11751
rect 69882 11717 70250 11751
rect 70470 11717 70838 11751
rect 71058 11717 71426 11751
rect 43422 11645 43790 11679
rect 44010 11645 44378 11679
rect 44598 11645 44966 11679
rect 45186 11645 45554 11679
rect 45774 11645 46142 11679
rect 46362 11645 46730 11679
rect 46950 11645 47318 11679
rect 47538 11645 47906 11679
rect 48126 11645 48494 11679
rect 48714 11645 49082 11679
rect 49302 11645 49670 11679
rect 49890 11645 50258 11679
rect 50478 11645 50846 11679
rect 51066 11645 51434 11679
rect 51654 11645 52022 11679
rect 52242 11645 52610 11679
rect 52830 11645 53198 11679
rect 53418 11645 53786 11679
rect 54006 11645 54374 11679
rect 54594 11645 54962 11679
rect 55182 11645 55550 11679
rect 55770 11645 56138 11679
rect 56358 11645 56726 11679
rect 56946 11645 57314 11679
rect 57534 11645 57902 11679
rect 58122 11645 58490 11679
rect 58710 11645 59078 11679
rect 59298 11645 59666 11679
rect 59886 11645 60254 11679
rect 60474 11645 60842 11679
rect 61062 11645 61430 11679
rect 61650 11645 62018 11679
rect 62238 11645 62606 11679
rect 62826 11645 63194 11679
rect 63414 11645 63782 11679
rect 64002 11645 64370 11679
rect 64590 11645 64958 11679
rect 65178 11645 65546 11679
rect 65766 11645 66134 11679
rect 66354 11645 66722 11679
rect 66942 11645 67310 11679
rect 67530 11645 67898 11679
rect 68118 11645 68486 11679
rect 68706 11645 69074 11679
rect 69294 11645 69662 11679
rect 69882 11645 70250 11679
rect 70470 11645 70838 11679
rect 71058 11645 71426 11679
rect 43360 10810 43394 11586
rect 43818 10810 43852 11586
rect 43948 10810 43982 11586
rect 44406 10810 44440 11586
rect 44536 10810 44570 11586
rect 44994 10810 45028 11586
rect 45124 10810 45158 11586
rect 45582 10810 45616 11586
rect 45712 10810 45746 11586
rect 46170 10810 46204 11586
rect 46300 10810 46334 11586
rect 46758 10810 46792 11586
rect 46888 10810 46922 11586
rect 47346 10810 47380 11586
rect 47476 10810 47510 11586
rect 47934 10810 47968 11586
rect 48064 10810 48098 11586
rect 48522 10810 48556 11586
rect 48652 10810 48686 11586
rect 49110 10810 49144 11586
rect 49240 10810 49274 11586
rect 49698 10810 49732 11586
rect 49828 10810 49862 11586
rect 50286 10810 50320 11586
rect 50416 10810 50450 11586
rect 50874 10810 50908 11586
rect 51004 10810 51038 11586
rect 51462 10810 51496 11586
rect 51592 10810 51626 11586
rect 52050 10810 52084 11586
rect 52180 10810 52214 11586
rect 52638 10810 52672 11586
rect 52768 10810 52802 11586
rect 53226 10810 53260 11586
rect 53356 10810 53390 11586
rect 53814 10810 53848 11586
rect 53944 10810 53978 11586
rect 54402 10810 54436 11586
rect 54532 10810 54566 11586
rect 54990 10810 55024 11586
rect 55120 10810 55154 11586
rect 55578 10810 55612 11586
rect 55708 10810 55742 11586
rect 56166 10810 56200 11586
rect 56296 10810 56330 11586
rect 56754 10810 56788 11586
rect 56884 10810 56918 11586
rect 57342 10810 57376 11586
rect 57472 10810 57506 11586
rect 57930 10810 57964 11586
rect 58060 10810 58094 11586
rect 58518 10810 58552 11586
rect 58648 10810 58682 11586
rect 59106 10810 59140 11586
rect 59236 10810 59270 11586
rect 59694 10810 59728 11586
rect 59824 10810 59858 11586
rect 60282 10810 60316 11586
rect 60412 10810 60446 11586
rect 60870 10810 60904 11586
rect 61000 10810 61034 11586
rect 61458 10810 61492 11586
rect 61588 10810 61622 11586
rect 62046 10810 62080 11586
rect 62176 10810 62210 11586
rect 62634 10810 62668 11586
rect 62764 10810 62798 11586
rect 63222 10810 63256 11586
rect 63352 10810 63386 11586
rect 63810 10810 63844 11586
rect 63940 10810 63974 11586
rect 64398 10810 64432 11586
rect 64528 10810 64562 11586
rect 64986 10810 65020 11586
rect 65116 10810 65150 11586
rect 65574 10810 65608 11586
rect 65704 10810 65738 11586
rect 66162 10810 66196 11586
rect 66292 10810 66326 11586
rect 66750 10810 66784 11586
rect 66880 10810 66914 11586
rect 67338 10810 67372 11586
rect 67468 10810 67502 11586
rect 67926 10810 67960 11586
rect 68056 10810 68090 11586
rect 68514 10810 68548 11586
rect 68644 10810 68678 11586
rect 69102 10810 69136 11586
rect 69232 10810 69266 11586
rect 69690 10810 69724 11586
rect 69820 10810 69854 11586
rect 70278 10810 70312 11586
rect 70408 10810 70442 11586
rect 70866 10810 70900 11586
rect 70996 10810 71030 11586
rect 71454 10810 71488 11586
rect 43422 10717 43790 10751
rect 44010 10717 44378 10751
rect 44598 10717 44966 10751
rect 45186 10717 45554 10751
rect 45774 10717 46142 10751
rect 46362 10717 46730 10751
rect 46950 10717 47318 10751
rect 47538 10717 47906 10751
rect 48126 10717 48494 10751
rect 48714 10717 49082 10751
rect 49302 10717 49670 10751
rect 49890 10717 50258 10751
rect 50478 10717 50846 10751
rect 51066 10717 51434 10751
rect 51654 10717 52022 10751
rect 52242 10717 52610 10751
rect 52830 10717 53198 10751
rect 53418 10717 53786 10751
rect 54006 10717 54374 10751
rect 54594 10717 54962 10751
rect 55182 10717 55550 10751
rect 55770 10717 56138 10751
rect 56358 10717 56726 10751
rect 56946 10717 57314 10751
rect 57534 10717 57902 10751
rect 58122 10717 58490 10751
rect 58710 10717 59078 10751
rect 59298 10717 59666 10751
rect 59886 10717 60254 10751
rect 60474 10717 60842 10751
rect 61062 10717 61430 10751
rect 61650 10717 62018 10751
rect 62238 10717 62606 10751
rect 62826 10717 63194 10751
rect 63414 10717 63782 10751
rect 64002 10717 64370 10751
rect 64590 10717 64958 10751
rect 65178 10717 65546 10751
rect 65766 10717 66134 10751
rect 66354 10717 66722 10751
rect 66942 10717 67310 10751
rect 67530 10717 67898 10751
rect 68118 10717 68486 10751
rect 68706 10717 69074 10751
rect 69294 10717 69662 10751
rect 69882 10717 70250 10751
rect 70470 10717 70838 10751
rect 71058 10717 71426 10751
rect 43422 10645 43790 10679
rect 44010 10645 44378 10679
rect 44598 10645 44966 10679
rect 45186 10645 45554 10679
rect 45774 10645 46142 10679
rect 46362 10645 46730 10679
rect 46950 10645 47318 10679
rect 47538 10645 47906 10679
rect 48126 10645 48494 10679
rect 48714 10645 49082 10679
rect 49302 10645 49670 10679
rect 49890 10645 50258 10679
rect 50478 10645 50846 10679
rect 51066 10645 51434 10679
rect 51654 10645 52022 10679
rect 52242 10645 52610 10679
rect 52830 10645 53198 10679
rect 53418 10645 53786 10679
rect 54006 10645 54374 10679
rect 54594 10645 54962 10679
rect 55182 10645 55550 10679
rect 55770 10645 56138 10679
rect 56358 10645 56726 10679
rect 56946 10645 57314 10679
rect 57534 10645 57902 10679
rect 58122 10645 58490 10679
rect 58710 10645 59078 10679
rect 59298 10645 59666 10679
rect 59886 10645 60254 10679
rect 60474 10645 60842 10679
rect 61062 10645 61430 10679
rect 61650 10645 62018 10679
rect 62238 10645 62606 10679
rect 62826 10645 63194 10679
rect 63414 10645 63782 10679
rect 64002 10645 64370 10679
rect 64590 10645 64958 10679
rect 65178 10645 65546 10679
rect 65766 10645 66134 10679
rect 66354 10645 66722 10679
rect 66942 10645 67310 10679
rect 67530 10645 67898 10679
rect 68118 10645 68486 10679
rect 68706 10645 69074 10679
rect 69294 10645 69662 10679
rect 69882 10645 70250 10679
rect 70470 10645 70838 10679
rect 71058 10645 71426 10679
rect 43360 9810 43394 10586
rect 43818 9810 43852 10586
rect 43948 9810 43982 10586
rect 44406 9810 44440 10586
rect 44536 9810 44570 10586
rect 44994 9810 45028 10586
rect 45124 9810 45158 10586
rect 45582 9810 45616 10586
rect 45712 9810 45746 10586
rect 46170 9810 46204 10586
rect 46300 9810 46334 10586
rect 46758 9810 46792 10586
rect 46888 9810 46922 10586
rect 47346 9810 47380 10586
rect 47476 9810 47510 10586
rect 47934 9810 47968 10586
rect 48064 9810 48098 10586
rect 48522 9810 48556 10586
rect 48652 9810 48686 10586
rect 49110 9810 49144 10586
rect 49240 9810 49274 10586
rect 49698 9810 49732 10586
rect 49828 9810 49862 10586
rect 50286 9810 50320 10586
rect 50416 9810 50450 10586
rect 50874 9810 50908 10586
rect 51004 9810 51038 10586
rect 51462 9810 51496 10586
rect 51592 9810 51626 10586
rect 52050 9810 52084 10586
rect 52180 9810 52214 10586
rect 52638 9810 52672 10586
rect 52768 9810 52802 10586
rect 53226 9810 53260 10586
rect 53356 9810 53390 10586
rect 53814 9810 53848 10586
rect 53944 9810 53978 10586
rect 54402 9810 54436 10586
rect 54532 9810 54566 10586
rect 54990 9810 55024 10586
rect 55120 9810 55154 10586
rect 55578 9810 55612 10586
rect 55708 9810 55742 10586
rect 56166 9810 56200 10586
rect 56296 9810 56330 10586
rect 56754 9810 56788 10586
rect 56884 9810 56918 10586
rect 57342 9810 57376 10586
rect 57472 9810 57506 10586
rect 57930 9810 57964 10586
rect 58060 9810 58094 10586
rect 58518 9810 58552 10586
rect 58648 9810 58682 10586
rect 59106 9810 59140 10586
rect 59236 9810 59270 10586
rect 59694 9810 59728 10586
rect 59824 9810 59858 10586
rect 60282 9810 60316 10586
rect 60412 9810 60446 10586
rect 60870 9810 60904 10586
rect 61000 9810 61034 10586
rect 61458 9810 61492 10586
rect 61588 9810 61622 10586
rect 62046 9810 62080 10586
rect 62176 9810 62210 10586
rect 62634 9810 62668 10586
rect 62764 9810 62798 10586
rect 63222 9810 63256 10586
rect 63352 9810 63386 10586
rect 63810 9810 63844 10586
rect 63940 9810 63974 10586
rect 64398 9810 64432 10586
rect 64528 9810 64562 10586
rect 64986 9810 65020 10586
rect 65116 9810 65150 10586
rect 65574 9810 65608 10586
rect 65704 9810 65738 10586
rect 66162 9810 66196 10586
rect 66292 9810 66326 10586
rect 66750 9810 66784 10586
rect 66880 9810 66914 10586
rect 67338 9810 67372 10586
rect 67468 9810 67502 10586
rect 67926 9810 67960 10586
rect 68056 9810 68090 10586
rect 68514 9810 68548 10586
rect 68644 9810 68678 10586
rect 69102 9810 69136 10586
rect 69232 9810 69266 10586
rect 69690 9810 69724 10586
rect 69820 9810 69854 10586
rect 70278 9810 70312 10586
rect 70408 9810 70442 10586
rect 70866 9810 70900 10586
rect 70996 9810 71030 10586
rect 71454 9810 71488 10586
rect 43422 9717 43790 9751
rect 44010 9717 44378 9751
rect 44598 9717 44966 9751
rect 45186 9717 45554 9751
rect 45774 9717 46142 9751
rect 46362 9717 46730 9751
rect 46950 9717 47318 9751
rect 47538 9717 47906 9751
rect 48126 9717 48494 9751
rect 48714 9717 49082 9751
rect 49302 9717 49670 9751
rect 49890 9717 50258 9751
rect 50478 9717 50846 9751
rect 51066 9717 51434 9751
rect 51654 9717 52022 9751
rect 52242 9717 52610 9751
rect 52830 9717 53198 9751
rect 53418 9717 53786 9751
rect 54006 9717 54374 9751
rect 54594 9717 54962 9751
rect 55182 9717 55550 9751
rect 55770 9717 56138 9751
rect 56358 9717 56726 9751
rect 56946 9717 57314 9751
rect 57534 9717 57902 9751
rect 58122 9717 58490 9751
rect 58710 9717 59078 9751
rect 59298 9717 59666 9751
rect 59886 9717 60254 9751
rect 60474 9717 60842 9751
rect 61062 9717 61430 9751
rect 61650 9717 62018 9751
rect 62238 9717 62606 9751
rect 62826 9717 63194 9751
rect 63414 9717 63782 9751
rect 64002 9717 64370 9751
rect 64590 9717 64958 9751
rect 65178 9717 65546 9751
rect 65766 9717 66134 9751
rect 66354 9717 66722 9751
rect 66942 9717 67310 9751
rect 67530 9717 67898 9751
rect 68118 9717 68486 9751
rect 68706 9717 69074 9751
rect 69294 9717 69662 9751
rect 69882 9717 70250 9751
rect 70470 9717 70838 9751
rect 71058 9717 71426 9751
rect 43806 9400 43994 9448
rect 44982 9400 45170 9448
rect 46158 9400 46346 9448
rect 47334 9400 47522 9448
rect 48510 9400 48698 9448
rect 49686 9400 49874 9448
rect 50862 9400 51050 9448
rect 52038 9400 52226 9448
rect 53214 9400 53402 9448
rect 54390 9400 54578 9448
rect 55566 9400 55754 9448
rect 56742 9400 56930 9448
rect 57918 9400 58106 9448
rect 59094 9400 59282 9448
rect 60270 9400 60458 9448
rect 61446 9400 61634 9448
rect 62622 9400 62810 9458
rect 63798 9400 63986 9448
rect 64974 9400 65162 9448
rect 66150 9400 66338 9448
rect 67312 9400 67524 9458
rect 68502 9400 68690 9448
rect 69678 9400 69866 9448
rect 70854 9400 71042 9448
rect 43806 9366 43994 9400
rect 44982 9366 45170 9400
rect 46158 9366 46346 9400
rect 47334 9366 47522 9400
rect 48510 9366 48698 9400
rect 49686 9366 49874 9400
rect 50862 9366 51050 9400
rect 52038 9366 52226 9400
rect 53214 9366 53402 9400
rect 54390 9366 54578 9400
rect 55566 9366 55754 9400
rect 56742 9366 56930 9400
rect 57918 9366 58106 9400
rect 59094 9366 59282 9400
rect 60270 9366 60458 9400
rect 61446 9366 61634 9400
rect 62622 9366 62810 9400
rect 63798 9366 63986 9400
rect 64974 9366 65162 9400
rect 66150 9366 66338 9400
rect 67312 9366 67524 9400
rect 68502 9366 68690 9400
rect 69678 9366 69866 9400
rect 70854 9366 71042 9400
rect 43806 9338 43994 9366
rect 44982 9338 45170 9366
rect 46158 9338 46346 9366
rect 47334 9338 47522 9366
rect 48510 9338 48698 9366
rect 49686 9338 49874 9366
rect 50862 9338 51050 9366
rect 52038 9338 52226 9366
rect 53214 9338 53402 9366
rect 54390 9338 54578 9366
rect 55566 9338 55754 9366
rect 56742 9338 56930 9366
rect 57918 9338 58106 9366
rect 59094 9338 59282 9366
rect 60270 9338 60458 9366
rect 61446 9338 61634 9366
rect 62622 9348 62810 9366
rect 63798 9338 63986 9366
rect 64974 9338 65162 9366
rect 66150 9338 66338 9366
rect 67312 9336 67524 9366
rect 68502 9338 68690 9366
rect 69678 9338 69866 9366
rect 70854 9338 71042 9366
rect 56474 8190 56512 8322
rect 56740 8190 56778 8322
rect 57006 8190 57044 8322
rect 57272 8190 57310 8322
rect 57538 8190 57576 8322
rect 57804 8190 57842 8322
rect 58070 8190 58108 8322
rect 58336 8190 58374 8322
rect 56412 7364 56446 8140
rect 56540 7364 56574 8140
rect 56678 7364 56712 8140
rect 56806 7364 56840 8140
rect 56944 7364 56978 8140
rect 57072 7364 57106 8140
rect 57210 7364 57244 8140
rect 57338 7364 57372 8140
rect 57476 7364 57510 8140
rect 57604 7364 57638 8140
rect 57742 7364 57776 8140
rect 57870 7364 57904 8140
rect 58008 7364 58042 8140
rect 58136 7364 58170 8140
rect 58274 7364 58308 8140
rect 58402 7364 58436 8140
rect 56474 7180 56512 7312
rect 56740 7180 56778 7312
rect 57006 7180 57044 7312
rect 57272 7180 57310 7312
rect 57538 7180 57576 7312
rect 57804 7180 57842 7312
rect 58070 7180 58108 7312
rect 58336 7180 58374 7312
rect 56412 6354 56446 7130
rect 56540 6354 56574 7130
rect 56678 6354 56712 7130
rect 56806 6354 56840 7130
rect 56944 6354 56978 7130
rect 57072 6354 57106 7130
rect 57210 6354 57244 7130
rect 57338 6354 57372 7130
rect 57476 6354 57510 7130
rect 57604 6354 57638 7130
rect 57742 6354 57776 7130
rect 57870 6354 57904 7130
rect 58008 6354 58042 7130
rect 58136 6354 58170 7130
rect 58274 6354 58308 7130
rect 58402 6354 58436 7130
rect 56474 6170 56512 6302
rect 56740 6170 56778 6302
rect 57006 6170 57044 6302
rect 57272 6170 57310 6302
rect 57538 6170 57576 6302
rect 57804 6170 57842 6302
rect 58070 6170 58108 6302
rect 58336 6170 58374 6302
rect 56412 5344 56446 6120
rect 56540 5344 56574 6120
rect 56678 5344 56712 6120
rect 56806 5344 56840 6120
rect 56944 5344 56978 6120
rect 57072 5344 57106 6120
rect 57210 5344 57244 6120
rect 57338 5344 57372 6120
rect 57476 5344 57510 6120
rect 57604 5344 57638 6120
rect 57742 5344 57776 6120
rect 57870 5344 57904 6120
rect 58008 5344 58042 6120
rect 58136 5344 58170 6120
rect 58274 5344 58308 6120
rect 58402 5344 58436 6120
rect 56474 5160 56512 5292
rect 56740 5160 56778 5292
rect 57006 5160 57044 5292
rect 57272 5160 57310 5292
rect 57538 5160 57576 5292
rect 57804 5160 57842 5292
rect 58070 5160 58108 5292
rect 58336 5160 58374 5292
rect 57046 3998 57084 4124
rect 57286 3998 57324 4124
rect 57526 3998 57564 4124
rect 57766 3998 57804 4124
rect 56984 3372 57018 3948
rect 57112 3372 57146 3948
rect 57224 3372 57258 3948
rect 57352 3372 57386 3948
rect 57464 3372 57498 3948
rect 57592 3372 57626 3948
rect 57704 3372 57738 3948
rect 57832 3372 57866 3948
rect 57046 3190 57084 3322
rect 57286 3190 57324 3322
rect 57526 3190 57564 3322
rect 57766 3190 57804 3322
rect 56984 2564 57018 3140
rect 57112 2564 57146 3140
rect 57224 2564 57258 3140
rect 57352 2564 57386 3140
rect 57464 2564 57498 3140
rect 57592 2564 57626 3140
rect 57704 2564 57738 3140
rect 57832 2564 57866 3140
rect 57046 2382 57084 2514
rect 57286 2382 57324 2514
rect 57526 2382 57564 2514
rect 57766 2382 57804 2514
rect 56736 2082 58088 2130
rect 56736 2048 56796 2082
rect 56796 2048 58006 2082
rect 58006 2048 58088 2082
rect 56736 2018 58088 2048
<< metal1 >>
rect 52798 17186 52932 17192
rect 52798 17114 52810 17186
rect 52920 17114 52932 17186
rect 52798 17108 52932 17114
rect 53278 17186 53412 17192
rect 53278 17114 53290 17186
rect 53400 17114 53412 17186
rect 53278 17108 53412 17114
rect 53758 17186 53892 17192
rect 53758 17114 53770 17186
rect 53880 17114 53892 17186
rect 53758 17108 53892 17114
rect 54238 17186 54372 17192
rect 54238 17114 54250 17186
rect 54360 17114 54372 17186
rect 54238 17108 54372 17114
rect 54718 17186 54852 17192
rect 54718 17114 54730 17186
rect 54840 17114 54852 17186
rect 54718 17108 54852 17114
rect 55198 17186 55332 17192
rect 55198 17114 55210 17186
rect 55320 17114 55332 17186
rect 55198 17108 55332 17114
rect 55678 17186 55812 17192
rect 55678 17114 55690 17186
rect 55800 17114 55812 17186
rect 55678 17108 55812 17114
rect 56158 17186 56292 17192
rect 56158 17114 56170 17186
rect 56280 17114 56292 17186
rect 56158 17108 56292 17114
rect 56638 17186 56772 17192
rect 56638 17114 56650 17186
rect 56760 17114 56772 17186
rect 56638 17108 56772 17114
rect 57118 17186 57252 17192
rect 57118 17114 57130 17186
rect 57240 17114 57252 17186
rect 57118 17108 57252 17114
rect 57598 17186 57732 17192
rect 57598 17114 57610 17186
rect 57720 17114 57732 17186
rect 57598 17108 57732 17114
rect 58078 17186 58212 17192
rect 58078 17114 58090 17186
rect 58200 17114 58212 17186
rect 58078 17108 58212 17114
rect 58558 17186 58692 17192
rect 58558 17114 58570 17186
rect 58680 17114 58692 17186
rect 58558 17108 58692 17114
rect 59038 17186 59172 17192
rect 59038 17114 59050 17186
rect 59160 17114 59172 17186
rect 59038 17108 59172 17114
rect 59518 17186 59652 17192
rect 59518 17114 59530 17186
rect 59640 17114 59652 17186
rect 59518 17108 59652 17114
rect 59998 17186 60132 17192
rect 59998 17114 60010 17186
rect 60120 17114 60132 17186
rect 59998 17108 60132 17114
rect 60478 17186 60612 17192
rect 60478 17114 60490 17186
rect 60600 17114 60612 17186
rect 60478 17108 60612 17114
rect 60958 17186 61092 17192
rect 60958 17114 60970 17186
rect 61080 17114 61092 17186
rect 60958 17108 61092 17114
rect 61438 17186 61572 17192
rect 61438 17114 61450 17186
rect 61560 17114 61572 17186
rect 61438 17108 61572 17114
rect 61918 17186 62052 17192
rect 61918 17114 61930 17186
rect 62040 17114 62052 17186
rect 61918 17108 62052 17114
rect 52710 16842 52780 16848
rect 52700 16710 52710 16842
rect 52780 16710 52790 16842
rect 52710 16704 52780 16710
rect 52838 16672 52892 17108
rect 52950 16842 53020 16848
rect 52940 16710 52950 16842
rect 53020 16710 53030 16842
rect 52950 16704 53020 16710
rect 53078 16700 53132 16852
rect 53190 16842 53260 16848
rect 53180 16710 53190 16842
rect 53260 16710 53270 16842
rect 53190 16704 53260 16710
rect 53318 16672 53372 17108
rect 53430 16842 53500 16848
rect 53420 16710 53430 16842
rect 53500 16710 53510 16842
rect 53430 16704 53500 16710
rect 53558 16700 53612 16852
rect 53670 16842 53740 16848
rect 53660 16710 53670 16842
rect 53740 16710 53750 16842
rect 53670 16704 53740 16710
rect 53798 16672 53852 17108
rect 53910 16842 53980 16848
rect 53900 16710 53910 16842
rect 53980 16710 53990 16842
rect 53910 16704 53980 16710
rect 54038 16700 54092 16852
rect 54150 16842 54220 16848
rect 54140 16710 54150 16842
rect 54220 16710 54230 16842
rect 54150 16704 54220 16710
rect 54278 16672 54332 17108
rect 54390 16842 54460 16848
rect 54380 16710 54390 16842
rect 54460 16710 54470 16842
rect 54390 16704 54460 16710
rect 54518 16700 54572 16852
rect 54630 16842 54700 16848
rect 54620 16710 54630 16842
rect 54700 16710 54710 16842
rect 54630 16704 54700 16710
rect 54758 16672 54812 17108
rect 54870 16842 54940 16848
rect 54860 16710 54870 16842
rect 54940 16710 54950 16842
rect 54870 16704 54940 16710
rect 54998 16700 55052 16852
rect 55110 16842 55180 16848
rect 55100 16710 55110 16842
rect 55180 16710 55190 16842
rect 55110 16704 55180 16710
rect 55238 16672 55292 17108
rect 55350 16842 55420 16848
rect 55340 16710 55350 16842
rect 55420 16710 55430 16842
rect 55350 16704 55420 16710
rect 55478 16700 55532 16852
rect 55590 16842 55660 16848
rect 55580 16710 55590 16842
rect 55660 16710 55670 16842
rect 55590 16704 55660 16710
rect 55718 16672 55772 17108
rect 55830 16842 55900 16848
rect 55820 16710 55830 16842
rect 55900 16710 55910 16842
rect 55830 16704 55900 16710
rect 55958 16700 56012 16852
rect 56070 16842 56140 16848
rect 56060 16710 56070 16842
rect 56140 16710 56150 16842
rect 56070 16704 56140 16710
rect 56198 16672 56252 17108
rect 56310 16842 56380 16848
rect 56300 16710 56310 16842
rect 56380 16710 56390 16842
rect 56310 16704 56380 16710
rect 56438 16700 56492 16852
rect 56550 16842 56620 16848
rect 56540 16710 56550 16842
rect 56620 16710 56630 16842
rect 56550 16704 56620 16710
rect 56678 16672 56732 17108
rect 56790 16842 56860 16848
rect 56780 16710 56790 16842
rect 56860 16710 56870 16842
rect 56790 16704 56860 16710
rect 56918 16700 56972 16852
rect 57030 16842 57100 16848
rect 57020 16710 57030 16842
rect 57100 16710 57110 16842
rect 57030 16704 57100 16710
rect 57158 16672 57212 17108
rect 57270 16842 57340 16848
rect 57260 16710 57270 16842
rect 57340 16710 57350 16842
rect 57270 16704 57340 16710
rect 57398 16700 57452 16852
rect 57510 16842 57580 16848
rect 57500 16710 57510 16842
rect 57580 16710 57590 16842
rect 57510 16704 57580 16710
rect 57638 16672 57692 17108
rect 57750 16842 57820 16848
rect 57740 16710 57750 16842
rect 57820 16710 57830 16842
rect 57750 16704 57820 16710
rect 57878 16700 57932 16852
rect 57990 16842 58060 16848
rect 57980 16710 57990 16842
rect 58060 16710 58070 16842
rect 57990 16704 58060 16710
rect 58118 16672 58172 17108
rect 58230 16842 58300 16848
rect 58220 16710 58230 16842
rect 58300 16710 58310 16842
rect 58230 16704 58300 16710
rect 58358 16700 58412 16852
rect 58470 16842 58540 16848
rect 58460 16710 58470 16842
rect 58540 16710 58550 16842
rect 58470 16704 58540 16710
rect 58598 16672 58652 17108
rect 58710 16842 58780 16848
rect 58700 16710 58710 16842
rect 58780 16710 58790 16842
rect 58710 16704 58780 16710
rect 58838 16700 58892 16852
rect 58950 16842 59020 16848
rect 58940 16710 58950 16842
rect 59020 16710 59030 16842
rect 58950 16704 59020 16710
rect 59078 16672 59132 17108
rect 59190 16842 59260 16848
rect 59180 16710 59190 16842
rect 59260 16710 59270 16842
rect 59190 16704 59260 16710
rect 59318 16700 59372 16852
rect 59430 16842 59500 16848
rect 59420 16710 59430 16842
rect 59500 16710 59510 16842
rect 59430 16704 59500 16710
rect 59558 16672 59612 17108
rect 59670 16842 59740 16848
rect 59660 16710 59670 16842
rect 59740 16710 59750 16842
rect 59670 16704 59740 16710
rect 59798 16700 59852 16852
rect 59910 16842 59980 16848
rect 59900 16710 59910 16842
rect 59980 16710 59990 16842
rect 59910 16704 59980 16710
rect 60038 16672 60092 17108
rect 60150 16842 60220 16848
rect 60140 16710 60150 16842
rect 60220 16710 60230 16842
rect 60150 16704 60220 16710
rect 60278 16700 60332 16852
rect 60390 16842 60460 16848
rect 60380 16710 60390 16842
rect 60460 16710 60470 16842
rect 60390 16704 60460 16710
rect 60518 16672 60572 17108
rect 60630 16842 60700 16848
rect 60620 16710 60630 16842
rect 60700 16710 60710 16842
rect 60630 16704 60700 16710
rect 60758 16700 60812 16852
rect 60870 16842 60940 16848
rect 60860 16710 60870 16842
rect 60940 16710 60950 16842
rect 60870 16704 60940 16710
rect 60998 16672 61052 17108
rect 61110 16842 61180 16848
rect 61100 16710 61110 16842
rect 61180 16710 61190 16842
rect 61110 16704 61180 16710
rect 61238 16700 61292 16852
rect 61350 16842 61420 16848
rect 61340 16710 61350 16842
rect 61420 16710 61430 16842
rect 61350 16704 61420 16710
rect 61478 16672 61532 17108
rect 61590 16842 61660 16848
rect 61580 16710 61590 16842
rect 61660 16710 61670 16842
rect 61590 16704 61660 16710
rect 61718 16700 61772 16852
rect 61830 16842 61900 16848
rect 61820 16710 61830 16842
rect 61900 16710 61910 16842
rect 61830 16704 61900 16710
rect 61958 16672 62012 17108
rect 62070 16842 62140 16848
rect 62060 16710 62070 16842
rect 62140 16710 62150 16842
rect 62070 16704 62140 16710
rect 52586 16660 52704 16672
rect 52586 16084 52664 16660
rect 52698 16084 52704 16660
rect 52586 16072 52704 16084
rect 52786 16660 52944 16672
rect 52786 16084 52792 16660
rect 52826 16084 52904 16660
rect 52938 16084 52944 16660
rect 52786 16072 52944 16084
rect 53026 16660 53184 16672
rect 53026 16084 53032 16660
rect 53066 16084 53144 16660
rect 53178 16084 53184 16660
rect 53026 16072 53184 16084
rect 53266 16660 53424 16672
rect 53266 16084 53272 16660
rect 53306 16084 53384 16660
rect 53418 16084 53424 16660
rect 53266 16072 53424 16084
rect 53506 16660 53664 16672
rect 53506 16084 53512 16660
rect 53546 16084 53624 16660
rect 53658 16084 53664 16660
rect 53506 16072 53664 16084
rect 53746 16660 53904 16672
rect 53746 16084 53752 16660
rect 53786 16084 53864 16660
rect 53898 16084 53904 16660
rect 53746 16072 53904 16084
rect 53986 16660 54144 16672
rect 53986 16084 53992 16660
rect 54026 16084 54104 16660
rect 54138 16084 54144 16660
rect 53986 16072 54144 16084
rect 54226 16660 54384 16672
rect 54226 16084 54232 16660
rect 54266 16084 54344 16660
rect 54378 16084 54384 16660
rect 54226 16072 54384 16084
rect 54466 16660 54624 16672
rect 54466 16084 54472 16660
rect 54506 16084 54584 16660
rect 54618 16084 54624 16660
rect 54466 16072 54624 16084
rect 54706 16660 54864 16672
rect 54706 16084 54712 16660
rect 54746 16084 54824 16660
rect 54858 16084 54864 16660
rect 54706 16072 54864 16084
rect 54946 16660 55104 16672
rect 54946 16084 54952 16660
rect 54986 16084 55064 16660
rect 55098 16084 55104 16660
rect 54946 16072 55104 16084
rect 55186 16660 55344 16672
rect 55186 16084 55192 16660
rect 55226 16084 55304 16660
rect 55338 16084 55344 16660
rect 55186 16072 55344 16084
rect 55426 16660 55584 16672
rect 55426 16084 55432 16660
rect 55466 16084 55544 16660
rect 55578 16084 55584 16660
rect 55426 16072 55584 16084
rect 55666 16660 55824 16672
rect 55666 16084 55672 16660
rect 55706 16084 55784 16660
rect 55818 16084 55824 16660
rect 55666 16072 55824 16084
rect 55906 16660 56064 16672
rect 55906 16084 55912 16660
rect 55946 16084 56024 16660
rect 56058 16084 56064 16660
rect 55906 16072 56064 16084
rect 56146 16660 56304 16672
rect 56146 16084 56152 16660
rect 56186 16084 56264 16660
rect 56298 16084 56304 16660
rect 56146 16072 56304 16084
rect 56386 16660 56544 16672
rect 56386 16084 56392 16660
rect 56426 16084 56504 16660
rect 56538 16084 56544 16660
rect 56386 16072 56544 16084
rect 56626 16660 56784 16672
rect 56626 16084 56632 16660
rect 56666 16084 56744 16660
rect 56778 16084 56784 16660
rect 56626 16072 56784 16084
rect 56866 16660 57024 16672
rect 56866 16084 56872 16660
rect 56906 16084 56984 16660
rect 57018 16084 57024 16660
rect 56866 16072 57024 16084
rect 57106 16660 57264 16672
rect 57106 16084 57112 16660
rect 57146 16084 57224 16660
rect 57258 16084 57264 16660
rect 57106 16072 57264 16084
rect 57346 16660 57504 16672
rect 57346 16084 57352 16660
rect 57386 16084 57464 16660
rect 57498 16084 57504 16660
rect 57346 16072 57504 16084
rect 57586 16660 57744 16672
rect 57586 16084 57592 16660
rect 57626 16084 57704 16660
rect 57738 16084 57744 16660
rect 57586 16072 57744 16084
rect 57826 16660 57984 16672
rect 57826 16084 57832 16660
rect 57866 16084 57944 16660
rect 57978 16084 57984 16660
rect 57826 16072 57984 16084
rect 58066 16660 58224 16672
rect 58066 16084 58072 16660
rect 58106 16084 58184 16660
rect 58218 16084 58224 16660
rect 58066 16072 58224 16084
rect 58306 16660 58464 16672
rect 58306 16084 58312 16660
rect 58346 16084 58424 16660
rect 58458 16084 58464 16660
rect 58306 16072 58464 16084
rect 58546 16660 58704 16672
rect 58546 16084 58552 16660
rect 58586 16084 58664 16660
rect 58698 16084 58704 16660
rect 58546 16072 58704 16084
rect 58786 16660 58944 16672
rect 58786 16084 58792 16660
rect 58826 16084 58904 16660
rect 58938 16084 58944 16660
rect 58786 16072 58944 16084
rect 59026 16660 59184 16672
rect 59026 16084 59032 16660
rect 59066 16084 59144 16660
rect 59178 16084 59184 16660
rect 59026 16072 59184 16084
rect 59266 16660 59424 16672
rect 59266 16084 59272 16660
rect 59306 16084 59384 16660
rect 59418 16084 59424 16660
rect 59266 16072 59424 16084
rect 59506 16660 59664 16672
rect 59506 16084 59512 16660
rect 59546 16084 59624 16660
rect 59658 16084 59664 16660
rect 59506 16072 59664 16084
rect 59746 16660 59904 16672
rect 59746 16084 59752 16660
rect 59786 16084 59864 16660
rect 59898 16084 59904 16660
rect 59746 16072 59904 16084
rect 59986 16660 60144 16672
rect 59986 16084 59992 16660
rect 60026 16084 60104 16660
rect 60138 16084 60144 16660
rect 59986 16072 60144 16084
rect 60226 16660 60384 16672
rect 60226 16084 60232 16660
rect 60266 16084 60344 16660
rect 60378 16084 60384 16660
rect 60226 16072 60384 16084
rect 60466 16660 60624 16672
rect 60466 16084 60472 16660
rect 60506 16084 60584 16660
rect 60618 16084 60624 16660
rect 60466 16072 60624 16084
rect 60706 16660 60864 16672
rect 60706 16084 60712 16660
rect 60746 16084 60824 16660
rect 60858 16084 60864 16660
rect 60706 16072 60864 16084
rect 60946 16660 61104 16672
rect 60946 16084 60952 16660
rect 60986 16084 61064 16660
rect 61098 16084 61104 16660
rect 60946 16072 61104 16084
rect 61186 16660 61344 16672
rect 61186 16084 61192 16660
rect 61226 16084 61304 16660
rect 61338 16084 61344 16660
rect 61186 16072 61344 16084
rect 61426 16660 61584 16672
rect 61426 16084 61432 16660
rect 61466 16084 61544 16660
rect 61578 16084 61584 16660
rect 61426 16072 61584 16084
rect 61666 16660 61824 16672
rect 61666 16084 61672 16660
rect 61706 16084 61784 16660
rect 61818 16084 61824 16660
rect 61666 16072 61824 16084
rect 61906 16660 62064 16672
rect 61906 16084 61912 16660
rect 61946 16084 62024 16660
rect 62058 16084 62064 16660
rect 61906 16072 62064 16084
rect 62146 16660 62264 16672
rect 62146 16084 62152 16660
rect 62186 16084 62264 16660
rect 62146 16072 62264 16084
rect 52586 15864 52664 16072
rect 52710 16034 52780 16040
rect 52700 15902 52710 16034
rect 52780 15902 52790 16034
rect 52710 15896 52780 15902
rect 52832 15864 52898 16072
rect 52950 16034 53020 16040
rect 52940 15902 52950 16034
rect 53020 15902 53030 16034
rect 52950 15896 53020 15902
rect 53072 15864 53138 16072
rect 53190 16034 53260 16040
rect 53180 15902 53190 16034
rect 53260 15902 53270 16034
rect 53190 15896 53260 15902
rect 53312 15864 53378 16072
rect 53430 16034 53500 16040
rect 53420 15902 53430 16034
rect 53500 15902 53510 16034
rect 53430 15896 53500 15902
rect 53546 15864 53624 16072
rect 53670 16034 53740 16040
rect 53660 15902 53670 16034
rect 53740 15902 53750 16034
rect 53670 15896 53740 15902
rect 53792 15864 53858 16072
rect 53910 16034 53980 16040
rect 53900 15902 53910 16034
rect 53980 15902 53990 16034
rect 53910 15896 53980 15902
rect 54032 15864 54098 16072
rect 54150 16034 54220 16040
rect 54140 15902 54150 16034
rect 54220 15902 54230 16034
rect 54150 15896 54220 15902
rect 54272 15864 54338 16072
rect 54390 16034 54460 16040
rect 54380 15902 54390 16034
rect 54460 15902 54470 16034
rect 54390 15896 54460 15902
rect 54506 15864 54584 16072
rect 54630 16034 54700 16040
rect 54620 15902 54630 16034
rect 54700 15902 54710 16034
rect 54630 15896 54700 15902
rect 54752 15864 54818 16072
rect 54870 16034 54940 16040
rect 54860 15902 54870 16034
rect 54940 15902 54950 16034
rect 54870 15896 54940 15902
rect 54992 15864 55058 16072
rect 55110 16034 55180 16040
rect 55100 15902 55110 16034
rect 55180 15902 55190 16034
rect 55110 15896 55180 15902
rect 55232 15864 55298 16072
rect 55350 16034 55420 16040
rect 55340 15902 55350 16034
rect 55420 15902 55430 16034
rect 55350 15896 55420 15902
rect 55466 15864 55544 16072
rect 55590 16034 55660 16040
rect 55580 15902 55590 16034
rect 55660 15902 55670 16034
rect 55590 15896 55660 15902
rect 55712 15864 55778 16072
rect 55830 16034 55900 16040
rect 55820 15902 55830 16034
rect 55900 15902 55910 16034
rect 55830 15896 55900 15902
rect 55952 15864 56018 16072
rect 56070 16034 56140 16040
rect 56060 15902 56070 16034
rect 56140 15902 56150 16034
rect 56070 15896 56140 15902
rect 56192 15864 56258 16072
rect 56310 16034 56380 16040
rect 56300 15902 56310 16034
rect 56380 15902 56390 16034
rect 56310 15896 56380 15902
rect 56426 15864 56504 16072
rect 56550 16034 56620 16040
rect 56540 15902 56550 16034
rect 56620 15902 56630 16034
rect 56550 15896 56620 15902
rect 56672 15864 56738 16072
rect 56790 16034 56860 16040
rect 56780 15902 56790 16034
rect 56860 15902 56870 16034
rect 56790 15896 56860 15902
rect 56912 15864 56978 16072
rect 57030 16034 57100 16040
rect 57020 15902 57030 16034
rect 57100 15902 57110 16034
rect 57030 15896 57100 15902
rect 57152 15864 57218 16072
rect 57270 16034 57340 16040
rect 57260 15902 57270 16034
rect 57340 15902 57350 16034
rect 57270 15896 57340 15902
rect 57386 15864 57464 16072
rect 57510 16034 57580 16040
rect 57500 15902 57510 16034
rect 57580 15902 57590 16034
rect 57510 15896 57580 15902
rect 57632 15864 57698 16072
rect 57750 16034 57820 16040
rect 57740 15902 57750 16034
rect 57820 15902 57830 16034
rect 57750 15896 57820 15902
rect 57872 15864 57938 16072
rect 57990 16034 58060 16040
rect 57980 15902 57990 16034
rect 58060 15902 58070 16034
rect 57990 15896 58060 15902
rect 58112 15864 58178 16072
rect 58230 16034 58300 16040
rect 58220 15902 58230 16034
rect 58300 15902 58310 16034
rect 58230 15896 58300 15902
rect 58346 15864 58424 16072
rect 58470 16034 58540 16040
rect 58460 15902 58470 16034
rect 58540 15902 58550 16034
rect 58470 15896 58540 15902
rect 58592 15864 58658 16072
rect 58710 16034 58780 16040
rect 58700 15902 58710 16034
rect 58780 15902 58790 16034
rect 58710 15896 58780 15902
rect 58832 15864 58898 16072
rect 58950 16034 59020 16040
rect 58940 15902 58950 16034
rect 59020 15902 59030 16034
rect 58950 15896 59020 15902
rect 59072 15864 59138 16072
rect 59190 16034 59260 16040
rect 59180 15902 59190 16034
rect 59260 15902 59270 16034
rect 59190 15896 59260 15902
rect 59306 15864 59384 16072
rect 59430 16034 59500 16040
rect 59420 15902 59430 16034
rect 59500 15902 59510 16034
rect 59430 15896 59500 15902
rect 59552 15864 59618 16072
rect 59670 16034 59740 16040
rect 59660 15902 59670 16034
rect 59740 15902 59750 16034
rect 59670 15896 59740 15902
rect 59792 15864 59858 16072
rect 59910 16034 59980 16040
rect 59900 15902 59910 16034
rect 59980 15902 59990 16034
rect 59910 15896 59980 15902
rect 60032 15864 60098 16072
rect 60150 16034 60220 16040
rect 60140 15902 60150 16034
rect 60220 15902 60230 16034
rect 60150 15896 60220 15902
rect 60266 15864 60344 16072
rect 60390 16034 60460 16040
rect 60380 15902 60390 16034
rect 60460 15902 60470 16034
rect 60390 15896 60460 15902
rect 60512 15864 60578 16072
rect 60630 16034 60700 16040
rect 60620 15902 60630 16034
rect 60700 15902 60710 16034
rect 60630 15896 60700 15902
rect 60752 15864 60818 16072
rect 60870 16034 60940 16040
rect 60860 15902 60870 16034
rect 60940 15902 60950 16034
rect 60870 15896 60940 15902
rect 60992 15864 61058 16072
rect 61110 16034 61180 16040
rect 61100 15902 61110 16034
rect 61180 15902 61190 16034
rect 61110 15896 61180 15902
rect 61226 15864 61304 16072
rect 61350 16034 61420 16040
rect 61340 15902 61350 16034
rect 61420 15902 61430 16034
rect 61350 15896 61420 15902
rect 61472 15864 61538 16072
rect 61590 16034 61660 16040
rect 61580 15902 61590 16034
rect 61660 15902 61670 16034
rect 61590 15896 61660 15902
rect 61712 15864 61778 16072
rect 61830 16034 61900 16040
rect 61820 15902 61830 16034
rect 61900 15902 61910 16034
rect 61830 15896 61900 15902
rect 61952 15864 62018 16072
rect 62070 16034 62140 16040
rect 62060 15902 62070 16034
rect 62140 15902 62150 16034
rect 62070 15896 62140 15902
rect 62186 15864 62264 16072
rect 52586 15852 52704 15864
rect 52586 15276 52664 15852
rect 52698 15276 52704 15852
rect 52586 15264 52704 15276
rect 52786 15852 52944 15864
rect 52786 15276 52792 15852
rect 52826 15276 52904 15852
rect 52938 15276 52944 15852
rect 52786 15264 52944 15276
rect 53026 15852 53184 15864
rect 53026 15276 53032 15852
rect 53066 15276 53144 15852
rect 53178 15276 53184 15852
rect 53026 15264 53184 15276
rect 53266 15852 53424 15864
rect 53266 15276 53272 15852
rect 53306 15276 53384 15852
rect 53418 15276 53424 15852
rect 53266 15264 53424 15276
rect 53506 15852 53664 15864
rect 53506 15276 53512 15852
rect 53546 15276 53624 15852
rect 53658 15276 53664 15852
rect 53506 15264 53664 15276
rect 53746 15852 53904 15864
rect 53746 15276 53752 15852
rect 53786 15276 53864 15852
rect 53898 15276 53904 15852
rect 53746 15264 53904 15276
rect 53986 15852 54144 15864
rect 53986 15276 53992 15852
rect 54026 15276 54104 15852
rect 54138 15276 54144 15852
rect 53986 15264 54144 15276
rect 54226 15852 54384 15864
rect 54226 15276 54232 15852
rect 54266 15276 54344 15852
rect 54378 15276 54384 15852
rect 54226 15264 54384 15276
rect 54466 15852 54624 15864
rect 54466 15276 54472 15852
rect 54506 15276 54584 15852
rect 54618 15276 54624 15852
rect 54466 15264 54624 15276
rect 54706 15852 54864 15864
rect 54706 15276 54712 15852
rect 54746 15276 54824 15852
rect 54858 15276 54864 15852
rect 54706 15264 54864 15276
rect 54946 15852 55104 15864
rect 54946 15276 54952 15852
rect 54986 15276 55064 15852
rect 55098 15276 55104 15852
rect 54946 15264 55104 15276
rect 55186 15852 55344 15864
rect 55186 15276 55192 15852
rect 55226 15276 55304 15852
rect 55338 15276 55344 15852
rect 55186 15264 55344 15276
rect 55426 15852 55584 15864
rect 55426 15276 55432 15852
rect 55466 15276 55544 15852
rect 55578 15276 55584 15852
rect 55426 15264 55584 15276
rect 55666 15852 55824 15864
rect 55666 15276 55672 15852
rect 55706 15276 55784 15852
rect 55818 15276 55824 15852
rect 55666 15264 55824 15276
rect 55906 15852 56064 15864
rect 55906 15276 55912 15852
rect 55946 15276 56024 15852
rect 56058 15276 56064 15852
rect 55906 15264 56064 15276
rect 56146 15852 56304 15864
rect 56146 15276 56152 15852
rect 56186 15276 56264 15852
rect 56298 15276 56304 15852
rect 56146 15264 56304 15276
rect 56386 15852 56544 15864
rect 56386 15276 56392 15852
rect 56426 15276 56504 15852
rect 56538 15276 56544 15852
rect 56386 15264 56544 15276
rect 56626 15852 56784 15864
rect 56626 15276 56632 15852
rect 56666 15276 56744 15852
rect 56778 15276 56784 15852
rect 56626 15264 56784 15276
rect 56866 15852 57024 15864
rect 56866 15276 56872 15852
rect 56906 15276 56984 15852
rect 57018 15276 57024 15852
rect 56866 15264 57024 15276
rect 57106 15852 57264 15864
rect 57106 15276 57112 15852
rect 57146 15276 57224 15852
rect 57258 15276 57264 15852
rect 57106 15264 57264 15276
rect 57346 15852 57504 15864
rect 57346 15276 57352 15852
rect 57386 15276 57464 15852
rect 57498 15276 57504 15852
rect 57346 15264 57504 15276
rect 57586 15852 57744 15864
rect 57586 15276 57592 15852
rect 57626 15276 57704 15852
rect 57738 15276 57744 15852
rect 57586 15264 57744 15276
rect 57826 15852 57984 15864
rect 57826 15276 57832 15852
rect 57866 15276 57944 15852
rect 57978 15276 57984 15852
rect 57826 15264 57984 15276
rect 58066 15852 58224 15864
rect 58066 15276 58072 15852
rect 58106 15276 58184 15852
rect 58218 15276 58224 15852
rect 58066 15264 58224 15276
rect 58306 15852 58464 15864
rect 58306 15276 58312 15852
rect 58346 15276 58424 15852
rect 58458 15276 58464 15852
rect 58306 15264 58464 15276
rect 58546 15852 58704 15864
rect 58546 15276 58552 15852
rect 58586 15276 58664 15852
rect 58698 15276 58704 15852
rect 58546 15264 58704 15276
rect 58786 15852 58944 15864
rect 58786 15276 58792 15852
rect 58826 15276 58904 15852
rect 58938 15276 58944 15852
rect 58786 15264 58944 15276
rect 59026 15852 59184 15864
rect 59026 15276 59032 15852
rect 59066 15276 59144 15852
rect 59178 15276 59184 15852
rect 59026 15264 59184 15276
rect 59266 15852 59424 15864
rect 59266 15276 59272 15852
rect 59306 15276 59384 15852
rect 59418 15276 59424 15852
rect 59266 15264 59424 15276
rect 59506 15852 59664 15864
rect 59506 15276 59512 15852
rect 59546 15276 59624 15852
rect 59658 15276 59664 15852
rect 59506 15264 59664 15276
rect 59746 15852 59904 15864
rect 59746 15276 59752 15852
rect 59786 15276 59864 15852
rect 59898 15276 59904 15852
rect 59746 15264 59904 15276
rect 59986 15852 60144 15864
rect 59986 15276 59992 15852
rect 60026 15276 60104 15852
rect 60138 15276 60144 15852
rect 59986 15264 60144 15276
rect 60226 15852 60384 15864
rect 60226 15276 60232 15852
rect 60266 15276 60344 15852
rect 60378 15276 60384 15852
rect 60226 15264 60384 15276
rect 60466 15852 60624 15864
rect 60466 15276 60472 15852
rect 60506 15276 60584 15852
rect 60618 15276 60624 15852
rect 60466 15264 60624 15276
rect 60706 15852 60864 15864
rect 60706 15276 60712 15852
rect 60746 15276 60824 15852
rect 60858 15276 60864 15852
rect 60706 15264 60864 15276
rect 60946 15852 61104 15864
rect 60946 15276 60952 15852
rect 60986 15276 61064 15852
rect 61098 15276 61104 15852
rect 60946 15264 61104 15276
rect 61186 15852 61344 15864
rect 61186 15276 61192 15852
rect 61226 15276 61304 15852
rect 61338 15276 61344 15852
rect 61186 15264 61344 15276
rect 61426 15852 61584 15864
rect 61426 15276 61432 15852
rect 61466 15276 61544 15852
rect 61578 15276 61584 15852
rect 61426 15264 61584 15276
rect 61666 15852 61824 15864
rect 61666 15276 61672 15852
rect 61706 15276 61784 15852
rect 61818 15276 61824 15852
rect 61666 15264 61824 15276
rect 61906 15852 62064 15864
rect 61906 15276 61912 15852
rect 61946 15276 62024 15852
rect 62058 15276 62064 15852
rect 61906 15264 62064 15276
rect 62146 15852 62264 15864
rect 62146 15276 62152 15852
rect 62186 15276 62264 15852
rect 62146 15264 62264 15276
rect 52586 14398 52652 15264
rect 52710 15226 52780 15232
rect 52950 15226 53020 15232
rect 52700 15094 52710 15226
rect 52780 15094 52790 15226
rect 52940 15094 52950 15226
rect 53020 15094 53030 15226
rect 52710 15088 52780 15094
rect 52950 15088 53020 15094
rect 53078 14398 53132 15264
rect 53190 15226 53260 15232
rect 53430 15226 53500 15232
rect 53180 15094 53190 15226
rect 53260 15094 53270 15226
rect 53420 15094 53430 15226
rect 53500 15094 53510 15226
rect 53190 15088 53260 15094
rect 53430 15088 53500 15094
rect 53558 14398 53612 15264
rect 53670 15226 53740 15232
rect 53910 15226 53980 15232
rect 53660 15094 53670 15226
rect 53740 15094 53750 15226
rect 53900 15094 53910 15226
rect 53980 15094 53990 15226
rect 53670 15088 53740 15094
rect 53910 15088 53980 15094
rect 54038 14398 54092 15264
rect 54150 15226 54220 15232
rect 54390 15226 54460 15232
rect 54140 15094 54150 15226
rect 54220 15094 54230 15226
rect 54380 15094 54390 15226
rect 54460 15094 54470 15226
rect 54150 15088 54220 15094
rect 54390 15088 54460 15094
rect 54518 14398 54572 15264
rect 54630 15226 54700 15232
rect 54870 15226 54940 15232
rect 54620 15094 54630 15226
rect 54700 15094 54710 15226
rect 54860 15094 54870 15226
rect 54940 15094 54950 15226
rect 54630 15088 54700 15094
rect 54870 15088 54940 15094
rect 54998 14398 55052 15264
rect 55110 15226 55180 15232
rect 55350 15226 55420 15232
rect 55100 15094 55110 15226
rect 55180 15094 55190 15226
rect 55340 15094 55350 15226
rect 55420 15094 55430 15226
rect 55110 15088 55180 15094
rect 55350 15088 55420 15094
rect 55478 14398 55532 15264
rect 55590 15226 55660 15232
rect 55830 15226 55900 15232
rect 55580 15094 55590 15226
rect 55660 15094 55670 15226
rect 55820 15094 55830 15226
rect 55900 15094 55910 15226
rect 55590 15088 55660 15094
rect 55830 15088 55900 15094
rect 55958 14398 56012 15264
rect 56070 15226 56140 15232
rect 56310 15226 56380 15232
rect 56060 15094 56070 15226
rect 56140 15094 56150 15226
rect 56300 15094 56310 15226
rect 56380 15094 56390 15226
rect 56070 15088 56140 15094
rect 56310 15088 56380 15094
rect 56438 14398 56492 15264
rect 56550 15226 56620 15232
rect 56790 15226 56860 15232
rect 56540 15094 56550 15226
rect 56620 15094 56630 15226
rect 56780 15094 56790 15226
rect 56860 15094 56870 15226
rect 56550 15088 56620 15094
rect 56790 15088 56860 15094
rect 56918 14398 56972 15264
rect 57030 15226 57100 15232
rect 57270 15226 57340 15232
rect 57020 15094 57030 15226
rect 57100 15094 57110 15226
rect 57260 15094 57270 15226
rect 57340 15094 57350 15226
rect 57030 15088 57100 15094
rect 57270 15088 57340 15094
rect 57398 14398 57452 15264
rect 57510 15226 57580 15232
rect 57750 15226 57820 15232
rect 57500 15094 57510 15226
rect 57580 15094 57590 15226
rect 57740 15094 57750 15226
rect 57820 15094 57830 15226
rect 57510 15088 57580 15094
rect 57750 15088 57820 15094
rect 57878 14398 57932 15264
rect 57990 15226 58060 15232
rect 58230 15226 58300 15232
rect 57980 15094 57990 15226
rect 58060 15094 58070 15226
rect 58220 15094 58230 15226
rect 58300 15094 58310 15226
rect 57990 15088 58060 15094
rect 58230 15088 58300 15094
rect 58358 14398 58412 15264
rect 58470 15226 58540 15232
rect 58710 15226 58780 15232
rect 58460 15094 58470 15226
rect 58540 15094 58550 15226
rect 58700 15094 58710 15226
rect 58780 15094 58790 15226
rect 58470 15088 58540 15094
rect 58710 15088 58780 15094
rect 58838 14398 58892 15264
rect 58950 15226 59020 15232
rect 59190 15226 59260 15232
rect 58940 15094 58950 15226
rect 59020 15094 59030 15226
rect 59180 15094 59190 15226
rect 59260 15094 59270 15226
rect 58950 15088 59020 15094
rect 59190 15088 59260 15094
rect 59318 14398 59372 15264
rect 59430 15226 59500 15232
rect 59670 15226 59740 15232
rect 59420 15094 59430 15226
rect 59500 15094 59510 15226
rect 59660 15094 59670 15226
rect 59740 15094 59750 15226
rect 59430 15088 59500 15094
rect 59670 15088 59740 15094
rect 59798 14398 59852 15264
rect 59910 15226 59980 15232
rect 60150 15226 60220 15232
rect 59900 15094 59910 15226
rect 59980 15094 59990 15226
rect 60140 15094 60150 15226
rect 60220 15094 60230 15226
rect 59910 15088 59980 15094
rect 60150 15088 60220 15094
rect 60278 14398 60332 15264
rect 60390 15226 60460 15232
rect 60630 15226 60700 15232
rect 60380 15094 60390 15226
rect 60460 15094 60470 15226
rect 60620 15094 60630 15226
rect 60700 15094 60710 15226
rect 60390 15088 60460 15094
rect 60630 15088 60700 15094
rect 60758 14398 60812 15264
rect 60870 15226 60940 15232
rect 61110 15226 61180 15232
rect 60860 15094 60870 15226
rect 60940 15094 60950 15226
rect 61100 15094 61110 15226
rect 61180 15094 61190 15226
rect 60870 15088 60940 15094
rect 61110 15088 61180 15094
rect 61238 14398 61292 15264
rect 61350 15226 61420 15232
rect 61590 15226 61660 15232
rect 61340 15094 61350 15226
rect 61420 15094 61430 15226
rect 61580 15094 61590 15226
rect 61660 15094 61670 15226
rect 61350 15088 61420 15094
rect 61590 15088 61660 15094
rect 61718 14398 61772 15264
rect 61830 15226 61900 15232
rect 62070 15226 62140 15232
rect 61820 15094 61830 15226
rect 61900 15094 61910 15226
rect 62060 15094 62070 15226
rect 62140 15094 62150 15226
rect 61830 15088 61900 15094
rect 62070 15088 62140 15094
rect 62198 14398 62264 15264
rect 43270 13536 71578 14398
rect 43270 12598 43348 13536
rect 43410 12679 43802 12685
rect 43410 12645 43422 12679
rect 43790 12645 43802 12679
rect 43410 12639 43802 12645
rect 43998 12679 44390 12685
rect 43998 12645 44010 12679
rect 44378 12645 44390 12679
rect 43998 12639 44390 12645
rect 44452 12598 44524 13536
rect 44586 12679 44978 12685
rect 44586 12645 44598 12679
rect 44966 12645 44978 12679
rect 44586 12639 44978 12645
rect 45174 12679 45566 12685
rect 45174 12645 45186 12679
rect 45554 12645 45566 12679
rect 45174 12639 45566 12645
rect 45628 12598 45700 13536
rect 45762 12679 46154 12685
rect 45762 12645 45774 12679
rect 46142 12645 46154 12679
rect 45762 12639 46154 12645
rect 46350 12679 46742 12685
rect 46350 12645 46362 12679
rect 46730 12645 46742 12679
rect 46350 12639 46742 12645
rect 46804 12598 46876 13536
rect 46938 12679 47330 12685
rect 46938 12645 46950 12679
rect 47318 12645 47330 12679
rect 46938 12639 47330 12645
rect 47526 12679 47918 12685
rect 47526 12645 47538 12679
rect 47906 12645 47918 12679
rect 47526 12639 47918 12645
rect 47980 12598 48052 13536
rect 48114 12679 48506 12685
rect 48114 12645 48126 12679
rect 48494 12645 48506 12679
rect 48114 12639 48506 12645
rect 48702 12679 49094 12685
rect 48702 12645 48714 12679
rect 49082 12645 49094 12679
rect 48702 12639 49094 12645
rect 49156 12598 49228 13536
rect 49290 12679 49682 12685
rect 49290 12645 49302 12679
rect 49670 12645 49682 12679
rect 49290 12639 49682 12645
rect 49878 12679 50270 12685
rect 49878 12645 49890 12679
rect 50258 12645 50270 12679
rect 49878 12639 50270 12645
rect 50332 12598 50404 13536
rect 50466 12679 50858 12685
rect 50466 12645 50478 12679
rect 50846 12645 50858 12679
rect 50466 12639 50858 12645
rect 51054 12679 51446 12685
rect 51054 12645 51066 12679
rect 51434 12645 51446 12679
rect 51054 12639 51446 12645
rect 51508 12598 51580 13536
rect 51642 12679 52034 12685
rect 51642 12645 51654 12679
rect 52022 12645 52034 12679
rect 51642 12639 52034 12645
rect 52230 12679 52622 12685
rect 52230 12645 52242 12679
rect 52610 12645 52622 12679
rect 52230 12639 52622 12645
rect 52684 12598 52756 13536
rect 52818 12679 53210 12685
rect 52818 12645 52830 12679
rect 53198 12645 53210 12679
rect 52818 12639 53210 12645
rect 53406 12679 53798 12685
rect 53406 12645 53418 12679
rect 53786 12645 53798 12679
rect 53406 12639 53798 12645
rect 53860 12598 53932 13536
rect 53994 12679 54386 12685
rect 53994 12645 54006 12679
rect 54374 12645 54386 12679
rect 53994 12639 54386 12645
rect 54582 12679 54974 12685
rect 54582 12645 54594 12679
rect 54962 12645 54974 12679
rect 54582 12639 54974 12645
rect 55008 12598 55080 13536
rect 55170 12679 55562 12685
rect 55170 12645 55182 12679
rect 55550 12645 55562 12679
rect 55170 12639 55562 12645
rect 55758 12679 56150 12685
rect 55758 12645 55770 12679
rect 56138 12645 56150 12679
rect 55758 12639 56150 12645
rect 56346 12679 56738 12685
rect 56346 12645 56358 12679
rect 56726 12645 56738 12679
rect 56346 12639 56738 12645
rect 56934 12679 57326 12685
rect 56934 12645 56946 12679
rect 57314 12645 57326 12679
rect 56934 12639 57326 12645
rect 57522 12679 57914 12685
rect 57522 12645 57534 12679
rect 57902 12645 57914 12679
rect 57522 12639 57914 12645
rect 58110 12679 58502 12685
rect 58110 12645 58122 12679
rect 58490 12645 58502 12679
rect 58110 12639 58502 12645
rect 58698 12679 59090 12685
rect 58698 12645 58710 12679
rect 59078 12645 59090 12679
rect 58698 12639 59090 12645
rect 59286 12679 59678 12685
rect 59286 12645 59298 12679
rect 59666 12645 59678 12679
rect 59286 12639 59678 12645
rect 59768 12598 59840 13536
rect 59874 12679 60266 12685
rect 59874 12645 59886 12679
rect 60254 12645 60266 12679
rect 59874 12639 60266 12645
rect 60462 12679 60854 12685
rect 60462 12645 60474 12679
rect 60842 12645 60854 12679
rect 60462 12639 60854 12645
rect 60916 12598 60988 13536
rect 61050 12679 61442 12685
rect 61050 12645 61062 12679
rect 61430 12645 61442 12679
rect 61050 12639 61442 12645
rect 61638 12679 62030 12685
rect 61638 12645 61650 12679
rect 62018 12645 62030 12679
rect 61638 12639 62030 12645
rect 62092 12598 62164 13536
rect 62226 12679 62618 12685
rect 62226 12645 62238 12679
rect 62606 12645 62618 12679
rect 62226 12639 62618 12645
rect 62814 12679 63206 12685
rect 62814 12645 62826 12679
rect 63194 12645 63206 12679
rect 62814 12639 63206 12645
rect 63268 12598 63340 13536
rect 63402 12679 63794 12685
rect 63402 12645 63414 12679
rect 63782 12645 63794 12679
rect 63402 12639 63794 12645
rect 63990 12679 64382 12685
rect 63990 12645 64002 12679
rect 64370 12645 64382 12679
rect 63990 12639 64382 12645
rect 64444 12598 64516 13536
rect 64578 12679 64970 12685
rect 64578 12645 64590 12679
rect 64958 12645 64970 12679
rect 64578 12639 64970 12645
rect 65166 12679 65558 12685
rect 65166 12645 65178 12679
rect 65546 12645 65558 12679
rect 65166 12639 65558 12645
rect 65620 12598 65692 13536
rect 65754 12679 66146 12685
rect 65754 12645 65766 12679
rect 66134 12645 66146 12679
rect 65754 12639 66146 12645
rect 66342 12679 66734 12685
rect 66342 12645 66354 12679
rect 66722 12645 66734 12679
rect 66342 12639 66734 12645
rect 66796 12598 66868 13536
rect 66930 12679 67322 12685
rect 66930 12645 66942 12679
rect 67310 12645 67322 12679
rect 66930 12639 67322 12645
rect 67518 12679 67910 12685
rect 67518 12645 67530 12679
rect 67898 12645 67910 12679
rect 67518 12639 67910 12645
rect 67972 12598 68044 13536
rect 68106 12679 68498 12685
rect 68106 12645 68118 12679
rect 68486 12645 68498 12679
rect 68106 12639 68498 12645
rect 68694 12679 69086 12685
rect 68694 12645 68706 12679
rect 69074 12645 69086 12679
rect 68694 12639 69086 12645
rect 69148 12598 69220 13536
rect 69282 12679 69674 12685
rect 69282 12645 69294 12679
rect 69662 12645 69674 12679
rect 69282 12639 69674 12645
rect 69870 12679 70262 12685
rect 69870 12645 69882 12679
rect 70250 12645 70262 12679
rect 69870 12639 70262 12645
rect 70324 12598 70396 13536
rect 70458 12679 70850 12685
rect 70458 12645 70470 12679
rect 70838 12645 70850 12679
rect 70458 12639 70850 12645
rect 71046 12679 71438 12685
rect 71046 12645 71058 12679
rect 71426 12645 71438 12679
rect 71046 12639 71438 12645
rect 71500 12598 71578 13536
rect 43270 12586 43400 12598
rect 43270 11810 43360 12586
rect 43394 11810 43400 12586
rect 43270 11798 43400 11810
rect 43812 12586 43988 12598
rect 43812 11810 43818 12586
rect 43852 11810 43948 12586
rect 43982 11810 43988 12586
rect 43812 11798 43988 11810
rect 44400 12586 44576 12598
rect 44400 11810 44406 12586
rect 44440 11810 44536 12586
rect 44570 11810 44576 12586
rect 44400 11798 44576 11810
rect 44988 12586 45164 12598
rect 44988 11810 44994 12586
rect 45028 11810 45124 12586
rect 45158 11810 45164 12586
rect 44988 11798 45164 11810
rect 45576 12586 45752 12598
rect 45576 11810 45582 12586
rect 45616 11810 45712 12586
rect 45746 11810 45752 12586
rect 45576 11798 45752 11810
rect 46164 12586 46340 12598
rect 46164 11810 46170 12586
rect 46204 11810 46300 12586
rect 46334 11810 46340 12586
rect 46164 11798 46340 11810
rect 46752 12586 46928 12598
rect 46752 11810 46758 12586
rect 46792 11810 46888 12586
rect 46922 11810 46928 12586
rect 46752 11798 46928 11810
rect 47340 12586 47516 12598
rect 47340 11810 47346 12586
rect 47380 11810 47476 12586
rect 47510 11810 47516 12586
rect 47340 11798 47516 11810
rect 47928 12586 48104 12598
rect 47928 11810 47934 12586
rect 47968 11810 48064 12586
rect 48098 11810 48104 12586
rect 47928 11798 48104 11810
rect 48516 12586 48692 12598
rect 48516 11810 48522 12586
rect 48556 11810 48652 12586
rect 48686 11810 48692 12586
rect 48516 11798 48692 11810
rect 49104 12586 49280 12598
rect 49104 11810 49110 12586
rect 49144 11810 49240 12586
rect 49274 11810 49280 12586
rect 49104 11798 49280 11810
rect 49692 12586 49868 12598
rect 49692 11810 49698 12586
rect 49732 11810 49828 12586
rect 49862 11810 49868 12586
rect 49692 11798 49868 11810
rect 50280 12586 50456 12598
rect 50280 11810 50286 12586
rect 50320 11810 50416 12586
rect 50450 11810 50456 12586
rect 50280 11798 50456 11810
rect 50868 12586 51044 12598
rect 50868 11810 50874 12586
rect 50908 11810 51004 12586
rect 51038 11810 51044 12586
rect 50868 11798 51044 11810
rect 51456 12586 51632 12598
rect 51456 11810 51462 12586
rect 51496 11810 51592 12586
rect 51626 11810 51632 12586
rect 51456 11798 51632 11810
rect 52044 12586 52220 12598
rect 52044 11810 52050 12586
rect 52084 11810 52180 12586
rect 52214 11810 52220 12586
rect 52044 11798 52220 11810
rect 52632 12586 52808 12598
rect 52632 11810 52638 12586
rect 52672 11810 52768 12586
rect 52802 11810 52808 12586
rect 52632 11798 52808 11810
rect 53220 12586 53396 12598
rect 53220 11810 53226 12586
rect 53260 11810 53356 12586
rect 53390 11810 53396 12586
rect 53220 11798 53396 11810
rect 53808 12586 53984 12598
rect 53808 11810 53814 12586
rect 53848 11810 53944 12586
rect 53978 11810 53984 12586
rect 53808 11798 53984 11810
rect 54396 12586 54572 12598
rect 54396 11810 54402 12586
rect 54436 11810 54532 12586
rect 54566 11810 54572 12586
rect 54396 11798 54572 11810
rect 54984 12586 55080 12598
rect 54984 11810 54990 12586
rect 55024 11862 55080 12586
rect 55114 12586 55160 12598
rect 55024 11810 55082 11862
rect 54984 11798 55082 11810
rect 55114 11810 55120 12586
rect 55154 11810 55160 12586
rect 55114 11798 55160 11810
rect 55572 12586 55748 12598
rect 55572 11810 55578 12586
rect 55612 11810 55708 12586
rect 55742 11810 55748 12586
rect 55572 11798 55748 11810
rect 56160 12586 56336 12598
rect 56160 11810 56166 12586
rect 56200 11810 56296 12586
rect 56330 11810 56336 12586
rect 56160 11798 56336 11810
rect 56748 12586 56924 12598
rect 56748 11810 56754 12586
rect 56788 11810 56884 12586
rect 56918 11810 56924 12586
rect 56748 11798 56924 11810
rect 57336 12586 57382 12598
rect 57336 11810 57342 12586
rect 57376 11810 57382 12586
rect 57336 11798 57382 11810
rect 57466 12586 57512 12598
rect 57466 11810 57472 12586
rect 57506 11810 57512 12586
rect 57466 11798 57512 11810
rect 57924 12586 58100 12598
rect 57924 11810 57930 12586
rect 57964 11810 58060 12586
rect 58094 11810 58100 12586
rect 57924 11798 58100 11810
rect 58512 12586 58688 12598
rect 58512 11810 58518 12586
rect 58552 11810 58648 12586
rect 58682 11810 58688 12586
rect 58512 11798 58688 11810
rect 59100 12586 59276 12598
rect 59100 11810 59106 12586
rect 59140 11810 59236 12586
rect 59270 11810 59276 12586
rect 59100 11798 59276 11810
rect 59688 12586 59734 12598
rect 59688 11810 59694 12586
rect 59728 11810 59734 12586
rect 59688 11798 59734 11810
rect 59768 12586 59864 12598
rect 59768 11810 59824 12586
rect 59858 11810 59864 12586
rect 59768 11798 59864 11810
rect 60276 12586 60452 12598
rect 60276 11810 60282 12586
rect 60316 11810 60412 12586
rect 60446 11810 60452 12586
rect 60276 11798 60452 11810
rect 60864 12586 61040 12598
rect 60864 11810 60870 12586
rect 60904 11810 61000 12586
rect 61034 11810 61040 12586
rect 60864 11798 61040 11810
rect 61452 12586 61628 12598
rect 61452 11810 61458 12586
rect 61492 11810 61588 12586
rect 61622 11810 61628 12586
rect 61452 11798 61628 11810
rect 62040 12586 62216 12598
rect 62040 11810 62046 12586
rect 62080 11810 62176 12586
rect 62210 11810 62216 12586
rect 62040 11798 62216 11810
rect 62628 12586 62804 12598
rect 62628 11810 62634 12586
rect 62668 11810 62764 12586
rect 62798 11810 62804 12586
rect 62628 11798 62804 11810
rect 63216 12586 63392 12598
rect 63216 11810 63222 12586
rect 63256 11810 63352 12586
rect 63386 11810 63392 12586
rect 63216 11798 63392 11810
rect 63804 12586 63980 12598
rect 63804 11810 63810 12586
rect 63844 11810 63940 12586
rect 63974 11810 63980 12586
rect 63804 11798 63980 11810
rect 64392 12586 64568 12598
rect 64392 11810 64398 12586
rect 64432 11810 64528 12586
rect 64562 11810 64568 12586
rect 64392 11798 64568 11810
rect 64980 12586 65156 12598
rect 64980 11810 64986 12586
rect 65020 11810 65116 12586
rect 65150 11810 65156 12586
rect 64980 11798 65156 11810
rect 65568 12586 65744 12598
rect 65568 11810 65574 12586
rect 65608 11810 65704 12586
rect 65738 11810 65744 12586
rect 65568 11798 65744 11810
rect 66156 12586 66332 12598
rect 66156 11810 66162 12586
rect 66196 11810 66292 12586
rect 66326 11810 66332 12586
rect 66156 11798 66332 11810
rect 66744 12586 66920 12598
rect 66744 11810 66750 12586
rect 66784 11810 66880 12586
rect 66914 11810 66920 12586
rect 66744 11798 66920 11810
rect 67332 12586 67508 12598
rect 67332 11810 67338 12586
rect 67372 11810 67468 12586
rect 67502 11810 67508 12586
rect 67332 11798 67508 11810
rect 67920 12586 68096 12598
rect 67920 11810 67926 12586
rect 67960 11810 68056 12586
rect 68090 11810 68096 12586
rect 67920 11798 68096 11810
rect 68508 12586 68684 12598
rect 68508 11810 68514 12586
rect 68548 11810 68644 12586
rect 68678 11810 68684 12586
rect 68508 11798 68684 11810
rect 69096 12586 69272 12598
rect 69096 11810 69102 12586
rect 69136 11810 69232 12586
rect 69266 11810 69272 12586
rect 69096 11798 69272 11810
rect 69684 12586 69860 12598
rect 69684 11810 69690 12586
rect 69724 11810 69820 12586
rect 69854 11810 69860 12586
rect 69684 11798 69860 11810
rect 70272 12586 70448 12598
rect 70272 11810 70278 12586
rect 70312 11810 70408 12586
rect 70442 11810 70448 12586
rect 70272 11798 70448 11810
rect 70860 12586 71036 12598
rect 70860 11810 70866 12586
rect 70900 11810 70996 12586
rect 71030 11810 71036 12586
rect 70860 11798 71036 11810
rect 71448 12586 71578 12598
rect 71448 11810 71454 12586
rect 71488 11810 71578 12586
rect 71448 11798 71578 11810
rect 43270 11598 43354 11798
rect 43410 11751 43802 11757
rect 43410 11717 43422 11751
rect 43790 11717 43802 11751
rect 43410 11679 43802 11717
rect 43410 11645 43422 11679
rect 43790 11645 43802 11679
rect 43410 11639 43802 11645
rect 43858 11598 43942 11798
rect 43998 11751 44390 11757
rect 43998 11717 44010 11751
rect 44378 11717 44390 11751
rect 43998 11679 44390 11717
rect 43998 11645 44010 11679
rect 44378 11645 44390 11679
rect 43998 11639 44390 11645
rect 44446 11598 44530 11798
rect 44586 11751 44978 11757
rect 44586 11717 44598 11751
rect 44966 11717 44978 11751
rect 44586 11679 44978 11717
rect 44586 11645 44598 11679
rect 44966 11645 44978 11679
rect 44586 11639 44978 11645
rect 45034 11598 45118 11798
rect 45174 11751 45566 11757
rect 45174 11717 45186 11751
rect 45554 11717 45566 11751
rect 45174 11679 45566 11717
rect 45174 11645 45186 11679
rect 45554 11645 45566 11679
rect 45174 11639 45566 11645
rect 45622 11598 45706 11798
rect 45762 11751 46154 11757
rect 45762 11717 45774 11751
rect 46142 11717 46154 11751
rect 45762 11679 46154 11717
rect 45762 11645 45774 11679
rect 46142 11645 46154 11679
rect 45762 11639 46154 11645
rect 46210 11598 46294 11798
rect 46350 11751 46742 11757
rect 46350 11717 46362 11751
rect 46730 11717 46742 11751
rect 46350 11679 46742 11717
rect 46350 11645 46362 11679
rect 46730 11645 46742 11679
rect 46350 11639 46742 11645
rect 46798 11598 46882 11798
rect 46938 11751 47330 11757
rect 46938 11717 46950 11751
rect 47318 11717 47330 11751
rect 46938 11679 47330 11717
rect 46938 11645 46950 11679
rect 47318 11645 47330 11679
rect 46938 11639 47330 11645
rect 47386 11598 47470 11798
rect 47526 11751 47918 11757
rect 47526 11717 47538 11751
rect 47906 11717 47918 11751
rect 47526 11679 47918 11717
rect 47526 11645 47538 11679
rect 47906 11645 47918 11679
rect 47526 11639 47918 11645
rect 47974 11598 48058 11798
rect 48114 11751 48506 11757
rect 48114 11717 48126 11751
rect 48494 11717 48506 11751
rect 48114 11679 48506 11717
rect 48114 11645 48126 11679
rect 48494 11645 48506 11679
rect 48114 11639 48506 11645
rect 48562 11598 48646 11798
rect 48702 11751 49094 11757
rect 48702 11717 48714 11751
rect 49082 11717 49094 11751
rect 48702 11679 49094 11717
rect 48702 11645 48714 11679
rect 49082 11645 49094 11679
rect 48702 11639 49094 11645
rect 49150 11598 49234 11798
rect 49290 11751 49682 11757
rect 49290 11717 49302 11751
rect 49670 11717 49682 11751
rect 49290 11679 49682 11717
rect 49290 11645 49302 11679
rect 49670 11645 49682 11679
rect 49290 11639 49682 11645
rect 49738 11598 49822 11798
rect 49878 11751 50270 11757
rect 49878 11717 49890 11751
rect 50258 11717 50270 11751
rect 49878 11679 50270 11717
rect 49878 11645 49890 11679
rect 50258 11645 50270 11679
rect 49878 11639 50270 11645
rect 50326 11598 50410 11798
rect 50466 11751 50858 11757
rect 50466 11717 50478 11751
rect 50846 11717 50858 11751
rect 50466 11679 50858 11717
rect 50466 11645 50478 11679
rect 50846 11645 50858 11679
rect 50466 11639 50858 11645
rect 50914 11598 50998 11798
rect 51054 11751 51446 11757
rect 51054 11717 51066 11751
rect 51434 11717 51446 11751
rect 51054 11679 51446 11717
rect 51054 11645 51066 11679
rect 51434 11645 51446 11679
rect 51054 11639 51446 11645
rect 51502 11598 51586 11798
rect 51642 11751 52034 11757
rect 51642 11717 51654 11751
rect 52022 11717 52034 11751
rect 51642 11679 52034 11717
rect 51642 11645 51654 11679
rect 52022 11645 52034 11679
rect 51642 11639 52034 11645
rect 52090 11598 52174 11798
rect 52230 11751 52622 11757
rect 52230 11717 52242 11751
rect 52610 11717 52622 11751
rect 52230 11679 52622 11717
rect 52230 11645 52242 11679
rect 52610 11645 52622 11679
rect 52230 11639 52622 11645
rect 52678 11598 52762 11798
rect 52818 11751 53210 11757
rect 52818 11717 52830 11751
rect 53198 11717 53210 11751
rect 52818 11679 53210 11717
rect 52818 11645 52830 11679
rect 53198 11645 53210 11679
rect 52818 11639 53210 11645
rect 53266 11598 53350 11798
rect 53406 11751 53798 11757
rect 53406 11717 53418 11751
rect 53786 11717 53798 11751
rect 53406 11679 53798 11717
rect 53406 11645 53418 11679
rect 53786 11645 53798 11679
rect 53406 11639 53798 11645
rect 53854 11598 53938 11798
rect 53994 11751 54386 11757
rect 53994 11717 54006 11751
rect 54374 11717 54386 11751
rect 53994 11679 54386 11717
rect 53994 11645 54006 11679
rect 54374 11645 54386 11679
rect 53994 11639 54386 11645
rect 54442 11598 54526 11798
rect 54582 11751 54974 11757
rect 54582 11717 54594 11751
rect 54962 11717 54974 11751
rect 54582 11679 54974 11717
rect 54582 11645 54594 11679
rect 54962 11645 54974 11679
rect 54582 11639 54974 11645
rect 55024 11598 55082 11798
rect 55170 11751 55562 11757
rect 55170 11717 55182 11751
rect 55550 11717 55562 11751
rect 55170 11679 55562 11717
rect 55170 11645 55182 11679
rect 55550 11645 55562 11679
rect 55170 11639 55562 11645
rect 55618 11598 55702 11798
rect 55758 11751 56150 11757
rect 55758 11717 55770 11751
rect 56138 11717 56150 11751
rect 55758 11679 56150 11717
rect 55758 11645 55770 11679
rect 56138 11645 56150 11679
rect 55758 11639 56150 11645
rect 56206 11598 56290 11798
rect 56346 11751 56738 11757
rect 56346 11717 56358 11751
rect 56726 11717 56738 11751
rect 56346 11679 56738 11717
rect 56346 11645 56358 11679
rect 56726 11645 56738 11679
rect 56346 11639 56738 11645
rect 56794 11598 56878 11798
rect 56934 11751 57326 11757
rect 56934 11717 56946 11751
rect 57314 11717 57326 11751
rect 56934 11679 57326 11717
rect 56934 11645 56946 11679
rect 57314 11645 57326 11679
rect 56934 11639 57326 11645
rect 57522 11751 57914 11757
rect 57522 11717 57534 11751
rect 57902 11717 57914 11751
rect 57522 11679 57914 11717
rect 57522 11645 57534 11679
rect 57902 11645 57914 11679
rect 57522 11639 57914 11645
rect 57970 11598 58054 11798
rect 58110 11751 58502 11757
rect 58110 11717 58122 11751
rect 58490 11717 58502 11751
rect 58110 11679 58502 11717
rect 58110 11645 58122 11679
rect 58490 11645 58502 11679
rect 58110 11639 58502 11645
rect 58558 11598 58642 11798
rect 58698 11751 59090 11757
rect 58698 11717 58710 11751
rect 59078 11717 59090 11751
rect 58698 11679 59090 11717
rect 58698 11645 58710 11679
rect 59078 11645 59090 11679
rect 58698 11639 59090 11645
rect 59146 11598 59230 11798
rect 59286 11751 59678 11757
rect 59286 11717 59298 11751
rect 59666 11717 59678 11751
rect 59286 11679 59678 11717
rect 59286 11645 59298 11679
rect 59666 11645 59678 11679
rect 59286 11639 59678 11645
rect 59768 11598 59824 11798
rect 59874 11751 60266 11757
rect 59874 11717 59886 11751
rect 60254 11717 60266 11751
rect 59874 11679 60266 11717
rect 59874 11645 59886 11679
rect 60254 11645 60266 11679
rect 59874 11639 60266 11645
rect 60322 11598 60406 11798
rect 60462 11751 60854 11757
rect 60462 11717 60474 11751
rect 60842 11717 60854 11751
rect 60462 11679 60854 11717
rect 60462 11645 60474 11679
rect 60842 11645 60854 11679
rect 60462 11639 60854 11645
rect 60910 11598 60994 11798
rect 61050 11751 61442 11757
rect 61050 11717 61062 11751
rect 61430 11717 61442 11751
rect 61050 11679 61442 11717
rect 61050 11645 61062 11679
rect 61430 11645 61442 11679
rect 61050 11639 61442 11645
rect 61498 11598 61582 11798
rect 61638 11751 62030 11757
rect 61638 11717 61650 11751
rect 62018 11717 62030 11751
rect 61638 11679 62030 11717
rect 61638 11645 61650 11679
rect 62018 11645 62030 11679
rect 61638 11639 62030 11645
rect 62086 11598 62170 11798
rect 62226 11751 62618 11757
rect 62226 11717 62238 11751
rect 62606 11717 62618 11751
rect 62226 11679 62618 11717
rect 62226 11645 62238 11679
rect 62606 11645 62618 11679
rect 62226 11639 62618 11645
rect 62674 11598 62758 11798
rect 62814 11751 63206 11757
rect 62814 11717 62826 11751
rect 63194 11717 63206 11751
rect 62814 11679 63206 11717
rect 62814 11645 62826 11679
rect 63194 11645 63206 11679
rect 62814 11639 63206 11645
rect 63262 11598 63346 11798
rect 63402 11751 63794 11757
rect 63402 11717 63414 11751
rect 63782 11717 63794 11751
rect 63402 11679 63794 11717
rect 63402 11645 63414 11679
rect 63782 11645 63794 11679
rect 63402 11639 63794 11645
rect 63850 11598 63934 11798
rect 63990 11751 64382 11757
rect 63990 11717 64002 11751
rect 64370 11717 64382 11751
rect 63990 11679 64382 11717
rect 63990 11645 64002 11679
rect 64370 11645 64382 11679
rect 63990 11639 64382 11645
rect 64438 11598 64522 11798
rect 64578 11751 64970 11757
rect 64578 11717 64590 11751
rect 64958 11717 64970 11751
rect 64578 11679 64970 11717
rect 64578 11645 64590 11679
rect 64958 11645 64970 11679
rect 64578 11639 64970 11645
rect 65026 11598 65110 11798
rect 65166 11751 65558 11757
rect 65166 11717 65178 11751
rect 65546 11717 65558 11751
rect 65166 11679 65558 11717
rect 65166 11645 65178 11679
rect 65546 11645 65558 11679
rect 65166 11639 65558 11645
rect 65614 11598 65698 11798
rect 65754 11751 66146 11757
rect 65754 11717 65766 11751
rect 66134 11717 66146 11751
rect 65754 11679 66146 11717
rect 65754 11645 65766 11679
rect 66134 11645 66146 11679
rect 65754 11639 66146 11645
rect 66202 11598 66286 11798
rect 66342 11751 66734 11757
rect 66342 11717 66354 11751
rect 66722 11717 66734 11751
rect 66342 11679 66734 11717
rect 66342 11645 66354 11679
rect 66722 11645 66734 11679
rect 66342 11639 66734 11645
rect 66790 11598 66874 11798
rect 66930 11751 67322 11757
rect 66930 11717 66942 11751
rect 67310 11717 67322 11751
rect 66930 11679 67322 11717
rect 66930 11645 66942 11679
rect 67310 11645 67322 11679
rect 66930 11639 67322 11645
rect 67378 11598 67462 11798
rect 67518 11751 67910 11757
rect 67518 11717 67530 11751
rect 67898 11717 67910 11751
rect 67518 11679 67910 11717
rect 67518 11645 67530 11679
rect 67898 11645 67910 11679
rect 67518 11639 67910 11645
rect 67966 11598 68050 11798
rect 68106 11751 68498 11757
rect 68106 11717 68118 11751
rect 68486 11717 68498 11751
rect 68106 11679 68498 11717
rect 68106 11645 68118 11679
rect 68486 11645 68498 11679
rect 68106 11639 68498 11645
rect 68554 11598 68638 11798
rect 68694 11751 69086 11757
rect 68694 11717 68706 11751
rect 69074 11717 69086 11751
rect 68694 11679 69086 11717
rect 68694 11645 68706 11679
rect 69074 11645 69086 11679
rect 68694 11639 69086 11645
rect 69142 11598 69226 11798
rect 69282 11751 69674 11757
rect 69282 11717 69294 11751
rect 69662 11717 69674 11751
rect 69282 11679 69674 11717
rect 69282 11645 69294 11679
rect 69662 11645 69674 11679
rect 69282 11639 69674 11645
rect 69730 11598 69814 11798
rect 69870 11751 70262 11757
rect 69870 11717 69882 11751
rect 70250 11717 70262 11751
rect 69870 11679 70262 11717
rect 69870 11645 69882 11679
rect 70250 11645 70262 11679
rect 69870 11639 70262 11645
rect 70318 11598 70402 11798
rect 70458 11751 70850 11757
rect 70458 11717 70470 11751
rect 70838 11717 70850 11751
rect 70458 11679 70850 11717
rect 70458 11645 70470 11679
rect 70838 11645 70850 11679
rect 70458 11639 70850 11645
rect 70906 11598 70990 11798
rect 71046 11751 71438 11757
rect 71046 11717 71058 11751
rect 71426 11717 71438 11751
rect 71046 11679 71438 11717
rect 71046 11645 71058 11679
rect 71426 11645 71438 11679
rect 71046 11639 71438 11645
rect 71494 11598 71578 11798
rect 43270 11586 43400 11598
rect 43270 10810 43360 11586
rect 43394 10810 43400 11586
rect 43270 10798 43400 10810
rect 43812 11586 43988 11598
rect 43812 10810 43818 11586
rect 43852 10810 43948 11586
rect 43982 10810 43988 11586
rect 43812 10798 43988 10810
rect 44400 11586 44576 11598
rect 44400 10810 44406 11586
rect 44440 10810 44536 11586
rect 44570 10810 44576 11586
rect 44400 10798 44576 10810
rect 44988 11586 45164 11598
rect 44988 10810 44994 11586
rect 45028 10810 45124 11586
rect 45158 10810 45164 11586
rect 44988 10798 45164 10810
rect 45576 11586 45752 11598
rect 45576 10810 45582 11586
rect 45616 10810 45712 11586
rect 45746 10810 45752 11586
rect 45576 10798 45752 10810
rect 46164 11586 46340 11598
rect 46164 10810 46170 11586
rect 46204 10810 46300 11586
rect 46334 10810 46340 11586
rect 46164 10798 46340 10810
rect 46752 11586 46928 11598
rect 46752 10810 46758 11586
rect 46792 10810 46888 11586
rect 46922 10810 46928 11586
rect 46752 10798 46928 10810
rect 47340 11586 47516 11598
rect 47340 10810 47346 11586
rect 47380 10810 47476 11586
rect 47510 10810 47516 11586
rect 47340 10798 47516 10810
rect 47928 11586 48104 11598
rect 47928 10810 47934 11586
rect 47968 10810 48064 11586
rect 48098 10810 48104 11586
rect 47928 10798 48104 10810
rect 48516 11586 48692 11598
rect 48516 10810 48522 11586
rect 48556 10810 48652 11586
rect 48686 10810 48692 11586
rect 48516 10798 48692 10810
rect 49104 11586 49280 11598
rect 49104 10810 49110 11586
rect 49144 10810 49240 11586
rect 49274 10810 49280 11586
rect 49104 10798 49280 10810
rect 49692 11586 49868 11598
rect 49692 10810 49698 11586
rect 49732 10810 49828 11586
rect 49862 10810 49868 11586
rect 49692 10798 49868 10810
rect 50280 11586 50456 11598
rect 50280 10810 50286 11586
rect 50320 10810 50416 11586
rect 50450 10810 50456 11586
rect 50280 10798 50456 10810
rect 50868 11586 51044 11598
rect 50868 10810 50874 11586
rect 50908 10810 51004 11586
rect 51038 10810 51044 11586
rect 50868 10798 51044 10810
rect 51456 11586 51632 11598
rect 51456 10810 51462 11586
rect 51496 10810 51592 11586
rect 51626 10810 51632 11586
rect 51456 10798 51632 10810
rect 52044 11586 52220 11598
rect 52044 10810 52050 11586
rect 52084 10810 52180 11586
rect 52214 10810 52220 11586
rect 52044 10798 52220 10810
rect 52632 11586 52808 11598
rect 52632 10810 52638 11586
rect 52672 10810 52768 11586
rect 52802 10810 52808 11586
rect 52632 10798 52808 10810
rect 53220 11586 53396 11598
rect 53220 10810 53226 11586
rect 53260 10810 53356 11586
rect 53390 10810 53396 11586
rect 53220 10798 53396 10810
rect 53808 11586 53984 11598
rect 53808 10810 53814 11586
rect 53848 10810 53944 11586
rect 53978 10810 53984 11586
rect 53808 10798 53984 10810
rect 54396 11586 54572 11598
rect 54396 10810 54402 11586
rect 54436 10810 54532 11586
rect 54566 10810 54572 11586
rect 54396 10798 54572 10810
rect 54984 11586 55082 11598
rect 54984 10810 54990 11586
rect 55024 10810 55082 11586
rect 54984 10798 55082 10810
rect 55114 11586 55160 11598
rect 55114 10810 55120 11586
rect 55154 10810 55160 11586
rect 55114 10798 55160 10810
rect 55572 11586 55748 11598
rect 55572 10810 55578 11586
rect 55612 10810 55708 11586
rect 55742 10810 55748 11586
rect 55572 10798 55748 10810
rect 56160 11586 56336 11598
rect 56160 10810 56166 11586
rect 56200 10810 56296 11586
rect 56330 10810 56336 11586
rect 56160 10798 56336 10810
rect 56748 11586 56924 11598
rect 56748 10810 56754 11586
rect 56788 10810 56884 11586
rect 56918 10810 56924 11586
rect 56748 10798 56924 10810
rect 57336 11586 57382 11598
rect 57336 10810 57342 11586
rect 57376 10810 57382 11586
rect 57336 10798 57382 10810
rect 57466 11586 57512 11598
rect 57466 10810 57472 11586
rect 57506 10810 57512 11586
rect 57466 10798 57512 10810
rect 57924 11586 58100 11598
rect 57924 10810 57930 11586
rect 57964 10810 58060 11586
rect 58094 10810 58100 11586
rect 57924 10798 58100 10810
rect 58512 11586 58688 11598
rect 58512 10810 58518 11586
rect 58552 10810 58648 11586
rect 58682 10810 58688 11586
rect 58512 10798 58688 10810
rect 59100 11586 59276 11598
rect 59100 10810 59106 11586
rect 59140 10810 59236 11586
rect 59270 10810 59276 11586
rect 59100 10798 59276 10810
rect 59688 11586 59734 11598
rect 59688 10810 59694 11586
rect 59728 10810 59734 11586
rect 59688 10798 59734 10810
rect 59768 11586 59864 11598
rect 59768 10810 59824 11586
rect 59858 10810 59864 11586
rect 59768 10798 59864 10810
rect 60276 11586 60452 11598
rect 60276 10810 60282 11586
rect 60316 10810 60412 11586
rect 60446 10810 60452 11586
rect 60276 10798 60452 10810
rect 60864 11586 61040 11598
rect 60864 10810 60870 11586
rect 60904 10810 61000 11586
rect 61034 10810 61040 11586
rect 60864 10798 61040 10810
rect 61452 11586 61628 11598
rect 61452 10810 61458 11586
rect 61492 10810 61588 11586
rect 61622 10810 61628 11586
rect 61452 10798 61628 10810
rect 62040 11586 62216 11598
rect 62040 10810 62046 11586
rect 62080 10810 62176 11586
rect 62210 10810 62216 11586
rect 62040 10798 62216 10810
rect 62628 11586 62804 11598
rect 62628 10810 62634 11586
rect 62668 10810 62764 11586
rect 62798 10810 62804 11586
rect 62628 10798 62804 10810
rect 63216 11586 63392 11598
rect 63216 10810 63222 11586
rect 63256 10810 63352 11586
rect 63386 10810 63392 11586
rect 63216 10798 63392 10810
rect 63804 11586 63980 11598
rect 63804 10810 63810 11586
rect 63844 10810 63940 11586
rect 63974 10810 63980 11586
rect 63804 10798 63980 10810
rect 64392 11586 64568 11598
rect 64392 10810 64398 11586
rect 64432 10810 64528 11586
rect 64562 10810 64568 11586
rect 64392 10798 64568 10810
rect 64980 11586 65156 11598
rect 64980 10810 64986 11586
rect 65020 10810 65116 11586
rect 65150 10810 65156 11586
rect 64980 10798 65156 10810
rect 65568 11586 65744 11598
rect 65568 10810 65574 11586
rect 65608 10810 65704 11586
rect 65738 10810 65744 11586
rect 65568 10798 65744 10810
rect 66156 11586 66332 11598
rect 66156 10810 66162 11586
rect 66196 10810 66292 11586
rect 66326 10810 66332 11586
rect 66156 10798 66332 10810
rect 66744 11586 66920 11598
rect 66744 10810 66750 11586
rect 66784 10810 66880 11586
rect 66914 10810 66920 11586
rect 66744 10798 66920 10810
rect 67332 11586 67508 11598
rect 67332 10810 67338 11586
rect 67372 10810 67468 11586
rect 67502 10810 67508 11586
rect 67332 10798 67508 10810
rect 67920 11586 68096 11598
rect 67920 10810 67926 11586
rect 67960 10810 68056 11586
rect 68090 10810 68096 11586
rect 67920 10798 68096 10810
rect 68508 11586 68684 11598
rect 68508 10810 68514 11586
rect 68548 10810 68644 11586
rect 68678 10810 68684 11586
rect 68508 10798 68684 10810
rect 69096 11586 69272 11598
rect 69096 10810 69102 11586
rect 69136 10810 69232 11586
rect 69266 10810 69272 11586
rect 69096 10798 69272 10810
rect 69684 11586 69860 11598
rect 69684 10810 69690 11586
rect 69724 10810 69820 11586
rect 69854 10810 69860 11586
rect 69684 10798 69860 10810
rect 70272 11586 70448 11598
rect 70272 10810 70278 11586
rect 70312 10810 70408 11586
rect 70442 10810 70448 11586
rect 70272 10798 70448 10810
rect 70860 11586 71036 11598
rect 70860 10810 70866 11586
rect 70900 10810 70996 11586
rect 71030 10810 71036 11586
rect 70860 10798 71036 10810
rect 71448 11586 71578 11598
rect 71448 10810 71454 11586
rect 71488 10810 71578 11586
rect 71448 10798 71578 10810
rect 43270 10598 43354 10798
rect 43410 10751 43802 10757
rect 43410 10717 43422 10751
rect 43790 10717 43802 10751
rect 43410 10679 43802 10717
rect 43410 10645 43422 10679
rect 43790 10645 43802 10679
rect 43410 10639 43802 10645
rect 43858 10598 43942 10798
rect 43998 10751 44390 10757
rect 43998 10717 44010 10751
rect 44378 10717 44390 10751
rect 43998 10679 44390 10717
rect 43998 10645 44010 10679
rect 44378 10645 44390 10679
rect 43998 10639 44390 10645
rect 44446 10598 44530 10798
rect 44586 10751 44978 10757
rect 44586 10717 44598 10751
rect 44966 10717 44978 10751
rect 44586 10679 44978 10717
rect 44586 10645 44598 10679
rect 44966 10645 44978 10679
rect 44586 10639 44978 10645
rect 45034 10598 45118 10798
rect 45174 10751 45566 10757
rect 45174 10717 45186 10751
rect 45554 10717 45566 10751
rect 45174 10679 45566 10717
rect 45174 10645 45186 10679
rect 45554 10645 45566 10679
rect 45174 10639 45566 10645
rect 45622 10598 45706 10798
rect 45762 10751 46154 10757
rect 45762 10717 45774 10751
rect 46142 10717 46154 10751
rect 45762 10679 46154 10717
rect 45762 10645 45774 10679
rect 46142 10645 46154 10679
rect 45762 10639 46154 10645
rect 46210 10598 46294 10798
rect 46350 10751 46742 10757
rect 46350 10717 46362 10751
rect 46730 10717 46742 10751
rect 46350 10679 46742 10717
rect 46350 10645 46362 10679
rect 46730 10645 46742 10679
rect 46350 10639 46742 10645
rect 46798 10598 46882 10798
rect 46938 10751 47330 10757
rect 46938 10717 46950 10751
rect 47318 10717 47330 10751
rect 46938 10679 47330 10717
rect 46938 10645 46950 10679
rect 47318 10645 47330 10679
rect 46938 10639 47330 10645
rect 47386 10598 47470 10798
rect 47526 10751 47918 10757
rect 47526 10717 47538 10751
rect 47906 10717 47918 10751
rect 47526 10679 47918 10717
rect 47526 10645 47538 10679
rect 47906 10645 47918 10679
rect 47526 10639 47918 10645
rect 47974 10598 48058 10798
rect 48114 10751 48506 10757
rect 48114 10717 48126 10751
rect 48494 10717 48506 10751
rect 48114 10679 48506 10717
rect 48114 10645 48126 10679
rect 48494 10645 48506 10679
rect 48114 10639 48506 10645
rect 48562 10598 48646 10798
rect 48702 10751 49094 10757
rect 48702 10717 48714 10751
rect 49082 10717 49094 10751
rect 48702 10679 49094 10717
rect 48702 10645 48714 10679
rect 49082 10645 49094 10679
rect 48702 10639 49094 10645
rect 49150 10598 49234 10798
rect 49290 10751 49682 10757
rect 49290 10717 49302 10751
rect 49670 10717 49682 10751
rect 49290 10679 49682 10717
rect 49290 10645 49302 10679
rect 49670 10645 49682 10679
rect 49290 10639 49682 10645
rect 49738 10598 49822 10798
rect 49878 10751 50270 10757
rect 49878 10717 49890 10751
rect 50258 10717 50270 10751
rect 49878 10679 50270 10717
rect 49878 10645 49890 10679
rect 50258 10645 50270 10679
rect 49878 10639 50270 10645
rect 50326 10598 50410 10798
rect 50466 10751 50858 10757
rect 50466 10717 50478 10751
rect 50846 10717 50858 10751
rect 50466 10679 50858 10717
rect 50466 10645 50478 10679
rect 50846 10645 50858 10679
rect 50466 10639 50858 10645
rect 50914 10598 50998 10798
rect 51054 10751 51446 10757
rect 51054 10717 51066 10751
rect 51434 10717 51446 10751
rect 51054 10679 51446 10717
rect 51054 10645 51066 10679
rect 51434 10645 51446 10679
rect 51054 10639 51446 10645
rect 51502 10598 51586 10798
rect 51642 10751 52034 10757
rect 51642 10717 51654 10751
rect 52022 10717 52034 10751
rect 51642 10679 52034 10717
rect 51642 10645 51654 10679
rect 52022 10645 52034 10679
rect 51642 10639 52034 10645
rect 52090 10598 52174 10798
rect 52230 10751 52622 10757
rect 52230 10717 52242 10751
rect 52610 10717 52622 10751
rect 52230 10679 52622 10717
rect 52230 10645 52242 10679
rect 52610 10645 52622 10679
rect 52230 10639 52622 10645
rect 52678 10598 52762 10798
rect 52818 10751 53210 10757
rect 52818 10717 52830 10751
rect 53198 10717 53210 10751
rect 52818 10679 53210 10717
rect 52818 10645 52830 10679
rect 53198 10645 53210 10679
rect 52818 10639 53210 10645
rect 53266 10598 53350 10798
rect 53406 10751 53798 10757
rect 53406 10717 53418 10751
rect 53786 10717 53798 10751
rect 53406 10679 53798 10717
rect 53406 10645 53418 10679
rect 53786 10645 53798 10679
rect 53406 10639 53798 10645
rect 53854 10598 53938 10798
rect 53994 10751 54386 10757
rect 53994 10717 54006 10751
rect 54374 10717 54386 10751
rect 53994 10679 54386 10717
rect 53994 10645 54006 10679
rect 54374 10645 54386 10679
rect 53994 10639 54386 10645
rect 54442 10598 54526 10798
rect 54582 10751 54974 10757
rect 54582 10717 54594 10751
rect 54962 10717 54974 10751
rect 54582 10679 54974 10717
rect 54582 10645 54594 10679
rect 54962 10645 54974 10679
rect 54582 10639 54974 10645
rect 55024 10598 55082 10798
rect 55170 10751 55562 10757
rect 55170 10717 55182 10751
rect 55550 10717 55562 10751
rect 55170 10679 55562 10717
rect 55170 10645 55182 10679
rect 55550 10645 55562 10679
rect 55170 10639 55562 10645
rect 55618 10598 55702 10798
rect 55758 10751 56150 10757
rect 55758 10717 55770 10751
rect 56138 10717 56150 10751
rect 55758 10679 56150 10717
rect 55758 10645 55770 10679
rect 56138 10645 56150 10679
rect 55758 10639 56150 10645
rect 56206 10598 56290 10798
rect 56346 10751 56738 10757
rect 56346 10717 56358 10751
rect 56726 10717 56738 10751
rect 56346 10679 56738 10717
rect 56346 10645 56358 10679
rect 56726 10645 56738 10679
rect 56346 10639 56738 10645
rect 56794 10598 56878 10798
rect 56934 10751 57326 10757
rect 56934 10717 56946 10751
rect 57314 10717 57326 10751
rect 56934 10679 57326 10717
rect 56934 10645 56946 10679
rect 57314 10645 57326 10679
rect 56934 10639 57326 10645
rect 57522 10751 57914 10757
rect 57522 10717 57534 10751
rect 57902 10717 57914 10751
rect 57522 10679 57914 10717
rect 57522 10645 57534 10679
rect 57902 10645 57914 10679
rect 57522 10639 57914 10645
rect 57970 10598 58054 10798
rect 58110 10751 58502 10757
rect 58110 10717 58122 10751
rect 58490 10717 58502 10751
rect 58110 10679 58502 10717
rect 58110 10645 58122 10679
rect 58490 10645 58502 10679
rect 58110 10639 58502 10645
rect 58558 10598 58642 10798
rect 58698 10751 59090 10757
rect 58698 10717 58710 10751
rect 59078 10717 59090 10751
rect 58698 10679 59090 10717
rect 58698 10645 58710 10679
rect 59078 10645 59090 10679
rect 58698 10639 59090 10645
rect 59146 10598 59230 10798
rect 59286 10751 59678 10757
rect 59286 10717 59298 10751
rect 59666 10717 59678 10751
rect 59286 10679 59678 10717
rect 59286 10645 59298 10679
rect 59666 10645 59678 10679
rect 59286 10639 59678 10645
rect 59768 10598 59824 10798
rect 59874 10751 60266 10757
rect 59874 10717 59886 10751
rect 60254 10717 60266 10751
rect 59874 10679 60266 10717
rect 59874 10645 59886 10679
rect 60254 10645 60266 10679
rect 59874 10639 60266 10645
rect 60322 10598 60406 10798
rect 60462 10751 60854 10757
rect 60462 10717 60474 10751
rect 60842 10717 60854 10751
rect 60462 10679 60854 10717
rect 60462 10645 60474 10679
rect 60842 10645 60854 10679
rect 60462 10639 60854 10645
rect 60910 10598 60994 10798
rect 61050 10751 61442 10757
rect 61050 10717 61062 10751
rect 61430 10717 61442 10751
rect 61050 10679 61442 10717
rect 61050 10645 61062 10679
rect 61430 10645 61442 10679
rect 61050 10639 61442 10645
rect 61498 10598 61582 10798
rect 61638 10751 62030 10757
rect 61638 10717 61650 10751
rect 62018 10717 62030 10751
rect 61638 10679 62030 10717
rect 61638 10645 61650 10679
rect 62018 10645 62030 10679
rect 61638 10639 62030 10645
rect 62086 10598 62170 10798
rect 62226 10751 62618 10757
rect 62226 10717 62238 10751
rect 62606 10717 62618 10751
rect 62226 10679 62618 10717
rect 62226 10645 62238 10679
rect 62606 10645 62618 10679
rect 62226 10639 62618 10645
rect 62674 10598 62758 10798
rect 62814 10751 63206 10757
rect 62814 10717 62826 10751
rect 63194 10717 63206 10751
rect 62814 10679 63206 10717
rect 62814 10645 62826 10679
rect 63194 10645 63206 10679
rect 62814 10639 63206 10645
rect 63262 10598 63346 10798
rect 63402 10751 63794 10757
rect 63402 10717 63414 10751
rect 63782 10717 63794 10751
rect 63402 10679 63794 10717
rect 63402 10645 63414 10679
rect 63782 10645 63794 10679
rect 63402 10639 63794 10645
rect 63850 10598 63934 10798
rect 63990 10751 64382 10757
rect 63990 10717 64002 10751
rect 64370 10717 64382 10751
rect 63990 10679 64382 10717
rect 63990 10645 64002 10679
rect 64370 10645 64382 10679
rect 63990 10639 64382 10645
rect 64438 10598 64522 10798
rect 64578 10751 64970 10757
rect 64578 10717 64590 10751
rect 64958 10717 64970 10751
rect 64578 10679 64970 10717
rect 64578 10645 64590 10679
rect 64958 10645 64970 10679
rect 64578 10639 64970 10645
rect 65026 10598 65110 10798
rect 65166 10751 65558 10757
rect 65166 10717 65178 10751
rect 65546 10717 65558 10751
rect 65166 10679 65558 10717
rect 65166 10645 65178 10679
rect 65546 10645 65558 10679
rect 65166 10639 65558 10645
rect 65614 10598 65698 10798
rect 65754 10751 66146 10757
rect 65754 10717 65766 10751
rect 66134 10717 66146 10751
rect 65754 10679 66146 10717
rect 65754 10645 65766 10679
rect 66134 10645 66146 10679
rect 65754 10639 66146 10645
rect 66202 10598 66286 10798
rect 66342 10751 66734 10757
rect 66342 10717 66354 10751
rect 66722 10717 66734 10751
rect 66342 10679 66734 10717
rect 66342 10645 66354 10679
rect 66722 10645 66734 10679
rect 66342 10639 66734 10645
rect 66790 10598 66874 10798
rect 66930 10751 67322 10757
rect 66930 10717 66942 10751
rect 67310 10717 67322 10751
rect 66930 10679 67322 10717
rect 66930 10645 66942 10679
rect 67310 10645 67322 10679
rect 66930 10639 67322 10645
rect 67378 10598 67462 10798
rect 67518 10751 67910 10757
rect 67518 10717 67530 10751
rect 67898 10717 67910 10751
rect 67518 10679 67910 10717
rect 67518 10645 67530 10679
rect 67898 10645 67910 10679
rect 67518 10639 67910 10645
rect 67966 10598 68050 10798
rect 68106 10751 68498 10757
rect 68106 10717 68118 10751
rect 68486 10717 68498 10751
rect 68106 10679 68498 10717
rect 68106 10645 68118 10679
rect 68486 10645 68498 10679
rect 68106 10639 68498 10645
rect 68554 10598 68638 10798
rect 68694 10751 69086 10757
rect 68694 10717 68706 10751
rect 69074 10717 69086 10751
rect 68694 10679 69086 10717
rect 68694 10645 68706 10679
rect 69074 10645 69086 10679
rect 68694 10639 69086 10645
rect 69142 10598 69226 10798
rect 69282 10751 69674 10757
rect 69282 10717 69294 10751
rect 69662 10717 69674 10751
rect 69282 10679 69674 10717
rect 69282 10645 69294 10679
rect 69662 10645 69674 10679
rect 69282 10639 69674 10645
rect 69730 10598 69814 10798
rect 69870 10751 70262 10757
rect 69870 10717 69882 10751
rect 70250 10717 70262 10751
rect 69870 10679 70262 10717
rect 69870 10645 69882 10679
rect 70250 10645 70262 10679
rect 69870 10639 70262 10645
rect 70318 10598 70402 10798
rect 70458 10751 70850 10757
rect 70458 10717 70470 10751
rect 70838 10717 70850 10751
rect 70458 10679 70850 10717
rect 70458 10645 70470 10679
rect 70838 10645 70850 10679
rect 70458 10639 70850 10645
rect 70906 10598 70990 10798
rect 71046 10751 71438 10757
rect 71046 10717 71058 10751
rect 71426 10717 71438 10751
rect 71046 10679 71438 10717
rect 71046 10645 71058 10679
rect 71426 10645 71438 10679
rect 71046 10639 71438 10645
rect 71494 10598 71578 10798
rect 43270 10586 43400 10598
rect 43270 9810 43360 10586
rect 43394 9810 43400 10586
rect 43270 9798 43400 9810
rect 43812 10586 43988 10598
rect 43812 9810 43818 10586
rect 43852 9810 43948 10586
rect 43982 9810 43988 10586
rect 43812 9798 43988 9810
rect 44400 10586 44576 10598
rect 44400 9810 44406 10586
rect 44440 9810 44536 10586
rect 44570 9810 44576 10586
rect 44400 9798 44576 9810
rect 44988 10586 45164 10598
rect 44988 9810 44994 10586
rect 45028 9810 45124 10586
rect 45158 9810 45164 10586
rect 44988 9798 45164 9810
rect 45576 10586 45752 10598
rect 45576 9810 45582 10586
rect 45616 9810 45712 10586
rect 45746 9810 45752 10586
rect 45576 9798 45752 9810
rect 46164 10586 46340 10598
rect 46164 9810 46170 10586
rect 46204 9810 46300 10586
rect 46334 9810 46340 10586
rect 46164 9798 46340 9810
rect 46752 10586 46928 10598
rect 46752 9810 46758 10586
rect 46792 9810 46888 10586
rect 46922 9810 46928 10586
rect 46752 9798 46928 9810
rect 47340 10586 47516 10598
rect 47340 9810 47346 10586
rect 47380 9810 47476 10586
rect 47510 9810 47516 10586
rect 47340 9798 47516 9810
rect 47928 10586 48104 10598
rect 47928 9810 47934 10586
rect 47968 9810 48064 10586
rect 48098 9810 48104 10586
rect 47928 9798 48104 9810
rect 48516 10586 48692 10598
rect 48516 9810 48522 10586
rect 48556 9810 48652 10586
rect 48686 9810 48692 10586
rect 48516 9798 48692 9810
rect 49104 10586 49280 10598
rect 49104 9810 49110 10586
rect 49144 9810 49240 10586
rect 49274 9810 49280 10586
rect 49104 9798 49280 9810
rect 49692 10586 49868 10598
rect 49692 9810 49698 10586
rect 49732 9810 49828 10586
rect 49862 9810 49868 10586
rect 49692 9798 49868 9810
rect 50280 10586 50456 10598
rect 50280 9810 50286 10586
rect 50320 9810 50416 10586
rect 50450 9810 50456 10586
rect 50280 9798 50456 9810
rect 50868 10586 51044 10598
rect 50868 9810 50874 10586
rect 50908 9810 51004 10586
rect 51038 9810 51044 10586
rect 50868 9798 51044 9810
rect 51456 10586 51632 10598
rect 51456 9810 51462 10586
rect 51496 9810 51592 10586
rect 51626 9810 51632 10586
rect 51456 9798 51632 9810
rect 52044 10586 52220 10598
rect 52044 9810 52050 10586
rect 52084 9810 52180 10586
rect 52214 9810 52220 10586
rect 52044 9798 52220 9810
rect 52632 10586 52808 10598
rect 52632 9810 52638 10586
rect 52672 9810 52768 10586
rect 52802 9810 52808 10586
rect 52632 9798 52808 9810
rect 53220 10586 53396 10598
rect 53220 9810 53226 10586
rect 53260 9810 53356 10586
rect 53390 9810 53396 10586
rect 53220 9798 53396 9810
rect 53808 10586 53984 10598
rect 53808 9810 53814 10586
rect 53848 9810 53944 10586
rect 53978 9810 53984 10586
rect 53808 9798 53984 9810
rect 54396 10586 54572 10598
rect 54396 9810 54402 10586
rect 54436 9810 54532 10586
rect 54566 9810 54572 10586
rect 54396 9798 54572 9810
rect 54984 10586 55082 10598
rect 54984 9810 54990 10586
rect 55024 9810 55082 10586
rect 54984 9798 55082 9810
rect 55114 10586 55160 10598
rect 55114 9810 55120 10586
rect 55154 9810 55160 10586
rect 55114 9798 55160 9810
rect 55572 10586 55748 10598
rect 55572 9810 55578 10586
rect 55612 9810 55708 10586
rect 55742 9810 55748 10586
rect 55572 9798 55748 9810
rect 56160 10586 56336 10598
rect 56160 9810 56166 10586
rect 56200 9810 56296 10586
rect 56330 9810 56336 10586
rect 56160 9798 56336 9810
rect 56748 10586 56924 10598
rect 56748 9810 56754 10586
rect 56788 9810 56884 10586
rect 56918 9810 56924 10586
rect 56748 9798 56924 9810
rect 57336 10586 57382 10598
rect 57336 9810 57342 10586
rect 57376 9810 57382 10586
rect 57336 9798 57382 9810
rect 57466 10586 57512 10598
rect 57466 9810 57472 10586
rect 57506 9810 57512 10586
rect 57466 9798 57512 9810
rect 57924 10586 58100 10598
rect 57924 9810 57930 10586
rect 57964 9810 58060 10586
rect 58094 9810 58100 10586
rect 57924 9798 58100 9810
rect 58512 10586 58688 10598
rect 58512 9810 58518 10586
rect 58552 9810 58648 10586
rect 58682 9810 58688 10586
rect 58512 9798 58688 9810
rect 59100 10586 59276 10598
rect 59100 9810 59106 10586
rect 59140 9810 59236 10586
rect 59270 9810 59276 10586
rect 59100 9798 59276 9810
rect 59688 10586 59734 10598
rect 59688 9810 59694 10586
rect 59728 9810 59734 10586
rect 59688 9798 59734 9810
rect 59768 10586 59864 10598
rect 59768 9810 59824 10586
rect 59858 9810 59864 10586
rect 59768 9798 59864 9810
rect 60276 10586 60452 10598
rect 60276 9810 60282 10586
rect 60316 9810 60412 10586
rect 60446 9810 60452 10586
rect 60276 9798 60452 9810
rect 60864 10586 61040 10598
rect 60864 9810 60870 10586
rect 60904 9810 61000 10586
rect 61034 9810 61040 10586
rect 60864 9798 61040 9810
rect 61452 10586 61628 10598
rect 61452 9810 61458 10586
rect 61492 9810 61588 10586
rect 61622 9810 61628 10586
rect 61452 9798 61628 9810
rect 62040 10586 62216 10598
rect 62040 9810 62046 10586
rect 62080 9810 62176 10586
rect 62210 9810 62216 10586
rect 62040 9798 62216 9810
rect 62628 10586 62804 10598
rect 62628 9810 62634 10586
rect 62668 9810 62764 10586
rect 62798 9810 62804 10586
rect 62628 9798 62804 9810
rect 63216 10586 63392 10598
rect 63216 9810 63222 10586
rect 63256 9810 63352 10586
rect 63386 9810 63392 10586
rect 63216 9798 63392 9810
rect 63804 10586 63980 10598
rect 63804 9810 63810 10586
rect 63844 9810 63940 10586
rect 63974 9810 63980 10586
rect 63804 9798 63980 9810
rect 64392 10586 64568 10598
rect 64392 9810 64398 10586
rect 64432 9810 64528 10586
rect 64562 9810 64568 10586
rect 64392 9798 64568 9810
rect 64980 10586 65156 10598
rect 64980 9810 64986 10586
rect 65020 9810 65116 10586
rect 65150 9810 65156 10586
rect 64980 9798 65156 9810
rect 65568 10586 65744 10598
rect 65568 9810 65574 10586
rect 65608 9810 65704 10586
rect 65738 9810 65744 10586
rect 65568 9798 65744 9810
rect 66156 10586 66332 10598
rect 66156 9810 66162 10586
rect 66196 9810 66292 10586
rect 66326 9810 66332 10586
rect 66156 9798 66332 9810
rect 66744 10586 66920 10598
rect 66744 9810 66750 10586
rect 66784 9810 66880 10586
rect 66914 9810 66920 10586
rect 66744 9798 66920 9810
rect 67332 10586 67508 10598
rect 67332 9810 67338 10586
rect 67372 9810 67468 10586
rect 67502 9810 67508 10586
rect 67332 9798 67508 9810
rect 67920 10586 68096 10598
rect 67920 9810 67926 10586
rect 67960 9810 68056 10586
rect 68090 9810 68096 10586
rect 67920 9798 68096 9810
rect 68508 10586 68684 10598
rect 68508 9810 68514 10586
rect 68548 9810 68644 10586
rect 68678 9810 68684 10586
rect 68508 9798 68684 9810
rect 69096 10586 69272 10598
rect 69096 9810 69102 10586
rect 69136 9810 69232 10586
rect 69266 9810 69272 10586
rect 69096 9798 69272 9810
rect 69684 10586 69860 10598
rect 69684 9810 69690 10586
rect 69724 9810 69820 10586
rect 69854 9810 69860 10586
rect 69684 9798 69860 9810
rect 70272 10586 70448 10598
rect 70272 9810 70278 10586
rect 70312 9810 70408 10586
rect 70442 9810 70448 10586
rect 70272 9798 70448 9810
rect 70860 10586 71036 10598
rect 70860 9810 70866 10586
rect 70900 9810 70996 10586
rect 71030 9810 71036 10586
rect 70860 9798 71036 9810
rect 71448 10586 71578 10598
rect 71448 9810 71454 10586
rect 71488 9810 71578 10586
rect 71448 9798 71578 9810
rect 43410 9751 43802 9757
rect 43410 9717 43422 9751
rect 43790 9717 43802 9751
rect 43410 9711 43802 9717
rect 43864 9454 43936 9798
rect 43998 9751 44390 9757
rect 43998 9717 44010 9751
rect 44378 9717 44390 9751
rect 43998 9711 44390 9717
rect 44586 9751 44978 9757
rect 44586 9717 44598 9751
rect 44966 9717 44978 9751
rect 44586 9711 44978 9717
rect 45040 9454 45112 9798
rect 45174 9751 45566 9757
rect 45174 9717 45186 9751
rect 45554 9717 45566 9751
rect 45174 9711 45566 9717
rect 45762 9751 46154 9757
rect 45762 9717 45774 9751
rect 46142 9717 46154 9751
rect 45762 9711 46154 9717
rect 46216 9454 46288 9798
rect 46350 9751 46742 9757
rect 46350 9717 46362 9751
rect 46730 9717 46742 9751
rect 46350 9711 46742 9717
rect 46938 9751 47330 9757
rect 46938 9717 46950 9751
rect 47318 9717 47330 9751
rect 46938 9711 47330 9717
rect 47392 9454 47464 9798
rect 47526 9751 47918 9757
rect 47526 9717 47538 9751
rect 47906 9717 47918 9751
rect 47526 9711 47918 9717
rect 48114 9751 48506 9757
rect 48114 9717 48126 9751
rect 48494 9717 48506 9751
rect 48114 9711 48506 9717
rect 48568 9454 48640 9798
rect 48702 9751 49094 9757
rect 48702 9717 48714 9751
rect 49082 9717 49094 9751
rect 48702 9711 49094 9717
rect 49290 9751 49682 9757
rect 49290 9717 49302 9751
rect 49670 9717 49682 9751
rect 49290 9711 49682 9717
rect 49744 9454 49816 9798
rect 49878 9751 50270 9757
rect 49878 9717 49890 9751
rect 50258 9717 50270 9751
rect 49878 9711 50270 9717
rect 50466 9751 50858 9757
rect 50466 9717 50478 9751
rect 50846 9717 50858 9751
rect 50466 9711 50858 9717
rect 50920 9454 50992 9798
rect 51054 9751 51446 9757
rect 51054 9717 51066 9751
rect 51434 9717 51446 9751
rect 51054 9711 51446 9717
rect 51642 9751 52034 9757
rect 51642 9717 51654 9751
rect 52022 9717 52034 9751
rect 51642 9711 52034 9717
rect 52096 9454 52168 9798
rect 52230 9751 52622 9757
rect 52230 9717 52242 9751
rect 52610 9717 52622 9751
rect 52230 9711 52622 9717
rect 52818 9751 53210 9757
rect 52818 9717 52830 9751
rect 53198 9717 53210 9751
rect 52818 9711 53210 9717
rect 53272 9454 53344 9798
rect 53406 9751 53798 9757
rect 53406 9717 53418 9751
rect 53786 9717 53798 9751
rect 53406 9711 53798 9717
rect 53994 9751 54386 9757
rect 53994 9717 54006 9751
rect 54374 9717 54386 9751
rect 53994 9711 54386 9717
rect 54448 9454 54520 9798
rect 54582 9751 54974 9757
rect 54582 9717 54594 9751
rect 54962 9717 54974 9751
rect 54582 9711 54974 9717
rect 55170 9751 55562 9757
rect 55170 9717 55182 9751
rect 55550 9717 55562 9751
rect 55170 9711 55562 9717
rect 55624 9454 55696 9798
rect 55758 9751 56150 9757
rect 55758 9717 55770 9751
rect 56138 9717 56150 9751
rect 55758 9711 56150 9717
rect 43794 9448 44006 9454
rect 43794 9338 43806 9448
rect 43994 9338 44006 9448
rect 43794 9332 44006 9338
rect 44970 9448 45182 9454
rect 44970 9338 44982 9448
rect 45170 9338 45182 9448
rect 44970 9332 45182 9338
rect 46146 9448 46358 9454
rect 46146 9338 46158 9448
rect 46346 9338 46358 9448
rect 46146 9332 46358 9338
rect 47322 9448 47534 9454
rect 47322 9338 47334 9448
rect 47522 9338 47534 9448
rect 47322 9332 47534 9338
rect 48498 9448 48710 9454
rect 48498 9338 48510 9448
rect 48698 9338 48710 9448
rect 48498 9332 48710 9338
rect 49674 9448 49886 9454
rect 49674 9338 49686 9448
rect 49874 9338 49886 9448
rect 49674 9332 49886 9338
rect 50850 9448 51062 9454
rect 50850 9338 50862 9448
rect 51050 9338 51062 9448
rect 50850 9332 51062 9338
rect 52026 9448 52238 9454
rect 52026 9338 52038 9448
rect 52226 9338 52238 9448
rect 52026 9332 52238 9338
rect 53202 9448 53414 9454
rect 53202 9338 53214 9448
rect 53402 9338 53414 9448
rect 53202 9332 53414 9338
rect 54378 9448 54590 9454
rect 54378 9338 54390 9448
rect 54578 9338 54590 9448
rect 54378 9332 54590 9338
rect 55554 9448 55766 9454
rect 55554 9338 55566 9448
rect 55754 9338 55766 9448
rect 55554 9332 55766 9338
rect 56212 8946 56284 9798
rect 56346 9751 56738 9757
rect 56346 9717 56358 9751
rect 56726 9717 56738 9751
rect 56346 9711 56738 9717
rect 56800 9454 56872 9798
rect 56934 9751 57326 9757
rect 56934 9717 56946 9751
rect 57314 9717 57326 9751
rect 56934 9711 57326 9717
rect 57522 9751 57914 9757
rect 57522 9717 57534 9751
rect 57902 9717 57914 9751
rect 57522 9711 57914 9717
rect 57976 9454 58048 9798
rect 58110 9751 58502 9757
rect 58110 9717 58122 9751
rect 58490 9717 58502 9751
rect 58110 9711 58502 9717
rect 56730 9448 56942 9454
rect 56730 9338 56742 9448
rect 56930 9338 56942 9448
rect 56730 9332 56942 9338
rect 57906 9448 58118 9454
rect 57906 9338 57918 9448
rect 58106 9338 58118 9448
rect 57906 9332 58118 9338
rect 58564 8946 58636 9798
rect 58698 9751 59090 9757
rect 58698 9717 58710 9751
rect 59078 9717 59090 9751
rect 58698 9711 59090 9717
rect 59152 9454 59224 9798
rect 59286 9751 59678 9757
rect 59286 9717 59298 9751
rect 59666 9717 59678 9751
rect 59286 9711 59678 9717
rect 59874 9751 60266 9757
rect 59874 9717 59886 9751
rect 60254 9717 60266 9751
rect 59874 9711 60266 9717
rect 60328 9454 60400 9798
rect 60462 9751 60854 9757
rect 60462 9717 60474 9751
rect 60842 9717 60854 9751
rect 60462 9711 60854 9717
rect 61050 9751 61442 9757
rect 61050 9717 61062 9751
rect 61430 9717 61442 9751
rect 61050 9711 61442 9717
rect 61504 9454 61576 9798
rect 61638 9751 62030 9757
rect 61638 9717 61650 9751
rect 62018 9717 62030 9751
rect 61638 9711 62030 9717
rect 62226 9751 62618 9757
rect 62226 9717 62238 9751
rect 62606 9717 62618 9751
rect 62226 9711 62618 9717
rect 62680 9464 62752 9798
rect 62814 9751 63206 9757
rect 62814 9717 62826 9751
rect 63194 9717 63206 9751
rect 62814 9711 63206 9717
rect 63402 9751 63794 9757
rect 63402 9717 63414 9751
rect 63782 9717 63794 9751
rect 63402 9711 63794 9717
rect 62610 9458 62822 9464
rect 59082 9448 59294 9454
rect 59082 9338 59094 9448
rect 59282 9338 59294 9448
rect 59082 9332 59294 9338
rect 60258 9448 60470 9454
rect 60258 9338 60270 9448
rect 60458 9338 60470 9448
rect 60258 9332 60470 9338
rect 61434 9448 61646 9454
rect 61434 9338 61446 9448
rect 61634 9338 61646 9448
rect 62610 9348 62622 9458
rect 62810 9348 62822 9458
rect 63856 9454 63928 9798
rect 63990 9751 64382 9757
rect 63990 9717 64002 9751
rect 64370 9717 64382 9751
rect 63990 9711 64382 9717
rect 64578 9751 64970 9757
rect 64578 9717 64590 9751
rect 64958 9717 64970 9751
rect 64578 9711 64970 9717
rect 65032 9454 65104 9798
rect 65166 9751 65558 9757
rect 65166 9717 65178 9751
rect 65546 9717 65558 9751
rect 65166 9711 65558 9717
rect 65754 9751 66146 9757
rect 65754 9717 65766 9751
rect 66134 9717 66146 9751
rect 65754 9711 66146 9717
rect 66208 9454 66280 9798
rect 66342 9751 66734 9757
rect 66342 9717 66354 9751
rect 66722 9717 66734 9751
rect 66342 9711 66734 9717
rect 66930 9751 67322 9757
rect 66930 9717 66942 9751
rect 67310 9717 67322 9751
rect 66930 9711 67322 9717
rect 67384 9464 67456 9798
rect 67518 9751 67910 9757
rect 67518 9717 67530 9751
rect 67898 9717 67910 9751
rect 67518 9711 67910 9717
rect 68106 9751 68498 9757
rect 68106 9717 68118 9751
rect 68486 9717 68498 9751
rect 68106 9711 68498 9717
rect 67300 9458 67536 9464
rect 62610 9342 62822 9348
rect 63786 9448 63998 9454
rect 61434 9332 61646 9338
rect 63786 9338 63798 9448
rect 63986 9338 63998 9448
rect 63786 9332 63998 9338
rect 64962 9448 65174 9454
rect 64962 9338 64974 9448
rect 65162 9338 65174 9448
rect 64962 9332 65174 9338
rect 66138 9448 66350 9454
rect 66138 9338 66150 9448
rect 66338 9338 66350 9448
rect 66138 9332 66350 9338
rect 67300 9336 67312 9458
rect 67524 9336 67536 9458
rect 68560 9454 68632 9798
rect 68694 9751 69086 9757
rect 68694 9717 68706 9751
rect 69074 9717 69086 9751
rect 68694 9711 69086 9717
rect 69282 9751 69674 9757
rect 69282 9717 69294 9751
rect 69662 9717 69674 9751
rect 69282 9711 69674 9717
rect 69736 9454 69808 9798
rect 69870 9751 70262 9757
rect 69870 9717 69882 9751
rect 70250 9717 70262 9751
rect 69870 9711 70262 9717
rect 70458 9751 70850 9757
rect 70458 9717 70470 9751
rect 70838 9717 70850 9751
rect 70458 9711 70850 9717
rect 70912 9454 70984 9798
rect 71046 9751 71438 9757
rect 71046 9717 71058 9751
rect 71426 9717 71438 9751
rect 71046 9711 71438 9717
rect 67300 9330 67536 9336
rect 68490 9448 68702 9454
rect 68490 9338 68502 9448
rect 68690 9338 68702 9448
rect 68490 9332 68702 9338
rect 69666 9448 69878 9454
rect 69666 9338 69678 9448
rect 69866 9338 69878 9448
rect 69666 9332 69878 9338
rect 70842 9448 71054 9454
rect 70842 9338 70854 9448
rect 71042 9338 71054 9448
rect 70842 9332 71054 9338
rect 56212 8866 58636 8946
rect 56320 8152 56400 8866
rect 56456 8322 56530 8328
rect 56456 8190 56466 8322
rect 56520 8190 56530 8322
rect 56456 8184 56530 8190
rect 56722 8322 56796 8328
rect 56722 8190 56732 8322
rect 56786 8190 56796 8322
rect 56722 8184 56796 8190
rect 56852 8152 56932 8866
rect 56988 8322 57062 8328
rect 56988 8190 56998 8322
rect 57052 8190 57062 8322
rect 56988 8184 57062 8190
rect 57254 8322 57328 8328
rect 57254 8190 57264 8322
rect 57318 8190 57328 8322
rect 57254 8184 57328 8190
rect 57384 8152 57464 8866
rect 57520 8322 57594 8328
rect 57520 8190 57530 8322
rect 57584 8190 57594 8322
rect 57520 8184 57594 8190
rect 57786 8322 57860 8328
rect 57786 8190 57796 8322
rect 57850 8190 57860 8322
rect 57786 8184 57860 8190
rect 57916 8152 57996 8866
rect 58052 8322 58126 8328
rect 58052 8190 58062 8322
rect 58116 8190 58126 8322
rect 58052 8184 58126 8190
rect 58318 8322 58392 8328
rect 58318 8190 58328 8322
rect 58382 8190 58392 8322
rect 58318 8184 58392 8190
rect 58448 8152 58528 8866
rect 56320 8140 56452 8152
rect 56320 7364 56412 8140
rect 56446 7364 56452 8140
rect 56320 7352 56452 7364
rect 56534 8140 56718 8152
rect 56534 7364 56540 8140
rect 56574 7364 56678 8140
rect 56712 7364 56718 8140
rect 56534 7352 56718 7364
rect 56800 8140 56984 8152
rect 56800 7364 56806 8140
rect 56840 7364 56944 8140
rect 56978 7364 56984 8140
rect 56800 7352 56984 7364
rect 57066 8140 57250 8152
rect 57066 7364 57072 8140
rect 57106 7364 57210 8140
rect 57244 7364 57250 8140
rect 57066 7352 57250 7364
rect 57332 8140 57516 8152
rect 57332 7364 57338 8140
rect 57372 7364 57476 8140
rect 57510 7364 57516 8140
rect 57332 7352 57516 7364
rect 57598 8140 57782 8152
rect 57598 7364 57604 8140
rect 57638 7364 57742 8140
rect 57776 7364 57782 8140
rect 57598 7352 57782 7364
rect 57864 8140 58048 8152
rect 57864 7364 57870 8140
rect 57904 7364 58008 8140
rect 58042 7364 58048 8140
rect 57864 7352 58048 7364
rect 58130 8140 58314 8152
rect 58130 7364 58136 8140
rect 58170 7364 58274 8140
rect 58308 7364 58314 8140
rect 58130 7352 58314 7364
rect 58396 8140 58528 8152
rect 58396 7364 58402 8140
rect 58436 7364 58528 8140
rect 58396 7352 58528 7364
rect 56320 7142 56406 7352
rect 56456 7312 56530 7318
rect 56456 7180 56466 7312
rect 56520 7180 56530 7312
rect 56456 7174 56530 7180
rect 56580 7142 56672 7352
rect 56722 7312 56796 7318
rect 56722 7180 56732 7312
rect 56786 7180 56796 7312
rect 56722 7174 56796 7180
rect 56846 7142 56938 7352
rect 56988 7312 57062 7318
rect 56988 7180 56998 7312
rect 57052 7180 57062 7312
rect 56988 7174 57062 7180
rect 57112 7142 57204 7352
rect 57254 7312 57328 7318
rect 57254 7180 57264 7312
rect 57318 7180 57328 7312
rect 57254 7174 57328 7180
rect 57378 7142 57470 7352
rect 57520 7312 57594 7318
rect 57520 7180 57530 7312
rect 57584 7180 57594 7312
rect 57520 7174 57594 7180
rect 57644 7142 57736 7352
rect 57786 7312 57860 7318
rect 57786 7180 57796 7312
rect 57850 7180 57860 7312
rect 57786 7174 57860 7180
rect 57910 7142 58002 7352
rect 58052 7312 58126 7318
rect 58052 7180 58062 7312
rect 58116 7180 58126 7312
rect 58052 7174 58126 7180
rect 58176 7142 58268 7352
rect 58318 7312 58392 7318
rect 58318 7180 58328 7312
rect 58382 7180 58392 7312
rect 58318 7174 58392 7180
rect 58442 7142 58528 7352
rect 56320 7130 56452 7142
rect 56320 6354 56412 7130
rect 56446 6354 56452 7130
rect 56320 6342 56452 6354
rect 56534 7130 56718 7142
rect 56534 6354 56540 7130
rect 56574 6354 56678 7130
rect 56712 6354 56718 7130
rect 56534 6342 56718 6354
rect 56800 7130 56984 7142
rect 56800 6354 56806 7130
rect 56840 6354 56944 7130
rect 56978 6354 56984 7130
rect 56800 6342 56984 6354
rect 57066 7130 57250 7142
rect 57066 6354 57072 7130
rect 57106 6354 57210 7130
rect 57244 6354 57250 7130
rect 57066 6342 57250 6354
rect 57332 7130 57516 7142
rect 57332 6354 57338 7130
rect 57372 6354 57476 7130
rect 57510 6354 57516 7130
rect 57332 6342 57516 6354
rect 57598 7130 57782 7142
rect 57598 6354 57604 7130
rect 57638 6354 57742 7130
rect 57776 6354 57782 7130
rect 57598 6342 57782 6354
rect 57864 7130 58048 7142
rect 57864 6354 57870 7130
rect 57904 6354 58008 7130
rect 58042 6354 58048 7130
rect 57864 6342 58048 6354
rect 58130 7130 58314 7142
rect 58130 6354 58136 7130
rect 58170 6354 58274 7130
rect 58308 6354 58314 7130
rect 58130 6342 58314 6354
rect 58396 7130 58528 7142
rect 58396 6354 58402 7130
rect 58436 6354 58528 7130
rect 58396 6342 58528 6354
rect 56320 6132 56406 6342
rect 56456 6302 56530 6308
rect 56456 6170 56466 6302
rect 56520 6170 56530 6302
rect 56456 6164 56530 6170
rect 56580 6132 56672 6342
rect 56722 6302 56796 6308
rect 56722 6170 56732 6302
rect 56786 6170 56796 6302
rect 56722 6164 56796 6170
rect 56846 6132 56938 6342
rect 56988 6302 57062 6308
rect 56988 6170 56998 6302
rect 57052 6170 57062 6302
rect 56988 6164 57062 6170
rect 57112 6132 57204 6342
rect 57254 6302 57328 6308
rect 57254 6170 57264 6302
rect 57318 6170 57328 6302
rect 57254 6164 57328 6170
rect 57378 6132 57470 6342
rect 57520 6302 57594 6308
rect 57520 6170 57530 6302
rect 57584 6170 57594 6302
rect 57520 6164 57594 6170
rect 57644 6132 57736 6342
rect 57786 6302 57860 6308
rect 57786 6170 57796 6302
rect 57850 6170 57860 6302
rect 57786 6164 57860 6170
rect 57910 6132 58002 6342
rect 58052 6302 58126 6308
rect 58052 6170 58062 6302
rect 58116 6170 58126 6302
rect 58052 6164 58126 6170
rect 58176 6132 58268 6342
rect 58318 6302 58392 6308
rect 58318 6170 58328 6302
rect 58382 6170 58392 6302
rect 58318 6164 58392 6170
rect 58442 6132 58528 6342
rect 56320 6120 56452 6132
rect 56320 5344 56412 6120
rect 56446 5344 56452 6120
rect 56320 5332 56452 5344
rect 56534 6120 56718 6132
rect 56534 5344 56540 6120
rect 56574 5344 56678 6120
rect 56712 5344 56718 6120
rect 56534 5332 56718 5344
rect 56800 6120 56984 6132
rect 56800 5344 56806 6120
rect 56840 5344 56944 6120
rect 56978 5344 56984 6120
rect 56800 5332 56984 5344
rect 57066 6120 57250 6132
rect 57066 5344 57072 6120
rect 57106 5344 57210 6120
rect 57244 5344 57250 6120
rect 57066 5332 57250 5344
rect 57332 6120 57516 6132
rect 57332 5344 57338 6120
rect 57372 5344 57476 6120
rect 57510 5344 57516 6120
rect 57332 5332 57516 5344
rect 57598 6120 57782 6132
rect 57598 5344 57604 6120
rect 57638 5344 57742 6120
rect 57776 5344 57782 6120
rect 57598 5332 57782 5344
rect 57864 6120 58048 6132
rect 57864 5344 57870 6120
rect 57904 5344 58008 6120
rect 58042 5344 58048 6120
rect 57864 5332 58048 5344
rect 58130 6120 58314 6132
rect 58130 5344 58136 6120
rect 58170 5344 58274 6120
rect 58308 5344 58314 6120
rect 58130 5332 58314 5344
rect 58396 6120 58528 6132
rect 58396 5344 58402 6120
rect 58436 5344 58528 6120
rect 58396 5332 58528 5344
rect 56456 5292 56530 5298
rect 56456 5160 56466 5292
rect 56520 5160 56530 5292
rect 56456 5154 56530 5160
rect 56586 3960 56666 5332
rect 56722 5292 56796 5298
rect 56722 5160 56732 5292
rect 56786 5160 56796 5292
rect 56722 5154 56796 5160
rect 56988 5292 57062 5298
rect 56988 5160 56998 5292
rect 57052 5160 57062 5292
rect 56988 5154 57062 5160
rect 57118 4776 57198 5332
rect 57254 5292 57328 5298
rect 57254 5160 57264 5292
rect 57318 5160 57328 5292
rect 57254 5154 57328 5160
rect 57520 5292 57594 5298
rect 57520 5160 57530 5292
rect 57584 5160 57594 5292
rect 57520 5154 57594 5160
rect 57650 4776 57730 5332
rect 57786 5292 57860 5298
rect 57786 5160 57796 5292
rect 57850 5160 57860 5292
rect 57786 5154 57860 5160
rect 58052 5292 58126 5298
rect 58052 5160 58062 5292
rect 58116 5160 58126 5292
rect 58052 5154 58126 5160
rect 57118 4744 57730 4776
rect 57118 4616 57164 4744
rect 57658 4616 57730 4744
rect 57118 4586 57730 4616
rect 57030 4124 57340 4130
rect 57030 3998 57046 4124
rect 57084 3998 57286 4124
rect 57324 3998 57340 4124
rect 57030 3992 57100 3998
rect 57270 3992 57340 3998
rect 57398 3960 57452 4586
rect 57510 4124 57820 4130
rect 57510 3998 57526 4124
rect 57564 3998 57766 4124
rect 57804 3998 57820 4124
rect 57510 3992 57580 3998
rect 57750 3992 57820 3998
rect 58182 3960 58262 5332
rect 58318 5292 58392 5298
rect 58318 5160 58328 5292
rect 58382 5160 58392 5292
rect 58318 5154 58392 5160
rect 56586 3948 57024 3960
rect 56586 3890 56984 3948
rect 56934 3372 56984 3890
rect 57018 3372 57024 3948
rect 56934 3360 57024 3372
rect 57106 3948 57264 3960
rect 57106 3372 57112 3948
rect 57146 3372 57224 3948
rect 57258 3372 57264 3948
rect 57106 3360 57264 3372
rect 57346 3948 57504 3960
rect 57346 3372 57352 3948
rect 57386 3372 57464 3948
rect 57498 3372 57504 3948
rect 57346 3360 57504 3372
rect 57586 3948 57744 3960
rect 57586 3372 57592 3948
rect 57626 3372 57704 3948
rect 57738 3372 57744 3948
rect 57586 3360 57744 3372
rect 57826 3948 58262 3960
rect 57826 3372 57832 3948
rect 57866 3890 58262 3948
rect 57866 3372 57922 3890
rect 57826 3360 57922 3372
rect 56934 3152 56984 3360
rect 57030 3322 57100 3328
rect 57030 3190 57046 3322
rect 57084 3190 57100 3322
rect 57030 3184 57100 3190
rect 57152 3152 57218 3360
rect 57270 3322 57340 3328
rect 57270 3190 57286 3322
rect 57324 3190 57340 3322
rect 57270 3184 57340 3190
rect 57392 3152 57458 3360
rect 57510 3322 57580 3328
rect 57510 3190 57526 3322
rect 57564 3190 57580 3322
rect 57510 3184 57580 3190
rect 57632 3152 57698 3360
rect 57750 3322 57820 3328
rect 57750 3190 57766 3322
rect 57804 3190 57820 3322
rect 57750 3184 57820 3190
rect 57872 3152 57922 3360
rect 56934 3140 57024 3152
rect 56934 2564 56984 3140
rect 57018 2564 57024 3140
rect 56934 2552 57024 2564
rect 57106 3140 57264 3152
rect 57106 2564 57112 3140
rect 57146 2564 57224 3140
rect 57258 2564 57264 3140
rect 57106 2552 57264 2564
rect 57346 3140 57504 3152
rect 57346 2564 57352 3140
rect 57386 2564 57464 3140
rect 57498 2564 57504 3140
rect 57346 2552 57504 2564
rect 57586 3140 57744 3152
rect 57586 2564 57592 3140
rect 57626 2564 57704 3140
rect 57738 2564 57744 3140
rect 57586 2552 57744 2564
rect 57826 3140 57922 3152
rect 57826 2564 57832 3140
rect 57866 2564 57922 3140
rect 57826 2552 57922 2564
rect 57030 2514 57100 2520
rect 57030 2382 57046 2514
rect 57084 2382 57100 2514
rect 57030 2376 57100 2382
rect 57158 2136 57212 2552
rect 57270 2514 57340 2520
rect 57270 2382 57286 2514
rect 57324 2382 57340 2514
rect 57270 2376 57340 2382
rect 57510 2514 57580 2520
rect 57510 2382 57526 2514
rect 57564 2382 57580 2514
rect 57510 2376 57580 2382
rect 57638 2136 57692 2552
rect 57750 2514 57820 2520
rect 57750 2382 57766 2514
rect 57804 2382 57820 2514
rect 57750 2376 57820 2382
rect 56724 2130 58100 2136
rect 56724 2018 56736 2130
rect 58088 2018 58100 2130
rect 56724 2012 58100 2018
<< via1 >>
rect 52810 17114 52920 17186
rect 53290 17114 53400 17186
rect 53770 17114 53880 17186
rect 54250 17114 54360 17186
rect 54730 17114 54840 17186
rect 55210 17114 55320 17186
rect 55690 17114 55800 17186
rect 56170 17114 56280 17186
rect 56650 17114 56760 17186
rect 57130 17114 57240 17186
rect 57610 17114 57720 17186
rect 58090 17114 58200 17186
rect 58570 17114 58680 17186
rect 59050 17114 59160 17186
rect 59530 17114 59640 17186
rect 60010 17114 60120 17186
rect 60490 17114 60600 17186
rect 60970 17114 61080 17186
rect 61450 17114 61560 17186
rect 61930 17114 62040 17186
rect 52710 16710 52726 16842
rect 52726 16710 52764 16842
rect 52764 16710 52780 16842
rect 52950 16710 52966 16842
rect 52966 16710 53004 16842
rect 53004 16710 53020 16842
rect 53190 16710 53206 16842
rect 53206 16710 53244 16842
rect 53244 16710 53260 16842
rect 53430 16710 53446 16842
rect 53446 16710 53484 16842
rect 53484 16710 53500 16842
rect 53670 16710 53686 16842
rect 53686 16710 53724 16842
rect 53724 16710 53740 16842
rect 53910 16710 53926 16842
rect 53926 16710 53964 16842
rect 53964 16710 53980 16842
rect 54150 16710 54166 16842
rect 54166 16710 54204 16842
rect 54204 16710 54220 16842
rect 54390 16710 54406 16842
rect 54406 16710 54444 16842
rect 54444 16710 54460 16842
rect 54630 16710 54646 16842
rect 54646 16710 54684 16842
rect 54684 16710 54700 16842
rect 54870 16710 54886 16842
rect 54886 16710 54924 16842
rect 54924 16710 54940 16842
rect 55110 16710 55126 16842
rect 55126 16710 55164 16842
rect 55164 16710 55180 16842
rect 55350 16710 55366 16842
rect 55366 16710 55404 16842
rect 55404 16710 55420 16842
rect 55590 16710 55606 16842
rect 55606 16710 55644 16842
rect 55644 16710 55660 16842
rect 55830 16710 55846 16842
rect 55846 16710 55884 16842
rect 55884 16710 55900 16842
rect 56070 16710 56086 16842
rect 56086 16710 56124 16842
rect 56124 16710 56140 16842
rect 56310 16710 56326 16842
rect 56326 16710 56364 16842
rect 56364 16710 56380 16842
rect 56550 16710 56566 16842
rect 56566 16710 56604 16842
rect 56604 16710 56620 16842
rect 56790 16710 56806 16842
rect 56806 16710 56844 16842
rect 56844 16710 56860 16842
rect 57030 16710 57046 16842
rect 57046 16710 57084 16842
rect 57084 16710 57100 16842
rect 57270 16710 57286 16842
rect 57286 16710 57324 16842
rect 57324 16710 57340 16842
rect 57510 16710 57526 16842
rect 57526 16710 57564 16842
rect 57564 16710 57580 16842
rect 57750 16710 57766 16842
rect 57766 16710 57804 16842
rect 57804 16710 57820 16842
rect 57990 16710 58006 16842
rect 58006 16710 58044 16842
rect 58044 16710 58060 16842
rect 58230 16710 58246 16842
rect 58246 16710 58284 16842
rect 58284 16710 58300 16842
rect 58470 16710 58486 16842
rect 58486 16710 58524 16842
rect 58524 16710 58540 16842
rect 58710 16710 58726 16842
rect 58726 16710 58764 16842
rect 58764 16710 58780 16842
rect 58950 16710 58966 16842
rect 58966 16710 59004 16842
rect 59004 16710 59020 16842
rect 59190 16710 59206 16842
rect 59206 16710 59244 16842
rect 59244 16710 59260 16842
rect 59430 16710 59446 16842
rect 59446 16710 59484 16842
rect 59484 16710 59500 16842
rect 59670 16710 59686 16842
rect 59686 16710 59724 16842
rect 59724 16710 59740 16842
rect 59910 16710 59926 16842
rect 59926 16710 59964 16842
rect 59964 16710 59980 16842
rect 60150 16710 60166 16842
rect 60166 16710 60204 16842
rect 60204 16710 60220 16842
rect 60390 16710 60406 16842
rect 60406 16710 60444 16842
rect 60444 16710 60460 16842
rect 60630 16710 60646 16842
rect 60646 16710 60684 16842
rect 60684 16710 60700 16842
rect 60870 16710 60886 16842
rect 60886 16710 60924 16842
rect 60924 16710 60940 16842
rect 61110 16710 61126 16842
rect 61126 16710 61164 16842
rect 61164 16710 61180 16842
rect 61350 16710 61366 16842
rect 61366 16710 61404 16842
rect 61404 16710 61420 16842
rect 61590 16710 61606 16842
rect 61606 16710 61644 16842
rect 61644 16710 61660 16842
rect 61830 16710 61846 16842
rect 61846 16710 61884 16842
rect 61884 16710 61900 16842
rect 62070 16710 62086 16842
rect 62086 16710 62124 16842
rect 62124 16710 62140 16842
rect 52710 15902 52726 16034
rect 52726 15902 52764 16034
rect 52764 15902 52780 16034
rect 52950 15902 52966 16034
rect 52966 15902 53004 16034
rect 53004 15902 53020 16034
rect 53190 15902 53206 16034
rect 53206 15902 53244 16034
rect 53244 15902 53260 16034
rect 53430 15902 53446 16034
rect 53446 15902 53484 16034
rect 53484 15902 53500 16034
rect 53670 15902 53686 16034
rect 53686 15902 53724 16034
rect 53724 15902 53740 16034
rect 53910 15902 53926 16034
rect 53926 15902 53964 16034
rect 53964 15902 53980 16034
rect 54150 15902 54166 16034
rect 54166 15902 54204 16034
rect 54204 15902 54220 16034
rect 54390 15902 54406 16034
rect 54406 15902 54444 16034
rect 54444 15902 54460 16034
rect 54630 15902 54646 16034
rect 54646 15902 54684 16034
rect 54684 15902 54700 16034
rect 54870 15902 54886 16034
rect 54886 15902 54924 16034
rect 54924 15902 54940 16034
rect 55110 15902 55126 16034
rect 55126 15902 55164 16034
rect 55164 15902 55180 16034
rect 55350 15902 55366 16034
rect 55366 15902 55404 16034
rect 55404 15902 55420 16034
rect 55590 15902 55606 16034
rect 55606 15902 55644 16034
rect 55644 15902 55660 16034
rect 55830 15902 55846 16034
rect 55846 15902 55884 16034
rect 55884 15902 55900 16034
rect 56070 15902 56086 16034
rect 56086 15902 56124 16034
rect 56124 15902 56140 16034
rect 56310 15902 56326 16034
rect 56326 15902 56364 16034
rect 56364 15902 56380 16034
rect 56550 15902 56566 16034
rect 56566 15902 56604 16034
rect 56604 15902 56620 16034
rect 56790 15902 56806 16034
rect 56806 15902 56844 16034
rect 56844 15902 56860 16034
rect 57030 15902 57046 16034
rect 57046 15902 57084 16034
rect 57084 15902 57100 16034
rect 57270 15902 57286 16034
rect 57286 15902 57324 16034
rect 57324 15902 57340 16034
rect 57510 15902 57526 16034
rect 57526 15902 57564 16034
rect 57564 15902 57580 16034
rect 57750 15902 57766 16034
rect 57766 15902 57804 16034
rect 57804 15902 57820 16034
rect 57990 15902 58006 16034
rect 58006 15902 58044 16034
rect 58044 15902 58060 16034
rect 58230 15902 58246 16034
rect 58246 15902 58284 16034
rect 58284 15902 58300 16034
rect 58470 15902 58486 16034
rect 58486 15902 58524 16034
rect 58524 15902 58540 16034
rect 58710 15902 58726 16034
rect 58726 15902 58764 16034
rect 58764 15902 58780 16034
rect 58950 15902 58966 16034
rect 58966 15902 59004 16034
rect 59004 15902 59020 16034
rect 59190 15902 59206 16034
rect 59206 15902 59244 16034
rect 59244 15902 59260 16034
rect 59430 15902 59446 16034
rect 59446 15902 59484 16034
rect 59484 15902 59500 16034
rect 59670 15902 59686 16034
rect 59686 15902 59724 16034
rect 59724 15902 59740 16034
rect 59910 15902 59926 16034
rect 59926 15902 59964 16034
rect 59964 15902 59980 16034
rect 60150 15902 60166 16034
rect 60166 15902 60204 16034
rect 60204 15902 60220 16034
rect 60390 15902 60406 16034
rect 60406 15902 60444 16034
rect 60444 15902 60460 16034
rect 60630 15902 60646 16034
rect 60646 15902 60684 16034
rect 60684 15902 60700 16034
rect 60870 15902 60886 16034
rect 60886 15902 60924 16034
rect 60924 15902 60940 16034
rect 61110 15902 61126 16034
rect 61126 15902 61164 16034
rect 61164 15902 61180 16034
rect 61350 15902 61366 16034
rect 61366 15902 61404 16034
rect 61404 15902 61420 16034
rect 61590 15902 61606 16034
rect 61606 15902 61644 16034
rect 61644 15902 61660 16034
rect 61830 15902 61846 16034
rect 61846 15902 61884 16034
rect 61884 15902 61900 16034
rect 62070 15902 62086 16034
rect 62086 15902 62124 16034
rect 62124 15902 62140 16034
rect 52710 15094 52726 15226
rect 52726 15094 52764 15226
rect 52764 15094 52780 15226
rect 52950 15094 52966 15226
rect 52966 15094 53004 15226
rect 53004 15094 53020 15226
rect 53190 15094 53206 15226
rect 53206 15094 53244 15226
rect 53244 15094 53260 15226
rect 53430 15094 53446 15226
rect 53446 15094 53484 15226
rect 53484 15094 53500 15226
rect 53670 15094 53686 15226
rect 53686 15094 53724 15226
rect 53724 15094 53740 15226
rect 53910 15094 53926 15226
rect 53926 15094 53964 15226
rect 53964 15094 53980 15226
rect 54150 15094 54166 15226
rect 54166 15094 54204 15226
rect 54204 15094 54220 15226
rect 54390 15094 54406 15226
rect 54406 15094 54444 15226
rect 54444 15094 54460 15226
rect 54630 15094 54646 15226
rect 54646 15094 54684 15226
rect 54684 15094 54700 15226
rect 54870 15094 54886 15226
rect 54886 15094 54924 15226
rect 54924 15094 54940 15226
rect 55110 15094 55126 15226
rect 55126 15094 55164 15226
rect 55164 15094 55180 15226
rect 55350 15094 55366 15226
rect 55366 15094 55404 15226
rect 55404 15094 55420 15226
rect 55590 15094 55606 15226
rect 55606 15094 55644 15226
rect 55644 15094 55660 15226
rect 55830 15094 55846 15226
rect 55846 15094 55884 15226
rect 55884 15094 55900 15226
rect 56070 15094 56086 15226
rect 56086 15094 56124 15226
rect 56124 15094 56140 15226
rect 56310 15094 56326 15226
rect 56326 15094 56364 15226
rect 56364 15094 56380 15226
rect 56550 15094 56566 15226
rect 56566 15094 56604 15226
rect 56604 15094 56620 15226
rect 56790 15094 56806 15226
rect 56806 15094 56844 15226
rect 56844 15094 56860 15226
rect 57030 15094 57046 15226
rect 57046 15094 57084 15226
rect 57084 15094 57100 15226
rect 57270 15094 57286 15226
rect 57286 15094 57324 15226
rect 57324 15094 57340 15226
rect 57510 15094 57526 15226
rect 57526 15094 57564 15226
rect 57564 15094 57580 15226
rect 57750 15094 57766 15226
rect 57766 15094 57804 15226
rect 57804 15094 57820 15226
rect 57990 15094 58006 15226
rect 58006 15094 58044 15226
rect 58044 15094 58060 15226
rect 58230 15094 58246 15226
rect 58246 15094 58284 15226
rect 58284 15094 58300 15226
rect 58470 15094 58486 15226
rect 58486 15094 58524 15226
rect 58524 15094 58540 15226
rect 58710 15094 58726 15226
rect 58726 15094 58764 15226
rect 58764 15094 58780 15226
rect 58950 15094 58966 15226
rect 58966 15094 59004 15226
rect 59004 15094 59020 15226
rect 59190 15094 59206 15226
rect 59206 15094 59244 15226
rect 59244 15094 59260 15226
rect 59430 15094 59446 15226
rect 59446 15094 59484 15226
rect 59484 15094 59500 15226
rect 59670 15094 59686 15226
rect 59686 15094 59724 15226
rect 59724 15094 59740 15226
rect 59910 15094 59926 15226
rect 59926 15094 59964 15226
rect 59964 15094 59980 15226
rect 60150 15094 60166 15226
rect 60166 15094 60204 15226
rect 60204 15094 60220 15226
rect 60390 15094 60406 15226
rect 60406 15094 60444 15226
rect 60444 15094 60460 15226
rect 60630 15094 60646 15226
rect 60646 15094 60684 15226
rect 60684 15094 60700 15226
rect 60870 15094 60886 15226
rect 60886 15094 60924 15226
rect 60924 15094 60940 15226
rect 61110 15094 61126 15226
rect 61126 15094 61164 15226
rect 61164 15094 61180 15226
rect 61350 15094 61366 15226
rect 61366 15094 61404 15226
rect 61404 15094 61420 15226
rect 61590 15094 61606 15226
rect 61606 15094 61644 15226
rect 61644 15094 61660 15226
rect 61830 15094 61846 15226
rect 61846 15094 61884 15226
rect 61884 15094 61900 15226
rect 62070 15094 62086 15226
rect 62086 15094 62124 15226
rect 62124 15094 62140 15226
rect 43806 9338 43994 9448
rect 44982 9338 45170 9448
rect 46158 9338 46346 9448
rect 47334 9338 47522 9448
rect 48510 9338 48698 9448
rect 49686 9338 49874 9448
rect 50862 9338 51050 9448
rect 52038 9338 52226 9448
rect 53214 9338 53402 9448
rect 54390 9338 54578 9448
rect 55566 9338 55754 9448
rect 56742 9338 56930 9448
rect 57918 9338 58106 9448
rect 59094 9338 59282 9448
rect 60270 9338 60458 9448
rect 61446 9338 61634 9448
rect 63798 9338 63986 9448
rect 64974 9338 65162 9448
rect 66150 9338 66338 9448
rect 68502 9338 68690 9448
rect 69678 9338 69866 9448
rect 70854 9338 71042 9448
rect 56466 8190 56474 8322
rect 56474 8190 56512 8322
rect 56512 8190 56520 8322
rect 56732 8190 56740 8322
rect 56740 8190 56778 8322
rect 56778 8190 56786 8322
rect 56998 8190 57006 8322
rect 57006 8190 57044 8322
rect 57044 8190 57052 8322
rect 57264 8190 57272 8322
rect 57272 8190 57310 8322
rect 57310 8190 57318 8322
rect 57530 8190 57538 8322
rect 57538 8190 57576 8322
rect 57576 8190 57584 8322
rect 57796 8190 57804 8322
rect 57804 8190 57842 8322
rect 57842 8190 57850 8322
rect 58062 8190 58070 8322
rect 58070 8190 58108 8322
rect 58108 8190 58116 8322
rect 58328 8190 58336 8322
rect 58336 8190 58374 8322
rect 58374 8190 58382 8322
rect 56466 7180 56474 7312
rect 56474 7180 56512 7312
rect 56512 7180 56520 7312
rect 56732 7180 56740 7312
rect 56740 7180 56778 7312
rect 56778 7180 56786 7312
rect 56998 7180 57006 7312
rect 57006 7180 57044 7312
rect 57044 7180 57052 7312
rect 57264 7180 57272 7312
rect 57272 7180 57310 7312
rect 57310 7180 57318 7312
rect 57530 7180 57538 7312
rect 57538 7180 57576 7312
rect 57576 7180 57584 7312
rect 57796 7180 57804 7312
rect 57804 7180 57842 7312
rect 57842 7180 57850 7312
rect 58062 7180 58070 7312
rect 58070 7180 58108 7312
rect 58108 7180 58116 7312
rect 58328 7180 58336 7312
rect 58336 7180 58374 7312
rect 58374 7180 58382 7312
rect 56466 6170 56474 6302
rect 56474 6170 56512 6302
rect 56512 6170 56520 6302
rect 56732 6170 56740 6302
rect 56740 6170 56778 6302
rect 56778 6170 56786 6302
rect 56998 6170 57006 6302
rect 57006 6170 57044 6302
rect 57044 6170 57052 6302
rect 57264 6170 57272 6302
rect 57272 6170 57310 6302
rect 57310 6170 57318 6302
rect 57530 6170 57538 6302
rect 57538 6170 57576 6302
rect 57576 6170 57584 6302
rect 57796 6170 57804 6302
rect 57804 6170 57842 6302
rect 57842 6170 57850 6302
rect 58062 6170 58070 6302
rect 58070 6170 58108 6302
rect 58108 6170 58116 6302
rect 58328 6170 58336 6302
rect 58336 6170 58374 6302
rect 58374 6170 58382 6302
rect 56466 5160 56474 5292
rect 56474 5160 56512 5292
rect 56512 5160 56520 5292
rect 56732 5160 56740 5292
rect 56740 5160 56778 5292
rect 56778 5160 56786 5292
rect 56998 5160 57006 5292
rect 57006 5160 57044 5292
rect 57044 5160 57052 5292
rect 57264 5160 57272 5292
rect 57272 5160 57310 5292
rect 57310 5160 57318 5292
rect 57530 5160 57538 5292
rect 57538 5160 57576 5292
rect 57576 5160 57584 5292
rect 57796 5160 57804 5292
rect 57804 5160 57842 5292
rect 57842 5160 57850 5292
rect 58062 5160 58070 5292
rect 58070 5160 58108 5292
rect 58108 5160 58116 5292
rect 57164 4616 57658 4744
rect 58328 5160 58336 5292
rect 58336 5160 58374 5292
rect 58374 5160 58382 5292
rect 56736 2018 58088 2130
<< metal2 >>
rect 52810 17186 52920 17196
rect 52810 17104 52920 17114
rect 53290 17186 53400 17196
rect 53290 17104 53400 17114
rect 53770 17186 53880 17196
rect 53770 17104 53880 17114
rect 54250 17186 54360 17196
rect 54250 17104 54360 17114
rect 54730 17186 54840 17196
rect 54730 17104 54840 17114
rect 55210 17186 55320 17196
rect 55210 17104 55320 17114
rect 55690 17186 55800 17196
rect 55690 17104 55800 17114
rect 56170 17186 56280 17196
rect 56170 17104 56280 17114
rect 56650 17186 56760 17196
rect 56650 17104 56760 17114
rect 57130 17186 57240 17196
rect 57130 17104 57240 17114
rect 57610 17186 57720 17196
rect 57610 17104 57720 17114
rect 58090 17186 58200 17196
rect 58090 17104 58200 17114
rect 58570 17186 58680 17196
rect 58570 17104 58680 17114
rect 59050 17186 59160 17196
rect 59050 17104 59160 17114
rect 59530 17186 59640 17196
rect 59530 17104 59640 17114
rect 60010 17186 60120 17196
rect 60010 17104 60120 17114
rect 60490 17186 60600 17196
rect 60490 17104 60600 17114
rect 60970 17186 61080 17196
rect 60970 17104 61080 17114
rect 61450 17186 61560 17196
rect 61450 17104 61560 17114
rect 61930 17186 62040 17196
rect 61930 17104 62040 17114
rect 62748 17000 63048 17010
rect 52700 16842 62748 16852
rect 52700 16710 52710 16842
rect 52780 16710 52950 16842
rect 53020 16710 53190 16842
rect 53260 16710 53430 16842
rect 53500 16710 53670 16842
rect 53740 16710 53910 16842
rect 53980 16710 54150 16842
rect 54220 16710 54390 16842
rect 54460 16710 54630 16842
rect 54700 16710 54870 16842
rect 54940 16710 55110 16842
rect 55180 16710 55350 16842
rect 55420 16710 55590 16842
rect 55660 16710 55830 16842
rect 55900 16710 56070 16842
rect 56140 16710 56310 16842
rect 56380 16710 56550 16842
rect 56620 16710 56790 16842
rect 56860 16710 57030 16842
rect 57100 16710 57270 16842
rect 57340 16710 57510 16842
rect 57580 16710 57750 16842
rect 57820 16710 57990 16842
rect 58060 16710 58230 16842
rect 58300 16710 58470 16842
rect 58540 16710 58710 16842
rect 58780 16710 58950 16842
rect 59020 16710 59190 16842
rect 59260 16710 59430 16842
rect 59500 16710 59670 16842
rect 59740 16710 59910 16842
rect 59980 16710 60150 16842
rect 60220 16710 60390 16842
rect 60460 16710 60630 16842
rect 60700 16710 60870 16842
rect 60940 16710 61110 16842
rect 61180 16710 61350 16842
rect 61420 16710 61590 16842
rect 61660 16710 61830 16842
rect 61900 16710 62070 16842
rect 62140 16710 62748 16842
rect 52700 16700 62748 16710
rect 62748 16690 63048 16700
rect 62748 16192 63048 16202
rect 52700 16034 62748 16044
rect 52700 15902 52710 16034
rect 52780 15902 52950 16034
rect 53020 15902 53190 16034
rect 53260 15902 53430 16034
rect 53500 15902 53670 16034
rect 53740 15902 53910 16034
rect 53980 15902 54150 16034
rect 54220 15902 54390 16034
rect 54460 15902 54630 16034
rect 54700 15902 54870 16034
rect 54940 15902 55110 16034
rect 55180 15902 55350 16034
rect 55420 15902 55590 16034
rect 55660 15902 55830 16034
rect 55900 15902 56070 16034
rect 56140 15902 56310 16034
rect 56380 15902 56550 16034
rect 56620 15902 56790 16034
rect 56860 15902 57030 16034
rect 57100 15902 57270 16034
rect 57340 15902 57510 16034
rect 57580 15902 57750 16034
rect 57820 15902 57990 16034
rect 58060 15902 58230 16034
rect 58300 15902 58470 16034
rect 58540 15902 58710 16034
rect 58780 15902 58950 16034
rect 59020 15902 59190 16034
rect 59260 15902 59430 16034
rect 59500 15902 59670 16034
rect 59740 15902 59910 16034
rect 59980 15902 60150 16034
rect 60220 15902 60390 16034
rect 60460 15902 60630 16034
rect 60700 15902 60870 16034
rect 60940 15902 61110 16034
rect 61180 15902 61350 16034
rect 61420 15902 61590 16034
rect 61660 15902 61830 16034
rect 61900 15902 62070 16034
rect 62140 15902 62748 16034
rect 52700 15892 62748 15902
rect 62748 15882 63048 15892
rect 62748 15384 63048 15394
rect 52700 15226 62748 15236
rect 52700 15094 52710 15226
rect 52780 15094 52950 15226
rect 53020 15094 53190 15226
rect 53260 15094 53430 15226
rect 53500 15094 53670 15226
rect 53740 15094 53910 15226
rect 53980 15094 54150 15226
rect 54220 15094 54390 15226
rect 54460 15094 54630 15226
rect 54700 15094 54870 15226
rect 54940 15094 55110 15226
rect 55180 15094 55350 15226
rect 55420 15094 55590 15226
rect 55660 15094 55830 15226
rect 55900 15094 56070 15226
rect 56140 15094 56310 15226
rect 56380 15094 56550 15226
rect 56620 15094 56790 15226
rect 56860 15094 57030 15226
rect 57100 15094 57270 15226
rect 57340 15094 57510 15226
rect 57580 15094 57750 15226
rect 57820 15094 57990 15226
rect 58060 15094 58230 15226
rect 58300 15094 58470 15226
rect 58540 15094 58710 15226
rect 58780 15094 58950 15226
rect 59020 15094 59190 15226
rect 59260 15094 59430 15226
rect 59500 15094 59670 15226
rect 59740 15094 59910 15226
rect 59980 15094 60150 15226
rect 60220 15094 60390 15226
rect 60460 15094 60630 15226
rect 60700 15094 60870 15226
rect 60940 15094 61110 15226
rect 61180 15094 61350 15226
rect 61420 15094 61590 15226
rect 61660 15094 61830 15226
rect 61900 15094 62070 15226
rect 62140 15094 62748 15226
rect 52700 15084 62748 15094
rect 62748 15074 63048 15084
rect 43806 9448 43994 9458
rect 43806 9328 43994 9338
rect 44982 9448 45170 9458
rect 44982 9328 45170 9338
rect 46158 9448 46346 9458
rect 46158 9328 46346 9338
rect 47334 9448 47522 9458
rect 47334 9328 47522 9338
rect 48510 9448 48698 9458
rect 48510 9328 48698 9338
rect 49686 9448 49874 9458
rect 49686 9328 49874 9338
rect 50862 9448 51050 9458
rect 50862 9328 51050 9338
rect 52038 9448 52226 9458
rect 52038 9328 52226 9338
rect 53214 9448 53402 9458
rect 53214 9328 53402 9338
rect 54390 9448 54578 9458
rect 54390 9328 54578 9338
rect 55566 9448 55754 9458
rect 55566 9328 55754 9338
rect 56742 9448 56930 9458
rect 56742 9328 56930 9338
rect 57918 9448 58106 9458
rect 57918 9328 58106 9338
rect 59094 9448 59282 9458
rect 59094 9328 59282 9338
rect 60270 9448 60458 9458
rect 60270 9328 60458 9338
rect 61446 9448 61634 9458
rect 61446 9328 61634 9338
rect 63798 9448 63986 9458
rect 63798 9328 63986 9338
rect 64974 9448 65162 9458
rect 64974 9328 65162 9338
rect 66150 9448 66338 9458
rect 66150 9328 66338 9338
rect 68502 9448 68690 9458
rect 68502 9328 68690 9338
rect 69678 9448 69866 9458
rect 69678 9328 69866 9338
rect 70854 9448 71042 9458
rect 70854 9328 71042 9338
rect 56998 8446 59176 8572
rect 56998 8332 57318 8446
rect 56466 8322 56786 8332
rect 56520 8190 56732 8322
rect 56466 8066 56786 8190
rect 56998 8322 57052 8332
rect 56998 8180 57052 8190
rect 57264 8322 57318 8332
rect 57264 8180 57318 8190
rect 57530 8322 57850 8446
rect 57584 8190 57796 8322
rect 57530 8184 57850 8190
rect 58062 8322 58116 8332
rect 58062 8184 58116 8190
rect 58328 8322 58382 8332
rect 58328 8184 58382 8190
rect 58062 8066 58382 8184
rect 55672 7940 58382 8066
rect 55672 7056 55920 7940
rect 58928 7562 59176 8446
rect 56998 7436 59176 7562
rect 56998 7322 57318 7436
rect 57538 7322 57858 7436
rect 56466 7312 56520 7322
rect 56466 7170 56520 7180
rect 56732 7312 56786 7322
rect 56732 7170 56786 7180
rect 56998 7312 57052 7322
rect 56998 7170 57052 7180
rect 57264 7312 57318 7322
rect 57264 7170 57318 7180
rect 57530 7312 57584 7322
rect 57530 7170 57584 7180
rect 57796 7312 57850 7322
rect 57796 7170 57850 7180
rect 58062 7312 58116 7322
rect 58062 7170 58116 7180
rect 58328 7312 58382 7322
rect 58328 7170 58382 7180
rect 56466 7056 56786 7170
rect 58062 7056 58382 7170
rect 55672 6930 58382 7056
rect 55672 6046 55920 6930
rect 58928 6552 59176 7436
rect 56998 6426 59176 6552
rect 56998 6312 57318 6426
rect 56466 6302 56520 6312
rect 56466 6160 56520 6170
rect 56732 6302 56786 6312
rect 56732 6160 56786 6170
rect 56998 6302 57052 6312
rect 56998 6160 57052 6170
rect 57264 6302 57318 6312
rect 57264 6160 57318 6170
rect 57530 6308 57850 6426
rect 57530 6302 57584 6308
rect 57530 6160 57584 6170
rect 57796 6302 57850 6308
rect 57796 6160 57850 6170
rect 58062 6302 58116 6312
rect 58062 6160 58116 6170
rect 58328 6302 58382 6312
rect 58328 6160 58382 6170
rect 56466 6046 56786 6160
rect 58062 6046 58382 6160
rect 55672 5920 58382 6046
rect 55672 5036 55920 5920
rect 58928 5542 59176 6426
rect 56998 5416 59176 5542
rect 56998 5302 57318 5416
rect 56466 5292 56520 5302
rect 56466 5150 56520 5160
rect 56732 5292 56786 5302
rect 56732 5150 56786 5160
rect 56998 5292 57052 5302
rect 56998 5150 57052 5160
rect 57264 5292 57318 5302
rect 57264 5150 57318 5160
rect 57530 5302 57850 5416
rect 57530 5292 57584 5302
rect 57530 5150 57584 5160
rect 57796 5292 57850 5302
rect 57796 5150 57850 5160
rect 58062 5292 58116 5302
rect 58062 5150 58116 5160
rect 58328 5292 58382 5302
rect 58328 5150 58382 5160
rect 56466 5036 56786 5150
rect 58062 5036 58382 5150
rect 55672 4910 58382 5036
rect 62758 4906 63058 4916
rect 57164 4744 62758 4754
rect 57658 4616 62758 4744
rect 57164 4606 62758 4616
rect 63058 4606 63068 4754
rect 62758 4596 63058 4606
rect 56736 2130 58088 2140
rect 56736 2008 58088 2018
<< via2 >>
rect 52810 17114 52920 17186
rect 53290 17114 53400 17186
rect 53770 17114 53880 17186
rect 54250 17114 54360 17186
rect 54730 17114 54840 17186
rect 55210 17114 55320 17186
rect 55690 17114 55800 17186
rect 56170 17114 56280 17186
rect 56650 17114 56760 17186
rect 57130 17114 57240 17186
rect 57610 17114 57720 17186
rect 58090 17114 58200 17186
rect 58570 17114 58680 17186
rect 59050 17114 59160 17186
rect 59530 17114 59640 17186
rect 60010 17114 60120 17186
rect 60490 17114 60600 17186
rect 60970 17114 61080 17186
rect 61450 17114 61560 17186
rect 61930 17114 62040 17186
rect 62748 16700 63048 17000
rect 62748 15892 63048 16192
rect 62748 15084 63048 15384
rect 43806 9338 43994 9448
rect 44982 9338 45170 9448
rect 46158 9338 46346 9448
rect 47334 9338 47522 9448
rect 48510 9338 48698 9448
rect 49686 9338 49874 9448
rect 50862 9338 51050 9448
rect 52038 9338 52226 9448
rect 53214 9338 53402 9448
rect 54390 9338 54578 9448
rect 55566 9338 55754 9448
rect 56742 9338 56930 9448
rect 57918 9338 58106 9448
rect 59094 9338 59282 9448
rect 60270 9338 60458 9448
rect 61446 9338 61634 9448
rect 63798 9338 63986 9448
rect 64974 9338 65162 9448
rect 66150 9338 66338 9448
rect 68502 9338 68690 9448
rect 69678 9338 69866 9448
rect 70854 9338 71042 9448
rect 62758 4606 63058 4906
rect 56736 2018 58088 2130
<< metal3 >>
rect 52800 17186 52930 17191
rect 52800 17114 52810 17186
rect 52920 17114 52930 17186
rect 52800 17109 52930 17114
rect 53280 17186 53410 17191
rect 53280 17114 53290 17186
rect 53400 17114 53410 17186
rect 53280 17109 53410 17114
rect 53760 17186 53890 17191
rect 53760 17114 53770 17186
rect 53880 17114 53890 17186
rect 53760 17109 53890 17114
rect 54240 17186 54370 17191
rect 54240 17114 54250 17186
rect 54360 17114 54370 17186
rect 54240 17109 54370 17114
rect 54720 17186 54850 17191
rect 54720 17114 54730 17186
rect 54840 17114 54850 17186
rect 54720 17109 54850 17114
rect 55200 17186 55330 17191
rect 55200 17114 55210 17186
rect 55320 17114 55330 17186
rect 55200 17109 55330 17114
rect 55680 17186 55810 17191
rect 55680 17114 55690 17186
rect 55800 17114 55810 17186
rect 55680 17109 55810 17114
rect 56160 17186 56290 17191
rect 56160 17114 56170 17186
rect 56280 17114 56290 17186
rect 56160 17109 56290 17114
rect 56640 17186 56770 17191
rect 56640 17114 56650 17186
rect 56760 17114 56770 17186
rect 56640 17109 56770 17114
rect 57120 17186 57250 17191
rect 57120 17114 57130 17186
rect 57240 17114 57250 17186
rect 57120 17109 57250 17114
rect 57600 17186 57730 17191
rect 57600 17114 57610 17186
rect 57720 17114 57730 17186
rect 57600 17109 57730 17114
rect 58080 17186 58210 17191
rect 58080 17114 58090 17186
rect 58200 17114 58210 17186
rect 58080 17109 58210 17114
rect 58560 17186 58690 17191
rect 58560 17114 58570 17186
rect 58680 17114 58690 17186
rect 58560 17109 58690 17114
rect 59040 17186 59170 17191
rect 59040 17114 59050 17186
rect 59160 17114 59170 17186
rect 59040 17109 59170 17114
rect 59520 17186 59650 17191
rect 59520 17114 59530 17186
rect 59640 17114 59650 17186
rect 59520 17109 59650 17114
rect 60000 17186 60130 17191
rect 60000 17114 60010 17186
rect 60120 17114 60130 17186
rect 60000 17109 60130 17114
rect 60480 17186 60610 17191
rect 60480 17114 60490 17186
rect 60600 17114 60610 17186
rect 60480 17109 60610 17114
rect 60960 17186 61090 17191
rect 60960 17114 60970 17186
rect 61080 17114 61090 17186
rect 60960 17109 61090 17114
rect 61440 17186 61570 17191
rect 61440 17114 61450 17186
rect 61560 17114 61570 17186
rect 61440 17109 61570 17114
rect 61920 17186 62050 17191
rect 61920 17114 61930 17186
rect 62040 17114 62050 17186
rect 61920 17109 62050 17114
rect 62738 17004 63058 17005
rect 62738 17000 63068 17004
rect 62738 16700 62748 17000
rect 63048 16700 63068 17000
rect 62738 16695 63068 16700
rect 62748 16197 63068 16695
rect 62738 16192 63068 16197
rect 62738 15892 62748 16192
rect 63048 15892 63068 16192
rect 62738 15887 63068 15892
rect 62748 15389 63068 15887
rect 62738 15384 63068 15389
rect 62738 15084 62748 15384
rect 63048 15084 63068 15384
rect 62738 15079 63068 15084
rect 43796 9448 44004 9453
rect 43796 9338 43806 9448
rect 43994 9338 44004 9448
rect 43796 9333 44004 9338
rect 44972 9448 45180 9453
rect 44972 9338 44982 9448
rect 45170 9338 45180 9448
rect 44972 9333 45180 9338
rect 46148 9448 46356 9453
rect 46148 9338 46158 9448
rect 46346 9338 46356 9448
rect 46148 9333 46356 9338
rect 47324 9448 47532 9453
rect 47324 9338 47334 9448
rect 47522 9338 47532 9448
rect 47324 9333 47532 9338
rect 48500 9448 48708 9453
rect 48500 9338 48510 9448
rect 48698 9338 48708 9448
rect 48500 9333 48708 9338
rect 49676 9448 49884 9453
rect 49676 9338 49686 9448
rect 49874 9338 49884 9448
rect 49676 9333 49884 9338
rect 50852 9448 51060 9453
rect 50852 9338 50862 9448
rect 51050 9338 51060 9448
rect 50852 9333 51060 9338
rect 52028 9448 52236 9453
rect 52028 9338 52038 9448
rect 52226 9338 52236 9448
rect 52028 9333 52236 9338
rect 53204 9448 53412 9453
rect 53204 9338 53214 9448
rect 53402 9338 53412 9448
rect 53204 9333 53412 9338
rect 54380 9448 54588 9453
rect 54380 9338 54390 9448
rect 54578 9338 54588 9448
rect 54380 9333 54588 9338
rect 55556 9448 55764 9453
rect 55556 9338 55566 9448
rect 55754 9338 55764 9448
rect 55556 9333 55764 9338
rect 56732 9448 56940 9453
rect 56732 9338 56742 9448
rect 56930 9338 56940 9448
rect 56732 9333 56940 9338
rect 57908 9448 58116 9453
rect 57908 9338 57918 9448
rect 58106 9338 58116 9448
rect 57908 9333 58116 9338
rect 59084 9448 59292 9453
rect 59084 9338 59094 9448
rect 59282 9338 59292 9448
rect 59084 9333 59292 9338
rect 60260 9448 60468 9453
rect 60260 9338 60270 9448
rect 60458 9338 60468 9448
rect 60260 9333 60468 9338
rect 61436 9448 61644 9453
rect 61436 9338 61446 9448
rect 61634 9338 61644 9448
rect 61436 9333 61644 9338
rect 62748 4906 63068 15079
rect 63788 9448 63996 9453
rect 63788 9338 63798 9448
rect 63986 9338 63996 9448
rect 63788 9333 63996 9338
rect 64964 9448 65172 9453
rect 64964 9338 64974 9448
rect 65162 9338 65172 9448
rect 64964 9333 65172 9338
rect 66140 9448 66348 9453
rect 66140 9338 66150 9448
rect 66338 9338 66348 9448
rect 66140 9333 66348 9338
rect 68492 9448 68700 9453
rect 68492 9338 68502 9448
rect 68690 9338 68700 9448
rect 68492 9333 68700 9338
rect 69668 9448 69876 9453
rect 69668 9338 69678 9448
rect 69866 9338 69876 9448
rect 69668 9333 69876 9338
rect 70844 9448 71052 9453
rect 70844 9338 70854 9448
rect 71042 9338 71052 9448
rect 70844 9333 71052 9338
rect 62748 4606 62758 4906
rect 63058 4606 63068 4906
rect 62748 4601 63068 4606
rect 56726 2130 58098 2135
rect 56726 2018 56736 2130
rect 58088 2018 58098 2130
rect 56726 2013 58098 2018
<< via3 >>
rect 52810 17114 52920 17186
rect 53290 17114 53400 17186
rect 53770 17114 53880 17186
rect 54250 17114 54360 17186
rect 54730 17114 54840 17186
rect 55210 17114 55320 17186
rect 55690 17114 55800 17186
rect 56170 17114 56280 17186
rect 56650 17114 56760 17186
rect 57130 17114 57240 17186
rect 57610 17114 57720 17186
rect 58090 17114 58200 17186
rect 58570 17114 58680 17186
rect 59050 17114 59160 17186
rect 59530 17114 59640 17186
rect 60010 17114 60120 17186
rect 60490 17114 60600 17186
rect 60970 17114 61080 17186
rect 61450 17114 61560 17186
rect 61930 17114 62040 17186
rect 43806 9338 43994 9448
rect 44982 9338 45170 9448
rect 46158 9338 46346 9448
rect 47334 9338 47522 9448
rect 48510 9338 48698 9448
rect 49686 9338 49874 9448
rect 50862 9338 51050 9448
rect 52038 9338 52226 9448
rect 53214 9338 53402 9448
rect 54390 9338 54578 9448
rect 55566 9338 55754 9448
rect 56742 9338 56930 9448
rect 57918 9338 58106 9448
rect 59094 9338 59282 9448
rect 60270 9338 60458 9448
rect 61446 9338 61634 9448
rect 63798 9338 63986 9448
rect 64974 9338 65162 9448
rect 66150 9338 66338 9448
rect 68502 9338 68690 9448
rect 69678 9338 69866 9448
rect 70854 9338 71042 9448
rect 56736 2018 58088 2130
<< metal4 >>
rect 41122 17818 68492 17892
rect 40040 17186 68492 17818
rect 40040 17114 52810 17186
rect 52920 17114 53290 17186
rect 53400 17114 53770 17186
rect 53880 17114 54250 17186
rect 54360 17114 54730 17186
rect 54840 17114 55210 17186
rect 55320 17114 55690 17186
rect 55800 17114 56170 17186
rect 56280 17114 56650 17186
rect 56760 17114 57130 17186
rect 57240 17114 57610 17186
rect 57720 17114 58090 17186
rect 58200 17114 58570 17186
rect 58680 17114 59050 17186
rect 59160 17114 59530 17186
rect 59640 17114 60010 17186
rect 60120 17114 60490 17186
rect 60600 17114 60970 17186
rect 61080 17114 61450 17186
rect 61560 17114 61930 17186
rect 62040 17114 68492 17186
rect 40040 16628 68492 17114
rect 40040 16626 46658 16628
rect 40040 3024 41422 16626
rect 41782 9448 72106 10312
rect 41782 9338 43806 9448
rect 43994 9338 44982 9448
rect 45170 9338 46158 9448
rect 46346 9338 47334 9448
rect 47522 9338 48510 9448
rect 48698 9338 49686 9448
rect 49874 9338 50862 9448
rect 51050 9338 52038 9448
rect 52226 9338 53214 9448
rect 53402 9338 54390 9448
rect 54578 9338 55566 9448
rect 55754 9338 56742 9448
rect 56930 9338 57918 9448
rect 58106 9338 59094 9448
rect 59282 9338 60270 9448
rect 60458 9338 61446 9448
rect 61634 9338 63798 9448
rect 63986 9338 64974 9448
rect 65162 9338 66150 9448
rect 66338 9338 68502 9448
rect 68690 9338 69678 9448
rect 69866 9338 70854 9448
rect 71042 9338 72106 9448
rect 41782 8780 72106 9338
rect 40040 2130 72106 3024
rect 40040 2018 56736 2130
rect 58088 2018 72106 2130
rect 40040 1492 72106 2018
rect 40040 1490 41422 1492
<< labels >>
flabel metal1 70056 13890 70056 13890 0 FreeSans 1600 0 0 0 vout
port 5 nsew
flabel metal1 43580 10694 43580 10694 0 FreeSans 1600 0 0 0 vbias
port 3 nsew
flabel metal2 55764 6712 55764 6712 0 FreeSans 1600 0 0 0 vn
port 2 nsew
flabel metal2 59012 7180 59012 7180 0 FreeSans 1600 0 0 0 vp
port 1 nsew
flabel metal4 42244 9298 42244 9298 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal4 42442 2164 42442 2164 0 FreeSans 1600 0 0 0 vss
port 4 nsew
<< end >>
