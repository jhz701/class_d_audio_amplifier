magic
tech sky130A
magscale 1 2
timestamp 1628692234
<< nwell >>
rect 19191 8743 31315 10853
rect 20679 4119 23875 8465
<< pwell >>
rect 20679 1897 29827 3771
<< pmoslvt >>
rect 19387 10234 19587 10634
rect 19759 10234 19959 10634
rect 20131 10234 20331 10634
rect 20503 10234 20703 10634
rect 20875 10234 21075 10634
rect 21247 10234 21447 10634
rect 21619 10234 21819 10634
rect 21991 10234 22191 10634
rect 22363 10234 22563 10634
rect 22735 10234 22935 10634
rect 23107 10234 23307 10634
rect 23479 10234 23679 10634
rect 23851 10234 24051 10634
rect 24223 10234 24423 10634
rect 24595 10234 24795 10634
rect 24967 10234 25167 10634
rect 25339 10234 25539 10634
rect 25711 10234 25911 10634
rect 26083 10234 26283 10634
rect 26455 10234 26655 10634
rect 26827 10234 27027 10634
rect 27199 10234 27399 10634
rect 27571 10234 27771 10634
rect 27943 10234 28143 10634
rect 28315 10234 28515 10634
rect 28687 10234 28887 10634
rect 29059 10234 29259 10634
rect 29431 10234 29631 10634
rect 29803 10234 30003 10634
rect 30175 10234 30375 10634
rect 30547 10234 30747 10634
rect 30919 10234 31119 10634
rect 19387 9598 19587 9998
rect 19759 9598 19959 9998
rect 20131 9598 20331 9998
rect 20503 9598 20703 9998
rect 20875 9598 21075 9998
rect 21247 9598 21447 9998
rect 21619 9598 21819 9998
rect 21991 9598 22191 9998
rect 22363 9598 22563 9998
rect 22735 9598 22935 9998
rect 23107 9598 23307 9998
rect 23479 9598 23679 9998
rect 23851 9598 24051 9998
rect 24223 9598 24423 9998
rect 24595 9598 24795 9998
rect 24967 9598 25167 9998
rect 25339 9598 25539 9998
rect 25711 9598 25911 9998
rect 26083 9598 26283 9998
rect 26455 9598 26655 9998
rect 26827 9598 27027 9998
rect 27199 9598 27399 9998
rect 27571 9598 27771 9998
rect 27943 9598 28143 9998
rect 28315 9598 28515 9998
rect 28687 9598 28887 9998
rect 29059 9598 29259 9998
rect 29431 9598 29631 9998
rect 29803 9598 30003 9998
rect 30175 9598 30375 9998
rect 30547 9598 30747 9998
rect 30919 9598 31119 9998
rect 19387 8962 19587 9362
rect 19759 8962 19959 9362
rect 20131 8962 20331 9362
rect 20503 8962 20703 9362
rect 20875 8962 21075 9362
rect 21247 8962 21447 9362
rect 21619 8962 21819 9362
rect 21991 8962 22191 9362
rect 22363 8962 22563 9362
rect 22735 8962 22935 9362
rect 23107 8962 23307 9362
rect 23479 8962 23679 9362
rect 23851 8962 24051 9362
rect 24223 8962 24423 9362
rect 24595 8962 24795 9362
rect 24967 8962 25167 9362
rect 25339 8962 25539 9362
rect 25711 8962 25911 9362
rect 26083 8962 26283 9362
rect 26455 8962 26655 9362
rect 26827 8962 27027 9362
rect 27199 8962 27399 9362
rect 27571 8962 27771 9362
rect 27943 8962 28143 9362
rect 28315 8962 28515 9362
rect 28687 8962 28887 9362
rect 29059 8962 29259 9362
rect 29431 8962 29631 9362
rect 29803 8962 30003 9362
rect 30175 8962 30375 9362
rect 30547 8962 30747 9362
rect 30919 8962 31119 9362
rect 20875 7446 21075 8246
rect 21247 7446 21447 8246
rect 21619 7446 21819 8246
rect 21991 7446 22191 8246
rect 22363 7446 22563 8246
rect 22735 7446 22935 8246
rect 23107 7446 23307 8246
rect 23479 7446 23679 8246
rect 20875 6410 21075 7210
rect 21247 6410 21447 7210
rect 21619 6410 21819 7210
rect 21991 6410 22191 7210
rect 22363 6410 22563 7210
rect 22735 6410 22935 7210
rect 23107 6410 23307 7210
rect 23479 6410 23679 7210
rect 20875 5374 21075 6174
rect 21247 5374 21447 6174
rect 21619 5374 21819 6174
rect 21991 5374 22191 6174
rect 22363 5374 22563 6174
rect 22735 5374 22935 6174
rect 23107 5374 23307 6174
rect 23479 5374 23679 6174
rect 20875 4338 21075 5138
rect 21247 4338 21447 5138
rect 21619 4338 21819 5138
rect 21991 4338 22191 5138
rect 22363 4338 22563 5138
rect 22735 4338 22935 5138
rect 23107 4338 23307 5138
rect 23479 4338 23679 5138
<< nmoslvt >>
rect 20875 3361 21075 3561
rect 21247 3361 21447 3561
rect 21619 3361 21819 3561
rect 21991 3361 22191 3561
rect 22363 3361 22563 3561
rect 22735 3361 22935 3561
rect 23107 3361 23307 3561
rect 23479 3361 23679 3561
rect 23851 3361 24051 3561
rect 24223 3361 24423 3561
rect 24595 3361 24795 3561
rect 24967 3361 25167 3561
rect 25339 3361 25539 3561
rect 25711 3361 25911 3561
rect 26083 3361 26283 3561
rect 26455 3361 26655 3561
rect 26827 3361 27027 3561
rect 27199 3361 27399 3561
rect 27571 3361 27771 3561
rect 27943 3361 28143 3561
rect 28315 3361 28515 3561
rect 28687 3361 28887 3561
rect 29059 3361 29259 3561
rect 29431 3361 29631 3561
rect 20875 2943 21075 3143
rect 21247 2943 21447 3143
rect 21619 2943 21819 3143
rect 21991 2943 22191 3143
rect 22363 2943 22563 3143
rect 22735 2943 22935 3143
rect 23107 2943 23307 3143
rect 23479 2943 23679 3143
rect 23851 2943 24051 3143
rect 24223 2943 24423 3143
rect 24595 2943 24795 3143
rect 24967 2943 25167 3143
rect 25339 2943 25539 3143
rect 25711 2943 25911 3143
rect 26083 2943 26283 3143
rect 26455 2943 26655 3143
rect 26827 2943 27027 3143
rect 27199 2943 27399 3143
rect 27571 2943 27771 3143
rect 27943 2943 28143 3143
rect 28315 2943 28515 3143
rect 28687 2943 28887 3143
rect 29059 2943 29259 3143
rect 29431 2943 29631 3143
rect 20875 2525 21075 2725
rect 21247 2525 21447 2725
rect 21619 2525 21819 2725
rect 21991 2525 22191 2725
rect 22363 2525 22563 2725
rect 22735 2525 22935 2725
rect 23107 2525 23307 2725
rect 23479 2525 23679 2725
rect 23851 2525 24051 2725
rect 24223 2525 24423 2725
rect 24595 2525 24795 2725
rect 24967 2525 25167 2725
rect 25339 2525 25539 2725
rect 25711 2525 25911 2725
rect 26083 2525 26283 2725
rect 26455 2525 26655 2725
rect 26827 2525 27027 2725
rect 27199 2525 27399 2725
rect 27571 2525 27771 2725
rect 27943 2525 28143 2725
rect 28315 2525 28515 2725
rect 28687 2525 28887 2725
rect 29059 2525 29259 2725
rect 29431 2525 29631 2725
rect 20875 2107 21075 2307
rect 21247 2107 21447 2307
rect 21619 2107 21819 2307
rect 21991 2107 22191 2307
rect 22363 2107 22563 2307
rect 22735 2107 22935 2307
rect 23107 2107 23307 2307
rect 23479 2107 23679 2307
rect 23851 2107 24051 2307
rect 24223 2107 24423 2307
rect 24595 2107 24795 2307
rect 24967 2107 25167 2307
rect 25339 2107 25539 2307
rect 25711 2107 25911 2307
rect 26083 2107 26283 2307
rect 26455 2107 26655 2307
rect 26827 2107 27027 2307
rect 27199 2107 27399 2307
rect 27571 2107 27771 2307
rect 27943 2107 28143 2307
rect 28315 2107 28515 2307
rect 28687 2107 28887 2307
rect 29059 2107 29259 2307
rect 29431 2107 29631 2307
<< ndiff >>
rect 20817 3549 20875 3561
rect 20817 3373 20829 3549
rect 20863 3373 20875 3549
rect 20817 3361 20875 3373
rect 21075 3549 21133 3561
rect 21075 3373 21087 3549
rect 21121 3373 21133 3549
rect 21075 3361 21133 3373
rect 21189 3549 21247 3561
rect 21189 3373 21201 3549
rect 21235 3373 21247 3549
rect 21189 3361 21247 3373
rect 21447 3549 21505 3561
rect 21447 3373 21459 3549
rect 21493 3373 21505 3549
rect 21447 3361 21505 3373
rect 21561 3549 21619 3561
rect 21561 3373 21573 3549
rect 21607 3373 21619 3549
rect 21561 3361 21619 3373
rect 21819 3549 21877 3561
rect 21819 3373 21831 3549
rect 21865 3373 21877 3549
rect 21819 3361 21877 3373
rect 21933 3549 21991 3561
rect 21933 3373 21945 3549
rect 21979 3373 21991 3549
rect 21933 3361 21991 3373
rect 22191 3549 22249 3561
rect 22191 3373 22203 3549
rect 22237 3373 22249 3549
rect 22191 3361 22249 3373
rect 22305 3549 22363 3561
rect 22305 3373 22317 3549
rect 22351 3373 22363 3549
rect 22305 3361 22363 3373
rect 22563 3549 22621 3561
rect 22563 3373 22575 3549
rect 22609 3373 22621 3549
rect 22563 3361 22621 3373
rect 22677 3549 22735 3561
rect 22677 3373 22689 3549
rect 22723 3373 22735 3549
rect 22677 3361 22735 3373
rect 22935 3549 22993 3561
rect 22935 3373 22947 3549
rect 22981 3373 22993 3549
rect 22935 3361 22993 3373
rect 23049 3549 23107 3561
rect 23049 3373 23061 3549
rect 23095 3373 23107 3549
rect 23049 3361 23107 3373
rect 23307 3549 23365 3561
rect 23307 3373 23319 3549
rect 23353 3373 23365 3549
rect 23307 3361 23365 3373
rect 23421 3549 23479 3561
rect 23421 3373 23433 3549
rect 23467 3373 23479 3549
rect 23421 3361 23479 3373
rect 23679 3549 23737 3561
rect 23679 3373 23691 3549
rect 23725 3373 23737 3549
rect 23679 3361 23737 3373
rect 23793 3549 23851 3561
rect 23793 3373 23805 3549
rect 23839 3373 23851 3549
rect 23793 3361 23851 3373
rect 24051 3549 24109 3561
rect 24051 3373 24063 3549
rect 24097 3373 24109 3549
rect 24051 3361 24109 3373
rect 24165 3549 24223 3561
rect 24165 3373 24177 3549
rect 24211 3373 24223 3549
rect 24165 3361 24223 3373
rect 24423 3549 24481 3561
rect 24423 3373 24435 3549
rect 24469 3373 24481 3549
rect 24423 3361 24481 3373
rect 24537 3549 24595 3561
rect 24537 3373 24549 3549
rect 24583 3373 24595 3549
rect 24537 3361 24595 3373
rect 24795 3549 24853 3561
rect 24795 3373 24807 3549
rect 24841 3373 24853 3549
rect 24795 3361 24853 3373
rect 24909 3549 24967 3561
rect 24909 3373 24921 3549
rect 24955 3373 24967 3549
rect 24909 3361 24967 3373
rect 25167 3549 25225 3561
rect 25167 3373 25179 3549
rect 25213 3373 25225 3549
rect 25167 3361 25225 3373
rect 25281 3549 25339 3561
rect 25281 3373 25293 3549
rect 25327 3373 25339 3549
rect 25281 3361 25339 3373
rect 25539 3549 25597 3561
rect 25539 3373 25551 3549
rect 25585 3373 25597 3549
rect 25539 3361 25597 3373
rect 25653 3549 25711 3561
rect 25653 3373 25665 3549
rect 25699 3373 25711 3549
rect 25653 3361 25711 3373
rect 25911 3549 25969 3561
rect 25911 3373 25923 3549
rect 25957 3373 25969 3549
rect 25911 3361 25969 3373
rect 26025 3549 26083 3561
rect 26025 3373 26037 3549
rect 26071 3373 26083 3549
rect 26025 3361 26083 3373
rect 26283 3549 26341 3561
rect 26283 3373 26295 3549
rect 26329 3373 26341 3549
rect 26283 3361 26341 3373
rect 26397 3549 26455 3561
rect 26397 3373 26409 3549
rect 26443 3373 26455 3549
rect 26397 3361 26455 3373
rect 26655 3549 26713 3561
rect 26655 3373 26667 3549
rect 26701 3373 26713 3549
rect 26655 3361 26713 3373
rect 26769 3549 26827 3561
rect 26769 3373 26781 3549
rect 26815 3373 26827 3549
rect 26769 3361 26827 3373
rect 27027 3549 27085 3561
rect 27027 3373 27039 3549
rect 27073 3373 27085 3549
rect 27027 3361 27085 3373
rect 27141 3549 27199 3561
rect 27141 3373 27153 3549
rect 27187 3373 27199 3549
rect 27141 3361 27199 3373
rect 27399 3549 27457 3561
rect 27399 3373 27411 3549
rect 27445 3373 27457 3549
rect 27399 3361 27457 3373
rect 27513 3549 27571 3561
rect 27513 3373 27525 3549
rect 27559 3373 27571 3549
rect 27513 3361 27571 3373
rect 27771 3549 27829 3561
rect 27771 3373 27783 3549
rect 27817 3373 27829 3549
rect 27771 3361 27829 3373
rect 27885 3549 27943 3561
rect 27885 3373 27897 3549
rect 27931 3373 27943 3549
rect 27885 3361 27943 3373
rect 28143 3549 28201 3561
rect 28143 3373 28155 3549
rect 28189 3373 28201 3549
rect 28143 3361 28201 3373
rect 28257 3549 28315 3561
rect 28257 3373 28269 3549
rect 28303 3373 28315 3549
rect 28257 3361 28315 3373
rect 28515 3549 28573 3561
rect 28515 3373 28527 3549
rect 28561 3373 28573 3549
rect 28515 3361 28573 3373
rect 28629 3549 28687 3561
rect 28629 3373 28641 3549
rect 28675 3373 28687 3549
rect 28629 3361 28687 3373
rect 28887 3549 28945 3561
rect 28887 3373 28899 3549
rect 28933 3373 28945 3549
rect 28887 3361 28945 3373
rect 29001 3549 29059 3561
rect 29001 3373 29013 3549
rect 29047 3373 29059 3549
rect 29001 3361 29059 3373
rect 29259 3549 29317 3561
rect 29259 3373 29271 3549
rect 29305 3373 29317 3549
rect 29259 3361 29317 3373
rect 29373 3549 29431 3561
rect 29373 3373 29385 3549
rect 29419 3373 29431 3549
rect 29373 3361 29431 3373
rect 29631 3549 29689 3561
rect 29631 3373 29643 3549
rect 29677 3373 29689 3549
rect 29631 3361 29689 3373
rect 20817 3131 20875 3143
rect 20817 2955 20829 3131
rect 20863 2955 20875 3131
rect 20817 2943 20875 2955
rect 21075 3131 21133 3143
rect 21075 2955 21087 3131
rect 21121 2955 21133 3131
rect 21075 2943 21133 2955
rect 21189 3131 21247 3143
rect 21189 2955 21201 3131
rect 21235 2955 21247 3131
rect 21189 2943 21247 2955
rect 21447 3131 21505 3143
rect 21447 2955 21459 3131
rect 21493 2955 21505 3131
rect 21447 2943 21505 2955
rect 21561 3131 21619 3143
rect 21561 2955 21573 3131
rect 21607 2955 21619 3131
rect 21561 2943 21619 2955
rect 21819 3131 21877 3143
rect 21819 2955 21831 3131
rect 21865 2955 21877 3131
rect 21819 2943 21877 2955
rect 21933 3131 21991 3143
rect 21933 2955 21945 3131
rect 21979 2955 21991 3131
rect 21933 2943 21991 2955
rect 22191 3131 22249 3143
rect 22191 2955 22203 3131
rect 22237 2955 22249 3131
rect 22191 2943 22249 2955
rect 22305 3131 22363 3143
rect 22305 2955 22317 3131
rect 22351 2955 22363 3131
rect 22305 2943 22363 2955
rect 22563 3131 22621 3143
rect 22563 2955 22575 3131
rect 22609 2955 22621 3131
rect 22563 2943 22621 2955
rect 22677 3131 22735 3143
rect 22677 2955 22689 3131
rect 22723 2955 22735 3131
rect 22677 2943 22735 2955
rect 22935 3131 22993 3143
rect 22935 2955 22947 3131
rect 22981 2955 22993 3131
rect 22935 2943 22993 2955
rect 23049 3131 23107 3143
rect 23049 2955 23061 3131
rect 23095 2955 23107 3131
rect 23049 2943 23107 2955
rect 23307 3131 23365 3143
rect 23307 2955 23319 3131
rect 23353 2955 23365 3131
rect 23307 2943 23365 2955
rect 23421 3131 23479 3143
rect 23421 2955 23433 3131
rect 23467 2955 23479 3131
rect 23421 2943 23479 2955
rect 23679 3131 23737 3143
rect 23679 2955 23691 3131
rect 23725 2955 23737 3131
rect 23679 2943 23737 2955
rect 23793 3131 23851 3143
rect 23793 2955 23805 3131
rect 23839 2955 23851 3131
rect 23793 2943 23851 2955
rect 24051 3131 24109 3143
rect 24051 2955 24063 3131
rect 24097 2955 24109 3131
rect 24051 2943 24109 2955
rect 24165 3131 24223 3143
rect 24165 2955 24177 3131
rect 24211 2955 24223 3131
rect 24165 2943 24223 2955
rect 24423 3131 24481 3143
rect 24423 2955 24435 3131
rect 24469 2955 24481 3131
rect 24423 2943 24481 2955
rect 24537 3131 24595 3143
rect 24537 2955 24549 3131
rect 24583 2955 24595 3131
rect 24537 2943 24595 2955
rect 24795 3131 24853 3143
rect 24795 2955 24807 3131
rect 24841 2955 24853 3131
rect 24795 2943 24853 2955
rect 24909 3131 24967 3143
rect 24909 2955 24921 3131
rect 24955 2955 24967 3131
rect 24909 2943 24967 2955
rect 25167 3131 25225 3143
rect 25167 2955 25179 3131
rect 25213 2955 25225 3131
rect 25167 2943 25225 2955
rect 25281 3131 25339 3143
rect 25281 2955 25293 3131
rect 25327 2955 25339 3131
rect 25281 2943 25339 2955
rect 25539 3131 25597 3143
rect 25539 2955 25551 3131
rect 25585 2955 25597 3131
rect 25539 2943 25597 2955
rect 25653 3131 25711 3143
rect 25653 2955 25665 3131
rect 25699 2955 25711 3131
rect 25653 2943 25711 2955
rect 25911 3131 25969 3143
rect 25911 2955 25923 3131
rect 25957 2955 25969 3131
rect 25911 2943 25969 2955
rect 26025 3131 26083 3143
rect 26025 2955 26037 3131
rect 26071 2955 26083 3131
rect 26025 2943 26083 2955
rect 26283 3131 26341 3143
rect 26283 2955 26295 3131
rect 26329 2955 26341 3131
rect 26283 2943 26341 2955
rect 26397 3131 26455 3143
rect 26397 2955 26409 3131
rect 26443 2955 26455 3131
rect 26397 2943 26455 2955
rect 26655 3131 26713 3143
rect 26655 2955 26667 3131
rect 26701 2955 26713 3131
rect 26655 2943 26713 2955
rect 26769 3131 26827 3143
rect 26769 2955 26781 3131
rect 26815 2955 26827 3131
rect 26769 2943 26827 2955
rect 27027 3131 27085 3143
rect 27027 2955 27039 3131
rect 27073 2955 27085 3131
rect 27027 2943 27085 2955
rect 27141 3131 27199 3143
rect 27141 2955 27153 3131
rect 27187 2955 27199 3131
rect 27141 2943 27199 2955
rect 27399 3131 27457 3143
rect 27399 2955 27411 3131
rect 27445 2955 27457 3131
rect 27399 2943 27457 2955
rect 27513 3131 27571 3143
rect 27513 2955 27525 3131
rect 27559 2955 27571 3131
rect 27513 2943 27571 2955
rect 27771 3131 27829 3143
rect 27771 2955 27783 3131
rect 27817 2955 27829 3131
rect 27771 2943 27829 2955
rect 27885 3131 27943 3143
rect 27885 2955 27897 3131
rect 27931 2955 27943 3131
rect 27885 2943 27943 2955
rect 28143 3131 28201 3143
rect 28143 2955 28155 3131
rect 28189 2955 28201 3131
rect 28143 2943 28201 2955
rect 28257 3131 28315 3143
rect 28257 2955 28269 3131
rect 28303 2955 28315 3131
rect 28257 2943 28315 2955
rect 28515 3131 28573 3143
rect 28515 2955 28527 3131
rect 28561 2955 28573 3131
rect 28515 2943 28573 2955
rect 28629 3131 28687 3143
rect 28629 2955 28641 3131
rect 28675 2955 28687 3131
rect 28629 2943 28687 2955
rect 28887 3131 28945 3143
rect 28887 2955 28899 3131
rect 28933 2955 28945 3131
rect 28887 2943 28945 2955
rect 29001 3131 29059 3143
rect 29001 2955 29013 3131
rect 29047 2955 29059 3131
rect 29001 2943 29059 2955
rect 29259 3131 29317 3143
rect 29259 2955 29271 3131
rect 29305 2955 29317 3131
rect 29259 2943 29317 2955
rect 29373 3131 29431 3143
rect 29373 2955 29385 3131
rect 29419 2955 29431 3131
rect 29373 2943 29431 2955
rect 29631 3131 29689 3143
rect 29631 2955 29643 3131
rect 29677 2955 29689 3131
rect 29631 2943 29689 2955
rect 20817 2713 20875 2725
rect 20817 2537 20829 2713
rect 20863 2537 20875 2713
rect 20817 2525 20875 2537
rect 21075 2713 21133 2725
rect 21075 2537 21087 2713
rect 21121 2537 21133 2713
rect 21075 2525 21133 2537
rect 21189 2713 21247 2725
rect 21189 2537 21201 2713
rect 21235 2537 21247 2713
rect 21189 2525 21247 2537
rect 21447 2713 21505 2725
rect 21447 2537 21459 2713
rect 21493 2537 21505 2713
rect 21447 2525 21505 2537
rect 21561 2713 21619 2725
rect 21561 2537 21573 2713
rect 21607 2537 21619 2713
rect 21561 2525 21619 2537
rect 21819 2713 21877 2725
rect 21819 2537 21831 2713
rect 21865 2537 21877 2713
rect 21819 2525 21877 2537
rect 21933 2713 21991 2725
rect 21933 2537 21945 2713
rect 21979 2537 21991 2713
rect 21933 2525 21991 2537
rect 22191 2713 22249 2725
rect 22191 2537 22203 2713
rect 22237 2537 22249 2713
rect 22191 2525 22249 2537
rect 22305 2713 22363 2725
rect 22305 2537 22317 2713
rect 22351 2537 22363 2713
rect 22305 2525 22363 2537
rect 22563 2713 22621 2725
rect 22563 2537 22575 2713
rect 22609 2537 22621 2713
rect 22563 2525 22621 2537
rect 22677 2713 22735 2725
rect 22677 2537 22689 2713
rect 22723 2537 22735 2713
rect 22677 2525 22735 2537
rect 22935 2713 22993 2725
rect 22935 2537 22947 2713
rect 22981 2537 22993 2713
rect 22935 2525 22993 2537
rect 23049 2713 23107 2725
rect 23049 2537 23061 2713
rect 23095 2537 23107 2713
rect 23049 2525 23107 2537
rect 23307 2713 23365 2725
rect 23307 2537 23319 2713
rect 23353 2537 23365 2713
rect 23307 2525 23365 2537
rect 23421 2713 23479 2725
rect 23421 2537 23433 2713
rect 23467 2537 23479 2713
rect 23421 2525 23479 2537
rect 23679 2713 23737 2725
rect 23679 2537 23691 2713
rect 23725 2537 23737 2713
rect 23679 2525 23737 2537
rect 23793 2713 23851 2725
rect 23793 2537 23805 2713
rect 23839 2537 23851 2713
rect 23793 2525 23851 2537
rect 24051 2713 24109 2725
rect 24051 2537 24063 2713
rect 24097 2537 24109 2713
rect 24051 2525 24109 2537
rect 24165 2713 24223 2725
rect 24165 2537 24177 2713
rect 24211 2537 24223 2713
rect 24165 2525 24223 2537
rect 24423 2713 24481 2725
rect 24423 2537 24435 2713
rect 24469 2537 24481 2713
rect 24423 2525 24481 2537
rect 24537 2713 24595 2725
rect 24537 2537 24549 2713
rect 24583 2537 24595 2713
rect 24537 2525 24595 2537
rect 24795 2713 24853 2725
rect 24795 2537 24807 2713
rect 24841 2537 24853 2713
rect 24795 2525 24853 2537
rect 24909 2713 24967 2725
rect 24909 2537 24921 2713
rect 24955 2537 24967 2713
rect 24909 2525 24967 2537
rect 25167 2713 25225 2725
rect 25167 2537 25179 2713
rect 25213 2537 25225 2713
rect 25167 2525 25225 2537
rect 25281 2713 25339 2725
rect 25281 2537 25293 2713
rect 25327 2537 25339 2713
rect 25281 2525 25339 2537
rect 25539 2713 25597 2725
rect 25539 2537 25551 2713
rect 25585 2537 25597 2713
rect 25539 2525 25597 2537
rect 25653 2713 25711 2725
rect 25653 2537 25665 2713
rect 25699 2537 25711 2713
rect 25653 2525 25711 2537
rect 25911 2713 25969 2725
rect 25911 2537 25923 2713
rect 25957 2537 25969 2713
rect 25911 2525 25969 2537
rect 26025 2713 26083 2725
rect 26025 2537 26037 2713
rect 26071 2537 26083 2713
rect 26025 2525 26083 2537
rect 26283 2713 26341 2725
rect 26283 2537 26295 2713
rect 26329 2537 26341 2713
rect 26283 2525 26341 2537
rect 26397 2713 26455 2725
rect 26397 2537 26409 2713
rect 26443 2537 26455 2713
rect 26397 2525 26455 2537
rect 26655 2713 26713 2725
rect 26655 2537 26667 2713
rect 26701 2537 26713 2713
rect 26655 2525 26713 2537
rect 26769 2713 26827 2725
rect 26769 2537 26781 2713
rect 26815 2537 26827 2713
rect 26769 2525 26827 2537
rect 27027 2713 27085 2725
rect 27027 2537 27039 2713
rect 27073 2537 27085 2713
rect 27027 2525 27085 2537
rect 27141 2713 27199 2725
rect 27141 2537 27153 2713
rect 27187 2537 27199 2713
rect 27141 2525 27199 2537
rect 27399 2713 27457 2725
rect 27399 2537 27411 2713
rect 27445 2537 27457 2713
rect 27399 2525 27457 2537
rect 27513 2713 27571 2725
rect 27513 2537 27525 2713
rect 27559 2537 27571 2713
rect 27513 2525 27571 2537
rect 27771 2713 27829 2725
rect 27771 2537 27783 2713
rect 27817 2537 27829 2713
rect 27771 2525 27829 2537
rect 27885 2713 27943 2725
rect 27885 2537 27897 2713
rect 27931 2537 27943 2713
rect 27885 2525 27943 2537
rect 28143 2713 28201 2725
rect 28143 2537 28155 2713
rect 28189 2537 28201 2713
rect 28143 2525 28201 2537
rect 28257 2713 28315 2725
rect 28257 2537 28269 2713
rect 28303 2537 28315 2713
rect 28257 2525 28315 2537
rect 28515 2713 28573 2725
rect 28515 2537 28527 2713
rect 28561 2537 28573 2713
rect 28515 2525 28573 2537
rect 28629 2713 28687 2725
rect 28629 2537 28641 2713
rect 28675 2537 28687 2713
rect 28629 2525 28687 2537
rect 28887 2713 28945 2725
rect 28887 2537 28899 2713
rect 28933 2537 28945 2713
rect 28887 2525 28945 2537
rect 29001 2713 29059 2725
rect 29001 2537 29013 2713
rect 29047 2537 29059 2713
rect 29001 2525 29059 2537
rect 29259 2713 29317 2725
rect 29259 2537 29271 2713
rect 29305 2537 29317 2713
rect 29259 2525 29317 2537
rect 29373 2713 29431 2725
rect 29373 2537 29385 2713
rect 29419 2537 29431 2713
rect 29373 2525 29431 2537
rect 29631 2713 29689 2725
rect 29631 2537 29643 2713
rect 29677 2537 29689 2713
rect 29631 2525 29689 2537
rect 20817 2295 20875 2307
rect 20817 2119 20829 2295
rect 20863 2119 20875 2295
rect 20817 2107 20875 2119
rect 21075 2295 21133 2307
rect 21075 2119 21087 2295
rect 21121 2119 21133 2295
rect 21075 2107 21133 2119
rect 21189 2295 21247 2307
rect 21189 2119 21201 2295
rect 21235 2119 21247 2295
rect 21189 2107 21247 2119
rect 21447 2295 21505 2307
rect 21447 2119 21459 2295
rect 21493 2119 21505 2295
rect 21447 2107 21505 2119
rect 21561 2295 21619 2307
rect 21561 2119 21573 2295
rect 21607 2119 21619 2295
rect 21561 2107 21619 2119
rect 21819 2295 21877 2307
rect 21819 2119 21831 2295
rect 21865 2119 21877 2295
rect 21819 2107 21877 2119
rect 21933 2295 21991 2307
rect 21933 2119 21945 2295
rect 21979 2119 21991 2295
rect 21933 2107 21991 2119
rect 22191 2295 22249 2307
rect 22191 2119 22203 2295
rect 22237 2119 22249 2295
rect 22191 2107 22249 2119
rect 22305 2295 22363 2307
rect 22305 2119 22317 2295
rect 22351 2119 22363 2295
rect 22305 2107 22363 2119
rect 22563 2295 22621 2307
rect 22563 2119 22575 2295
rect 22609 2119 22621 2295
rect 22563 2107 22621 2119
rect 22677 2295 22735 2307
rect 22677 2119 22689 2295
rect 22723 2119 22735 2295
rect 22677 2107 22735 2119
rect 22935 2295 22993 2307
rect 22935 2119 22947 2295
rect 22981 2119 22993 2295
rect 22935 2107 22993 2119
rect 23049 2295 23107 2307
rect 23049 2119 23061 2295
rect 23095 2119 23107 2295
rect 23049 2107 23107 2119
rect 23307 2295 23365 2307
rect 23307 2119 23319 2295
rect 23353 2119 23365 2295
rect 23307 2107 23365 2119
rect 23421 2295 23479 2307
rect 23421 2119 23433 2295
rect 23467 2119 23479 2295
rect 23421 2107 23479 2119
rect 23679 2295 23737 2307
rect 23679 2119 23691 2295
rect 23725 2119 23737 2295
rect 23679 2107 23737 2119
rect 23793 2295 23851 2307
rect 23793 2119 23805 2295
rect 23839 2119 23851 2295
rect 23793 2107 23851 2119
rect 24051 2295 24109 2307
rect 24051 2119 24063 2295
rect 24097 2119 24109 2295
rect 24051 2107 24109 2119
rect 24165 2295 24223 2307
rect 24165 2119 24177 2295
rect 24211 2119 24223 2295
rect 24165 2107 24223 2119
rect 24423 2295 24481 2307
rect 24423 2119 24435 2295
rect 24469 2119 24481 2295
rect 24423 2107 24481 2119
rect 24537 2295 24595 2307
rect 24537 2119 24549 2295
rect 24583 2119 24595 2295
rect 24537 2107 24595 2119
rect 24795 2295 24853 2307
rect 24795 2119 24807 2295
rect 24841 2119 24853 2295
rect 24795 2107 24853 2119
rect 24909 2295 24967 2307
rect 24909 2119 24921 2295
rect 24955 2119 24967 2295
rect 24909 2107 24967 2119
rect 25167 2295 25225 2307
rect 25167 2119 25179 2295
rect 25213 2119 25225 2295
rect 25167 2107 25225 2119
rect 25281 2295 25339 2307
rect 25281 2119 25293 2295
rect 25327 2119 25339 2295
rect 25281 2107 25339 2119
rect 25539 2295 25597 2307
rect 25539 2119 25551 2295
rect 25585 2119 25597 2295
rect 25539 2107 25597 2119
rect 25653 2295 25711 2307
rect 25653 2119 25665 2295
rect 25699 2119 25711 2295
rect 25653 2107 25711 2119
rect 25911 2295 25969 2307
rect 25911 2119 25923 2295
rect 25957 2119 25969 2295
rect 25911 2107 25969 2119
rect 26025 2295 26083 2307
rect 26025 2119 26037 2295
rect 26071 2119 26083 2295
rect 26025 2107 26083 2119
rect 26283 2295 26341 2307
rect 26283 2119 26295 2295
rect 26329 2119 26341 2295
rect 26283 2107 26341 2119
rect 26397 2295 26455 2307
rect 26397 2119 26409 2295
rect 26443 2119 26455 2295
rect 26397 2107 26455 2119
rect 26655 2295 26713 2307
rect 26655 2119 26667 2295
rect 26701 2119 26713 2295
rect 26655 2107 26713 2119
rect 26769 2295 26827 2307
rect 26769 2119 26781 2295
rect 26815 2119 26827 2295
rect 26769 2107 26827 2119
rect 27027 2295 27085 2307
rect 27027 2119 27039 2295
rect 27073 2119 27085 2295
rect 27027 2107 27085 2119
rect 27141 2295 27199 2307
rect 27141 2119 27153 2295
rect 27187 2119 27199 2295
rect 27141 2107 27199 2119
rect 27399 2295 27457 2307
rect 27399 2119 27411 2295
rect 27445 2119 27457 2295
rect 27399 2107 27457 2119
rect 27513 2295 27571 2307
rect 27513 2119 27525 2295
rect 27559 2119 27571 2295
rect 27513 2107 27571 2119
rect 27771 2295 27829 2307
rect 27771 2119 27783 2295
rect 27817 2119 27829 2295
rect 27771 2107 27829 2119
rect 27885 2295 27943 2307
rect 27885 2119 27897 2295
rect 27931 2119 27943 2295
rect 27885 2107 27943 2119
rect 28143 2295 28201 2307
rect 28143 2119 28155 2295
rect 28189 2119 28201 2295
rect 28143 2107 28201 2119
rect 28257 2295 28315 2307
rect 28257 2119 28269 2295
rect 28303 2119 28315 2295
rect 28257 2107 28315 2119
rect 28515 2295 28573 2307
rect 28515 2119 28527 2295
rect 28561 2119 28573 2295
rect 28515 2107 28573 2119
rect 28629 2295 28687 2307
rect 28629 2119 28641 2295
rect 28675 2119 28687 2295
rect 28629 2107 28687 2119
rect 28887 2295 28945 2307
rect 28887 2119 28899 2295
rect 28933 2119 28945 2295
rect 28887 2107 28945 2119
rect 29001 2295 29059 2307
rect 29001 2119 29013 2295
rect 29047 2119 29059 2295
rect 29001 2107 29059 2119
rect 29259 2295 29317 2307
rect 29259 2119 29271 2295
rect 29305 2119 29317 2295
rect 29259 2107 29317 2119
rect 29373 2295 29431 2307
rect 29373 2119 29385 2295
rect 29419 2119 29431 2295
rect 29373 2107 29431 2119
rect 29631 2295 29689 2307
rect 29631 2119 29643 2295
rect 29677 2119 29689 2295
rect 29631 2107 29689 2119
<< pdiff >>
rect 19329 10622 19387 10634
rect 19329 10246 19341 10622
rect 19375 10246 19387 10622
rect 19329 10234 19387 10246
rect 19587 10622 19645 10634
rect 19587 10246 19599 10622
rect 19633 10246 19645 10622
rect 19587 10234 19645 10246
rect 19701 10622 19759 10634
rect 19701 10246 19713 10622
rect 19747 10246 19759 10622
rect 19701 10234 19759 10246
rect 19959 10622 20017 10634
rect 19959 10246 19971 10622
rect 20005 10246 20017 10622
rect 19959 10234 20017 10246
rect 20073 10622 20131 10634
rect 20073 10246 20085 10622
rect 20119 10246 20131 10622
rect 20073 10234 20131 10246
rect 20331 10622 20389 10634
rect 20331 10246 20343 10622
rect 20377 10246 20389 10622
rect 20331 10234 20389 10246
rect 20445 10622 20503 10634
rect 20445 10246 20457 10622
rect 20491 10246 20503 10622
rect 20445 10234 20503 10246
rect 20703 10622 20761 10634
rect 20703 10246 20715 10622
rect 20749 10246 20761 10622
rect 20703 10234 20761 10246
rect 20817 10622 20875 10634
rect 20817 10246 20829 10622
rect 20863 10246 20875 10622
rect 20817 10234 20875 10246
rect 21075 10622 21133 10634
rect 21075 10246 21087 10622
rect 21121 10246 21133 10622
rect 21075 10234 21133 10246
rect 21189 10622 21247 10634
rect 21189 10246 21201 10622
rect 21235 10246 21247 10622
rect 21189 10234 21247 10246
rect 21447 10622 21505 10634
rect 21447 10246 21459 10622
rect 21493 10246 21505 10622
rect 21447 10234 21505 10246
rect 21561 10622 21619 10634
rect 21561 10246 21573 10622
rect 21607 10246 21619 10622
rect 21561 10234 21619 10246
rect 21819 10622 21877 10634
rect 21819 10246 21831 10622
rect 21865 10246 21877 10622
rect 21819 10234 21877 10246
rect 21933 10622 21991 10634
rect 21933 10246 21945 10622
rect 21979 10246 21991 10622
rect 21933 10234 21991 10246
rect 22191 10622 22249 10634
rect 22191 10246 22203 10622
rect 22237 10246 22249 10622
rect 22191 10234 22249 10246
rect 22305 10622 22363 10634
rect 22305 10246 22317 10622
rect 22351 10246 22363 10622
rect 22305 10234 22363 10246
rect 22563 10622 22621 10634
rect 22563 10246 22575 10622
rect 22609 10246 22621 10622
rect 22563 10234 22621 10246
rect 22677 10622 22735 10634
rect 22677 10246 22689 10622
rect 22723 10246 22735 10622
rect 22677 10234 22735 10246
rect 22935 10622 22993 10634
rect 22935 10246 22947 10622
rect 22981 10246 22993 10622
rect 22935 10234 22993 10246
rect 23049 10622 23107 10634
rect 23049 10246 23061 10622
rect 23095 10246 23107 10622
rect 23049 10234 23107 10246
rect 23307 10622 23365 10634
rect 23307 10246 23319 10622
rect 23353 10246 23365 10622
rect 23307 10234 23365 10246
rect 23421 10622 23479 10634
rect 23421 10246 23433 10622
rect 23467 10246 23479 10622
rect 23421 10234 23479 10246
rect 23679 10622 23737 10634
rect 23679 10246 23691 10622
rect 23725 10246 23737 10622
rect 23679 10234 23737 10246
rect 23793 10622 23851 10634
rect 23793 10246 23805 10622
rect 23839 10246 23851 10622
rect 23793 10234 23851 10246
rect 24051 10622 24109 10634
rect 24051 10246 24063 10622
rect 24097 10246 24109 10622
rect 24051 10234 24109 10246
rect 24165 10622 24223 10634
rect 24165 10246 24177 10622
rect 24211 10246 24223 10622
rect 24165 10234 24223 10246
rect 24423 10622 24481 10634
rect 24423 10246 24435 10622
rect 24469 10246 24481 10622
rect 24423 10234 24481 10246
rect 24537 10622 24595 10634
rect 24537 10246 24549 10622
rect 24583 10246 24595 10622
rect 24537 10234 24595 10246
rect 24795 10622 24853 10634
rect 24795 10246 24807 10622
rect 24841 10246 24853 10622
rect 24795 10234 24853 10246
rect 24909 10622 24967 10634
rect 24909 10246 24921 10622
rect 24955 10246 24967 10622
rect 24909 10234 24967 10246
rect 25167 10622 25225 10634
rect 25167 10246 25179 10622
rect 25213 10246 25225 10622
rect 25167 10234 25225 10246
rect 25281 10622 25339 10634
rect 25281 10246 25293 10622
rect 25327 10246 25339 10622
rect 25281 10234 25339 10246
rect 25539 10622 25597 10634
rect 25539 10246 25551 10622
rect 25585 10246 25597 10622
rect 25539 10234 25597 10246
rect 25653 10622 25711 10634
rect 25653 10246 25665 10622
rect 25699 10246 25711 10622
rect 25653 10234 25711 10246
rect 25911 10622 25969 10634
rect 25911 10246 25923 10622
rect 25957 10246 25969 10622
rect 25911 10234 25969 10246
rect 26025 10622 26083 10634
rect 26025 10246 26037 10622
rect 26071 10246 26083 10622
rect 26025 10234 26083 10246
rect 26283 10622 26341 10634
rect 26283 10246 26295 10622
rect 26329 10246 26341 10622
rect 26283 10234 26341 10246
rect 26397 10622 26455 10634
rect 26397 10246 26409 10622
rect 26443 10246 26455 10622
rect 26397 10234 26455 10246
rect 26655 10622 26713 10634
rect 26655 10246 26667 10622
rect 26701 10246 26713 10622
rect 26655 10234 26713 10246
rect 26769 10622 26827 10634
rect 26769 10246 26781 10622
rect 26815 10246 26827 10622
rect 26769 10234 26827 10246
rect 27027 10622 27085 10634
rect 27027 10246 27039 10622
rect 27073 10246 27085 10622
rect 27027 10234 27085 10246
rect 27141 10622 27199 10634
rect 27141 10246 27153 10622
rect 27187 10246 27199 10622
rect 27141 10234 27199 10246
rect 27399 10622 27457 10634
rect 27399 10246 27411 10622
rect 27445 10246 27457 10622
rect 27399 10234 27457 10246
rect 27513 10622 27571 10634
rect 27513 10246 27525 10622
rect 27559 10246 27571 10622
rect 27513 10234 27571 10246
rect 27771 10622 27829 10634
rect 27771 10246 27783 10622
rect 27817 10246 27829 10622
rect 27771 10234 27829 10246
rect 27885 10622 27943 10634
rect 27885 10246 27897 10622
rect 27931 10246 27943 10622
rect 27885 10234 27943 10246
rect 28143 10622 28201 10634
rect 28143 10246 28155 10622
rect 28189 10246 28201 10622
rect 28143 10234 28201 10246
rect 28257 10622 28315 10634
rect 28257 10246 28269 10622
rect 28303 10246 28315 10622
rect 28257 10234 28315 10246
rect 28515 10622 28573 10634
rect 28515 10246 28527 10622
rect 28561 10246 28573 10622
rect 28515 10234 28573 10246
rect 28629 10622 28687 10634
rect 28629 10246 28641 10622
rect 28675 10246 28687 10622
rect 28629 10234 28687 10246
rect 28887 10622 28945 10634
rect 28887 10246 28899 10622
rect 28933 10246 28945 10622
rect 28887 10234 28945 10246
rect 29001 10622 29059 10634
rect 29001 10246 29013 10622
rect 29047 10246 29059 10622
rect 29001 10234 29059 10246
rect 29259 10622 29317 10634
rect 29259 10246 29271 10622
rect 29305 10246 29317 10622
rect 29259 10234 29317 10246
rect 29373 10622 29431 10634
rect 29373 10246 29385 10622
rect 29419 10246 29431 10622
rect 29373 10234 29431 10246
rect 29631 10622 29689 10634
rect 29631 10246 29643 10622
rect 29677 10246 29689 10622
rect 29631 10234 29689 10246
rect 29745 10622 29803 10634
rect 29745 10246 29757 10622
rect 29791 10246 29803 10622
rect 29745 10234 29803 10246
rect 30003 10622 30061 10634
rect 30003 10246 30015 10622
rect 30049 10246 30061 10622
rect 30003 10234 30061 10246
rect 30117 10622 30175 10634
rect 30117 10246 30129 10622
rect 30163 10246 30175 10622
rect 30117 10234 30175 10246
rect 30375 10622 30433 10634
rect 30375 10246 30387 10622
rect 30421 10246 30433 10622
rect 30375 10234 30433 10246
rect 30489 10622 30547 10634
rect 30489 10246 30501 10622
rect 30535 10246 30547 10622
rect 30489 10234 30547 10246
rect 30747 10622 30805 10634
rect 30747 10246 30759 10622
rect 30793 10246 30805 10622
rect 30747 10234 30805 10246
rect 30861 10622 30919 10634
rect 30861 10246 30873 10622
rect 30907 10246 30919 10622
rect 30861 10234 30919 10246
rect 31119 10622 31177 10634
rect 31119 10246 31131 10622
rect 31165 10246 31177 10622
rect 31119 10234 31177 10246
rect 19329 9986 19387 9998
rect 19329 9610 19341 9986
rect 19375 9610 19387 9986
rect 19329 9598 19387 9610
rect 19587 9986 19645 9998
rect 19587 9610 19599 9986
rect 19633 9610 19645 9986
rect 19587 9598 19645 9610
rect 19701 9986 19759 9998
rect 19701 9610 19713 9986
rect 19747 9610 19759 9986
rect 19701 9598 19759 9610
rect 19959 9986 20017 9998
rect 19959 9610 19971 9986
rect 20005 9610 20017 9986
rect 19959 9598 20017 9610
rect 20073 9986 20131 9998
rect 20073 9610 20085 9986
rect 20119 9610 20131 9986
rect 20073 9598 20131 9610
rect 20331 9986 20389 9998
rect 20331 9610 20343 9986
rect 20377 9610 20389 9986
rect 20331 9598 20389 9610
rect 20445 9986 20503 9998
rect 20445 9610 20457 9986
rect 20491 9610 20503 9986
rect 20445 9598 20503 9610
rect 20703 9986 20761 9998
rect 20703 9610 20715 9986
rect 20749 9610 20761 9986
rect 20703 9598 20761 9610
rect 20817 9986 20875 9998
rect 20817 9610 20829 9986
rect 20863 9610 20875 9986
rect 20817 9598 20875 9610
rect 21075 9986 21133 9998
rect 21075 9610 21087 9986
rect 21121 9610 21133 9986
rect 21075 9598 21133 9610
rect 21189 9986 21247 9998
rect 21189 9610 21201 9986
rect 21235 9610 21247 9986
rect 21189 9598 21247 9610
rect 21447 9986 21505 9998
rect 21447 9610 21459 9986
rect 21493 9610 21505 9986
rect 21447 9598 21505 9610
rect 21561 9986 21619 9998
rect 21561 9610 21573 9986
rect 21607 9610 21619 9986
rect 21561 9598 21619 9610
rect 21819 9986 21877 9998
rect 21819 9610 21831 9986
rect 21865 9610 21877 9986
rect 21819 9598 21877 9610
rect 21933 9986 21991 9998
rect 21933 9610 21945 9986
rect 21979 9610 21991 9986
rect 21933 9598 21991 9610
rect 22191 9986 22249 9998
rect 22191 9610 22203 9986
rect 22237 9610 22249 9986
rect 22191 9598 22249 9610
rect 22305 9986 22363 9998
rect 22305 9610 22317 9986
rect 22351 9610 22363 9986
rect 22305 9598 22363 9610
rect 22563 9986 22621 9998
rect 22563 9610 22575 9986
rect 22609 9610 22621 9986
rect 22563 9598 22621 9610
rect 22677 9986 22735 9998
rect 22677 9610 22689 9986
rect 22723 9610 22735 9986
rect 22677 9598 22735 9610
rect 22935 9986 22993 9998
rect 22935 9610 22947 9986
rect 22981 9610 22993 9986
rect 22935 9598 22993 9610
rect 23049 9986 23107 9998
rect 23049 9610 23061 9986
rect 23095 9610 23107 9986
rect 23049 9598 23107 9610
rect 23307 9986 23365 9998
rect 23307 9610 23319 9986
rect 23353 9610 23365 9986
rect 23307 9598 23365 9610
rect 23421 9986 23479 9998
rect 23421 9610 23433 9986
rect 23467 9610 23479 9986
rect 23421 9598 23479 9610
rect 23679 9986 23737 9998
rect 23679 9610 23691 9986
rect 23725 9610 23737 9986
rect 23679 9598 23737 9610
rect 23793 9986 23851 9998
rect 23793 9610 23805 9986
rect 23839 9610 23851 9986
rect 23793 9598 23851 9610
rect 24051 9986 24109 9998
rect 24051 9610 24063 9986
rect 24097 9610 24109 9986
rect 24051 9598 24109 9610
rect 24165 9986 24223 9998
rect 24165 9610 24177 9986
rect 24211 9610 24223 9986
rect 24165 9598 24223 9610
rect 24423 9986 24481 9998
rect 24423 9610 24435 9986
rect 24469 9610 24481 9986
rect 24423 9598 24481 9610
rect 24537 9986 24595 9998
rect 24537 9610 24549 9986
rect 24583 9610 24595 9986
rect 24537 9598 24595 9610
rect 24795 9986 24853 9998
rect 24795 9610 24807 9986
rect 24841 9610 24853 9986
rect 24795 9598 24853 9610
rect 24909 9986 24967 9998
rect 24909 9610 24921 9986
rect 24955 9610 24967 9986
rect 24909 9598 24967 9610
rect 25167 9986 25225 9998
rect 25167 9610 25179 9986
rect 25213 9610 25225 9986
rect 25167 9598 25225 9610
rect 25281 9986 25339 9998
rect 25281 9610 25293 9986
rect 25327 9610 25339 9986
rect 25281 9598 25339 9610
rect 25539 9986 25597 9998
rect 25539 9610 25551 9986
rect 25585 9610 25597 9986
rect 25539 9598 25597 9610
rect 25653 9986 25711 9998
rect 25653 9610 25665 9986
rect 25699 9610 25711 9986
rect 25653 9598 25711 9610
rect 25911 9986 25969 9998
rect 25911 9610 25923 9986
rect 25957 9610 25969 9986
rect 25911 9598 25969 9610
rect 26025 9986 26083 9998
rect 26025 9610 26037 9986
rect 26071 9610 26083 9986
rect 26025 9598 26083 9610
rect 26283 9986 26341 9998
rect 26283 9610 26295 9986
rect 26329 9610 26341 9986
rect 26283 9598 26341 9610
rect 26397 9986 26455 9998
rect 26397 9610 26409 9986
rect 26443 9610 26455 9986
rect 26397 9598 26455 9610
rect 26655 9986 26713 9998
rect 26655 9610 26667 9986
rect 26701 9610 26713 9986
rect 26655 9598 26713 9610
rect 26769 9986 26827 9998
rect 26769 9610 26781 9986
rect 26815 9610 26827 9986
rect 26769 9598 26827 9610
rect 27027 9986 27085 9998
rect 27027 9610 27039 9986
rect 27073 9610 27085 9986
rect 27027 9598 27085 9610
rect 27141 9986 27199 9998
rect 27141 9610 27153 9986
rect 27187 9610 27199 9986
rect 27141 9598 27199 9610
rect 27399 9986 27457 9998
rect 27399 9610 27411 9986
rect 27445 9610 27457 9986
rect 27399 9598 27457 9610
rect 27513 9986 27571 9998
rect 27513 9610 27525 9986
rect 27559 9610 27571 9986
rect 27513 9598 27571 9610
rect 27771 9986 27829 9998
rect 27771 9610 27783 9986
rect 27817 9610 27829 9986
rect 27771 9598 27829 9610
rect 27885 9986 27943 9998
rect 27885 9610 27897 9986
rect 27931 9610 27943 9986
rect 27885 9598 27943 9610
rect 28143 9986 28201 9998
rect 28143 9610 28155 9986
rect 28189 9610 28201 9986
rect 28143 9598 28201 9610
rect 28257 9986 28315 9998
rect 28257 9610 28269 9986
rect 28303 9610 28315 9986
rect 28257 9598 28315 9610
rect 28515 9986 28573 9998
rect 28515 9610 28527 9986
rect 28561 9610 28573 9986
rect 28515 9598 28573 9610
rect 28629 9986 28687 9998
rect 28629 9610 28641 9986
rect 28675 9610 28687 9986
rect 28629 9598 28687 9610
rect 28887 9986 28945 9998
rect 28887 9610 28899 9986
rect 28933 9610 28945 9986
rect 28887 9598 28945 9610
rect 29001 9986 29059 9998
rect 29001 9610 29013 9986
rect 29047 9610 29059 9986
rect 29001 9598 29059 9610
rect 29259 9986 29317 9998
rect 29259 9610 29271 9986
rect 29305 9610 29317 9986
rect 29259 9598 29317 9610
rect 29373 9986 29431 9998
rect 29373 9610 29385 9986
rect 29419 9610 29431 9986
rect 29373 9598 29431 9610
rect 29631 9986 29689 9998
rect 29631 9610 29643 9986
rect 29677 9610 29689 9986
rect 29631 9598 29689 9610
rect 29745 9986 29803 9998
rect 29745 9610 29757 9986
rect 29791 9610 29803 9986
rect 29745 9598 29803 9610
rect 30003 9986 30061 9998
rect 30003 9610 30015 9986
rect 30049 9610 30061 9986
rect 30003 9598 30061 9610
rect 30117 9986 30175 9998
rect 30117 9610 30129 9986
rect 30163 9610 30175 9986
rect 30117 9598 30175 9610
rect 30375 9986 30433 9998
rect 30375 9610 30387 9986
rect 30421 9610 30433 9986
rect 30375 9598 30433 9610
rect 30489 9986 30547 9998
rect 30489 9610 30501 9986
rect 30535 9610 30547 9986
rect 30489 9598 30547 9610
rect 30747 9986 30805 9998
rect 30747 9610 30759 9986
rect 30793 9610 30805 9986
rect 30747 9598 30805 9610
rect 30861 9986 30919 9998
rect 30861 9610 30873 9986
rect 30907 9610 30919 9986
rect 30861 9598 30919 9610
rect 31119 9986 31177 9998
rect 31119 9610 31131 9986
rect 31165 9610 31177 9986
rect 31119 9598 31177 9610
rect 19329 9350 19387 9362
rect 19329 8974 19341 9350
rect 19375 8974 19387 9350
rect 19329 8962 19387 8974
rect 19587 9350 19645 9362
rect 19587 8974 19599 9350
rect 19633 8974 19645 9350
rect 19587 8962 19645 8974
rect 19701 9350 19759 9362
rect 19701 8974 19713 9350
rect 19747 8974 19759 9350
rect 19701 8962 19759 8974
rect 19959 9350 20017 9362
rect 19959 8974 19971 9350
rect 20005 8974 20017 9350
rect 19959 8962 20017 8974
rect 20073 9350 20131 9362
rect 20073 8974 20085 9350
rect 20119 8974 20131 9350
rect 20073 8962 20131 8974
rect 20331 9350 20389 9362
rect 20331 8974 20343 9350
rect 20377 8974 20389 9350
rect 20331 8962 20389 8974
rect 20445 9350 20503 9362
rect 20445 8974 20457 9350
rect 20491 8974 20503 9350
rect 20445 8962 20503 8974
rect 20703 9350 20761 9362
rect 20703 8974 20715 9350
rect 20749 8974 20761 9350
rect 20703 8962 20761 8974
rect 20817 9350 20875 9362
rect 20817 8974 20829 9350
rect 20863 8974 20875 9350
rect 20817 8962 20875 8974
rect 21075 9350 21133 9362
rect 21075 8974 21087 9350
rect 21121 8974 21133 9350
rect 21075 8962 21133 8974
rect 21189 9350 21247 9362
rect 21189 8974 21201 9350
rect 21235 8974 21247 9350
rect 21189 8962 21247 8974
rect 21447 9350 21505 9362
rect 21447 8974 21459 9350
rect 21493 8974 21505 9350
rect 21447 8962 21505 8974
rect 21561 9350 21619 9362
rect 21561 8974 21573 9350
rect 21607 8974 21619 9350
rect 21561 8962 21619 8974
rect 21819 9350 21877 9362
rect 21819 8974 21831 9350
rect 21865 8974 21877 9350
rect 21819 8962 21877 8974
rect 21933 9350 21991 9362
rect 21933 8974 21945 9350
rect 21979 8974 21991 9350
rect 21933 8962 21991 8974
rect 22191 9350 22249 9362
rect 22191 8974 22203 9350
rect 22237 8974 22249 9350
rect 22191 8962 22249 8974
rect 22305 9350 22363 9362
rect 22305 8974 22317 9350
rect 22351 8974 22363 9350
rect 22305 8962 22363 8974
rect 22563 9350 22621 9362
rect 22563 8974 22575 9350
rect 22609 8974 22621 9350
rect 22563 8962 22621 8974
rect 22677 9350 22735 9362
rect 22677 8974 22689 9350
rect 22723 8974 22735 9350
rect 22677 8962 22735 8974
rect 22935 9350 22993 9362
rect 22935 8974 22947 9350
rect 22981 8974 22993 9350
rect 22935 8962 22993 8974
rect 23049 9350 23107 9362
rect 23049 8974 23061 9350
rect 23095 8974 23107 9350
rect 23049 8962 23107 8974
rect 23307 9350 23365 9362
rect 23307 8974 23319 9350
rect 23353 8974 23365 9350
rect 23307 8962 23365 8974
rect 23421 9350 23479 9362
rect 23421 8974 23433 9350
rect 23467 8974 23479 9350
rect 23421 8962 23479 8974
rect 23679 9350 23737 9362
rect 23679 8974 23691 9350
rect 23725 8974 23737 9350
rect 23679 8962 23737 8974
rect 23793 9350 23851 9362
rect 23793 8974 23805 9350
rect 23839 8974 23851 9350
rect 23793 8962 23851 8974
rect 24051 9350 24109 9362
rect 24051 8974 24063 9350
rect 24097 8974 24109 9350
rect 24051 8962 24109 8974
rect 24165 9350 24223 9362
rect 24165 8974 24177 9350
rect 24211 8974 24223 9350
rect 24165 8962 24223 8974
rect 24423 9350 24481 9362
rect 24423 8974 24435 9350
rect 24469 8974 24481 9350
rect 24423 8962 24481 8974
rect 24537 9350 24595 9362
rect 24537 8974 24549 9350
rect 24583 8974 24595 9350
rect 24537 8962 24595 8974
rect 24795 9350 24853 9362
rect 24795 8974 24807 9350
rect 24841 8974 24853 9350
rect 24795 8962 24853 8974
rect 24909 9350 24967 9362
rect 24909 8974 24921 9350
rect 24955 8974 24967 9350
rect 24909 8962 24967 8974
rect 25167 9350 25225 9362
rect 25167 8974 25179 9350
rect 25213 8974 25225 9350
rect 25167 8962 25225 8974
rect 25281 9350 25339 9362
rect 25281 8974 25293 9350
rect 25327 8974 25339 9350
rect 25281 8962 25339 8974
rect 25539 9350 25597 9362
rect 25539 8974 25551 9350
rect 25585 8974 25597 9350
rect 25539 8962 25597 8974
rect 25653 9350 25711 9362
rect 25653 8974 25665 9350
rect 25699 8974 25711 9350
rect 25653 8962 25711 8974
rect 25911 9350 25969 9362
rect 25911 8974 25923 9350
rect 25957 8974 25969 9350
rect 25911 8962 25969 8974
rect 26025 9350 26083 9362
rect 26025 8974 26037 9350
rect 26071 8974 26083 9350
rect 26025 8962 26083 8974
rect 26283 9350 26341 9362
rect 26283 8974 26295 9350
rect 26329 8974 26341 9350
rect 26283 8962 26341 8974
rect 26397 9350 26455 9362
rect 26397 8974 26409 9350
rect 26443 8974 26455 9350
rect 26397 8962 26455 8974
rect 26655 9350 26713 9362
rect 26655 8974 26667 9350
rect 26701 8974 26713 9350
rect 26655 8962 26713 8974
rect 26769 9350 26827 9362
rect 26769 8974 26781 9350
rect 26815 8974 26827 9350
rect 26769 8962 26827 8974
rect 27027 9350 27085 9362
rect 27027 8974 27039 9350
rect 27073 8974 27085 9350
rect 27027 8962 27085 8974
rect 27141 9350 27199 9362
rect 27141 8974 27153 9350
rect 27187 8974 27199 9350
rect 27141 8962 27199 8974
rect 27399 9350 27457 9362
rect 27399 8974 27411 9350
rect 27445 8974 27457 9350
rect 27399 8962 27457 8974
rect 27513 9350 27571 9362
rect 27513 8974 27525 9350
rect 27559 8974 27571 9350
rect 27513 8962 27571 8974
rect 27771 9350 27829 9362
rect 27771 8974 27783 9350
rect 27817 8974 27829 9350
rect 27771 8962 27829 8974
rect 27885 9350 27943 9362
rect 27885 8974 27897 9350
rect 27931 8974 27943 9350
rect 27885 8962 27943 8974
rect 28143 9350 28201 9362
rect 28143 8974 28155 9350
rect 28189 8974 28201 9350
rect 28143 8962 28201 8974
rect 28257 9350 28315 9362
rect 28257 8974 28269 9350
rect 28303 8974 28315 9350
rect 28257 8962 28315 8974
rect 28515 9350 28573 9362
rect 28515 8974 28527 9350
rect 28561 8974 28573 9350
rect 28515 8962 28573 8974
rect 28629 9350 28687 9362
rect 28629 8974 28641 9350
rect 28675 8974 28687 9350
rect 28629 8962 28687 8974
rect 28887 9350 28945 9362
rect 28887 8974 28899 9350
rect 28933 8974 28945 9350
rect 28887 8962 28945 8974
rect 29001 9350 29059 9362
rect 29001 8974 29013 9350
rect 29047 8974 29059 9350
rect 29001 8962 29059 8974
rect 29259 9350 29317 9362
rect 29259 8974 29271 9350
rect 29305 8974 29317 9350
rect 29259 8962 29317 8974
rect 29373 9350 29431 9362
rect 29373 8974 29385 9350
rect 29419 8974 29431 9350
rect 29373 8962 29431 8974
rect 29631 9350 29689 9362
rect 29631 8974 29643 9350
rect 29677 8974 29689 9350
rect 29631 8962 29689 8974
rect 29745 9350 29803 9362
rect 29745 8974 29757 9350
rect 29791 8974 29803 9350
rect 29745 8962 29803 8974
rect 30003 9350 30061 9362
rect 30003 8974 30015 9350
rect 30049 8974 30061 9350
rect 30003 8962 30061 8974
rect 30117 9350 30175 9362
rect 30117 8974 30129 9350
rect 30163 8974 30175 9350
rect 30117 8962 30175 8974
rect 30375 9350 30433 9362
rect 30375 8974 30387 9350
rect 30421 8974 30433 9350
rect 30375 8962 30433 8974
rect 30489 9350 30547 9362
rect 30489 8974 30501 9350
rect 30535 8974 30547 9350
rect 30489 8962 30547 8974
rect 30747 9350 30805 9362
rect 30747 8974 30759 9350
rect 30793 8974 30805 9350
rect 30747 8962 30805 8974
rect 30861 9350 30919 9362
rect 30861 8974 30873 9350
rect 30907 8974 30919 9350
rect 30861 8962 30919 8974
rect 31119 9350 31177 9362
rect 31119 8974 31131 9350
rect 31165 8974 31177 9350
rect 31119 8962 31177 8974
rect 20817 8234 20875 8246
rect 20817 7458 20829 8234
rect 20863 7458 20875 8234
rect 20817 7446 20875 7458
rect 21075 8234 21133 8246
rect 21075 7458 21087 8234
rect 21121 7458 21133 8234
rect 21075 7446 21133 7458
rect 21189 8234 21247 8246
rect 21189 7458 21201 8234
rect 21235 7458 21247 8234
rect 21189 7446 21247 7458
rect 21447 8234 21505 8246
rect 21447 7458 21459 8234
rect 21493 7458 21505 8234
rect 21447 7446 21505 7458
rect 21561 8234 21619 8246
rect 21561 7458 21573 8234
rect 21607 7458 21619 8234
rect 21561 7446 21619 7458
rect 21819 8234 21877 8246
rect 21819 7458 21831 8234
rect 21865 7458 21877 8234
rect 21819 7446 21877 7458
rect 21933 8234 21991 8246
rect 21933 7458 21945 8234
rect 21979 7458 21991 8234
rect 21933 7446 21991 7458
rect 22191 8234 22249 8246
rect 22191 7458 22203 8234
rect 22237 7458 22249 8234
rect 22191 7446 22249 7458
rect 22305 8234 22363 8246
rect 22305 7458 22317 8234
rect 22351 7458 22363 8234
rect 22305 7446 22363 7458
rect 22563 8234 22621 8246
rect 22563 7458 22575 8234
rect 22609 7458 22621 8234
rect 22563 7446 22621 7458
rect 22677 8234 22735 8246
rect 22677 7458 22689 8234
rect 22723 7458 22735 8234
rect 22677 7446 22735 7458
rect 22935 8234 22993 8246
rect 22935 7458 22947 8234
rect 22981 7458 22993 8234
rect 22935 7446 22993 7458
rect 23049 8234 23107 8246
rect 23049 7458 23061 8234
rect 23095 7458 23107 8234
rect 23049 7446 23107 7458
rect 23307 8234 23365 8246
rect 23307 7458 23319 8234
rect 23353 7458 23365 8234
rect 23307 7446 23365 7458
rect 23421 8234 23479 8246
rect 23421 7458 23433 8234
rect 23467 7458 23479 8234
rect 23421 7446 23479 7458
rect 23679 8234 23737 8246
rect 23679 7458 23691 8234
rect 23725 7458 23737 8234
rect 23679 7446 23737 7458
rect 20817 7198 20875 7210
rect 20817 6422 20829 7198
rect 20863 6422 20875 7198
rect 20817 6410 20875 6422
rect 21075 7198 21133 7210
rect 21075 6422 21087 7198
rect 21121 6422 21133 7198
rect 21075 6410 21133 6422
rect 21189 7198 21247 7210
rect 21189 6422 21201 7198
rect 21235 6422 21247 7198
rect 21189 6410 21247 6422
rect 21447 7198 21505 7210
rect 21447 6422 21459 7198
rect 21493 6422 21505 7198
rect 21447 6410 21505 6422
rect 21561 7198 21619 7210
rect 21561 6422 21573 7198
rect 21607 6422 21619 7198
rect 21561 6410 21619 6422
rect 21819 7198 21877 7210
rect 21819 6422 21831 7198
rect 21865 6422 21877 7198
rect 21819 6410 21877 6422
rect 21933 7198 21991 7210
rect 21933 6422 21945 7198
rect 21979 6422 21991 7198
rect 21933 6410 21991 6422
rect 22191 7198 22249 7210
rect 22191 6422 22203 7198
rect 22237 6422 22249 7198
rect 22191 6410 22249 6422
rect 22305 7198 22363 7210
rect 22305 6422 22317 7198
rect 22351 6422 22363 7198
rect 22305 6410 22363 6422
rect 22563 7198 22621 7210
rect 22563 6422 22575 7198
rect 22609 6422 22621 7198
rect 22563 6410 22621 6422
rect 22677 7198 22735 7210
rect 22677 6422 22689 7198
rect 22723 6422 22735 7198
rect 22677 6410 22735 6422
rect 22935 7198 22993 7210
rect 22935 6422 22947 7198
rect 22981 6422 22993 7198
rect 22935 6410 22993 6422
rect 23049 7198 23107 7210
rect 23049 6422 23061 7198
rect 23095 6422 23107 7198
rect 23049 6410 23107 6422
rect 23307 7198 23365 7210
rect 23307 6422 23319 7198
rect 23353 6422 23365 7198
rect 23307 6410 23365 6422
rect 23421 7198 23479 7210
rect 23421 6422 23433 7198
rect 23467 6422 23479 7198
rect 23421 6410 23479 6422
rect 23679 7198 23737 7210
rect 23679 6422 23691 7198
rect 23725 6422 23737 7198
rect 23679 6410 23737 6422
rect 20817 6162 20875 6174
rect 20817 5386 20829 6162
rect 20863 5386 20875 6162
rect 20817 5374 20875 5386
rect 21075 6162 21133 6174
rect 21075 5386 21087 6162
rect 21121 5386 21133 6162
rect 21075 5374 21133 5386
rect 21189 6162 21247 6174
rect 21189 5386 21201 6162
rect 21235 5386 21247 6162
rect 21189 5374 21247 5386
rect 21447 6162 21505 6174
rect 21447 5386 21459 6162
rect 21493 5386 21505 6162
rect 21447 5374 21505 5386
rect 21561 6162 21619 6174
rect 21561 5386 21573 6162
rect 21607 5386 21619 6162
rect 21561 5374 21619 5386
rect 21819 6162 21877 6174
rect 21819 5386 21831 6162
rect 21865 5386 21877 6162
rect 21819 5374 21877 5386
rect 21933 6162 21991 6174
rect 21933 5386 21945 6162
rect 21979 5386 21991 6162
rect 21933 5374 21991 5386
rect 22191 6162 22249 6174
rect 22191 5386 22203 6162
rect 22237 5386 22249 6162
rect 22191 5374 22249 5386
rect 22305 6162 22363 6174
rect 22305 5386 22317 6162
rect 22351 5386 22363 6162
rect 22305 5374 22363 5386
rect 22563 6162 22621 6174
rect 22563 5386 22575 6162
rect 22609 5386 22621 6162
rect 22563 5374 22621 5386
rect 22677 6162 22735 6174
rect 22677 5386 22689 6162
rect 22723 5386 22735 6162
rect 22677 5374 22735 5386
rect 22935 6162 22993 6174
rect 22935 5386 22947 6162
rect 22981 5386 22993 6162
rect 22935 5374 22993 5386
rect 23049 6162 23107 6174
rect 23049 5386 23061 6162
rect 23095 5386 23107 6162
rect 23049 5374 23107 5386
rect 23307 6162 23365 6174
rect 23307 5386 23319 6162
rect 23353 5386 23365 6162
rect 23307 5374 23365 5386
rect 23421 6162 23479 6174
rect 23421 5386 23433 6162
rect 23467 5386 23479 6162
rect 23421 5374 23479 5386
rect 23679 6162 23737 6174
rect 23679 5386 23691 6162
rect 23725 5386 23737 6162
rect 23679 5374 23737 5386
rect 20817 5126 20875 5138
rect 20817 4350 20829 5126
rect 20863 4350 20875 5126
rect 20817 4338 20875 4350
rect 21075 5126 21133 5138
rect 21075 4350 21087 5126
rect 21121 4350 21133 5126
rect 21075 4338 21133 4350
rect 21189 5126 21247 5138
rect 21189 4350 21201 5126
rect 21235 4350 21247 5126
rect 21189 4338 21247 4350
rect 21447 5126 21505 5138
rect 21447 4350 21459 5126
rect 21493 4350 21505 5126
rect 21447 4338 21505 4350
rect 21561 5126 21619 5138
rect 21561 4350 21573 5126
rect 21607 4350 21619 5126
rect 21561 4338 21619 4350
rect 21819 5126 21877 5138
rect 21819 4350 21831 5126
rect 21865 4350 21877 5126
rect 21819 4338 21877 4350
rect 21933 5126 21991 5138
rect 21933 4350 21945 5126
rect 21979 4350 21991 5126
rect 21933 4338 21991 4350
rect 22191 5126 22249 5138
rect 22191 4350 22203 5126
rect 22237 4350 22249 5126
rect 22191 4338 22249 4350
rect 22305 5126 22363 5138
rect 22305 4350 22317 5126
rect 22351 4350 22363 5126
rect 22305 4338 22363 4350
rect 22563 5126 22621 5138
rect 22563 4350 22575 5126
rect 22609 4350 22621 5126
rect 22563 4338 22621 4350
rect 22677 5126 22735 5138
rect 22677 4350 22689 5126
rect 22723 4350 22735 5126
rect 22677 4338 22735 4350
rect 22935 5126 22993 5138
rect 22935 4350 22947 5126
rect 22981 4350 22993 5126
rect 22935 4338 22993 4350
rect 23049 5126 23107 5138
rect 23049 4350 23061 5126
rect 23095 4350 23107 5126
rect 23049 4338 23107 4350
rect 23307 5126 23365 5138
rect 23307 4350 23319 5126
rect 23353 4350 23365 5126
rect 23307 4338 23365 4350
rect 23421 5126 23479 5138
rect 23421 4350 23433 5126
rect 23467 4350 23479 5126
rect 23421 4338 23479 4350
rect 23679 5126 23737 5138
rect 23679 4350 23691 5126
rect 23725 4350 23737 5126
rect 23679 4338 23737 4350
<< ndiffc >>
rect 20829 3373 20863 3549
rect 21087 3373 21121 3549
rect 21201 3373 21235 3549
rect 21459 3373 21493 3549
rect 21573 3373 21607 3549
rect 21831 3373 21865 3549
rect 21945 3373 21979 3549
rect 22203 3373 22237 3549
rect 22317 3373 22351 3549
rect 22575 3373 22609 3549
rect 22689 3373 22723 3549
rect 22947 3373 22981 3549
rect 23061 3373 23095 3549
rect 23319 3373 23353 3549
rect 23433 3373 23467 3549
rect 23691 3373 23725 3549
rect 23805 3373 23839 3549
rect 24063 3373 24097 3549
rect 24177 3373 24211 3549
rect 24435 3373 24469 3549
rect 24549 3373 24583 3549
rect 24807 3373 24841 3549
rect 24921 3373 24955 3549
rect 25179 3373 25213 3549
rect 25293 3373 25327 3549
rect 25551 3373 25585 3549
rect 25665 3373 25699 3549
rect 25923 3373 25957 3549
rect 26037 3373 26071 3549
rect 26295 3373 26329 3549
rect 26409 3373 26443 3549
rect 26667 3373 26701 3549
rect 26781 3373 26815 3549
rect 27039 3373 27073 3549
rect 27153 3373 27187 3549
rect 27411 3373 27445 3549
rect 27525 3373 27559 3549
rect 27783 3373 27817 3549
rect 27897 3373 27931 3549
rect 28155 3373 28189 3549
rect 28269 3373 28303 3549
rect 28527 3373 28561 3549
rect 28641 3373 28675 3549
rect 28899 3373 28933 3549
rect 29013 3373 29047 3549
rect 29271 3373 29305 3549
rect 29385 3373 29419 3549
rect 29643 3373 29677 3549
rect 20829 2955 20863 3131
rect 21087 2955 21121 3131
rect 21201 2955 21235 3131
rect 21459 2955 21493 3131
rect 21573 2955 21607 3131
rect 21831 2955 21865 3131
rect 21945 2955 21979 3131
rect 22203 2955 22237 3131
rect 22317 2955 22351 3131
rect 22575 2955 22609 3131
rect 22689 2955 22723 3131
rect 22947 2955 22981 3131
rect 23061 2955 23095 3131
rect 23319 2955 23353 3131
rect 23433 2955 23467 3131
rect 23691 2955 23725 3131
rect 23805 2955 23839 3131
rect 24063 2955 24097 3131
rect 24177 2955 24211 3131
rect 24435 2955 24469 3131
rect 24549 2955 24583 3131
rect 24807 2955 24841 3131
rect 24921 2955 24955 3131
rect 25179 2955 25213 3131
rect 25293 2955 25327 3131
rect 25551 2955 25585 3131
rect 25665 2955 25699 3131
rect 25923 2955 25957 3131
rect 26037 2955 26071 3131
rect 26295 2955 26329 3131
rect 26409 2955 26443 3131
rect 26667 2955 26701 3131
rect 26781 2955 26815 3131
rect 27039 2955 27073 3131
rect 27153 2955 27187 3131
rect 27411 2955 27445 3131
rect 27525 2955 27559 3131
rect 27783 2955 27817 3131
rect 27897 2955 27931 3131
rect 28155 2955 28189 3131
rect 28269 2955 28303 3131
rect 28527 2955 28561 3131
rect 28641 2955 28675 3131
rect 28899 2955 28933 3131
rect 29013 2955 29047 3131
rect 29271 2955 29305 3131
rect 29385 2955 29419 3131
rect 29643 2955 29677 3131
rect 20829 2537 20863 2713
rect 21087 2537 21121 2713
rect 21201 2537 21235 2713
rect 21459 2537 21493 2713
rect 21573 2537 21607 2713
rect 21831 2537 21865 2713
rect 21945 2537 21979 2713
rect 22203 2537 22237 2713
rect 22317 2537 22351 2713
rect 22575 2537 22609 2713
rect 22689 2537 22723 2713
rect 22947 2537 22981 2713
rect 23061 2537 23095 2713
rect 23319 2537 23353 2713
rect 23433 2537 23467 2713
rect 23691 2537 23725 2713
rect 23805 2537 23839 2713
rect 24063 2537 24097 2713
rect 24177 2537 24211 2713
rect 24435 2537 24469 2713
rect 24549 2537 24583 2713
rect 24807 2537 24841 2713
rect 24921 2537 24955 2713
rect 25179 2537 25213 2713
rect 25293 2537 25327 2713
rect 25551 2537 25585 2713
rect 25665 2537 25699 2713
rect 25923 2537 25957 2713
rect 26037 2537 26071 2713
rect 26295 2537 26329 2713
rect 26409 2537 26443 2713
rect 26667 2537 26701 2713
rect 26781 2537 26815 2713
rect 27039 2537 27073 2713
rect 27153 2537 27187 2713
rect 27411 2537 27445 2713
rect 27525 2537 27559 2713
rect 27783 2537 27817 2713
rect 27897 2537 27931 2713
rect 28155 2537 28189 2713
rect 28269 2537 28303 2713
rect 28527 2537 28561 2713
rect 28641 2537 28675 2713
rect 28899 2537 28933 2713
rect 29013 2537 29047 2713
rect 29271 2537 29305 2713
rect 29385 2537 29419 2713
rect 29643 2537 29677 2713
rect 20829 2119 20863 2295
rect 21087 2119 21121 2295
rect 21201 2119 21235 2295
rect 21459 2119 21493 2295
rect 21573 2119 21607 2295
rect 21831 2119 21865 2295
rect 21945 2119 21979 2295
rect 22203 2119 22237 2295
rect 22317 2119 22351 2295
rect 22575 2119 22609 2295
rect 22689 2119 22723 2295
rect 22947 2119 22981 2295
rect 23061 2119 23095 2295
rect 23319 2119 23353 2295
rect 23433 2119 23467 2295
rect 23691 2119 23725 2295
rect 23805 2119 23839 2295
rect 24063 2119 24097 2295
rect 24177 2119 24211 2295
rect 24435 2119 24469 2295
rect 24549 2119 24583 2295
rect 24807 2119 24841 2295
rect 24921 2119 24955 2295
rect 25179 2119 25213 2295
rect 25293 2119 25327 2295
rect 25551 2119 25585 2295
rect 25665 2119 25699 2295
rect 25923 2119 25957 2295
rect 26037 2119 26071 2295
rect 26295 2119 26329 2295
rect 26409 2119 26443 2295
rect 26667 2119 26701 2295
rect 26781 2119 26815 2295
rect 27039 2119 27073 2295
rect 27153 2119 27187 2295
rect 27411 2119 27445 2295
rect 27525 2119 27559 2295
rect 27783 2119 27817 2295
rect 27897 2119 27931 2295
rect 28155 2119 28189 2295
rect 28269 2119 28303 2295
rect 28527 2119 28561 2295
rect 28641 2119 28675 2295
rect 28899 2119 28933 2295
rect 29013 2119 29047 2295
rect 29271 2119 29305 2295
rect 29385 2119 29419 2295
rect 29643 2119 29677 2295
<< pdiffc >>
rect 19341 10246 19375 10622
rect 19599 10246 19633 10622
rect 19713 10246 19747 10622
rect 19971 10246 20005 10622
rect 20085 10246 20119 10622
rect 20343 10246 20377 10622
rect 20457 10246 20491 10622
rect 20715 10246 20749 10622
rect 20829 10246 20863 10622
rect 21087 10246 21121 10622
rect 21201 10246 21235 10622
rect 21459 10246 21493 10622
rect 21573 10246 21607 10622
rect 21831 10246 21865 10622
rect 21945 10246 21979 10622
rect 22203 10246 22237 10622
rect 22317 10246 22351 10622
rect 22575 10246 22609 10622
rect 22689 10246 22723 10622
rect 22947 10246 22981 10622
rect 23061 10246 23095 10622
rect 23319 10246 23353 10622
rect 23433 10246 23467 10622
rect 23691 10246 23725 10622
rect 23805 10246 23839 10622
rect 24063 10246 24097 10622
rect 24177 10246 24211 10622
rect 24435 10246 24469 10622
rect 24549 10246 24583 10622
rect 24807 10246 24841 10622
rect 24921 10246 24955 10622
rect 25179 10246 25213 10622
rect 25293 10246 25327 10622
rect 25551 10246 25585 10622
rect 25665 10246 25699 10622
rect 25923 10246 25957 10622
rect 26037 10246 26071 10622
rect 26295 10246 26329 10622
rect 26409 10246 26443 10622
rect 26667 10246 26701 10622
rect 26781 10246 26815 10622
rect 27039 10246 27073 10622
rect 27153 10246 27187 10622
rect 27411 10246 27445 10622
rect 27525 10246 27559 10622
rect 27783 10246 27817 10622
rect 27897 10246 27931 10622
rect 28155 10246 28189 10622
rect 28269 10246 28303 10622
rect 28527 10246 28561 10622
rect 28641 10246 28675 10622
rect 28899 10246 28933 10622
rect 29013 10246 29047 10622
rect 29271 10246 29305 10622
rect 29385 10246 29419 10622
rect 29643 10246 29677 10622
rect 29757 10246 29791 10622
rect 30015 10246 30049 10622
rect 30129 10246 30163 10622
rect 30387 10246 30421 10622
rect 30501 10246 30535 10622
rect 30759 10246 30793 10622
rect 30873 10246 30907 10622
rect 31131 10246 31165 10622
rect 19341 9610 19375 9986
rect 19599 9610 19633 9986
rect 19713 9610 19747 9986
rect 19971 9610 20005 9986
rect 20085 9610 20119 9986
rect 20343 9610 20377 9986
rect 20457 9610 20491 9986
rect 20715 9610 20749 9986
rect 20829 9610 20863 9986
rect 21087 9610 21121 9986
rect 21201 9610 21235 9986
rect 21459 9610 21493 9986
rect 21573 9610 21607 9986
rect 21831 9610 21865 9986
rect 21945 9610 21979 9986
rect 22203 9610 22237 9986
rect 22317 9610 22351 9986
rect 22575 9610 22609 9986
rect 22689 9610 22723 9986
rect 22947 9610 22981 9986
rect 23061 9610 23095 9986
rect 23319 9610 23353 9986
rect 23433 9610 23467 9986
rect 23691 9610 23725 9986
rect 23805 9610 23839 9986
rect 24063 9610 24097 9986
rect 24177 9610 24211 9986
rect 24435 9610 24469 9986
rect 24549 9610 24583 9986
rect 24807 9610 24841 9986
rect 24921 9610 24955 9986
rect 25179 9610 25213 9986
rect 25293 9610 25327 9986
rect 25551 9610 25585 9986
rect 25665 9610 25699 9986
rect 25923 9610 25957 9986
rect 26037 9610 26071 9986
rect 26295 9610 26329 9986
rect 26409 9610 26443 9986
rect 26667 9610 26701 9986
rect 26781 9610 26815 9986
rect 27039 9610 27073 9986
rect 27153 9610 27187 9986
rect 27411 9610 27445 9986
rect 27525 9610 27559 9986
rect 27783 9610 27817 9986
rect 27897 9610 27931 9986
rect 28155 9610 28189 9986
rect 28269 9610 28303 9986
rect 28527 9610 28561 9986
rect 28641 9610 28675 9986
rect 28899 9610 28933 9986
rect 29013 9610 29047 9986
rect 29271 9610 29305 9986
rect 29385 9610 29419 9986
rect 29643 9610 29677 9986
rect 29757 9610 29791 9986
rect 30015 9610 30049 9986
rect 30129 9610 30163 9986
rect 30387 9610 30421 9986
rect 30501 9610 30535 9986
rect 30759 9610 30793 9986
rect 30873 9610 30907 9986
rect 31131 9610 31165 9986
rect 19341 8974 19375 9350
rect 19599 8974 19633 9350
rect 19713 8974 19747 9350
rect 19971 8974 20005 9350
rect 20085 8974 20119 9350
rect 20343 8974 20377 9350
rect 20457 8974 20491 9350
rect 20715 8974 20749 9350
rect 20829 8974 20863 9350
rect 21087 8974 21121 9350
rect 21201 8974 21235 9350
rect 21459 8974 21493 9350
rect 21573 8974 21607 9350
rect 21831 8974 21865 9350
rect 21945 8974 21979 9350
rect 22203 8974 22237 9350
rect 22317 8974 22351 9350
rect 22575 8974 22609 9350
rect 22689 8974 22723 9350
rect 22947 8974 22981 9350
rect 23061 8974 23095 9350
rect 23319 8974 23353 9350
rect 23433 8974 23467 9350
rect 23691 8974 23725 9350
rect 23805 8974 23839 9350
rect 24063 8974 24097 9350
rect 24177 8974 24211 9350
rect 24435 8974 24469 9350
rect 24549 8974 24583 9350
rect 24807 8974 24841 9350
rect 24921 8974 24955 9350
rect 25179 8974 25213 9350
rect 25293 8974 25327 9350
rect 25551 8974 25585 9350
rect 25665 8974 25699 9350
rect 25923 8974 25957 9350
rect 26037 8974 26071 9350
rect 26295 8974 26329 9350
rect 26409 8974 26443 9350
rect 26667 8974 26701 9350
rect 26781 8974 26815 9350
rect 27039 8974 27073 9350
rect 27153 8974 27187 9350
rect 27411 8974 27445 9350
rect 27525 8974 27559 9350
rect 27783 8974 27817 9350
rect 27897 8974 27931 9350
rect 28155 8974 28189 9350
rect 28269 8974 28303 9350
rect 28527 8974 28561 9350
rect 28641 8974 28675 9350
rect 28899 8974 28933 9350
rect 29013 8974 29047 9350
rect 29271 8974 29305 9350
rect 29385 8974 29419 9350
rect 29643 8974 29677 9350
rect 29757 8974 29791 9350
rect 30015 8974 30049 9350
rect 30129 8974 30163 9350
rect 30387 8974 30421 9350
rect 30501 8974 30535 9350
rect 30759 8974 30793 9350
rect 30873 8974 30907 9350
rect 31131 8974 31165 9350
rect 20829 7458 20863 8234
rect 21087 7458 21121 8234
rect 21201 7458 21235 8234
rect 21459 7458 21493 8234
rect 21573 7458 21607 8234
rect 21831 7458 21865 8234
rect 21945 7458 21979 8234
rect 22203 7458 22237 8234
rect 22317 7458 22351 8234
rect 22575 7458 22609 8234
rect 22689 7458 22723 8234
rect 22947 7458 22981 8234
rect 23061 7458 23095 8234
rect 23319 7458 23353 8234
rect 23433 7458 23467 8234
rect 23691 7458 23725 8234
rect 20829 6422 20863 7198
rect 21087 6422 21121 7198
rect 21201 6422 21235 7198
rect 21459 6422 21493 7198
rect 21573 6422 21607 7198
rect 21831 6422 21865 7198
rect 21945 6422 21979 7198
rect 22203 6422 22237 7198
rect 22317 6422 22351 7198
rect 22575 6422 22609 7198
rect 22689 6422 22723 7198
rect 22947 6422 22981 7198
rect 23061 6422 23095 7198
rect 23319 6422 23353 7198
rect 23433 6422 23467 7198
rect 23691 6422 23725 7198
rect 20829 5386 20863 6162
rect 21087 5386 21121 6162
rect 21201 5386 21235 6162
rect 21459 5386 21493 6162
rect 21573 5386 21607 6162
rect 21831 5386 21865 6162
rect 21945 5386 21979 6162
rect 22203 5386 22237 6162
rect 22317 5386 22351 6162
rect 22575 5386 22609 6162
rect 22689 5386 22723 6162
rect 22947 5386 22981 6162
rect 23061 5386 23095 6162
rect 23319 5386 23353 6162
rect 23433 5386 23467 6162
rect 23691 5386 23725 6162
rect 20829 4350 20863 5126
rect 21087 4350 21121 5126
rect 21201 4350 21235 5126
rect 21459 4350 21493 5126
rect 21573 4350 21607 5126
rect 21831 4350 21865 5126
rect 21945 4350 21979 5126
rect 22203 4350 22237 5126
rect 22317 4350 22351 5126
rect 22575 4350 22609 5126
rect 22689 4350 22723 5126
rect 22947 4350 22981 5126
rect 23061 4350 23095 5126
rect 23319 4350 23353 5126
rect 23433 4350 23467 5126
rect 23691 4350 23725 5126
<< psubdiff >>
rect 20715 3701 20811 3735
rect 29695 3701 29791 3735
rect 20715 3639 20749 3701
rect 29757 3639 29791 3701
rect 20715 1967 20749 2029
rect 29757 1967 29791 2029
rect 20715 1933 20811 1967
rect 29695 1933 29791 1967
<< nsubdiff >>
rect 19227 10783 19323 10817
rect 31183 10783 31279 10817
rect 19227 10721 19261 10783
rect 31245 10721 31279 10783
rect 19227 8813 19261 8875
rect 31245 8813 31279 8875
rect 19227 8779 19323 8813
rect 31183 8779 31279 8813
rect 20715 8395 20811 8429
rect 23743 8395 23839 8429
rect 20715 8333 20749 8395
rect 23805 8333 23839 8395
rect 20715 4189 20749 4251
rect 23805 4189 23839 4251
rect 20715 4155 20811 4189
rect 23743 4155 23839 4189
<< psubdiffcont >>
rect 20811 3701 29695 3735
rect 20715 2029 20749 3639
rect 29757 2029 29791 3639
rect 20811 1933 29695 1967
<< nsubdiffcont >>
rect 19323 10783 31183 10817
rect 19227 8875 19261 10721
rect 31245 8875 31279 10721
rect 19323 8779 31183 8813
rect 20811 8395 23743 8429
rect 20715 4251 20749 8333
rect 23805 4251 23839 8333
rect 20811 4155 23743 4189
<< poly >>
rect 19387 10715 19587 10731
rect 19387 10681 19403 10715
rect 19571 10681 19587 10715
rect 19387 10634 19587 10681
rect 19759 10715 19959 10731
rect 19759 10681 19775 10715
rect 19943 10681 19959 10715
rect 19759 10634 19959 10681
rect 20131 10715 20331 10731
rect 20131 10681 20147 10715
rect 20315 10681 20331 10715
rect 20131 10634 20331 10681
rect 20503 10715 20703 10731
rect 20503 10681 20519 10715
rect 20687 10681 20703 10715
rect 20503 10634 20703 10681
rect 20875 10715 21075 10731
rect 20875 10681 20891 10715
rect 21059 10681 21075 10715
rect 20875 10634 21075 10681
rect 21247 10715 21447 10731
rect 21247 10681 21263 10715
rect 21431 10681 21447 10715
rect 21247 10634 21447 10681
rect 21619 10715 21819 10731
rect 21619 10681 21635 10715
rect 21803 10681 21819 10715
rect 21619 10634 21819 10681
rect 21991 10715 22191 10731
rect 21991 10681 22007 10715
rect 22175 10681 22191 10715
rect 21991 10634 22191 10681
rect 22363 10715 22563 10731
rect 22363 10681 22379 10715
rect 22547 10681 22563 10715
rect 22363 10634 22563 10681
rect 22735 10715 22935 10731
rect 22735 10681 22751 10715
rect 22919 10681 22935 10715
rect 22735 10634 22935 10681
rect 23107 10715 23307 10731
rect 23107 10681 23123 10715
rect 23291 10681 23307 10715
rect 23107 10634 23307 10681
rect 23479 10715 23679 10731
rect 23479 10681 23495 10715
rect 23663 10681 23679 10715
rect 23479 10634 23679 10681
rect 23851 10715 24051 10731
rect 23851 10681 23867 10715
rect 24035 10681 24051 10715
rect 23851 10634 24051 10681
rect 24223 10715 24423 10731
rect 24223 10681 24239 10715
rect 24407 10681 24423 10715
rect 24223 10634 24423 10681
rect 24595 10715 24795 10731
rect 24595 10681 24611 10715
rect 24779 10681 24795 10715
rect 24595 10634 24795 10681
rect 24967 10715 25167 10731
rect 24967 10681 24983 10715
rect 25151 10681 25167 10715
rect 24967 10634 25167 10681
rect 25339 10715 25539 10731
rect 25339 10681 25355 10715
rect 25523 10681 25539 10715
rect 25339 10634 25539 10681
rect 25711 10715 25911 10731
rect 25711 10681 25727 10715
rect 25895 10681 25911 10715
rect 25711 10634 25911 10681
rect 26083 10715 26283 10731
rect 26083 10681 26099 10715
rect 26267 10681 26283 10715
rect 26083 10634 26283 10681
rect 26455 10715 26655 10731
rect 26455 10681 26471 10715
rect 26639 10681 26655 10715
rect 26455 10634 26655 10681
rect 26827 10715 27027 10731
rect 26827 10681 26843 10715
rect 27011 10681 27027 10715
rect 26827 10634 27027 10681
rect 27199 10715 27399 10731
rect 27199 10681 27215 10715
rect 27383 10681 27399 10715
rect 27199 10634 27399 10681
rect 27571 10715 27771 10731
rect 27571 10681 27587 10715
rect 27755 10681 27771 10715
rect 27571 10634 27771 10681
rect 27943 10715 28143 10731
rect 27943 10681 27959 10715
rect 28127 10681 28143 10715
rect 27943 10634 28143 10681
rect 28315 10715 28515 10731
rect 28315 10681 28331 10715
rect 28499 10681 28515 10715
rect 28315 10634 28515 10681
rect 28687 10715 28887 10731
rect 28687 10681 28703 10715
rect 28871 10681 28887 10715
rect 28687 10634 28887 10681
rect 29059 10715 29259 10731
rect 29059 10681 29075 10715
rect 29243 10681 29259 10715
rect 29059 10634 29259 10681
rect 29431 10715 29631 10731
rect 29431 10681 29447 10715
rect 29615 10681 29631 10715
rect 29431 10634 29631 10681
rect 29803 10715 30003 10731
rect 29803 10681 29819 10715
rect 29987 10681 30003 10715
rect 29803 10634 30003 10681
rect 30175 10715 30375 10731
rect 30175 10681 30191 10715
rect 30359 10681 30375 10715
rect 30175 10634 30375 10681
rect 30547 10715 30747 10731
rect 30547 10681 30563 10715
rect 30731 10681 30747 10715
rect 30547 10634 30747 10681
rect 30919 10715 31119 10731
rect 30919 10681 30935 10715
rect 31103 10681 31119 10715
rect 30919 10634 31119 10681
rect 19387 10187 19587 10234
rect 19387 10153 19403 10187
rect 19571 10153 19587 10187
rect 19387 10137 19587 10153
rect 19759 10187 19959 10234
rect 19759 10153 19775 10187
rect 19943 10153 19959 10187
rect 19759 10137 19959 10153
rect 20131 10187 20331 10234
rect 20131 10153 20147 10187
rect 20315 10153 20331 10187
rect 20131 10137 20331 10153
rect 20503 10187 20703 10234
rect 20503 10153 20519 10187
rect 20687 10153 20703 10187
rect 20503 10137 20703 10153
rect 20875 10187 21075 10234
rect 20875 10153 20891 10187
rect 21059 10153 21075 10187
rect 20875 10137 21075 10153
rect 21247 10187 21447 10234
rect 21247 10153 21263 10187
rect 21431 10153 21447 10187
rect 21247 10137 21447 10153
rect 21619 10187 21819 10234
rect 21619 10153 21635 10187
rect 21803 10153 21819 10187
rect 21619 10137 21819 10153
rect 21991 10187 22191 10234
rect 21991 10153 22007 10187
rect 22175 10153 22191 10187
rect 21991 10137 22191 10153
rect 22363 10187 22563 10234
rect 22363 10153 22379 10187
rect 22547 10153 22563 10187
rect 22363 10137 22563 10153
rect 22735 10187 22935 10234
rect 22735 10153 22751 10187
rect 22919 10153 22935 10187
rect 22735 10137 22935 10153
rect 23107 10187 23307 10234
rect 23107 10153 23123 10187
rect 23291 10153 23307 10187
rect 23107 10137 23307 10153
rect 23479 10187 23679 10234
rect 23479 10153 23495 10187
rect 23663 10153 23679 10187
rect 23479 10137 23679 10153
rect 23851 10187 24051 10234
rect 23851 10153 23867 10187
rect 24035 10153 24051 10187
rect 23851 10137 24051 10153
rect 24223 10187 24423 10234
rect 24223 10153 24239 10187
rect 24407 10153 24423 10187
rect 24223 10137 24423 10153
rect 24595 10187 24795 10234
rect 24595 10153 24611 10187
rect 24779 10153 24795 10187
rect 24595 10137 24795 10153
rect 24967 10187 25167 10234
rect 24967 10153 24983 10187
rect 25151 10153 25167 10187
rect 24967 10137 25167 10153
rect 25339 10187 25539 10234
rect 25339 10153 25355 10187
rect 25523 10153 25539 10187
rect 25339 10137 25539 10153
rect 25711 10187 25911 10234
rect 25711 10153 25727 10187
rect 25895 10153 25911 10187
rect 25711 10137 25911 10153
rect 26083 10187 26283 10234
rect 26083 10153 26099 10187
rect 26267 10153 26283 10187
rect 26083 10137 26283 10153
rect 26455 10187 26655 10234
rect 26455 10153 26471 10187
rect 26639 10153 26655 10187
rect 26455 10137 26655 10153
rect 26827 10187 27027 10234
rect 26827 10153 26843 10187
rect 27011 10153 27027 10187
rect 26827 10137 27027 10153
rect 27199 10187 27399 10234
rect 27199 10153 27215 10187
rect 27383 10153 27399 10187
rect 27199 10137 27399 10153
rect 27571 10187 27771 10234
rect 27571 10153 27587 10187
rect 27755 10153 27771 10187
rect 27571 10137 27771 10153
rect 27943 10187 28143 10234
rect 27943 10153 27959 10187
rect 28127 10153 28143 10187
rect 27943 10137 28143 10153
rect 28315 10187 28515 10234
rect 28315 10153 28331 10187
rect 28499 10153 28515 10187
rect 28315 10137 28515 10153
rect 28687 10187 28887 10234
rect 28687 10153 28703 10187
rect 28871 10153 28887 10187
rect 28687 10137 28887 10153
rect 29059 10187 29259 10234
rect 29059 10153 29075 10187
rect 29243 10153 29259 10187
rect 29059 10137 29259 10153
rect 29431 10187 29631 10234
rect 29431 10153 29447 10187
rect 29615 10153 29631 10187
rect 29431 10137 29631 10153
rect 29803 10187 30003 10234
rect 29803 10153 29819 10187
rect 29987 10153 30003 10187
rect 29803 10137 30003 10153
rect 30175 10187 30375 10234
rect 30175 10153 30191 10187
rect 30359 10153 30375 10187
rect 30175 10137 30375 10153
rect 30547 10187 30747 10234
rect 30547 10153 30563 10187
rect 30731 10153 30747 10187
rect 30547 10137 30747 10153
rect 30919 10187 31119 10234
rect 30919 10153 30935 10187
rect 31103 10153 31119 10187
rect 30919 10137 31119 10153
rect 19387 10079 19587 10095
rect 19387 10045 19403 10079
rect 19571 10045 19587 10079
rect 19387 9998 19587 10045
rect 19759 10079 19959 10095
rect 19759 10045 19775 10079
rect 19943 10045 19959 10079
rect 19759 9998 19959 10045
rect 20131 10079 20331 10095
rect 20131 10045 20147 10079
rect 20315 10045 20331 10079
rect 20131 9998 20331 10045
rect 20503 10079 20703 10095
rect 20503 10045 20519 10079
rect 20687 10045 20703 10079
rect 20503 9998 20703 10045
rect 20875 10079 21075 10095
rect 20875 10045 20891 10079
rect 21059 10045 21075 10079
rect 20875 9998 21075 10045
rect 21247 10079 21447 10095
rect 21247 10045 21263 10079
rect 21431 10045 21447 10079
rect 21247 9998 21447 10045
rect 21619 10079 21819 10095
rect 21619 10045 21635 10079
rect 21803 10045 21819 10079
rect 21619 9998 21819 10045
rect 21991 10079 22191 10095
rect 21991 10045 22007 10079
rect 22175 10045 22191 10079
rect 21991 9998 22191 10045
rect 22363 10079 22563 10095
rect 22363 10045 22379 10079
rect 22547 10045 22563 10079
rect 22363 9998 22563 10045
rect 22735 10079 22935 10095
rect 22735 10045 22751 10079
rect 22919 10045 22935 10079
rect 22735 9998 22935 10045
rect 23107 10079 23307 10095
rect 23107 10045 23123 10079
rect 23291 10045 23307 10079
rect 23107 9998 23307 10045
rect 23479 10079 23679 10095
rect 23479 10045 23495 10079
rect 23663 10045 23679 10079
rect 23479 9998 23679 10045
rect 23851 10079 24051 10095
rect 23851 10045 23867 10079
rect 24035 10045 24051 10079
rect 23851 9998 24051 10045
rect 24223 10079 24423 10095
rect 24223 10045 24239 10079
rect 24407 10045 24423 10079
rect 24223 9998 24423 10045
rect 24595 10079 24795 10095
rect 24595 10045 24611 10079
rect 24779 10045 24795 10079
rect 24595 9998 24795 10045
rect 24967 10079 25167 10095
rect 24967 10045 24983 10079
rect 25151 10045 25167 10079
rect 24967 9998 25167 10045
rect 25339 10079 25539 10095
rect 25339 10045 25355 10079
rect 25523 10045 25539 10079
rect 25339 9998 25539 10045
rect 25711 10079 25911 10095
rect 25711 10045 25727 10079
rect 25895 10045 25911 10079
rect 25711 9998 25911 10045
rect 26083 10079 26283 10095
rect 26083 10045 26099 10079
rect 26267 10045 26283 10079
rect 26083 9998 26283 10045
rect 26455 10079 26655 10095
rect 26455 10045 26471 10079
rect 26639 10045 26655 10079
rect 26455 9998 26655 10045
rect 26827 10079 27027 10095
rect 26827 10045 26843 10079
rect 27011 10045 27027 10079
rect 26827 9998 27027 10045
rect 27199 10079 27399 10095
rect 27199 10045 27215 10079
rect 27383 10045 27399 10079
rect 27199 9998 27399 10045
rect 27571 10079 27771 10095
rect 27571 10045 27587 10079
rect 27755 10045 27771 10079
rect 27571 9998 27771 10045
rect 27943 10079 28143 10095
rect 27943 10045 27959 10079
rect 28127 10045 28143 10079
rect 27943 9998 28143 10045
rect 28315 10079 28515 10095
rect 28315 10045 28331 10079
rect 28499 10045 28515 10079
rect 28315 9998 28515 10045
rect 28687 10079 28887 10095
rect 28687 10045 28703 10079
rect 28871 10045 28887 10079
rect 28687 9998 28887 10045
rect 29059 10079 29259 10095
rect 29059 10045 29075 10079
rect 29243 10045 29259 10079
rect 29059 9998 29259 10045
rect 29431 10079 29631 10095
rect 29431 10045 29447 10079
rect 29615 10045 29631 10079
rect 29431 9998 29631 10045
rect 29803 10079 30003 10095
rect 29803 10045 29819 10079
rect 29987 10045 30003 10079
rect 29803 9998 30003 10045
rect 30175 10079 30375 10095
rect 30175 10045 30191 10079
rect 30359 10045 30375 10079
rect 30175 9998 30375 10045
rect 30547 10079 30747 10095
rect 30547 10045 30563 10079
rect 30731 10045 30747 10079
rect 30547 9998 30747 10045
rect 30919 10079 31119 10095
rect 30919 10045 30935 10079
rect 31103 10045 31119 10079
rect 30919 9998 31119 10045
rect 19387 9551 19587 9598
rect 19387 9517 19403 9551
rect 19571 9517 19587 9551
rect 19387 9501 19587 9517
rect 19759 9551 19959 9598
rect 19759 9517 19775 9551
rect 19943 9517 19959 9551
rect 19759 9501 19959 9517
rect 20131 9551 20331 9598
rect 20131 9517 20147 9551
rect 20315 9517 20331 9551
rect 20131 9501 20331 9517
rect 20503 9551 20703 9598
rect 20503 9517 20519 9551
rect 20687 9517 20703 9551
rect 20503 9501 20703 9517
rect 20875 9551 21075 9598
rect 20875 9517 20891 9551
rect 21059 9517 21075 9551
rect 20875 9501 21075 9517
rect 21247 9551 21447 9598
rect 21247 9517 21263 9551
rect 21431 9517 21447 9551
rect 21247 9501 21447 9517
rect 21619 9551 21819 9598
rect 21619 9517 21635 9551
rect 21803 9517 21819 9551
rect 21619 9501 21819 9517
rect 21991 9551 22191 9598
rect 21991 9517 22007 9551
rect 22175 9517 22191 9551
rect 21991 9501 22191 9517
rect 22363 9551 22563 9598
rect 22363 9517 22379 9551
rect 22547 9517 22563 9551
rect 22363 9501 22563 9517
rect 22735 9551 22935 9598
rect 22735 9517 22751 9551
rect 22919 9517 22935 9551
rect 22735 9501 22935 9517
rect 23107 9551 23307 9598
rect 23107 9517 23123 9551
rect 23291 9517 23307 9551
rect 23107 9501 23307 9517
rect 23479 9551 23679 9598
rect 23479 9517 23495 9551
rect 23663 9517 23679 9551
rect 23479 9501 23679 9517
rect 23851 9551 24051 9598
rect 23851 9517 23867 9551
rect 24035 9517 24051 9551
rect 23851 9501 24051 9517
rect 24223 9551 24423 9598
rect 24223 9517 24239 9551
rect 24407 9517 24423 9551
rect 24223 9501 24423 9517
rect 24595 9551 24795 9598
rect 24595 9517 24611 9551
rect 24779 9517 24795 9551
rect 24595 9501 24795 9517
rect 24967 9551 25167 9598
rect 24967 9517 24983 9551
rect 25151 9517 25167 9551
rect 24967 9501 25167 9517
rect 25339 9551 25539 9598
rect 25339 9517 25355 9551
rect 25523 9517 25539 9551
rect 25339 9501 25539 9517
rect 25711 9551 25911 9598
rect 25711 9517 25727 9551
rect 25895 9517 25911 9551
rect 25711 9501 25911 9517
rect 26083 9551 26283 9598
rect 26083 9517 26099 9551
rect 26267 9517 26283 9551
rect 26083 9501 26283 9517
rect 26455 9551 26655 9598
rect 26455 9517 26471 9551
rect 26639 9517 26655 9551
rect 26455 9501 26655 9517
rect 26827 9551 27027 9598
rect 26827 9517 26843 9551
rect 27011 9517 27027 9551
rect 26827 9501 27027 9517
rect 27199 9551 27399 9598
rect 27199 9517 27215 9551
rect 27383 9517 27399 9551
rect 27199 9501 27399 9517
rect 27571 9551 27771 9598
rect 27571 9517 27587 9551
rect 27755 9517 27771 9551
rect 27571 9501 27771 9517
rect 27943 9551 28143 9598
rect 27943 9517 27959 9551
rect 28127 9517 28143 9551
rect 27943 9501 28143 9517
rect 28315 9551 28515 9598
rect 28315 9517 28331 9551
rect 28499 9517 28515 9551
rect 28315 9501 28515 9517
rect 28687 9551 28887 9598
rect 28687 9517 28703 9551
rect 28871 9517 28887 9551
rect 28687 9501 28887 9517
rect 29059 9551 29259 9598
rect 29059 9517 29075 9551
rect 29243 9517 29259 9551
rect 29059 9501 29259 9517
rect 29431 9551 29631 9598
rect 29431 9517 29447 9551
rect 29615 9517 29631 9551
rect 29431 9501 29631 9517
rect 29803 9551 30003 9598
rect 29803 9517 29819 9551
rect 29987 9517 30003 9551
rect 29803 9501 30003 9517
rect 30175 9551 30375 9598
rect 30175 9517 30191 9551
rect 30359 9517 30375 9551
rect 30175 9501 30375 9517
rect 30547 9551 30747 9598
rect 30547 9517 30563 9551
rect 30731 9517 30747 9551
rect 30547 9501 30747 9517
rect 30919 9551 31119 9598
rect 30919 9517 30935 9551
rect 31103 9517 31119 9551
rect 30919 9501 31119 9517
rect 19387 9443 19587 9459
rect 19387 9409 19403 9443
rect 19571 9409 19587 9443
rect 19387 9362 19587 9409
rect 19759 9443 19959 9459
rect 19759 9409 19775 9443
rect 19943 9409 19959 9443
rect 19759 9362 19959 9409
rect 20131 9443 20331 9459
rect 20131 9409 20147 9443
rect 20315 9409 20331 9443
rect 20131 9362 20331 9409
rect 20503 9443 20703 9459
rect 20503 9409 20519 9443
rect 20687 9409 20703 9443
rect 20503 9362 20703 9409
rect 20875 9443 21075 9459
rect 20875 9409 20891 9443
rect 21059 9409 21075 9443
rect 20875 9362 21075 9409
rect 21247 9443 21447 9459
rect 21247 9409 21263 9443
rect 21431 9409 21447 9443
rect 21247 9362 21447 9409
rect 21619 9443 21819 9459
rect 21619 9409 21635 9443
rect 21803 9409 21819 9443
rect 21619 9362 21819 9409
rect 21991 9443 22191 9459
rect 21991 9409 22007 9443
rect 22175 9409 22191 9443
rect 21991 9362 22191 9409
rect 22363 9443 22563 9459
rect 22363 9409 22379 9443
rect 22547 9409 22563 9443
rect 22363 9362 22563 9409
rect 22735 9443 22935 9459
rect 22735 9409 22751 9443
rect 22919 9409 22935 9443
rect 22735 9362 22935 9409
rect 23107 9443 23307 9459
rect 23107 9409 23123 9443
rect 23291 9409 23307 9443
rect 23107 9362 23307 9409
rect 23479 9443 23679 9459
rect 23479 9409 23495 9443
rect 23663 9409 23679 9443
rect 23479 9362 23679 9409
rect 23851 9443 24051 9459
rect 23851 9409 23867 9443
rect 24035 9409 24051 9443
rect 23851 9362 24051 9409
rect 24223 9443 24423 9459
rect 24223 9409 24239 9443
rect 24407 9409 24423 9443
rect 24223 9362 24423 9409
rect 24595 9443 24795 9459
rect 24595 9409 24611 9443
rect 24779 9409 24795 9443
rect 24595 9362 24795 9409
rect 24967 9443 25167 9459
rect 24967 9409 24983 9443
rect 25151 9409 25167 9443
rect 24967 9362 25167 9409
rect 25339 9443 25539 9459
rect 25339 9409 25355 9443
rect 25523 9409 25539 9443
rect 25339 9362 25539 9409
rect 25711 9443 25911 9459
rect 25711 9409 25727 9443
rect 25895 9409 25911 9443
rect 25711 9362 25911 9409
rect 26083 9443 26283 9459
rect 26083 9409 26099 9443
rect 26267 9409 26283 9443
rect 26083 9362 26283 9409
rect 26455 9443 26655 9459
rect 26455 9409 26471 9443
rect 26639 9409 26655 9443
rect 26455 9362 26655 9409
rect 26827 9443 27027 9459
rect 26827 9409 26843 9443
rect 27011 9409 27027 9443
rect 26827 9362 27027 9409
rect 27199 9443 27399 9459
rect 27199 9409 27215 9443
rect 27383 9409 27399 9443
rect 27199 9362 27399 9409
rect 27571 9443 27771 9459
rect 27571 9409 27587 9443
rect 27755 9409 27771 9443
rect 27571 9362 27771 9409
rect 27943 9443 28143 9459
rect 27943 9409 27959 9443
rect 28127 9409 28143 9443
rect 27943 9362 28143 9409
rect 28315 9443 28515 9459
rect 28315 9409 28331 9443
rect 28499 9409 28515 9443
rect 28315 9362 28515 9409
rect 28687 9443 28887 9459
rect 28687 9409 28703 9443
rect 28871 9409 28887 9443
rect 28687 9362 28887 9409
rect 29059 9443 29259 9459
rect 29059 9409 29075 9443
rect 29243 9409 29259 9443
rect 29059 9362 29259 9409
rect 29431 9443 29631 9459
rect 29431 9409 29447 9443
rect 29615 9409 29631 9443
rect 29431 9362 29631 9409
rect 29803 9443 30003 9459
rect 29803 9409 29819 9443
rect 29987 9409 30003 9443
rect 29803 9362 30003 9409
rect 30175 9443 30375 9459
rect 30175 9409 30191 9443
rect 30359 9409 30375 9443
rect 30175 9362 30375 9409
rect 30547 9443 30747 9459
rect 30547 9409 30563 9443
rect 30731 9409 30747 9443
rect 30547 9362 30747 9409
rect 30919 9443 31119 9459
rect 30919 9409 30935 9443
rect 31103 9409 31119 9443
rect 30919 9362 31119 9409
rect 19387 8915 19587 8962
rect 19387 8881 19403 8915
rect 19571 8881 19587 8915
rect 19387 8865 19587 8881
rect 19759 8915 19959 8962
rect 19759 8881 19775 8915
rect 19943 8881 19959 8915
rect 19759 8865 19959 8881
rect 20131 8915 20331 8962
rect 20131 8881 20147 8915
rect 20315 8881 20331 8915
rect 20131 8865 20331 8881
rect 20503 8915 20703 8962
rect 20503 8881 20519 8915
rect 20687 8881 20703 8915
rect 20503 8865 20703 8881
rect 20875 8915 21075 8962
rect 20875 8881 20891 8915
rect 21059 8881 21075 8915
rect 20875 8865 21075 8881
rect 21247 8915 21447 8962
rect 21247 8881 21263 8915
rect 21431 8881 21447 8915
rect 21247 8865 21447 8881
rect 21619 8915 21819 8962
rect 21619 8881 21635 8915
rect 21803 8881 21819 8915
rect 21619 8865 21819 8881
rect 21991 8915 22191 8962
rect 21991 8881 22007 8915
rect 22175 8881 22191 8915
rect 21991 8865 22191 8881
rect 22363 8915 22563 8962
rect 22363 8881 22379 8915
rect 22547 8881 22563 8915
rect 22363 8865 22563 8881
rect 22735 8915 22935 8962
rect 22735 8881 22751 8915
rect 22919 8881 22935 8915
rect 22735 8865 22935 8881
rect 23107 8915 23307 8962
rect 23107 8881 23123 8915
rect 23291 8881 23307 8915
rect 23107 8865 23307 8881
rect 23479 8915 23679 8962
rect 23479 8881 23495 8915
rect 23663 8881 23679 8915
rect 23479 8865 23679 8881
rect 23851 8915 24051 8962
rect 23851 8881 23867 8915
rect 24035 8881 24051 8915
rect 23851 8865 24051 8881
rect 24223 8915 24423 8962
rect 24223 8881 24239 8915
rect 24407 8881 24423 8915
rect 24223 8865 24423 8881
rect 24595 8915 24795 8962
rect 24595 8881 24611 8915
rect 24779 8881 24795 8915
rect 24595 8865 24795 8881
rect 24967 8915 25167 8962
rect 24967 8881 24983 8915
rect 25151 8881 25167 8915
rect 24967 8865 25167 8881
rect 25339 8915 25539 8962
rect 25339 8881 25355 8915
rect 25523 8881 25539 8915
rect 25339 8865 25539 8881
rect 25711 8915 25911 8962
rect 25711 8881 25727 8915
rect 25895 8881 25911 8915
rect 25711 8865 25911 8881
rect 26083 8915 26283 8962
rect 26083 8881 26099 8915
rect 26267 8881 26283 8915
rect 26083 8865 26283 8881
rect 26455 8915 26655 8962
rect 26455 8881 26471 8915
rect 26639 8881 26655 8915
rect 26455 8865 26655 8881
rect 26827 8915 27027 8962
rect 26827 8881 26843 8915
rect 27011 8881 27027 8915
rect 26827 8865 27027 8881
rect 27199 8915 27399 8962
rect 27199 8881 27215 8915
rect 27383 8881 27399 8915
rect 27199 8865 27399 8881
rect 27571 8915 27771 8962
rect 27571 8881 27587 8915
rect 27755 8881 27771 8915
rect 27571 8865 27771 8881
rect 27943 8915 28143 8962
rect 27943 8881 27959 8915
rect 28127 8881 28143 8915
rect 27943 8865 28143 8881
rect 28315 8915 28515 8962
rect 28315 8881 28331 8915
rect 28499 8881 28515 8915
rect 28315 8865 28515 8881
rect 28687 8915 28887 8962
rect 28687 8881 28703 8915
rect 28871 8881 28887 8915
rect 28687 8865 28887 8881
rect 29059 8915 29259 8962
rect 29059 8881 29075 8915
rect 29243 8881 29259 8915
rect 29059 8865 29259 8881
rect 29431 8915 29631 8962
rect 29431 8881 29447 8915
rect 29615 8881 29631 8915
rect 29431 8865 29631 8881
rect 29803 8915 30003 8962
rect 29803 8881 29819 8915
rect 29987 8881 30003 8915
rect 29803 8865 30003 8881
rect 30175 8915 30375 8962
rect 30175 8881 30191 8915
rect 30359 8881 30375 8915
rect 30175 8865 30375 8881
rect 30547 8915 30747 8962
rect 30547 8881 30563 8915
rect 30731 8881 30747 8915
rect 30547 8865 30747 8881
rect 30919 8915 31119 8962
rect 30919 8881 30935 8915
rect 31103 8881 31119 8915
rect 30919 8865 31119 8881
rect 20875 8327 21075 8343
rect 20875 8293 20891 8327
rect 21059 8293 21075 8327
rect 20875 8246 21075 8293
rect 21247 8327 21447 8343
rect 21247 8293 21263 8327
rect 21431 8293 21447 8327
rect 21247 8246 21447 8293
rect 21619 8327 21819 8343
rect 21619 8293 21635 8327
rect 21803 8293 21819 8327
rect 21619 8246 21819 8293
rect 21991 8327 22191 8343
rect 21991 8293 22007 8327
rect 22175 8293 22191 8327
rect 21991 8246 22191 8293
rect 22363 8327 22563 8343
rect 22363 8293 22379 8327
rect 22547 8293 22563 8327
rect 22363 8246 22563 8293
rect 22735 8327 22935 8343
rect 22735 8293 22751 8327
rect 22919 8293 22935 8327
rect 22735 8246 22935 8293
rect 23107 8327 23307 8343
rect 23107 8293 23123 8327
rect 23291 8293 23307 8327
rect 23107 8246 23307 8293
rect 23479 8327 23679 8343
rect 23479 8293 23495 8327
rect 23663 8293 23679 8327
rect 23479 8246 23679 8293
rect 20875 7399 21075 7446
rect 20875 7365 20891 7399
rect 21059 7365 21075 7399
rect 20875 7349 21075 7365
rect 21247 7399 21447 7446
rect 21247 7365 21263 7399
rect 21431 7365 21447 7399
rect 21247 7349 21447 7365
rect 21619 7399 21819 7446
rect 21619 7365 21635 7399
rect 21803 7365 21819 7399
rect 21619 7349 21819 7365
rect 21991 7399 22191 7446
rect 21991 7365 22007 7399
rect 22175 7365 22191 7399
rect 21991 7349 22191 7365
rect 22363 7399 22563 7446
rect 22363 7365 22379 7399
rect 22547 7365 22563 7399
rect 22363 7349 22563 7365
rect 22735 7399 22935 7446
rect 22735 7365 22751 7399
rect 22919 7365 22935 7399
rect 22735 7349 22935 7365
rect 23107 7399 23307 7446
rect 23107 7365 23123 7399
rect 23291 7365 23307 7399
rect 23107 7349 23307 7365
rect 23479 7399 23679 7446
rect 23479 7365 23495 7399
rect 23663 7365 23679 7399
rect 23479 7349 23679 7365
rect 20875 7291 21075 7307
rect 20875 7257 20891 7291
rect 21059 7257 21075 7291
rect 20875 7210 21075 7257
rect 21247 7291 21447 7307
rect 21247 7257 21263 7291
rect 21431 7257 21447 7291
rect 21247 7210 21447 7257
rect 21619 7291 21819 7307
rect 21619 7257 21635 7291
rect 21803 7257 21819 7291
rect 21619 7210 21819 7257
rect 21991 7291 22191 7307
rect 21991 7257 22007 7291
rect 22175 7257 22191 7291
rect 21991 7210 22191 7257
rect 22363 7291 22563 7307
rect 22363 7257 22379 7291
rect 22547 7257 22563 7291
rect 22363 7210 22563 7257
rect 22735 7291 22935 7307
rect 22735 7257 22751 7291
rect 22919 7257 22935 7291
rect 22735 7210 22935 7257
rect 23107 7291 23307 7307
rect 23107 7257 23123 7291
rect 23291 7257 23307 7291
rect 23107 7210 23307 7257
rect 23479 7291 23679 7307
rect 23479 7257 23495 7291
rect 23663 7257 23679 7291
rect 23479 7210 23679 7257
rect 20875 6363 21075 6410
rect 20875 6329 20891 6363
rect 21059 6329 21075 6363
rect 20875 6313 21075 6329
rect 21247 6363 21447 6410
rect 21247 6329 21263 6363
rect 21431 6329 21447 6363
rect 21247 6313 21447 6329
rect 21619 6363 21819 6410
rect 21619 6329 21635 6363
rect 21803 6329 21819 6363
rect 21619 6313 21819 6329
rect 21991 6363 22191 6410
rect 21991 6329 22007 6363
rect 22175 6329 22191 6363
rect 21991 6313 22191 6329
rect 22363 6363 22563 6410
rect 22363 6329 22379 6363
rect 22547 6329 22563 6363
rect 22363 6313 22563 6329
rect 22735 6363 22935 6410
rect 22735 6329 22751 6363
rect 22919 6329 22935 6363
rect 22735 6313 22935 6329
rect 23107 6363 23307 6410
rect 23107 6329 23123 6363
rect 23291 6329 23307 6363
rect 23107 6313 23307 6329
rect 23479 6363 23679 6410
rect 23479 6329 23495 6363
rect 23663 6329 23679 6363
rect 23479 6313 23679 6329
rect 20875 6255 21075 6271
rect 20875 6221 20891 6255
rect 21059 6221 21075 6255
rect 20875 6174 21075 6221
rect 21247 6255 21447 6271
rect 21247 6221 21263 6255
rect 21431 6221 21447 6255
rect 21247 6174 21447 6221
rect 21619 6255 21819 6271
rect 21619 6221 21635 6255
rect 21803 6221 21819 6255
rect 21619 6174 21819 6221
rect 21991 6255 22191 6271
rect 21991 6221 22007 6255
rect 22175 6221 22191 6255
rect 21991 6174 22191 6221
rect 22363 6255 22563 6271
rect 22363 6221 22379 6255
rect 22547 6221 22563 6255
rect 22363 6174 22563 6221
rect 22735 6255 22935 6271
rect 22735 6221 22751 6255
rect 22919 6221 22935 6255
rect 22735 6174 22935 6221
rect 23107 6255 23307 6271
rect 23107 6221 23123 6255
rect 23291 6221 23307 6255
rect 23107 6174 23307 6221
rect 23479 6255 23679 6271
rect 23479 6221 23495 6255
rect 23663 6221 23679 6255
rect 23479 6174 23679 6221
rect 20875 5327 21075 5374
rect 20875 5293 20891 5327
rect 21059 5293 21075 5327
rect 20875 5277 21075 5293
rect 21247 5327 21447 5374
rect 21247 5293 21263 5327
rect 21431 5293 21447 5327
rect 21247 5277 21447 5293
rect 21619 5327 21819 5374
rect 21619 5293 21635 5327
rect 21803 5293 21819 5327
rect 21619 5277 21819 5293
rect 21991 5327 22191 5374
rect 21991 5293 22007 5327
rect 22175 5293 22191 5327
rect 21991 5277 22191 5293
rect 22363 5327 22563 5374
rect 22363 5293 22379 5327
rect 22547 5293 22563 5327
rect 22363 5277 22563 5293
rect 22735 5327 22935 5374
rect 22735 5293 22751 5327
rect 22919 5293 22935 5327
rect 22735 5277 22935 5293
rect 23107 5327 23307 5374
rect 23107 5293 23123 5327
rect 23291 5293 23307 5327
rect 23107 5277 23307 5293
rect 23479 5327 23679 5374
rect 23479 5293 23495 5327
rect 23663 5293 23679 5327
rect 23479 5277 23679 5293
rect 20875 5219 21075 5235
rect 20875 5185 20891 5219
rect 21059 5185 21075 5219
rect 20875 5138 21075 5185
rect 21247 5219 21447 5235
rect 21247 5185 21263 5219
rect 21431 5185 21447 5219
rect 21247 5138 21447 5185
rect 21619 5219 21819 5235
rect 21619 5185 21635 5219
rect 21803 5185 21819 5219
rect 21619 5138 21819 5185
rect 21991 5219 22191 5235
rect 21991 5185 22007 5219
rect 22175 5185 22191 5219
rect 21991 5138 22191 5185
rect 22363 5219 22563 5235
rect 22363 5185 22379 5219
rect 22547 5185 22563 5219
rect 22363 5138 22563 5185
rect 22735 5219 22935 5235
rect 22735 5185 22751 5219
rect 22919 5185 22935 5219
rect 22735 5138 22935 5185
rect 23107 5219 23307 5235
rect 23107 5185 23123 5219
rect 23291 5185 23307 5219
rect 23107 5138 23307 5185
rect 23479 5219 23679 5235
rect 23479 5185 23495 5219
rect 23663 5185 23679 5219
rect 23479 5138 23679 5185
rect 20875 4291 21075 4338
rect 20875 4257 20891 4291
rect 21059 4257 21075 4291
rect 20875 4241 21075 4257
rect 21247 4291 21447 4338
rect 21247 4257 21263 4291
rect 21431 4257 21447 4291
rect 21247 4241 21447 4257
rect 21619 4291 21819 4338
rect 21619 4257 21635 4291
rect 21803 4257 21819 4291
rect 21619 4241 21819 4257
rect 21991 4291 22191 4338
rect 21991 4257 22007 4291
rect 22175 4257 22191 4291
rect 21991 4241 22191 4257
rect 22363 4291 22563 4338
rect 22363 4257 22379 4291
rect 22547 4257 22563 4291
rect 22363 4241 22563 4257
rect 22735 4291 22935 4338
rect 22735 4257 22751 4291
rect 22919 4257 22935 4291
rect 22735 4241 22935 4257
rect 23107 4291 23307 4338
rect 23107 4257 23123 4291
rect 23291 4257 23307 4291
rect 23107 4241 23307 4257
rect 23479 4291 23679 4338
rect 23479 4257 23495 4291
rect 23663 4257 23679 4291
rect 23479 4241 23679 4257
rect 20875 3633 21075 3649
rect 20875 3599 20891 3633
rect 21059 3599 21075 3633
rect 20875 3561 21075 3599
rect 21247 3633 21447 3649
rect 21247 3599 21263 3633
rect 21431 3599 21447 3633
rect 21247 3561 21447 3599
rect 21619 3633 21819 3649
rect 21619 3599 21635 3633
rect 21803 3599 21819 3633
rect 21619 3561 21819 3599
rect 21991 3633 22191 3649
rect 21991 3599 22007 3633
rect 22175 3599 22191 3633
rect 21991 3561 22191 3599
rect 22363 3633 22563 3649
rect 22363 3599 22379 3633
rect 22547 3599 22563 3633
rect 22363 3561 22563 3599
rect 22735 3633 22935 3649
rect 22735 3599 22751 3633
rect 22919 3599 22935 3633
rect 22735 3561 22935 3599
rect 23107 3633 23307 3649
rect 23107 3599 23123 3633
rect 23291 3599 23307 3633
rect 23107 3561 23307 3599
rect 23479 3633 23679 3649
rect 23479 3599 23495 3633
rect 23663 3599 23679 3633
rect 23479 3561 23679 3599
rect 23851 3633 24051 3649
rect 23851 3599 23867 3633
rect 24035 3599 24051 3633
rect 23851 3561 24051 3599
rect 24223 3633 24423 3649
rect 24223 3599 24239 3633
rect 24407 3599 24423 3633
rect 24223 3561 24423 3599
rect 24595 3633 24795 3649
rect 24595 3599 24611 3633
rect 24779 3599 24795 3633
rect 24595 3561 24795 3599
rect 24967 3633 25167 3649
rect 24967 3599 24983 3633
rect 25151 3599 25167 3633
rect 24967 3561 25167 3599
rect 25339 3633 25539 3649
rect 25339 3599 25355 3633
rect 25523 3599 25539 3633
rect 25339 3561 25539 3599
rect 25711 3633 25911 3649
rect 25711 3599 25727 3633
rect 25895 3599 25911 3633
rect 25711 3561 25911 3599
rect 26083 3633 26283 3649
rect 26083 3599 26099 3633
rect 26267 3599 26283 3633
rect 26083 3561 26283 3599
rect 26455 3633 26655 3649
rect 26455 3599 26471 3633
rect 26639 3599 26655 3633
rect 26455 3561 26655 3599
rect 26827 3633 27027 3649
rect 26827 3599 26843 3633
rect 27011 3599 27027 3633
rect 26827 3561 27027 3599
rect 27199 3633 27399 3649
rect 27199 3599 27215 3633
rect 27383 3599 27399 3633
rect 27199 3561 27399 3599
rect 27571 3633 27771 3649
rect 27571 3599 27587 3633
rect 27755 3599 27771 3633
rect 27571 3561 27771 3599
rect 27943 3633 28143 3649
rect 27943 3599 27959 3633
rect 28127 3599 28143 3633
rect 27943 3561 28143 3599
rect 28315 3633 28515 3649
rect 28315 3599 28331 3633
rect 28499 3599 28515 3633
rect 28315 3561 28515 3599
rect 28687 3633 28887 3649
rect 28687 3599 28703 3633
rect 28871 3599 28887 3633
rect 28687 3561 28887 3599
rect 29059 3633 29259 3649
rect 29059 3599 29075 3633
rect 29243 3599 29259 3633
rect 29059 3561 29259 3599
rect 29431 3633 29631 3649
rect 29431 3599 29447 3633
rect 29615 3599 29631 3633
rect 29431 3561 29631 3599
rect 20875 3323 21075 3361
rect 20875 3289 20891 3323
rect 21059 3289 21075 3323
rect 20875 3273 21075 3289
rect 21247 3323 21447 3361
rect 21247 3289 21263 3323
rect 21431 3289 21447 3323
rect 21247 3273 21447 3289
rect 21619 3323 21819 3361
rect 21619 3289 21635 3323
rect 21803 3289 21819 3323
rect 21619 3273 21819 3289
rect 21991 3323 22191 3361
rect 21991 3289 22007 3323
rect 22175 3289 22191 3323
rect 21991 3273 22191 3289
rect 22363 3323 22563 3361
rect 22363 3289 22379 3323
rect 22547 3289 22563 3323
rect 22363 3273 22563 3289
rect 22735 3323 22935 3361
rect 22735 3289 22751 3323
rect 22919 3289 22935 3323
rect 22735 3273 22935 3289
rect 23107 3323 23307 3361
rect 23107 3289 23123 3323
rect 23291 3289 23307 3323
rect 23107 3273 23307 3289
rect 23479 3323 23679 3361
rect 23479 3289 23495 3323
rect 23663 3289 23679 3323
rect 23479 3273 23679 3289
rect 23851 3323 24051 3361
rect 23851 3289 23867 3323
rect 24035 3289 24051 3323
rect 23851 3273 24051 3289
rect 24223 3323 24423 3361
rect 24223 3289 24239 3323
rect 24407 3289 24423 3323
rect 24223 3273 24423 3289
rect 24595 3323 24795 3361
rect 24595 3289 24611 3323
rect 24779 3289 24795 3323
rect 24595 3273 24795 3289
rect 24967 3323 25167 3361
rect 24967 3289 24983 3323
rect 25151 3289 25167 3323
rect 24967 3273 25167 3289
rect 25339 3323 25539 3361
rect 25339 3289 25355 3323
rect 25523 3289 25539 3323
rect 25339 3273 25539 3289
rect 25711 3323 25911 3361
rect 25711 3289 25727 3323
rect 25895 3289 25911 3323
rect 25711 3273 25911 3289
rect 26083 3323 26283 3361
rect 26083 3289 26099 3323
rect 26267 3289 26283 3323
rect 26083 3273 26283 3289
rect 26455 3323 26655 3361
rect 26455 3289 26471 3323
rect 26639 3289 26655 3323
rect 26455 3273 26655 3289
rect 26827 3323 27027 3361
rect 26827 3289 26843 3323
rect 27011 3289 27027 3323
rect 26827 3273 27027 3289
rect 27199 3323 27399 3361
rect 27199 3289 27215 3323
rect 27383 3289 27399 3323
rect 27199 3273 27399 3289
rect 27571 3323 27771 3361
rect 27571 3289 27587 3323
rect 27755 3289 27771 3323
rect 27571 3273 27771 3289
rect 27943 3323 28143 3361
rect 27943 3289 27959 3323
rect 28127 3289 28143 3323
rect 27943 3273 28143 3289
rect 28315 3323 28515 3361
rect 28315 3289 28331 3323
rect 28499 3289 28515 3323
rect 28315 3273 28515 3289
rect 28687 3323 28887 3361
rect 28687 3289 28703 3323
rect 28871 3289 28887 3323
rect 28687 3273 28887 3289
rect 29059 3323 29259 3361
rect 29059 3289 29075 3323
rect 29243 3289 29259 3323
rect 29059 3273 29259 3289
rect 29431 3323 29631 3361
rect 29431 3289 29447 3323
rect 29615 3289 29631 3323
rect 29431 3273 29631 3289
rect 20875 3215 21075 3231
rect 20875 3181 20891 3215
rect 21059 3181 21075 3215
rect 20875 3143 21075 3181
rect 21247 3215 21447 3231
rect 21247 3181 21263 3215
rect 21431 3181 21447 3215
rect 21247 3143 21447 3181
rect 21619 3215 21819 3231
rect 21619 3181 21635 3215
rect 21803 3181 21819 3215
rect 21619 3143 21819 3181
rect 21991 3215 22191 3231
rect 21991 3181 22007 3215
rect 22175 3181 22191 3215
rect 21991 3143 22191 3181
rect 22363 3215 22563 3231
rect 22363 3181 22379 3215
rect 22547 3181 22563 3215
rect 22363 3143 22563 3181
rect 22735 3215 22935 3231
rect 22735 3181 22751 3215
rect 22919 3181 22935 3215
rect 22735 3143 22935 3181
rect 23107 3215 23307 3231
rect 23107 3181 23123 3215
rect 23291 3181 23307 3215
rect 23107 3143 23307 3181
rect 23479 3215 23679 3231
rect 23479 3181 23495 3215
rect 23663 3181 23679 3215
rect 23479 3143 23679 3181
rect 23851 3215 24051 3231
rect 23851 3181 23867 3215
rect 24035 3181 24051 3215
rect 23851 3143 24051 3181
rect 24223 3215 24423 3231
rect 24223 3181 24239 3215
rect 24407 3181 24423 3215
rect 24223 3143 24423 3181
rect 24595 3215 24795 3231
rect 24595 3181 24611 3215
rect 24779 3181 24795 3215
rect 24595 3143 24795 3181
rect 24967 3215 25167 3231
rect 24967 3181 24983 3215
rect 25151 3181 25167 3215
rect 24967 3143 25167 3181
rect 25339 3215 25539 3231
rect 25339 3181 25355 3215
rect 25523 3181 25539 3215
rect 25339 3143 25539 3181
rect 25711 3215 25911 3231
rect 25711 3181 25727 3215
rect 25895 3181 25911 3215
rect 25711 3143 25911 3181
rect 26083 3215 26283 3231
rect 26083 3181 26099 3215
rect 26267 3181 26283 3215
rect 26083 3143 26283 3181
rect 26455 3215 26655 3231
rect 26455 3181 26471 3215
rect 26639 3181 26655 3215
rect 26455 3143 26655 3181
rect 26827 3215 27027 3231
rect 26827 3181 26843 3215
rect 27011 3181 27027 3215
rect 26827 3143 27027 3181
rect 27199 3215 27399 3231
rect 27199 3181 27215 3215
rect 27383 3181 27399 3215
rect 27199 3143 27399 3181
rect 27571 3215 27771 3231
rect 27571 3181 27587 3215
rect 27755 3181 27771 3215
rect 27571 3143 27771 3181
rect 27943 3215 28143 3231
rect 27943 3181 27959 3215
rect 28127 3181 28143 3215
rect 27943 3143 28143 3181
rect 28315 3215 28515 3231
rect 28315 3181 28331 3215
rect 28499 3181 28515 3215
rect 28315 3143 28515 3181
rect 28687 3215 28887 3231
rect 28687 3181 28703 3215
rect 28871 3181 28887 3215
rect 28687 3143 28887 3181
rect 29059 3215 29259 3231
rect 29059 3181 29075 3215
rect 29243 3181 29259 3215
rect 29059 3143 29259 3181
rect 29431 3215 29631 3231
rect 29431 3181 29447 3215
rect 29615 3181 29631 3215
rect 29431 3143 29631 3181
rect 20875 2905 21075 2943
rect 20875 2871 20891 2905
rect 21059 2871 21075 2905
rect 20875 2855 21075 2871
rect 21247 2905 21447 2943
rect 21247 2871 21263 2905
rect 21431 2871 21447 2905
rect 21247 2855 21447 2871
rect 21619 2905 21819 2943
rect 21619 2871 21635 2905
rect 21803 2871 21819 2905
rect 21619 2855 21819 2871
rect 21991 2905 22191 2943
rect 21991 2871 22007 2905
rect 22175 2871 22191 2905
rect 21991 2855 22191 2871
rect 22363 2905 22563 2943
rect 22363 2871 22379 2905
rect 22547 2871 22563 2905
rect 22363 2855 22563 2871
rect 22735 2905 22935 2943
rect 22735 2871 22751 2905
rect 22919 2871 22935 2905
rect 22735 2855 22935 2871
rect 23107 2905 23307 2943
rect 23107 2871 23123 2905
rect 23291 2871 23307 2905
rect 23107 2855 23307 2871
rect 23479 2905 23679 2943
rect 23479 2871 23495 2905
rect 23663 2871 23679 2905
rect 23479 2855 23679 2871
rect 23851 2905 24051 2943
rect 23851 2871 23867 2905
rect 24035 2871 24051 2905
rect 23851 2855 24051 2871
rect 24223 2905 24423 2943
rect 24223 2871 24239 2905
rect 24407 2871 24423 2905
rect 24223 2855 24423 2871
rect 24595 2905 24795 2943
rect 24595 2871 24611 2905
rect 24779 2871 24795 2905
rect 24595 2855 24795 2871
rect 24967 2905 25167 2943
rect 24967 2871 24983 2905
rect 25151 2871 25167 2905
rect 24967 2855 25167 2871
rect 25339 2905 25539 2943
rect 25339 2871 25355 2905
rect 25523 2871 25539 2905
rect 25339 2855 25539 2871
rect 25711 2905 25911 2943
rect 25711 2871 25727 2905
rect 25895 2871 25911 2905
rect 25711 2855 25911 2871
rect 26083 2905 26283 2943
rect 26083 2871 26099 2905
rect 26267 2871 26283 2905
rect 26083 2855 26283 2871
rect 26455 2905 26655 2943
rect 26455 2871 26471 2905
rect 26639 2871 26655 2905
rect 26455 2855 26655 2871
rect 26827 2905 27027 2943
rect 26827 2871 26843 2905
rect 27011 2871 27027 2905
rect 26827 2855 27027 2871
rect 27199 2905 27399 2943
rect 27199 2871 27215 2905
rect 27383 2871 27399 2905
rect 27199 2855 27399 2871
rect 27571 2905 27771 2943
rect 27571 2871 27587 2905
rect 27755 2871 27771 2905
rect 27571 2855 27771 2871
rect 27943 2905 28143 2943
rect 27943 2871 27959 2905
rect 28127 2871 28143 2905
rect 27943 2855 28143 2871
rect 28315 2905 28515 2943
rect 28315 2871 28331 2905
rect 28499 2871 28515 2905
rect 28315 2855 28515 2871
rect 28687 2905 28887 2943
rect 28687 2871 28703 2905
rect 28871 2871 28887 2905
rect 28687 2855 28887 2871
rect 29059 2905 29259 2943
rect 29059 2871 29075 2905
rect 29243 2871 29259 2905
rect 29059 2855 29259 2871
rect 29431 2905 29631 2943
rect 29431 2871 29447 2905
rect 29615 2871 29631 2905
rect 29431 2855 29631 2871
rect 20875 2797 21075 2813
rect 20875 2763 20891 2797
rect 21059 2763 21075 2797
rect 20875 2725 21075 2763
rect 21247 2797 21447 2813
rect 21247 2763 21263 2797
rect 21431 2763 21447 2797
rect 21247 2725 21447 2763
rect 21619 2797 21819 2813
rect 21619 2763 21635 2797
rect 21803 2763 21819 2797
rect 21619 2725 21819 2763
rect 21991 2797 22191 2813
rect 21991 2763 22007 2797
rect 22175 2763 22191 2797
rect 21991 2725 22191 2763
rect 22363 2797 22563 2813
rect 22363 2763 22379 2797
rect 22547 2763 22563 2797
rect 22363 2725 22563 2763
rect 22735 2797 22935 2813
rect 22735 2763 22751 2797
rect 22919 2763 22935 2797
rect 22735 2725 22935 2763
rect 23107 2797 23307 2813
rect 23107 2763 23123 2797
rect 23291 2763 23307 2797
rect 23107 2725 23307 2763
rect 23479 2797 23679 2813
rect 23479 2763 23495 2797
rect 23663 2763 23679 2797
rect 23479 2725 23679 2763
rect 23851 2797 24051 2813
rect 23851 2763 23867 2797
rect 24035 2763 24051 2797
rect 23851 2725 24051 2763
rect 24223 2797 24423 2813
rect 24223 2763 24239 2797
rect 24407 2763 24423 2797
rect 24223 2725 24423 2763
rect 24595 2797 24795 2813
rect 24595 2763 24611 2797
rect 24779 2763 24795 2797
rect 24595 2725 24795 2763
rect 24967 2797 25167 2813
rect 24967 2763 24983 2797
rect 25151 2763 25167 2797
rect 24967 2725 25167 2763
rect 25339 2797 25539 2813
rect 25339 2763 25355 2797
rect 25523 2763 25539 2797
rect 25339 2725 25539 2763
rect 25711 2797 25911 2813
rect 25711 2763 25727 2797
rect 25895 2763 25911 2797
rect 25711 2725 25911 2763
rect 26083 2797 26283 2813
rect 26083 2763 26099 2797
rect 26267 2763 26283 2797
rect 26083 2725 26283 2763
rect 26455 2797 26655 2813
rect 26455 2763 26471 2797
rect 26639 2763 26655 2797
rect 26455 2725 26655 2763
rect 26827 2797 27027 2813
rect 26827 2763 26843 2797
rect 27011 2763 27027 2797
rect 26827 2725 27027 2763
rect 27199 2797 27399 2813
rect 27199 2763 27215 2797
rect 27383 2763 27399 2797
rect 27199 2725 27399 2763
rect 27571 2797 27771 2813
rect 27571 2763 27587 2797
rect 27755 2763 27771 2797
rect 27571 2725 27771 2763
rect 27943 2797 28143 2813
rect 27943 2763 27959 2797
rect 28127 2763 28143 2797
rect 27943 2725 28143 2763
rect 28315 2797 28515 2813
rect 28315 2763 28331 2797
rect 28499 2763 28515 2797
rect 28315 2725 28515 2763
rect 28687 2797 28887 2813
rect 28687 2763 28703 2797
rect 28871 2763 28887 2797
rect 28687 2725 28887 2763
rect 29059 2797 29259 2813
rect 29059 2763 29075 2797
rect 29243 2763 29259 2797
rect 29059 2725 29259 2763
rect 29431 2797 29631 2813
rect 29431 2763 29447 2797
rect 29615 2763 29631 2797
rect 29431 2725 29631 2763
rect 20875 2487 21075 2525
rect 20875 2453 20891 2487
rect 21059 2453 21075 2487
rect 20875 2437 21075 2453
rect 21247 2487 21447 2525
rect 21247 2453 21263 2487
rect 21431 2453 21447 2487
rect 21247 2437 21447 2453
rect 21619 2487 21819 2525
rect 21619 2453 21635 2487
rect 21803 2453 21819 2487
rect 21619 2437 21819 2453
rect 21991 2487 22191 2525
rect 21991 2453 22007 2487
rect 22175 2453 22191 2487
rect 21991 2437 22191 2453
rect 22363 2487 22563 2525
rect 22363 2453 22379 2487
rect 22547 2453 22563 2487
rect 22363 2437 22563 2453
rect 22735 2487 22935 2525
rect 22735 2453 22751 2487
rect 22919 2453 22935 2487
rect 22735 2437 22935 2453
rect 23107 2487 23307 2525
rect 23107 2453 23123 2487
rect 23291 2453 23307 2487
rect 23107 2437 23307 2453
rect 23479 2487 23679 2525
rect 23479 2453 23495 2487
rect 23663 2453 23679 2487
rect 23479 2437 23679 2453
rect 23851 2487 24051 2525
rect 23851 2453 23867 2487
rect 24035 2453 24051 2487
rect 23851 2437 24051 2453
rect 24223 2487 24423 2525
rect 24223 2453 24239 2487
rect 24407 2453 24423 2487
rect 24223 2437 24423 2453
rect 24595 2487 24795 2525
rect 24595 2453 24611 2487
rect 24779 2453 24795 2487
rect 24595 2437 24795 2453
rect 24967 2487 25167 2525
rect 24967 2453 24983 2487
rect 25151 2453 25167 2487
rect 24967 2437 25167 2453
rect 25339 2487 25539 2525
rect 25339 2453 25355 2487
rect 25523 2453 25539 2487
rect 25339 2437 25539 2453
rect 25711 2487 25911 2525
rect 25711 2453 25727 2487
rect 25895 2453 25911 2487
rect 25711 2437 25911 2453
rect 26083 2487 26283 2525
rect 26083 2453 26099 2487
rect 26267 2453 26283 2487
rect 26083 2437 26283 2453
rect 26455 2487 26655 2525
rect 26455 2453 26471 2487
rect 26639 2453 26655 2487
rect 26455 2437 26655 2453
rect 26827 2487 27027 2525
rect 26827 2453 26843 2487
rect 27011 2453 27027 2487
rect 26827 2437 27027 2453
rect 27199 2487 27399 2525
rect 27199 2453 27215 2487
rect 27383 2453 27399 2487
rect 27199 2437 27399 2453
rect 27571 2487 27771 2525
rect 27571 2453 27587 2487
rect 27755 2453 27771 2487
rect 27571 2437 27771 2453
rect 27943 2487 28143 2525
rect 27943 2453 27959 2487
rect 28127 2453 28143 2487
rect 27943 2437 28143 2453
rect 28315 2487 28515 2525
rect 28315 2453 28331 2487
rect 28499 2453 28515 2487
rect 28315 2437 28515 2453
rect 28687 2487 28887 2525
rect 28687 2453 28703 2487
rect 28871 2453 28887 2487
rect 28687 2437 28887 2453
rect 29059 2487 29259 2525
rect 29059 2453 29075 2487
rect 29243 2453 29259 2487
rect 29059 2437 29259 2453
rect 29431 2487 29631 2525
rect 29431 2453 29447 2487
rect 29615 2453 29631 2487
rect 29431 2437 29631 2453
rect 20875 2379 21075 2395
rect 20875 2345 20891 2379
rect 21059 2345 21075 2379
rect 20875 2307 21075 2345
rect 21247 2379 21447 2395
rect 21247 2345 21263 2379
rect 21431 2345 21447 2379
rect 21247 2307 21447 2345
rect 21619 2379 21819 2395
rect 21619 2345 21635 2379
rect 21803 2345 21819 2379
rect 21619 2307 21819 2345
rect 21991 2379 22191 2395
rect 21991 2345 22007 2379
rect 22175 2345 22191 2379
rect 21991 2307 22191 2345
rect 22363 2379 22563 2395
rect 22363 2345 22379 2379
rect 22547 2345 22563 2379
rect 22363 2307 22563 2345
rect 22735 2379 22935 2395
rect 22735 2345 22751 2379
rect 22919 2345 22935 2379
rect 22735 2307 22935 2345
rect 23107 2379 23307 2395
rect 23107 2345 23123 2379
rect 23291 2345 23307 2379
rect 23107 2307 23307 2345
rect 23479 2379 23679 2395
rect 23479 2345 23495 2379
rect 23663 2345 23679 2379
rect 23479 2307 23679 2345
rect 23851 2379 24051 2395
rect 23851 2345 23867 2379
rect 24035 2345 24051 2379
rect 23851 2307 24051 2345
rect 24223 2379 24423 2395
rect 24223 2345 24239 2379
rect 24407 2345 24423 2379
rect 24223 2307 24423 2345
rect 24595 2379 24795 2395
rect 24595 2345 24611 2379
rect 24779 2345 24795 2379
rect 24595 2307 24795 2345
rect 24967 2379 25167 2395
rect 24967 2345 24983 2379
rect 25151 2345 25167 2379
rect 24967 2307 25167 2345
rect 25339 2379 25539 2395
rect 25339 2345 25355 2379
rect 25523 2345 25539 2379
rect 25339 2307 25539 2345
rect 25711 2379 25911 2395
rect 25711 2345 25727 2379
rect 25895 2345 25911 2379
rect 25711 2307 25911 2345
rect 26083 2379 26283 2395
rect 26083 2345 26099 2379
rect 26267 2345 26283 2379
rect 26083 2307 26283 2345
rect 26455 2379 26655 2395
rect 26455 2345 26471 2379
rect 26639 2345 26655 2379
rect 26455 2307 26655 2345
rect 26827 2379 27027 2395
rect 26827 2345 26843 2379
rect 27011 2345 27027 2379
rect 26827 2307 27027 2345
rect 27199 2379 27399 2395
rect 27199 2345 27215 2379
rect 27383 2345 27399 2379
rect 27199 2307 27399 2345
rect 27571 2379 27771 2395
rect 27571 2345 27587 2379
rect 27755 2345 27771 2379
rect 27571 2307 27771 2345
rect 27943 2379 28143 2395
rect 27943 2345 27959 2379
rect 28127 2345 28143 2379
rect 27943 2307 28143 2345
rect 28315 2379 28515 2395
rect 28315 2345 28331 2379
rect 28499 2345 28515 2379
rect 28315 2307 28515 2345
rect 28687 2379 28887 2395
rect 28687 2345 28703 2379
rect 28871 2345 28887 2379
rect 28687 2307 28887 2345
rect 29059 2379 29259 2395
rect 29059 2345 29075 2379
rect 29243 2345 29259 2379
rect 29059 2307 29259 2345
rect 29431 2379 29631 2395
rect 29431 2345 29447 2379
rect 29615 2345 29631 2379
rect 29431 2307 29631 2345
rect 20875 2069 21075 2107
rect 20875 2035 20891 2069
rect 21059 2035 21075 2069
rect 20875 2019 21075 2035
rect 21247 2069 21447 2107
rect 21247 2035 21263 2069
rect 21431 2035 21447 2069
rect 21247 2019 21447 2035
rect 21619 2069 21819 2107
rect 21619 2035 21635 2069
rect 21803 2035 21819 2069
rect 21619 2019 21819 2035
rect 21991 2069 22191 2107
rect 21991 2035 22007 2069
rect 22175 2035 22191 2069
rect 21991 2019 22191 2035
rect 22363 2069 22563 2107
rect 22363 2035 22379 2069
rect 22547 2035 22563 2069
rect 22363 2019 22563 2035
rect 22735 2069 22935 2107
rect 22735 2035 22751 2069
rect 22919 2035 22935 2069
rect 22735 2019 22935 2035
rect 23107 2069 23307 2107
rect 23107 2035 23123 2069
rect 23291 2035 23307 2069
rect 23107 2019 23307 2035
rect 23479 2069 23679 2107
rect 23479 2035 23495 2069
rect 23663 2035 23679 2069
rect 23479 2019 23679 2035
rect 23851 2069 24051 2107
rect 23851 2035 23867 2069
rect 24035 2035 24051 2069
rect 23851 2019 24051 2035
rect 24223 2069 24423 2107
rect 24223 2035 24239 2069
rect 24407 2035 24423 2069
rect 24223 2019 24423 2035
rect 24595 2069 24795 2107
rect 24595 2035 24611 2069
rect 24779 2035 24795 2069
rect 24595 2019 24795 2035
rect 24967 2069 25167 2107
rect 24967 2035 24983 2069
rect 25151 2035 25167 2069
rect 24967 2019 25167 2035
rect 25339 2069 25539 2107
rect 25339 2035 25355 2069
rect 25523 2035 25539 2069
rect 25339 2019 25539 2035
rect 25711 2069 25911 2107
rect 25711 2035 25727 2069
rect 25895 2035 25911 2069
rect 25711 2019 25911 2035
rect 26083 2069 26283 2107
rect 26083 2035 26099 2069
rect 26267 2035 26283 2069
rect 26083 2019 26283 2035
rect 26455 2069 26655 2107
rect 26455 2035 26471 2069
rect 26639 2035 26655 2069
rect 26455 2019 26655 2035
rect 26827 2069 27027 2107
rect 26827 2035 26843 2069
rect 27011 2035 27027 2069
rect 26827 2019 27027 2035
rect 27199 2069 27399 2107
rect 27199 2035 27215 2069
rect 27383 2035 27399 2069
rect 27199 2019 27399 2035
rect 27571 2069 27771 2107
rect 27571 2035 27587 2069
rect 27755 2035 27771 2069
rect 27571 2019 27771 2035
rect 27943 2069 28143 2107
rect 27943 2035 27959 2069
rect 28127 2035 28143 2069
rect 27943 2019 28143 2035
rect 28315 2069 28515 2107
rect 28315 2035 28331 2069
rect 28499 2035 28515 2069
rect 28315 2019 28515 2035
rect 28687 2069 28887 2107
rect 28687 2035 28703 2069
rect 28871 2035 28887 2069
rect 28687 2019 28887 2035
rect 29059 2069 29259 2107
rect 29059 2035 29075 2069
rect 29243 2035 29259 2069
rect 29059 2019 29259 2035
rect 29431 2069 29631 2107
rect 29431 2035 29447 2069
rect 29615 2035 29631 2069
rect 29431 2019 29631 2035
<< polycont >>
rect 19403 10681 19571 10715
rect 19775 10681 19943 10715
rect 20147 10681 20315 10715
rect 20519 10681 20687 10715
rect 20891 10681 21059 10715
rect 21263 10681 21431 10715
rect 21635 10681 21803 10715
rect 22007 10681 22175 10715
rect 22379 10681 22547 10715
rect 22751 10681 22919 10715
rect 23123 10681 23291 10715
rect 23495 10681 23663 10715
rect 23867 10681 24035 10715
rect 24239 10681 24407 10715
rect 24611 10681 24779 10715
rect 24983 10681 25151 10715
rect 25355 10681 25523 10715
rect 25727 10681 25895 10715
rect 26099 10681 26267 10715
rect 26471 10681 26639 10715
rect 26843 10681 27011 10715
rect 27215 10681 27383 10715
rect 27587 10681 27755 10715
rect 27959 10681 28127 10715
rect 28331 10681 28499 10715
rect 28703 10681 28871 10715
rect 29075 10681 29243 10715
rect 29447 10681 29615 10715
rect 29819 10681 29987 10715
rect 30191 10681 30359 10715
rect 30563 10681 30731 10715
rect 30935 10681 31103 10715
rect 19403 10153 19571 10187
rect 19775 10153 19943 10187
rect 20147 10153 20315 10187
rect 20519 10153 20687 10187
rect 20891 10153 21059 10187
rect 21263 10153 21431 10187
rect 21635 10153 21803 10187
rect 22007 10153 22175 10187
rect 22379 10153 22547 10187
rect 22751 10153 22919 10187
rect 23123 10153 23291 10187
rect 23495 10153 23663 10187
rect 23867 10153 24035 10187
rect 24239 10153 24407 10187
rect 24611 10153 24779 10187
rect 24983 10153 25151 10187
rect 25355 10153 25523 10187
rect 25727 10153 25895 10187
rect 26099 10153 26267 10187
rect 26471 10153 26639 10187
rect 26843 10153 27011 10187
rect 27215 10153 27383 10187
rect 27587 10153 27755 10187
rect 27959 10153 28127 10187
rect 28331 10153 28499 10187
rect 28703 10153 28871 10187
rect 29075 10153 29243 10187
rect 29447 10153 29615 10187
rect 29819 10153 29987 10187
rect 30191 10153 30359 10187
rect 30563 10153 30731 10187
rect 30935 10153 31103 10187
rect 19403 10045 19571 10079
rect 19775 10045 19943 10079
rect 20147 10045 20315 10079
rect 20519 10045 20687 10079
rect 20891 10045 21059 10079
rect 21263 10045 21431 10079
rect 21635 10045 21803 10079
rect 22007 10045 22175 10079
rect 22379 10045 22547 10079
rect 22751 10045 22919 10079
rect 23123 10045 23291 10079
rect 23495 10045 23663 10079
rect 23867 10045 24035 10079
rect 24239 10045 24407 10079
rect 24611 10045 24779 10079
rect 24983 10045 25151 10079
rect 25355 10045 25523 10079
rect 25727 10045 25895 10079
rect 26099 10045 26267 10079
rect 26471 10045 26639 10079
rect 26843 10045 27011 10079
rect 27215 10045 27383 10079
rect 27587 10045 27755 10079
rect 27959 10045 28127 10079
rect 28331 10045 28499 10079
rect 28703 10045 28871 10079
rect 29075 10045 29243 10079
rect 29447 10045 29615 10079
rect 29819 10045 29987 10079
rect 30191 10045 30359 10079
rect 30563 10045 30731 10079
rect 30935 10045 31103 10079
rect 19403 9517 19571 9551
rect 19775 9517 19943 9551
rect 20147 9517 20315 9551
rect 20519 9517 20687 9551
rect 20891 9517 21059 9551
rect 21263 9517 21431 9551
rect 21635 9517 21803 9551
rect 22007 9517 22175 9551
rect 22379 9517 22547 9551
rect 22751 9517 22919 9551
rect 23123 9517 23291 9551
rect 23495 9517 23663 9551
rect 23867 9517 24035 9551
rect 24239 9517 24407 9551
rect 24611 9517 24779 9551
rect 24983 9517 25151 9551
rect 25355 9517 25523 9551
rect 25727 9517 25895 9551
rect 26099 9517 26267 9551
rect 26471 9517 26639 9551
rect 26843 9517 27011 9551
rect 27215 9517 27383 9551
rect 27587 9517 27755 9551
rect 27959 9517 28127 9551
rect 28331 9517 28499 9551
rect 28703 9517 28871 9551
rect 29075 9517 29243 9551
rect 29447 9517 29615 9551
rect 29819 9517 29987 9551
rect 30191 9517 30359 9551
rect 30563 9517 30731 9551
rect 30935 9517 31103 9551
rect 19403 9409 19571 9443
rect 19775 9409 19943 9443
rect 20147 9409 20315 9443
rect 20519 9409 20687 9443
rect 20891 9409 21059 9443
rect 21263 9409 21431 9443
rect 21635 9409 21803 9443
rect 22007 9409 22175 9443
rect 22379 9409 22547 9443
rect 22751 9409 22919 9443
rect 23123 9409 23291 9443
rect 23495 9409 23663 9443
rect 23867 9409 24035 9443
rect 24239 9409 24407 9443
rect 24611 9409 24779 9443
rect 24983 9409 25151 9443
rect 25355 9409 25523 9443
rect 25727 9409 25895 9443
rect 26099 9409 26267 9443
rect 26471 9409 26639 9443
rect 26843 9409 27011 9443
rect 27215 9409 27383 9443
rect 27587 9409 27755 9443
rect 27959 9409 28127 9443
rect 28331 9409 28499 9443
rect 28703 9409 28871 9443
rect 29075 9409 29243 9443
rect 29447 9409 29615 9443
rect 29819 9409 29987 9443
rect 30191 9409 30359 9443
rect 30563 9409 30731 9443
rect 30935 9409 31103 9443
rect 19403 8881 19571 8915
rect 19775 8881 19943 8915
rect 20147 8881 20315 8915
rect 20519 8881 20687 8915
rect 20891 8881 21059 8915
rect 21263 8881 21431 8915
rect 21635 8881 21803 8915
rect 22007 8881 22175 8915
rect 22379 8881 22547 8915
rect 22751 8881 22919 8915
rect 23123 8881 23291 8915
rect 23495 8881 23663 8915
rect 23867 8881 24035 8915
rect 24239 8881 24407 8915
rect 24611 8881 24779 8915
rect 24983 8881 25151 8915
rect 25355 8881 25523 8915
rect 25727 8881 25895 8915
rect 26099 8881 26267 8915
rect 26471 8881 26639 8915
rect 26843 8881 27011 8915
rect 27215 8881 27383 8915
rect 27587 8881 27755 8915
rect 27959 8881 28127 8915
rect 28331 8881 28499 8915
rect 28703 8881 28871 8915
rect 29075 8881 29243 8915
rect 29447 8881 29615 8915
rect 29819 8881 29987 8915
rect 30191 8881 30359 8915
rect 30563 8881 30731 8915
rect 30935 8881 31103 8915
rect 20891 8293 21059 8327
rect 21263 8293 21431 8327
rect 21635 8293 21803 8327
rect 22007 8293 22175 8327
rect 22379 8293 22547 8327
rect 22751 8293 22919 8327
rect 23123 8293 23291 8327
rect 23495 8293 23663 8327
rect 20891 7365 21059 7399
rect 21263 7365 21431 7399
rect 21635 7365 21803 7399
rect 22007 7365 22175 7399
rect 22379 7365 22547 7399
rect 22751 7365 22919 7399
rect 23123 7365 23291 7399
rect 23495 7365 23663 7399
rect 20891 7257 21059 7291
rect 21263 7257 21431 7291
rect 21635 7257 21803 7291
rect 22007 7257 22175 7291
rect 22379 7257 22547 7291
rect 22751 7257 22919 7291
rect 23123 7257 23291 7291
rect 23495 7257 23663 7291
rect 20891 6329 21059 6363
rect 21263 6329 21431 6363
rect 21635 6329 21803 6363
rect 22007 6329 22175 6363
rect 22379 6329 22547 6363
rect 22751 6329 22919 6363
rect 23123 6329 23291 6363
rect 23495 6329 23663 6363
rect 20891 6221 21059 6255
rect 21263 6221 21431 6255
rect 21635 6221 21803 6255
rect 22007 6221 22175 6255
rect 22379 6221 22547 6255
rect 22751 6221 22919 6255
rect 23123 6221 23291 6255
rect 23495 6221 23663 6255
rect 20891 5293 21059 5327
rect 21263 5293 21431 5327
rect 21635 5293 21803 5327
rect 22007 5293 22175 5327
rect 22379 5293 22547 5327
rect 22751 5293 22919 5327
rect 23123 5293 23291 5327
rect 23495 5293 23663 5327
rect 20891 5185 21059 5219
rect 21263 5185 21431 5219
rect 21635 5185 21803 5219
rect 22007 5185 22175 5219
rect 22379 5185 22547 5219
rect 22751 5185 22919 5219
rect 23123 5185 23291 5219
rect 23495 5185 23663 5219
rect 20891 4257 21059 4291
rect 21263 4257 21431 4291
rect 21635 4257 21803 4291
rect 22007 4257 22175 4291
rect 22379 4257 22547 4291
rect 22751 4257 22919 4291
rect 23123 4257 23291 4291
rect 23495 4257 23663 4291
rect 20891 3599 21059 3633
rect 21263 3599 21431 3633
rect 21635 3599 21803 3633
rect 22007 3599 22175 3633
rect 22379 3599 22547 3633
rect 22751 3599 22919 3633
rect 23123 3599 23291 3633
rect 23495 3599 23663 3633
rect 23867 3599 24035 3633
rect 24239 3599 24407 3633
rect 24611 3599 24779 3633
rect 24983 3599 25151 3633
rect 25355 3599 25523 3633
rect 25727 3599 25895 3633
rect 26099 3599 26267 3633
rect 26471 3599 26639 3633
rect 26843 3599 27011 3633
rect 27215 3599 27383 3633
rect 27587 3599 27755 3633
rect 27959 3599 28127 3633
rect 28331 3599 28499 3633
rect 28703 3599 28871 3633
rect 29075 3599 29243 3633
rect 29447 3599 29615 3633
rect 20891 3289 21059 3323
rect 21263 3289 21431 3323
rect 21635 3289 21803 3323
rect 22007 3289 22175 3323
rect 22379 3289 22547 3323
rect 22751 3289 22919 3323
rect 23123 3289 23291 3323
rect 23495 3289 23663 3323
rect 23867 3289 24035 3323
rect 24239 3289 24407 3323
rect 24611 3289 24779 3323
rect 24983 3289 25151 3323
rect 25355 3289 25523 3323
rect 25727 3289 25895 3323
rect 26099 3289 26267 3323
rect 26471 3289 26639 3323
rect 26843 3289 27011 3323
rect 27215 3289 27383 3323
rect 27587 3289 27755 3323
rect 27959 3289 28127 3323
rect 28331 3289 28499 3323
rect 28703 3289 28871 3323
rect 29075 3289 29243 3323
rect 29447 3289 29615 3323
rect 20891 3181 21059 3215
rect 21263 3181 21431 3215
rect 21635 3181 21803 3215
rect 22007 3181 22175 3215
rect 22379 3181 22547 3215
rect 22751 3181 22919 3215
rect 23123 3181 23291 3215
rect 23495 3181 23663 3215
rect 23867 3181 24035 3215
rect 24239 3181 24407 3215
rect 24611 3181 24779 3215
rect 24983 3181 25151 3215
rect 25355 3181 25523 3215
rect 25727 3181 25895 3215
rect 26099 3181 26267 3215
rect 26471 3181 26639 3215
rect 26843 3181 27011 3215
rect 27215 3181 27383 3215
rect 27587 3181 27755 3215
rect 27959 3181 28127 3215
rect 28331 3181 28499 3215
rect 28703 3181 28871 3215
rect 29075 3181 29243 3215
rect 29447 3181 29615 3215
rect 20891 2871 21059 2905
rect 21263 2871 21431 2905
rect 21635 2871 21803 2905
rect 22007 2871 22175 2905
rect 22379 2871 22547 2905
rect 22751 2871 22919 2905
rect 23123 2871 23291 2905
rect 23495 2871 23663 2905
rect 23867 2871 24035 2905
rect 24239 2871 24407 2905
rect 24611 2871 24779 2905
rect 24983 2871 25151 2905
rect 25355 2871 25523 2905
rect 25727 2871 25895 2905
rect 26099 2871 26267 2905
rect 26471 2871 26639 2905
rect 26843 2871 27011 2905
rect 27215 2871 27383 2905
rect 27587 2871 27755 2905
rect 27959 2871 28127 2905
rect 28331 2871 28499 2905
rect 28703 2871 28871 2905
rect 29075 2871 29243 2905
rect 29447 2871 29615 2905
rect 20891 2763 21059 2797
rect 21263 2763 21431 2797
rect 21635 2763 21803 2797
rect 22007 2763 22175 2797
rect 22379 2763 22547 2797
rect 22751 2763 22919 2797
rect 23123 2763 23291 2797
rect 23495 2763 23663 2797
rect 23867 2763 24035 2797
rect 24239 2763 24407 2797
rect 24611 2763 24779 2797
rect 24983 2763 25151 2797
rect 25355 2763 25523 2797
rect 25727 2763 25895 2797
rect 26099 2763 26267 2797
rect 26471 2763 26639 2797
rect 26843 2763 27011 2797
rect 27215 2763 27383 2797
rect 27587 2763 27755 2797
rect 27959 2763 28127 2797
rect 28331 2763 28499 2797
rect 28703 2763 28871 2797
rect 29075 2763 29243 2797
rect 29447 2763 29615 2797
rect 20891 2453 21059 2487
rect 21263 2453 21431 2487
rect 21635 2453 21803 2487
rect 22007 2453 22175 2487
rect 22379 2453 22547 2487
rect 22751 2453 22919 2487
rect 23123 2453 23291 2487
rect 23495 2453 23663 2487
rect 23867 2453 24035 2487
rect 24239 2453 24407 2487
rect 24611 2453 24779 2487
rect 24983 2453 25151 2487
rect 25355 2453 25523 2487
rect 25727 2453 25895 2487
rect 26099 2453 26267 2487
rect 26471 2453 26639 2487
rect 26843 2453 27011 2487
rect 27215 2453 27383 2487
rect 27587 2453 27755 2487
rect 27959 2453 28127 2487
rect 28331 2453 28499 2487
rect 28703 2453 28871 2487
rect 29075 2453 29243 2487
rect 29447 2453 29615 2487
rect 20891 2345 21059 2379
rect 21263 2345 21431 2379
rect 21635 2345 21803 2379
rect 22007 2345 22175 2379
rect 22379 2345 22547 2379
rect 22751 2345 22919 2379
rect 23123 2345 23291 2379
rect 23495 2345 23663 2379
rect 23867 2345 24035 2379
rect 24239 2345 24407 2379
rect 24611 2345 24779 2379
rect 24983 2345 25151 2379
rect 25355 2345 25523 2379
rect 25727 2345 25895 2379
rect 26099 2345 26267 2379
rect 26471 2345 26639 2379
rect 26843 2345 27011 2379
rect 27215 2345 27383 2379
rect 27587 2345 27755 2379
rect 27959 2345 28127 2379
rect 28331 2345 28499 2379
rect 28703 2345 28871 2379
rect 29075 2345 29243 2379
rect 29447 2345 29615 2379
rect 20891 2035 21059 2069
rect 21263 2035 21431 2069
rect 21635 2035 21803 2069
rect 22007 2035 22175 2069
rect 22379 2035 22547 2069
rect 22751 2035 22919 2069
rect 23123 2035 23291 2069
rect 23495 2035 23663 2069
rect 23867 2035 24035 2069
rect 24239 2035 24407 2069
rect 24611 2035 24779 2069
rect 24983 2035 25151 2069
rect 25355 2035 25523 2069
rect 25727 2035 25895 2069
rect 26099 2035 26267 2069
rect 26471 2035 26639 2069
rect 26843 2035 27011 2069
rect 27215 2035 27383 2069
rect 27587 2035 27755 2069
rect 27959 2035 28127 2069
rect 28331 2035 28499 2069
rect 28703 2035 28871 2069
rect 29075 2035 29243 2069
rect 29447 2035 29615 2069
<< locali >>
rect 19227 10783 19323 10817
rect 31186 10783 31279 10817
rect 19227 10721 19261 10783
rect 31245 10721 31279 10783
rect 19387 10681 19403 10715
rect 19571 10681 19587 10715
rect 19759 10681 19775 10715
rect 19943 10681 19959 10715
rect 20131 10681 20147 10715
rect 20315 10681 20331 10715
rect 20503 10681 20519 10715
rect 20687 10681 20703 10715
rect 20875 10681 20891 10715
rect 21059 10681 21075 10715
rect 21247 10681 21263 10715
rect 21431 10681 21447 10715
rect 21619 10681 21635 10715
rect 21803 10681 21819 10715
rect 21991 10681 22007 10715
rect 22175 10681 22191 10715
rect 22363 10681 22379 10715
rect 22547 10681 22563 10715
rect 22735 10681 22751 10715
rect 22919 10681 22935 10715
rect 23107 10681 23123 10715
rect 23291 10681 23307 10715
rect 23479 10681 23495 10715
rect 23663 10681 23679 10715
rect 23851 10681 23867 10715
rect 24035 10681 24051 10715
rect 24223 10681 24239 10715
rect 24407 10681 24423 10715
rect 24595 10681 24611 10715
rect 24779 10681 24795 10715
rect 24967 10681 24983 10715
rect 25151 10681 25167 10715
rect 25339 10681 25355 10715
rect 25523 10681 25539 10715
rect 25711 10681 25727 10715
rect 25895 10681 25911 10715
rect 26083 10681 26099 10715
rect 26267 10681 26283 10715
rect 26455 10681 26471 10715
rect 26639 10681 26655 10715
rect 26827 10681 26843 10715
rect 27011 10681 27027 10715
rect 27199 10681 27215 10715
rect 27383 10681 27399 10715
rect 27571 10681 27587 10715
rect 27755 10681 27771 10715
rect 27943 10681 27959 10715
rect 28127 10681 28143 10715
rect 28315 10681 28331 10715
rect 28499 10681 28515 10715
rect 28687 10681 28703 10715
rect 28871 10681 28887 10715
rect 29059 10681 29075 10715
rect 29243 10681 29259 10715
rect 29431 10681 29447 10715
rect 29615 10681 29631 10715
rect 29803 10681 29819 10715
rect 29987 10681 30003 10715
rect 30175 10681 30191 10715
rect 30359 10681 30375 10715
rect 30547 10681 30563 10715
rect 30731 10681 30747 10715
rect 30919 10681 30935 10715
rect 31103 10681 31119 10715
rect 19341 10622 19375 10638
rect 19341 10230 19375 10246
rect 19599 10622 19633 10638
rect 19599 10230 19633 10246
rect 19713 10622 19747 10638
rect 19713 10230 19747 10246
rect 19971 10622 20005 10638
rect 19971 10230 20005 10246
rect 20085 10622 20119 10638
rect 20085 10230 20119 10246
rect 20343 10622 20377 10638
rect 20343 10230 20377 10246
rect 20457 10622 20491 10638
rect 20457 10230 20491 10246
rect 20715 10622 20749 10638
rect 20715 10230 20749 10246
rect 20829 10622 20863 10638
rect 20829 10230 20863 10246
rect 21087 10622 21121 10638
rect 21087 10230 21121 10246
rect 21201 10622 21235 10638
rect 21201 10230 21235 10246
rect 21459 10622 21493 10638
rect 21459 10230 21493 10246
rect 21573 10622 21607 10638
rect 21573 10230 21607 10246
rect 21831 10622 21865 10638
rect 21831 10230 21865 10246
rect 21945 10622 21979 10638
rect 21945 10230 21979 10246
rect 22203 10622 22237 10638
rect 22203 10230 22237 10246
rect 22317 10622 22351 10638
rect 22317 10230 22351 10246
rect 22575 10622 22609 10638
rect 22575 10230 22609 10246
rect 22689 10622 22723 10638
rect 22689 10230 22723 10246
rect 22947 10622 22981 10638
rect 22947 10230 22981 10246
rect 23061 10622 23095 10638
rect 23061 10230 23095 10246
rect 23319 10622 23353 10638
rect 23319 10230 23353 10246
rect 23433 10622 23467 10638
rect 23433 10230 23467 10246
rect 23691 10622 23725 10638
rect 23691 10230 23725 10246
rect 23805 10622 23839 10638
rect 23805 10230 23839 10246
rect 24063 10622 24097 10638
rect 24063 10230 24097 10246
rect 24177 10622 24211 10638
rect 24177 10230 24211 10246
rect 24435 10622 24469 10638
rect 24435 10230 24469 10246
rect 24549 10622 24583 10638
rect 24549 10230 24583 10246
rect 24807 10622 24841 10638
rect 24807 10230 24841 10246
rect 24921 10622 24955 10638
rect 24921 10230 24955 10246
rect 25179 10622 25213 10638
rect 25179 10230 25213 10246
rect 25293 10622 25327 10638
rect 25293 10230 25327 10246
rect 25551 10622 25585 10638
rect 25551 10230 25585 10246
rect 25665 10622 25699 10638
rect 25665 10230 25699 10246
rect 25923 10622 25957 10638
rect 25923 10230 25957 10246
rect 26037 10622 26071 10638
rect 26037 10230 26071 10246
rect 26295 10622 26329 10638
rect 26295 10230 26329 10246
rect 26409 10622 26443 10638
rect 26409 10230 26443 10246
rect 26667 10622 26701 10638
rect 26667 10230 26701 10246
rect 26781 10622 26815 10638
rect 26781 10230 26815 10246
rect 27039 10622 27073 10638
rect 27039 10230 27073 10246
rect 27153 10622 27187 10638
rect 27153 10230 27187 10246
rect 27411 10622 27445 10638
rect 27411 10230 27445 10246
rect 27525 10622 27559 10638
rect 27525 10230 27559 10246
rect 27783 10622 27817 10638
rect 27783 10230 27817 10246
rect 27897 10622 27931 10638
rect 27897 10230 27931 10246
rect 28155 10622 28189 10638
rect 28155 10230 28189 10246
rect 28269 10622 28303 10638
rect 28269 10230 28303 10246
rect 28527 10622 28561 10638
rect 28527 10230 28561 10246
rect 28641 10622 28675 10638
rect 28641 10230 28675 10246
rect 28899 10622 28933 10638
rect 28899 10230 28933 10246
rect 29013 10622 29047 10638
rect 29013 10230 29047 10246
rect 29271 10622 29305 10638
rect 29271 10230 29305 10246
rect 29385 10622 29419 10638
rect 29385 10230 29419 10246
rect 29643 10622 29677 10638
rect 29643 10230 29677 10246
rect 29757 10622 29791 10638
rect 29757 10230 29791 10246
rect 30015 10622 30049 10638
rect 30015 10230 30049 10246
rect 30129 10622 30163 10638
rect 30129 10230 30163 10246
rect 30387 10622 30421 10638
rect 30387 10230 30421 10246
rect 30501 10622 30535 10638
rect 30501 10230 30535 10246
rect 30759 10622 30793 10638
rect 30759 10230 30793 10246
rect 30873 10622 30907 10638
rect 30873 10230 30907 10246
rect 31131 10622 31165 10638
rect 31131 10230 31165 10246
rect 19387 10153 19403 10187
rect 19571 10153 19587 10187
rect 19759 10153 19775 10187
rect 19943 10153 19959 10187
rect 20131 10153 20147 10187
rect 20315 10153 20331 10187
rect 20503 10153 20519 10187
rect 20687 10153 20703 10187
rect 20875 10153 20891 10187
rect 21059 10153 21075 10187
rect 21247 10153 21263 10187
rect 21431 10153 21447 10187
rect 21619 10153 21635 10187
rect 21803 10153 21819 10187
rect 21991 10153 22007 10187
rect 22175 10153 22191 10187
rect 22363 10153 22379 10187
rect 22547 10153 22563 10187
rect 22735 10153 22751 10187
rect 22919 10153 22935 10187
rect 23107 10153 23123 10187
rect 23291 10153 23307 10187
rect 23479 10153 23495 10187
rect 23663 10153 23679 10187
rect 23851 10153 23867 10187
rect 24035 10153 24051 10187
rect 24223 10153 24239 10187
rect 24407 10153 24423 10187
rect 24595 10153 24611 10187
rect 24779 10153 24795 10187
rect 24967 10153 24983 10187
rect 25151 10153 25167 10187
rect 25339 10153 25355 10187
rect 25523 10153 25539 10187
rect 25711 10153 25727 10187
rect 25895 10153 25911 10187
rect 26083 10153 26099 10187
rect 26267 10153 26283 10187
rect 26455 10153 26471 10187
rect 26639 10153 26655 10187
rect 26827 10153 26843 10187
rect 27011 10153 27027 10187
rect 27199 10153 27215 10187
rect 27383 10153 27399 10187
rect 27571 10153 27587 10187
rect 27755 10153 27771 10187
rect 27943 10153 27959 10187
rect 28127 10153 28143 10187
rect 28315 10153 28331 10187
rect 28499 10153 28515 10187
rect 28687 10153 28703 10187
rect 28871 10153 28887 10187
rect 29059 10153 29075 10187
rect 29243 10153 29259 10187
rect 29431 10153 29447 10187
rect 29615 10153 29631 10187
rect 29803 10153 29819 10187
rect 29987 10153 30003 10187
rect 30175 10153 30191 10187
rect 30359 10153 30375 10187
rect 30547 10153 30563 10187
rect 30731 10153 30747 10187
rect 30919 10153 30935 10187
rect 31103 10153 31119 10187
rect 19387 10045 19403 10079
rect 19571 10045 19587 10079
rect 19759 10045 19775 10079
rect 19943 10045 19959 10079
rect 20131 10045 20147 10079
rect 20315 10045 20331 10079
rect 20503 10045 20519 10079
rect 20687 10045 20703 10079
rect 20875 10045 20891 10079
rect 21059 10045 21075 10079
rect 21247 10045 21263 10079
rect 21431 10045 21447 10079
rect 21619 10045 21635 10079
rect 21803 10045 21819 10079
rect 21991 10045 22007 10079
rect 22175 10045 22191 10079
rect 22363 10045 22379 10079
rect 22547 10045 22563 10079
rect 22735 10045 22751 10079
rect 22919 10045 22935 10079
rect 23107 10045 23123 10079
rect 23291 10045 23307 10079
rect 23479 10045 23495 10079
rect 23663 10045 23679 10079
rect 23851 10045 23867 10079
rect 24035 10045 24051 10079
rect 24223 10045 24239 10079
rect 24407 10045 24423 10079
rect 24595 10045 24611 10079
rect 24779 10045 24795 10079
rect 24967 10045 24983 10079
rect 25151 10045 25167 10079
rect 25339 10045 25355 10079
rect 25523 10045 25539 10079
rect 25711 10045 25727 10079
rect 25895 10045 25911 10079
rect 26083 10045 26099 10079
rect 26267 10045 26283 10079
rect 26455 10045 26471 10079
rect 26639 10045 26655 10079
rect 26827 10045 26843 10079
rect 27011 10045 27027 10079
rect 27199 10045 27215 10079
rect 27383 10045 27399 10079
rect 27571 10045 27587 10079
rect 27755 10045 27771 10079
rect 27943 10045 27959 10079
rect 28127 10045 28143 10079
rect 28315 10045 28331 10079
rect 28499 10045 28515 10079
rect 28687 10045 28703 10079
rect 28871 10045 28887 10079
rect 29059 10045 29075 10079
rect 29243 10045 29259 10079
rect 29431 10045 29447 10079
rect 29615 10045 29631 10079
rect 29803 10045 29819 10079
rect 29987 10045 30003 10079
rect 30175 10045 30191 10079
rect 30359 10045 30375 10079
rect 30547 10045 30563 10079
rect 30731 10045 30747 10079
rect 30919 10045 30935 10079
rect 31103 10045 31119 10079
rect 19341 9986 19375 10002
rect 19341 9594 19375 9610
rect 19599 9986 19633 10002
rect 19599 9594 19633 9610
rect 19713 9986 19747 10002
rect 19713 9594 19747 9610
rect 19971 9986 20005 10002
rect 19971 9594 20005 9610
rect 20085 9986 20119 10002
rect 20085 9594 20119 9610
rect 20343 9986 20377 10002
rect 20343 9594 20377 9610
rect 20457 9986 20491 10002
rect 20457 9594 20491 9610
rect 20715 9986 20749 10002
rect 20715 9594 20749 9610
rect 20829 9986 20863 10002
rect 20829 9594 20863 9610
rect 21087 9986 21121 10002
rect 21087 9594 21121 9610
rect 21201 9986 21235 10002
rect 21201 9594 21235 9610
rect 21459 9986 21493 10002
rect 21459 9594 21493 9610
rect 21573 9986 21607 10002
rect 21573 9594 21607 9610
rect 21831 9986 21865 10002
rect 21831 9594 21865 9610
rect 21945 9986 21979 10002
rect 21945 9594 21979 9610
rect 22203 9986 22237 10002
rect 22203 9594 22237 9610
rect 22317 9986 22351 10002
rect 22317 9594 22351 9610
rect 22575 9986 22609 10002
rect 22575 9594 22609 9610
rect 22689 9986 22723 10002
rect 22689 9594 22723 9610
rect 22947 9986 22981 10002
rect 22947 9594 22981 9610
rect 23061 9986 23095 10002
rect 23061 9594 23095 9610
rect 23319 9986 23353 10002
rect 23319 9594 23353 9610
rect 23433 9986 23467 10002
rect 23433 9594 23467 9610
rect 23691 9986 23725 10002
rect 23691 9594 23725 9610
rect 23805 9986 23839 10002
rect 23805 9594 23839 9610
rect 24063 9986 24097 10002
rect 24063 9594 24097 9610
rect 24177 9986 24211 10002
rect 24177 9594 24211 9610
rect 24435 9986 24469 10002
rect 24435 9594 24469 9610
rect 24549 9986 24583 10002
rect 24549 9594 24583 9610
rect 24807 9986 24841 10002
rect 24807 9594 24841 9610
rect 24921 9986 24955 10002
rect 24921 9594 24955 9610
rect 25179 9986 25213 10002
rect 25179 9594 25213 9610
rect 25293 9986 25327 10002
rect 25293 9594 25327 9610
rect 25551 9986 25585 10002
rect 25551 9594 25585 9610
rect 25665 9986 25699 10002
rect 25665 9594 25699 9610
rect 25923 9986 25957 10002
rect 25923 9594 25957 9610
rect 26037 9986 26071 10002
rect 26037 9594 26071 9610
rect 26295 9986 26329 10002
rect 26295 9594 26329 9610
rect 26409 9986 26443 10002
rect 26409 9594 26443 9610
rect 26667 9986 26701 10002
rect 26667 9594 26701 9610
rect 26781 9986 26815 10002
rect 26781 9594 26815 9610
rect 27039 9986 27073 10002
rect 27039 9594 27073 9610
rect 27153 9986 27187 10002
rect 27153 9594 27187 9610
rect 27411 9986 27445 10002
rect 27411 9594 27445 9610
rect 27525 9986 27559 10002
rect 27525 9594 27559 9610
rect 27783 9986 27817 10002
rect 27783 9594 27817 9610
rect 27897 9986 27931 10002
rect 27897 9594 27931 9610
rect 28155 9986 28189 10002
rect 28155 9594 28189 9610
rect 28269 9986 28303 10002
rect 28269 9594 28303 9610
rect 28527 9986 28561 10002
rect 28527 9594 28561 9610
rect 28641 9986 28675 10002
rect 28641 9594 28675 9610
rect 28899 9986 28933 10002
rect 28899 9594 28933 9610
rect 29013 9986 29047 10002
rect 29013 9594 29047 9610
rect 29271 9986 29305 10002
rect 29271 9594 29305 9610
rect 29385 9986 29419 10002
rect 29385 9594 29419 9610
rect 29643 9986 29677 10002
rect 29643 9594 29677 9610
rect 29757 9986 29791 10002
rect 29757 9594 29791 9610
rect 30015 9986 30049 10002
rect 30015 9594 30049 9610
rect 30129 9986 30163 10002
rect 30129 9594 30163 9610
rect 30387 9986 30421 10002
rect 30387 9594 30421 9610
rect 30501 9986 30535 10002
rect 30501 9594 30535 9610
rect 30759 9986 30793 10002
rect 30759 9594 30793 9610
rect 30873 9986 30907 10002
rect 30873 9594 30907 9610
rect 31131 9986 31165 10002
rect 31131 9594 31165 9610
rect 19387 9517 19403 9551
rect 19571 9517 19587 9551
rect 19759 9517 19775 9551
rect 19943 9517 19959 9551
rect 20131 9517 20147 9551
rect 20315 9517 20331 9551
rect 20503 9517 20519 9551
rect 20687 9517 20703 9551
rect 20875 9517 20891 9551
rect 21059 9517 21075 9551
rect 21247 9517 21263 9551
rect 21431 9517 21447 9551
rect 21619 9517 21635 9551
rect 21803 9517 21819 9551
rect 21991 9517 22007 9551
rect 22175 9517 22191 9551
rect 22363 9517 22379 9551
rect 22547 9517 22563 9551
rect 22735 9517 22751 9551
rect 22919 9517 22935 9551
rect 23107 9517 23123 9551
rect 23291 9517 23307 9551
rect 23479 9517 23495 9551
rect 23663 9517 23679 9551
rect 23851 9517 23867 9551
rect 24035 9517 24051 9551
rect 24223 9517 24239 9551
rect 24407 9517 24423 9551
rect 24595 9517 24611 9551
rect 24779 9517 24795 9551
rect 24967 9517 24983 9551
rect 25151 9517 25167 9551
rect 25339 9517 25355 9551
rect 25523 9517 25539 9551
rect 25711 9517 25727 9551
rect 25895 9517 25911 9551
rect 26083 9517 26099 9551
rect 26267 9517 26283 9551
rect 26455 9517 26471 9551
rect 26639 9517 26655 9551
rect 26827 9517 26843 9551
rect 27011 9517 27027 9551
rect 27199 9517 27215 9551
rect 27383 9517 27399 9551
rect 27571 9517 27587 9551
rect 27755 9517 27771 9551
rect 27943 9517 27959 9551
rect 28127 9517 28143 9551
rect 28315 9517 28331 9551
rect 28499 9517 28515 9551
rect 28687 9517 28703 9551
rect 28871 9517 28887 9551
rect 29059 9517 29075 9551
rect 29243 9517 29259 9551
rect 29431 9517 29447 9551
rect 29615 9517 29631 9551
rect 29803 9517 29819 9551
rect 29987 9517 30003 9551
rect 30175 9517 30191 9551
rect 30359 9517 30375 9551
rect 30547 9517 30563 9551
rect 30731 9517 30747 9551
rect 30919 9517 30935 9551
rect 31103 9517 31119 9551
rect 19387 9409 19403 9443
rect 19571 9409 19587 9443
rect 19759 9409 19775 9443
rect 19943 9409 19959 9443
rect 20131 9409 20147 9443
rect 20315 9409 20331 9443
rect 20503 9409 20519 9443
rect 20687 9409 20703 9443
rect 20875 9409 20891 9443
rect 21059 9409 21075 9443
rect 21247 9409 21263 9443
rect 21431 9409 21447 9443
rect 21619 9409 21635 9443
rect 21803 9409 21819 9443
rect 21991 9409 22007 9443
rect 22175 9409 22191 9443
rect 22363 9409 22379 9443
rect 22547 9409 22563 9443
rect 22735 9409 22751 9443
rect 22919 9409 22935 9443
rect 23107 9409 23123 9443
rect 23291 9409 23307 9443
rect 23479 9409 23495 9443
rect 23663 9409 23679 9443
rect 23851 9409 23867 9443
rect 24035 9409 24051 9443
rect 24223 9409 24239 9443
rect 24407 9409 24423 9443
rect 24595 9409 24611 9443
rect 24779 9409 24795 9443
rect 24967 9409 24983 9443
rect 25151 9409 25167 9443
rect 25339 9409 25355 9443
rect 25523 9409 25539 9443
rect 25711 9409 25727 9443
rect 25895 9409 25911 9443
rect 26083 9409 26099 9443
rect 26267 9409 26283 9443
rect 26455 9409 26471 9443
rect 26639 9409 26655 9443
rect 26827 9409 26843 9443
rect 27011 9409 27027 9443
rect 27199 9409 27215 9443
rect 27383 9409 27399 9443
rect 27571 9409 27587 9443
rect 27755 9409 27771 9443
rect 27943 9409 27959 9443
rect 28127 9409 28143 9443
rect 28315 9409 28331 9443
rect 28499 9409 28515 9443
rect 28687 9409 28703 9443
rect 28871 9409 28887 9443
rect 29059 9409 29075 9443
rect 29243 9409 29259 9443
rect 29431 9409 29447 9443
rect 29615 9409 29631 9443
rect 29803 9409 29819 9443
rect 29987 9409 30003 9443
rect 30175 9409 30191 9443
rect 30359 9409 30375 9443
rect 30547 9409 30563 9443
rect 30731 9409 30747 9443
rect 30919 9409 30935 9443
rect 31103 9409 31119 9443
rect 19341 9350 19375 9366
rect 19341 8958 19375 8974
rect 19599 9350 19633 9366
rect 19599 8958 19633 8974
rect 19713 9350 19747 9366
rect 19713 8958 19747 8974
rect 19971 9350 20005 9366
rect 19971 8958 20005 8974
rect 20085 9350 20119 9366
rect 20085 8958 20119 8974
rect 20343 9350 20377 9366
rect 20343 8958 20377 8974
rect 20457 9350 20491 9366
rect 20457 8958 20491 8974
rect 20715 9350 20749 9366
rect 20715 8958 20749 8974
rect 20829 9350 20863 9366
rect 20829 8958 20863 8974
rect 21087 9350 21121 9366
rect 21087 8958 21121 8974
rect 21201 9350 21235 9366
rect 21201 8958 21235 8974
rect 21459 9350 21493 9366
rect 21459 8958 21493 8974
rect 21573 9350 21607 9366
rect 21573 8958 21607 8974
rect 21831 9350 21865 9366
rect 21831 8958 21865 8974
rect 21945 9350 21979 9366
rect 21945 8958 21979 8974
rect 22203 9350 22237 9366
rect 22203 8958 22237 8974
rect 22317 9350 22351 9366
rect 22317 8958 22351 8974
rect 22575 9350 22609 9366
rect 22575 8958 22609 8974
rect 22689 9350 22723 9366
rect 22689 8958 22723 8974
rect 22947 9350 22981 9366
rect 22947 8958 22981 8974
rect 23061 9350 23095 9366
rect 23061 8958 23095 8974
rect 23319 9350 23353 9366
rect 23319 8958 23353 8974
rect 23433 9350 23467 9366
rect 23433 8958 23467 8974
rect 23691 9350 23725 9366
rect 23691 8958 23725 8974
rect 23805 9350 23839 9366
rect 23805 8958 23839 8974
rect 24063 9350 24097 9366
rect 24063 8958 24097 8974
rect 24177 9350 24211 9366
rect 24177 8958 24211 8974
rect 24435 9350 24469 9366
rect 24435 8958 24469 8974
rect 24549 9350 24583 9366
rect 24549 8958 24583 8974
rect 24807 9350 24841 9366
rect 24807 8958 24841 8974
rect 24921 9350 24955 9366
rect 24921 8958 24955 8974
rect 25179 9350 25213 9366
rect 25179 8958 25213 8974
rect 25293 9350 25327 9366
rect 25293 8958 25327 8974
rect 25551 9350 25585 9366
rect 25551 8958 25585 8974
rect 25665 9350 25699 9366
rect 25665 8958 25699 8974
rect 25923 9350 25957 9366
rect 25923 8958 25957 8974
rect 26037 9350 26071 9366
rect 26037 8958 26071 8974
rect 26295 9350 26329 9366
rect 26295 8958 26329 8974
rect 26409 9350 26443 9366
rect 26409 8958 26443 8974
rect 26667 9350 26701 9366
rect 26667 8958 26701 8974
rect 26781 9350 26815 9366
rect 26781 8958 26815 8974
rect 27039 9350 27073 9366
rect 27039 8958 27073 8974
rect 27153 9350 27187 9366
rect 27153 8958 27187 8974
rect 27411 9350 27445 9366
rect 27411 8958 27445 8974
rect 27525 9350 27559 9366
rect 27525 8958 27559 8974
rect 27783 9350 27817 9366
rect 27783 8958 27817 8974
rect 27897 9350 27931 9366
rect 27897 8958 27931 8974
rect 28155 9350 28189 9366
rect 28155 8958 28189 8974
rect 28269 9350 28303 9366
rect 28269 8958 28303 8974
rect 28527 9350 28561 9366
rect 28527 8958 28561 8974
rect 28641 9350 28675 9366
rect 28641 8958 28675 8974
rect 28899 9350 28933 9366
rect 28899 8958 28933 8974
rect 29013 9350 29047 9366
rect 29013 8958 29047 8974
rect 29271 9350 29305 9366
rect 29271 8958 29305 8974
rect 29385 9350 29419 9366
rect 29385 8958 29419 8974
rect 29643 9350 29677 9366
rect 29643 8958 29677 8974
rect 29757 9350 29791 9366
rect 29757 8958 29791 8974
rect 30015 9350 30049 9366
rect 30015 8958 30049 8974
rect 30129 9350 30163 9366
rect 30129 8958 30163 8974
rect 30387 9350 30421 9366
rect 30387 8958 30421 8974
rect 30501 9350 30535 9366
rect 30501 8958 30535 8974
rect 30759 9350 30793 9366
rect 30759 8958 30793 8974
rect 30873 9350 30907 9366
rect 30873 8958 30907 8974
rect 31131 9350 31165 9366
rect 31131 8958 31165 8974
rect 19387 8881 19403 8915
rect 19571 8881 19587 8915
rect 19759 8881 19775 8915
rect 19943 8881 19959 8915
rect 20131 8881 20147 8915
rect 20315 8881 20331 8915
rect 20503 8881 20519 8915
rect 20687 8881 20703 8915
rect 20875 8881 20891 8915
rect 21059 8881 21075 8915
rect 21247 8881 21263 8915
rect 21431 8881 21447 8915
rect 21619 8881 21635 8915
rect 21803 8881 21819 8915
rect 21991 8881 22007 8915
rect 22175 8881 22191 8915
rect 22363 8881 22379 8915
rect 22547 8881 22563 8915
rect 22735 8881 22751 8915
rect 22919 8881 22935 8915
rect 23107 8881 23123 8915
rect 23291 8881 23307 8915
rect 23479 8881 23495 8915
rect 23663 8881 23679 8915
rect 23851 8881 23867 8915
rect 24035 8881 24051 8915
rect 24223 8881 24239 8915
rect 24407 8881 24423 8915
rect 24595 8881 24611 8915
rect 24779 8881 24795 8915
rect 24967 8881 24983 8915
rect 25151 8881 25167 8915
rect 25339 8881 25355 8915
rect 25523 8881 25539 8915
rect 25711 8881 25727 8915
rect 25895 8881 25911 8915
rect 26083 8881 26099 8915
rect 26267 8881 26283 8915
rect 26455 8881 26471 8915
rect 26639 8881 26655 8915
rect 26827 8881 26843 8915
rect 27011 8881 27027 8915
rect 27199 8881 27215 8915
rect 27383 8881 27399 8915
rect 27571 8881 27587 8915
rect 27755 8881 27771 8915
rect 27943 8881 27959 8915
rect 28127 8881 28143 8915
rect 28315 8881 28331 8915
rect 28499 8881 28515 8915
rect 28687 8881 28703 8915
rect 28871 8881 28887 8915
rect 29059 8881 29075 8915
rect 29243 8881 29259 8915
rect 29431 8881 29447 8915
rect 29615 8881 29631 8915
rect 29803 8881 29819 8915
rect 29987 8881 30003 8915
rect 30175 8881 30191 8915
rect 30359 8881 30375 8915
rect 30547 8881 30563 8915
rect 30731 8881 30747 8915
rect 30919 8881 30935 8915
rect 31103 8881 31119 8915
rect 19227 8813 19261 8875
rect 31245 8813 31279 8875
rect 19227 8779 19323 8813
rect 31183 8779 31279 8813
rect 20715 8395 20800 8429
rect 23743 8395 23839 8429
rect 20715 8333 20749 8395
rect 23805 8333 23839 8395
rect 20875 8293 20891 8327
rect 21059 8293 21075 8327
rect 21247 8293 21263 8327
rect 21431 8293 21447 8327
rect 21619 8293 21635 8327
rect 21803 8293 21819 8327
rect 21991 8293 22007 8327
rect 22175 8293 22191 8327
rect 22363 8293 22379 8327
rect 22547 8293 22563 8327
rect 22735 8293 22751 8327
rect 22919 8293 22935 8327
rect 23107 8293 23123 8327
rect 23291 8293 23307 8327
rect 23479 8293 23495 8327
rect 23663 8293 23679 8327
rect 20829 8234 20863 8250
rect 20829 7442 20863 7458
rect 21087 8234 21121 8250
rect 21087 7442 21121 7458
rect 21201 8234 21235 8250
rect 21201 7442 21235 7458
rect 21459 8234 21493 8250
rect 21459 7442 21493 7458
rect 21573 8234 21607 8250
rect 21573 7442 21607 7458
rect 21831 8234 21865 8250
rect 21831 7442 21865 7458
rect 21945 8234 21979 8250
rect 21945 7442 21979 7458
rect 22203 8234 22237 8250
rect 22203 7442 22237 7458
rect 22317 8234 22351 8250
rect 22317 7442 22351 7458
rect 22575 8234 22609 8250
rect 22575 7442 22609 7458
rect 22689 8234 22723 8250
rect 22689 7442 22723 7458
rect 22947 8234 22981 8250
rect 22947 7442 22981 7458
rect 23061 8234 23095 8250
rect 23061 7442 23095 7458
rect 23319 8234 23353 8250
rect 23319 7442 23353 7458
rect 23433 8234 23467 8250
rect 23433 7442 23467 7458
rect 23691 8234 23725 8250
rect 23691 7442 23725 7458
rect 20875 7365 20891 7399
rect 21059 7365 21075 7399
rect 21247 7365 21263 7399
rect 21431 7365 21447 7399
rect 21619 7365 21635 7399
rect 21803 7365 21819 7399
rect 21991 7365 22007 7399
rect 22175 7365 22191 7399
rect 22363 7365 22379 7399
rect 22547 7365 22563 7399
rect 22735 7365 22751 7399
rect 22919 7365 22935 7399
rect 23107 7365 23123 7399
rect 23291 7365 23307 7399
rect 23479 7365 23495 7399
rect 23663 7365 23679 7399
rect 20875 7257 20891 7291
rect 21059 7257 21075 7291
rect 21247 7257 21263 7291
rect 21431 7257 21447 7291
rect 21619 7257 21635 7291
rect 21803 7257 21819 7291
rect 21991 7257 22007 7291
rect 22175 7257 22191 7291
rect 22363 7257 22379 7291
rect 22547 7257 22563 7291
rect 22735 7257 22751 7291
rect 22919 7257 22935 7291
rect 23107 7257 23123 7291
rect 23291 7257 23307 7291
rect 23479 7257 23495 7291
rect 23663 7257 23679 7291
rect 20829 7198 20863 7214
rect 20829 6406 20863 6422
rect 21087 7198 21121 7214
rect 21087 6406 21121 6422
rect 21201 7198 21235 7214
rect 21201 6406 21235 6422
rect 21459 7198 21493 7214
rect 21459 6406 21493 6422
rect 21573 7198 21607 7214
rect 21573 6406 21607 6422
rect 21831 7198 21865 7214
rect 21831 6406 21865 6422
rect 21945 7198 21979 7214
rect 21945 6406 21979 6422
rect 22203 7198 22237 7214
rect 22203 6406 22237 6422
rect 22317 7198 22351 7214
rect 22317 6406 22351 6422
rect 22575 7198 22609 7214
rect 22575 6406 22609 6422
rect 22689 7198 22723 7214
rect 22689 6406 22723 6422
rect 22947 7198 22981 7214
rect 22947 6406 22981 6422
rect 23061 7198 23095 7214
rect 23061 6406 23095 6422
rect 23319 7198 23353 7214
rect 23319 6406 23353 6422
rect 23433 7198 23467 7214
rect 23433 6406 23467 6422
rect 23691 7198 23725 7214
rect 23691 6406 23725 6422
rect 20875 6329 20891 6363
rect 21059 6329 21075 6363
rect 21247 6329 21263 6363
rect 21431 6329 21447 6363
rect 21619 6329 21635 6363
rect 21803 6329 21819 6363
rect 21991 6329 22007 6363
rect 22175 6329 22191 6363
rect 22363 6329 22379 6363
rect 22547 6329 22563 6363
rect 22735 6329 22751 6363
rect 22919 6329 22935 6363
rect 23107 6329 23123 6363
rect 23291 6329 23307 6363
rect 23479 6329 23495 6363
rect 23663 6329 23679 6363
rect 20875 6221 20891 6255
rect 21059 6221 21075 6255
rect 21247 6221 21263 6255
rect 21431 6221 21447 6255
rect 21619 6221 21635 6255
rect 21803 6221 21819 6255
rect 21991 6221 22007 6255
rect 22175 6221 22191 6255
rect 22363 6221 22379 6255
rect 22547 6221 22563 6255
rect 22735 6221 22751 6255
rect 22919 6221 22935 6255
rect 23107 6221 23123 6255
rect 23291 6221 23307 6255
rect 23479 6221 23495 6255
rect 23663 6221 23679 6255
rect 20829 6162 20863 6178
rect 20829 5370 20863 5386
rect 21087 6162 21121 6178
rect 21087 5370 21121 5386
rect 21201 6162 21235 6178
rect 21201 5370 21235 5386
rect 21459 6162 21493 6178
rect 21459 5370 21493 5386
rect 21573 6162 21607 6178
rect 21573 5370 21607 5386
rect 21831 6162 21865 6178
rect 21831 5370 21865 5386
rect 21945 6162 21979 6178
rect 21945 5370 21979 5386
rect 22203 6162 22237 6178
rect 22203 5370 22237 5386
rect 22317 6162 22351 6178
rect 22317 5370 22351 5386
rect 22575 6162 22609 6178
rect 22575 5370 22609 5386
rect 22689 6162 22723 6178
rect 22689 5370 22723 5386
rect 22947 6162 22981 6178
rect 22947 5370 22981 5386
rect 23061 6162 23095 6178
rect 23061 5370 23095 5386
rect 23319 6162 23353 6178
rect 23319 5370 23353 5386
rect 23433 6162 23467 6178
rect 23433 5370 23467 5386
rect 23691 6162 23725 6178
rect 23691 5370 23725 5386
rect 20875 5293 20891 5327
rect 21059 5293 21075 5327
rect 21247 5293 21263 5327
rect 21431 5293 21447 5327
rect 21619 5293 21635 5327
rect 21803 5293 21819 5327
rect 21991 5293 22007 5327
rect 22175 5293 22191 5327
rect 22363 5293 22379 5327
rect 22547 5293 22563 5327
rect 22735 5293 22751 5327
rect 22919 5293 22935 5327
rect 23107 5293 23123 5327
rect 23291 5293 23307 5327
rect 23479 5293 23495 5327
rect 23663 5293 23679 5327
rect 20875 5185 20891 5219
rect 21059 5185 21075 5219
rect 21247 5185 21263 5219
rect 21431 5185 21447 5219
rect 21619 5185 21635 5219
rect 21803 5185 21819 5219
rect 21991 5185 22007 5219
rect 22175 5185 22191 5219
rect 22363 5185 22379 5219
rect 22547 5185 22563 5219
rect 22735 5185 22751 5219
rect 22919 5185 22935 5219
rect 23107 5185 23123 5219
rect 23291 5185 23307 5219
rect 23479 5185 23495 5219
rect 23663 5185 23679 5219
rect 20829 5126 20863 5142
rect 20829 4334 20863 4350
rect 21087 5126 21121 5142
rect 21087 4334 21121 4350
rect 21201 5126 21235 5142
rect 21201 4334 21235 4350
rect 21459 5126 21493 5142
rect 21459 4334 21493 4350
rect 21573 5126 21607 5142
rect 21573 4334 21607 4350
rect 21831 5126 21865 5142
rect 21831 4334 21865 4350
rect 21945 5126 21979 5142
rect 21945 4334 21979 4350
rect 22203 5126 22237 5142
rect 22203 4334 22237 4350
rect 22317 5126 22351 5142
rect 22317 4334 22351 4350
rect 22575 5126 22609 5142
rect 22575 4334 22609 4350
rect 22689 5126 22723 5142
rect 22689 4334 22723 4350
rect 22947 5126 22981 5142
rect 22947 4334 22981 4350
rect 23061 5126 23095 5142
rect 23061 4334 23095 4350
rect 23319 5126 23353 5142
rect 23319 4334 23353 4350
rect 23433 5126 23467 5142
rect 23433 4334 23467 4350
rect 23691 5126 23725 5142
rect 23691 4334 23725 4350
rect 20875 4257 20891 4291
rect 21059 4257 21075 4291
rect 21247 4257 21263 4291
rect 21431 4257 21447 4291
rect 21619 4257 21635 4291
rect 21803 4257 21819 4291
rect 21991 4257 22007 4291
rect 22175 4257 22191 4291
rect 22363 4257 22379 4291
rect 22547 4257 22563 4291
rect 22735 4257 22751 4291
rect 22919 4257 22935 4291
rect 23107 4257 23123 4291
rect 23291 4257 23307 4291
rect 23479 4257 23495 4291
rect 23663 4257 23679 4291
rect 20715 4189 20749 4251
rect 23805 4189 23839 4251
rect 20715 4155 20811 4189
rect 23743 4155 23839 4189
rect 20715 3701 20811 3735
rect 29695 3701 29791 3735
rect 20715 3639 20749 3701
rect 29757 3639 29791 3701
rect 20875 3599 20891 3633
rect 21059 3599 21075 3633
rect 21247 3599 21263 3633
rect 21431 3599 21447 3633
rect 21619 3599 21635 3633
rect 21803 3599 21819 3633
rect 21991 3599 22007 3633
rect 22175 3599 22191 3633
rect 22363 3599 22379 3633
rect 22547 3599 22563 3633
rect 22735 3599 22751 3633
rect 22919 3599 22935 3633
rect 23107 3599 23123 3633
rect 23291 3599 23307 3633
rect 23479 3599 23495 3633
rect 23663 3599 23679 3633
rect 23851 3599 23867 3633
rect 24035 3599 24051 3633
rect 24223 3599 24239 3633
rect 24407 3599 24423 3633
rect 24595 3599 24611 3633
rect 24779 3599 24795 3633
rect 24967 3599 24983 3633
rect 25151 3599 25167 3633
rect 25339 3599 25355 3633
rect 25523 3599 25539 3633
rect 25711 3599 25727 3633
rect 25895 3599 25911 3633
rect 26083 3599 26099 3633
rect 26267 3599 26283 3633
rect 26455 3599 26471 3633
rect 26639 3599 26655 3633
rect 26827 3599 26843 3633
rect 27011 3599 27027 3633
rect 27199 3599 27215 3633
rect 27383 3599 27399 3633
rect 27571 3599 27587 3633
rect 27755 3599 27771 3633
rect 27943 3599 27959 3633
rect 28127 3599 28143 3633
rect 28315 3599 28331 3633
rect 28499 3599 28515 3633
rect 28687 3599 28703 3633
rect 28871 3599 28887 3633
rect 29059 3599 29075 3633
rect 29243 3599 29259 3633
rect 29431 3599 29447 3633
rect 29615 3599 29631 3633
rect 20829 3549 20863 3565
rect 20829 3357 20863 3373
rect 21087 3549 21121 3565
rect 21087 3357 21121 3373
rect 21201 3549 21235 3565
rect 21201 3357 21235 3373
rect 21459 3549 21493 3565
rect 21459 3357 21493 3373
rect 21573 3549 21607 3565
rect 21573 3357 21607 3373
rect 21831 3549 21865 3565
rect 21831 3357 21865 3373
rect 21945 3549 21979 3565
rect 21945 3357 21979 3373
rect 22203 3549 22237 3565
rect 22203 3357 22237 3373
rect 22317 3549 22351 3565
rect 22317 3357 22351 3373
rect 22575 3549 22609 3565
rect 22575 3357 22609 3373
rect 22689 3549 22723 3565
rect 22689 3357 22723 3373
rect 22947 3549 22981 3565
rect 22947 3357 22981 3373
rect 23061 3549 23095 3565
rect 23061 3357 23095 3373
rect 23319 3549 23353 3565
rect 23319 3357 23353 3373
rect 23433 3549 23467 3565
rect 23433 3357 23467 3373
rect 23691 3549 23725 3565
rect 23691 3357 23725 3373
rect 23805 3549 23839 3565
rect 23805 3357 23839 3373
rect 24063 3549 24097 3565
rect 24063 3357 24097 3373
rect 24177 3549 24211 3565
rect 24177 3357 24211 3373
rect 24435 3549 24469 3565
rect 24435 3357 24469 3373
rect 24549 3549 24583 3565
rect 24549 3357 24583 3373
rect 24807 3549 24841 3565
rect 24807 3357 24841 3373
rect 24921 3549 24955 3565
rect 24921 3357 24955 3373
rect 25179 3549 25213 3565
rect 25179 3357 25213 3373
rect 25293 3549 25327 3565
rect 25293 3357 25327 3373
rect 25551 3549 25585 3565
rect 25551 3357 25585 3373
rect 25665 3549 25699 3565
rect 25665 3357 25699 3373
rect 25923 3549 25957 3565
rect 25923 3357 25957 3373
rect 26037 3549 26071 3565
rect 26037 3357 26071 3373
rect 26295 3549 26329 3565
rect 26295 3357 26329 3373
rect 26409 3549 26443 3565
rect 26409 3357 26443 3373
rect 26667 3549 26701 3565
rect 26667 3357 26701 3373
rect 26781 3549 26815 3565
rect 26781 3357 26815 3373
rect 27039 3549 27073 3565
rect 27039 3357 27073 3373
rect 27153 3549 27187 3565
rect 27153 3357 27187 3373
rect 27411 3549 27445 3565
rect 27411 3357 27445 3373
rect 27525 3549 27559 3565
rect 27525 3357 27559 3373
rect 27783 3549 27817 3565
rect 27783 3357 27817 3373
rect 27897 3549 27931 3565
rect 27897 3357 27931 3373
rect 28155 3549 28189 3565
rect 28155 3357 28189 3373
rect 28269 3549 28303 3565
rect 28269 3357 28303 3373
rect 28527 3549 28561 3565
rect 28527 3357 28561 3373
rect 28641 3549 28675 3565
rect 28641 3357 28675 3373
rect 28899 3549 28933 3565
rect 28899 3357 28933 3373
rect 29013 3549 29047 3565
rect 29013 3357 29047 3373
rect 29271 3549 29305 3565
rect 29271 3357 29305 3373
rect 29385 3549 29419 3565
rect 29385 3357 29419 3373
rect 29643 3549 29677 3565
rect 29643 3357 29677 3373
rect 20875 3289 20891 3323
rect 21059 3289 21075 3323
rect 21247 3289 21263 3323
rect 21431 3289 21447 3323
rect 21619 3289 21635 3323
rect 21803 3289 21819 3323
rect 21991 3289 22007 3323
rect 22175 3289 22191 3323
rect 22363 3289 22379 3323
rect 22547 3289 22563 3323
rect 22735 3289 22751 3323
rect 22919 3289 22935 3323
rect 23107 3289 23123 3323
rect 23291 3289 23307 3323
rect 23479 3289 23495 3323
rect 23663 3289 23679 3323
rect 23851 3289 23867 3323
rect 24035 3289 24051 3323
rect 24223 3289 24239 3323
rect 24407 3289 24423 3323
rect 24595 3289 24611 3323
rect 24779 3289 24795 3323
rect 24967 3289 24983 3323
rect 25151 3289 25167 3323
rect 25339 3289 25355 3323
rect 25523 3289 25539 3323
rect 25711 3289 25727 3323
rect 25895 3289 25911 3323
rect 26083 3289 26099 3323
rect 26267 3289 26283 3323
rect 26455 3289 26471 3323
rect 26639 3289 26655 3323
rect 26827 3289 26843 3323
rect 27011 3289 27027 3323
rect 27199 3289 27215 3323
rect 27383 3289 27399 3323
rect 27571 3289 27587 3323
rect 27755 3289 27771 3323
rect 27943 3289 27959 3323
rect 28127 3289 28143 3323
rect 28315 3289 28331 3323
rect 28499 3289 28515 3323
rect 28687 3289 28703 3323
rect 28871 3289 28887 3323
rect 29059 3289 29075 3323
rect 29243 3289 29259 3323
rect 29431 3289 29447 3323
rect 29615 3289 29631 3323
rect 20875 3181 20891 3215
rect 21059 3181 21075 3215
rect 21247 3181 21263 3215
rect 21431 3181 21447 3215
rect 21619 3181 21635 3215
rect 21803 3181 21819 3215
rect 21991 3181 22007 3215
rect 22175 3181 22191 3215
rect 22363 3181 22379 3215
rect 22547 3181 22563 3215
rect 22735 3181 22751 3215
rect 22919 3181 22935 3215
rect 23107 3181 23123 3215
rect 23291 3181 23307 3215
rect 23479 3181 23495 3215
rect 23663 3181 23679 3215
rect 23851 3181 23867 3215
rect 24035 3181 24051 3215
rect 24223 3181 24239 3215
rect 24407 3181 24423 3215
rect 24595 3181 24611 3215
rect 24779 3181 24795 3215
rect 24967 3181 24983 3215
rect 25151 3181 25167 3215
rect 25339 3181 25355 3215
rect 25523 3181 25539 3215
rect 25711 3181 25727 3215
rect 25895 3181 25911 3215
rect 26083 3181 26099 3215
rect 26267 3181 26283 3215
rect 26455 3181 26471 3215
rect 26639 3181 26655 3215
rect 26827 3181 26843 3215
rect 27011 3181 27027 3215
rect 27199 3181 27215 3215
rect 27383 3181 27399 3215
rect 27571 3181 27587 3215
rect 27755 3181 27771 3215
rect 27943 3181 27959 3215
rect 28127 3181 28143 3215
rect 28315 3181 28331 3215
rect 28499 3181 28515 3215
rect 28687 3181 28703 3215
rect 28871 3181 28887 3215
rect 29059 3181 29075 3215
rect 29243 3181 29259 3215
rect 29431 3181 29447 3215
rect 29615 3181 29631 3215
rect 20829 3131 20863 3147
rect 20829 2939 20863 2955
rect 21087 3131 21121 3147
rect 21087 2939 21121 2955
rect 21201 3131 21235 3147
rect 21201 2939 21235 2955
rect 21459 3131 21493 3147
rect 21459 2939 21493 2955
rect 21573 3131 21607 3147
rect 21573 2939 21607 2955
rect 21831 3131 21865 3147
rect 21831 2939 21865 2955
rect 21945 3131 21979 3147
rect 21945 2939 21979 2955
rect 22203 3131 22237 3147
rect 22203 2939 22237 2955
rect 22317 3131 22351 3147
rect 22317 2939 22351 2955
rect 22575 3131 22609 3147
rect 22575 2939 22609 2955
rect 22689 3131 22723 3147
rect 22689 2939 22723 2955
rect 22947 3131 22981 3147
rect 22947 2939 22981 2955
rect 23061 3131 23095 3147
rect 23061 2939 23095 2955
rect 23319 3131 23353 3147
rect 23319 2939 23353 2955
rect 23433 3131 23467 3147
rect 23433 2939 23467 2955
rect 23691 3131 23725 3147
rect 23691 2939 23725 2955
rect 23805 3131 23839 3147
rect 23805 2939 23839 2955
rect 24063 3131 24097 3147
rect 24063 2939 24097 2955
rect 24177 3131 24211 3147
rect 24177 2939 24211 2955
rect 24435 3131 24469 3147
rect 24435 2939 24469 2955
rect 24549 3131 24583 3147
rect 24549 2939 24583 2955
rect 24807 3131 24841 3147
rect 24807 2939 24841 2955
rect 24921 3131 24955 3147
rect 24921 2939 24955 2955
rect 25179 3131 25213 3147
rect 25179 2939 25213 2955
rect 25293 3131 25327 3147
rect 25293 2939 25327 2955
rect 25551 3131 25585 3147
rect 25551 2939 25585 2955
rect 25665 3131 25699 3147
rect 25665 2939 25699 2955
rect 25923 3131 25957 3147
rect 25923 2939 25957 2955
rect 26037 3131 26071 3147
rect 26037 2939 26071 2955
rect 26295 3131 26329 3147
rect 26295 2939 26329 2955
rect 26409 3131 26443 3147
rect 26409 2939 26443 2955
rect 26667 3131 26701 3147
rect 26667 2939 26701 2955
rect 26781 3131 26815 3147
rect 26781 2939 26815 2955
rect 27039 3131 27073 3147
rect 27039 2939 27073 2955
rect 27153 3131 27187 3147
rect 27153 2939 27187 2955
rect 27411 3131 27445 3147
rect 27411 2939 27445 2955
rect 27525 3131 27559 3147
rect 27525 2939 27559 2955
rect 27783 3131 27817 3147
rect 27783 2939 27817 2955
rect 27897 3131 27931 3147
rect 27897 2939 27931 2955
rect 28155 3131 28189 3147
rect 28155 2939 28189 2955
rect 28269 3131 28303 3147
rect 28269 2939 28303 2955
rect 28527 3131 28561 3147
rect 28527 2939 28561 2955
rect 28641 3131 28675 3147
rect 28641 2939 28675 2955
rect 28899 3131 28933 3147
rect 28899 2939 28933 2955
rect 29013 3131 29047 3147
rect 29013 2939 29047 2955
rect 29271 3131 29305 3147
rect 29271 2939 29305 2955
rect 29385 3131 29419 3147
rect 29385 2939 29419 2955
rect 29643 3131 29677 3147
rect 29643 2939 29677 2955
rect 20875 2871 20891 2905
rect 21059 2871 21075 2905
rect 21247 2871 21263 2905
rect 21431 2871 21447 2905
rect 21619 2871 21635 2905
rect 21803 2871 21819 2905
rect 21991 2871 22007 2905
rect 22175 2871 22191 2905
rect 22363 2871 22379 2905
rect 22547 2871 22563 2905
rect 22735 2871 22751 2905
rect 22919 2871 22935 2905
rect 23107 2871 23123 2905
rect 23291 2871 23307 2905
rect 23479 2871 23495 2905
rect 23663 2871 23679 2905
rect 23851 2871 23867 2905
rect 24035 2871 24051 2905
rect 24223 2871 24239 2905
rect 24407 2871 24423 2905
rect 24595 2871 24611 2905
rect 24779 2871 24795 2905
rect 24967 2871 24983 2905
rect 25151 2871 25167 2905
rect 25339 2871 25355 2905
rect 25523 2871 25539 2905
rect 25711 2871 25727 2905
rect 25895 2871 25911 2905
rect 26083 2871 26099 2905
rect 26267 2871 26283 2905
rect 26455 2871 26471 2905
rect 26639 2871 26655 2905
rect 26827 2871 26843 2905
rect 27011 2871 27027 2905
rect 27199 2871 27215 2905
rect 27383 2871 27399 2905
rect 27571 2871 27587 2905
rect 27755 2871 27771 2905
rect 27943 2871 27959 2905
rect 28127 2871 28143 2905
rect 28315 2871 28331 2905
rect 28499 2871 28515 2905
rect 28687 2871 28703 2905
rect 28871 2871 28887 2905
rect 29059 2871 29075 2905
rect 29243 2871 29259 2905
rect 29431 2871 29447 2905
rect 29615 2871 29631 2905
rect 20875 2763 20891 2797
rect 21059 2763 21075 2797
rect 21247 2763 21263 2797
rect 21431 2763 21447 2797
rect 21619 2763 21635 2797
rect 21803 2763 21819 2797
rect 21991 2763 22007 2797
rect 22175 2763 22191 2797
rect 22363 2763 22379 2797
rect 22547 2763 22563 2797
rect 22735 2763 22751 2797
rect 22919 2763 22935 2797
rect 23107 2763 23123 2797
rect 23291 2763 23307 2797
rect 23479 2763 23495 2797
rect 23663 2763 23679 2797
rect 23851 2763 23867 2797
rect 24035 2763 24051 2797
rect 24223 2763 24239 2797
rect 24407 2763 24423 2797
rect 24595 2763 24611 2797
rect 24779 2763 24795 2797
rect 24967 2763 24983 2797
rect 25151 2763 25167 2797
rect 25339 2763 25355 2797
rect 25523 2763 25539 2797
rect 25711 2763 25727 2797
rect 25895 2763 25911 2797
rect 26083 2763 26099 2797
rect 26267 2763 26283 2797
rect 26455 2763 26471 2797
rect 26639 2763 26655 2797
rect 26827 2763 26843 2797
rect 27011 2763 27027 2797
rect 27199 2763 27215 2797
rect 27383 2763 27399 2797
rect 27571 2763 27587 2797
rect 27755 2763 27771 2797
rect 27943 2763 27959 2797
rect 28127 2763 28143 2797
rect 28315 2763 28331 2797
rect 28499 2763 28515 2797
rect 28687 2763 28703 2797
rect 28871 2763 28887 2797
rect 29059 2763 29075 2797
rect 29243 2763 29259 2797
rect 29431 2763 29447 2797
rect 29615 2763 29631 2797
rect 20829 2713 20863 2729
rect 20829 2521 20863 2537
rect 21087 2713 21121 2729
rect 21087 2521 21121 2537
rect 21201 2713 21235 2729
rect 21201 2521 21235 2537
rect 21459 2713 21493 2729
rect 21459 2521 21493 2537
rect 21573 2713 21607 2729
rect 21573 2521 21607 2537
rect 21831 2713 21865 2729
rect 21831 2521 21865 2537
rect 21945 2713 21979 2729
rect 21945 2521 21979 2537
rect 22203 2713 22237 2729
rect 22203 2521 22237 2537
rect 22317 2713 22351 2729
rect 22317 2521 22351 2537
rect 22575 2713 22609 2729
rect 22575 2521 22609 2537
rect 22689 2713 22723 2729
rect 22689 2521 22723 2537
rect 22947 2713 22981 2729
rect 22947 2521 22981 2537
rect 23061 2713 23095 2729
rect 23061 2521 23095 2537
rect 23319 2713 23353 2729
rect 23319 2521 23353 2537
rect 23433 2713 23467 2729
rect 23433 2521 23467 2537
rect 23691 2713 23725 2729
rect 23691 2521 23725 2537
rect 23805 2713 23839 2729
rect 23805 2521 23839 2537
rect 24063 2713 24097 2729
rect 24063 2521 24097 2537
rect 24177 2713 24211 2729
rect 24177 2521 24211 2537
rect 24435 2713 24469 2729
rect 24435 2521 24469 2537
rect 24549 2713 24583 2729
rect 24549 2521 24583 2537
rect 24807 2713 24841 2729
rect 24807 2521 24841 2537
rect 24921 2713 24955 2729
rect 24921 2521 24955 2537
rect 25179 2713 25213 2729
rect 25179 2521 25213 2537
rect 25293 2713 25327 2729
rect 25293 2521 25327 2537
rect 25551 2713 25585 2729
rect 25551 2521 25585 2537
rect 25665 2713 25699 2729
rect 25665 2521 25699 2537
rect 25923 2713 25957 2729
rect 25923 2521 25957 2537
rect 26037 2713 26071 2729
rect 26037 2521 26071 2537
rect 26295 2713 26329 2729
rect 26295 2521 26329 2537
rect 26409 2713 26443 2729
rect 26409 2521 26443 2537
rect 26667 2713 26701 2729
rect 26667 2521 26701 2537
rect 26781 2713 26815 2729
rect 26781 2521 26815 2537
rect 27039 2713 27073 2729
rect 27039 2521 27073 2537
rect 27153 2713 27187 2729
rect 27153 2521 27187 2537
rect 27411 2713 27445 2729
rect 27411 2521 27445 2537
rect 27525 2713 27559 2729
rect 27525 2521 27559 2537
rect 27783 2713 27817 2729
rect 27783 2521 27817 2537
rect 27897 2713 27931 2729
rect 27897 2521 27931 2537
rect 28155 2713 28189 2729
rect 28155 2521 28189 2537
rect 28269 2713 28303 2729
rect 28269 2521 28303 2537
rect 28527 2713 28561 2729
rect 28527 2521 28561 2537
rect 28641 2713 28675 2729
rect 28641 2521 28675 2537
rect 28899 2713 28933 2729
rect 28899 2521 28933 2537
rect 29013 2713 29047 2729
rect 29013 2521 29047 2537
rect 29271 2713 29305 2729
rect 29271 2521 29305 2537
rect 29385 2713 29419 2729
rect 29385 2521 29419 2537
rect 29643 2713 29677 2729
rect 29643 2521 29677 2537
rect 20875 2453 20891 2487
rect 21059 2453 21075 2487
rect 21247 2453 21263 2487
rect 21431 2453 21447 2487
rect 21619 2453 21635 2487
rect 21803 2453 21819 2487
rect 21991 2453 22007 2487
rect 22175 2453 22191 2487
rect 22363 2453 22379 2487
rect 22547 2453 22563 2487
rect 22735 2453 22751 2487
rect 22919 2453 22935 2487
rect 23107 2453 23123 2487
rect 23291 2453 23307 2487
rect 23479 2453 23495 2487
rect 23663 2453 23679 2487
rect 23851 2453 23867 2487
rect 24035 2453 24051 2487
rect 24223 2453 24239 2487
rect 24407 2453 24423 2487
rect 24595 2453 24611 2487
rect 24779 2453 24795 2487
rect 24967 2453 24983 2487
rect 25151 2453 25167 2487
rect 25339 2453 25355 2487
rect 25523 2453 25539 2487
rect 25711 2453 25727 2487
rect 25895 2453 25911 2487
rect 26083 2453 26099 2487
rect 26267 2453 26283 2487
rect 26455 2453 26471 2487
rect 26639 2453 26655 2487
rect 26827 2453 26843 2487
rect 27011 2453 27027 2487
rect 27199 2453 27215 2487
rect 27383 2453 27399 2487
rect 27571 2453 27587 2487
rect 27755 2453 27771 2487
rect 27943 2453 27959 2487
rect 28127 2453 28143 2487
rect 28315 2453 28331 2487
rect 28499 2453 28515 2487
rect 28687 2453 28703 2487
rect 28871 2453 28887 2487
rect 29059 2453 29075 2487
rect 29243 2453 29259 2487
rect 29431 2453 29447 2487
rect 29615 2453 29631 2487
rect 20875 2345 20891 2379
rect 21059 2345 21075 2379
rect 21247 2345 21263 2379
rect 21431 2345 21447 2379
rect 21619 2345 21635 2379
rect 21803 2345 21819 2379
rect 21991 2345 22007 2379
rect 22175 2345 22191 2379
rect 22363 2345 22379 2379
rect 22547 2345 22563 2379
rect 22735 2345 22751 2379
rect 22919 2345 22935 2379
rect 23107 2345 23123 2379
rect 23291 2345 23307 2379
rect 23479 2345 23495 2379
rect 23663 2345 23679 2379
rect 23851 2345 23867 2379
rect 24035 2345 24051 2379
rect 24223 2345 24239 2379
rect 24407 2345 24423 2379
rect 24595 2345 24611 2379
rect 24779 2345 24795 2379
rect 24967 2345 24983 2379
rect 25151 2345 25167 2379
rect 25339 2345 25355 2379
rect 25523 2345 25539 2379
rect 25711 2345 25727 2379
rect 25895 2345 25911 2379
rect 26083 2345 26099 2379
rect 26267 2345 26283 2379
rect 26455 2345 26471 2379
rect 26639 2345 26655 2379
rect 26827 2345 26843 2379
rect 27011 2345 27027 2379
rect 27199 2345 27215 2379
rect 27383 2345 27399 2379
rect 27571 2345 27587 2379
rect 27755 2345 27771 2379
rect 27943 2345 27959 2379
rect 28127 2345 28143 2379
rect 28315 2345 28331 2379
rect 28499 2345 28515 2379
rect 28687 2345 28703 2379
rect 28871 2345 28887 2379
rect 29059 2345 29075 2379
rect 29243 2345 29259 2379
rect 29431 2345 29447 2379
rect 29615 2345 29631 2379
rect 20829 2295 20863 2311
rect 20829 2103 20863 2119
rect 21087 2295 21121 2311
rect 21087 2103 21121 2119
rect 21201 2295 21235 2311
rect 21201 2103 21235 2119
rect 21459 2295 21493 2311
rect 21459 2103 21493 2119
rect 21573 2295 21607 2311
rect 21573 2103 21607 2119
rect 21831 2295 21865 2311
rect 21831 2103 21865 2119
rect 21945 2295 21979 2311
rect 21945 2103 21979 2119
rect 22203 2295 22237 2311
rect 22203 2103 22237 2119
rect 22317 2295 22351 2311
rect 22317 2103 22351 2119
rect 22575 2295 22609 2311
rect 22575 2103 22609 2119
rect 22689 2295 22723 2311
rect 22689 2103 22723 2119
rect 22947 2295 22981 2311
rect 22947 2103 22981 2119
rect 23061 2295 23095 2311
rect 23061 2103 23095 2119
rect 23319 2295 23353 2311
rect 23319 2103 23353 2119
rect 23433 2295 23467 2311
rect 23433 2103 23467 2119
rect 23691 2295 23725 2311
rect 23691 2103 23725 2119
rect 23805 2295 23839 2311
rect 23805 2103 23839 2119
rect 24063 2295 24097 2311
rect 24063 2103 24097 2119
rect 24177 2295 24211 2311
rect 24177 2103 24211 2119
rect 24435 2295 24469 2311
rect 24435 2103 24469 2119
rect 24549 2295 24583 2311
rect 24549 2103 24583 2119
rect 24807 2295 24841 2311
rect 24807 2103 24841 2119
rect 24921 2295 24955 2311
rect 24921 2103 24955 2119
rect 25179 2295 25213 2311
rect 25179 2103 25213 2119
rect 25293 2295 25327 2311
rect 25293 2103 25327 2119
rect 25551 2295 25585 2311
rect 25551 2103 25585 2119
rect 25665 2295 25699 2311
rect 25665 2103 25699 2119
rect 25923 2295 25957 2311
rect 25923 2103 25957 2119
rect 26037 2295 26071 2311
rect 26037 2103 26071 2119
rect 26295 2295 26329 2311
rect 26295 2103 26329 2119
rect 26409 2295 26443 2311
rect 26409 2103 26443 2119
rect 26667 2295 26701 2311
rect 26667 2103 26701 2119
rect 26781 2295 26815 2311
rect 26781 2103 26815 2119
rect 27039 2295 27073 2311
rect 27039 2103 27073 2119
rect 27153 2295 27187 2311
rect 27153 2103 27187 2119
rect 27411 2295 27445 2311
rect 27411 2103 27445 2119
rect 27525 2295 27559 2311
rect 27525 2103 27559 2119
rect 27783 2295 27817 2311
rect 27783 2103 27817 2119
rect 27897 2295 27931 2311
rect 27897 2103 27931 2119
rect 28155 2295 28189 2311
rect 28155 2103 28189 2119
rect 28269 2295 28303 2311
rect 28269 2103 28303 2119
rect 28527 2295 28561 2311
rect 28527 2103 28561 2119
rect 28641 2295 28675 2311
rect 28641 2103 28675 2119
rect 28899 2295 28933 2311
rect 28899 2103 28933 2119
rect 29013 2295 29047 2311
rect 29013 2103 29047 2119
rect 29271 2295 29305 2311
rect 29271 2103 29305 2119
rect 29385 2295 29419 2311
rect 29385 2103 29419 2119
rect 29643 2295 29677 2311
rect 29643 2103 29677 2119
rect 20875 2035 20891 2069
rect 21059 2035 21075 2069
rect 21247 2035 21263 2069
rect 21431 2035 21447 2069
rect 21619 2035 21635 2069
rect 21803 2035 21819 2069
rect 21991 2035 22007 2069
rect 22175 2035 22191 2069
rect 22363 2035 22379 2069
rect 22547 2035 22563 2069
rect 22735 2035 22751 2069
rect 22919 2035 22935 2069
rect 23107 2035 23123 2069
rect 23291 2035 23307 2069
rect 23479 2035 23495 2069
rect 23663 2035 23679 2069
rect 23851 2035 23867 2069
rect 24035 2035 24051 2069
rect 24223 2035 24239 2069
rect 24407 2035 24423 2069
rect 24595 2035 24611 2069
rect 24779 2035 24795 2069
rect 24967 2035 24983 2069
rect 25151 2035 25167 2069
rect 25339 2035 25355 2069
rect 25523 2035 25539 2069
rect 25711 2035 25727 2069
rect 25895 2035 25911 2069
rect 26083 2035 26099 2069
rect 26267 2035 26283 2069
rect 26455 2035 26471 2069
rect 26639 2035 26655 2069
rect 26827 2035 26843 2069
rect 27011 2035 27027 2069
rect 27199 2035 27215 2069
rect 27383 2035 27399 2069
rect 27571 2035 27587 2069
rect 27755 2035 27771 2069
rect 27943 2035 27959 2069
rect 28127 2035 28143 2069
rect 28315 2035 28331 2069
rect 28499 2035 28515 2069
rect 28687 2035 28703 2069
rect 28871 2035 28887 2069
rect 29059 2035 29075 2069
rect 29243 2035 29259 2069
rect 29431 2035 29447 2069
rect 29615 2035 29631 2069
rect 20715 1967 20749 2029
rect 29757 1967 29791 2029
rect 20715 1933 20811 1967
rect 29695 1933 29791 1967
<< viali >>
rect 19638 10817 19708 10834
rect 20382 10817 20452 10834
rect 21126 10817 21196 10834
rect 21870 10817 21940 10834
rect 22614 10817 22684 10834
rect 23358 10817 23428 10834
rect 24102 10817 24172 10834
rect 24846 10817 24916 10834
rect 25218 10817 25288 10834
rect 25962 10817 26032 10834
rect 26706 10817 26776 10834
rect 27450 10817 27520 10834
rect 28194 10817 28264 10834
rect 28938 10817 29008 10834
rect 29682 10817 29752 10834
rect 30426 10817 30496 10834
rect 31116 10817 31186 10834
rect 19638 10783 19708 10817
rect 20382 10783 20452 10817
rect 21126 10783 21196 10817
rect 21870 10783 21940 10817
rect 22614 10783 22684 10817
rect 23358 10783 23428 10817
rect 24102 10783 24172 10817
rect 24846 10783 24916 10817
rect 25218 10783 25288 10817
rect 25962 10783 26032 10817
rect 26706 10783 26776 10817
rect 27450 10783 27520 10817
rect 28194 10783 28264 10817
rect 28938 10783 29008 10817
rect 29682 10783 29752 10817
rect 30426 10783 30496 10817
rect 31116 10783 31183 10817
rect 31183 10783 31186 10817
rect 19638 10764 19708 10783
rect 20382 10764 20452 10783
rect 21126 10764 21196 10783
rect 21870 10764 21940 10783
rect 22614 10764 22684 10783
rect 23358 10764 23428 10783
rect 24102 10764 24172 10783
rect 24846 10764 24916 10783
rect 25218 10764 25288 10783
rect 25962 10764 26032 10783
rect 26706 10764 26776 10783
rect 27450 10764 27520 10783
rect 28194 10764 28264 10783
rect 28938 10764 29008 10783
rect 29682 10764 29752 10783
rect 30426 10764 30496 10783
rect 31116 10764 31186 10783
rect 19403 10681 19571 10715
rect 19775 10681 19943 10715
rect 20147 10681 20315 10715
rect 20519 10681 20687 10715
rect 20891 10681 21059 10715
rect 21263 10681 21431 10715
rect 21635 10681 21803 10715
rect 22007 10681 22175 10715
rect 22379 10681 22547 10715
rect 22751 10681 22919 10715
rect 23123 10681 23291 10715
rect 23495 10681 23663 10715
rect 23867 10681 24035 10715
rect 24239 10681 24407 10715
rect 24611 10681 24779 10715
rect 24983 10681 25151 10715
rect 25355 10681 25523 10715
rect 25727 10681 25895 10715
rect 26099 10681 26267 10715
rect 26471 10681 26639 10715
rect 26843 10681 27011 10715
rect 27215 10681 27383 10715
rect 27587 10681 27755 10715
rect 27959 10681 28127 10715
rect 28331 10681 28499 10715
rect 28703 10681 28871 10715
rect 29075 10681 29243 10715
rect 29447 10681 29615 10715
rect 29819 10681 29987 10715
rect 30191 10681 30359 10715
rect 30563 10681 30731 10715
rect 30935 10681 31103 10715
rect 19341 10246 19375 10622
rect 19599 10246 19633 10622
rect 19713 10246 19747 10622
rect 19971 10246 20005 10622
rect 20085 10246 20119 10622
rect 20343 10246 20377 10622
rect 20457 10246 20491 10622
rect 20715 10246 20749 10622
rect 20829 10246 20863 10622
rect 21087 10246 21121 10622
rect 21201 10246 21235 10622
rect 21459 10246 21493 10622
rect 21573 10246 21607 10622
rect 21831 10246 21865 10622
rect 21945 10246 21979 10622
rect 22203 10246 22237 10622
rect 22317 10246 22351 10622
rect 22575 10246 22609 10622
rect 22689 10246 22723 10622
rect 22947 10246 22981 10622
rect 23061 10246 23095 10622
rect 23319 10246 23353 10622
rect 23433 10246 23467 10622
rect 23691 10246 23725 10622
rect 23805 10246 23839 10622
rect 24063 10246 24097 10622
rect 24177 10246 24211 10622
rect 24435 10246 24469 10622
rect 24549 10246 24583 10622
rect 24807 10246 24841 10622
rect 24921 10246 24955 10622
rect 25179 10246 25213 10622
rect 25293 10246 25327 10622
rect 25551 10246 25585 10622
rect 25665 10246 25699 10622
rect 25923 10246 25957 10622
rect 26037 10246 26071 10622
rect 26295 10246 26329 10622
rect 26409 10246 26443 10622
rect 26667 10246 26701 10622
rect 26781 10246 26815 10622
rect 27039 10246 27073 10622
rect 27153 10246 27187 10622
rect 27411 10246 27445 10622
rect 27525 10246 27559 10622
rect 27783 10246 27817 10622
rect 27897 10246 27931 10622
rect 28155 10246 28189 10622
rect 28269 10246 28303 10622
rect 28527 10246 28561 10622
rect 28641 10246 28675 10622
rect 28899 10246 28933 10622
rect 29013 10246 29047 10622
rect 29271 10246 29305 10622
rect 29385 10246 29419 10622
rect 29643 10246 29677 10622
rect 29757 10246 29791 10622
rect 30015 10246 30049 10622
rect 30129 10246 30163 10622
rect 30387 10246 30421 10622
rect 30501 10246 30535 10622
rect 30759 10246 30793 10622
rect 30873 10246 30907 10622
rect 31131 10246 31165 10622
rect 19403 10153 19571 10187
rect 19775 10153 19943 10187
rect 20147 10153 20315 10187
rect 20519 10153 20687 10187
rect 20891 10153 21059 10187
rect 21263 10153 21431 10187
rect 21635 10153 21803 10187
rect 22007 10153 22175 10187
rect 22379 10153 22547 10187
rect 22751 10153 22919 10187
rect 23123 10153 23291 10187
rect 23495 10153 23663 10187
rect 23867 10153 24035 10187
rect 24239 10153 24407 10187
rect 24611 10153 24779 10187
rect 24983 10153 25151 10187
rect 25355 10153 25523 10187
rect 25727 10153 25895 10187
rect 26099 10153 26267 10187
rect 26471 10153 26639 10187
rect 26843 10153 27011 10187
rect 27215 10153 27383 10187
rect 27587 10153 27755 10187
rect 27959 10153 28127 10187
rect 28331 10153 28499 10187
rect 28703 10153 28871 10187
rect 29075 10153 29243 10187
rect 29447 10153 29615 10187
rect 29819 10153 29987 10187
rect 30191 10153 30359 10187
rect 30563 10153 30731 10187
rect 30935 10153 31103 10187
rect 19403 10045 19571 10079
rect 19775 10045 19943 10079
rect 20147 10045 20315 10079
rect 20519 10045 20687 10079
rect 20891 10045 21059 10079
rect 21263 10045 21431 10079
rect 21635 10045 21803 10079
rect 22007 10045 22175 10079
rect 22379 10045 22547 10079
rect 22751 10045 22919 10079
rect 23123 10045 23291 10079
rect 23495 10045 23663 10079
rect 23867 10045 24035 10079
rect 24239 10045 24407 10079
rect 24611 10045 24779 10079
rect 24983 10045 25151 10079
rect 25355 10045 25523 10079
rect 25727 10045 25895 10079
rect 26099 10045 26267 10079
rect 26471 10045 26639 10079
rect 26843 10045 27011 10079
rect 27215 10045 27383 10079
rect 27587 10045 27755 10079
rect 27959 10045 28127 10079
rect 28331 10045 28499 10079
rect 28703 10045 28871 10079
rect 29075 10045 29243 10079
rect 29447 10045 29615 10079
rect 29819 10045 29987 10079
rect 30191 10045 30359 10079
rect 30563 10045 30731 10079
rect 30935 10045 31103 10079
rect 19341 9610 19375 9986
rect 19599 9610 19633 9986
rect 19713 9610 19747 9986
rect 19971 9610 20005 9986
rect 20085 9610 20119 9986
rect 20343 9610 20377 9986
rect 20457 9610 20491 9986
rect 20715 9610 20749 9986
rect 20829 9610 20863 9986
rect 21087 9610 21121 9986
rect 21201 9610 21235 9986
rect 21459 9610 21493 9986
rect 21573 9610 21607 9986
rect 21831 9610 21865 9986
rect 21945 9610 21979 9986
rect 22203 9610 22237 9986
rect 22317 9610 22351 9986
rect 22575 9610 22609 9986
rect 22689 9610 22723 9986
rect 22947 9610 22981 9986
rect 23061 9610 23095 9986
rect 23319 9610 23353 9986
rect 23433 9610 23467 9986
rect 23691 9610 23725 9986
rect 23805 9610 23839 9986
rect 24063 9610 24097 9986
rect 24177 9610 24211 9986
rect 24435 9610 24469 9986
rect 24549 9610 24583 9986
rect 24807 9610 24841 9986
rect 24921 9610 24955 9986
rect 25179 9610 25213 9986
rect 25293 9610 25327 9986
rect 25551 9610 25585 9986
rect 25665 9610 25699 9986
rect 25923 9610 25957 9986
rect 26037 9610 26071 9986
rect 26295 9610 26329 9986
rect 26409 9610 26443 9986
rect 26667 9610 26701 9986
rect 26781 9610 26815 9986
rect 27039 9610 27073 9986
rect 27153 9610 27187 9986
rect 27411 9610 27445 9986
rect 27525 9610 27559 9986
rect 27783 9610 27817 9986
rect 27897 9610 27931 9986
rect 28155 9610 28189 9986
rect 28269 9610 28303 9986
rect 28527 9610 28561 9986
rect 28641 9610 28675 9986
rect 28899 9610 28933 9986
rect 29013 9610 29047 9986
rect 29271 9610 29305 9986
rect 29385 9610 29419 9986
rect 29643 9610 29677 9986
rect 29757 9610 29791 9986
rect 30015 9610 30049 9986
rect 30129 9610 30163 9986
rect 30387 9610 30421 9986
rect 30501 9610 30535 9986
rect 30759 9610 30793 9986
rect 30873 9610 30907 9986
rect 31131 9610 31165 9986
rect 19403 9517 19571 9551
rect 19775 9517 19943 9551
rect 20147 9517 20315 9551
rect 20519 9517 20687 9551
rect 20891 9517 21059 9551
rect 21263 9517 21431 9551
rect 21635 9517 21803 9551
rect 22007 9517 22175 9551
rect 22379 9517 22547 9551
rect 22751 9517 22919 9551
rect 23123 9517 23291 9551
rect 23495 9517 23663 9551
rect 23867 9517 24035 9551
rect 24239 9517 24407 9551
rect 24611 9517 24779 9551
rect 24983 9517 25151 9551
rect 25355 9517 25523 9551
rect 25727 9517 25895 9551
rect 26099 9517 26267 9551
rect 26471 9517 26639 9551
rect 26843 9517 27011 9551
rect 27215 9517 27383 9551
rect 27587 9517 27755 9551
rect 27959 9517 28127 9551
rect 28331 9517 28499 9551
rect 28703 9517 28871 9551
rect 29075 9517 29243 9551
rect 29447 9517 29615 9551
rect 29819 9517 29987 9551
rect 30191 9517 30359 9551
rect 30563 9517 30731 9551
rect 30935 9517 31103 9551
rect 19403 9409 19571 9443
rect 19775 9409 19943 9443
rect 20147 9409 20315 9443
rect 20519 9409 20687 9443
rect 20891 9409 21059 9443
rect 21263 9409 21431 9443
rect 21635 9409 21803 9443
rect 22007 9409 22175 9443
rect 22379 9409 22547 9443
rect 22751 9409 22919 9443
rect 23123 9409 23291 9443
rect 23495 9409 23663 9443
rect 23867 9409 24035 9443
rect 24239 9409 24407 9443
rect 24611 9409 24779 9443
rect 24983 9409 25151 9443
rect 25355 9409 25523 9443
rect 25727 9409 25895 9443
rect 26099 9409 26267 9443
rect 26471 9409 26639 9443
rect 26843 9409 27011 9443
rect 27215 9409 27383 9443
rect 27587 9409 27755 9443
rect 27959 9409 28127 9443
rect 28331 9409 28499 9443
rect 28703 9409 28871 9443
rect 29075 9409 29243 9443
rect 29447 9409 29615 9443
rect 29819 9409 29987 9443
rect 30191 9409 30359 9443
rect 30563 9409 30731 9443
rect 30935 9409 31103 9443
rect 19341 8974 19375 9350
rect 19599 8974 19633 9350
rect 19713 8974 19747 9350
rect 19971 8974 20005 9350
rect 20085 8974 20119 9350
rect 20343 8974 20377 9350
rect 20457 8974 20491 9350
rect 20715 8974 20749 9350
rect 20829 8974 20863 9350
rect 21087 8974 21121 9350
rect 21201 8974 21235 9350
rect 21459 8974 21493 9350
rect 21573 8974 21607 9350
rect 21831 8974 21865 9350
rect 21945 8974 21979 9350
rect 22203 8974 22237 9350
rect 22317 8974 22351 9350
rect 22575 8974 22609 9350
rect 22689 8974 22723 9350
rect 22947 8974 22981 9350
rect 23061 8974 23095 9350
rect 23319 8974 23353 9350
rect 23433 8974 23467 9350
rect 23691 8974 23725 9350
rect 23805 8974 23839 9350
rect 24063 8974 24097 9350
rect 24177 8974 24211 9350
rect 24435 8974 24469 9350
rect 24549 8974 24583 9350
rect 24807 8974 24841 9350
rect 24921 8974 24955 9350
rect 25179 8974 25213 9350
rect 25293 8974 25327 9350
rect 25551 8974 25585 9350
rect 25665 8974 25699 9350
rect 25923 8974 25957 9350
rect 26037 8974 26071 9350
rect 26295 8974 26329 9350
rect 26409 8974 26443 9350
rect 26667 8974 26701 9350
rect 26781 8974 26815 9350
rect 27039 8974 27073 9350
rect 27153 8974 27187 9350
rect 27411 8974 27445 9350
rect 27525 8974 27559 9350
rect 27783 8974 27817 9350
rect 27897 8974 27931 9350
rect 28155 8974 28189 9350
rect 28269 8974 28303 9350
rect 28527 8974 28561 9350
rect 28641 8974 28675 9350
rect 28899 8974 28933 9350
rect 29013 8974 29047 9350
rect 29271 8974 29305 9350
rect 29385 8974 29419 9350
rect 29643 8974 29677 9350
rect 29757 8974 29791 9350
rect 30015 8974 30049 9350
rect 30129 8974 30163 9350
rect 30387 8974 30421 9350
rect 30501 8974 30535 9350
rect 30759 8974 30793 9350
rect 30873 8974 30907 9350
rect 31131 8974 31165 9350
rect 19403 8881 19571 8915
rect 19775 8881 19943 8915
rect 20147 8881 20315 8915
rect 20519 8881 20687 8915
rect 20891 8881 21059 8915
rect 21263 8881 21431 8915
rect 21635 8881 21803 8915
rect 22007 8881 22175 8915
rect 22379 8881 22547 8915
rect 22751 8881 22919 8915
rect 23123 8881 23291 8915
rect 23495 8881 23663 8915
rect 23867 8881 24035 8915
rect 24239 8881 24407 8915
rect 24611 8881 24779 8915
rect 24983 8881 25151 8915
rect 25355 8881 25523 8915
rect 25727 8881 25895 8915
rect 26099 8881 26267 8915
rect 26471 8881 26639 8915
rect 26843 8881 27011 8915
rect 27215 8881 27383 8915
rect 27587 8881 27755 8915
rect 27959 8881 28127 8915
rect 28331 8881 28499 8915
rect 28703 8881 28871 8915
rect 29075 8881 29243 8915
rect 29447 8881 29615 8915
rect 29819 8881 29987 8915
rect 30191 8881 30359 8915
rect 30563 8881 30731 8915
rect 30935 8881 31103 8915
rect 20800 8429 20870 8446
rect 21172 8429 21242 8446
rect 21544 8429 21614 8446
rect 21916 8429 21986 8446
rect 22288 8429 22358 8446
rect 22660 8429 22730 8446
rect 23032 8429 23102 8446
rect 23404 8429 23474 8446
rect 23666 8429 23736 8446
rect 20800 8395 20811 8429
rect 20811 8395 20870 8429
rect 21172 8395 21242 8429
rect 21544 8395 21614 8429
rect 21916 8395 21986 8429
rect 22288 8395 22358 8429
rect 22660 8395 22730 8429
rect 23032 8395 23102 8429
rect 23404 8395 23474 8429
rect 23666 8395 23736 8429
rect 20800 8376 20870 8395
rect 21172 8376 21242 8395
rect 21544 8376 21614 8395
rect 21916 8376 21986 8395
rect 22288 8376 22358 8395
rect 22660 8376 22730 8395
rect 23032 8376 23102 8395
rect 23404 8376 23474 8395
rect 23666 8376 23736 8395
rect 20891 8293 21059 8327
rect 21263 8293 21431 8327
rect 21635 8293 21803 8327
rect 22007 8293 22175 8327
rect 22379 8293 22547 8327
rect 22751 8293 22919 8327
rect 23123 8293 23291 8327
rect 23495 8293 23663 8327
rect 20829 7458 20863 8234
rect 21087 7458 21121 8234
rect 21201 7458 21235 8234
rect 21459 7458 21493 8234
rect 21573 7458 21607 8234
rect 21831 7458 21865 8234
rect 21945 7458 21979 8234
rect 22203 7458 22237 8234
rect 22317 7458 22351 8234
rect 22575 7458 22609 8234
rect 22689 7458 22723 8234
rect 22947 7458 22981 8234
rect 23061 7458 23095 8234
rect 23319 7458 23353 8234
rect 23433 7458 23467 8234
rect 23691 7458 23725 8234
rect 20891 7365 21059 7399
rect 21263 7365 21431 7399
rect 21635 7365 21803 7399
rect 22007 7365 22175 7399
rect 22379 7365 22547 7399
rect 22751 7365 22919 7399
rect 23123 7365 23291 7399
rect 23495 7365 23663 7399
rect 20891 7257 21059 7291
rect 21263 7257 21431 7291
rect 21635 7257 21803 7291
rect 22007 7257 22175 7291
rect 22379 7257 22547 7291
rect 22751 7257 22919 7291
rect 23123 7257 23291 7291
rect 23495 7257 23663 7291
rect 20829 6422 20863 7198
rect 21087 6422 21121 7198
rect 21201 6422 21235 7198
rect 21459 6422 21493 7198
rect 21573 6422 21607 7198
rect 21831 6422 21865 7198
rect 21945 6422 21979 7198
rect 22203 6422 22237 7198
rect 22317 6422 22351 7198
rect 22575 6422 22609 7198
rect 22689 6422 22723 7198
rect 22947 6422 22981 7198
rect 23061 6422 23095 7198
rect 23319 6422 23353 7198
rect 23433 6422 23467 7198
rect 23691 6422 23725 7198
rect 20891 6329 21059 6363
rect 21263 6329 21431 6363
rect 21635 6329 21803 6363
rect 22007 6329 22175 6363
rect 22379 6329 22547 6363
rect 22751 6329 22919 6363
rect 23123 6329 23291 6363
rect 23495 6329 23663 6363
rect 20891 6221 21059 6255
rect 21263 6221 21431 6255
rect 21635 6221 21803 6255
rect 22007 6221 22175 6255
rect 22379 6221 22547 6255
rect 22751 6221 22919 6255
rect 23123 6221 23291 6255
rect 23495 6221 23663 6255
rect 20829 5386 20863 6162
rect 21087 5386 21121 6162
rect 21201 5386 21235 6162
rect 21459 5386 21493 6162
rect 21573 5386 21607 6162
rect 21831 5386 21865 6162
rect 21945 5386 21979 6162
rect 22203 5386 22237 6162
rect 22317 5386 22351 6162
rect 22575 5386 22609 6162
rect 22689 5386 22723 6162
rect 22947 5386 22981 6162
rect 23061 5386 23095 6162
rect 23319 5386 23353 6162
rect 23433 5386 23467 6162
rect 23691 5386 23725 6162
rect 20891 5293 21059 5327
rect 21263 5293 21431 5327
rect 21635 5293 21803 5327
rect 22007 5293 22175 5327
rect 22379 5293 22547 5327
rect 22751 5293 22919 5327
rect 23123 5293 23291 5327
rect 23495 5293 23663 5327
rect 20891 5185 21059 5219
rect 21263 5185 21431 5219
rect 21635 5185 21803 5219
rect 22007 5185 22175 5219
rect 22379 5185 22547 5219
rect 22751 5185 22919 5219
rect 23123 5185 23291 5219
rect 23495 5185 23663 5219
rect 20829 4350 20863 5126
rect 21087 4350 21121 5126
rect 21201 4350 21235 5126
rect 21459 4350 21493 5126
rect 21573 4350 21607 5126
rect 21831 4350 21865 5126
rect 21945 4350 21979 5126
rect 22203 4350 22237 5126
rect 22317 4350 22351 5126
rect 22575 4350 22609 5126
rect 22689 4350 22723 5126
rect 22947 4350 22981 5126
rect 23061 4350 23095 5126
rect 23319 4350 23353 5126
rect 23433 4350 23467 5126
rect 23691 4350 23725 5126
rect 20891 4257 21059 4291
rect 21263 4257 21431 4291
rect 21635 4257 21803 4291
rect 22007 4257 22175 4291
rect 22379 4257 22547 4291
rect 22751 4257 22919 4291
rect 23123 4257 23291 4291
rect 23495 4257 23663 4291
rect 20891 3599 21059 3633
rect 21263 3599 21431 3633
rect 21635 3599 21803 3633
rect 22007 3599 22175 3633
rect 22379 3599 22547 3633
rect 22751 3599 22919 3633
rect 23123 3599 23291 3633
rect 23495 3599 23663 3633
rect 23867 3599 24035 3633
rect 24239 3599 24407 3633
rect 24611 3599 24779 3633
rect 24983 3599 25151 3633
rect 25355 3599 25523 3633
rect 25727 3599 25895 3633
rect 26099 3599 26267 3633
rect 26471 3599 26639 3633
rect 26843 3599 27011 3633
rect 27215 3599 27383 3633
rect 27587 3599 27755 3633
rect 27959 3599 28127 3633
rect 28331 3599 28499 3633
rect 28703 3599 28871 3633
rect 29075 3599 29243 3633
rect 29447 3599 29615 3633
rect 20829 3373 20863 3549
rect 21087 3373 21121 3549
rect 21201 3373 21235 3549
rect 21459 3373 21493 3549
rect 21573 3373 21607 3549
rect 21831 3373 21865 3549
rect 21945 3373 21979 3549
rect 22203 3373 22237 3549
rect 22317 3373 22351 3549
rect 22575 3373 22609 3549
rect 22689 3373 22723 3549
rect 22947 3373 22981 3549
rect 23061 3373 23095 3549
rect 23319 3373 23353 3549
rect 23433 3373 23467 3549
rect 23691 3373 23725 3549
rect 23805 3373 23839 3549
rect 24063 3373 24097 3549
rect 24177 3373 24211 3549
rect 24435 3373 24469 3549
rect 24549 3373 24583 3549
rect 24807 3373 24841 3549
rect 24921 3373 24955 3549
rect 25179 3373 25213 3549
rect 25293 3373 25327 3549
rect 25551 3373 25585 3549
rect 25665 3373 25699 3549
rect 25923 3373 25957 3549
rect 26037 3373 26071 3549
rect 26295 3373 26329 3549
rect 26409 3373 26443 3549
rect 26667 3373 26701 3549
rect 26781 3373 26815 3549
rect 27039 3373 27073 3549
rect 27153 3373 27187 3549
rect 27411 3373 27445 3549
rect 27525 3373 27559 3549
rect 27783 3373 27817 3549
rect 27897 3373 27931 3549
rect 28155 3373 28189 3549
rect 28269 3373 28303 3549
rect 28527 3373 28561 3549
rect 28641 3373 28675 3549
rect 28899 3373 28933 3549
rect 29013 3373 29047 3549
rect 29271 3373 29305 3549
rect 29385 3373 29419 3549
rect 29643 3373 29677 3549
rect 20891 3289 21059 3323
rect 21263 3289 21431 3323
rect 21635 3289 21803 3323
rect 22007 3289 22175 3323
rect 22379 3289 22547 3323
rect 22751 3289 22919 3323
rect 23123 3289 23291 3323
rect 23495 3289 23663 3323
rect 23867 3289 24035 3323
rect 24239 3289 24407 3323
rect 24611 3289 24779 3323
rect 24983 3289 25151 3323
rect 25355 3289 25523 3323
rect 25727 3289 25895 3323
rect 26099 3289 26267 3323
rect 26471 3289 26639 3323
rect 26843 3289 27011 3323
rect 27215 3289 27383 3323
rect 27587 3289 27755 3323
rect 27959 3289 28127 3323
rect 28331 3289 28499 3323
rect 28703 3289 28871 3323
rect 29075 3289 29243 3323
rect 29447 3289 29615 3323
rect 20891 3181 21059 3215
rect 21263 3181 21431 3215
rect 21635 3181 21803 3215
rect 22007 3181 22175 3215
rect 22379 3181 22547 3215
rect 22751 3181 22919 3215
rect 23123 3181 23291 3215
rect 23495 3181 23663 3215
rect 23867 3181 24035 3215
rect 24239 3181 24407 3215
rect 24611 3181 24779 3215
rect 24983 3181 25151 3215
rect 25355 3181 25523 3215
rect 25727 3181 25895 3215
rect 26099 3181 26267 3215
rect 26471 3181 26639 3215
rect 26843 3181 27011 3215
rect 27215 3181 27383 3215
rect 27587 3181 27755 3215
rect 27959 3181 28127 3215
rect 28331 3181 28499 3215
rect 28703 3181 28871 3215
rect 29075 3181 29243 3215
rect 29447 3181 29615 3215
rect 20829 2955 20863 3131
rect 21087 2955 21121 3131
rect 21201 2955 21235 3131
rect 21459 2955 21493 3131
rect 21573 2955 21607 3131
rect 21831 2955 21865 3131
rect 21945 2955 21979 3131
rect 22203 2955 22237 3131
rect 22317 2955 22351 3131
rect 22575 2955 22609 3131
rect 22689 2955 22723 3131
rect 22947 2955 22981 3131
rect 23061 2955 23095 3131
rect 23319 2955 23353 3131
rect 23433 2955 23467 3131
rect 23691 2955 23725 3131
rect 23805 2955 23839 3131
rect 24063 2955 24097 3131
rect 24177 2955 24211 3131
rect 24435 2955 24469 3131
rect 24549 2955 24583 3131
rect 24807 2955 24841 3131
rect 24921 2955 24955 3131
rect 25179 2955 25213 3131
rect 25293 2955 25327 3131
rect 25551 2955 25585 3131
rect 25665 2955 25699 3131
rect 25923 2955 25957 3131
rect 26037 2955 26071 3131
rect 26295 2955 26329 3131
rect 26409 2955 26443 3131
rect 26667 2955 26701 3131
rect 26781 2955 26815 3131
rect 27039 2955 27073 3131
rect 27153 2955 27187 3131
rect 27411 2955 27445 3131
rect 27525 2955 27559 3131
rect 27783 2955 27817 3131
rect 27897 2955 27931 3131
rect 28155 2955 28189 3131
rect 28269 2955 28303 3131
rect 28527 2955 28561 3131
rect 28641 2955 28675 3131
rect 28899 2955 28933 3131
rect 29013 2955 29047 3131
rect 29271 2955 29305 3131
rect 29385 2955 29419 3131
rect 29643 2955 29677 3131
rect 20891 2871 21059 2905
rect 21263 2871 21431 2905
rect 21635 2871 21803 2905
rect 22007 2871 22175 2905
rect 22379 2871 22547 2905
rect 22751 2871 22919 2905
rect 23123 2871 23291 2905
rect 23495 2871 23663 2905
rect 23867 2871 24035 2905
rect 24239 2871 24407 2905
rect 24611 2871 24779 2905
rect 24983 2871 25151 2905
rect 25355 2871 25523 2905
rect 25727 2871 25895 2905
rect 26099 2871 26267 2905
rect 26471 2871 26639 2905
rect 26843 2871 27011 2905
rect 27215 2871 27383 2905
rect 27587 2871 27755 2905
rect 27959 2871 28127 2905
rect 28331 2871 28499 2905
rect 28703 2871 28871 2905
rect 29075 2871 29243 2905
rect 29447 2871 29615 2905
rect 20891 2763 21059 2797
rect 21263 2763 21431 2797
rect 21635 2763 21803 2797
rect 22007 2763 22175 2797
rect 22379 2763 22547 2797
rect 22751 2763 22919 2797
rect 23123 2763 23291 2797
rect 23495 2763 23663 2797
rect 23867 2763 24035 2797
rect 24239 2763 24407 2797
rect 24611 2763 24779 2797
rect 24983 2763 25151 2797
rect 25355 2763 25523 2797
rect 25727 2763 25895 2797
rect 26099 2763 26267 2797
rect 26471 2763 26639 2797
rect 26843 2763 27011 2797
rect 27215 2763 27383 2797
rect 27587 2763 27755 2797
rect 27959 2763 28127 2797
rect 28331 2763 28499 2797
rect 28703 2763 28871 2797
rect 29075 2763 29243 2797
rect 29447 2763 29615 2797
rect 20829 2537 20863 2713
rect 21087 2537 21121 2713
rect 21201 2537 21235 2713
rect 21459 2537 21493 2713
rect 21573 2537 21607 2713
rect 21831 2537 21865 2713
rect 21945 2537 21979 2713
rect 22203 2537 22237 2713
rect 22317 2537 22351 2713
rect 22575 2537 22609 2713
rect 22689 2537 22723 2713
rect 22947 2537 22981 2713
rect 23061 2537 23095 2713
rect 23319 2537 23353 2713
rect 23433 2537 23467 2713
rect 23691 2537 23725 2713
rect 23805 2537 23839 2713
rect 24063 2537 24097 2713
rect 24177 2537 24211 2713
rect 24435 2537 24469 2713
rect 24549 2537 24583 2713
rect 24807 2537 24841 2713
rect 24921 2537 24955 2713
rect 25179 2537 25213 2713
rect 25293 2537 25327 2713
rect 25551 2537 25585 2713
rect 25665 2537 25699 2713
rect 25923 2537 25957 2713
rect 26037 2537 26071 2713
rect 26295 2537 26329 2713
rect 26409 2537 26443 2713
rect 26667 2537 26701 2713
rect 26781 2537 26815 2713
rect 27039 2537 27073 2713
rect 27153 2537 27187 2713
rect 27411 2537 27445 2713
rect 27525 2537 27559 2713
rect 27783 2537 27817 2713
rect 27897 2537 27931 2713
rect 28155 2537 28189 2713
rect 28269 2537 28303 2713
rect 28527 2537 28561 2713
rect 28641 2537 28675 2713
rect 28899 2537 28933 2713
rect 29013 2537 29047 2713
rect 29271 2537 29305 2713
rect 29385 2537 29419 2713
rect 29643 2537 29677 2713
rect 20891 2453 21059 2487
rect 21263 2453 21431 2487
rect 21635 2453 21803 2487
rect 22007 2453 22175 2487
rect 22379 2453 22547 2487
rect 22751 2453 22919 2487
rect 23123 2453 23291 2487
rect 23495 2453 23663 2487
rect 23867 2453 24035 2487
rect 24239 2453 24407 2487
rect 24611 2453 24779 2487
rect 24983 2453 25151 2487
rect 25355 2453 25523 2487
rect 25727 2453 25895 2487
rect 26099 2453 26267 2487
rect 26471 2453 26639 2487
rect 26843 2453 27011 2487
rect 27215 2453 27383 2487
rect 27587 2453 27755 2487
rect 27959 2453 28127 2487
rect 28331 2453 28499 2487
rect 28703 2453 28871 2487
rect 29075 2453 29243 2487
rect 29447 2453 29615 2487
rect 20891 2345 21059 2379
rect 21263 2345 21431 2379
rect 21635 2345 21803 2379
rect 22007 2345 22175 2379
rect 22379 2345 22547 2379
rect 22751 2345 22919 2379
rect 23123 2345 23291 2379
rect 23495 2345 23663 2379
rect 23867 2345 24035 2379
rect 24239 2345 24407 2379
rect 24611 2345 24779 2379
rect 24983 2345 25151 2379
rect 25355 2345 25523 2379
rect 25727 2345 25895 2379
rect 26099 2345 26267 2379
rect 26471 2345 26639 2379
rect 26843 2345 27011 2379
rect 27215 2345 27383 2379
rect 27587 2345 27755 2379
rect 27959 2345 28127 2379
rect 28331 2345 28499 2379
rect 28703 2345 28871 2379
rect 29075 2345 29243 2379
rect 29447 2345 29615 2379
rect 20829 2119 20863 2295
rect 21087 2119 21121 2295
rect 21201 2119 21235 2295
rect 21459 2119 21493 2295
rect 21573 2119 21607 2295
rect 21831 2119 21865 2295
rect 21945 2119 21979 2295
rect 22203 2119 22237 2295
rect 22317 2119 22351 2295
rect 22575 2119 22609 2295
rect 22689 2119 22723 2295
rect 22947 2119 22981 2295
rect 23061 2119 23095 2295
rect 23319 2119 23353 2295
rect 23433 2119 23467 2295
rect 23691 2119 23725 2295
rect 23805 2119 23839 2295
rect 24063 2119 24097 2295
rect 24177 2119 24211 2295
rect 24435 2119 24469 2295
rect 24549 2119 24583 2295
rect 24807 2119 24841 2295
rect 24921 2119 24955 2295
rect 25179 2119 25213 2295
rect 25293 2119 25327 2295
rect 25551 2119 25585 2295
rect 25665 2119 25699 2295
rect 25923 2119 25957 2295
rect 26037 2119 26071 2295
rect 26295 2119 26329 2295
rect 26409 2119 26443 2295
rect 26667 2119 26701 2295
rect 26781 2119 26815 2295
rect 27039 2119 27073 2295
rect 27153 2119 27187 2295
rect 27411 2119 27445 2295
rect 27525 2119 27559 2295
rect 27783 2119 27817 2295
rect 27897 2119 27931 2295
rect 28155 2119 28189 2295
rect 28269 2119 28303 2295
rect 28527 2119 28561 2295
rect 28641 2119 28675 2295
rect 28899 2119 28933 2295
rect 29013 2119 29047 2295
rect 29271 2119 29305 2295
rect 29385 2119 29419 2295
rect 29643 2119 29677 2295
rect 20891 2035 21059 2069
rect 21263 2035 21431 2069
rect 21635 2035 21803 2069
rect 22007 2035 22175 2069
rect 22379 2035 22547 2069
rect 22751 2035 22919 2069
rect 23123 2035 23291 2069
rect 23495 2035 23663 2069
rect 23867 2035 24035 2069
rect 24239 2035 24407 2069
rect 24611 2035 24779 2069
rect 24983 2035 25151 2069
rect 25355 2035 25523 2069
rect 25727 2035 25895 2069
rect 26099 2035 26267 2069
rect 26471 2035 26639 2069
rect 26843 2035 27011 2069
rect 27215 2035 27383 2069
rect 27587 2035 27755 2069
rect 27959 2035 28127 2069
rect 28331 2035 28499 2069
rect 28703 2035 28871 2069
rect 29075 2035 29243 2069
rect 29447 2035 29615 2069
rect 20830 1967 20900 1978
rect 21498 1967 21568 1986
rect 22242 1967 22312 1986
rect 22986 1967 23056 1986
rect 23730 1967 23800 1986
rect 24474 1967 24544 1986
rect 25218 1967 25288 1986
rect 25962 1967 26032 1986
rect 26706 1967 26776 1986
rect 27450 1967 27520 1986
rect 28194 1967 28264 1986
rect 28938 1967 29008 1986
rect 29600 1967 29670 1982
rect 20830 1933 20900 1967
rect 21498 1933 21568 1967
rect 22242 1933 22312 1967
rect 22986 1933 23056 1967
rect 23730 1933 23800 1967
rect 24474 1933 24544 1967
rect 25218 1933 25288 1967
rect 25962 1933 26032 1967
rect 26706 1933 26776 1967
rect 27450 1933 27520 1967
rect 28194 1933 28264 1967
rect 28938 1933 29008 1967
rect 29600 1933 29670 1967
rect 20830 1908 20900 1933
rect 21498 1916 21568 1933
rect 22242 1916 22312 1933
rect 22986 1916 23056 1933
rect 23730 1916 23800 1933
rect 24474 1916 24544 1933
rect 25218 1916 25288 1933
rect 25962 1916 26032 1933
rect 26706 1916 26776 1933
rect 27450 1916 27520 1933
rect 28194 1916 28264 1933
rect 28938 1916 29008 1933
rect 29600 1912 29670 1933
<< metal1 >>
rect 19562 10916 19572 11116
rect 19772 10916 19782 11116
rect 20306 10916 20316 11116
rect 20516 10916 20526 11116
rect 21050 10916 21060 11116
rect 21260 10916 21270 11116
rect 21794 10916 21804 11116
rect 22004 10916 22014 11116
rect 22538 10916 22548 11116
rect 22748 10916 22758 11116
rect 23282 10916 23292 11116
rect 23492 10916 23502 11116
rect 24026 10916 24036 11116
rect 24236 10916 24246 11116
rect 24770 10916 24780 11116
rect 24980 10916 24990 11116
rect 25142 10916 25152 11116
rect 25352 10916 25362 11116
rect 25886 10916 25896 11116
rect 26096 10916 26106 11116
rect 26630 10916 26640 11116
rect 26840 10916 26850 11116
rect 27374 10916 27384 11116
rect 27584 10916 27594 11116
rect 28118 10916 28128 11116
rect 28328 10916 28338 11116
rect 28862 10916 28872 11116
rect 29072 10916 29082 11116
rect 29606 10916 29616 11116
rect 29816 10916 29826 11116
rect 30350 10916 30360 11116
rect 30560 10916 30570 11116
rect 31094 10916 31104 11116
rect 31304 10916 31314 11116
rect 19644 10840 19702 10916
rect 20388 10840 20446 10916
rect 21132 10840 21190 10916
rect 21876 10840 21934 10916
rect 22620 10840 22678 10916
rect 23364 10840 23422 10916
rect 24108 10840 24166 10916
rect 24832 10906 24910 10916
rect 24852 10840 24910 10906
rect 25262 10840 25314 10916
rect 25968 10840 26026 10916
rect 26712 10840 26770 10916
rect 27456 10840 27514 10916
rect 28200 10840 28258 10916
rect 28944 10840 29002 10916
rect 29688 10840 29746 10916
rect 30432 10840 30490 10916
rect 31158 10900 31234 10916
rect 31158 10840 31216 10900
rect 19626 10834 19720 10840
rect 19626 10764 19638 10834
rect 19708 10764 19720 10834
rect 19626 10758 19720 10764
rect 20370 10834 20464 10840
rect 20370 10764 20382 10834
rect 20452 10764 20464 10834
rect 20370 10758 20464 10764
rect 21114 10834 21208 10840
rect 21114 10764 21126 10834
rect 21196 10764 21208 10834
rect 21114 10758 21208 10764
rect 21858 10834 21952 10840
rect 21858 10764 21870 10834
rect 21940 10764 21952 10834
rect 21858 10758 21952 10764
rect 22602 10834 22696 10840
rect 22602 10764 22614 10834
rect 22684 10764 22696 10834
rect 22602 10758 22696 10764
rect 23346 10834 23440 10840
rect 23346 10764 23358 10834
rect 23428 10764 23440 10834
rect 23346 10758 23440 10764
rect 24090 10834 24184 10840
rect 24090 10764 24102 10834
rect 24172 10764 24184 10834
rect 24090 10758 24184 10764
rect 24834 10834 24928 10840
rect 24834 10764 24846 10834
rect 24916 10764 24928 10834
rect 24834 10758 24928 10764
rect 25206 10834 25314 10840
rect 25206 10764 25218 10834
rect 25288 10764 25314 10834
rect 25206 10758 25314 10764
rect 25950 10834 26044 10840
rect 25950 10764 25962 10834
rect 26032 10764 26044 10834
rect 25950 10758 26044 10764
rect 26694 10834 26788 10840
rect 26694 10764 26706 10834
rect 26776 10764 26788 10834
rect 26694 10758 26788 10764
rect 27438 10834 27532 10840
rect 27438 10764 27450 10834
rect 27520 10764 27532 10834
rect 27438 10758 27532 10764
rect 28182 10834 28276 10840
rect 28182 10764 28194 10834
rect 28264 10764 28276 10834
rect 28182 10758 28276 10764
rect 28926 10834 29020 10840
rect 28926 10764 28938 10834
rect 29008 10764 29020 10834
rect 28926 10758 29020 10764
rect 29670 10834 29764 10840
rect 29670 10764 29682 10834
rect 29752 10764 29764 10834
rect 29670 10758 29764 10764
rect 30414 10834 30508 10840
rect 30414 10764 30426 10834
rect 30496 10764 30508 10834
rect 30414 10758 30508 10764
rect 31104 10834 31216 10840
rect 31104 10764 31116 10834
rect 31186 10764 31216 10834
rect 31104 10758 31216 10764
rect 19334 10668 19402 10728
rect 19572 10721 19582 10728
rect 19572 10675 19583 10721
rect 19572 10668 19582 10675
rect 19334 10622 19382 10668
rect 19644 10634 19702 10758
rect 19764 10721 19774 10728
rect 19763 10675 19774 10721
rect 19944 10721 19954 10728
rect 20136 10721 20146 10728
rect 19764 10668 19774 10675
rect 19944 10675 19955 10721
rect 20135 10675 20146 10721
rect 20316 10721 20326 10728
rect 19944 10668 19954 10675
rect 20136 10668 20146 10675
rect 20316 10675 20327 10721
rect 20316 10668 20326 10675
rect 20388 10634 20446 10758
rect 20508 10721 20518 10728
rect 20507 10675 20518 10721
rect 20508 10668 20518 10675
rect 20688 10668 20890 10728
rect 21060 10721 21070 10728
rect 21060 10675 21071 10721
rect 21060 10668 21070 10675
rect 20760 10634 20818 10668
rect 21132 10634 21190 10758
rect 21252 10721 21262 10728
rect 21251 10675 21262 10721
rect 21432 10721 21442 10728
rect 21624 10721 21634 10728
rect 21252 10668 21262 10675
rect 21432 10675 21443 10721
rect 21623 10675 21634 10721
rect 21804 10721 21814 10728
rect 21432 10668 21442 10675
rect 21624 10668 21634 10675
rect 21804 10675 21815 10721
rect 21804 10668 21814 10675
rect 21876 10634 21934 10758
rect 21996 10721 22006 10728
rect 21995 10675 22006 10721
rect 21996 10668 22006 10675
rect 22176 10668 22378 10728
rect 22548 10721 22558 10728
rect 22548 10675 22559 10721
rect 22548 10668 22558 10675
rect 22248 10634 22306 10668
rect 22620 10634 22678 10758
rect 22740 10721 22750 10728
rect 22739 10675 22750 10721
rect 22920 10721 22930 10728
rect 23112 10721 23122 10728
rect 22740 10668 22750 10675
rect 22920 10675 22931 10721
rect 23111 10675 23122 10721
rect 23292 10721 23302 10728
rect 22920 10668 22930 10675
rect 23112 10668 23122 10675
rect 23292 10675 23303 10721
rect 23292 10668 23302 10675
rect 23364 10634 23422 10758
rect 23484 10721 23494 10728
rect 23483 10675 23494 10721
rect 23484 10668 23494 10675
rect 23664 10668 23866 10728
rect 24036 10721 24046 10728
rect 24036 10675 24047 10721
rect 24036 10668 24046 10675
rect 23736 10634 23794 10668
rect 24108 10634 24166 10758
rect 24228 10721 24238 10728
rect 24227 10675 24238 10721
rect 24408 10721 24418 10728
rect 24600 10721 24610 10728
rect 24228 10668 24238 10675
rect 24408 10675 24419 10721
rect 24599 10675 24610 10721
rect 24780 10721 24790 10728
rect 24408 10668 24418 10675
rect 24600 10668 24610 10675
rect 24780 10675 24791 10721
rect 24780 10668 24790 10675
rect 24852 10634 24910 10758
rect 24972 10721 24982 10728
rect 24971 10675 24982 10721
rect 24972 10668 24982 10675
rect 25152 10668 25224 10728
rect 19334 10246 19341 10622
rect 19375 10246 19382 10622
rect 19334 10194 19382 10246
rect 19593 10622 19753 10634
rect 19593 10246 19599 10622
rect 19633 10246 19713 10622
rect 19747 10246 19753 10622
rect 19593 10234 19753 10246
rect 19965 10622 20125 10634
rect 19965 10246 19971 10622
rect 20005 10246 20085 10622
rect 20119 10246 20125 10622
rect 19965 10234 20125 10246
rect 20337 10622 20497 10634
rect 20337 10246 20343 10622
rect 20377 10246 20457 10622
rect 20491 10246 20497 10622
rect 20337 10234 20497 10246
rect 20709 10622 20869 10634
rect 20709 10246 20715 10622
rect 20749 10246 20829 10622
rect 20863 10246 20869 10622
rect 20709 10234 20869 10246
rect 21081 10622 21241 10634
rect 21081 10246 21087 10622
rect 21121 10246 21201 10622
rect 21235 10246 21241 10622
rect 21081 10234 21241 10246
rect 21453 10622 21613 10634
rect 21453 10246 21459 10622
rect 21493 10246 21573 10622
rect 21607 10246 21613 10622
rect 21453 10234 21613 10246
rect 21825 10622 21985 10634
rect 21825 10246 21831 10622
rect 21865 10246 21945 10622
rect 21979 10246 21985 10622
rect 21825 10234 21985 10246
rect 22197 10622 22357 10634
rect 22197 10246 22203 10622
rect 22237 10246 22317 10622
rect 22351 10246 22357 10622
rect 22197 10234 22357 10246
rect 22569 10622 22729 10634
rect 22569 10246 22575 10622
rect 22609 10246 22689 10622
rect 22723 10246 22729 10622
rect 22569 10234 22729 10246
rect 22941 10622 23101 10634
rect 22941 10246 22947 10622
rect 22981 10246 23061 10622
rect 23095 10246 23101 10622
rect 22941 10234 23101 10246
rect 23313 10622 23473 10634
rect 23313 10246 23319 10622
rect 23353 10246 23433 10622
rect 23467 10246 23473 10622
rect 23313 10234 23473 10246
rect 23685 10622 23845 10634
rect 23685 10246 23691 10622
rect 23725 10246 23805 10622
rect 23839 10246 23845 10622
rect 23685 10234 23845 10246
rect 24057 10622 24217 10634
rect 24057 10246 24063 10622
rect 24097 10246 24177 10622
rect 24211 10246 24217 10622
rect 24057 10234 24217 10246
rect 24429 10622 24589 10634
rect 24429 10246 24435 10622
rect 24469 10246 24549 10622
rect 24583 10246 24589 10622
rect 24429 10234 24589 10246
rect 24801 10622 24961 10634
rect 24801 10246 24807 10622
rect 24841 10246 24921 10622
rect 24955 10246 24961 10622
rect 24801 10234 24961 10246
rect 25172 10622 25224 10668
rect 25172 10246 25179 10622
rect 25213 10246 25224 10622
rect 19334 10193 19422 10194
rect 19334 10188 19583 10193
rect 19334 10044 19402 10188
rect 19572 10147 19583 10188
rect 19572 10085 19582 10147
rect 19572 10044 19583 10085
rect 19334 10039 19583 10044
rect 19334 10038 19420 10039
rect 19334 9986 19382 10038
rect 19638 9998 19708 10234
rect 19763 10188 19955 10193
rect 19763 10147 19774 10188
rect 19764 10085 19774 10147
rect 19763 10044 19774 10085
rect 19944 10147 19955 10188
rect 19944 10085 19954 10147
rect 19944 10044 19955 10085
rect 19763 10039 19955 10044
rect 20010 9998 20080 10234
rect 20135 10188 20327 10193
rect 20135 10147 20146 10188
rect 20136 10085 20146 10147
rect 20135 10044 20146 10085
rect 20316 10147 20327 10188
rect 20316 10085 20326 10147
rect 20316 10044 20327 10085
rect 20135 10039 20327 10044
rect 20382 9998 20452 10234
rect 20507 10192 20699 10193
rect 20754 10192 20824 10234
rect 20879 10192 21071 10193
rect 20507 10188 21071 10192
rect 20507 10147 20518 10188
rect 20508 10085 20518 10147
rect 20507 10044 20518 10085
rect 20688 10044 20890 10188
rect 21060 10147 21071 10188
rect 21060 10085 21070 10147
rect 21060 10044 21071 10085
rect 20507 10040 21071 10044
rect 20507 10039 20699 10040
rect 20754 9998 20824 10040
rect 20879 10039 21071 10040
rect 21126 9998 21196 10234
rect 21251 10188 21443 10193
rect 21251 10147 21262 10188
rect 21252 10085 21262 10147
rect 21251 10044 21262 10085
rect 21432 10147 21443 10188
rect 21432 10085 21442 10147
rect 21432 10044 21443 10085
rect 21251 10039 21443 10044
rect 21498 9998 21568 10234
rect 21623 10188 21815 10193
rect 21623 10147 21634 10188
rect 21624 10085 21634 10147
rect 21623 10044 21634 10085
rect 21804 10147 21815 10188
rect 21804 10085 21814 10147
rect 21804 10044 21815 10085
rect 21623 10039 21815 10044
rect 21870 9998 21940 10234
rect 22242 10194 22312 10234
rect 22050 10193 22468 10194
rect 21995 10188 22559 10193
rect 21995 10147 22006 10188
rect 21996 10085 22006 10147
rect 21995 10044 22006 10085
rect 22176 10044 22378 10188
rect 22548 10147 22559 10188
rect 22548 10085 22558 10147
rect 22548 10044 22559 10085
rect 21995 10039 22559 10044
rect 22050 10038 22468 10039
rect 22242 9998 22312 10038
rect 22614 9998 22684 10234
rect 22739 10188 22931 10193
rect 22739 10147 22750 10188
rect 22740 10085 22750 10147
rect 22739 10044 22750 10085
rect 22920 10147 22931 10188
rect 22920 10085 22930 10147
rect 22920 10044 22931 10085
rect 22739 10039 22931 10044
rect 22986 9998 23056 10234
rect 23111 10188 23303 10193
rect 23111 10147 23122 10188
rect 23112 10085 23122 10147
rect 23111 10044 23122 10085
rect 23292 10147 23303 10188
rect 23292 10085 23302 10147
rect 23292 10044 23303 10085
rect 23111 10039 23303 10044
rect 23358 9998 23428 10234
rect 23730 10194 23800 10234
rect 23578 10193 23954 10194
rect 23483 10188 24047 10193
rect 23483 10147 23494 10188
rect 23484 10085 23494 10147
rect 23483 10044 23494 10085
rect 23664 10044 23866 10188
rect 24036 10147 24047 10188
rect 24036 10085 24046 10147
rect 24036 10044 24047 10085
rect 23483 10039 24047 10044
rect 23578 10038 23954 10039
rect 23730 9998 23800 10038
rect 24102 9998 24172 10234
rect 24227 10188 24419 10193
rect 24227 10147 24238 10188
rect 24228 10085 24238 10147
rect 24227 10044 24238 10085
rect 24408 10147 24419 10188
rect 24408 10085 24418 10147
rect 24408 10044 24419 10085
rect 24227 10039 24419 10044
rect 24474 9998 24544 10234
rect 24599 10188 24791 10193
rect 24599 10147 24610 10188
rect 24600 10085 24610 10147
rect 24599 10044 24610 10085
rect 24780 10147 24791 10188
rect 24780 10085 24790 10147
rect 24780 10044 24791 10085
rect 24599 10039 24791 10044
rect 24846 9998 24916 10234
rect 25172 10194 25224 10246
rect 25066 10193 25224 10194
rect 24971 10188 25224 10193
rect 24971 10147 24982 10188
rect 24972 10085 24982 10147
rect 24971 10044 24982 10085
rect 25152 10044 25224 10188
rect 24971 10039 25224 10044
rect 25066 10038 25224 10039
rect 19334 9610 19341 9986
rect 19375 9610 19382 9986
rect 19334 9558 19382 9610
rect 19593 9986 19753 9998
rect 19593 9610 19599 9986
rect 19633 9610 19713 9986
rect 19747 9610 19753 9986
rect 19593 9598 19753 9610
rect 19965 9986 20125 9998
rect 19965 9610 19971 9986
rect 20005 9610 20085 9986
rect 20119 9610 20125 9986
rect 19965 9598 20125 9610
rect 20337 9986 20497 9998
rect 20337 9610 20343 9986
rect 20377 9610 20457 9986
rect 20491 9610 20497 9986
rect 20337 9598 20497 9610
rect 20709 9986 20869 9998
rect 20709 9610 20715 9986
rect 20749 9610 20829 9986
rect 20863 9610 20869 9986
rect 20709 9598 20869 9610
rect 21081 9986 21241 9998
rect 21081 9610 21087 9986
rect 21121 9610 21201 9986
rect 21235 9610 21241 9986
rect 21081 9598 21241 9610
rect 21453 9986 21613 9998
rect 21453 9610 21459 9986
rect 21493 9610 21573 9986
rect 21607 9610 21613 9986
rect 21453 9598 21613 9610
rect 21825 9986 21985 9998
rect 21825 9610 21831 9986
rect 21865 9610 21945 9986
rect 21979 9610 21985 9986
rect 21825 9598 21985 9610
rect 22197 9986 22357 9998
rect 22197 9610 22203 9986
rect 22237 9610 22317 9986
rect 22351 9610 22357 9986
rect 22197 9598 22357 9610
rect 22569 9986 22729 9998
rect 22569 9610 22575 9986
rect 22609 9610 22689 9986
rect 22723 9610 22729 9986
rect 22569 9598 22729 9610
rect 22941 9986 23101 9998
rect 22941 9610 22947 9986
rect 22981 9610 23061 9986
rect 23095 9610 23101 9986
rect 22941 9598 23101 9610
rect 23313 9986 23473 9998
rect 23313 9610 23319 9986
rect 23353 9610 23433 9986
rect 23467 9610 23473 9986
rect 23313 9598 23473 9610
rect 23685 9986 23845 9998
rect 23685 9610 23691 9986
rect 23725 9610 23805 9986
rect 23839 9610 23845 9986
rect 23685 9598 23845 9610
rect 24057 9986 24217 9998
rect 24057 9610 24063 9986
rect 24097 9610 24177 9986
rect 24211 9610 24217 9986
rect 24057 9598 24217 9610
rect 24429 9986 24589 9998
rect 24429 9610 24435 9986
rect 24469 9610 24549 9986
rect 24583 9610 24589 9986
rect 24429 9598 24589 9610
rect 24801 9986 24961 9998
rect 24801 9610 24807 9986
rect 24841 9610 24921 9986
rect 24955 9610 24961 9986
rect 24801 9598 24961 9610
rect 25172 9986 25224 10038
rect 25172 9610 25179 9986
rect 25213 9610 25224 9986
rect 19334 9557 19424 9558
rect 19334 9552 19583 9557
rect 19334 9408 19402 9552
rect 19572 9511 19583 9552
rect 19572 9449 19582 9511
rect 19572 9408 19583 9449
rect 19334 9403 19583 9408
rect 19334 9398 19424 9403
rect 19334 9350 19382 9398
rect 19638 9362 19708 9598
rect 19763 9552 19955 9557
rect 19763 9511 19774 9552
rect 19764 9449 19774 9511
rect 19763 9408 19774 9449
rect 19944 9511 19955 9552
rect 19944 9449 19954 9511
rect 19944 9408 19955 9449
rect 19763 9403 19955 9408
rect 20010 9362 20080 9598
rect 20135 9552 20327 9557
rect 20135 9511 20146 9552
rect 20136 9449 20146 9511
rect 20135 9408 20146 9449
rect 20316 9511 20327 9552
rect 20316 9449 20326 9511
rect 20316 9408 20327 9449
rect 20135 9403 20327 9408
rect 20382 9362 20452 9598
rect 20507 9554 20699 9557
rect 20754 9554 20824 9598
rect 20879 9554 21071 9557
rect 20507 9552 21071 9554
rect 20507 9511 20518 9552
rect 20508 9449 20518 9511
rect 20507 9408 20518 9449
rect 20688 9408 20890 9552
rect 21060 9511 21071 9552
rect 21060 9449 21070 9511
rect 21060 9408 21071 9449
rect 20507 9403 21071 9408
rect 20548 9402 21024 9403
rect 20754 9362 20824 9402
rect 21126 9362 21196 9598
rect 21251 9552 21443 9557
rect 21251 9511 21262 9552
rect 21252 9449 21262 9511
rect 21251 9408 21262 9449
rect 21432 9511 21443 9552
rect 21432 9449 21442 9511
rect 21432 9408 21443 9449
rect 21251 9403 21443 9408
rect 21498 9362 21568 9598
rect 21623 9552 21815 9557
rect 21623 9511 21634 9552
rect 21624 9449 21634 9511
rect 21623 9408 21634 9449
rect 21804 9511 21815 9552
rect 21804 9449 21814 9511
rect 21804 9408 21815 9449
rect 21623 9403 21815 9408
rect 21870 9362 21940 9598
rect 22242 9558 22312 9598
rect 22070 9557 22488 9558
rect 21995 9552 22559 9557
rect 21995 9511 22006 9552
rect 21996 9449 22006 9511
rect 21995 9408 22006 9449
rect 22176 9408 22378 9552
rect 22548 9511 22559 9552
rect 22548 9449 22558 9511
rect 22548 9408 22559 9449
rect 21995 9403 22559 9408
rect 22070 9402 22488 9403
rect 22242 9362 22312 9402
rect 22614 9362 22684 9598
rect 22739 9552 22931 9557
rect 22739 9511 22750 9552
rect 22740 9449 22750 9511
rect 22739 9408 22750 9449
rect 22920 9511 22931 9552
rect 22920 9449 22930 9511
rect 22920 9408 22931 9449
rect 22739 9403 22931 9408
rect 22986 9362 23056 9598
rect 23111 9552 23303 9557
rect 23111 9511 23122 9552
rect 23112 9449 23122 9511
rect 23111 9408 23122 9449
rect 23292 9511 23303 9552
rect 23292 9449 23302 9511
rect 23292 9408 23303 9449
rect 23111 9403 23303 9408
rect 23358 9362 23428 9598
rect 23730 9558 23800 9598
rect 23566 9557 23942 9558
rect 23483 9552 24047 9557
rect 23483 9511 23494 9552
rect 23484 9449 23494 9511
rect 23483 9408 23494 9449
rect 23664 9408 23866 9552
rect 24036 9511 24047 9552
rect 24036 9449 24046 9511
rect 24036 9408 24047 9449
rect 23483 9403 24047 9408
rect 23566 9402 23942 9403
rect 23730 9362 23800 9402
rect 24102 9362 24172 9598
rect 24227 9552 24419 9557
rect 24227 9511 24238 9552
rect 24228 9449 24238 9511
rect 24227 9408 24238 9449
rect 24408 9511 24419 9552
rect 24408 9449 24418 9511
rect 24408 9408 24419 9449
rect 24227 9403 24419 9408
rect 24474 9362 24544 9598
rect 24599 9552 24791 9557
rect 24599 9511 24610 9552
rect 24600 9449 24610 9511
rect 24599 9408 24610 9449
rect 24780 9511 24791 9552
rect 24780 9449 24790 9511
rect 24780 9408 24791 9449
rect 24599 9403 24791 9408
rect 24846 9362 24916 9598
rect 25172 9558 25224 9610
rect 25082 9557 25224 9558
rect 24971 9552 25224 9557
rect 24971 9511 24982 9552
rect 24972 9449 24982 9511
rect 24971 9408 24982 9449
rect 25152 9408 25224 9552
rect 24971 9403 25224 9408
rect 25082 9402 25224 9403
rect 19334 8974 19341 9350
rect 19375 8974 19382 9350
rect 19334 8928 19382 8974
rect 19593 9350 19753 9362
rect 19593 8974 19599 9350
rect 19633 8974 19713 9350
rect 19747 8974 19753 9350
rect 19593 8962 19753 8974
rect 19965 9350 20125 9362
rect 19965 8974 19971 9350
rect 20005 8974 20085 9350
rect 20119 8974 20125 9350
rect 19965 8962 20125 8974
rect 20337 9350 20497 9362
rect 20337 8974 20343 9350
rect 20377 8974 20457 9350
rect 20491 8974 20497 9350
rect 20337 8962 20497 8974
rect 20709 9350 20869 9362
rect 20709 8974 20715 9350
rect 20749 8974 20829 9350
rect 20863 8974 20869 9350
rect 20709 8962 20869 8974
rect 21081 9350 21241 9362
rect 21081 8974 21087 9350
rect 21121 8974 21201 9350
rect 21235 8974 21241 9350
rect 21081 8962 21241 8974
rect 21453 9350 21613 9362
rect 21453 8974 21459 9350
rect 21493 8974 21573 9350
rect 21607 8974 21613 9350
rect 21453 8962 21613 8974
rect 21825 9350 21985 9362
rect 21825 8974 21831 9350
rect 21865 8974 21945 9350
rect 21979 8974 21985 9350
rect 21825 8962 21985 8974
rect 22197 9350 22357 9362
rect 22197 8974 22203 9350
rect 22237 8974 22317 9350
rect 22351 8974 22357 9350
rect 22197 8962 22357 8974
rect 22569 9350 22729 9362
rect 22569 8974 22575 9350
rect 22609 8974 22689 9350
rect 22723 8974 22729 9350
rect 22569 8962 22729 8974
rect 22941 9350 23101 9362
rect 22941 8974 22947 9350
rect 22981 8974 23061 9350
rect 23095 8974 23101 9350
rect 22941 8962 23101 8974
rect 23313 9350 23473 9362
rect 23313 8974 23319 9350
rect 23353 8974 23433 9350
rect 23467 8974 23473 9350
rect 23313 8962 23473 8974
rect 23685 9350 23845 9362
rect 23685 8974 23691 9350
rect 23725 8974 23805 9350
rect 23839 8974 23845 9350
rect 23685 8962 23845 8974
rect 24057 9350 24217 9362
rect 24057 8974 24063 9350
rect 24097 8974 24177 9350
rect 24211 8974 24217 9350
rect 24057 8962 24217 8974
rect 24429 9350 24589 9362
rect 24429 8974 24435 9350
rect 24469 8974 24549 9350
rect 24583 8974 24589 9350
rect 24429 8962 24589 8974
rect 24801 9350 24961 9362
rect 24801 8974 24807 9350
rect 24841 8974 24921 9350
rect 24955 8974 24961 9350
rect 24801 8962 24961 8974
rect 25172 9350 25224 9402
rect 25172 8974 25179 9350
rect 25213 8974 25224 9350
rect 19334 8868 19402 8928
rect 19572 8921 19582 8928
rect 19764 8921 19774 8928
rect 19572 8875 19583 8921
rect 19763 8875 19774 8921
rect 19944 8921 19954 8928
rect 19572 8868 19582 8875
rect 19764 8868 19774 8875
rect 19944 8875 19955 8921
rect 19944 8868 19954 8875
rect 20016 8620 20074 8962
rect 20760 8928 20818 8962
rect 20136 8921 20146 8928
rect 20135 8875 20146 8921
rect 20316 8921 20326 8928
rect 20508 8921 20518 8928
rect 20136 8868 20146 8875
rect 20316 8875 20327 8921
rect 20507 8875 20518 8921
rect 20316 8868 20326 8875
rect 20508 8868 20518 8875
rect 20688 8868 20890 8928
rect 21060 8921 21070 8928
rect 21252 8921 21262 8928
rect 21060 8875 21071 8921
rect 21251 8875 21262 8921
rect 21432 8921 21442 8928
rect 21060 8868 21070 8875
rect 21252 8868 21262 8875
rect 21432 8875 21443 8921
rect 21432 8868 21442 8875
rect 20634 8866 20964 8868
rect 21504 8620 21562 8962
rect 22248 8928 22306 8962
rect 21624 8921 21634 8928
rect 21623 8875 21634 8921
rect 21804 8921 21814 8928
rect 21996 8921 22006 8928
rect 21624 8868 21634 8875
rect 21804 8875 21815 8921
rect 21995 8875 22006 8921
rect 21804 8868 21814 8875
rect 21996 8868 22006 8875
rect 22176 8868 22378 8928
rect 22548 8921 22558 8928
rect 22740 8921 22750 8928
rect 22548 8875 22559 8921
rect 22739 8875 22750 8921
rect 22920 8921 22930 8928
rect 22548 8868 22558 8875
rect 22740 8868 22750 8875
rect 22920 8875 22931 8921
rect 22920 8868 22930 8875
rect 22992 8620 23050 8962
rect 23736 8928 23794 8962
rect 23112 8921 23122 8928
rect 23111 8875 23122 8921
rect 23292 8921 23302 8928
rect 23484 8921 23494 8928
rect 23112 8868 23122 8875
rect 23292 8875 23303 8921
rect 23483 8875 23494 8921
rect 23292 8868 23302 8875
rect 23484 8868 23494 8875
rect 23664 8868 23866 8928
rect 24036 8921 24046 8928
rect 24228 8921 24238 8928
rect 24036 8875 24047 8921
rect 24227 8875 24238 8921
rect 24408 8921 24418 8928
rect 24036 8868 24046 8875
rect 24228 8868 24238 8875
rect 24408 8875 24419 8921
rect 24408 8868 24418 8875
rect 24480 8620 24538 8962
rect 25172 8928 25224 8974
rect 25262 10634 25314 10758
rect 25348 10668 25354 10728
rect 25524 10721 25534 10728
rect 25716 10721 25726 10728
rect 25524 10675 25535 10721
rect 25715 10675 25726 10721
rect 25896 10721 25906 10728
rect 25524 10668 25534 10675
rect 25716 10668 25726 10675
rect 25896 10675 25907 10721
rect 25896 10668 25906 10675
rect 25968 10634 26026 10758
rect 26088 10721 26098 10728
rect 26087 10675 26098 10721
rect 26268 10721 26278 10728
rect 26460 10721 26470 10728
rect 26088 10668 26098 10675
rect 26268 10675 26279 10721
rect 26459 10675 26470 10721
rect 26640 10721 26650 10728
rect 26268 10668 26278 10675
rect 26460 10668 26470 10675
rect 26640 10675 26651 10721
rect 26640 10668 26650 10675
rect 26712 10634 26770 10758
rect 26832 10721 26842 10728
rect 26831 10675 26842 10721
rect 27012 10721 27022 10728
rect 27204 10721 27214 10728
rect 26832 10668 26842 10675
rect 27012 10675 27023 10721
rect 27203 10675 27214 10721
rect 27384 10721 27394 10728
rect 27012 10668 27022 10675
rect 27204 10668 27214 10675
rect 27384 10675 27395 10721
rect 27384 10668 27394 10675
rect 27456 10634 27514 10758
rect 27576 10721 27586 10728
rect 27575 10675 27586 10721
rect 27756 10721 27766 10728
rect 27948 10721 27958 10728
rect 27576 10668 27586 10675
rect 27756 10675 27767 10721
rect 27947 10675 27958 10721
rect 28128 10721 28138 10728
rect 27756 10668 27766 10675
rect 27948 10668 27958 10675
rect 28128 10675 28139 10721
rect 28128 10668 28138 10675
rect 28200 10634 28258 10758
rect 28320 10721 28330 10728
rect 28319 10675 28330 10721
rect 28500 10721 28510 10728
rect 28692 10721 28702 10728
rect 28320 10668 28330 10675
rect 28500 10675 28511 10721
rect 28691 10675 28702 10721
rect 28872 10721 28882 10728
rect 28500 10668 28510 10675
rect 28692 10668 28702 10675
rect 28872 10675 28883 10721
rect 28872 10668 28882 10675
rect 28944 10634 29002 10758
rect 29064 10721 29074 10728
rect 29063 10675 29074 10721
rect 29244 10721 29254 10728
rect 29436 10721 29446 10728
rect 29064 10668 29074 10675
rect 29244 10675 29255 10721
rect 29435 10675 29446 10721
rect 29616 10721 29626 10728
rect 29244 10668 29254 10675
rect 29436 10668 29446 10675
rect 29616 10675 29627 10721
rect 29616 10668 29626 10675
rect 29688 10634 29746 10758
rect 29808 10721 29818 10728
rect 29807 10675 29818 10721
rect 29988 10721 29998 10728
rect 30180 10721 30190 10728
rect 29808 10668 29818 10675
rect 29988 10675 29999 10721
rect 30179 10675 30190 10721
rect 30360 10721 30370 10728
rect 29988 10668 29998 10675
rect 30180 10668 30190 10675
rect 30360 10675 30371 10721
rect 30360 10668 30370 10675
rect 30432 10634 30490 10758
rect 30552 10721 30562 10728
rect 30551 10675 30562 10721
rect 30732 10721 30742 10728
rect 30924 10721 30934 10728
rect 30552 10668 30562 10675
rect 30732 10675 30743 10721
rect 30923 10675 30934 10721
rect 31104 10721 31114 10728
rect 30732 10668 30742 10675
rect 30924 10668 30934 10675
rect 31104 10675 31115 10721
rect 31104 10668 31114 10675
rect 31158 10634 31216 10758
rect 25262 10622 25333 10634
rect 25262 10246 25293 10622
rect 25327 10246 25333 10622
rect 25262 10234 25333 10246
rect 25545 10622 25705 10634
rect 25545 10246 25551 10622
rect 25585 10246 25665 10622
rect 25699 10246 25705 10622
rect 25545 10234 25705 10246
rect 25917 10622 26077 10634
rect 25917 10246 25923 10622
rect 25957 10246 26037 10622
rect 26071 10246 26077 10622
rect 25917 10234 26077 10246
rect 26289 10622 26449 10634
rect 26289 10246 26295 10622
rect 26329 10246 26409 10622
rect 26443 10246 26449 10622
rect 26289 10234 26449 10246
rect 26661 10622 26821 10634
rect 26661 10246 26667 10622
rect 26701 10246 26781 10622
rect 26815 10246 26821 10622
rect 26661 10234 26821 10246
rect 27033 10622 27193 10634
rect 27033 10246 27039 10622
rect 27073 10246 27153 10622
rect 27187 10246 27193 10622
rect 27033 10234 27193 10246
rect 27405 10622 27565 10634
rect 27405 10246 27411 10622
rect 27445 10246 27525 10622
rect 27559 10246 27565 10622
rect 27405 10234 27565 10246
rect 27777 10622 27937 10634
rect 27777 10246 27783 10622
rect 27817 10246 27897 10622
rect 27931 10246 27937 10622
rect 27777 10234 27937 10246
rect 28149 10622 28309 10634
rect 28149 10246 28155 10622
rect 28189 10246 28269 10622
rect 28303 10246 28309 10622
rect 28149 10234 28309 10246
rect 28521 10622 28681 10634
rect 28521 10246 28527 10622
rect 28561 10246 28641 10622
rect 28675 10246 28681 10622
rect 28521 10234 28681 10246
rect 28893 10622 29053 10634
rect 28893 10246 28899 10622
rect 28933 10246 29013 10622
rect 29047 10246 29053 10622
rect 28893 10234 29053 10246
rect 29265 10622 29425 10634
rect 29265 10246 29271 10622
rect 29305 10246 29385 10622
rect 29419 10246 29425 10622
rect 29265 10234 29425 10246
rect 29637 10622 29797 10634
rect 29637 10246 29643 10622
rect 29677 10246 29757 10622
rect 29791 10246 29797 10622
rect 29637 10234 29797 10246
rect 30009 10622 30169 10634
rect 30009 10246 30015 10622
rect 30049 10246 30129 10622
rect 30163 10246 30169 10622
rect 30009 10234 30169 10246
rect 30381 10622 30541 10634
rect 30381 10246 30387 10622
rect 30421 10246 30501 10622
rect 30535 10246 30541 10622
rect 30381 10234 30541 10246
rect 30753 10622 30913 10634
rect 30753 10246 30759 10622
rect 30793 10246 30873 10622
rect 30907 10246 30913 10622
rect 30753 10234 30913 10246
rect 31125 10622 31216 10634
rect 31125 10246 31131 10622
rect 31165 10246 31216 10622
rect 31125 10234 31216 10246
rect 25262 9998 25314 10234
rect 25342 10193 25468 10194
rect 25342 10188 25535 10193
rect 25342 10044 25354 10188
rect 25524 10147 25535 10188
rect 25524 10085 25534 10147
rect 25524 10044 25535 10085
rect 25342 10039 25535 10044
rect 25342 10038 25468 10039
rect 25590 9998 25660 10234
rect 25715 10188 25907 10193
rect 25715 10147 25726 10188
rect 25716 10085 25726 10147
rect 25715 10044 25726 10085
rect 25896 10147 25907 10188
rect 25896 10085 25906 10147
rect 25896 10044 25907 10085
rect 25715 10039 25907 10044
rect 25962 9998 26032 10234
rect 26087 10188 26279 10193
rect 26087 10147 26098 10188
rect 26088 10085 26098 10147
rect 26087 10044 26098 10085
rect 26268 10147 26279 10188
rect 26268 10085 26278 10147
rect 26268 10044 26279 10085
rect 26087 10039 26279 10044
rect 26334 9998 26404 10234
rect 26459 10188 26651 10193
rect 26459 10147 26470 10188
rect 26460 10085 26470 10147
rect 26459 10044 26470 10085
rect 26640 10147 26651 10188
rect 26640 10085 26650 10147
rect 26640 10044 26651 10085
rect 26459 10039 26651 10044
rect 26706 9998 26776 10234
rect 26831 10188 27023 10193
rect 26831 10147 26842 10188
rect 26832 10085 26842 10147
rect 26831 10044 26842 10085
rect 27012 10147 27023 10188
rect 27012 10085 27022 10147
rect 27012 10044 27023 10085
rect 26831 10039 27023 10044
rect 27078 9998 27148 10234
rect 27203 10188 27395 10193
rect 27203 10147 27214 10188
rect 27204 10085 27214 10147
rect 27203 10044 27214 10085
rect 27384 10147 27395 10188
rect 27384 10085 27394 10147
rect 27384 10044 27395 10085
rect 27203 10039 27395 10044
rect 27450 9998 27520 10234
rect 27575 10188 27767 10193
rect 27575 10147 27586 10188
rect 27576 10085 27586 10147
rect 27575 10044 27586 10085
rect 27756 10147 27767 10188
rect 27756 10085 27766 10147
rect 27756 10044 27767 10085
rect 27575 10039 27767 10044
rect 27822 9998 27892 10234
rect 27947 10188 28139 10193
rect 27947 10147 27958 10188
rect 27948 10085 27958 10147
rect 27947 10044 27958 10085
rect 28128 10147 28139 10188
rect 28128 10085 28138 10147
rect 28128 10044 28139 10085
rect 27947 10039 28139 10044
rect 28194 9998 28264 10234
rect 28319 10188 28511 10193
rect 28319 10147 28330 10188
rect 28320 10085 28330 10147
rect 28319 10044 28330 10085
rect 28500 10147 28511 10188
rect 28500 10085 28510 10147
rect 28500 10044 28511 10085
rect 28319 10039 28511 10044
rect 28566 9998 28636 10234
rect 28691 10188 28883 10193
rect 28691 10147 28702 10188
rect 28692 10085 28702 10147
rect 28691 10044 28702 10085
rect 28872 10147 28883 10188
rect 28872 10085 28882 10147
rect 28872 10044 28883 10085
rect 28691 10039 28883 10044
rect 28938 9998 29008 10234
rect 29063 10188 29255 10193
rect 29063 10147 29074 10188
rect 29064 10085 29074 10147
rect 29063 10044 29074 10085
rect 29244 10147 29255 10188
rect 29244 10085 29254 10147
rect 29244 10044 29255 10085
rect 29063 10039 29255 10044
rect 29310 9998 29380 10234
rect 29435 10188 29627 10193
rect 29435 10147 29446 10188
rect 29436 10085 29446 10147
rect 29435 10044 29446 10085
rect 29616 10147 29627 10188
rect 29616 10085 29626 10147
rect 29616 10044 29627 10085
rect 29435 10039 29627 10044
rect 29682 9998 29752 10234
rect 29807 10188 29999 10193
rect 29807 10147 29818 10188
rect 29808 10085 29818 10147
rect 29807 10044 29818 10085
rect 29988 10147 29999 10188
rect 29988 10085 29998 10147
rect 29988 10044 29999 10085
rect 29807 10039 29999 10044
rect 30054 9998 30124 10234
rect 30179 10188 30371 10193
rect 30179 10147 30190 10188
rect 30180 10085 30190 10147
rect 30179 10044 30190 10085
rect 30360 10147 30371 10188
rect 30360 10085 30370 10147
rect 30360 10044 30371 10085
rect 30179 10039 30371 10044
rect 30426 9998 30496 10234
rect 30551 10188 30743 10193
rect 30551 10147 30562 10188
rect 30552 10085 30562 10147
rect 30551 10044 30562 10085
rect 30732 10147 30743 10188
rect 30732 10085 30742 10147
rect 30732 10044 30743 10085
rect 30551 10039 30743 10044
rect 30798 9998 30868 10234
rect 30923 10188 31115 10193
rect 30923 10147 30934 10188
rect 30924 10085 30934 10147
rect 30923 10044 30934 10085
rect 31104 10147 31115 10188
rect 31104 10085 31114 10147
rect 31104 10044 31115 10085
rect 30923 10039 31115 10044
rect 31158 9998 31216 10234
rect 25262 9986 25333 9998
rect 25262 9610 25293 9986
rect 25327 9610 25333 9986
rect 25262 9598 25333 9610
rect 25545 9986 25705 9998
rect 25545 9610 25551 9986
rect 25585 9610 25665 9986
rect 25699 9610 25705 9986
rect 25545 9598 25705 9610
rect 25917 9986 26077 9998
rect 25917 9610 25923 9986
rect 25957 9610 26037 9986
rect 26071 9610 26077 9986
rect 25917 9598 26077 9610
rect 26289 9986 26449 9998
rect 26289 9610 26295 9986
rect 26329 9610 26409 9986
rect 26443 9610 26449 9986
rect 26289 9598 26449 9610
rect 26661 9986 26821 9998
rect 26661 9610 26667 9986
rect 26701 9610 26781 9986
rect 26815 9610 26821 9986
rect 26661 9598 26821 9610
rect 27033 9986 27193 9998
rect 27033 9610 27039 9986
rect 27073 9610 27153 9986
rect 27187 9610 27193 9986
rect 27033 9598 27193 9610
rect 27405 9986 27565 9998
rect 27405 9610 27411 9986
rect 27445 9610 27525 9986
rect 27559 9610 27565 9986
rect 27405 9598 27565 9610
rect 27777 9986 27937 9998
rect 27777 9610 27783 9986
rect 27817 9610 27897 9986
rect 27931 9610 27937 9986
rect 27777 9598 27937 9610
rect 28149 9986 28309 9998
rect 28149 9610 28155 9986
rect 28189 9610 28269 9986
rect 28303 9610 28309 9986
rect 28149 9598 28309 9610
rect 28521 9986 28681 9998
rect 28521 9610 28527 9986
rect 28561 9610 28641 9986
rect 28675 9610 28681 9986
rect 28521 9598 28681 9610
rect 28893 9986 29053 9998
rect 28893 9610 28899 9986
rect 28933 9610 29013 9986
rect 29047 9610 29053 9986
rect 28893 9598 29053 9610
rect 29265 9986 29425 9998
rect 29265 9610 29271 9986
rect 29305 9610 29385 9986
rect 29419 9610 29425 9986
rect 29265 9598 29425 9610
rect 29637 9986 29797 9998
rect 29637 9610 29643 9986
rect 29677 9610 29757 9986
rect 29791 9610 29797 9986
rect 29637 9598 29797 9610
rect 30009 9986 30169 9998
rect 30009 9610 30015 9986
rect 30049 9610 30129 9986
rect 30163 9610 30169 9986
rect 30009 9598 30169 9610
rect 30381 9986 30541 9998
rect 30381 9610 30387 9986
rect 30421 9610 30501 9986
rect 30535 9610 30541 9986
rect 30381 9598 30541 9610
rect 30753 9986 30913 9998
rect 30753 9610 30759 9986
rect 30793 9610 30873 9986
rect 30907 9610 30913 9986
rect 30753 9598 30913 9610
rect 31125 9986 31216 9998
rect 31125 9610 31131 9986
rect 31165 9610 31216 9986
rect 31125 9598 31216 9610
rect 25262 9362 25314 9598
rect 25342 9557 25484 9558
rect 25342 9552 25535 9557
rect 25342 9408 25354 9552
rect 25524 9511 25535 9552
rect 25524 9449 25534 9511
rect 25524 9408 25535 9449
rect 25342 9403 25535 9408
rect 25342 9402 25484 9403
rect 25590 9362 25660 9598
rect 25715 9552 25907 9557
rect 25715 9511 25726 9552
rect 25716 9449 25726 9511
rect 25715 9408 25726 9449
rect 25896 9511 25907 9552
rect 25896 9449 25906 9511
rect 25896 9408 25907 9449
rect 25715 9403 25907 9408
rect 25962 9362 26032 9598
rect 26087 9552 26279 9557
rect 26087 9511 26098 9552
rect 26088 9449 26098 9511
rect 26087 9408 26098 9449
rect 26268 9511 26279 9552
rect 26268 9449 26278 9511
rect 26268 9408 26279 9449
rect 26087 9403 26279 9408
rect 26334 9362 26404 9598
rect 26459 9552 26651 9557
rect 26459 9511 26470 9552
rect 26460 9449 26470 9511
rect 26459 9408 26470 9449
rect 26640 9511 26651 9552
rect 26640 9449 26650 9511
rect 26640 9408 26651 9449
rect 26459 9403 26651 9408
rect 26706 9362 26776 9598
rect 26831 9552 27023 9557
rect 26831 9511 26842 9552
rect 26832 9449 26842 9511
rect 26831 9408 26842 9449
rect 27012 9511 27023 9552
rect 27012 9449 27022 9511
rect 27012 9408 27023 9449
rect 26831 9403 27023 9408
rect 27078 9362 27148 9598
rect 27203 9552 27395 9557
rect 27203 9511 27214 9552
rect 27204 9449 27214 9511
rect 27203 9408 27214 9449
rect 27384 9511 27395 9552
rect 27384 9449 27394 9511
rect 27384 9408 27395 9449
rect 27203 9403 27395 9408
rect 27450 9362 27520 9598
rect 27575 9552 27767 9557
rect 27575 9511 27586 9552
rect 27576 9449 27586 9511
rect 27575 9408 27586 9449
rect 27756 9511 27767 9552
rect 27756 9449 27766 9511
rect 27756 9408 27767 9449
rect 27575 9403 27767 9408
rect 27822 9362 27892 9598
rect 27947 9552 28139 9557
rect 27947 9511 27958 9552
rect 27948 9449 27958 9511
rect 27947 9408 27958 9449
rect 28128 9511 28139 9552
rect 28128 9449 28138 9511
rect 28128 9408 28139 9449
rect 27947 9403 28139 9408
rect 28194 9362 28264 9598
rect 28319 9552 28511 9557
rect 28319 9511 28330 9552
rect 28320 9449 28330 9511
rect 28319 9408 28330 9449
rect 28500 9511 28511 9552
rect 28500 9449 28510 9511
rect 28500 9408 28511 9449
rect 28319 9403 28511 9408
rect 28566 9362 28636 9598
rect 28691 9552 28883 9557
rect 28691 9511 28702 9552
rect 28692 9449 28702 9511
rect 28691 9408 28702 9449
rect 28872 9511 28883 9552
rect 28872 9449 28882 9511
rect 28872 9408 28883 9449
rect 28691 9403 28883 9408
rect 28938 9362 29008 9598
rect 29063 9552 29255 9557
rect 29063 9511 29074 9552
rect 29064 9449 29074 9511
rect 29063 9408 29074 9449
rect 29244 9511 29255 9552
rect 29244 9449 29254 9511
rect 29244 9408 29255 9449
rect 29063 9403 29255 9408
rect 29310 9362 29380 9598
rect 29435 9552 29627 9557
rect 29435 9511 29446 9552
rect 29436 9449 29446 9511
rect 29435 9408 29446 9449
rect 29616 9511 29627 9552
rect 29616 9449 29626 9511
rect 29616 9408 29627 9449
rect 29435 9403 29627 9408
rect 29682 9362 29752 9598
rect 29807 9552 29999 9557
rect 29807 9511 29818 9552
rect 29808 9449 29818 9511
rect 29807 9408 29818 9449
rect 29988 9511 29999 9552
rect 29988 9449 29998 9511
rect 29988 9408 29999 9449
rect 29807 9403 29999 9408
rect 30054 9362 30124 9598
rect 30179 9552 30371 9557
rect 30179 9511 30190 9552
rect 30180 9449 30190 9511
rect 30179 9408 30190 9449
rect 30360 9511 30371 9552
rect 30360 9449 30370 9511
rect 30360 9408 30371 9449
rect 30179 9403 30371 9408
rect 30426 9362 30496 9598
rect 30551 9552 30743 9557
rect 30551 9511 30562 9552
rect 30552 9449 30562 9511
rect 30551 9408 30562 9449
rect 30732 9511 30743 9552
rect 30732 9449 30742 9511
rect 30732 9408 30743 9449
rect 30551 9403 30743 9408
rect 30798 9362 30868 9598
rect 30923 9552 31115 9557
rect 30923 9511 30934 9552
rect 30924 9449 30934 9511
rect 30923 9408 30934 9449
rect 31104 9511 31115 9552
rect 31104 9449 31114 9511
rect 31104 9408 31115 9449
rect 30923 9403 31115 9408
rect 31158 9362 31216 9598
rect 25262 9350 25333 9362
rect 25262 8974 25293 9350
rect 25327 8974 25333 9350
rect 25262 8962 25333 8974
rect 25545 9350 25705 9362
rect 25545 8974 25551 9350
rect 25585 8974 25665 9350
rect 25699 8974 25705 9350
rect 25545 8962 25705 8974
rect 25917 9350 26077 9362
rect 25917 8974 25923 9350
rect 25957 8974 26037 9350
rect 26071 8974 26077 9350
rect 25917 8962 26077 8974
rect 26289 9350 26449 9362
rect 26289 8974 26295 9350
rect 26329 8974 26409 9350
rect 26443 8974 26449 9350
rect 26289 8962 26449 8974
rect 26661 9350 26821 9362
rect 26661 8974 26667 9350
rect 26701 8974 26781 9350
rect 26815 8974 26821 9350
rect 26661 8962 26821 8974
rect 27033 9350 27193 9362
rect 27033 8974 27039 9350
rect 27073 8974 27153 9350
rect 27187 8974 27193 9350
rect 27033 8962 27193 8974
rect 27405 9350 27565 9362
rect 27405 8974 27411 9350
rect 27445 8974 27525 9350
rect 27559 8974 27565 9350
rect 27405 8962 27565 8974
rect 27777 9350 27937 9362
rect 27777 8974 27783 9350
rect 27817 8974 27897 9350
rect 27931 8974 27937 9350
rect 27777 8962 27937 8974
rect 28149 9350 28309 9362
rect 28149 8974 28155 9350
rect 28189 8974 28269 9350
rect 28303 8974 28309 9350
rect 28149 8962 28309 8974
rect 28521 9350 28681 9362
rect 28521 8974 28527 9350
rect 28561 8974 28641 9350
rect 28675 8974 28681 9350
rect 28521 8962 28681 8974
rect 28893 9350 29053 9362
rect 28893 8974 28899 9350
rect 28933 8974 29013 9350
rect 29047 8974 29053 9350
rect 28893 8962 29053 8974
rect 29265 9350 29425 9362
rect 29265 8974 29271 9350
rect 29305 8974 29385 9350
rect 29419 8974 29425 9350
rect 29265 8962 29425 8974
rect 29637 9350 29797 9362
rect 29637 8974 29643 9350
rect 29677 8974 29757 9350
rect 29791 8974 29797 9350
rect 29637 8962 29797 8974
rect 30009 9350 30169 9362
rect 30009 8974 30015 9350
rect 30049 8974 30129 9350
rect 30163 8974 30169 9350
rect 30009 8962 30169 8974
rect 30381 9350 30541 9362
rect 30381 8974 30387 9350
rect 30421 8974 30501 9350
rect 30535 8974 30541 9350
rect 30381 8962 30541 8974
rect 30753 9350 30913 9362
rect 30753 8974 30759 9350
rect 30793 8974 30873 9350
rect 30907 8974 30913 9350
rect 30753 8962 30913 8974
rect 31125 9350 31216 9362
rect 31125 8974 31131 9350
rect 31165 8974 31216 9350
rect 31125 8962 31216 8974
rect 24600 8921 24610 8928
rect 24599 8875 24610 8921
rect 24780 8921 24790 8928
rect 24972 8921 24982 8928
rect 24600 8868 24610 8875
rect 24780 8875 24791 8921
rect 24971 8875 24982 8921
rect 24780 8868 24790 8875
rect 24972 8868 24982 8875
rect 25152 8868 25224 8928
rect 25340 8868 25354 8928
rect 25524 8921 25534 8928
rect 25524 8875 25535 8921
rect 25524 8868 25534 8875
rect 20016 8556 24538 8620
rect 25590 8720 25660 8962
rect 25716 8921 25726 8928
rect 25715 8875 25726 8921
rect 25896 8921 25906 8928
rect 26088 8921 26098 8928
rect 25716 8868 25726 8875
rect 25896 8875 25907 8921
rect 26087 8875 26098 8921
rect 26268 8921 26278 8928
rect 25896 8868 25906 8875
rect 26088 8868 26098 8875
rect 26268 8875 26279 8921
rect 26268 8868 26278 8875
rect 26334 8720 26404 8962
rect 26460 8921 26470 8928
rect 26459 8875 26470 8921
rect 26640 8921 26650 8928
rect 26832 8921 26842 8928
rect 26460 8868 26470 8875
rect 26640 8875 26651 8921
rect 26831 8875 26842 8921
rect 27012 8921 27022 8928
rect 26640 8868 26650 8875
rect 26832 8868 26842 8875
rect 27012 8875 27023 8921
rect 27012 8868 27022 8875
rect 27078 8720 27148 8962
rect 27204 8921 27214 8928
rect 27203 8875 27214 8921
rect 27384 8921 27394 8928
rect 27576 8921 27586 8928
rect 27204 8868 27214 8875
rect 27384 8875 27395 8921
rect 27575 8875 27586 8921
rect 27756 8921 27766 8928
rect 27384 8868 27394 8875
rect 27576 8868 27586 8875
rect 27756 8875 27767 8921
rect 27756 8868 27766 8875
rect 27822 8720 27892 8962
rect 27948 8921 27958 8928
rect 27947 8875 27958 8921
rect 28128 8921 28138 8928
rect 28320 8921 28330 8928
rect 27948 8868 27958 8875
rect 28128 8875 28139 8921
rect 28319 8875 28330 8921
rect 28500 8921 28510 8928
rect 28128 8868 28138 8875
rect 28320 8868 28330 8875
rect 28500 8875 28511 8921
rect 28500 8868 28510 8875
rect 28566 8720 28636 8962
rect 28692 8921 28702 8928
rect 28691 8875 28702 8921
rect 28872 8921 28882 8928
rect 29064 8921 29074 8928
rect 28692 8868 28702 8875
rect 28872 8875 28883 8921
rect 29063 8875 29074 8921
rect 29244 8921 29254 8928
rect 28872 8868 28882 8875
rect 29064 8868 29074 8875
rect 29244 8875 29255 8921
rect 29244 8868 29254 8875
rect 29310 8720 29380 8962
rect 29436 8921 29446 8928
rect 29435 8875 29446 8921
rect 29616 8921 29626 8928
rect 29808 8921 29818 8928
rect 29436 8868 29446 8875
rect 29616 8875 29627 8921
rect 29807 8875 29818 8921
rect 29988 8921 29998 8928
rect 29616 8868 29626 8875
rect 29808 8868 29818 8875
rect 29988 8875 29999 8921
rect 29988 8868 29998 8875
rect 30054 8720 30124 8962
rect 30180 8921 30190 8928
rect 30179 8875 30190 8921
rect 30360 8921 30370 8928
rect 30552 8921 30562 8928
rect 30180 8868 30190 8875
rect 30360 8875 30371 8921
rect 30551 8875 30562 8921
rect 30732 8921 30742 8928
rect 30360 8868 30370 8875
rect 30552 8868 30562 8875
rect 30732 8875 30743 8921
rect 30732 8868 30742 8875
rect 30798 8720 30868 8962
rect 30924 8921 30934 8928
rect 30923 8875 30934 8921
rect 31104 8921 31114 8928
rect 30924 8868 30934 8875
rect 31104 8875 31115 8921
rect 31104 8868 31114 8875
rect 25590 8572 30868 8720
rect 20776 8452 20830 8556
rect 21172 8452 21242 8556
rect 21504 8452 21562 8556
rect 21916 8452 21986 8556
rect 22248 8452 22306 8556
rect 22660 8452 22730 8556
rect 22992 8452 23050 8556
rect 23404 8452 23474 8556
rect 23724 8452 23778 8556
rect 20776 8446 20882 8452
rect 20776 8376 20800 8446
rect 20870 8376 20882 8446
rect 20776 8370 20882 8376
rect 21160 8446 21254 8452
rect 21160 8376 21172 8446
rect 21242 8376 21254 8446
rect 21160 8370 21254 8376
rect 21504 8446 21626 8452
rect 21504 8376 21544 8446
rect 21614 8376 21626 8446
rect 21504 8370 21626 8376
rect 21904 8446 21998 8452
rect 21904 8376 21916 8446
rect 21986 8376 21998 8446
rect 21904 8370 21998 8376
rect 22248 8446 22370 8452
rect 22248 8376 22288 8446
rect 22358 8376 22370 8446
rect 22248 8370 22370 8376
rect 22648 8446 22742 8452
rect 22648 8376 22660 8446
rect 22730 8376 22742 8446
rect 22648 8370 22742 8376
rect 22992 8446 23114 8452
rect 22992 8376 23032 8446
rect 23102 8376 23114 8446
rect 22992 8370 23114 8376
rect 23392 8446 23486 8452
rect 23392 8376 23404 8446
rect 23474 8376 23486 8446
rect 23392 8370 23486 8376
rect 23654 8446 23778 8452
rect 23654 8376 23666 8446
rect 23736 8376 23778 8446
rect 23654 8370 23778 8376
rect 20776 8246 20830 8370
rect 20880 8333 20890 8342
rect 20879 8287 20890 8333
rect 21060 8333 21070 8342
rect 21252 8333 21262 8342
rect 20880 8278 20890 8287
rect 21060 8287 21071 8333
rect 21251 8287 21262 8333
rect 21432 8333 21442 8342
rect 21060 8278 21070 8287
rect 21252 8278 21262 8287
rect 21432 8287 21443 8333
rect 21432 8278 21442 8287
rect 21504 8246 21562 8370
rect 21624 8333 21634 8342
rect 21623 8287 21634 8333
rect 21804 8333 21814 8342
rect 21996 8333 22006 8342
rect 21624 8278 21634 8287
rect 21804 8287 21815 8333
rect 21995 8287 22006 8333
rect 22176 8333 22186 8342
rect 21804 8278 21814 8287
rect 21996 8278 22006 8287
rect 22176 8287 22187 8333
rect 22176 8278 22186 8287
rect 22248 8246 22306 8370
rect 22368 8333 22378 8342
rect 22367 8287 22378 8333
rect 22548 8333 22558 8342
rect 22740 8333 22750 8342
rect 22368 8278 22378 8287
rect 22548 8287 22559 8333
rect 22739 8287 22750 8333
rect 22920 8333 22930 8342
rect 22548 8278 22558 8287
rect 22740 8278 22750 8287
rect 22920 8287 22931 8333
rect 22920 8278 22930 8287
rect 22992 8246 23050 8370
rect 23112 8333 23122 8342
rect 23111 8287 23122 8333
rect 23292 8333 23302 8342
rect 23484 8333 23494 8342
rect 23112 8278 23122 8287
rect 23292 8287 23303 8333
rect 23483 8287 23494 8333
rect 23664 8333 23674 8342
rect 23292 8278 23302 8287
rect 23484 8278 23494 8287
rect 23664 8287 23675 8333
rect 23664 8278 23674 8287
rect 23724 8246 23778 8370
rect 20776 8234 20869 8246
rect 20776 7458 20829 8234
rect 20863 7458 20869 8234
rect 20776 7446 20869 7458
rect 21081 8234 21241 8246
rect 21081 7458 21087 8234
rect 21121 7458 21201 8234
rect 21235 7458 21241 8234
rect 21081 7446 21241 7458
rect 21453 8234 21613 8246
rect 21453 7458 21459 8234
rect 21493 7458 21573 8234
rect 21607 7458 21613 8234
rect 21453 7446 21613 7458
rect 21825 8234 21985 8246
rect 21825 7458 21831 8234
rect 21865 7458 21945 8234
rect 21979 7458 21985 8234
rect 21825 7446 21985 7458
rect 22197 8234 22357 8246
rect 22197 7458 22203 8234
rect 22237 7458 22317 8234
rect 22351 7458 22357 8234
rect 22197 7446 22357 7458
rect 22569 8234 22729 8246
rect 22569 7458 22575 8234
rect 22609 7458 22689 8234
rect 22723 7458 22729 8234
rect 22569 7446 22729 7458
rect 22941 8234 23101 8246
rect 22941 7458 22947 8234
rect 22981 7458 23061 8234
rect 23095 7458 23101 8234
rect 22941 7446 23101 7458
rect 23313 8234 23473 8246
rect 23313 7458 23319 8234
rect 23353 7458 23433 8234
rect 23467 7458 23473 8234
rect 23313 7446 23473 7458
rect 23685 8234 23778 8246
rect 23685 7458 23691 8234
rect 23725 7458 23778 8234
rect 23685 7446 23778 7458
rect 20776 7210 20824 7446
rect 20879 7400 21071 7405
rect 20879 7359 20890 7400
rect 20880 7297 20890 7359
rect 20879 7256 20890 7297
rect 21060 7359 21071 7400
rect 21060 7297 21070 7359
rect 21060 7256 21071 7297
rect 20879 7251 21071 7256
rect 21126 7210 21196 7446
rect 21251 7400 21443 7405
rect 21251 7359 21262 7400
rect 21252 7297 21262 7359
rect 21251 7256 21262 7297
rect 21432 7359 21443 7400
rect 21432 7297 21442 7359
rect 21432 7256 21443 7297
rect 21251 7251 21443 7256
rect 21498 7210 21568 7446
rect 21623 7400 21815 7405
rect 21623 7359 21634 7400
rect 21624 7297 21634 7359
rect 21623 7256 21634 7297
rect 21804 7359 21815 7400
rect 21804 7297 21814 7359
rect 21804 7256 21815 7297
rect 21623 7251 21815 7256
rect 21870 7210 21940 7446
rect 21995 7400 22187 7405
rect 21995 7359 22006 7400
rect 21996 7297 22006 7359
rect 21995 7256 22006 7297
rect 22176 7359 22187 7400
rect 22176 7297 22186 7359
rect 22176 7256 22187 7297
rect 21995 7251 22187 7256
rect 22242 7210 22312 7446
rect 22367 7400 22559 7405
rect 22367 7359 22378 7400
rect 22368 7297 22378 7359
rect 22367 7256 22378 7297
rect 22548 7359 22559 7400
rect 22548 7297 22558 7359
rect 22548 7256 22559 7297
rect 22367 7251 22559 7256
rect 22614 7210 22684 7446
rect 22739 7400 22931 7405
rect 22739 7359 22750 7400
rect 22740 7297 22750 7359
rect 22739 7256 22750 7297
rect 22920 7359 22931 7400
rect 22920 7297 22930 7359
rect 22920 7256 22931 7297
rect 22739 7251 22931 7256
rect 22986 7210 23056 7446
rect 23111 7400 23303 7405
rect 23111 7359 23122 7400
rect 23112 7297 23122 7359
rect 23111 7256 23122 7297
rect 23292 7359 23303 7400
rect 23292 7297 23302 7359
rect 23292 7256 23303 7297
rect 23111 7251 23303 7256
rect 23358 7210 23428 7446
rect 23483 7400 23675 7405
rect 23483 7359 23494 7400
rect 23484 7297 23494 7359
rect 23483 7256 23494 7297
rect 23664 7359 23675 7400
rect 23664 7297 23674 7359
rect 23664 7256 23675 7297
rect 23483 7251 23675 7256
rect 23724 7210 23778 7446
rect 20776 7198 20869 7210
rect 20776 6422 20829 7198
rect 20863 6422 20869 7198
rect 20776 6410 20869 6422
rect 21081 7198 21241 7210
rect 21081 6422 21087 7198
rect 21121 6422 21201 7198
rect 21235 6422 21241 7198
rect 21081 6410 21241 6422
rect 21453 7198 21613 7210
rect 21453 6422 21459 7198
rect 21493 6422 21573 7198
rect 21607 6422 21613 7198
rect 21453 6410 21613 6422
rect 21825 7198 21985 7210
rect 21825 6422 21831 7198
rect 21865 6422 21945 7198
rect 21979 6422 21985 7198
rect 21825 6410 21985 6422
rect 22197 7198 22357 7210
rect 22197 6422 22203 7198
rect 22237 6422 22317 7198
rect 22351 6422 22357 7198
rect 22197 6410 22357 6422
rect 22569 7198 22729 7210
rect 22569 6422 22575 7198
rect 22609 6422 22689 7198
rect 22723 6422 22729 7198
rect 22569 6410 22729 6422
rect 22941 7198 23101 7210
rect 22941 6422 22947 7198
rect 22981 6422 23061 7198
rect 23095 6422 23101 7198
rect 22941 6410 23101 6422
rect 23313 7198 23473 7210
rect 23313 6422 23319 7198
rect 23353 6422 23433 7198
rect 23467 6422 23473 7198
rect 23313 6410 23473 6422
rect 23685 7198 23778 7210
rect 23685 6422 23691 7198
rect 23725 6422 23778 7198
rect 23685 6410 23778 6422
rect 20776 6174 20824 6410
rect 20879 6364 21071 6369
rect 20879 6323 20890 6364
rect 20880 6261 20890 6323
rect 20879 6220 20890 6261
rect 21060 6323 21071 6364
rect 21060 6261 21070 6323
rect 21060 6220 21071 6261
rect 20879 6215 21071 6220
rect 21126 6174 21196 6410
rect 21251 6364 21443 6369
rect 21251 6323 21262 6364
rect 21252 6261 21262 6323
rect 21251 6220 21262 6261
rect 21432 6323 21443 6364
rect 21432 6261 21442 6323
rect 21432 6220 21443 6261
rect 21251 6215 21443 6220
rect 21498 6174 21568 6410
rect 21623 6364 21815 6369
rect 21623 6323 21634 6364
rect 21624 6261 21634 6323
rect 21623 6220 21634 6261
rect 21804 6323 21815 6364
rect 21804 6261 21814 6323
rect 21804 6220 21815 6261
rect 21623 6215 21815 6220
rect 21870 6174 21940 6410
rect 21995 6364 22187 6369
rect 21995 6323 22006 6364
rect 21996 6261 22006 6323
rect 21995 6220 22006 6261
rect 22176 6323 22187 6364
rect 22176 6261 22186 6323
rect 22176 6220 22187 6261
rect 21995 6215 22187 6220
rect 22242 6174 22312 6410
rect 22367 6364 22559 6369
rect 22367 6323 22378 6364
rect 22368 6261 22378 6323
rect 22367 6220 22378 6261
rect 22548 6323 22559 6364
rect 22548 6261 22558 6323
rect 22548 6220 22559 6261
rect 22367 6215 22559 6220
rect 22614 6174 22684 6410
rect 22739 6364 22931 6369
rect 22739 6323 22750 6364
rect 22740 6261 22750 6323
rect 22739 6220 22750 6261
rect 22920 6323 22931 6364
rect 22920 6261 22930 6323
rect 22920 6220 22931 6261
rect 22739 6215 22931 6220
rect 22986 6174 23056 6410
rect 23111 6364 23303 6369
rect 23111 6323 23122 6364
rect 23112 6261 23122 6323
rect 23111 6220 23122 6261
rect 23292 6323 23303 6364
rect 23292 6261 23302 6323
rect 23292 6220 23303 6261
rect 23111 6215 23303 6220
rect 23358 6174 23428 6410
rect 23483 6364 23675 6369
rect 23483 6323 23494 6364
rect 23484 6261 23494 6323
rect 23483 6220 23494 6261
rect 23664 6323 23675 6364
rect 23664 6261 23674 6323
rect 23664 6220 23675 6261
rect 23483 6215 23675 6220
rect 23724 6174 23778 6410
rect 20776 6162 20869 6174
rect 20776 5386 20829 6162
rect 20863 5386 20869 6162
rect 20776 5374 20869 5386
rect 21081 6162 21241 6174
rect 21081 5386 21087 6162
rect 21121 5386 21201 6162
rect 21235 5386 21241 6162
rect 21081 5374 21241 5386
rect 21453 6162 21613 6174
rect 21453 5386 21459 6162
rect 21493 5386 21573 6162
rect 21607 5386 21613 6162
rect 21453 5374 21613 5386
rect 21825 6162 21985 6174
rect 21825 5386 21831 6162
rect 21865 5386 21945 6162
rect 21979 5386 21985 6162
rect 21825 5374 21985 5386
rect 22197 6162 22357 6174
rect 22197 5386 22203 6162
rect 22237 5386 22317 6162
rect 22351 5386 22357 6162
rect 22197 5374 22357 5386
rect 22569 6162 22729 6174
rect 22569 5386 22575 6162
rect 22609 5386 22689 6162
rect 22723 5386 22729 6162
rect 22569 5374 22729 5386
rect 22941 6162 23101 6174
rect 22941 5386 22947 6162
rect 22981 5386 23061 6162
rect 23095 5386 23101 6162
rect 22941 5374 23101 5386
rect 23313 6162 23473 6174
rect 23313 5386 23319 6162
rect 23353 5386 23433 6162
rect 23467 5386 23473 6162
rect 23313 5374 23473 5386
rect 23685 6162 23778 6174
rect 23685 5386 23691 6162
rect 23725 5386 23778 6162
rect 23685 5374 23778 5386
rect 20776 5138 20824 5374
rect 20879 5328 21071 5333
rect 20879 5287 20890 5328
rect 20880 5225 20890 5287
rect 20879 5184 20890 5225
rect 21060 5287 21071 5328
rect 21060 5225 21070 5287
rect 21060 5184 21071 5225
rect 20879 5179 21071 5184
rect 21126 5138 21196 5374
rect 21251 5328 21443 5333
rect 21251 5287 21262 5328
rect 21252 5225 21262 5287
rect 21251 5184 21262 5225
rect 21432 5287 21443 5328
rect 21432 5225 21442 5287
rect 21432 5184 21443 5225
rect 21251 5179 21443 5184
rect 21498 5138 21568 5374
rect 21623 5328 21815 5333
rect 21623 5287 21634 5328
rect 21624 5225 21634 5287
rect 21623 5184 21634 5225
rect 21804 5287 21815 5328
rect 21804 5225 21814 5287
rect 21804 5184 21815 5225
rect 21623 5179 21815 5184
rect 21870 5138 21940 5374
rect 21995 5328 22187 5333
rect 21995 5287 22006 5328
rect 21996 5225 22006 5287
rect 21995 5184 22006 5225
rect 22176 5287 22187 5328
rect 22176 5225 22186 5287
rect 22176 5184 22187 5225
rect 21995 5179 22187 5184
rect 22242 5138 22312 5374
rect 22367 5328 22559 5333
rect 22367 5287 22378 5328
rect 22368 5225 22378 5287
rect 22367 5184 22378 5225
rect 22548 5287 22559 5328
rect 22548 5225 22558 5287
rect 22548 5184 22559 5225
rect 22367 5179 22559 5184
rect 22614 5138 22684 5374
rect 22739 5328 22931 5333
rect 22739 5287 22750 5328
rect 22740 5225 22750 5287
rect 22739 5184 22750 5225
rect 22920 5287 22931 5328
rect 22920 5225 22930 5287
rect 22920 5184 22931 5225
rect 22739 5179 22931 5184
rect 22986 5138 23056 5374
rect 23111 5328 23303 5333
rect 23111 5287 23122 5328
rect 23112 5225 23122 5287
rect 23111 5184 23122 5225
rect 23292 5287 23303 5328
rect 23292 5225 23302 5287
rect 23292 5184 23303 5225
rect 23111 5179 23303 5184
rect 23358 5138 23428 5374
rect 23483 5328 23675 5333
rect 23483 5287 23494 5328
rect 23484 5225 23494 5287
rect 23483 5184 23494 5225
rect 23664 5287 23675 5328
rect 23664 5225 23674 5287
rect 23664 5184 23675 5225
rect 23483 5179 23675 5184
rect 23724 5138 23778 5374
rect 20776 5126 20869 5138
rect 20776 4350 20829 5126
rect 20863 4350 20869 5126
rect 20776 4338 20869 4350
rect 21081 5126 21241 5138
rect 21081 4350 21087 5126
rect 21121 4350 21201 5126
rect 21235 4350 21241 5126
rect 21081 4338 21241 4350
rect 21453 5126 21613 5138
rect 21453 4350 21459 5126
rect 21493 4350 21573 5126
rect 21607 4350 21613 5126
rect 21453 4338 21613 4350
rect 21825 5126 21985 5138
rect 21825 4350 21831 5126
rect 21865 4350 21945 5126
rect 21979 4350 21985 5126
rect 21825 4338 21985 4350
rect 22197 5126 22357 5138
rect 22197 4350 22203 5126
rect 22237 4350 22317 5126
rect 22351 4350 22357 5126
rect 22197 4338 22357 4350
rect 22569 5126 22729 5138
rect 22569 4350 22575 5126
rect 22609 4350 22689 5126
rect 22723 4350 22729 5126
rect 22569 4338 22729 4350
rect 22941 5126 23101 5138
rect 22941 4350 22947 5126
rect 22981 4350 23061 5126
rect 23095 4350 23101 5126
rect 22941 4338 23101 4350
rect 23313 5126 23473 5138
rect 23313 4350 23319 5126
rect 23353 4350 23433 5126
rect 23467 4350 23473 5126
rect 23313 4338 23473 4350
rect 23685 5126 23778 5138
rect 23685 4350 23691 5126
rect 23725 4350 23778 5126
rect 23685 4338 23778 4350
rect 20880 4297 20890 4302
rect 20879 4251 20890 4297
rect 21060 4297 21070 4302
rect 20880 4248 20890 4251
rect 21060 4251 21071 4297
rect 21060 4248 21070 4251
rect 21126 3654 21196 4338
rect 21252 4297 21262 4302
rect 21251 4251 21262 4297
rect 21432 4297 21442 4302
rect 21624 4297 21634 4302
rect 21252 4248 21262 4251
rect 21432 4251 21443 4297
rect 21623 4251 21634 4297
rect 21804 4297 21814 4302
rect 21432 4248 21442 4251
rect 21624 4248 21634 4251
rect 21804 4251 21815 4297
rect 21804 4248 21814 4251
rect 21870 3962 21940 4338
rect 21996 4297 22006 4302
rect 21995 4251 22006 4297
rect 22176 4297 22186 4302
rect 22368 4297 22378 4302
rect 21996 4248 22006 4251
rect 22176 4251 22187 4297
rect 22367 4251 22378 4297
rect 22548 4297 22558 4302
rect 22176 4248 22186 4251
rect 22368 4248 22378 4251
rect 22548 4251 22559 4297
rect 22548 4248 22558 4251
rect 22614 3962 22684 4338
rect 22740 4297 22750 4302
rect 22739 4251 22750 4297
rect 22920 4297 22930 4302
rect 23112 4297 23122 4302
rect 22740 4248 22750 4251
rect 22920 4251 22931 4297
rect 23111 4251 23122 4297
rect 23292 4297 23302 4302
rect 22920 4248 22930 4251
rect 23112 4248 23122 4251
rect 23292 4251 23303 4297
rect 23292 4248 23302 4251
rect 21860 3782 21870 3962
rect 22684 3782 22694 3962
rect 20878 3644 21444 3654
rect 20878 3598 20890 3644
rect 20879 3593 20890 3598
rect 20880 3588 20890 3593
rect 21060 3598 21262 3644
rect 21060 3593 21071 3598
rect 21060 3588 21070 3593
rect 20774 3561 20848 3562
rect 21126 3561 21196 3598
rect 21251 3593 21262 3598
rect 21252 3588 21262 3593
rect 21432 3598 21444 3644
rect 21624 3639 21634 3644
rect 21432 3593 21443 3598
rect 21623 3593 21634 3639
rect 21804 3639 21814 3644
rect 21432 3588 21442 3593
rect 21624 3588 21634 3593
rect 21804 3593 21815 3639
rect 21804 3588 21814 3593
rect 21498 3561 21568 3562
rect 21870 3561 21940 3782
rect 21996 3639 22006 3644
rect 21995 3593 22006 3639
rect 22176 3639 22186 3644
rect 22368 3639 22378 3644
rect 21996 3588 22006 3593
rect 22176 3593 22187 3639
rect 22367 3593 22378 3639
rect 22548 3639 22558 3644
rect 22176 3588 22186 3593
rect 22368 3588 22378 3593
rect 22548 3593 22559 3639
rect 22548 3588 22558 3593
rect 22242 3561 22312 3562
rect 22614 3561 22684 3782
rect 23358 3654 23428 4338
rect 23484 4297 23494 4302
rect 23483 4251 23494 4297
rect 23664 4297 23674 4302
rect 23484 4248 23494 4251
rect 23664 4251 23675 4297
rect 23664 4248 23674 4251
rect 27858 4080 28088 8572
rect 24102 3932 29380 4080
rect 23110 3644 23676 3654
rect 22740 3639 22750 3644
rect 22739 3593 22750 3639
rect 22920 3639 22930 3644
rect 22740 3588 22750 3593
rect 22920 3593 22931 3639
rect 23110 3598 23122 3644
rect 23111 3593 23122 3598
rect 22920 3588 22930 3593
rect 23112 3588 23122 3593
rect 23292 3598 23494 3644
rect 23292 3593 23303 3598
rect 23292 3588 23302 3593
rect 22986 3561 23056 3562
rect 23358 3561 23428 3598
rect 23483 3593 23494 3598
rect 23484 3588 23494 3593
rect 23664 3598 23676 3644
rect 23856 3639 23866 3644
rect 23664 3593 23675 3598
rect 23855 3593 23866 3639
rect 24036 3639 24046 3644
rect 23664 3588 23674 3593
rect 23856 3588 23866 3593
rect 24036 3593 24047 3639
rect 24036 3588 24046 3593
rect 23730 3561 23800 3562
rect 24102 3561 24172 3932
rect 24228 3639 24238 3644
rect 24227 3593 24238 3639
rect 24408 3639 24418 3644
rect 24600 3639 24610 3644
rect 24228 3588 24238 3593
rect 24408 3593 24419 3639
rect 24599 3593 24610 3639
rect 24780 3639 24790 3644
rect 24408 3588 24418 3593
rect 24600 3588 24610 3593
rect 24780 3593 24791 3639
rect 24780 3588 24790 3593
rect 24474 3561 24544 3562
rect 24846 3561 24916 3932
rect 24972 3639 24982 3644
rect 24971 3593 24982 3639
rect 25152 3639 25162 3644
rect 25344 3639 25354 3644
rect 24972 3588 24982 3593
rect 25152 3593 25163 3639
rect 25343 3593 25354 3639
rect 25524 3639 25534 3644
rect 25152 3588 25162 3593
rect 25344 3588 25354 3593
rect 25524 3593 25535 3639
rect 25524 3588 25534 3593
rect 25218 3561 25288 3562
rect 25590 3561 25660 3932
rect 25716 3639 25726 3644
rect 25715 3593 25726 3639
rect 25896 3639 25906 3644
rect 26088 3639 26098 3644
rect 25716 3588 25726 3593
rect 25896 3593 25907 3639
rect 26087 3593 26098 3639
rect 26268 3639 26278 3644
rect 25896 3588 25906 3593
rect 26088 3588 26098 3593
rect 26268 3593 26279 3639
rect 26268 3588 26278 3593
rect 25962 3561 26032 3562
rect 26334 3561 26404 3932
rect 26460 3639 26470 3644
rect 26459 3593 26470 3639
rect 26640 3639 26650 3644
rect 26832 3639 26842 3644
rect 26460 3588 26470 3593
rect 26640 3593 26651 3639
rect 26831 3593 26842 3639
rect 27012 3639 27022 3644
rect 26640 3588 26650 3593
rect 26832 3588 26842 3593
rect 27012 3593 27023 3639
rect 27012 3588 27022 3593
rect 26706 3561 26776 3562
rect 27078 3561 27148 3932
rect 27204 3639 27214 3644
rect 27203 3593 27214 3639
rect 27384 3639 27394 3644
rect 27576 3639 27586 3644
rect 27204 3588 27214 3593
rect 27384 3593 27395 3639
rect 27575 3593 27586 3639
rect 27756 3639 27766 3644
rect 27384 3588 27394 3593
rect 27576 3588 27586 3593
rect 27756 3593 27767 3639
rect 27756 3588 27766 3593
rect 27450 3561 27520 3562
rect 27822 3561 27892 3932
rect 27948 3639 27958 3644
rect 27947 3593 27958 3639
rect 28128 3639 28138 3644
rect 28320 3639 28330 3644
rect 27948 3588 27958 3593
rect 28128 3593 28139 3639
rect 28319 3593 28330 3639
rect 28500 3639 28510 3644
rect 28128 3588 28138 3593
rect 28320 3588 28330 3593
rect 28500 3593 28511 3639
rect 28500 3588 28510 3593
rect 28194 3561 28264 3562
rect 28566 3561 28636 3932
rect 28692 3639 28702 3644
rect 28691 3593 28702 3639
rect 28872 3639 28882 3644
rect 29064 3639 29074 3644
rect 28692 3588 28702 3593
rect 28872 3593 28883 3639
rect 29063 3593 29074 3639
rect 29244 3639 29254 3644
rect 28872 3588 28882 3593
rect 29064 3588 29074 3593
rect 29244 3593 29255 3639
rect 29244 3588 29254 3593
rect 28938 3561 29008 3562
rect 29310 3561 29380 3932
rect 29436 3639 29446 3644
rect 29435 3593 29446 3639
rect 29616 3639 29626 3644
rect 29436 3588 29446 3593
rect 29616 3593 29627 3639
rect 29616 3588 29626 3593
rect 29658 3561 29732 3574
rect 20774 3549 20869 3561
rect 20774 3373 20829 3549
rect 20863 3373 20869 3549
rect 20774 3361 20869 3373
rect 21081 3549 21241 3561
rect 21081 3373 21087 3549
rect 21121 3373 21201 3549
rect 21235 3373 21241 3549
rect 21081 3361 21241 3373
rect 21453 3549 21613 3561
rect 21453 3373 21459 3549
rect 21493 3373 21573 3549
rect 21607 3373 21613 3549
rect 21453 3361 21613 3373
rect 21825 3549 21985 3561
rect 21825 3373 21831 3549
rect 21865 3373 21945 3549
rect 21979 3373 21985 3549
rect 21825 3361 21985 3373
rect 22197 3549 22357 3561
rect 22197 3373 22203 3549
rect 22237 3373 22317 3549
rect 22351 3373 22357 3549
rect 22197 3361 22357 3373
rect 22569 3549 22729 3561
rect 22569 3373 22575 3549
rect 22609 3373 22689 3549
rect 22723 3373 22729 3549
rect 22569 3361 22729 3373
rect 22941 3549 23101 3561
rect 22941 3373 22947 3549
rect 22981 3373 23061 3549
rect 23095 3373 23101 3549
rect 22941 3361 23101 3373
rect 23313 3549 23473 3561
rect 23313 3373 23319 3549
rect 23353 3373 23433 3549
rect 23467 3373 23473 3549
rect 23313 3361 23473 3373
rect 23685 3549 23845 3561
rect 23685 3373 23691 3549
rect 23725 3373 23805 3549
rect 23839 3373 23845 3549
rect 23685 3361 23845 3373
rect 24057 3549 24217 3561
rect 24057 3373 24063 3549
rect 24097 3373 24177 3549
rect 24211 3373 24217 3549
rect 24057 3361 24217 3373
rect 24429 3549 24589 3561
rect 24429 3373 24435 3549
rect 24469 3373 24549 3549
rect 24583 3373 24589 3549
rect 24429 3361 24589 3373
rect 24801 3549 24961 3561
rect 24801 3373 24807 3549
rect 24841 3373 24921 3549
rect 24955 3373 24961 3549
rect 24801 3361 24961 3373
rect 25173 3549 25333 3561
rect 25173 3373 25179 3549
rect 25213 3373 25293 3549
rect 25327 3373 25333 3549
rect 25173 3361 25333 3373
rect 25545 3549 25705 3561
rect 25545 3373 25551 3549
rect 25585 3373 25665 3549
rect 25699 3373 25705 3549
rect 25545 3361 25705 3373
rect 25917 3549 26077 3561
rect 25917 3373 25923 3549
rect 25957 3373 26037 3549
rect 26071 3373 26077 3549
rect 25917 3361 26077 3373
rect 26289 3549 26449 3561
rect 26289 3373 26295 3549
rect 26329 3373 26409 3549
rect 26443 3373 26449 3549
rect 26289 3361 26449 3373
rect 26661 3549 26821 3561
rect 26661 3373 26667 3549
rect 26701 3373 26781 3549
rect 26815 3373 26821 3549
rect 26661 3361 26821 3373
rect 27033 3549 27193 3561
rect 27033 3373 27039 3549
rect 27073 3373 27153 3549
rect 27187 3373 27193 3549
rect 27033 3361 27193 3373
rect 27405 3549 27565 3561
rect 27405 3373 27411 3549
rect 27445 3373 27525 3549
rect 27559 3373 27565 3549
rect 27405 3361 27565 3373
rect 27777 3549 27937 3561
rect 27777 3373 27783 3549
rect 27817 3373 27897 3549
rect 27931 3373 27937 3549
rect 27777 3361 27937 3373
rect 28149 3549 28309 3561
rect 28149 3373 28155 3549
rect 28189 3373 28269 3549
rect 28303 3373 28309 3549
rect 28149 3361 28309 3373
rect 28521 3549 28681 3561
rect 28521 3373 28527 3549
rect 28561 3373 28641 3549
rect 28675 3373 28681 3549
rect 28521 3361 28681 3373
rect 28893 3549 29053 3561
rect 28893 3373 28899 3549
rect 28933 3373 29013 3549
rect 29047 3373 29053 3549
rect 28893 3361 29053 3373
rect 29265 3549 29425 3561
rect 29265 3373 29271 3549
rect 29305 3373 29385 3549
rect 29419 3373 29425 3549
rect 29265 3361 29425 3373
rect 29637 3549 29732 3561
rect 29637 3373 29643 3549
rect 29677 3373 29732 3549
rect 29637 3361 29732 3373
rect 20774 3143 20848 3361
rect 21126 3330 21196 3361
rect 20878 3324 21444 3330
rect 20878 3180 20890 3324
rect 21060 3180 21262 3324
rect 21432 3180 21444 3324
rect 20878 3174 21444 3180
rect 21126 3143 21196 3174
rect 21498 3143 21568 3361
rect 21623 3324 21815 3329
rect 21623 3283 21634 3324
rect 21624 3221 21634 3283
rect 21623 3180 21634 3221
rect 21804 3283 21815 3324
rect 21804 3221 21814 3283
rect 21804 3180 21815 3221
rect 21623 3175 21815 3180
rect 21870 3143 21940 3361
rect 21995 3324 22187 3329
rect 21995 3283 22006 3324
rect 21996 3221 22006 3283
rect 21995 3180 22006 3221
rect 22176 3283 22187 3324
rect 22176 3221 22186 3283
rect 22176 3180 22187 3221
rect 21995 3175 22187 3180
rect 22242 3143 22312 3361
rect 22367 3324 22559 3329
rect 22367 3283 22378 3324
rect 22368 3221 22378 3283
rect 22367 3180 22378 3221
rect 22548 3283 22559 3324
rect 22548 3221 22558 3283
rect 22548 3180 22559 3221
rect 22367 3175 22559 3180
rect 22614 3143 22684 3361
rect 22739 3324 22931 3329
rect 22739 3283 22750 3324
rect 22740 3221 22750 3283
rect 22739 3180 22750 3221
rect 22920 3283 22931 3324
rect 22920 3221 22930 3283
rect 22920 3180 22931 3221
rect 22739 3175 22931 3180
rect 22986 3143 23056 3361
rect 23358 3330 23428 3361
rect 23110 3324 23676 3330
rect 23110 3180 23122 3324
rect 23292 3180 23494 3324
rect 23664 3180 23676 3324
rect 23110 3174 23676 3180
rect 23358 3143 23428 3174
rect 23730 3143 23800 3361
rect 23855 3324 24047 3329
rect 23855 3283 23866 3324
rect 23856 3221 23866 3283
rect 23855 3180 23866 3221
rect 24036 3283 24047 3324
rect 24036 3221 24046 3283
rect 24036 3180 24047 3221
rect 23855 3175 24047 3180
rect 24102 3143 24172 3361
rect 24227 3324 24419 3329
rect 24227 3283 24238 3324
rect 24228 3221 24238 3283
rect 24227 3180 24238 3221
rect 24408 3283 24419 3324
rect 24408 3221 24418 3283
rect 24408 3180 24419 3221
rect 24227 3175 24419 3180
rect 24474 3143 24544 3361
rect 24599 3324 24791 3329
rect 24599 3283 24610 3324
rect 24600 3221 24610 3283
rect 24599 3180 24610 3221
rect 24780 3283 24791 3324
rect 24780 3221 24790 3283
rect 24780 3180 24791 3221
rect 24599 3175 24791 3180
rect 24846 3143 24916 3361
rect 24971 3324 25163 3329
rect 24971 3283 24982 3324
rect 24972 3221 24982 3283
rect 24971 3180 24982 3221
rect 25152 3283 25163 3324
rect 25152 3221 25162 3283
rect 25152 3180 25163 3221
rect 24971 3175 25163 3180
rect 25218 3143 25288 3361
rect 25343 3324 25535 3329
rect 25343 3283 25354 3324
rect 25344 3221 25354 3283
rect 25343 3180 25354 3221
rect 25524 3283 25535 3324
rect 25524 3221 25534 3283
rect 25524 3180 25535 3221
rect 25343 3175 25535 3180
rect 25590 3143 25660 3361
rect 25715 3324 25907 3329
rect 25715 3283 25726 3324
rect 25716 3221 25726 3283
rect 25715 3180 25726 3221
rect 25896 3283 25907 3324
rect 25896 3221 25906 3283
rect 25896 3180 25907 3221
rect 25715 3175 25907 3180
rect 25962 3143 26032 3361
rect 26087 3324 26279 3329
rect 26087 3283 26098 3324
rect 26088 3221 26098 3283
rect 26087 3180 26098 3221
rect 26268 3283 26279 3324
rect 26268 3221 26278 3283
rect 26268 3180 26279 3221
rect 26087 3175 26279 3180
rect 26334 3143 26404 3361
rect 26459 3324 26651 3329
rect 26459 3283 26470 3324
rect 26460 3221 26470 3283
rect 26459 3180 26470 3221
rect 26640 3283 26651 3324
rect 26640 3221 26650 3283
rect 26640 3180 26651 3221
rect 26459 3175 26651 3180
rect 26706 3143 26776 3361
rect 26831 3324 27023 3329
rect 26831 3283 26842 3324
rect 26832 3221 26842 3283
rect 26831 3180 26842 3221
rect 27012 3283 27023 3324
rect 27012 3221 27022 3283
rect 27012 3180 27023 3221
rect 26831 3175 27023 3180
rect 27078 3143 27148 3361
rect 27203 3324 27395 3329
rect 27203 3283 27214 3324
rect 27204 3221 27214 3283
rect 27203 3180 27214 3221
rect 27384 3283 27395 3324
rect 27384 3221 27394 3283
rect 27384 3180 27395 3221
rect 27203 3175 27395 3180
rect 27450 3143 27520 3361
rect 27575 3324 27767 3329
rect 27575 3283 27586 3324
rect 27576 3221 27586 3283
rect 27575 3180 27586 3221
rect 27756 3283 27767 3324
rect 27756 3221 27766 3283
rect 27756 3180 27767 3221
rect 27575 3175 27767 3180
rect 27822 3143 27892 3361
rect 27947 3324 28139 3329
rect 27947 3283 27958 3324
rect 27948 3221 27958 3283
rect 27947 3180 27958 3221
rect 28128 3283 28139 3324
rect 28128 3221 28138 3283
rect 28128 3180 28139 3221
rect 27947 3175 28139 3180
rect 28194 3143 28264 3361
rect 28319 3324 28511 3329
rect 28319 3283 28330 3324
rect 28320 3221 28330 3283
rect 28319 3180 28330 3221
rect 28500 3283 28511 3324
rect 28500 3221 28510 3283
rect 28500 3180 28511 3221
rect 28319 3175 28511 3180
rect 28566 3143 28636 3361
rect 28691 3324 28883 3329
rect 28691 3283 28702 3324
rect 28692 3221 28702 3283
rect 28691 3180 28702 3221
rect 28872 3283 28883 3324
rect 28872 3221 28882 3283
rect 28872 3180 28883 3221
rect 28691 3175 28883 3180
rect 28938 3143 29008 3361
rect 29063 3324 29255 3329
rect 29063 3283 29074 3324
rect 29064 3221 29074 3283
rect 29063 3180 29074 3221
rect 29244 3283 29255 3324
rect 29244 3221 29254 3283
rect 29244 3180 29255 3221
rect 29063 3175 29255 3180
rect 29310 3143 29380 3361
rect 29435 3324 29627 3329
rect 29435 3283 29446 3324
rect 29436 3221 29446 3283
rect 29435 3180 29446 3221
rect 29616 3283 29627 3324
rect 29616 3221 29626 3283
rect 29616 3180 29627 3221
rect 29435 3175 29627 3180
rect 29658 3143 29732 3361
rect 20774 3131 20869 3143
rect 20774 2955 20829 3131
rect 20863 2955 20869 3131
rect 20774 2943 20869 2955
rect 21081 3131 21241 3143
rect 21081 2955 21087 3131
rect 21121 2955 21201 3131
rect 21235 2955 21241 3131
rect 21081 2943 21241 2955
rect 21453 3131 21613 3143
rect 21453 2955 21459 3131
rect 21493 2955 21573 3131
rect 21607 2955 21613 3131
rect 21453 2943 21613 2955
rect 21825 3131 21985 3143
rect 21825 2955 21831 3131
rect 21865 2955 21945 3131
rect 21979 2955 21985 3131
rect 21825 2943 21985 2955
rect 22197 3131 22357 3143
rect 22197 2955 22203 3131
rect 22237 2955 22317 3131
rect 22351 2955 22357 3131
rect 22197 2943 22357 2955
rect 22569 3131 22729 3143
rect 22569 2955 22575 3131
rect 22609 2955 22689 3131
rect 22723 2955 22729 3131
rect 22569 2943 22729 2955
rect 22941 3131 23101 3143
rect 22941 2955 22947 3131
rect 22981 2955 23061 3131
rect 23095 2955 23101 3131
rect 22941 2943 23101 2955
rect 23313 3131 23473 3143
rect 23313 2955 23319 3131
rect 23353 2955 23433 3131
rect 23467 2955 23473 3131
rect 23313 2943 23473 2955
rect 23685 3131 23845 3143
rect 23685 2955 23691 3131
rect 23725 2955 23805 3131
rect 23839 2955 23845 3131
rect 23685 2943 23845 2955
rect 24057 3131 24217 3143
rect 24057 2955 24063 3131
rect 24097 2955 24177 3131
rect 24211 2955 24217 3131
rect 24057 2943 24217 2955
rect 24429 3131 24589 3143
rect 24429 2955 24435 3131
rect 24469 2955 24549 3131
rect 24583 2955 24589 3131
rect 24429 2943 24589 2955
rect 24801 3131 24961 3143
rect 24801 2955 24807 3131
rect 24841 2955 24921 3131
rect 24955 2955 24961 3131
rect 24801 2943 24961 2955
rect 25173 3131 25333 3143
rect 25173 2955 25179 3131
rect 25213 2955 25293 3131
rect 25327 2955 25333 3131
rect 25173 2943 25333 2955
rect 25545 3131 25705 3143
rect 25545 2955 25551 3131
rect 25585 2955 25665 3131
rect 25699 2955 25705 3131
rect 25545 2943 25705 2955
rect 25917 3131 26077 3143
rect 25917 2955 25923 3131
rect 25957 2955 26037 3131
rect 26071 2955 26077 3131
rect 25917 2943 26077 2955
rect 26289 3131 26449 3143
rect 26289 2955 26295 3131
rect 26329 2955 26409 3131
rect 26443 2955 26449 3131
rect 26289 2943 26449 2955
rect 26661 3131 26821 3143
rect 26661 2955 26667 3131
rect 26701 2955 26781 3131
rect 26815 2955 26821 3131
rect 26661 2943 26821 2955
rect 27033 3131 27193 3143
rect 27033 2955 27039 3131
rect 27073 2955 27153 3131
rect 27187 2955 27193 3131
rect 27033 2943 27193 2955
rect 27405 3131 27565 3143
rect 27405 2955 27411 3131
rect 27445 2955 27525 3131
rect 27559 2955 27565 3131
rect 27405 2943 27565 2955
rect 27777 3131 27937 3143
rect 27777 2955 27783 3131
rect 27817 2955 27897 3131
rect 27931 2955 27937 3131
rect 27777 2943 27937 2955
rect 28149 3131 28309 3143
rect 28149 2955 28155 3131
rect 28189 2955 28269 3131
rect 28303 2955 28309 3131
rect 28149 2943 28309 2955
rect 28521 3131 28681 3143
rect 28521 2955 28527 3131
rect 28561 2955 28641 3131
rect 28675 2955 28681 3131
rect 28521 2943 28681 2955
rect 28893 3131 29053 3143
rect 28893 2955 28899 3131
rect 28933 2955 29013 3131
rect 29047 2955 29053 3131
rect 28893 2943 29053 2955
rect 29265 3131 29425 3143
rect 29265 2955 29271 3131
rect 29305 2955 29385 3131
rect 29419 2955 29425 3131
rect 29265 2943 29425 2955
rect 29637 3131 29732 3143
rect 29637 2955 29643 3131
rect 29677 2955 29732 3131
rect 29637 2943 29732 2955
rect 20774 2725 20848 2943
rect 21126 2912 21196 2943
rect 20878 2906 21444 2912
rect 20878 2762 20890 2906
rect 21060 2762 21262 2906
rect 21432 2762 21444 2906
rect 20878 2756 21444 2762
rect 21126 2725 21196 2756
rect 21498 2725 21568 2943
rect 21623 2906 21815 2911
rect 21623 2865 21634 2906
rect 21624 2803 21634 2865
rect 21623 2762 21634 2803
rect 21804 2865 21815 2906
rect 21804 2803 21814 2865
rect 21804 2762 21815 2803
rect 21623 2757 21815 2762
rect 21870 2725 21940 2943
rect 21995 2906 22187 2911
rect 21995 2865 22006 2906
rect 21996 2803 22006 2865
rect 21995 2762 22006 2803
rect 22176 2865 22187 2906
rect 22176 2803 22186 2865
rect 22176 2762 22187 2803
rect 21995 2757 22187 2762
rect 22242 2725 22312 2943
rect 22367 2906 22559 2911
rect 22367 2865 22378 2906
rect 22368 2803 22378 2865
rect 22367 2762 22378 2803
rect 22548 2865 22559 2906
rect 22548 2803 22558 2865
rect 22548 2762 22559 2803
rect 22367 2757 22559 2762
rect 22614 2725 22684 2943
rect 22739 2906 22931 2911
rect 22739 2865 22750 2906
rect 22740 2803 22750 2865
rect 22739 2762 22750 2803
rect 22920 2865 22931 2906
rect 22920 2803 22930 2865
rect 22920 2762 22931 2803
rect 22739 2757 22931 2762
rect 22986 2725 23056 2943
rect 23358 2912 23428 2943
rect 23110 2906 23676 2912
rect 23110 2762 23122 2906
rect 23292 2762 23494 2906
rect 23664 2762 23676 2906
rect 23110 2756 23676 2762
rect 23358 2725 23428 2756
rect 23730 2725 23800 2943
rect 23855 2906 24047 2911
rect 23855 2865 23866 2906
rect 23856 2803 23866 2865
rect 23855 2762 23866 2803
rect 24036 2865 24047 2906
rect 24036 2803 24046 2865
rect 24036 2762 24047 2803
rect 23855 2757 24047 2762
rect 24102 2725 24172 2943
rect 24227 2906 24419 2911
rect 24227 2865 24238 2906
rect 24228 2803 24238 2865
rect 24227 2762 24238 2803
rect 24408 2865 24419 2906
rect 24408 2803 24418 2865
rect 24408 2762 24419 2803
rect 24227 2757 24419 2762
rect 24474 2725 24544 2943
rect 24599 2906 24791 2911
rect 24599 2865 24610 2906
rect 24600 2803 24610 2865
rect 24599 2762 24610 2803
rect 24780 2865 24791 2906
rect 24780 2803 24790 2865
rect 24780 2762 24791 2803
rect 24599 2757 24791 2762
rect 24846 2725 24916 2943
rect 24971 2906 25163 2911
rect 24971 2865 24982 2906
rect 24972 2803 24982 2865
rect 24971 2762 24982 2803
rect 25152 2865 25163 2906
rect 25152 2803 25162 2865
rect 25152 2762 25163 2803
rect 24971 2757 25163 2762
rect 25218 2725 25288 2943
rect 25343 2906 25535 2911
rect 25343 2865 25354 2906
rect 25344 2803 25354 2865
rect 25343 2762 25354 2803
rect 25524 2865 25535 2906
rect 25524 2803 25534 2865
rect 25524 2762 25535 2803
rect 25343 2757 25535 2762
rect 25590 2725 25660 2943
rect 25715 2906 25907 2911
rect 25715 2865 25726 2906
rect 25716 2803 25726 2865
rect 25715 2762 25726 2803
rect 25896 2865 25907 2906
rect 25896 2803 25906 2865
rect 25896 2762 25907 2803
rect 25715 2757 25907 2762
rect 25962 2725 26032 2943
rect 26087 2906 26279 2911
rect 26087 2865 26098 2906
rect 26088 2803 26098 2865
rect 26087 2762 26098 2803
rect 26268 2865 26279 2906
rect 26268 2803 26278 2865
rect 26268 2762 26279 2803
rect 26087 2757 26279 2762
rect 26334 2725 26404 2943
rect 26459 2906 26651 2911
rect 26459 2865 26470 2906
rect 26460 2803 26470 2865
rect 26459 2762 26470 2803
rect 26640 2865 26651 2906
rect 26640 2803 26650 2865
rect 26640 2762 26651 2803
rect 26459 2757 26651 2762
rect 26706 2725 26776 2943
rect 26831 2906 27023 2911
rect 26831 2865 26842 2906
rect 26832 2803 26842 2865
rect 26831 2762 26842 2803
rect 27012 2865 27023 2906
rect 27012 2803 27022 2865
rect 27012 2762 27023 2803
rect 26831 2757 27023 2762
rect 27078 2725 27148 2943
rect 27203 2906 27395 2911
rect 27203 2865 27214 2906
rect 27204 2803 27214 2865
rect 27203 2762 27214 2803
rect 27384 2865 27395 2906
rect 27384 2803 27394 2865
rect 27384 2762 27395 2803
rect 27203 2757 27395 2762
rect 27450 2725 27520 2943
rect 27575 2906 27767 2911
rect 27575 2865 27586 2906
rect 27576 2803 27586 2865
rect 27575 2762 27586 2803
rect 27756 2865 27767 2906
rect 27756 2803 27766 2865
rect 27756 2762 27767 2803
rect 27575 2757 27767 2762
rect 27822 2725 27892 2943
rect 27947 2906 28139 2911
rect 27947 2865 27958 2906
rect 27948 2803 27958 2865
rect 27947 2762 27958 2803
rect 28128 2865 28139 2906
rect 28128 2803 28138 2865
rect 28128 2762 28139 2803
rect 27947 2757 28139 2762
rect 28194 2725 28264 2943
rect 28319 2906 28511 2911
rect 28319 2865 28330 2906
rect 28320 2803 28330 2865
rect 28319 2762 28330 2803
rect 28500 2865 28511 2906
rect 28500 2803 28510 2865
rect 28500 2762 28511 2803
rect 28319 2757 28511 2762
rect 28566 2725 28636 2943
rect 28691 2906 28883 2911
rect 28691 2865 28702 2906
rect 28692 2803 28702 2865
rect 28691 2762 28702 2803
rect 28872 2865 28883 2906
rect 28872 2803 28882 2865
rect 28872 2762 28883 2803
rect 28691 2757 28883 2762
rect 28938 2725 29008 2943
rect 29063 2906 29255 2911
rect 29063 2865 29074 2906
rect 29064 2803 29074 2865
rect 29063 2762 29074 2803
rect 29244 2865 29255 2906
rect 29244 2803 29254 2865
rect 29244 2762 29255 2803
rect 29063 2757 29255 2762
rect 29310 2725 29380 2943
rect 29435 2906 29627 2911
rect 29435 2865 29446 2906
rect 29436 2803 29446 2865
rect 29435 2762 29446 2803
rect 29616 2865 29627 2906
rect 29616 2803 29626 2865
rect 29616 2762 29627 2803
rect 29435 2757 29627 2762
rect 29658 2725 29732 2943
rect 20774 2713 20869 2725
rect 20774 2537 20829 2713
rect 20863 2537 20869 2713
rect 20774 2525 20869 2537
rect 21081 2713 21241 2725
rect 21081 2537 21087 2713
rect 21121 2537 21201 2713
rect 21235 2537 21241 2713
rect 21081 2525 21241 2537
rect 21453 2713 21613 2725
rect 21453 2537 21459 2713
rect 21493 2537 21573 2713
rect 21607 2537 21613 2713
rect 21453 2525 21613 2537
rect 21825 2713 21985 2725
rect 21825 2537 21831 2713
rect 21865 2537 21945 2713
rect 21979 2537 21985 2713
rect 21825 2525 21985 2537
rect 22197 2713 22357 2725
rect 22197 2537 22203 2713
rect 22237 2537 22317 2713
rect 22351 2537 22357 2713
rect 22197 2525 22357 2537
rect 22569 2713 22729 2725
rect 22569 2537 22575 2713
rect 22609 2537 22689 2713
rect 22723 2537 22729 2713
rect 22569 2525 22729 2537
rect 22941 2713 23101 2725
rect 22941 2537 22947 2713
rect 22981 2537 23061 2713
rect 23095 2537 23101 2713
rect 22941 2525 23101 2537
rect 23313 2713 23473 2725
rect 23313 2537 23319 2713
rect 23353 2537 23433 2713
rect 23467 2537 23473 2713
rect 23313 2525 23473 2537
rect 23685 2713 23845 2725
rect 23685 2537 23691 2713
rect 23725 2537 23805 2713
rect 23839 2537 23845 2713
rect 23685 2525 23845 2537
rect 24057 2713 24217 2725
rect 24057 2537 24063 2713
rect 24097 2537 24177 2713
rect 24211 2537 24217 2713
rect 24057 2525 24217 2537
rect 24429 2713 24589 2725
rect 24429 2537 24435 2713
rect 24469 2537 24549 2713
rect 24583 2537 24589 2713
rect 24429 2525 24589 2537
rect 24801 2713 24961 2725
rect 24801 2537 24807 2713
rect 24841 2537 24921 2713
rect 24955 2537 24961 2713
rect 24801 2525 24961 2537
rect 25173 2713 25333 2725
rect 25173 2537 25179 2713
rect 25213 2537 25293 2713
rect 25327 2537 25333 2713
rect 25173 2525 25333 2537
rect 25545 2713 25705 2725
rect 25545 2537 25551 2713
rect 25585 2537 25665 2713
rect 25699 2537 25705 2713
rect 25545 2525 25705 2537
rect 25917 2713 26077 2725
rect 25917 2537 25923 2713
rect 25957 2537 26037 2713
rect 26071 2537 26077 2713
rect 25917 2525 26077 2537
rect 26289 2713 26449 2725
rect 26289 2537 26295 2713
rect 26329 2537 26409 2713
rect 26443 2537 26449 2713
rect 26289 2525 26449 2537
rect 26661 2713 26821 2725
rect 26661 2537 26667 2713
rect 26701 2537 26781 2713
rect 26815 2537 26821 2713
rect 26661 2525 26821 2537
rect 27033 2713 27193 2725
rect 27033 2537 27039 2713
rect 27073 2537 27153 2713
rect 27187 2537 27193 2713
rect 27033 2525 27193 2537
rect 27405 2713 27565 2725
rect 27405 2537 27411 2713
rect 27445 2537 27525 2713
rect 27559 2537 27565 2713
rect 27405 2525 27565 2537
rect 27777 2713 27937 2725
rect 27777 2537 27783 2713
rect 27817 2537 27897 2713
rect 27931 2537 27937 2713
rect 27777 2525 27937 2537
rect 28149 2713 28309 2725
rect 28149 2537 28155 2713
rect 28189 2537 28269 2713
rect 28303 2537 28309 2713
rect 28149 2525 28309 2537
rect 28521 2713 28681 2725
rect 28521 2537 28527 2713
rect 28561 2537 28641 2713
rect 28675 2537 28681 2713
rect 28521 2525 28681 2537
rect 28893 2713 29053 2725
rect 28893 2537 28899 2713
rect 28933 2537 29013 2713
rect 29047 2537 29053 2713
rect 28893 2525 29053 2537
rect 29265 2713 29425 2725
rect 29265 2537 29271 2713
rect 29305 2537 29385 2713
rect 29419 2537 29425 2713
rect 29265 2525 29425 2537
rect 29637 2713 29732 2725
rect 29637 2537 29643 2713
rect 29677 2537 29732 2713
rect 29637 2525 29732 2537
rect 20774 2307 20848 2525
rect 21126 2494 21196 2525
rect 20878 2488 21444 2494
rect 20878 2344 20890 2488
rect 21060 2344 21262 2488
rect 21432 2344 21444 2488
rect 20878 2338 21444 2344
rect 21126 2307 21196 2338
rect 21498 2307 21568 2525
rect 21623 2488 21815 2493
rect 21623 2447 21634 2488
rect 21624 2385 21634 2447
rect 21623 2344 21634 2385
rect 21804 2447 21815 2488
rect 21804 2385 21814 2447
rect 21804 2344 21815 2385
rect 21623 2339 21815 2344
rect 21870 2307 21940 2525
rect 21995 2488 22187 2493
rect 21995 2447 22006 2488
rect 21996 2385 22006 2447
rect 21995 2344 22006 2385
rect 22176 2447 22187 2488
rect 22176 2385 22186 2447
rect 22176 2344 22187 2385
rect 21995 2339 22187 2344
rect 22242 2307 22312 2525
rect 22367 2488 22559 2493
rect 22367 2447 22378 2488
rect 22368 2385 22378 2447
rect 22367 2344 22378 2385
rect 22548 2447 22559 2488
rect 22548 2385 22558 2447
rect 22548 2344 22559 2385
rect 22367 2339 22559 2344
rect 22614 2307 22684 2525
rect 22739 2488 22931 2493
rect 22739 2447 22750 2488
rect 22740 2385 22750 2447
rect 22739 2344 22750 2385
rect 22920 2447 22931 2488
rect 22920 2385 22930 2447
rect 22920 2344 22931 2385
rect 22739 2339 22931 2344
rect 22986 2307 23056 2525
rect 23358 2494 23428 2525
rect 23110 2488 23676 2494
rect 23110 2344 23122 2488
rect 23292 2344 23494 2488
rect 23664 2344 23676 2488
rect 23110 2338 23676 2344
rect 23358 2307 23428 2338
rect 23730 2307 23800 2525
rect 23855 2488 24047 2493
rect 23855 2447 23866 2488
rect 23856 2385 23866 2447
rect 23855 2344 23866 2385
rect 24036 2447 24047 2488
rect 24036 2385 24046 2447
rect 24036 2344 24047 2385
rect 23855 2339 24047 2344
rect 24102 2307 24172 2525
rect 24227 2488 24419 2493
rect 24227 2447 24238 2488
rect 24228 2385 24238 2447
rect 24227 2344 24238 2385
rect 24408 2447 24419 2488
rect 24408 2385 24418 2447
rect 24408 2344 24419 2385
rect 24227 2339 24419 2344
rect 24474 2307 24544 2525
rect 24599 2488 24791 2493
rect 24599 2447 24610 2488
rect 24600 2385 24610 2447
rect 24599 2344 24610 2385
rect 24780 2447 24791 2488
rect 24780 2385 24790 2447
rect 24780 2344 24791 2385
rect 24599 2339 24791 2344
rect 24846 2307 24916 2525
rect 24971 2488 25163 2493
rect 24971 2447 24982 2488
rect 24972 2385 24982 2447
rect 24971 2344 24982 2385
rect 25152 2447 25163 2488
rect 25152 2385 25162 2447
rect 25152 2344 25163 2385
rect 24971 2339 25163 2344
rect 25218 2307 25288 2525
rect 25343 2488 25535 2493
rect 25343 2447 25354 2488
rect 25344 2385 25354 2447
rect 25343 2344 25354 2385
rect 25524 2447 25535 2488
rect 25524 2385 25534 2447
rect 25524 2344 25535 2385
rect 25343 2339 25535 2344
rect 25590 2307 25660 2525
rect 25715 2488 25907 2493
rect 25715 2447 25726 2488
rect 25716 2385 25726 2447
rect 25715 2344 25726 2385
rect 25896 2447 25907 2488
rect 25896 2385 25906 2447
rect 25896 2344 25907 2385
rect 25715 2339 25907 2344
rect 25962 2307 26032 2525
rect 26087 2488 26279 2493
rect 26087 2447 26098 2488
rect 26088 2385 26098 2447
rect 26087 2344 26098 2385
rect 26268 2447 26279 2488
rect 26268 2385 26278 2447
rect 26268 2344 26279 2385
rect 26087 2339 26279 2344
rect 26334 2307 26404 2525
rect 26459 2488 26651 2493
rect 26459 2447 26470 2488
rect 26460 2385 26470 2447
rect 26459 2344 26470 2385
rect 26640 2447 26651 2488
rect 26640 2385 26650 2447
rect 26640 2344 26651 2385
rect 26459 2339 26651 2344
rect 26706 2307 26776 2525
rect 26831 2488 27023 2493
rect 26831 2447 26842 2488
rect 26832 2385 26842 2447
rect 26831 2344 26842 2385
rect 27012 2447 27023 2488
rect 27012 2385 27022 2447
rect 27012 2344 27023 2385
rect 26831 2339 27023 2344
rect 27078 2307 27148 2525
rect 27203 2488 27395 2493
rect 27203 2447 27214 2488
rect 27204 2385 27214 2447
rect 27203 2344 27214 2385
rect 27384 2447 27395 2488
rect 27384 2385 27394 2447
rect 27384 2344 27395 2385
rect 27203 2339 27395 2344
rect 27450 2307 27520 2525
rect 27575 2488 27767 2493
rect 27575 2447 27586 2488
rect 27576 2385 27586 2447
rect 27575 2344 27586 2385
rect 27756 2447 27767 2488
rect 27756 2385 27766 2447
rect 27756 2344 27767 2385
rect 27575 2339 27767 2344
rect 27822 2307 27892 2525
rect 27947 2488 28139 2493
rect 27947 2447 27958 2488
rect 27948 2385 27958 2447
rect 27947 2344 27958 2385
rect 28128 2447 28139 2488
rect 28128 2385 28138 2447
rect 28128 2344 28139 2385
rect 27947 2339 28139 2344
rect 28194 2307 28264 2525
rect 28319 2488 28511 2493
rect 28319 2447 28330 2488
rect 28320 2385 28330 2447
rect 28319 2344 28330 2385
rect 28500 2447 28511 2488
rect 28500 2385 28510 2447
rect 28500 2344 28511 2385
rect 28319 2339 28511 2344
rect 28566 2307 28636 2525
rect 28691 2488 28883 2493
rect 28691 2447 28702 2488
rect 28692 2385 28702 2447
rect 28691 2344 28702 2385
rect 28872 2447 28883 2488
rect 28872 2385 28882 2447
rect 28872 2344 28883 2385
rect 28691 2339 28883 2344
rect 28938 2307 29008 2525
rect 29063 2488 29255 2493
rect 29063 2447 29074 2488
rect 29064 2385 29074 2447
rect 29063 2344 29074 2385
rect 29244 2447 29255 2488
rect 29244 2385 29254 2447
rect 29244 2344 29255 2385
rect 29063 2339 29255 2344
rect 29310 2307 29380 2525
rect 29435 2488 29627 2493
rect 29435 2447 29446 2488
rect 29436 2385 29446 2447
rect 29435 2344 29446 2385
rect 29616 2447 29627 2488
rect 29616 2385 29626 2447
rect 29616 2344 29627 2385
rect 29435 2339 29627 2344
rect 29658 2307 29732 2525
rect 20774 2295 20869 2307
rect 20774 2119 20829 2295
rect 20863 2119 20869 2295
rect 20774 2107 20869 2119
rect 21081 2295 21241 2307
rect 21081 2119 21087 2295
rect 21121 2119 21201 2295
rect 21235 2119 21241 2295
rect 21081 2107 21241 2119
rect 21453 2295 21613 2307
rect 21453 2119 21459 2295
rect 21493 2119 21573 2295
rect 21607 2119 21613 2295
rect 21453 2107 21613 2119
rect 21825 2295 21985 2307
rect 21825 2119 21831 2295
rect 21865 2119 21945 2295
rect 21979 2119 21985 2295
rect 21825 2107 21985 2119
rect 22197 2295 22357 2307
rect 22197 2119 22203 2295
rect 22237 2119 22317 2295
rect 22351 2119 22357 2295
rect 22197 2107 22357 2119
rect 22569 2295 22729 2307
rect 22569 2119 22575 2295
rect 22609 2119 22689 2295
rect 22723 2119 22729 2295
rect 22569 2107 22729 2119
rect 22941 2295 23101 2307
rect 22941 2119 22947 2295
rect 22981 2119 23061 2295
rect 23095 2119 23101 2295
rect 22941 2107 23101 2119
rect 23313 2295 23473 2307
rect 23313 2119 23319 2295
rect 23353 2119 23433 2295
rect 23467 2119 23473 2295
rect 23313 2107 23473 2119
rect 23685 2295 23845 2307
rect 23685 2119 23691 2295
rect 23725 2119 23805 2295
rect 23839 2119 23845 2295
rect 23685 2107 23845 2119
rect 24057 2295 24217 2307
rect 24057 2119 24063 2295
rect 24097 2119 24177 2295
rect 24211 2119 24217 2295
rect 24057 2107 24217 2119
rect 24429 2295 24589 2307
rect 24429 2119 24435 2295
rect 24469 2119 24549 2295
rect 24583 2119 24589 2295
rect 24429 2107 24589 2119
rect 24801 2295 24961 2307
rect 24801 2119 24807 2295
rect 24841 2119 24921 2295
rect 24955 2119 24961 2295
rect 24801 2107 24961 2119
rect 25173 2295 25333 2307
rect 25173 2119 25179 2295
rect 25213 2119 25293 2295
rect 25327 2119 25333 2295
rect 25173 2107 25333 2119
rect 25545 2295 25705 2307
rect 25545 2119 25551 2295
rect 25585 2119 25665 2295
rect 25699 2119 25705 2295
rect 25545 2107 25705 2119
rect 25917 2295 26077 2307
rect 25917 2119 25923 2295
rect 25957 2119 26037 2295
rect 26071 2119 26077 2295
rect 25917 2107 26077 2119
rect 26289 2295 26449 2307
rect 26289 2119 26295 2295
rect 26329 2119 26409 2295
rect 26443 2119 26449 2295
rect 26289 2107 26449 2119
rect 26661 2295 26821 2307
rect 26661 2119 26667 2295
rect 26701 2119 26781 2295
rect 26815 2119 26821 2295
rect 26661 2107 26821 2119
rect 27033 2295 27193 2307
rect 27033 2119 27039 2295
rect 27073 2119 27153 2295
rect 27187 2119 27193 2295
rect 27033 2107 27193 2119
rect 27405 2295 27565 2307
rect 27405 2119 27411 2295
rect 27445 2119 27525 2295
rect 27559 2119 27565 2295
rect 27405 2107 27565 2119
rect 27777 2295 27937 2307
rect 27777 2119 27783 2295
rect 27817 2119 27897 2295
rect 27931 2119 27937 2295
rect 27777 2107 27937 2119
rect 28149 2295 28309 2307
rect 28149 2119 28155 2295
rect 28189 2119 28269 2295
rect 28303 2119 28309 2295
rect 28149 2107 28309 2119
rect 28521 2295 28681 2307
rect 28521 2119 28527 2295
rect 28561 2119 28641 2295
rect 28675 2119 28681 2295
rect 28521 2107 28681 2119
rect 28893 2295 29053 2307
rect 28893 2119 28899 2295
rect 28933 2119 29013 2295
rect 29047 2119 29053 2295
rect 28893 2107 29053 2119
rect 29265 2295 29425 2307
rect 29265 2119 29271 2295
rect 29305 2119 29385 2295
rect 29419 2119 29425 2295
rect 29265 2107 29425 2119
rect 29637 2295 29732 2307
rect 29637 2119 29643 2295
rect 29677 2119 29732 2295
rect 29637 2107 29732 2119
rect 20774 1984 20848 2107
rect 20880 2075 20890 2080
rect 20879 2070 20890 2075
rect 20878 2024 20890 2070
rect 21060 2075 21070 2080
rect 21060 2070 21071 2075
rect 21126 2070 21196 2107
rect 21498 2106 21568 2107
rect 21870 2106 21940 2107
rect 22242 2106 22312 2107
rect 22614 2106 22684 2107
rect 22986 2106 23056 2107
rect 21252 2075 21262 2080
rect 21251 2070 21262 2075
rect 21060 2024 21262 2070
rect 21432 2075 21442 2080
rect 21432 2070 21443 2075
rect 21432 2024 21444 2070
rect 20878 2012 21444 2024
rect 21504 1992 21562 2106
rect 21624 2075 21634 2080
rect 21623 2029 21634 2075
rect 21804 2075 21814 2080
rect 21996 2075 22006 2080
rect 21624 2024 21634 2029
rect 21804 2029 21815 2075
rect 21995 2029 22006 2075
rect 22176 2075 22186 2080
rect 21804 2024 21814 2029
rect 21996 2024 22006 2029
rect 22176 2029 22187 2075
rect 22176 2024 22186 2029
rect 22248 1992 22306 2106
rect 22368 2075 22378 2080
rect 22367 2029 22378 2075
rect 22548 2075 22558 2080
rect 22740 2075 22750 2080
rect 22368 2024 22378 2029
rect 22548 2029 22559 2075
rect 22739 2029 22750 2075
rect 22920 2075 22930 2080
rect 22548 2024 22558 2029
rect 22740 2024 22750 2029
rect 22920 2029 22931 2075
rect 22920 2024 22930 2029
rect 22992 1992 23050 2106
rect 23112 2075 23122 2080
rect 23111 2070 23122 2075
rect 23110 2024 23122 2070
rect 23292 2075 23302 2080
rect 23292 2070 23303 2075
rect 23358 2070 23428 2107
rect 23730 2106 23800 2107
rect 24102 2106 24172 2107
rect 24474 2106 24544 2107
rect 24846 2106 24916 2107
rect 25218 2106 25288 2107
rect 25590 2106 25660 2107
rect 25962 2106 26032 2107
rect 26334 2106 26404 2107
rect 26706 2106 26776 2107
rect 27078 2106 27148 2107
rect 27450 2106 27520 2107
rect 27822 2106 27892 2107
rect 28194 2106 28264 2107
rect 28566 2106 28636 2107
rect 28938 2106 29008 2107
rect 29310 2106 29380 2107
rect 23484 2075 23494 2080
rect 23483 2070 23494 2075
rect 23292 2024 23494 2070
rect 23664 2075 23674 2080
rect 23664 2070 23675 2075
rect 23664 2024 23676 2070
rect 23110 2012 23676 2024
rect 23736 1992 23794 2106
rect 23856 2075 23866 2080
rect 23855 2029 23866 2075
rect 24036 2075 24046 2080
rect 24228 2075 24238 2080
rect 23856 2024 23866 2029
rect 24036 2029 24047 2075
rect 24227 2029 24238 2075
rect 24408 2075 24418 2080
rect 24036 2024 24046 2029
rect 24228 2024 24238 2029
rect 24408 2029 24419 2075
rect 24408 2024 24418 2029
rect 24480 1992 24538 2106
rect 24600 2075 24610 2080
rect 24599 2029 24610 2075
rect 24780 2075 24790 2080
rect 24972 2075 24982 2080
rect 24600 2024 24610 2029
rect 24780 2029 24791 2075
rect 24971 2029 24982 2075
rect 25152 2075 25162 2080
rect 24780 2024 24790 2029
rect 24972 2024 24982 2029
rect 25152 2029 25163 2075
rect 25152 2024 25162 2029
rect 25224 1992 25282 2106
rect 25344 2075 25354 2080
rect 25343 2029 25354 2075
rect 25524 2075 25534 2080
rect 25716 2075 25726 2080
rect 25344 2024 25354 2029
rect 25524 2029 25535 2075
rect 25715 2029 25726 2075
rect 25896 2075 25906 2080
rect 25524 2024 25534 2029
rect 25716 2024 25726 2029
rect 25896 2029 25907 2075
rect 25896 2024 25906 2029
rect 25968 1992 26026 2106
rect 26088 2075 26098 2080
rect 26087 2029 26098 2075
rect 26268 2075 26278 2080
rect 26460 2075 26470 2080
rect 26088 2024 26098 2029
rect 26268 2029 26279 2075
rect 26459 2029 26470 2075
rect 26640 2075 26650 2080
rect 26268 2024 26278 2029
rect 26460 2024 26470 2029
rect 26640 2029 26651 2075
rect 26640 2024 26650 2029
rect 26712 1992 26770 2106
rect 26832 2075 26842 2080
rect 26831 2029 26842 2075
rect 27012 2075 27022 2080
rect 27204 2075 27214 2080
rect 26832 2024 26842 2029
rect 27012 2029 27023 2075
rect 27203 2029 27214 2075
rect 27384 2075 27394 2080
rect 27012 2024 27022 2029
rect 27204 2024 27214 2029
rect 27384 2029 27395 2075
rect 27384 2024 27394 2029
rect 27456 1992 27514 2106
rect 27576 2075 27586 2080
rect 27575 2029 27586 2075
rect 27756 2075 27766 2080
rect 27948 2075 27958 2080
rect 27576 2024 27586 2029
rect 27756 2029 27767 2075
rect 27947 2029 27958 2075
rect 28128 2075 28138 2080
rect 27756 2024 27766 2029
rect 27948 2024 27958 2029
rect 28128 2029 28139 2075
rect 28128 2024 28138 2029
rect 28200 1992 28258 2106
rect 28320 2075 28330 2080
rect 28319 2029 28330 2075
rect 28500 2075 28510 2080
rect 28692 2075 28702 2080
rect 28320 2024 28330 2029
rect 28500 2029 28511 2075
rect 28691 2029 28702 2075
rect 28872 2075 28882 2080
rect 28500 2024 28510 2029
rect 28692 2024 28702 2029
rect 28872 2029 28883 2075
rect 28872 2024 28882 2029
rect 28944 1992 29002 2106
rect 29064 2075 29074 2080
rect 29063 2029 29074 2075
rect 29244 2075 29254 2080
rect 29436 2075 29446 2080
rect 29064 2024 29074 2029
rect 29244 2029 29255 2075
rect 29435 2029 29446 2075
rect 29616 2075 29626 2080
rect 29244 2024 29254 2029
rect 29436 2024 29446 2029
rect 29616 2029 29627 2075
rect 29616 2024 29626 2029
rect 21486 1986 21580 1992
rect 20774 1978 20912 1984
rect 20774 1908 20830 1978
rect 20900 1908 20912 1978
rect 21486 1916 21498 1986
rect 21568 1916 21580 1986
rect 21486 1910 21580 1916
rect 22230 1986 22324 1992
rect 22230 1916 22242 1986
rect 22312 1916 22324 1986
rect 22230 1910 22324 1916
rect 22974 1986 23068 1992
rect 22974 1916 22986 1986
rect 23056 1916 23068 1986
rect 22974 1910 23068 1916
rect 23718 1986 23812 1992
rect 23718 1916 23730 1986
rect 23800 1916 23812 1986
rect 23718 1910 23812 1916
rect 24462 1986 24556 1992
rect 24462 1916 24474 1986
rect 24544 1916 24556 1986
rect 24462 1910 24556 1916
rect 25206 1986 25300 1992
rect 25206 1916 25218 1986
rect 25288 1916 25300 1986
rect 25206 1910 25300 1916
rect 25950 1986 26044 1992
rect 25950 1916 25962 1986
rect 26032 1916 26044 1986
rect 25950 1910 26044 1916
rect 26694 1986 26788 1992
rect 26694 1916 26706 1986
rect 26776 1916 26788 1986
rect 26694 1910 26788 1916
rect 27438 1986 27532 1992
rect 27438 1916 27450 1986
rect 27520 1916 27532 1986
rect 27438 1910 27532 1916
rect 28182 1986 28276 1992
rect 28182 1916 28194 1986
rect 28264 1916 28276 1986
rect 28182 1910 28276 1916
rect 28926 1986 29020 1992
rect 29658 1988 29732 2107
rect 28926 1916 28938 1986
rect 29008 1916 29020 1986
rect 28926 1910 29020 1916
rect 29588 1982 29732 1988
rect 29588 1912 29600 1982
rect 29670 1912 29732 1982
rect 20774 1902 20912 1908
rect 20774 1870 20848 1902
rect 21504 1870 21562 1910
rect 22248 1870 22306 1910
rect 22992 1870 23050 1910
rect 23736 1870 23794 1910
rect 24480 1870 24538 1910
rect 25224 1870 25282 1910
rect 25968 1870 26026 1910
rect 26712 1870 26770 1910
rect 27456 1870 27514 1910
rect 28200 1870 28258 1910
rect 28944 1870 29002 1910
rect 29588 1906 29732 1912
rect 29658 1882 29732 1906
rect 29658 1870 29746 1882
rect 20700 1670 20710 1870
rect 20910 1670 20920 1870
rect 21424 1670 21434 1870
rect 21634 1670 21644 1870
rect 22168 1670 22178 1870
rect 22378 1670 22388 1870
rect 22912 1670 22922 1870
rect 23122 1670 23132 1870
rect 23656 1670 23666 1870
rect 23866 1670 23876 1870
rect 24400 1670 24410 1870
rect 24610 1670 24620 1870
rect 25144 1670 25154 1870
rect 25354 1670 25364 1870
rect 25888 1670 25898 1870
rect 26098 1670 26108 1870
rect 26632 1670 26642 1870
rect 26842 1670 26852 1870
rect 27376 1670 27386 1870
rect 27586 1670 27596 1870
rect 28120 1670 28130 1870
rect 28330 1670 28340 1870
rect 28864 1670 28874 1870
rect 29074 1670 29084 1870
rect 29608 1670 29618 1870
rect 29818 1670 29828 1870
<< via1 >>
rect 19572 10916 19772 11116
rect 20316 10916 20516 11116
rect 21060 10916 21260 11116
rect 21804 10916 22004 11116
rect 22548 10916 22748 11116
rect 23292 10916 23492 11116
rect 24036 10916 24236 11116
rect 24780 10916 24980 11116
rect 25152 10916 25352 11116
rect 25896 10916 26096 11116
rect 26640 10916 26840 11116
rect 27384 10916 27584 11116
rect 28128 10916 28328 11116
rect 28872 10916 29072 11116
rect 29616 10916 29816 11116
rect 30360 10916 30560 11116
rect 31104 10916 31304 11116
rect 19402 10715 19572 10728
rect 19402 10681 19403 10715
rect 19403 10681 19571 10715
rect 19571 10681 19572 10715
rect 19402 10668 19572 10681
rect 19774 10715 19944 10728
rect 19774 10681 19775 10715
rect 19775 10681 19943 10715
rect 19943 10681 19944 10715
rect 19774 10668 19944 10681
rect 20146 10715 20316 10728
rect 20146 10681 20147 10715
rect 20147 10681 20315 10715
rect 20315 10681 20316 10715
rect 20146 10668 20316 10681
rect 20518 10715 20688 10728
rect 20518 10681 20519 10715
rect 20519 10681 20687 10715
rect 20687 10681 20688 10715
rect 20518 10668 20688 10681
rect 20890 10715 21060 10728
rect 20890 10681 20891 10715
rect 20891 10681 21059 10715
rect 21059 10681 21060 10715
rect 20890 10668 21060 10681
rect 21262 10715 21432 10728
rect 21262 10681 21263 10715
rect 21263 10681 21431 10715
rect 21431 10681 21432 10715
rect 21262 10668 21432 10681
rect 21634 10715 21804 10728
rect 21634 10681 21635 10715
rect 21635 10681 21803 10715
rect 21803 10681 21804 10715
rect 21634 10668 21804 10681
rect 22006 10715 22176 10728
rect 22006 10681 22007 10715
rect 22007 10681 22175 10715
rect 22175 10681 22176 10715
rect 22006 10668 22176 10681
rect 22378 10715 22548 10728
rect 22378 10681 22379 10715
rect 22379 10681 22547 10715
rect 22547 10681 22548 10715
rect 22378 10668 22548 10681
rect 22750 10715 22920 10728
rect 22750 10681 22751 10715
rect 22751 10681 22919 10715
rect 22919 10681 22920 10715
rect 22750 10668 22920 10681
rect 23122 10715 23292 10728
rect 23122 10681 23123 10715
rect 23123 10681 23291 10715
rect 23291 10681 23292 10715
rect 23122 10668 23292 10681
rect 23494 10715 23664 10728
rect 23494 10681 23495 10715
rect 23495 10681 23663 10715
rect 23663 10681 23664 10715
rect 23494 10668 23664 10681
rect 23866 10715 24036 10728
rect 23866 10681 23867 10715
rect 23867 10681 24035 10715
rect 24035 10681 24036 10715
rect 23866 10668 24036 10681
rect 24238 10715 24408 10728
rect 24238 10681 24239 10715
rect 24239 10681 24407 10715
rect 24407 10681 24408 10715
rect 24238 10668 24408 10681
rect 24610 10715 24780 10728
rect 24610 10681 24611 10715
rect 24611 10681 24779 10715
rect 24779 10681 24780 10715
rect 24610 10668 24780 10681
rect 24982 10715 25152 10728
rect 24982 10681 24983 10715
rect 24983 10681 25151 10715
rect 25151 10681 25152 10715
rect 24982 10668 25152 10681
rect 19402 10187 19572 10188
rect 19402 10153 19403 10187
rect 19403 10153 19571 10187
rect 19571 10153 19572 10187
rect 19402 10079 19572 10153
rect 19402 10045 19403 10079
rect 19403 10045 19571 10079
rect 19571 10045 19572 10079
rect 19402 10044 19572 10045
rect 19774 10187 19944 10188
rect 19774 10153 19775 10187
rect 19775 10153 19943 10187
rect 19943 10153 19944 10187
rect 19774 10079 19944 10153
rect 19774 10045 19775 10079
rect 19775 10045 19943 10079
rect 19943 10045 19944 10079
rect 19774 10044 19944 10045
rect 20146 10187 20316 10188
rect 20146 10153 20147 10187
rect 20147 10153 20315 10187
rect 20315 10153 20316 10187
rect 20146 10079 20316 10153
rect 20146 10045 20147 10079
rect 20147 10045 20315 10079
rect 20315 10045 20316 10079
rect 20146 10044 20316 10045
rect 20518 10187 20688 10188
rect 20518 10153 20519 10187
rect 20519 10153 20687 10187
rect 20687 10153 20688 10187
rect 20518 10079 20688 10153
rect 20518 10045 20519 10079
rect 20519 10045 20687 10079
rect 20687 10045 20688 10079
rect 20518 10044 20688 10045
rect 20890 10187 21060 10188
rect 20890 10153 20891 10187
rect 20891 10153 21059 10187
rect 21059 10153 21060 10187
rect 20890 10079 21060 10153
rect 20890 10045 20891 10079
rect 20891 10045 21059 10079
rect 21059 10045 21060 10079
rect 20890 10044 21060 10045
rect 21262 10187 21432 10188
rect 21262 10153 21263 10187
rect 21263 10153 21431 10187
rect 21431 10153 21432 10187
rect 21262 10079 21432 10153
rect 21262 10045 21263 10079
rect 21263 10045 21431 10079
rect 21431 10045 21432 10079
rect 21262 10044 21432 10045
rect 21634 10187 21804 10188
rect 21634 10153 21635 10187
rect 21635 10153 21803 10187
rect 21803 10153 21804 10187
rect 21634 10079 21804 10153
rect 21634 10045 21635 10079
rect 21635 10045 21803 10079
rect 21803 10045 21804 10079
rect 21634 10044 21804 10045
rect 22006 10187 22176 10188
rect 22006 10153 22007 10187
rect 22007 10153 22175 10187
rect 22175 10153 22176 10187
rect 22006 10079 22176 10153
rect 22006 10045 22007 10079
rect 22007 10045 22175 10079
rect 22175 10045 22176 10079
rect 22006 10044 22176 10045
rect 22378 10187 22548 10188
rect 22378 10153 22379 10187
rect 22379 10153 22547 10187
rect 22547 10153 22548 10187
rect 22378 10079 22548 10153
rect 22378 10045 22379 10079
rect 22379 10045 22547 10079
rect 22547 10045 22548 10079
rect 22378 10044 22548 10045
rect 22750 10187 22920 10188
rect 22750 10153 22751 10187
rect 22751 10153 22919 10187
rect 22919 10153 22920 10187
rect 22750 10079 22920 10153
rect 22750 10045 22751 10079
rect 22751 10045 22919 10079
rect 22919 10045 22920 10079
rect 22750 10044 22920 10045
rect 23122 10187 23292 10188
rect 23122 10153 23123 10187
rect 23123 10153 23291 10187
rect 23291 10153 23292 10187
rect 23122 10079 23292 10153
rect 23122 10045 23123 10079
rect 23123 10045 23291 10079
rect 23291 10045 23292 10079
rect 23122 10044 23292 10045
rect 23494 10187 23664 10188
rect 23494 10153 23495 10187
rect 23495 10153 23663 10187
rect 23663 10153 23664 10187
rect 23494 10079 23664 10153
rect 23494 10045 23495 10079
rect 23495 10045 23663 10079
rect 23663 10045 23664 10079
rect 23494 10044 23664 10045
rect 23866 10187 24036 10188
rect 23866 10153 23867 10187
rect 23867 10153 24035 10187
rect 24035 10153 24036 10187
rect 23866 10079 24036 10153
rect 23866 10045 23867 10079
rect 23867 10045 24035 10079
rect 24035 10045 24036 10079
rect 23866 10044 24036 10045
rect 24238 10187 24408 10188
rect 24238 10153 24239 10187
rect 24239 10153 24407 10187
rect 24407 10153 24408 10187
rect 24238 10079 24408 10153
rect 24238 10045 24239 10079
rect 24239 10045 24407 10079
rect 24407 10045 24408 10079
rect 24238 10044 24408 10045
rect 24610 10187 24780 10188
rect 24610 10153 24611 10187
rect 24611 10153 24779 10187
rect 24779 10153 24780 10187
rect 24610 10079 24780 10153
rect 24610 10045 24611 10079
rect 24611 10045 24779 10079
rect 24779 10045 24780 10079
rect 24610 10044 24780 10045
rect 24982 10187 25152 10188
rect 24982 10153 24983 10187
rect 24983 10153 25151 10187
rect 25151 10153 25152 10187
rect 24982 10079 25152 10153
rect 24982 10045 24983 10079
rect 24983 10045 25151 10079
rect 25151 10045 25152 10079
rect 24982 10044 25152 10045
rect 19402 9551 19572 9552
rect 19402 9517 19403 9551
rect 19403 9517 19571 9551
rect 19571 9517 19572 9551
rect 19402 9443 19572 9517
rect 19402 9409 19403 9443
rect 19403 9409 19571 9443
rect 19571 9409 19572 9443
rect 19402 9408 19572 9409
rect 19774 9551 19944 9552
rect 19774 9517 19775 9551
rect 19775 9517 19943 9551
rect 19943 9517 19944 9551
rect 19774 9443 19944 9517
rect 19774 9409 19775 9443
rect 19775 9409 19943 9443
rect 19943 9409 19944 9443
rect 19774 9408 19944 9409
rect 20146 9551 20316 9552
rect 20146 9517 20147 9551
rect 20147 9517 20315 9551
rect 20315 9517 20316 9551
rect 20146 9443 20316 9517
rect 20146 9409 20147 9443
rect 20147 9409 20315 9443
rect 20315 9409 20316 9443
rect 20146 9408 20316 9409
rect 20518 9551 20688 9552
rect 20518 9517 20519 9551
rect 20519 9517 20687 9551
rect 20687 9517 20688 9551
rect 20518 9443 20688 9517
rect 20518 9409 20519 9443
rect 20519 9409 20687 9443
rect 20687 9409 20688 9443
rect 20518 9408 20688 9409
rect 20890 9551 21060 9552
rect 20890 9517 20891 9551
rect 20891 9517 21059 9551
rect 21059 9517 21060 9551
rect 20890 9443 21060 9517
rect 20890 9409 20891 9443
rect 20891 9409 21059 9443
rect 21059 9409 21060 9443
rect 20890 9408 21060 9409
rect 21262 9551 21432 9552
rect 21262 9517 21263 9551
rect 21263 9517 21431 9551
rect 21431 9517 21432 9551
rect 21262 9443 21432 9517
rect 21262 9409 21263 9443
rect 21263 9409 21431 9443
rect 21431 9409 21432 9443
rect 21262 9408 21432 9409
rect 21634 9551 21804 9552
rect 21634 9517 21635 9551
rect 21635 9517 21803 9551
rect 21803 9517 21804 9551
rect 21634 9443 21804 9517
rect 21634 9409 21635 9443
rect 21635 9409 21803 9443
rect 21803 9409 21804 9443
rect 21634 9408 21804 9409
rect 22006 9551 22176 9552
rect 22006 9517 22007 9551
rect 22007 9517 22175 9551
rect 22175 9517 22176 9551
rect 22006 9443 22176 9517
rect 22006 9409 22007 9443
rect 22007 9409 22175 9443
rect 22175 9409 22176 9443
rect 22006 9408 22176 9409
rect 22378 9551 22548 9552
rect 22378 9517 22379 9551
rect 22379 9517 22547 9551
rect 22547 9517 22548 9551
rect 22378 9443 22548 9517
rect 22378 9409 22379 9443
rect 22379 9409 22547 9443
rect 22547 9409 22548 9443
rect 22378 9408 22548 9409
rect 22750 9551 22920 9552
rect 22750 9517 22751 9551
rect 22751 9517 22919 9551
rect 22919 9517 22920 9551
rect 22750 9443 22920 9517
rect 22750 9409 22751 9443
rect 22751 9409 22919 9443
rect 22919 9409 22920 9443
rect 22750 9408 22920 9409
rect 23122 9551 23292 9552
rect 23122 9517 23123 9551
rect 23123 9517 23291 9551
rect 23291 9517 23292 9551
rect 23122 9443 23292 9517
rect 23122 9409 23123 9443
rect 23123 9409 23291 9443
rect 23291 9409 23292 9443
rect 23122 9408 23292 9409
rect 23494 9551 23664 9552
rect 23494 9517 23495 9551
rect 23495 9517 23663 9551
rect 23663 9517 23664 9551
rect 23494 9443 23664 9517
rect 23494 9409 23495 9443
rect 23495 9409 23663 9443
rect 23663 9409 23664 9443
rect 23494 9408 23664 9409
rect 23866 9551 24036 9552
rect 23866 9517 23867 9551
rect 23867 9517 24035 9551
rect 24035 9517 24036 9551
rect 23866 9443 24036 9517
rect 23866 9409 23867 9443
rect 23867 9409 24035 9443
rect 24035 9409 24036 9443
rect 23866 9408 24036 9409
rect 24238 9551 24408 9552
rect 24238 9517 24239 9551
rect 24239 9517 24407 9551
rect 24407 9517 24408 9551
rect 24238 9443 24408 9517
rect 24238 9409 24239 9443
rect 24239 9409 24407 9443
rect 24407 9409 24408 9443
rect 24238 9408 24408 9409
rect 24610 9551 24780 9552
rect 24610 9517 24611 9551
rect 24611 9517 24779 9551
rect 24779 9517 24780 9551
rect 24610 9443 24780 9517
rect 24610 9409 24611 9443
rect 24611 9409 24779 9443
rect 24779 9409 24780 9443
rect 24610 9408 24780 9409
rect 24982 9551 25152 9552
rect 24982 9517 24983 9551
rect 24983 9517 25151 9551
rect 25151 9517 25152 9551
rect 24982 9443 25152 9517
rect 24982 9409 24983 9443
rect 24983 9409 25151 9443
rect 25151 9409 25152 9443
rect 24982 9408 25152 9409
rect 19402 8915 19572 8928
rect 19402 8881 19403 8915
rect 19403 8881 19571 8915
rect 19571 8881 19572 8915
rect 19402 8868 19572 8881
rect 19774 8915 19944 8928
rect 19774 8881 19775 8915
rect 19775 8881 19943 8915
rect 19943 8881 19944 8915
rect 19774 8868 19944 8881
rect 20146 8915 20316 8928
rect 20146 8881 20147 8915
rect 20147 8881 20315 8915
rect 20315 8881 20316 8915
rect 20146 8868 20316 8881
rect 20518 8915 20688 8928
rect 20518 8881 20519 8915
rect 20519 8881 20687 8915
rect 20687 8881 20688 8915
rect 20518 8868 20688 8881
rect 20890 8915 21060 8928
rect 20890 8881 20891 8915
rect 20891 8881 21059 8915
rect 21059 8881 21060 8915
rect 20890 8868 21060 8881
rect 21262 8915 21432 8928
rect 21262 8881 21263 8915
rect 21263 8881 21431 8915
rect 21431 8881 21432 8915
rect 21262 8868 21432 8881
rect 21634 8915 21804 8928
rect 21634 8881 21635 8915
rect 21635 8881 21803 8915
rect 21803 8881 21804 8915
rect 21634 8868 21804 8881
rect 22006 8915 22176 8928
rect 22006 8881 22007 8915
rect 22007 8881 22175 8915
rect 22175 8881 22176 8915
rect 22006 8868 22176 8881
rect 22378 8915 22548 8928
rect 22378 8881 22379 8915
rect 22379 8881 22547 8915
rect 22547 8881 22548 8915
rect 22378 8868 22548 8881
rect 22750 8915 22920 8928
rect 22750 8881 22751 8915
rect 22751 8881 22919 8915
rect 22919 8881 22920 8915
rect 22750 8868 22920 8881
rect 23122 8915 23292 8928
rect 23122 8881 23123 8915
rect 23123 8881 23291 8915
rect 23291 8881 23292 8915
rect 23122 8868 23292 8881
rect 23494 8915 23664 8928
rect 23494 8881 23495 8915
rect 23495 8881 23663 8915
rect 23663 8881 23664 8915
rect 23494 8868 23664 8881
rect 23866 8915 24036 8928
rect 23866 8881 23867 8915
rect 23867 8881 24035 8915
rect 24035 8881 24036 8915
rect 23866 8868 24036 8881
rect 24238 8915 24408 8928
rect 24238 8881 24239 8915
rect 24239 8881 24407 8915
rect 24407 8881 24408 8915
rect 24238 8868 24408 8881
rect 25354 10715 25524 10728
rect 25354 10681 25355 10715
rect 25355 10681 25523 10715
rect 25523 10681 25524 10715
rect 25354 10668 25524 10681
rect 25726 10715 25896 10728
rect 25726 10681 25727 10715
rect 25727 10681 25895 10715
rect 25895 10681 25896 10715
rect 25726 10668 25896 10681
rect 26098 10715 26268 10728
rect 26098 10681 26099 10715
rect 26099 10681 26267 10715
rect 26267 10681 26268 10715
rect 26098 10668 26268 10681
rect 26470 10715 26640 10728
rect 26470 10681 26471 10715
rect 26471 10681 26639 10715
rect 26639 10681 26640 10715
rect 26470 10668 26640 10681
rect 26842 10715 27012 10728
rect 26842 10681 26843 10715
rect 26843 10681 27011 10715
rect 27011 10681 27012 10715
rect 26842 10668 27012 10681
rect 27214 10715 27384 10728
rect 27214 10681 27215 10715
rect 27215 10681 27383 10715
rect 27383 10681 27384 10715
rect 27214 10668 27384 10681
rect 27586 10715 27756 10728
rect 27586 10681 27587 10715
rect 27587 10681 27755 10715
rect 27755 10681 27756 10715
rect 27586 10668 27756 10681
rect 27958 10715 28128 10728
rect 27958 10681 27959 10715
rect 27959 10681 28127 10715
rect 28127 10681 28128 10715
rect 27958 10668 28128 10681
rect 28330 10715 28500 10728
rect 28330 10681 28331 10715
rect 28331 10681 28499 10715
rect 28499 10681 28500 10715
rect 28330 10668 28500 10681
rect 28702 10715 28872 10728
rect 28702 10681 28703 10715
rect 28703 10681 28871 10715
rect 28871 10681 28872 10715
rect 28702 10668 28872 10681
rect 29074 10715 29244 10728
rect 29074 10681 29075 10715
rect 29075 10681 29243 10715
rect 29243 10681 29244 10715
rect 29074 10668 29244 10681
rect 29446 10715 29616 10728
rect 29446 10681 29447 10715
rect 29447 10681 29615 10715
rect 29615 10681 29616 10715
rect 29446 10668 29616 10681
rect 29818 10715 29988 10728
rect 29818 10681 29819 10715
rect 29819 10681 29987 10715
rect 29987 10681 29988 10715
rect 29818 10668 29988 10681
rect 30190 10715 30360 10728
rect 30190 10681 30191 10715
rect 30191 10681 30359 10715
rect 30359 10681 30360 10715
rect 30190 10668 30360 10681
rect 30562 10715 30732 10728
rect 30562 10681 30563 10715
rect 30563 10681 30731 10715
rect 30731 10681 30732 10715
rect 30562 10668 30732 10681
rect 30934 10715 31104 10728
rect 30934 10681 30935 10715
rect 30935 10681 31103 10715
rect 31103 10681 31104 10715
rect 30934 10668 31104 10681
rect 25354 10187 25524 10188
rect 25354 10153 25355 10187
rect 25355 10153 25523 10187
rect 25523 10153 25524 10187
rect 25354 10079 25524 10153
rect 25354 10045 25355 10079
rect 25355 10045 25523 10079
rect 25523 10045 25524 10079
rect 25354 10044 25524 10045
rect 25726 10187 25896 10188
rect 25726 10153 25727 10187
rect 25727 10153 25895 10187
rect 25895 10153 25896 10187
rect 25726 10079 25896 10153
rect 25726 10045 25727 10079
rect 25727 10045 25895 10079
rect 25895 10045 25896 10079
rect 25726 10044 25896 10045
rect 26098 10187 26268 10188
rect 26098 10153 26099 10187
rect 26099 10153 26267 10187
rect 26267 10153 26268 10187
rect 26098 10079 26268 10153
rect 26098 10045 26099 10079
rect 26099 10045 26267 10079
rect 26267 10045 26268 10079
rect 26098 10044 26268 10045
rect 26470 10187 26640 10188
rect 26470 10153 26471 10187
rect 26471 10153 26639 10187
rect 26639 10153 26640 10187
rect 26470 10079 26640 10153
rect 26470 10045 26471 10079
rect 26471 10045 26639 10079
rect 26639 10045 26640 10079
rect 26470 10044 26640 10045
rect 26842 10187 27012 10188
rect 26842 10153 26843 10187
rect 26843 10153 27011 10187
rect 27011 10153 27012 10187
rect 26842 10079 27012 10153
rect 26842 10045 26843 10079
rect 26843 10045 27011 10079
rect 27011 10045 27012 10079
rect 26842 10044 27012 10045
rect 27214 10187 27384 10188
rect 27214 10153 27215 10187
rect 27215 10153 27383 10187
rect 27383 10153 27384 10187
rect 27214 10079 27384 10153
rect 27214 10045 27215 10079
rect 27215 10045 27383 10079
rect 27383 10045 27384 10079
rect 27214 10044 27384 10045
rect 27586 10187 27756 10188
rect 27586 10153 27587 10187
rect 27587 10153 27755 10187
rect 27755 10153 27756 10187
rect 27586 10079 27756 10153
rect 27586 10045 27587 10079
rect 27587 10045 27755 10079
rect 27755 10045 27756 10079
rect 27586 10044 27756 10045
rect 27958 10187 28128 10188
rect 27958 10153 27959 10187
rect 27959 10153 28127 10187
rect 28127 10153 28128 10187
rect 27958 10079 28128 10153
rect 27958 10045 27959 10079
rect 27959 10045 28127 10079
rect 28127 10045 28128 10079
rect 27958 10044 28128 10045
rect 28330 10187 28500 10188
rect 28330 10153 28331 10187
rect 28331 10153 28499 10187
rect 28499 10153 28500 10187
rect 28330 10079 28500 10153
rect 28330 10045 28331 10079
rect 28331 10045 28499 10079
rect 28499 10045 28500 10079
rect 28330 10044 28500 10045
rect 28702 10187 28872 10188
rect 28702 10153 28703 10187
rect 28703 10153 28871 10187
rect 28871 10153 28872 10187
rect 28702 10079 28872 10153
rect 28702 10045 28703 10079
rect 28703 10045 28871 10079
rect 28871 10045 28872 10079
rect 28702 10044 28872 10045
rect 29074 10187 29244 10188
rect 29074 10153 29075 10187
rect 29075 10153 29243 10187
rect 29243 10153 29244 10187
rect 29074 10079 29244 10153
rect 29074 10045 29075 10079
rect 29075 10045 29243 10079
rect 29243 10045 29244 10079
rect 29074 10044 29244 10045
rect 29446 10187 29616 10188
rect 29446 10153 29447 10187
rect 29447 10153 29615 10187
rect 29615 10153 29616 10187
rect 29446 10079 29616 10153
rect 29446 10045 29447 10079
rect 29447 10045 29615 10079
rect 29615 10045 29616 10079
rect 29446 10044 29616 10045
rect 29818 10187 29988 10188
rect 29818 10153 29819 10187
rect 29819 10153 29987 10187
rect 29987 10153 29988 10187
rect 29818 10079 29988 10153
rect 29818 10045 29819 10079
rect 29819 10045 29987 10079
rect 29987 10045 29988 10079
rect 29818 10044 29988 10045
rect 30190 10187 30360 10188
rect 30190 10153 30191 10187
rect 30191 10153 30359 10187
rect 30359 10153 30360 10187
rect 30190 10079 30360 10153
rect 30190 10045 30191 10079
rect 30191 10045 30359 10079
rect 30359 10045 30360 10079
rect 30190 10044 30360 10045
rect 30562 10187 30732 10188
rect 30562 10153 30563 10187
rect 30563 10153 30731 10187
rect 30731 10153 30732 10187
rect 30562 10079 30732 10153
rect 30562 10045 30563 10079
rect 30563 10045 30731 10079
rect 30731 10045 30732 10079
rect 30562 10044 30732 10045
rect 30934 10187 31104 10188
rect 30934 10153 30935 10187
rect 30935 10153 31103 10187
rect 31103 10153 31104 10187
rect 30934 10079 31104 10153
rect 30934 10045 30935 10079
rect 30935 10045 31103 10079
rect 31103 10045 31104 10079
rect 30934 10044 31104 10045
rect 25354 9551 25524 9552
rect 25354 9517 25355 9551
rect 25355 9517 25523 9551
rect 25523 9517 25524 9551
rect 25354 9443 25524 9517
rect 25354 9409 25355 9443
rect 25355 9409 25523 9443
rect 25523 9409 25524 9443
rect 25354 9408 25524 9409
rect 25726 9551 25896 9552
rect 25726 9517 25727 9551
rect 25727 9517 25895 9551
rect 25895 9517 25896 9551
rect 25726 9443 25896 9517
rect 25726 9409 25727 9443
rect 25727 9409 25895 9443
rect 25895 9409 25896 9443
rect 25726 9408 25896 9409
rect 26098 9551 26268 9552
rect 26098 9517 26099 9551
rect 26099 9517 26267 9551
rect 26267 9517 26268 9551
rect 26098 9443 26268 9517
rect 26098 9409 26099 9443
rect 26099 9409 26267 9443
rect 26267 9409 26268 9443
rect 26098 9408 26268 9409
rect 26470 9551 26640 9552
rect 26470 9517 26471 9551
rect 26471 9517 26639 9551
rect 26639 9517 26640 9551
rect 26470 9443 26640 9517
rect 26470 9409 26471 9443
rect 26471 9409 26639 9443
rect 26639 9409 26640 9443
rect 26470 9408 26640 9409
rect 26842 9551 27012 9552
rect 26842 9517 26843 9551
rect 26843 9517 27011 9551
rect 27011 9517 27012 9551
rect 26842 9443 27012 9517
rect 26842 9409 26843 9443
rect 26843 9409 27011 9443
rect 27011 9409 27012 9443
rect 26842 9408 27012 9409
rect 27214 9551 27384 9552
rect 27214 9517 27215 9551
rect 27215 9517 27383 9551
rect 27383 9517 27384 9551
rect 27214 9443 27384 9517
rect 27214 9409 27215 9443
rect 27215 9409 27383 9443
rect 27383 9409 27384 9443
rect 27214 9408 27384 9409
rect 27586 9551 27756 9552
rect 27586 9517 27587 9551
rect 27587 9517 27755 9551
rect 27755 9517 27756 9551
rect 27586 9443 27756 9517
rect 27586 9409 27587 9443
rect 27587 9409 27755 9443
rect 27755 9409 27756 9443
rect 27586 9408 27756 9409
rect 27958 9551 28128 9552
rect 27958 9517 27959 9551
rect 27959 9517 28127 9551
rect 28127 9517 28128 9551
rect 27958 9443 28128 9517
rect 27958 9409 27959 9443
rect 27959 9409 28127 9443
rect 28127 9409 28128 9443
rect 27958 9408 28128 9409
rect 28330 9551 28500 9552
rect 28330 9517 28331 9551
rect 28331 9517 28499 9551
rect 28499 9517 28500 9551
rect 28330 9443 28500 9517
rect 28330 9409 28331 9443
rect 28331 9409 28499 9443
rect 28499 9409 28500 9443
rect 28330 9408 28500 9409
rect 28702 9551 28872 9552
rect 28702 9517 28703 9551
rect 28703 9517 28871 9551
rect 28871 9517 28872 9551
rect 28702 9443 28872 9517
rect 28702 9409 28703 9443
rect 28703 9409 28871 9443
rect 28871 9409 28872 9443
rect 28702 9408 28872 9409
rect 29074 9551 29244 9552
rect 29074 9517 29075 9551
rect 29075 9517 29243 9551
rect 29243 9517 29244 9551
rect 29074 9443 29244 9517
rect 29074 9409 29075 9443
rect 29075 9409 29243 9443
rect 29243 9409 29244 9443
rect 29074 9408 29244 9409
rect 29446 9551 29616 9552
rect 29446 9517 29447 9551
rect 29447 9517 29615 9551
rect 29615 9517 29616 9551
rect 29446 9443 29616 9517
rect 29446 9409 29447 9443
rect 29447 9409 29615 9443
rect 29615 9409 29616 9443
rect 29446 9408 29616 9409
rect 29818 9551 29988 9552
rect 29818 9517 29819 9551
rect 29819 9517 29987 9551
rect 29987 9517 29988 9551
rect 29818 9443 29988 9517
rect 29818 9409 29819 9443
rect 29819 9409 29987 9443
rect 29987 9409 29988 9443
rect 29818 9408 29988 9409
rect 30190 9551 30360 9552
rect 30190 9517 30191 9551
rect 30191 9517 30359 9551
rect 30359 9517 30360 9551
rect 30190 9443 30360 9517
rect 30190 9409 30191 9443
rect 30191 9409 30359 9443
rect 30359 9409 30360 9443
rect 30190 9408 30360 9409
rect 30562 9551 30732 9552
rect 30562 9517 30563 9551
rect 30563 9517 30731 9551
rect 30731 9517 30732 9551
rect 30562 9443 30732 9517
rect 30562 9409 30563 9443
rect 30563 9409 30731 9443
rect 30731 9409 30732 9443
rect 30562 9408 30732 9409
rect 30934 9551 31104 9552
rect 30934 9517 30935 9551
rect 30935 9517 31103 9551
rect 31103 9517 31104 9551
rect 30934 9443 31104 9517
rect 30934 9409 30935 9443
rect 30935 9409 31103 9443
rect 31103 9409 31104 9443
rect 30934 9408 31104 9409
rect 24610 8915 24780 8928
rect 24610 8881 24611 8915
rect 24611 8881 24779 8915
rect 24779 8881 24780 8915
rect 24610 8868 24780 8881
rect 24982 8915 25152 8928
rect 24982 8881 24983 8915
rect 24983 8881 25151 8915
rect 25151 8881 25152 8915
rect 24982 8868 25152 8881
rect 25354 8915 25524 8928
rect 25354 8881 25355 8915
rect 25355 8881 25523 8915
rect 25523 8881 25524 8915
rect 25354 8868 25524 8881
rect 25726 8915 25896 8928
rect 25726 8881 25727 8915
rect 25727 8881 25895 8915
rect 25895 8881 25896 8915
rect 25726 8868 25896 8881
rect 26098 8915 26268 8928
rect 26098 8881 26099 8915
rect 26099 8881 26267 8915
rect 26267 8881 26268 8915
rect 26098 8868 26268 8881
rect 26470 8915 26640 8928
rect 26470 8881 26471 8915
rect 26471 8881 26639 8915
rect 26639 8881 26640 8915
rect 26470 8868 26640 8881
rect 26842 8915 27012 8928
rect 26842 8881 26843 8915
rect 26843 8881 27011 8915
rect 27011 8881 27012 8915
rect 26842 8868 27012 8881
rect 27214 8915 27384 8928
rect 27214 8881 27215 8915
rect 27215 8881 27383 8915
rect 27383 8881 27384 8915
rect 27214 8868 27384 8881
rect 27586 8915 27756 8928
rect 27586 8881 27587 8915
rect 27587 8881 27755 8915
rect 27755 8881 27756 8915
rect 27586 8868 27756 8881
rect 27958 8915 28128 8928
rect 27958 8881 27959 8915
rect 27959 8881 28127 8915
rect 28127 8881 28128 8915
rect 27958 8868 28128 8881
rect 28330 8915 28500 8928
rect 28330 8881 28331 8915
rect 28331 8881 28499 8915
rect 28499 8881 28500 8915
rect 28330 8868 28500 8881
rect 28702 8915 28872 8928
rect 28702 8881 28703 8915
rect 28703 8881 28871 8915
rect 28871 8881 28872 8915
rect 28702 8868 28872 8881
rect 29074 8915 29244 8928
rect 29074 8881 29075 8915
rect 29075 8881 29243 8915
rect 29243 8881 29244 8915
rect 29074 8868 29244 8881
rect 29446 8915 29616 8928
rect 29446 8881 29447 8915
rect 29447 8881 29615 8915
rect 29615 8881 29616 8915
rect 29446 8868 29616 8881
rect 29818 8915 29988 8928
rect 29818 8881 29819 8915
rect 29819 8881 29987 8915
rect 29987 8881 29988 8915
rect 29818 8868 29988 8881
rect 30190 8915 30360 8928
rect 30190 8881 30191 8915
rect 30191 8881 30359 8915
rect 30359 8881 30360 8915
rect 30190 8868 30360 8881
rect 30562 8915 30732 8928
rect 30562 8881 30563 8915
rect 30563 8881 30731 8915
rect 30731 8881 30732 8915
rect 30562 8868 30732 8881
rect 30934 8915 31104 8928
rect 30934 8881 30935 8915
rect 30935 8881 31103 8915
rect 31103 8881 31104 8915
rect 30934 8868 31104 8881
rect 20890 8327 21060 8342
rect 20890 8293 20891 8327
rect 20891 8293 21059 8327
rect 21059 8293 21060 8327
rect 20890 8278 21060 8293
rect 21262 8327 21432 8342
rect 21262 8293 21263 8327
rect 21263 8293 21431 8327
rect 21431 8293 21432 8327
rect 21262 8278 21432 8293
rect 21634 8327 21804 8342
rect 21634 8293 21635 8327
rect 21635 8293 21803 8327
rect 21803 8293 21804 8327
rect 21634 8278 21804 8293
rect 22006 8327 22176 8342
rect 22006 8293 22007 8327
rect 22007 8293 22175 8327
rect 22175 8293 22176 8327
rect 22006 8278 22176 8293
rect 22378 8327 22548 8342
rect 22378 8293 22379 8327
rect 22379 8293 22547 8327
rect 22547 8293 22548 8327
rect 22378 8278 22548 8293
rect 22750 8327 22920 8342
rect 22750 8293 22751 8327
rect 22751 8293 22919 8327
rect 22919 8293 22920 8327
rect 22750 8278 22920 8293
rect 23122 8327 23292 8342
rect 23122 8293 23123 8327
rect 23123 8293 23291 8327
rect 23291 8293 23292 8327
rect 23122 8278 23292 8293
rect 23494 8327 23664 8342
rect 23494 8293 23495 8327
rect 23495 8293 23663 8327
rect 23663 8293 23664 8327
rect 23494 8278 23664 8293
rect 20890 7399 21060 7400
rect 20890 7365 20891 7399
rect 20891 7365 21059 7399
rect 21059 7365 21060 7399
rect 20890 7291 21060 7365
rect 20890 7257 20891 7291
rect 20891 7257 21059 7291
rect 21059 7257 21060 7291
rect 20890 7256 21060 7257
rect 21262 7399 21432 7400
rect 21262 7365 21263 7399
rect 21263 7365 21431 7399
rect 21431 7365 21432 7399
rect 21262 7291 21432 7365
rect 21262 7257 21263 7291
rect 21263 7257 21431 7291
rect 21431 7257 21432 7291
rect 21262 7256 21432 7257
rect 21634 7399 21804 7400
rect 21634 7365 21635 7399
rect 21635 7365 21803 7399
rect 21803 7365 21804 7399
rect 21634 7291 21804 7365
rect 21634 7257 21635 7291
rect 21635 7257 21803 7291
rect 21803 7257 21804 7291
rect 21634 7256 21804 7257
rect 22006 7399 22176 7400
rect 22006 7365 22007 7399
rect 22007 7365 22175 7399
rect 22175 7365 22176 7399
rect 22006 7291 22176 7365
rect 22006 7257 22007 7291
rect 22007 7257 22175 7291
rect 22175 7257 22176 7291
rect 22006 7256 22176 7257
rect 22378 7399 22548 7400
rect 22378 7365 22379 7399
rect 22379 7365 22547 7399
rect 22547 7365 22548 7399
rect 22378 7291 22548 7365
rect 22378 7257 22379 7291
rect 22379 7257 22547 7291
rect 22547 7257 22548 7291
rect 22378 7256 22548 7257
rect 22750 7399 22920 7400
rect 22750 7365 22751 7399
rect 22751 7365 22919 7399
rect 22919 7365 22920 7399
rect 22750 7291 22920 7365
rect 22750 7257 22751 7291
rect 22751 7257 22919 7291
rect 22919 7257 22920 7291
rect 22750 7256 22920 7257
rect 23122 7399 23292 7400
rect 23122 7365 23123 7399
rect 23123 7365 23291 7399
rect 23291 7365 23292 7399
rect 23122 7291 23292 7365
rect 23122 7257 23123 7291
rect 23123 7257 23291 7291
rect 23291 7257 23292 7291
rect 23122 7256 23292 7257
rect 23494 7399 23664 7400
rect 23494 7365 23495 7399
rect 23495 7365 23663 7399
rect 23663 7365 23664 7399
rect 23494 7291 23664 7365
rect 23494 7257 23495 7291
rect 23495 7257 23663 7291
rect 23663 7257 23664 7291
rect 23494 7256 23664 7257
rect 20890 6363 21060 6364
rect 20890 6329 20891 6363
rect 20891 6329 21059 6363
rect 21059 6329 21060 6363
rect 20890 6255 21060 6329
rect 20890 6221 20891 6255
rect 20891 6221 21059 6255
rect 21059 6221 21060 6255
rect 20890 6220 21060 6221
rect 21262 6363 21432 6364
rect 21262 6329 21263 6363
rect 21263 6329 21431 6363
rect 21431 6329 21432 6363
rect 21262 6255 21432 6329
rect 21262 6221 21263 6255
rect 21263 6221 21431 6255
rect 21431 6221 21432 6255
rect 21262 6220 21432 6221
rect 21634 6363 21804 6364
rect 21634 6329 21635 6363
rect 21635 6329 21803 6363
rect 21803 6329 21804 6363
rect 21634 6255 21804 6329
rect 21634 6221 21635 6255
rect 21635 6221 21803 6255
rect 21803 6221 21804 6255
rect 21634 6220 21804 6221
rect 22006 6363 22176 6364
rect 22006 6329 22007 6363
rect 22007 6329 22175 6363
rect 22175 6329 22176 6363
rect 22006 6255 22176 6329
rect 22006 6221 22007 6255
rect 22007 6221 22175 6255
rect 22175 6221 22176 6255
rect 22006 6220 22176 6221
rect 22378 6363 22548 6364
rect 22378 6329 22379 6363
rect 22379 6329 22547 6363
rect 22547 6329 22548 6363
rect 22378 6255 22548 6329
rect 22378 6221 22379 6255
rect 22379 6221 22547 6255
rect 22547 6221 22548 6255
rect 22378 6220 22548 6221
rect 22750 6363 22920 6364
rect 22750 6329 22751 6363
rect 22751 6329 22919 6363
rect 22919 6329 22920 6363
rect 22750 6255 22920 6329
rect 22750 6221 22751 6255
rect 22751 6221 22919 6255
rect 22919 6221 22920 6255
rect 22750 6220 22920 6221
rect 23122 6363 23292 6364
rect 23122 6329 23123 6363
rect 23123 6329 23291 6363
rect 23291 6329 23292 6363
rect 23122 6255 23292 6329
rect 23122 6221 23123 6255
rect 23123 6221 23291 6255
rect 23291 6221 23292 6255
rect 23122 6220 23292 6221
rect 23494 6363 23664 6364
rect 23494 6329 23495 6363
rect 23495 6329 23663 6363
rect 23663 6329 23664 6363
rect 23494 6255 23664 6329
rect 23494 6221 23495 6255
rect 23495 6221 23663 6255
rect 23663 6221 23664 6255
rect 23494 6220 23664 6221
rect 20890 5327 21060 5328
rect 20890 5293 20891 5327
rect 20891 5293 21059 5327
rect 21059 5293 21060 5327
rect 20890 5219 21060 5293
rect 20890 5185 20891 5219
rect 20891 5185 21059 5219
rect 21059 5185 21060 5219
rect 20890 5184 21060 5185
rect 21262 5327 21432 5328
rect 21262 5293 21263 5327
rect 21263 5293 21431 5327
rect 21431 5293 21432 5327
rect 21262 5219 21432 5293
rect 21262 5185 21263 5219
rect 21263 5185 21431 5219
rect 21431 5185 21432 5219
rect 21262 5184 21432 5185
rect 21634 5327 21804 5328
rect 21634 5293 21635 5327
rect 21635 5293 21803 5327
rect 21803 5293 21804 5327
rect 21634 5219 21804 5293
rect 21634 5185 21635 5219
rect 21635 5185 21803 5219
rect 21803 5185 21804 5219
rect 21634 5184 21804 5185
rect 22006 5327 22176 5328
rect 22006 5293 22007 5327
rect 22007 5293 22175 5327
rect 22175 5293 22176 5327
rect 22006 5219 22176 5293
rect 22006 5185 22007 5219
rect 22007 5185 22175 5219
rect 22175 5185 22176 5219
rect 22006 5184 22176 5185
rect 22378 5327 22548 5328
rect 22378 5293 22379 5327
rect 22379 5293 22547 5327
rect 22547 5293 22548 5327
rect 22378 5219 22548 5293
rect 22378 5185 22379 5219
rect 22379 5185 22547 5219
rect 22547 5185 22548 5219
rect 22378 5184 22548 5185
rect 22750 5327 22920 5328
rect 22750 5293 22751 5327
rect 22751 5293 22919 5327
rect 22919 5293 22920 5327
rect 22750 5219 22920 5293
rect 22750 5185 22751 5219
rect 22751 5185 22919 5219
rect 22919 5185 22920 5219
rect 22750 5184 22920 5185
rect 23122 5327 23292 5328
rect 23122 5293 23123 5327
rect 23123 5293 23291 5327
rect 23291 5293 23292 5327
rect 23122 5219 23292 5293
rect 23122 5185 23123 5219
rect 23123 5185 23291 5219
rect 23291 5185 23292 5219
rect 23122 5184 23292 5185
rect 23494 5327 23664 5328
rect 23494 5293 23495 5327
rect 23495 5293 23663 5327
rect 23663 5293 23664 5327
rect 23494 5219 23664 5293
rect 23494 5185 23495 5219
rect 23495 5185 23663 5219
rect 23663 5185 23664 5219
rect 23494 5184 23664 5185
rect 20890 4291 21060 4302
rect 20890 4257 20891 4291
rect 20891 4257 21059 4291
rect 21059 4257 21060 4291
rect 20890 4248 21060 4257
rect 21262 4291 21432 4302
rect 21262 4257 21263 4291
rect 21263 4257 21431 4291
rect 21431 4257 21432 4291
rect 21262 4248 21432 4257
rect 21634 4291 21804 4302
rect 21634 4257 21635 4291
rect 21635 4257 21803 4291
rect 21803 4257 21804 4291
rect 21634 4248 21804 4257
rect 22006 4291 22176 4302
rect 22006 4257 22007 4291
rect 22007 4257 22175 4291
rect 22175 4257 22176 4291
rect 22006 4248 22176 4257
rect 22378 4291 22548 4302
rect 22378 4257 22379 4291
rect 22379 4257 22547 4291
rect 22547 4257 22548 4291
rect 22378 4248 22548 4257
rect 22750 4291 22920 4302
rect 22750 4257 22751 4291
rect 22751 4257 22919 4291
rect 22919 4257 22920 4291
rect 22750 4248 22920 4257
rect 23122 4291 23292 4302
rect 23122 4257 23123 4291
rect 23123 4257 23291 4291
rect 23291 4257 23292 4291
rect 23122 4248 23292 4257
rect 21870 3782 22684 3962
rect 20890 3633 21060 3644
rect 20890 3599 20891 3633
rect 20891 3599 21059 3633
rect 21059 3599 21060 3633
rect 20890 3588 21060 3599
rect 21262 3633 21432 3644
rect 21262 3599 21263 3633
rect 21263 3599 21431 3633
rect 21431 3599 21432 3633
rect 21262 3588 21432 3599
rect 21634 3633 21804 3644
rect 21634 3599 21635 3633
rect 21635 3599 21803 3633
rect 21803 3599 21804 3633
rect 21634 3588 21804 3599
rect 22006 3633 22176 3644
rect 22006 3599 22007 3633
rect 22007 3599 22175 3633
rect 22175 3599 22176 3633
rect 22006 3588 22176 3599
rect 22378 3633 22548 3644
rect 22378 3599 22379 3633
rect 22379 3599 22547 3633
rect 22547 3599 22548 3633
rect 22378 3588 22548 3599
rect 23494 4291 23664 4302
rect 23494 4257 23495 4291
rect 23495 4257 23663 4291
rect 23663 4257 23664 4291
rect 23494 4248 23664 4257
rect 22750 3633 22920 3644
rect 22750 3599 22751 3633
rect 22751 3599 22919 3633
rect 22919 3599 22920 3633
rect 22750 3588 22920 3599
rect 23122 3633 23292 3644
rect 23122 3599 23123 3633
rect 23123 3599 23291 3633
rect 23291 3599 23292 3633
rect 23122 3588 23292 3599
rect 23494 3633 23664 3644
rect 23494 3599 23495 3633
rect 23495 3599 23663 3633
rect 23663 3599 23664 3633
rect 23494 3588 23664 3599
rect 23866 3633 24036 3644
rect 23866 3599 23867 3633
rect 23867 3599 24035 3633
rect 24035 3599 24036 3633
rect 23866 3588 24036 3599
rect 24238 3633 24408 3644
rect 24238 3599 24239 3633
rect 24239 3599 24407 3633
rect 24407 3599 24408 3633
rect 24238 3588 24408 3599
rect 24610 3633 24780 3644
rect 24610 3599 24611 3633
rect 24611 3599 24779 3633
rect 24779 3599 24780 3633
rect 24610 3588 24780 3599
rect 24982 3633 25152 3644
rect 24982 3599 24983 3633
rect 24983 3599 25151 3633
rect 25151 3599 25152 3633
rect 24982 3588 25152 3599
rect 25354 3633 25524 3644
rect 25354 3599 25355 3633
rect 25355 3599 25523 3633
rect 25523 3599 25524 3633
rect 25354 3588 25524 3599
rect 25726 3633 25896 3644
rect 25726 3599 25727 3633
rect 25727 3599 25895 3633
rect 25895 3599 25896 3633
rect 25726 3588 25896 3599
rect 26098 3633 26268 3644
rect 26098 3599 26099 3633
rect 26099 3599 26267 3633
rect 26267 3599 26268 3633
rect 26098 3588 26268 3599
rect 26470 3633 26640 3644
rect 26470 3599 26471 3633
rect 26471 3599 26639 3633
rect 26639 3599 26640 3633
rect 26470 3588 26640 3599
rect 26842 3633 27012 3644
rect 26842 3599 26843 3633
rect 26843 3599 27011 3633
rect 27011 3599 27012 3633
rect 26842 3588 27012 3599
rect 27214 3633 27384 3644
rect 27214 3599 27215 3633
rect 27215 3599 27383 3633
rect 27383 3599 27384 3633
rect 27214 3588 27384 3599
rect 27586 3633 27756 3644
rect 27586 3599 27587 3633
rect 27587 3599 27755 3633
rect 27755 3599 27756 3633
rect 27586 3588 27756 3599
rect 27958 3633 28128 3644
rect 27958 3599 27959 3633
rect 27959 3599 28127 3633
rect 28127 3599 28128 3633
rect 27958 3588 28128 3599
rect 28330 3633 28500 3644
rect 28330 3599 28331 3633
rect 28331 3599 28499 3633
rect 28499 3599 28500 3633
rect 28330 3588 28500 3599
rect 28702 3633 28872 3644
rect 28702 3599 28703 3633
rect 28703 3599 28871 3633
rect 28871 3599 28872 3633
rect 28702 3588 28872 3599
rect 29074 3633 29244 3644
rect 29074 3599 29075 3633
rect 29075 3599 29243 3633
rect 29243 3599 29244 3633
rect 29074 3588 29244 3599
rect 29446 3633 29616 3644
rect 29446 3599 29447 3633
rect 29447 3599 29615 3633
rect 29615 3599 29616 3633
rect 29446 3588 29616 3599
rect 20890 3323 21060 3324
rect 20890 3289 20891 3323
rect 20891 3289 21059 3323
rect 21059 3289 21060 3323
rect 20890 3215 21060 3289
rect 20890 3181 20891 3215
rect 20891 3181 21059 3215
rect 21059 3181 21060 3215
rect 20890 3180 21060 3181
rect 21262 3323 21432 3324
rect 21262 3289 21263 3323
rect 21263 3289 21431 3323
rect 21431 3289 21432 3323
rect 21262 3215 21432 3289
rect 21262 3181 21263 3215
rect 21263 3181 21431 3215
rect 21431 3181 21432 3215
rect 21262 3180 21432 3181
rect 21634 3323 21804 3324
rect 21634 3289 21635 3323
rect 21635 3289 21803 3323
rect 21803 3289 21804 3323
rect 21634 3215 21804 3289
rect 21634 3181 21635 3215
rect 21635 3181 21803 3215
rect 21803 3181 21804 3215
rect 21634 3180 21804 3181
rect 22006 3323 22176 3324
rect 22006 3289 22007 3323
rect 22007 3289 22175 3323
rect 22175 3289 22176 3323
rect 22006 3215 22176 3289
rect 22006 3181 22007 3215
rect 22007 3181 22175 3215
rect 22175 3181 22176 3215
rect 22006 3180 22176 3181
rect 22378 3323 22548 3324
rect 22378 3289 22379 3323
rect 22379 3289 22547 3323
rect 22547 3289 22548 3323
rect 22378 3215 22548 3289
rect 22378 3181 22379 3215
rect 22379 3181 22547 3215
rect 22547 3181 22548 3215
rect 22378 3180 22548 3181
rect 22750 3323 22920 3324
rect 22750 3289 22751 3323
rect 22751 3289 22919 3323
rect 22919 3289 22920 3323
rect 22750 3215 22920 3289
rect 22750 3181 22751 3215
rect 22751 3181 22919 3215
rect 22919 3181 22920 3215
rect 22750 3180 22920 3181
rect 23122 3323 23292 3324
rect 23122 3289 23123 3323
rect 23123 3289 23291 3323
rect 23291 3289 23292 3323
rect 23122 3215 23292 3289
rect 23122 3181 23123 3215
rect 23123 3181 23291 3215
rect 23291 3181 23292 3215
rect 23122 3180 23292 3181
rect 23494 3323 23664 3324
rect 23494 3289 23495 3323
rect 23495 3289 23663 3323
rect 23663 3289 23664 3323
rect 23494 3215 23664 3289
rect 23494 3181 23495 3215
rect 23495 3181 23663 3215
rect 23663 3181 23664 3215
rect 23494 3180 23664 3181
rect 23866 3323 24036 3324
rect 23866 3289 23867 3323
rect 23867 3289 24035 3323
rect 24035 3289 24036 3323
rect 23866 3215 24036 3289
rect 23866 3181 23867 3215
rect 23867 3181 24035 3215
rect 24035 3181 24036 3215
rect 23866 3180 24036 3181
rect 24238 3323 24408 3324
rect 24238 3289 24239 3323
rect 24239 3289 24407 3323
rect 24407 3289 24408 3323
rect 24238 3215 24408 3289
rect 24238 3181 24239 3215
rect 24239 3181 24407 3215
rect 24407 3181 24408 3215
rect 24238 3180 24408 3181
rect 24610 3323 24780 3324
rect 24610 3289 24611 3323
rect 24611 3289 24779 3323
rect 24779 3289 24780 3323
rect 24610 3215 24780 3289
rect 24610 3181 24611 3215
rect 24611 3181 24779 3215
rect 24779 3181 24780 3215
rect 24610 3180 24780 3181
rect 24982 3323 25152 3324
rect 24982 3289 24983 3323
rect 24983 3289 25151 3323
rect 25151 3289 25152 3323
rect 24982 3215 25152 3289
rect 24982 3181 24983 3215
rect 24983 3181 25151 3215
rect 25151 3181 25152 3215
rect 24982 3180 25152 3181
rect 25354 3323 25524 3324
rect 25354 3289 25355 3323
rect 25355 3289 25523 3323
rect 25523 3289 25524 3323
rect 25354 3215 25524 3289
rect 25354 3181 25355 3215
rect 25355 3181 25523 3215
rect 25523 3181 25524 3215
rect 25354 3180 25524 3181
rect 25726 3323 25896 3324
rect 25726 3289 25727 3323
rect 25727 3289 25895 3323
rect 25895 3289 25896 3323
rect 25726 3215 25896 3289
rect 25726 3181 25727 3215
rect 25727 3181 25895 3215
rect 25895 3181 25896 3215
rect 25726 3180 25896 3181
rect 26098 3323 26268 3324
rect 26098 3289 26099 3323
rect 26099 3289 26267 3323
rect 26267 3289 26268 3323
rect 26098 3215 26268 3289
rect 26098 3181 26099 3215
rect 26099 3181 26267 3215
rect 26267 3181 26268 3215
rect 26098 3180 26268 3181
rect 26470 3323 26640 3324
rect 26470 3289 26471 3323
rect 26471 3289 26639 3323
rect 26639 3289 26640 3323
rect 26470 3215 26640 3289
rect 26470 3181 26471 3215
rect 26471 3181 26639 3215
rect 26639 3181 26640 3215
rect 26470 3180 26640 3181
rect 26842 3323 27012 3324
rect 26842 3289 26843 3323
rect 26843 3289 27011 3323
rect 27011 3289 27012 3323
rect 26842 3215 27012 3289
rect 26842 3181 26843 3215
rect 26843 3181 27011 3215
rect 27011 3181 27012 3215
rect 26842 3180 27012 3181
rect 27214 3323 27384 3324
rect 27214 3289 27215 3323
rect 27215 3289 27383 3323
rect 27383 3289 27384 3323
rect 27214 3215 27384 3289
rect 27214 3181 27215 3215
rect 27215 3181 27383 3215
rect 27383 3181 27384 3215
rect 27214 3180 27384 3181
rect 27586 3323 27756 3324
rect 27586 3289 27587 3323
rect 27587 3289 27755 3323
rect 27755 3289 27756 3323
rect 27586 3215 27756 3289
rect 27586 3181 27587 3215
rect 27587 3181 27755 3215
rect 27755 3181 27756 3215
rect 27586 3180 27756 3181
rect 27958 3323 28128 3324
rect 27958 3289 27959 3323
rect 27959 3289 28127 3323
rect 28127 3289 28128 3323
rect 27958 3215 28128 3289
rect 27958 3181 27959 3215
rect 27959 3181 28127 3215
rect 28127 3181 28128 3215
rect 27958 3180 28128 3181
rect 28330 3323 28500 3324
rect 28330 3289 28331 3323
rect 28331 3289 28499 3323
rect 28499 3289 28500 3323
rect 28330 3215 28500 3289
rect 28330 3181 28331 3215
rect 28331 3181 28499 3215
rect 28499 3181 28500 3215
rect 28330 3180 28500 3181
rect 28702 3323 28872 3324
rect 28702 3289 28703 3323
rect 28703 3289 28871 3323
rect 28871 3289 28872 3323
rect 28702 3215 28872 3289
rect 28702 3181 28703 3215
rect 28703 3181 28871 3215
rect 28871 3181 28872 3215
rect 28702 3180 28872 3181
rect 29074 3323 29244 3324
rect 29074 3289 29075 3323
rect 29075 3289 29243 3323
rect 29243 3289 29244 3323
rect 29074 3215 29244 3289
rect 29074 3181 29075 3215
rect 29075 3181 29243 3215
rect 29243 3181 29244 3215
rect 29074 3180 29244 3181
rect 29446 3323 29616 3324
rect 29446 3289 29447 3323
rect 29447 3289 29615 3323
rect 29615 3289 29616 3323
rect 29446 3215 29616 3289
rect 29446 3181 29447 3215
rect 29447 3181 29615 3215
rect 29615 3181 29616 3215
rect 29446 3180 29616 3181
rect 20890 2905 21060 2906
rect 20890 2871 20891 2905
rect 20891 2871 21059 2905
rect 21059 2871 21060 2905
rect 20890 2797 21060 2871
rect 20890 2763 20891 2797
rect 20891 2763 21059 2797
rect 21059 2763 21060 2797
rect 20890 2762 21060 2763
rect 21262 2905 21432 2906
rect 21262 2871 21263 2905
rect 21263 2871 21431 2905
rect 21431 2871 21432 2905
rect 21262 2797 21432 2871
rect 21262 2763 21263 2797
rect 21263 2763 21431 2797
rect 21431 2763 21432 2797
rect 21262 2762 21432 2763
rect 21634 2905 21804 2906
rect 21634 2871 21635 2905
rect 21635 2871 21803 2905
rect 21803 2871 21804 2905
rect 21634 2797 21804 2871
rect 21634 2763 21635 2797
rect 21635 2763 21803 2797
rect 21803 2763 21804 2797
rect 21634 2762 21804 2763
rect 22006 2905 22176 2906
rect 22006 2871 22007 2905
rect 22007 2871 22175 2905
rect 22175 2871 22176 2905
rect 22006 2797 22176 2871
rect 22006 2763 22007 2797
rect 22007 2763 22175 2797
rect 22175 2763 22176 2797
rect 22006 2762 22176 2763
rect 22378 2905 22548 2906
rect 22378 2871 22379 2905
rect 22379 2871 22547 2905
rect 22547 2871 22548 2905
rect 22378 2797 22548 2871
rect 22378 2763 22379 2797
rect 22379 2763 22547 2797
rect 22547 2763 22548 2797
rect 22378 2762 22548 2763
rect 22750 2905 22920 2906
rect 22750 2871 22751 2905
rect 22751 2871 22919 2905
rect 22919 2871 22920 2905
rect 22750 2797 22920 2871
rect 22750 2763 22751 2797
rect 22751 2763 22919 2797
rect 22919 2763 22920 2797
rect 22750 2762 22920 2763
rect 23122 2905 23292 2906
rect 23122 2871 23123 2905
rect 23123 2871 23291 2905
rect 23291 2871 23292 2905
rect 23122 2797 23292 2871
rect 23122 2763 23123 2797
rect 23123 2763 23291 2797
rect 23291 2763 23292 2797
rect 23122 2762 23292 2763
rect 23494 2905 23664 2906
rect 23494 2871 23495 2905
rect 23495 2871 23663 2905
rect 23663 2871 23664 2905
rect 23494 2797 23664 2871
rect 23494 2763 23495 2797
rect 23495 2763 23663 2797
rect 23663 2763 23664 2797
rect 23494 2762 23664 2763
rect 23866 2905 24036 2906
rect 23866 2871 23867 2905
rect 23867 2871 24035 2905
rect 24035 2871 24036 2905
rect 23866 2797 24036 2871
rect 23866 2763 23867 2797
rect 23867 2763 24035 2797
rect 24035 2763 24036 2797
rect 23866 2762 24036 2763
rect 24238 2905 24408 2906
rect 24238 2871 24239 2905
rect 24239 2871 24407 2905
rect 24407 2871 24408 2905
rect 24238 2797 24408 2871
rect 24238 2763 24239 2797
rect 24239 2763 24407 2797
rect 24407 2763 24408 2797
rect 24238 2762 24408 2763
rect 24610 2905 24780 2906
rect 24610 2871 24611 2905
rect 24611 2871 24779 2905
rect 24779 2871 24780 2905
rect 24610 2797 24780 2871
rect 24610 2763 24611 2797
rect 24611 2763 24779 2797
rect 24779 2763 24780 2797
rect 24610 2762 24780 2763
rect 24982 2905 25152 2906
rect 24982 2871 24983 2905
rect 24983 2871 25151 2905
rect 25151 2871 25152 2905
rect 24982 2797 25152 2871
rect 24982 2763 24983 2797
rect 24983 2763 25151 2797
rect 25151 2763 25152 2797
rect 24982 2762 25152 2763
rect 25354 2905 25524 2906
rect 25354 2871 25355 2905
rect 25355 2871 25523 2905
rect 25523 2871 25524 2905
rect 25354 2797 25524 2871
rect 25354 2763 25355 2797
rect 25355 2763 25523 2797
rect 25523 2763 25524 2797
rect 25354 2762 25524 2763
rect 25726 2905 25896 2906
rect 25726 2871 25727 2905
rect 25727 2871 25895 2905
rect 25895 2871 25896 2905
rect 25726 2797 25896 2871
rect 25726 2763 25727 2797
rect 25727 2763 25895 2797
rect 25895 2763 25896 2797
rect 25726 2762 25896 2763
rect 26098 2905 26268 2906
rect 26098 2871 26099 2905
rect 26099 2871 26267 2905
rect 26267 2871 26268 2905
rect 26098 2797 26268 2871
rect 26098 2763 26099 2797
rect 26099 2763 26267 2797
rect 26267 2763 26268 2797
rect 26098 2762 26268 2763
rect 26470 2905 26640 2906
rect 26470 2871 26471 2905
rect 26471 2871 26639 2905
rect 26639 2871 26640 2905
rect 26470 2797 26640 2871
rect 26470 2763 26471 2797
rect 26471 2763 26639 2797
rect 26639 2763 26640 2797
rect 26470 2762 26640 2763
rect 26842 2905 27012 2906
rect 26842 2871 26843 2905
rect 26843 2871 27011 2905
rect 27011 2871 27012 2905
rect 26842 2797 27012 2871
rect 26842 2763 26843 2797
rect 26843 2763 27011 2797
rect 27011 2763 27012 2797
rect 26842 2762 27012 2763
rect 27214 2905 27384 2906
rect 27214 2871 27215 2905
rect 27215 2871 27383 2905
rect 27383 2871 27384 2905
rect 27214 2797 27384 2871
rect 27214 2763 27215 2797
rect 27215 2763 27383 2797
rect 27383 2763 27384 2797
rect 27214 2762 27384 2763
rect 27586 2905 27756 2906
rect 27586 2871 27587 2905
rect 27587 2871 27755 2905
rect 27755 2871 27756 2905
rect 27586 2797 27756 2871
rect 27586 2763 27587 2797
rect 27587 2763 27755 2797
rect 27755 2763 27756 2797
rect 27586 2762 27756 2763
rect 27958 2905 28128 2906
rect 27958 2871 27959 2905
rect 27959 2871 28127 2905
rect 28127 2871 28128 2905
rect 27958 2797 28128 2871
rect 27958 2763 27959 2797
rect 27959 2763 28127 2797
rect 28127 2763 28128 2797
rect 27958 2762 28128 2763
rect 28330 2905 28500 2906
rect 28330 2871 28331 2905
rect 28331 2871 28499 2905
rect 28499 2871 28500 2905
rect 28330 2797 28500 2871
rect 28330 2763 28331 2797
rect 28331 2763 28499 2797
rect 28499 2763 28500 2797
rect 28330 2762 28500 2763
rect 28702 2905 28872 2906
rect 28702 2871 28703 2905
rect 28703 2871 28871 2905
rect 28871 2871 28872 2905
rect 28702 2797 28872 2871
rect 28702 2763 28703 2797
rect 28703 2763 28871 2797
rect 28871 2763 28872 2797
rect 28702 2762 28872 2763
rect 29074 2905 29244 2906
rect 29074 2871 29075 2905
rect 29075 2871 29243 2905
rect 29243 2871 29244 2905
rect 29074 2797 29244 2871
rect 29074 2763 29075 2797
rect 29075 2763 29243 2797
rect 29243 2763 29244 2797
rect 29074 2762 29244 2763
rect 29446 2905 29616 2906
rect 29446 2871 29447 2905
rect 29447 2871 29615 2905
rect 29615 2871 29616 2905
rect 29446 2797 29616 2871
rect 29446 2763 29447 2797
rect 29447 2763 29615 2797
rect 29615 2763 29616 2797
rect 29446 2762 29616 2763
rect 20890 2487 21060 2488
rect 20890 2453 20891 2487
rect 20891 2453 21059 2487
rect 21059 2453 21060 2487
rect 20890 2379 21060 2453
rect 20890 2345 20891 2379
rect 20891 2345 21059 2379
rect 21059 2345 21060 2379
rect 20890 2344 21060 2345
rect 21262 2487 21432 2488
rect 21262 2453 21263 2487
rect 21263 2453 21431 2487
rect 21431 2453 21432 2487
rect 21262 2379 21432 2453
rect 21262 2345 21263 2379
rect 21263 2345 21431 2379
rect 21431 2345 21432 2379
rect 21262 2344 21432 2345
rect 21634 2487 21804 2488
rect 21634 2453 21635 2487
rect 21635 2453 21803 2487
rect 21803 2453 21804 2487
rect 21634 2379 21804 2453
rect 21634 2345 21635 2379
rect 21635 2345 21803 2379
rect 21803 2345 21804 2379
rect 21634 2344 21804 2345
rect 22006 2487 22176 2488
rect 22006 2453 22007 2487
rect 22007 2453 22175 2487
rect 22175 2453 22176 2487
rect 22006 2379 22176 2453
rect 22006 2345 22007 2379
rect 22007 2345 22175 2379
rect 22175 2345 22176 2379
rect 22006 2344 22176 2345
rect 22378 2487 22548 2488
rect 22378 2453 22379 2487
rect 22379 2453 22547 2487
rect 22547 2453 22548 2487
rect 22378 2379 22548 2453
rect 22378 2345 22379 2379
rect 22379 2345 22547 2379
rect 22547 2345 22548 2379
rect 22378 2344 22548 2345
rect 22750 2487 22920 2488
rect 22750 2453 22751 2487
rect 22751 2453 22919 2487
rect 22919 2453 22920 2487
rect 22750 2379 22920 2453
rect 22750 2345 22751 2379
rect 22751 2345 22919 2379
rect 22919 2345 22920 2379
rect 22750 2344 22920 2345
rect 23122 2487 23292 2488
rect 23122 2453 23123 2487
rect 23123 2453 23291 2487
rect 23291 2453 23292 2487
rect 23122 2379 23292 2453
rect 23122 2345 23123 2379
rect 23123 2345 23291 2379
rect 23291 2345 23292 2379
rect 23122 2344 23292 2345
rect 23494 2487 23664 2488
rect 23494 2453 23495 2487
rect 23495 2453 23663 2487
rect 23663 2453 23664 2487
rect 23494 2379 23664 2453
rect 23494 2345 23495 2379
rect 23495 2345 23663 2379
rect 23663 2345 23664 2379
rect 23494 2344 23664 2345
rect 23866 2487 24036 2488
rect 23866 2453 23867 2487
rect 23867 2453 24035 2487
rect 24035 2453 24036 2487
rect 23866 2379 24036 2453
rect 23866 2345 23867 2379
rect 23867 2345 24035 2379
rect 24035 2345 24036 2379
rect 23866 2344 24036 2345
rect 24238 2487 24408 2488
rect 24238 2453 24239 2487
rect 24239 2453 24407 2487
rect 24407 2453 24408 2487
rect 24238 2379 24408 2453
rect 24238 2345 24239 2379
rect 24239 2345 24407 2379
rect 24407 2345 24408 2379
rect 24238 2344 24408 2345
rect 24610 2487 24780 2488
rect 24610 2453 24611 2487
rect 24611 2453 24779 2487
rect 24779 2453 24780 2487
rect 24610 2379 24780 2453
rect 24610 2345 24611 2379
rect 24611 2345 24779 2379
rect 24779 2345 24780 2379
rect 24610 2344 24780 2345
rect 24982 2487 25152 2488
rect 24982 2453 24983 2487
rect 24983 2453 25151 2487
rect 25151 2453 25152 2487
rect 24982 2379 25152 2453
rect 24982 2345 24983 2379
rect 24983 2345 25151 2379
rect 25151 2345 25152 2379
rect 24982 2344 25152 2345
rect 25354 2487 25524 2488
rect 25354 2453 25355 2487
rect 25355 2453 25523 2487
rect 25523 2453 25524 2487
rect 25354 2379 25524 2453
rect 25354 2345 25355 2379
rect 25355 2345 25523 2379
rect 25523 2345 25524 2379
rect 25354 2344 25524 2345
rect 25726 2487 25896 2488
rect 25726 2453 25727 2487
rect 25727 2453 25895 2487
rect 25895 2453 25896 2487
rect 25726 2379 25896 2453
rect 25726 2345 25727 2379
rect 25727 2345 25895 2379
rect 25895 2345 25896 2379
rect 25726 2344 25896 2345
rect 26098 2487 26268 2488
rect 26098 2453 26099 2487
rect 26099 2453 26267 2487
rect 26267 2453 26268 2487
rect 26098 2379 26268 2453
rect 26098 2345 26099 2379
rect 26099 2345 26267 2379
rect 26267 2345 26268 2379
rect 26098 2344 26268 2345
rect 26470 2487 26640 2488
rect 26470 2453 26471 2487
rect 26471 2453 26639 2487
rect 26639 2453 26640 2487
rect 26470 2379 26640 2453
rect 26470 2345 26471 2379
rect 26471 2345 26639 2379
rect 26639 2345 26640 2379
rect 26470 2344 26640 2345
rect 26842 2487 27012 2488
rect 26842 2453 26843 2487
rect 26843 2453 27011 2487
rect 27011 2453 27012 2487
rect 26842 2379 27012 2453
rect 26842 2345 26843 2379
rect 26843 2345 27011 2379
rect 27011 2345 27012 2379
rect 26842 2344 27012 2345
rect 27214 2487 27384 2488
rect 27214 2453 27215 2487
rect 27215 2453 27383 2487
rect 27383 2453 27384 2487
rect 27214 2379 27384 2453
rect 27214 2345 27215 2379
rect 27215 2345 27383 2379
rect 27383 2345 27384 2379
rect 27214 2344 27384 2345
rect 27586 2487 27756 2488
rect 27586 2453 27587 2487
rect 27587 2453 27755 2487
rect 27755 2453 27756 2487
rect 27586 2379 27756 2453
rect 27586 2345 27587 2379
rect 27587 2345 27755 2379
rect 27755 2345 27756 2379
rect 27586 2344 27756 2345
rect 27958 2487 28128 2488
rect 27958 2453 27959 2487
rect 27959 2453 28127 2487
rect 28127 2453 28128 2487
rect 27958 2379 28128 2453
rect 27958 2345 27959 2379
rect 27959 2345 28127 2379
rect 28127 2345 28128 2379
rect 27958 2344 28128 2345
rect 28330 2487 28500 2488
rect 28330 2453 28331 2487
rect 28331 2453 28499 2487
rect 28499 2453 28500 2487
rect 28330 2379 28500 2453
rect 28330 2345 28331 2379
rect 28331 2345 28499 2379
rect 28499 2345 28500 2379
rect 28330 2344 28500 2345
rect 28702 2487 28872 2488
rect 28702 2453 28703 2487
rect 28703 2453 28871 2487
rect 28871 2453 28872 2487
rect 28702 2379 28872 2453
rect 28702 2345 28703 2379
rect 28703 2345 28871 2379
rect 28871 2345 28872 2379
rect 28702 2344 28872 2345
rect 29074 2487 29244 2488
rect 29074 2453 29075 2487
rect 29075 2453 29243 2487
rect 29243 2453 29244 2487
rect 29074 2379 29244 2453
rect 29074 2345 29075 2379
rect 29075 2345 29243 2379
rect 29243 2345 29244 2379
rect 29074 2344 29244 2345
rect 29446 2487 29616 2488
rect 29446 2453 29447 2487
rect 29447 2453 29615 2487
rect 29615 2453 29616 2487
rect 29446 2379 29616 2453
rect 29446 2345 29447 2379
rect 29447 2345 29615 2379
rect 29615 2345 29616 2379
rect 29446 2344 29616 2345
rect 20890 2069 21060 2080
rect 20890 2035 20891 2069
rect 20891 2035 21059 2069
rect 21059 2035 21060 2069
rect 20890 2024 21060 2035
rect 21262 2069 21432 2080
rect 21262 2035 21263 2069
rect 21263 2035 21431 2069
rect 21431 2035 21432 2069
rect 21262 2024 21432 2035
rect 21634 2069 21804 2080
rect 21634 2035 21635 2069
rect 21635 2035 21803 2069
rect 21803 2035 21804 2069
rect 21634 2024 21804 2035
rect 22006 2069 22176 2080
rect 22006 2035 22007 2069
rect 22007 2035 22175 2069
rect 22175 2035 22176 2069
rect 22006 2024 22176 2035
rect 22378 2069 22548 2080
rect 22378 2035 22379 2069
rect 22379 2035 22547 2069
rect 22547 2035 22548 2069
rect 22378 2024 22548 2035
rect 22750 2069 22920 2080
rect 22750 2035 22751 2069
rect 22751 2035 22919 2069
rect 22919 2035 22920 2069
rect 22750 2024 22920 2035
rect 23122 2069 23292 2080
rect 23122 2035 23123 2069
rect 23123 2035 23291 2069
rect 23291 2035 23292 2069
rect 23122 2024 23292 2035
rect 23494 2069 23664 2080
rect 23494 2035 23495 2069
rect 23495 2035 23663 2069
rect 23663 2035 23664 2069
rect 23494 2024 23664 2035
rect 23866 2069 24036 2080
rect 23866 2035 23867 2069
rect 23867 2035 24035 2069
rect 24035 2035 24036 2069
rect 23866 2024 24036 2035
rect 24238 2069 24408 2080
rect 24238 2035 24239 2069
rect 24239 2035 24407 2069
rect 24407 2035 24408 2069
rect 24238 2024 24408 2035
rect 24610 2069 24780 2080
rect 24610 2035 24611 2069
rect 24611 2035 24779 2069
rect 24779 2035 24780 2069
rect 24610 2024 24780 2035
rect 24982 2069 25152 2080
rect 24982 2035 24983 2069
rect 24983 2035 25151 2069
rect 25151 2035 25152 2069
rect 24982 2024 25152 2035
rect 25354 2069 25524 2080
rect 25354 2035 25355 2069
rect 25355 2035 25523 2069
rect 25523 2035 25524 2069
rect 25354 2024 25524 2035
rect 25726 2069 25896 2080
rect 25726 2035 25727 2069
rect 25727 2035 25895 2069
rect 25895 2035 25896 2069
rect 25726 2024 25896 2035
rect 26098 2069 26268 2080
rect 26098 2035 26099 2069
rect 26099 2035 26267 2069
rect 26267 2035 26268 2069
rect 26098 2024 26268 2035
rect 26470 2069 26640 2080
rect 26470 2035 26471 2069
rect 26471 2035 26639 2069
rect 26639 2035 26640 2069
rect 26470 2024 26640 2035
rect 26842 2069 27012 2080
rect 26842 2035 26843 2069
rect 26843 2035 27011 2069
rect 27011 2035 27012 2069
rect 26842 2024 27012 2035
rect 27214 2069 27384 2080
rect 27214 2035 27215 2069
rect 27215 2035 27383 2069
rect 27383 2035 27384 2069
rect 27214 2024 27384 2035
rect 27586 2069 27756 2080
rect 27586 2035 27587 2069
rect 27587 2035 27755 2069
rect 27755 2035 27756 2069
rect 27586 2024 27756 2035
rect 27958 2069 28128 2080
rect 27958 2035 27959 2069
rect 27959 2035 28127 2069
rect 28127 2035 28128 2069
rect 27958 2024 28128 2035
rect 28330 2069 28500 2080
rect 28330 2035 28331 2069
rect 28331 2035 28499 2069
rect 28499 2035 28500 2069
rect 28330 2024 28500 2035
rect 28702 2069 28872 2080
rect 28702 2035 28703 2069
rect 28703 2035 28871 2069
rect 28871 2035 28872 2069
rect 28702 2024 28872 2035
rect 29074 2069 29244 2080
rect 29074 2035 29075 2069
rect 29075 2035 29243 2069
rect 29243 2035 29244 2069
rect 29074 2024 29244 2035
rect 29446 2069 29616 2080
rect 29446 2035 29447 2069
rect 29447 2035 29615 2069
rect 29615 2035 29616 2069
rect 29446 2024 29616 2035
rect 20710 1670 20910 1870
rect 21434 1670 21634 1870
rect 22178 1670 22378 1870
rect 22922 1670 23122 1870
rect 23666 1670 23866 1870
rect 24410 1670 24610 1870
rect 25154 1670 25354 1870
rect 25898 1670 26098 1870
rect 26642 1670 26842 1870
rect 27386 1670 27586 1870
rect 28130 1670 28330 1870
rect 28874 1670 29074 1870
rect 29618 1670 29818 1870
<< metal2 >>
rect 19572 11116 19772 11126
rect 19572 10906 19772 10916
rect 20316 11116 20516 11126
rect 20316 10906 20516 10916
rect 21060 11116 21260 11126
rect 21060 10906 21260 10916
rect 21804 11116 22004 11126
rect 21804 10906 22004 10916
rect 22548 11116 22748 11126
rect 22548 10906 22748 10916
rect 23292 11116 23492 11126
rect 23292 10906 23492 10916
rect 24036 11116 24236 11126
rect 24036 10906 24236 10916
rect 24780 11116 24980 11126
rect 24780 10906 24980 10916
rect 25152 11116 25352 11126
rect 25152 10906 25352 10916
rect 25896 11116 26096 11126
rect 25896 10906 26096 10916
rect 26640 11116 26840 11126
rect 26640 10906 26840 10916
rect 27384 11116 27584 11126
rect 27384 10906 27584 10916
rect 28128 11116 28328 11126
rect 28128 10906 28328 10916
rect 28872 11116 29072 11126
rect 28872 10906 29072 10916
rect 29616 11116 29816 11126
rect 29616 10906 29816 10916
rect 30360 11116 30560 11126
rect 30360 10906 30560 10916
rect 31104 11116 31304 11126
rect 31104 10906 31304 10916
rect 19402 10728 31114 10738
rect 19572 10668 19774 10728
rect 19944 10668 20146 10728
rect 20316 10668 20518 10728
rect 20688 10668 20890 10728
rect 21060 10668 21262 10728
rect 21432 10668 21634 10728
rect 21804 10668 22006 10728
rect 22176 10668 22378 10728
rect 22548 10668 22750 10728
rect 22920 10668 23122 10728
rect 23292 10668 23494 10728
rect 23664 10668 23866 10728
rect 24036 10668 24238 10728
rect 24408 10668 24610 10728
rect 24780 10668 24982 10728
rect 25152 10668 25354 10728
rect 25524 10668 25726 10728
rect 25896 10668 26098 10728
rect 26268 10668 26470 10728
rect 26640 10668 26842 10728
rect 27012 10668 27214 10728
rect 27384 10668 27586 10728
rect 27756 10668 27958 10728
rect 28128 10668 28330 10728
rect 28500 10668 28702 10728
rect 28872 10668 29074 10728
rect 29244 10668 29446 10728
rect 29616 10668 29818 10728
rect 29988 10668 30190 10728
rect 30360 10668 30562 10728
rect 30732 10668 30934 10728
rect 31104 10668 31114 10728
rect 19402 10658 31114 10668
rect 19402 10188 31104 10198
rect 19572 10044 19774 10188
rect 19944 10044 20146 10188
rect 20316 10044 20518 10188
rect 20688 10044 20890 10188
rect 21060 10044 21262 10188
rect 21432 10044 21634 10188
rect 21804 10044 22006 10188
rect 22176 10044 22378 10188
rect 22548 10044 22750 10188
rect 22920 10044 23122 10188
rect 23292 10044 23494 10188
rect 23664 10044 23866 10188
rect 24036 10044 24238 10188
rect 24408 10044 24610 10188
rect 24780 10044 24982 10188
rect 25152 10044 25354 10188
rect 25524 10044 25726 10188
rect 25896 10044 26098 10188
rect 26268 10044 26470 10188
rect 26640 10044 26842 10188
rect 27012 10044 27214 10188
rect 27384 10044 27586 10188
rect 27756 10044 27958 10188
rect 28128 10044 28330 10188
rect 28500 10044 28702 10188
rect 28872 10044 29074 10188
rect 29244 10044 29446 10188
rect 29616 10044 29818 10188
rect 29988 10044 30190 10188
rect 30360 10044 30562 10188
rect 30732 10044 30934 10188
rect 19402 10034 31104 10044
rect 19402 9552 31104 9562
rect 19572 9408 19774 9552
rect 19944 9408 20146 9552
rect 20316 9408 20518 9552
rect 20688 9408 20890 9552
rect 21060 9408 21262 9552
rect 21432 9408 21634 9552
rect 21804 9408 22006 9552
rect 22176 9408 22378 9552
rect 22548 9408 22750 9552
rect 22920 9408 23122 9552
rect 23292 9408 23494 9552
rect 23664 9408 23866 9552
rect 24036 9408 24238 9552
rect 24408 9408 24610 9552
rect 24780 9408 24982 9552
rect 25152 9408 25354 9552
rect 25524 9408 25726 9552
rect 25896 9408 26098 9552
rect 26268 9408 26470 9552
rect 26640 9408 26842 9552
rect 27012 9408 27214 9552
rect 27384 9408 27586 9552
rect 27756 9408 27958 9552
rect 28128 9408 28330 9552
rect 28500 9408 28702 9552
rect 28872 9408 29074 9552
rect 29244 9408 29446 9552
rect 29616 9408 29818 9552
rect 29988 9408 30190 9552
rect 30360 9408 30562 9552
rect 30732 9408 30934 9552
rect 19402 9398 31104 9408
rect 19402 8928 31104 8938
rect 19572 8868 19774 8928
rect 19944 8868 20146 8928
rect 20316 8868 20518 8928
rect 20688 8868 20890 8928
rect 21060 8868 21262 8928
rect 21432 8868 21634 8928
rect 21804 8868 22006 8928
rect 22176 8868 22378 8928
rect 22548 8868 22750 8928
rect 22920 8868 23122 8928
rect 23292 8868 23494 8928
rect 23664 8868 23866 8928
rect 24036 8868 24238 8928
rect 24408 8868 24610 8928
rect 24780 8868 24982 8928
rect 25152 8868 25354 8928
rect 25524 8868 25726 8928
rect 25896 8868 26098 8928
rect 26268 8868 26470 8928
rect 26640 8868 26842 8928
rect 27012 8868 27214 8928
rect 27384 8868 27586 8928
rect 27756 8868 27958 8928
rect 28128 8868 28330 8928
rect 28500 8868 28702 8928
rect 28872 8868 29074 8928
rect 29244 8868 29446 8928
rect 29616 8868 29818 8928
rect 29988 8868 30190 8928
rect 30360 8868 30562 8928
rect 30732 8868 30934 8928
rect 19402 8858 31104 8868
rect 20410 8442 23478 8540
rect 21076 8352 21246 8442
rect 23308 8352 23478 8442
rect 20890 8342 21432 8352
rect 21060 8278 21262 8342
rect 20890 8268 21432 8278
rect 21634 8342 22920 8352
rect 21804 8278 22006 8342
rect 22176 8278 22378 8342
rect 22548 8278 22750 8342
rect 21634 8268 22920 8278
rect 23122 8342 23664 8352
rect 23292 8278 23494 8342
rect 23122 8268 23664 8278
rect 21134 7410 21188 8268
rect 21878 7410 21932 8268
rect 22622 7410 22676 8268
rect 23366 7410 23420 8268
rect 20890 7400 21432 7410
rect 21060 7256 21262 7400
rect 20890 7246 21432 7256
rect 21634 7400 22920 7410
rect 21804 7256 22006 7400
rect 22176 7256 22378 7400
rect 22548 7256 22750 7400
rect 21634 7246 22920 7256
rect 23122 7400 23664 7410
rect 23292 7256 23494 7400
rect 23122 7246 23664 7256
rect 21134 6374 21188 7246
rect 21878 6374 21932 7246
rect 22622 6374 22676 7246
rect 23366 6374 23420 7246
rect 20890 6364 21432 6374
rect 21060 6220 21262 6364
rect 20890 6210 21432 6220
rect 21634 6364 22920 6374
rect 21804 6220 22006 6364
rect 22176 6220 22378 6364
rect 22548 6220 22750 6364
rect 21634 6210 22920 6220
rect 23122 6364 23664 6374
rect 23292 6220 23494 6364
rect 23122 6210 23664 6220
rect 21134 5338 21188 6210
rect 21878 5338 21932 6210
rect 22622 5338 22676 6210
rect 23366 5338 23420 6210
rect 20890 5328 21432 5338
rect 21060 5184 21262 5328
rect 20890 5174 21432 5184
rect 21634 5328 22920 5338
rect 21804 5184 22006 5328
rect 22176 5184 22378 5328
rect 22548 5184 22750 5328
rect 21634 5174 22920 5184
rect 23122 5328 23664 5338
rect 23292 5184 23494 5328
rect 23122 5174 23664 5184
rect 21134 4312 21188 5174
rect 21878 4312 21932 5174
rect 22622 4312 22676 5174
rect 23366 4312 23420 5174
rect 20890 4302 21432 4312
rect 21060 4248 21262 4302
rect 20890 4238 21432 4248
rect 21634 4302 22920 4312
rect 21804 4248 22006 4302
rect 22176 4248 22378 4302
rect 22548 4248 22750 4302
rect 21634 4238 22920 4248
rect 23122 4302 23664 4312
rect 23292 4248 23494 4302
rect 23122 4238 23664 4248
rect 21820 4138 21990 4238
rect 22564 4138 22734 4238
rect 20410 4040 22734 4138
rect 21870 3962 23850 3972
rect 22684 3782 23850 3962
rect 21870 3772 23850 3782
rect 23724 3654 23850 3772
rect 20890 3644 23676 3654
rect 21060 3588 21262 3644
rect 21432 3588 21634 3644
rect 21804 3588 22006 3644
rect 22176 3588 22378 3644
rect 22548 3588 22750 3644
rect 22920 3588 23122 3644
rect 23292 3588 23494 3644
rect 23664 3588 23676 3644
rect 20890 3578 23676 3588
rect 23724 3644 29616 3654
rect 23724 3588 23866 3644
rect 24036 3588 24238 3644
rect 24408 3588 24610 3644
rect 24780 3588 24982 3644
rect 25152 3588 25354 3644
rect 25524 3588 25726 3644
rect 25896 3588 26098 3644
rect 26268 3588 26470 3644
rect 26640 3588 26842 3644
rect 27012 3588 27214 3644
rect 27384 3588 27586 3644
rect 27756 3588 27958 3644
rect 28128 3588 28330 3644
rect 28500 3588 28702 3644
rect 28872 3588 29074 3644
rect 29244 3588 29446 3644
rect 23724 3578 29616 3588
rect 23724 3334 23850 3578
rect 20890 3324 23676 3334
rect 21060 3180 21262 3324
rect 21432 3180 21634 3324
rect 21804 3180 22006 3324
rect 22176 3180 22378 3324
rect 22548 3180 22750 3324
rect 22920 3180 23122 3324
rect 23292 3180 23494 3324
rect 23664 3180 23676 3324
rect 20890 3170 23676 3180
rect 23724 3324 29616 3334
rect 23724 3180 23866 3324
rect 24036 3180 24238 3324
rect 24408 3180 24610 3324
rect 24780 3180 24982 3324
rect 25152 3180 25354 3324
rect 25524 3180 25726 3324
rect 25896 3180 26098 3324
rect 26268 3180 26470 3324
rect 26640 3180 26842 3324
rect 27012 3180 27214 3324
rect 27384 3180 27586 3324
rect 27756 3180 27958 3324
rect 28128 3180 28330 3324
rect 28500 3180 28702 3324
rect 28872 3180 29074 3324
rect 29244 3180 29446 3324
rect 23724 3170 29616 3180
rect 23724 2916 23850 3170
rect 20890 2906 23676 2916
rect 21060 2762 21262 2906
rect 21432 2762 21634 2906
rect 21804 2762 22006 2906
rect 22176 2762 22378 2906
rect 22548 2762 22750 2906
rect 22920 2762 23122 2906
rect 23292 2762 23494 2906
rect 23664 2762 23676 2906
rect 20890 2752 23676 2762
rect 23724 2906 29616 2916
rect 23724 2762 23866 2906
rect 24036 2762 24238 2906
rect 24408 2762 24610 2906
rect 24780 2762 24982 2906
rect 25152 2762 25354 2906
rect 25524 2762 25726 2906
rect 25896 2762 26098 2906
rect 26268 2762 26470 2906
rect 26640 2762 26842 2906
rect 27012 2762 27214 2906
rect 27384 2762 27586 2906
rect 27756 2762 27958 2906
rect 28128 2762 28330 2906
rect 28500 2762 28702 2906
rect 28872 2762 29074 2906
rect 29244 2762 29446 2906
rect 23724 2752 29616 2762
rect 23724 2498 23850 2752
rect 20890 2488 23676 2498
rect 21060 2344 21262 2488
rect 21432 2344 21634 2488
rect 21804 2344 22006 2488
rect 22176 2344 22378 2488
rect 22548 2344 22750 2488
rect 22920 2344 23122 2488
rect 23292 2344 23494 2488
rect 23664 2344 23676 2488
rect 20890 2334 23676 2344
rect 23724 2488 29616 2498
rect 23724 2344 23866 2488
rect 24036 2344 24238 2488
rect 24408 2344 24610 2488
rect 24780 2344 24982 2488
rect 25152 2344 25354 2488
rect 25524 2344 25726 2488
rect 25896 2344 26098 2488
rect 26268 2344 26470 2488
rect 26640 2344 26842 2488
rect 27012 2344 27214 2488
rect 27384 2344 27586 2488
rect 27756 2344 27958 2488
rect 28128 2344 28330 2488
rect 28500 2344 28702 2488
rect 28872 2344 29074 2488
rect 29244 2344 29446 2488
rect 23724 2334 29616 2344
rect 23724 2090 23850 2334
rect 20890 2080 23676 2090
rect 21060 2024 21262 2080
rect 21432 2024 21634 2080
rect 21804 2024 22006 2080
rect 22176 2024 22378 2080
rect 22548 2024 22750 2080
rect 22920 2024 23122 2080
rect 23292 2024 23494 2080
rect 23664 2024 23676 2080
rect 20890 2014 23676 2024
rect 23724 2080 29616 2090
rect 23724 2024 23866 2080
rect 24036 2024 24238 2080
rect 24408 2024 24610 2080
rect 24780 2024 24982 2080
rect 25152 2024 25354 2080
rect 25524 2024 25726 2080
rect 25896 2024 26098 2080
rect 26268 2024 26470 2080
rect 26640 2024 26842 2080
rect 27012 2024 27214 2080
rect 27384 2024 27586 2080
rect 27756 2024 27958 2080
rect 28128 2024 28330 2080
rect 28500 2024 28702 2080
rect 28872 2024 29074 2080
rect 29244 2024 29446 2080
rect 23724 2014 29616 2024
rect 20710 1870 20910 1880
rect 20710 1660 20910 1670
rect 21434 1870 21634 1880
rect 21434 1660 21634 1670
rect 22178 1870 22378 1880
rect 22178 1660 22378 1670
rect 22922 1870 23122 1880
rect 22922 1660 23122 1670
rect 23666 1870 23866 1880
rect 23666 1660 23866 1670
rect 24410 1870 24610 1880
rect 24410 1660 24610 1670
rect 25154 1870 25354 1880
rect 25154 1660 25354 1670
rect 25898 1870 26098 1880
rect 25898 1660 26098 1670
rect 26642 1870 26842 1880
rect 26642 1660 26842 1670
rect 27386 1870 27586 1880
rect 27386 1660 27586 1670
rect 28130 1870 28330 1880
rect 28130 1660 28330 1670
rect 28874 1870 29074 1880
rect 28874 1660 29074 1670
rect 29618 1870 29818 1880
rect 29618 1660 29818 1670
<< via2 >>
rect 19572 10916 19772 11116
rect 20316 10916 20516 11116
rect 21060 10916 21260 11116
rect 21804 10916 22004 11116
rect 22548 10916 22748 11116
rect 23292 10916 23492 11116
rect 24036 10916 24236 11116
rect 24780 10916 24980 11116
rect 25152 10916 25352 11116
rect 25896 10916 26096 11116
rect 26640 10916 26840 11116
rect 27384 10916 27584 11116
rect 28128 10916 28328 11116
rect 28872 10916 29072 11116
rect 29616 10916 29816 11116
rect 30360 10916 30560 11116
rect 31104 10916 31304 11116
rect 20710 1670 20910 1870
rect 21434 1670 21634 1870
rect 22178 1670 22378 1870
rect 22922 1670 23122 1870
rect 23666 1670 23866 1870
rect 24410 1670 24610 1870
rect 25154 1670 25354 1870
rect 25898 1670 26098 1870
rect 26642 1670 26842 1870
rect 27386 1670 27586 1870
rect 28130 1670 28330 1870
rect 28874 1670 29074 1870
rect 29618 1670 29818 1870
<< metal3 >>
rect 19562 11116 19782 11121
rect 19562 10916 19572 11116
rect 19772 10916 19782 11116
rect 19562 10911 19782 10916
rect 20306 11116 20526 11121
rect 20306 10916 20316 11116
rect 20516 10916 20526 11116
rect 20306 10911 20526 10916
rect 21050 11116 21270 11121
rect 21050 10916 21060 11116
rect 21260 10916 21270 11116
rect 21050 10911 21270 10916
rect 21794 11116 22014 11121
rect 21794 10916 21804 11116
rect 22004 10916 22014 11116
rect 21794 10911 22014 10916
rect 22538 11116 22758 11121
rect 22538 10916 22548 11116
rect 22748 10916 22758 11116
rect 22538 10911 22758 10916
rect 23282 11116 23502 11121
rect 23282 10916 23292 11116
rect 23492 10916 23502 11116
rect 23282 10911 23502 10916
rect 24026 11116 24246 11121
rect 24026 10916 24036 11116
rect 24236 10916 24246 11116
rect 24026 10911 24246 10916
rect 24770 11116 24990 11121
rect 24770 10916 24780 11116
rect 24980 10916 24990 11116
rect 24770 10911 24990 10916
rect 25142 11116 25362 11121
rect 25142 10916 25152 11116
rect 25352 10916 25362 11116
rect 25142 10911 25362 10916
rect 25886 11116 26106 11121
rect 25886 10916 25896 11116
rect 26096 10916 26106 11116
rect 25886 10911 26106 10916
rect 26630 11116 26850 11121
rect 26630 10916 26640 11116
rect 26840 10916 26850 11116
rect 26630 10911 26850 10916
rect 27374 11116 27594 11121
rect 27374 10916 27384 11116
rect 27584 10916 27594 11116
rect 27374 10911 27594 10916
rect 28118 11116 28338 11121
rect 28118 10916 28128 11116
rect 28328 10916 28338 11116
rect 28118 10911 28338 10916
rect 28862 11116 29082 11121
rect 28862 10916 28872 11116
rect 29072 10916 29082 11116
rect 28862 10911 29082 10916
rect 29606 11116 29826 11121
rect 29606 10916 29616 11116
rect 29816 10916 29826 11116
rect 29606 10911 29826 10916
rect 30350 11116 30570 11121
rect 30350 10916 30360 11116
rect 30560 10916 30570 11116
rect 30350 10911 30570 10916
rect 31094 11116 31314 11121
rect 31094 10916 31104 11116
rect 31304 10916 31314 11116
rect 31094 10911 31314 10916
rect 20700 1870 20920 1875
rect 20700 1670 20710 1870
rect 20910 1670 20920 1870
rect 20700 1665 20920 1670
rect 21424 1870 21644 1875
rect 21424 1670 21434 1870
rect 21634 1670 21644 1870
rect 21424 1665 21644 1670
rect 22168 1870 22388 1875
rect 22168 1670 22178 1870
rect 22378 1670 22388 1870
rect 22168 1665 22388 1670
rect 22912 1870 23132 1875
rect 22912 1670 22922 1870
rect 23122 1670 23132 1870
rect 22912 1665 23132 1670
rect 23656 1870 23876 1875
rect 23656 1670 23666 1870
rect 23866 1670 23876 1870
rect 23656 1665 23876 1670
rect 24400 1870 24620 1875
rect 24400 1670 24410 1870
rect 24610 1670 24620 1870
rect 24400 1665 24620 1670
rect 25144 1870 25364 1875
rect 25144 1670 25154 1870
rect 25354 1670 25364 1870
rect 25144 1665 25364 1670
rect 25888 1870 26108 1875
rect 25888 1670 25898 1870
rect 26098 1670 26108 1870
rect 25888 1665 26108 1670
rect 26632 1870 26852 1875
rect 26632 1670 26642 1870
rect 26842 1670 26852 1870
rect 26632 1665 26852 1670
rect 27376 1870 27596 1875
rect 27376 1670 27386 1870
rect 27586 1670 27596 1870
rect 27376 1665 27596 1670
rect 28120 1870 28340 1875
rect 28120 1670 28130 1870
rect 28330 1670 28340 1870
rect 28120 1665 28340 1670
rect 28864 1870 29084 1875
rect 28864 1670 28874 1870
rect 29074 1670 29084 1870
rect 28864 1665 29084 1670
rect 29608 1870 29828 1875
rect 29608 1670 29618 1870
rect 29818 1670 29828 1870
rect 29608 1665 29828 1670
<< via3 >>
rect 19572 10916 19772 11116
rect 20316 10916 20516 11116
rect 21060 10916 21260 11116
rect 21804 10916 22004 11116
rect 22548 10916 22748 11116
rect 23292 10916 23492 11116
rect 24036 10916 24236 11116
rect 24780 10916 24980 11116
rect 25152 10916 25352 11116
rect 25896 10916 26096 11116
rect 26640 10916 26840 11116
rect 27384 10916 27584 11116
rect 28128 10916 28328 11116
rect 28872 10916 29072 11116
rect 29616 10916 29816 11116
rect 30360 10916 30560 11116
rect 31104 10916 31304 11116
rect 20710 1670 20910 1870
rect 21434 1670 21634 1870
rect 22178 1670 22378 1870
rect 22922 1670 23122 1870
rect 23666 1670 23866 1870
rect 24410 1670 24610 1870
rect 25154 1670 25354 1870
rect 25898 1670 26098 1870
rect 26642 1670 26842 1870
rect 27386 1670 27586 1870
rect 28130 1670 28330 1870
rect 28874 1670 29074 1870
rect 29618 1670 29818 1870
<< metal4 >>
rect 18966 11116 31490 11894
rect 18966 10916 19572 11116
rect 19772 10916 20316 11116
rect 20516 10916 21060 11116
rect 21260 10916 21804 11116
rect 22004 10916 22548 11116
rect 22748 10916 23292 11116
rect 23492 10916 24036 11116
rect 24236 10916 24780 11116
rect 24980 10916 25152 11116
rect 25352 10916 25896 11116
rect 26096 10916 26640 11116
rect 26840 10916 27384 11116
rect 27584 10916 28128 11116
rect 28328 10916 28872 11116
rect 29072 10916 29616 11116
rect 29816 10916 30360 11116
rect 30560 10916 31104 11116
rect 31304 10916 31490 11116
rect 18966 10890 31490 10916
rect 18966 1870 31490 1894
rect 18966 1670 20710 1870
rect 20910 1670 21434 1870
rect 21634 1670 22178 1870
rect 22378 1670 22922 1870
rect 23122 1670 23666 1870
rect 23866 1670 24410 1870
rect 24610 1670 25154 1870
rect 25354 1670 25898 1870
rect 26098 1670 26642 1870
rect 26842 1670 27386 1870
rect 27586 1670 28130 1870
rect 28330 1670 28874 1870
rect 29074 1670 29618 1870
rect 29818 1670 31490 1870
rect 18966 890 31490 1670
<< labels >>
flabel metal4 20162 11568 20162 11568 0 FreeSans 8000 0 0 0 vdd
port 0 nsew
flabel metal4 19728 1054 19728 1054 0 FreeSans 8000 0 0 0 vss
port 4 nsew
flabel metal2 20440 8472 20440 8472 0 FreeSans 8000 0 0 0 vn
port 2 nsew
flabel metal2 20476 4072 20476 4072 0 FreeSans 8000 0 0 0 vp
port 1 nsew
flabel metal1 19352 9472 19352 9472 0 FreeSans 8000 0 0 0 vbias
port 3 nsew
flabel metal1 27980 6420 27980 6420 0 FreeSans 8000 0 0 0 vout
port 5 nsew
<< end >>
