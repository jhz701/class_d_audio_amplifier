magic
tech sky130A
magscale 1 2
timestamp 1629295110
<< pwell >>
rect -4232 70922 -3540 70952
rect -68881 56799 -66685 59109
rect -68881 24641 -68774 24642
rect -68881 22331 -66685 24641
<< psubdiff >>
rect -68845 59039 -68749 59073
rect -66817 59039 -66721 59073
rect -68845 58977 -68811 59039
rect -66755 58977 -66721 59039
rect -68845 56869 -68811 56931
rect -66755 56869 -66721 56931
rect -68845 56835 -68749 56869
rect -66817 56835 -66721 56869
rect -68845 24605 -68774 24606
rect -68845 24571 -68749 24605
rect -66817 24571 -66721 24605
rect -68845 24510 -68811 24571
rect -66755 24509 -66721 24571
rect -68845 22402 -68811 22463
rect -68845 22401 -68774 22402
rect -66755 22401 -66721 22463
rect -68845 22367 -68749 22401
rect -66817 22367 -66721 22401
<< psubdiffcont >>
rect -68749 59039 -66817 59073
rect -68845 56931 -68811 58977
rect -66755 56931 -66721 58977
rect -68749 56835 -66817 56869
rect -68749 24571 -66817 24605
rect -68845 22463 -68811 24510
rect -66755 22463 -66721 24509
rect -68749 22367 -66817 22401
<< xpolycontact >>
rect -68715 58873 -68283 58943
rect -67283 58873 -66851 58943
rect -68715 58555 -68283 58625
rect -67283 58555 -66851 58625
rect -68715 58237 -68283 58307
rect -67283 58237 -66851 58307
rect -68715 57919 -68283 57989
rect -67283 57919 -66851 57989
rect -68715 57601 -68283 57671
rect -67283 57601 -66851 57671
rect -68715 57283 -68283 57353
rect -67283 57283 -66851 57353
rect -68715 56965 -68283 57035
rect -67283 56965 -66851 57035
rect -68715 24405 -68283 24475
rect -67283 24405 -66851 24475
rect -68715 24087 -68283 24157
rect -67283 24087 -66851 24157
rect -68715 23769 -68283 23839
rect -67283 23769 -66851 23839
rect -68715 23451 -68283 23521
rect -67283 23451 -66851 23521
rect -68715 23133 -68283 23203
rect -67283 23133 -66851 23203
rect -68715 22815 -68283 22885
rect -67283 22815 -66851 22885
rect -68715 22497 -68283 22567
rect -67283 22497 -66851 22567
<< xpolyres >>
rect -68283 58873 -67283 58943
rect -68283 58555 -67283 58625
rect -68283 58237 -67283 58307
rect -68283 57919 -67283 57989
rect -68283 57601 -67283 57671
rect -68283 57283 -67283 57353
rect -68283 56965 -67283 57035
rect -68283 24405 -67283 24475
rect -68283 24087 -67283 24157
rect -68283 23769 -67283 23839
rect -68283 23451 -67283 23521
rect -68283 23133 -67283 23203
rect -68283 22815 -67283 22885
rect -68283 22497 -67283 22567
<< locali >>
rect -68845 59039 -68749 59073
rect -66817 59039 -66721 59073
rect -68845 58977 -68811 59039
rect -66755 58977 -66721 59039
rect -68845 56869 -68811 56931
rect -66755 56869 -66721 56931
rect -68845 56835 -68749 56869
rect -66817 56835 -66721 56869
rect -68845 24605 -68774 24606
rect -68845 24571 -68749 24605
rect -66817 24571 -66721 24605
rect -68845 24510 -68811 24571
rect -66755 24509 -66721 24571
rect -68845 22402 -68811 22463
rect -68845 22401 -68774 22402
rect -66755 22401 -66721 22463
rect -68845 22367 -68749 22401
rect -66817 22367 -66721 22401
<< viali >>
rect -68697 58889 -68300 58927
rect -67266 58889 -66869 58927
rect -68862 58542 -68845 58612
rect -68845 58542 -68811 58612
rect -68811 58542 -68792 58612
rect -68697 58571 -68300 58609
rect -67266 58571 -66869 58609
rect -68697 58253 -68300 58291
rect -67266 58253 -66869 58291
rect -68862 58142 -68845 58212
rect -68845 58142 -68811 58212
rect -68811 58142 -68792 58212
rect -68697 57935 -68300 57973
rect -67266 57935 -66869 57973
rect -68862 57742 -68845 57812
rect -68845 57742 -68811 57812
rect -68811 57742 -68792 57812
rect -68697 57617 -68300 57655
rect -67266 57617 -66869 57655
rect -68862 57342 -68845 57412
rect -68845 57342 -68811 57412
rect -68811 57342 -68792 57412
rect -68697 57299 -68300 57337
rect -67266 57299 -66869 57337
rect -68862 56942 -68845 57012
rect -68845 56942 -68811 57012
rect -68811 56942 -68792 57012
rect -68697 56981 -68300 57019
rect -67266 56981 -66869 57019
rect -68862 24429 -68845 24499
rect -68845 24429 -68811 24499
rect -68811 24429 -68792 24499
rect -68697 24421 -68300 24459
rect -67266 24421 -66869 24459
rect -68697 24103 -68300 24141
rect -68862 24029 -68845 24099
rect -68845 24029 -68811 24099
rect -68811 24029 -68792 24099
rect -67266 24103 -66869 24141
rect -68697 23785 -68300 23823
rect -67266 23785 -66869 23823
rect -68862 23629 -68845 23699
rect -68845 23629 -68811 23699
rect -68811 23629 -68792 23699
rect -68697 23467 -68300 23505
rect -67266 23467 -66869 23505
rect -68862 23229 -68845 23299
rect -68845 23229 -68811 23299
rect -68811 23229 -68792 23299
rect -68697 23149 -68300 23187
rect -67266 23149 -66869 23187
rect -68862 22829 -68845 22899
rect -68845 22829 -68811 22899
rect -68811 22829 -68792 22899
rect -68697 22831 -68300 22869
rect -67266 22831 -66869 22869
rect -68697 22513 -68300 22551
rect -67266 22513 -66869 22551
<< metal1 >>
rect 1326 68986 1336 70952
rect 2712 68986 2722 70952
rect -65934 64918 -65898 65052
rect -49854 64934 -49824 65074
rect -68716 63090 -68246 63712
rect -68716 58927 -68282 63090
rect -41240 61932 -41112 62038
rect -23170 61932 -23130 62038
rect -41240 61088 -23130 61932
rect -41112 60982 -23170 61088
rect -68716 58889 -68697 58927
rect -68300 58889 -68282 58927
rect -68716 58872 -68282 58889
rect -67284 58927 -66850 58944
rect -67284 58889 -67266 58927
rect -66869 58889 -66850 58927
rect -69500 58482 -69490 58682
rect -69290 58618 -69280 58682
rect -69290 58612 -68780 58618
rect -69290 58542 -68862 58612
rect -68792 58542 -68780 58612
rect -69290 58536 -68780 58542
rect -68716 58609 -68282 58626
rect -68716 58571 -68697 58609
rect -68300 58571 -68282 58609
rect -69290 58482 -69280 58536
rect -68716 58291 -68282 58571
rect -67284 58609 -66850 58889
rect -67284 58571 -67266 58609
rect -66869 58571 -66850 58609
rect -67284 58554 -66850 58571
rect -69500 58082 -69490 58282
rect -69290 58218 -69280 58282
rect -68716 58253 -68697 58291
rect -68300 58253 -68282 58291
rect -68716 58236 -68282 58253
rect -67284 58291 -66850 58308
rect -67284 58253 -67266 58291
rect -66869 58253 -66850 58291
rect -69290 58212 -68780 58218
rect -69290 58142 -68862 58212
rect -68792 58142 -68780 58212
rect -69290 58136 -68780 58142
rect -69290 58082 -69280 58136
rect -68716 57973 -68282 57990
rect -68716 57935 -68697 57973
rect -68300 57935 -68282 57973
rect -69500 57682 -69490 57882
rect -69290 57818 -69280 57882
rect -69290 57812 -68780 57818
rect -69290 57742 -68862 57812
rect -68792 57742 -68780 57812
rect -69290 57736 -68780 57742
rect -69290 57682 -69280 57736
rect -68716 57655 -68282 57935
rect -67284 57973 -66850 58253
rect -67284 57935 -67266 57973
rect -66869 57935 -66850 57973
rect -67284 57918 -66850 57935
rect -68716 57617 -68697 57655
rect -68300 57617 -68282 57655
rect -68716 57600 -68282 57617
rect -67284 57655 -66850 57672
rect -67284 57617 -67266 57655
rect -66869 57617 -66850 57655
rect -69500 57282 -69490 57482
rect -69290 57418 -69280 57482
rect -69290 57412 -68780 57418
rect -69290 57342 -68862 57412
rect -68792 57342 -68780 57412
rect -69290 57336 -68780 57342
rect -68716 57337 -68282 57354
rect -69290 57282 -69280 57336
rect -68716 57299 -68697 57337
rect -68300 57299 -68282 57337
rect -69500 56882 -69490 57082
rect -69290 57018 -69280 57082
rect -68716 57019 -68282 57299
rect -67284 57337 -66850 57617
rect -67284 57299 -67266 57337
rect -66869 57299 -66850 57337
rect -67284 57282 -66850 57299
rect -69290 57012 -68780 57018
rect -69290 56942 -68862 57012
rect -68792 56942 -68780 57012
rect -68716 56981 -68697 57019
rect -68300 56981 -68282 57019
rect -68716 56964 -68282 56981
rect -67284 57019 -66850 57036
rect -67284 56981 -67266 57019
rect -66869 56981 -66850 57019
rect -69290 56936 -68780 56942
rect -69290 56882 -69280 56936
rect -67284 55404 -66850 56981
rect 2084 56656 2094 57440
rect 2858 56656 2868 57440
rect -67772 54436 -67762 55404
rect -66844 54436 -66834 55404
rect 2094 53520 2858 56656
rect -64550 43324 -64514 43476
rect -51022 43298 -50988 43410
rect -79996 42872 -79958 42992
rect -79996 39076 -79962 39198
rect -67772 26036 -67762 27004
rect -66844 26036 -66834 27004
rect -69500 24359 -69490 24559
rect -69290 24505 -69280 24559
rect -69290 24499 -68780 24505
rect -69290 24429 -68862 24499
rect -68792 24429 -68780 24499
rect -69290 24423 -68780 24429
rect -68716 24459 -68282 24476
rect -69290 24359 -69280 24423
rect -68716 24421 -68697 24459
rect -68300 24421 -68282 24459
rect -69500 23959 -69490 24159
rect -69290 24105 -69280 24159
rect -68716 24141 -68282 24421
rect -67284 24459 -66850 26036
rect 2094 24782 2858 28518
rect -67284 24421 -67266 24459
rect -66869 24421 -66850 24459
rect -67284 24404 -66850 24421
rect -69290 24099 -68780 24105
rect -69290 24029 -68862 24099
rect -68792 24029 -68780 24099
rect -68716 24103 -68697 24141
rect -68300 24103 -68282 24141
rect -68716 24086 -68282 24103
rect -67284 24141 -66850 24158
rect -67284 24103 -67266 24141
rect -66869 24103 -66850 24141
rect -69290 24023 -68780 24029
rect -69290 23959 -69280 24023
rect -68716 23823 -68282 23840
rect -68716 23785 -68697 23823
rect -68300 23785 -68282 23823
rect -69500 23559 -69490 23759
rect -69290 23705 -69280 23759
rect -69290 23699 -68780 23705
rect -69290 23629 -68862 23699
rect -68792 23629 -68780 23699
rect -69290 23623 -68780 23629
rect -69290 23559 -69280 23623
rect -68716 23505 -68282 23785
rect -67284 23823 -66850 24103
rect 2084 23998 2094 24782
rect 2858 23998 2868 24782
rect -67284 23785 -67266 23823
rect -66869 23785 -66850 23823
rect -67284 23768 -66850 23785
rect -68716 23467 -68697 23505
rect -68300 23467 -68282 23505
rect -68716 23450 -68282 23467
rect -67284 23505 -66850 23522
rect -67284 23467 -67266 23505
rect -66869 23467 -66850 23505
rect -69500 23159 -69490 23359
rect -69290 23305 -69280 23359
rect -69290 23299 -68780 23305
rect -69290 23229 -68862 23299
rect -68792 23229 -68780 23299
rect -69290 23223 -68780 23229
rect -69290 23159 -69280 23223
rect -68716 23187 -68282 23204
rect -68716 23149 -68697 23187
rect -68300 23149 -68282 23187
rect -69500 22759 -69490 22959
rect -69290 22905 -69280 22959
rect -69290 22899 -68780 22905
rect -69290 22829 -68862 22899
rect -68792 22829 -68780 22899
rect -69290 22823 -68780 22829
rect -68716 22869 -68282 23149
rect -67284 23187 -66850 23467
rect -67284 23149 -67266 23187
rect -66869 23149 -66850 23187
rect -67284 23132 -66850 23149
rect -68716 22831 -68697 22869
rect -68300 22831 -68282 22869
rect -69290 22759 -69280 22823
rect -68716 22814 -68282 22831
rect -67284 22869 -66850 22886
rect -67284 22831 -67266 22869
rect -66869 22831 -66850 22869
rect -68716 22551 -68282 22568
rect -68716 22513 -68697 22551
rect -68300 22513 -68282 22551
rect -68716 18350 -68282 22513
rect -67284 22551 -66850 22831
rect -67284 22513 -67266 22551
rect -66869 22513 -66850 22551
rect -67284 22496 -66850 22513
rect -41112 19506 -23170 20456
rect -68716 17728 -68238 18350
rect -67632 17728 -67622 18350
rect -68090 17682 -67814 17728
rect -65930 16348 -65896 16488
rect -49860 16330 -49830 16496
rect 1326 10486 1336 12452
rect 2712 10486 2722 12452
<< via1 >>
rect 1336 68986 2712 70952
rect -69490 58482 -69290 58682
rect -69490 58082 -69290 58282
rect -69490 57682 -69290 57882
rect -69490 57282 -69290 57482
rect -69490 56882 -69290 57082
rect 2094 56656 2858 57440
rect -67762 54436 -66844 55404
rect -67762 26036 -66844 27004
rect -69490 24359 -69290 24559
rect -69490 23959 -69290 24159
rect -69490 23559 -69290 23759
rect 2094 23998 2858 24782
rect -69490 23159 -69290 23359
rect -69490 22759 -69290 22959
rect -68238 17728 -67632 18350
rect 1336 10486 2712 12452
<< metal2 >>
rect 1336 70952 2712 70962
rect -4232 68986 1336 70952
rect 1336 68976 2712 68986
rect -84678 66636 -83760 66646
rect -83760 66116 -50150 66636
rect -84678 65658 -83760 65668
rect -50468 65102 -50150 66116
rect -50468 64938 -49614 65102
rect -83216 64872 -82298 64882
rect -82298 64302 -65686 64466
rect -83216 63894 -82298 63904
rect -50082 63572 -49434 63582
rect -49434 63346 -48746 63444
rect -50082 62888 -49434 62898
rect -50730 61118 -50082 61128
rect -50082 60574 -48710 60914
rect -50730 60434 -50082 60444
rect -81112 59480 -80194 59490
rect -80194 58944 -64790 59042
rect -48982 58944 -48710 60574
rect -81112 58502 -80194 58512
rect -69490 58682 -69290 58692
rect -69490 58472 -69290 58482
rect -69490 58282 -69290 58292
rect -69490 58072 -69290 58082
rect -69490 57882 -69290 57892
rect -69490 57672 -69290 57682
rect -69490 57482 -69290 57492
rect -69490 57272 -69290 57282
rect 2094 57440 2858 57450
rect -69490 57082 -69290 57092
rect -69490 56872 -69290 56882
rect -12924 56656 2094 57036
rect 2094 56646 2858 56656
rect -67762 55404 -66844 55414
rect -67762 54426 -66844 54436
rect -84680 46174 -83762 46184
rect -87618 45206 -84680 45388
rect -84680 45196 -83762 45206
rect -83188 44648 -82270 44658
rect -87618 44062 -83188 44244
rect -67752 44518 -50860 44676
rect -82270 44062 -82260 44244
rect -83188 43670 -82270 43680
rect -87618 43022 -80426 43100
rect -87618 42918 -79752 43022
rect -80618 42856 -79752 42918
rect -87626 41774 -82948 41956
rect -83148 41158 -82948 41774
rect -67752 41158 -67524 44518
rect -50958 43966 -50860 44518
rect -83148 40978 -67524 41158
rect -67184 42136 -64304 42216
rect -67184 40464 -66956 42136
rect -83148 40284 -66956 40464
rect -83148 39668 -82948 40284
rect -87620 39486 -82948 39668
rect -80618 38524 -79754 38584
rect -87618 38420 -79754 38524
rect -87618 38342 -80430 38420
rect -83184 37760 -82266 37770
rect -87618 37198 -83184 37380
rect -83184 36782 -82266 36792
rect -66306 37318 -63270 37416
rect -84678 36236 -83760 36246
rect -87618 36054 -84678 36236
rect -84678 35258 -83760 35268
rect -81112 33944 -80194 33954
rect -66306 33716 -66080 37318
rect -75540 33524 -66080 33716
rect -75540 33184 -75422 33524
rect -80194 33062 -78730 33160
rect -76604 33062 -75422 33184
rect -81112 32966 -80194 32976
rect -67762 27004 -66844 27014
rect -67762 26026 -66844 26036
rect 2094 24782 2858 24792
rect -69490 24559 -69290 24569
rect -12898 24402 2094 24782
rect -69490 24349 -69290 24359
rect -69490 24159 -69290 24169
rect 2094 23988 2858 23998
rect -69490 23949 -69290 23959
rect -69490 23759 -69290 23769
rect -69490 23549 -69290 23559
rect -69490 23359 -69290 23369
rect -69490 23149 -69290 23159
rect -69490 22959 -69290 22969
rect -81112 22944 -80194 22954
rect -69490 22749 -69290 22759
rect -80194 22398 -65138 22496
rect -48982 22398 -48644 22496
rect -81112 21966 -80194 21976
rect -50730 20996 -50082 21006
rect -48982 20866 -48710 22398
rect -50082 20526 -48710 20866
rect -50730 20312 -50082 20322
rect -49962 18554 -49314 18564
rect -68238 18350 -67632 18360
rect -67632 17996 -66650 18094
rect -49314 17994 -48716 18094
rect -49962 17870 -49314 17880
rect -68238 17718 -67632 17728
rect -83216 17566 -82298 17576
rect -82298 16974 -65686 17138
rect -83216 16588 -82298 16598
rect -50470 16338 -49616 16502
rect -84678 15772 -83760 15782
rect -50470 15324 -50152 16338
rect -83760 14804 -50152 15324
rect -84678 14794 -83760 14804
rect 1336 12452 2712 12462
rect -3792 10486 1336 12452
rect 1336 10476 2712 10486
<< via2 >>
rect -84678 65668 -83760 66636
rect -83216 63904 -82298 64872
rect -50082 62898 -49434 63572
rect -50730 60444 -50082 61118
rect -81112 58512 -80194 59480
rect -69490 58482 -69290 58682
rect -69490 58082 -69290 58282
rect -69490 57682 -69290 57882
rect -69490 57282 -69290 57482
rect -69490 56882 -69290 57082
rect -67762 54436 -66844 55404
rect -84680 45206 -83762 46174
rect -83188 43680 -82270 44648
rect -83184 36792 -82266 37760
rect -84678 35268 -83760 36236
rect -81112 32976 -80194 33944
rect -67762 26036 -66844 27004
rect -69490 24359 -69290 24559
rect -69490 23959 -69290 24159
rect -69490 23559 -69290 23759
rect -69490 23159 -69290 23359
rect -81112 21976 -80194 22944
rect -69490 22759 -69290 22959
rect -50730 20322 -50082 20996
rect -49962 17880 -49314 18554
rect -83216 16598 -82298 17566
rect -84678 14804 -83760 15772
<< metal3 >>
rect -2674 72970 -2664 74522
rect -1112 72970 -1102 74522
rect -84688 66636 -83750 66641
rect -84688 65668 -84678 66636
rect -83760 65668 -83750 66636
rect -84688 65663 -83750 65668
rect -92940 50526 -92930 51530
rect -92040 50526 -92030 51530
rect -92930 45936 -92040 50526
rect -84680 46179 -84016 65663
rect -83226 64872 -82288 64877
rect -83226 63904 -83216 64872
rect -82298 63904 -82288 64872
rect -83226 63899 -82288 63904
rect -84690 46174 -83752 46179
rect -84690 45206 -84680 46174
rect -83762 45206 -83752 46174
rect -84690 45201 -83752 45206
rect -82904 44653 -82542 63899
rect -50092 63572 -49424 63577
rect -50092 62898 -50082 63572
rect -49434 62898 -49424 63572
rect -50092 62893 -49424 62898
rect -50740 61118 -50072 61123
rect -50740 60444 -50730 61118
rect -50082 60444 -50072 61118
rect -50740 60439 -50072 60444
rect -81122 59480 -80184 59485
rect -81122 58512 -81112 59480
rect -80194 58512 -80184 59480
rect -81122 58507 -80184 58512
rect -69500 58682 -69280 58687
rect -83198 44648 -82260 44653
rect -83198 43680 -83188 44648
rect -82270 43680 -82260 44648
rect -83198 43675 -82260 43680
rect -83194 37760 -82256 37765
rect -83194 36792 -83184 37760
rect -82266 36792 -82256 37760
rect -83194 36787 -82256 36792
rect -84688 36236 -83750 36241
rect -92930 30916 -92040 35580
rect -84688 35268 -84678 36236
rect -83760 35268 -83750 36236
rect -84688 35263 -83750 35268
rect -92938 29912 -92928 30916
rect -92038 29912 -92028 30916
rect -84678 15777 -84014 35263
rect -82904 17571 -82542 36787
rect -80982 33949 -80284 58507
rect -69500 58482 -69490 58682
rect -69290 58482 -69280 58682
rect -69500 58477 -69280 58482
rect -69500 58282 -69280 58287
rect -69500 58082 -69490 58282
rect -69290 58082 -69280 58282
rect -69500 58077 -69280 58082
rect -69500 57882 -69280 57887
rect -69500 57682 -69490 57882
rect -69290 57682 -69280 57882
rect -69500 57677 -69280 57682
rect -69500 57482 -69280 57487
rect -69500 57282 -69490 57482
rect -69290 57282 -69280 57482
rect -69500 57277 -69280 57282
rect -69500 57082 -69280 57087
rect -69500 56882 -69490 57082
rect -69290 56882 -69280 57082
rect -69500 56877 -69280 56882
rect -67772 55404 -66834 55409
rect -67772 54912 -67762 55404
rect -67818 54436 -67762 54912
rect -66844 54912 -66834 55404
rect -66844 54436 -66794 54912
rect -67818 46272 -66794 54436
rect -49962 47756 -49532 62893
rect -2664 50516 -1112 72970
rect -2674 48964 -2664 50516
rect -1112 48964 -1102 50516
rect -2664 48962 -1112 48964
rect -69140 45530 -66794 46272
rect -69140 35168 -66794 35910
rect -81122 33944 -80184 33949
rect -81122 32976 -81112 33944
rect -80194 32976 -80184 33944
rect -81122 32971 -80184 32976
rect -80982 22949 -80284 32971
rect -67818 27004 -66794 35168
rect -53042 32278 -49532 32852
rect -2664 32474 -1112 32476
rect -67818 26528 -67762 27004
rect -67772 26036 -67762 26528
rect -66844 26528 -66794 27004
rect -66844 26036 -66834 26528
rect -67772 26031 -66834 26036
rect -69500 24559 -69280 24564
rect -69500 24359 -69490 24559
rect -69290 24359 -69280 24559
rect -69500 24354 -69280 24359
rect -69500 24159 -69280 24164
rect -69500 23959 -69490 24159
rect -69290 23959 -69280 24159
rect -69500 23954 -69280 23959
rect -69500 23759 -69280 23764
rect -69500 23559 -69490 23759
rect -69290 23559 -69280 23759
rect -69500 23554 -69280 23559
rect -69500 23359 -69280 23364
rect -69500 23159 -69490 23359
rect -69290 23159 -69280 23359
rect -69500 23154 -69280 23159
rect -69500 22959 -69280 22964
rect -81122 22944 -80184 22949
rect -81122 21976 -81112 22944
rect -80194 21976 -80184 22944
rect -69500 22759 -69490 22959
rect -69290 22759 -69280 22959
rect -69500 22754 -69280 22759
rect -81122 21971 -80184 21976
rect -50740 20996 -50072 21001
rect -50740 20916 -50730 20996
rect -50792 20430 -50730 20916
rect -50740 20322 -50730 20430
rect -50082 20322 -50072 20996
rect -50740 20317 -50072 20322
rect -49962 18559 -49532 32278
rect -2674 30922 -2664 32474
rect -1112 30922 -1102 32474
rect -49972 18554 -49304 18559
rect -49972 17880 -49962 18554
rect -49314 17880 -49304 18554
rect -49972 17875 -49304 17880
rect -83226 17566 -82288 17571
rect -83226 16598 -83216 17566
rect -82298 16598 -82288 17566
rect -83226 16593 -82288 16598
rect -84688 15772 -83750 15777
rect -84688 14804 -84678 15772
rect -83760 14804 -83750 15772
rect -84688 14799 -83750 14804
rect -2664 8468 -1112 30922
rect -2674 6916 -2664 8468
rect -1112 6916 -1102 8468
<< via3 >>
rect -2664 72970 -1112 74522
rect -92930 50526 -92040 51530
rect -92928 29912 -92038 30916
rect -69490 58482 -69290 58682
rect -69490 58082 -69290 58282
rect -69490 57682 -69290 57882
rect -69490 57282 -69290 57482
rect -69490 56882 -69290 57082
rect -2664 48964 -1112 50516
rect -69490 24359 -69290 24559
rect -69490 23959 -69290 24159
rect -69490 23559 -69290 23759
rect -69490 23159 -69290 23359
rect -69490 22759 -69290 22959
rect -2664 30922 -1112 32474
rect -2664 6916 -1112 8468
<< metal4 >>
rect -2665 74522 -1111 74523
rect -2665 72970 -2664 74522
rect -1112 72970 -1111 74522
rect -2665 72969 -1111 72970
rect -83908 65794 -66306 66798
rect -53782 65794 -50234 66798
rect 1546 64004 6068 79052
rect -3148 59482 6068 64004
rect -69686 58682 -69272 58724
rect -69686 58482 -69490 58682
rect -69290 58482 -69272 58682
rect -69686 58282 -69272 58482
rect -69686 58082 -69490 58282
rect -69290 58082 -69272 58282
rect -69686 57882 -69272 58082
rect -69686 57682 -69490 57882
rect -69290 57682 -69272 57882
rect -69686 57482 -69272 57682
rect -69686 57282 -69490 57482
rect -69290 57282 -69272 57482
rect -69686 57082 -69272 57282
rect -69686 56882 -69490 57082
rect -69290 56882 -69272 57082
rect -92931 51530 -92039 51531
rect -94876 50526 -92930 51530
rect -92040 50526 -80372 51530
rect -69686 51160 -69272 56882
rect -66306 51528 -65514 56798
rect -53782 55794 -50234 56798
rect -92931 50525 -92039 50526
rect -67946 50524 -65514 51528
rect -2665 50516 -1111 50517
rect -12766 48964 -2664 50516
rect -1112 48964 3234 50516
rect -2665 48963 -1111 48964
rect -67848 44168 -64772 45172
rect -83908 39912 -80278 41530
rect -67848 39912 -66824 44168
rect 2922 38364 34622 43482
rect -66564 34168 -64592 35172
rect -66564 30918 -65514 34168
rect -2665 32474 -1111 32475
rect -12770 30922 -2664 32474
rect -1112 30922 3230 32474
rect -2665 30921 -1111 30922
rect -67848 30917 -65514 30918
rect -92929 30916 -92037 30917
rect -94876 29912 -92928 30916
rect -92038 29912 -79394 30916
rect -67950 30915 -65514 30917
rect -69140 29914 -65514 30915
rect -69140 29912 -66650 29914
rect -92929 29911 -92037 29912
rect -69686 24559 -69272 29912
rect -69140 29911 -67848 29912
rect -66306 25648 -65514 29914
rect -66306 24644 -65146 25648
rect -53782 24642 -50168 25646
rect -69686 24359 -69490 24559
rect -69290 24359 -69272 24559
rect -69686 24159 -69272 24359
rect -69686 23959 -69490 24159
rect -69290 23959 -69272 24159
rect -69686 23759 -69272 23959
rect -69686 23559 -69490 23759
rect -69290 23559 -69272 23759
rect -69686 23359 -69272 23559
rect -69686 23159 -69490 23359
rect -69290 23159 -69272 23359
rect -69686 22959 -69272 23159
rect -69686 22759 -69490 22959
rect -69290 22759 -69272 22959
rect -69686 22717 -69272 22759
rect -3148 17434 6068 21956
rect -86606 17192 -83908 17246
rect -83908 14642 -66188 15646
rect -53782 14642 -50168 15646
rect -2665 8468 -1111 8469
rect -2665 6916 -2664 8468
rect -1112 6916 -1111 8468
rect -2665 6915 -1111 6916
rect 1546 2386 6068 17434
<< via4 >>
rect -86606 64194 -83908 66798
rect -97574 48980 -94876 51530
rect -86606 39462 -83908 42012
rect -97574 29912 -94876 32462
rect -86606 14642 -83908 17192
<< metal5 >>
rect -86630 66798 -83884 66822
rect -86630 64194 -86606 66798
rect -83908 64194 -83884 66798
rect -86630 64170 -83884 64194
rect -97598 51530 -94852 51554
rect -97598 48980 -97574 51530
rect -94876 48980 -94852 51530
rect -97598 48956 -94852 48980
rect -97574 32486 -94876 48956
rect -86606 42036 -83908 64170
rect -86630 42012 -83884 42036
rect -86630 39462 -86606 42012
rect -83908 39462 -83884 42012
rect -86630 39438 -83884 39462
rect -97598 32462 -94852 32486
rect -97598 29912 -97574 32462
rect -94876 29912 -94852 32462
rect -97598 29888 -94852 29912
rect -86606 17270 -83908 39438
rect -86630 17192 -83884 17270
rect -86630 14642 -86606 17192
rect -83908 14642 -83884 17192
rect -86630 14618 -83884 14642
use biasing_network  biasing_network_0
timestamp 1629274976
transform 0 1 -88634 -1 0 41178
box -4801 -4684 5802 1016
use S_to_D_final  S_to_D_final_0 ~/magic/class_d_audio_amplifier/S_to_D
timestamp 1629190088
transform 1 0 -119284 0 1 30788
box 38304 -876 51436 20741
use integrator  integrator_0 ~/magic/class_d_audio_amplifier/integrator
timestamp 1629189639
transform 1 0 -103940 0 1 56496
box 35518 -702 55900 26032
use integrator  integrator_1
timestamp 1629189639
transform 1 0 -103940 0 -1 24944
box 35518 -702 55900 26032
use triangle_revised  triangle_revised_0 ~/magic/class_d_audio_amplifier/triang
timestamp 1629189331
transform 1 0 -64913 0 1 34158
box -1869 -1600 26228 14688
use comparator_revised  comparator_revised_0 ~/magic/class_d_audio_amplifier/comparator
timestamp 1628692234
transform 1 0 -69200 0 1 54904
box 18966 890 31490 11894
use comparator_revised  comparator_revised_1
timestamp 1628692234
transform 1 0 -69200 0 -1 26535
box 18966 890 31490 11894
use dead_time_final  dead_time_final_1 ~/magic/class_d_audio_amplifier/dead_time
timestamp 1629091460
transform 1 0 -94234 0 -1 37760
box 57308 806 91570 35374
use dead_time_final  dead_time_final_0
timestamp 1629091460
transform 1 0 -94234 0 1 43678
box 57308 806 91570 35374
use output_driver_final  output_driver_final_0 ~/magic/class_d_audio_amplifier/output_driver
timestamp 1629091687
transform 1 0 -114276 0 1 -1168
box 116370 3554 149002 80219
<< labels >>
flabel metal5 -86368 36130 -86368 36130 0 FreeSans 16000 0 0 0 avdd
flabel metal4 22812 41026 22812 41026 0 FreeSans 16000 0 0 0 dvss
flabel space 27436 74066 27436 74066 0 FreeSans 16000 0 0 0 dvdd1
flabel space 21046 4722 21046 4722 0 FreeSans 16000 0 0 0 dvdd2
flabel metal3 -80704 46694 -80704 46694 0 FreeSans 16000 0 0 0 vin
flabel metal3 -49706 50138 -49706 50138 0 FreeSans 16000 0 0 0 vtriang
flabel metal3 -67224 48050 -67224 48050 0 FreeSans 16000 0 0 0 vin_p
flabel metal3 -67224 32814 -67224 32814 0 FreeSans 16000 0 0 0 vin_n
flabel metal2 -49170 60680 -49170 60680 0 FreeSans 16000 0 0 0 error_p
flabel metal2 -49214 20614 -49214 20614 0 FreeSans 16000 0 0 0 error_n
flabel metal1 -37988 61218 -37988 61218 0 FreeSans 16000 0 0 0 vcmp_p
flabel metal1 -38868 19748 -38868 19748 0 FreeSans 16000 0 0 0 vcmp_n
flabel metal2 128 69622 128 69622 0 FreeSans 16000 0 0 0 vp_p
flabel metal2 778 56776 778 56776 0 FreeSans 16000 0 0 0 vp_n
flabel metal2 1050 24596 1050 24596 0 FreeSans 16000 0 0 0 vn_n
flabel metal2 30 11592 30 11592 0 FreeSans 16000 0 0 0 vn_p
flabel space 23806 24106 23806 24106 0 FreeSans 16000 0 0 0 out_n
flabel space 29186 57864 29186 57864 0 FreeSans 16000 0 0 0 out_p
flabel metal1 -64534 43406 -64534 43406 0 FreeSans 16000 0 0 0 vbias1
flabel metal1 -51006 43350 -51006 43350 0 FreeSans 16000 0 0 0 vbias2
flabel metal1 -79980 42928 -79980 42928 0 FreeSans 16000 0 0 0 vbias3
flabel metal1 -79982 39148 -79982 39148 0 FreeSans 16000 0 0 0 vbias4
flabel metal1 -65916 64974 -65916 64974 0 FreeSans 16000 0 0 0 vbias5
flabel metal1 -65920 16400 -65920 16400 0 FreeSans 16000 0 0 0 vbias6
flabel metal1 -49840 64998 -49840 64998 0 FreeSans 16000 0 0 0 vbias7
flabel metal1 -49852 16424 -49852 16424 0 FreeSans 16000 0 0 0 vbias8
flabel space -93064 40710 -93064 40710 0 FreeSans 16000 0 0 0 iin
flabel metal5 -96730 35142 -96730 35142 0 FreeSans 16000 0 0 0 avss
flabel metal3 -80608 26478 -80608 26478 0 FreeSans 16000 0 0 0 vref
<< end >>
