magic
tech sky130A
magscale 1 2
timestamp 1630397679
<< nwell >>
rect 9878 5638 18876 8168
rect 5006 4212 18876 5638
rect 2404 2786 18876 4212
rect -832 110 -376 622
rect 2404 -2686 9446 -1260
rect 5006 -4112 9446 -2686
<< pwell >>
rect 9908 10402 19232 13484
rect 5234 5752 9434 7280
rect 2450 4306 4424 5480
rect 2450 -3954 4424 -2780
rect 5234 -7154 9434 -5626
<< nmos >>
rect 10394 12048 10424 13048
rect 10604 12048 10634 13048
rect 10814 12048 10844 13048
rect 11024 12048 11054 13048
rect 11234 12048 11264 13048
rect 11444 12048 11474 13048
rect 11654 12048 11684 13048
rect 11864 12048 11894 13048
rect 12074 12048 12104 13048
rect 12284 12048 12314 13048
rect 12494 12048 12524 13048
rect 12704 12048 12734 13048
rect 12914 12048 12944 13048
rect 13124 12048 13154 13048
rect 13334 12048 13364 13048
rect 13544 12048 13574 13048
rect 13754 12048 13784 13048
rect 13964 12048 13994 13048
rect 14174 12048 14204 13048
rect 14384 12048 14414 13048
rect 14594 12048 14624 13048
rect 14804 12048 14834 13048
rect 15014 12048 15044 13048
rect 15224 12048 15254 13048
rect 15434 12048 15464 13048
rect 15644 12048 15674 13048
rect 15854 12048 15884 13048
rect 16064 12048 16094 13048
rect 16274 12048 16304 13048
rect 16484 12048 16514 13048
rect 16694 12048 16724 13048
rect 16904 12048 16934 13048
rect 17114 12048 17144 13048
rect 17324 12048 17354 13048
rect 17534 12048 17564 13048
rect 17744 12048 17774 13048
rect 17954 12048 17984 13048
rect 18164 12048 18194 13048
rect 18374 12048 18404 13048
rect 18584 12048 18614 13048
rect 10394 10830 10424 11830
rect 10604 10830 10634 11830
rect 10814 10830 10844 11830
rect 11024 10830 11054 11830
rect 11234 10830 11264 11830
rect 11444 10830 11474 11830
rect 11654 10830 11684 11830
rect 11864 10830 11894 11830
rect 12074 10830 12104 11830
rect 12284 10830 12314 11830
rect 12494 10830 12524 11830
rect 12704 10830 12734 11830
rect 12914 10830 12944 11830
rect 13124 10830 13154 11830
rect 13334 10830 13364 11830
rect 13544 10830 13574 11830
rect 13754 10830 13784 11830
rect 13964 10830 13994 11830
rect 14174 10830 14204 11830
rect 14384 10830 14414 11830
rect 14594 10830 14624 11830
rect 14804 10830 14834 11830
rect 15014 10830 15044 11830
rect 15224 10830 15254 11830
rect 15434 10830 15464 11830
rect 15644 10830 15674 11830
rect 15854 10830 15884 11830
rect 16064 10830 16094 11830
rect 16274 10830 16304 11830
rect 16484 10830 16514 11830
rect 16694 10830 16724 11830
rect 16904 10830 16934 11830
rect 17114 10830 17144 11830
rect 17324 10830 17354 11830
rect 17534 10830 17564 11830
rect 17744 10830 17774 11830
rect 17954 10830 17984 11830
rect 18164 10830 18194 11830
rect 18374 10830 18404 11830
rect 18584 10830 18614 11830
rect 5544 5964 5574 6964
rect 5754 5964 5784 6964
rect 5964 5964 5994 6964
rect 6174 5964 6204 6964
rect 6384 5964 6414 6964
rect 6594 5964 6624 6964
rect 6804 5964 6834 6964
rect 7014 5964 7044 6964
rect 7224 5964 7254 6964
rect 7434 5964 7464 6964
rect 7644 5964 7674 6964
rect 7854 5964 7884 6964
rect 8064 5964 8094 6964
rect 8274 5964 8304 6964
rect 8484 5964 8514 6964
rect 8694 5964 8724 6964
rect 8904 5964 8934 6964
rect 9114 5964 9144 6964
rect 2632 4340 2662 5340
rect 3580 4340 3610 5340
rect 3790 4340 3820 5340
rect 4000 4340 4030 5340
rect 4210 4340 4240 5340
rect 2632 -3814 2662 -2814
rect 3580 -3814 3610 -2814
rect 3790 -3814 3820 -2814
rect 4000 -3814 4030 -2814
rect 4210 -3814 4240 -2814
rect 5544 -6838 5574 -5838
rect 5754 -6838 5784 -5838
rect 5964 -6838 5994 -5838
rect 6174 -6838 6204 -5838
rect 6384 -6838 6414 -5838
rect 6594 -6838 6624 -5838
rect 6804 -6838 6834 -5838
rect 7014 -6838 7044 -5838
rect 7224 -6838 7254 -5838
rect 7434 -6838 7464 -5838
rect 7644 -6838 7674 -5838
rect 7854 -6838 7884 -5838
rect 8064 -6838 8094 -5838
rect 8274 -6838 8304 -5838
rect 8484 -6838 8514 -5838
rect 8694 -6838 8724 -5838
rect 8904 -6838 8934 -5838
rect 9114 -6838 9144 -5838
<< pmos >>
rect 2632 3112 2662 4112
rect 2728 3112 2758 4112
rect 3370 3112 3400 4112
rect 3580 3112 3610 4112
rect 3790 3112 3820 4112
rect 4000 3112 4030 4112
rect 4210 3112 4240 4112
rect 4420 3112 4450 4112
rect 4630 3112 4660 4112
rect 4840 3112 4870 4112
rect 5544 4348 5574 5348
rect 5754 4348 5784 5348
rect 5964 4348 5994 5348
rect 6174 4348 6204 5348
rect 6384 4348 6414 5348
rect 6594 4348 6624 5348
rect 6804 4348 6834 5348
rect 7014 4348 7044 5348
rect 7224 4348 7254 5348
rect 7434 4348 7464 5348
rect 7644 4348 7674 5348
rect 7854 4348 7884 5348
rect 8064 4348 8094 5348
rect 8274 4348 8304 5348
rect 8484 4348 8514 5348
rect 8694 4348 8724 5348
rect 8904 4348 8934 5348
rect 9114 4348 9144 5348
rect 5544 3112 5574 4112
rect 5754 3112 5784 4112
rect 5964 3112 5994 4112
rect 6174 3112 6204 4112
rect 6384 3112 6414 4112
rect 6594 3112 6624 4112
rect 6804 3112 6834 4112
rect 7014 3112 7044 4112
rect 7224 3112 7254 4112
rect 7434 3112 7464 4112
rect 7644 3112 7674 4112
rect 7854 3112 7884 4112
rect 8064 3112 8094 4112
rect 8274 3112 8304 4112
rect 8484 3112 8514 4112
rect 8694 3112 8724 4112
rect 8904 3112 8934 4112
rect 9114 3112 9144 4112
rect 10394 6820 10424 7820
rect 10604 6820 10634 7820
rect 10814 6820 10844 7820
rect 11024 6820 11054 7820
rect 11234 6820 11264 7820
rect 11444 6820 11474 7820
rect 11654 6820 11684 7820
rect 11864 6820 11894 7820
rect 12074 6820 12104 7820
rect 12284 6820 12314 7820
rect 12494 6820 12524 7820
rect 12704 6820 12734 7820
rect 12914 6820 12944 7820
rect 13124 6820 13154 7820
rect 13334 6820 13364 7820
rect 13544 6820 13574 7820
rect 13754 6820 13784 7820
rect 13964 6820 13994 7820
rect 14174 6820 14204 7820
rect 14384 6820 14414 7820
rect 14594 6820 14624 7820
rect 14804 6820 14834 7820
rect 15014 6820 15044 7820
rect 15224 6820 15254 7820
rect 15434 6820 15464 7820
rect 15644 6820 15674 7820
rect 15854 6820 15884 7820
rect 16064 6820 16094 7820
rect 16274 6820 16304 7820
rect 16484 6820 16514 7820
rect 16694 6820 16724 7820
rect 16904 6820 16934 7820
rect 17114 6820 17144 7820
rect 17324 6820 17354 7820
rect 17534 6820 17564 7820
rect 17744 6820 17774 7820
rect 17954 6820 17984 7820
rect 18164 6820 18194 7820
rect 18374 6820 18404 7820
rect 18584 6820 18614 7820
rect 10394 5584 10424 6584
rect 10604 5584 10634 6584
rect 10814 5584 10844 6584
rect 11024 5584 11054 6584
rect 11234 5584 11264 6584
rect 11444 5584 11474 6584
rect 11654 5584 11684 6584
rect 11864 5584 11894 6584
rect 12074 5584 12104 6584
rect 12284 5584 12314 6584
rect 12494 5584 12524 6584
rect 12704 5584 12734 6584
rect 12914 5584 12944 6584
rect 13124 5584 13154 6584
rect 13334 5584 13364 6584
rect 13544 5584 13574 6584
rect 13754 5584 13784 6584
rect 13964 5584 13994 6584
rect 14174 5584 14204 6584
rect 14384 5584 14414 6584
rect 14594 5584 14624 6584
rect 14804 5584 14834 6584
rect 15014 5584 15044 6584
rect 15224 5584 15254 6584
rect 15434 5584 15464 6584
rect 15644 5584 15674 6584
rect 15854 5584 15884 6584
rect 16064 5584 16094 6584
rect 16274 5584 16304 6584
rect 16484 5584 16514 6584
rect 16694 5584 16724 6584
rect 16904 5584 16934 6584
rect 17114 5584 17144 6584
rect 17324 5584 17354 6584
rect 17534 5584 17564 6584
rect 17744 5584 17774 6584
rect 17954 5584 17984 6584
rect 18164 5584 18194 6584
rect 18374 5584 18404 6584
rect 18584 5584 18614 6584
rect 10394 4348 10424 5348
rect 10604 4348 10634 5348
rect 10814 4348 10844 5348
rect 11024 4348 11054 5348
rect 11234 4348 11264 5348
rect 11444 4348 11474 5348
rect 11654 4348 11684 5348
rect 11864 4348 11894 5348
rect 12074 4348 12104 5348
rect 12284 4348 12314 5348
rect 12494 4348 12524 5348
rect 12704 4348 12734 5348
rect 12914 4348 12944 5348
rect 13124 4348 13154 5348
rect 13334 4348 13364 5348
rect 13544 4348 13574 5348
rect 13754 4348 13784 5348
rect 13964 4348 13994 5348
rect 14174 4348 14204 5348
rect 14384 4348 14414 5348
rect 14594 4348 14624 5348
rect 14804 4348 14834 5348
rect 15014 4348 15044 5348
rect 15224 4348 15254 5348
rect 15434 4348 15464 5348
rect 15644 4348 15674 5348
rect 15854 4348 15884 5348
rect 16064 4348 16094 5348
rect 16274 4348 16304 5348
rect 16484 4348 16514 5348
rect 16694 4348 16724 5348
rect 16904 4348 16934 5348
rect 17114 4348 17144 5348
rect 17324 4348 17354 5348
rect 17534 4348 17564 5348
rect 17744 4348 17774 5348
rect 17954 4348 17984 5348
rect 18164 4348 18194 5348
rect 18374 4348 18404 5348
rect 18584 4348 18614 5348
rect 10394 3112 10424 4112
rect 10604 3112 10634 4112
rect 10814 3112 10844 4112
rect 11024 3112 11054 4112
rect 11234 3112 11264 4112
rect 11444 3112 11474 4112
rect 11654 3112 11684 4112
rect 11864 3112 11894 4112
rect 12074 3112 12104 4112
rect 12284 3112 12314 4112
rect 12494 3112 12524 4112
rect 12704 3112 12734 4112
rect 12914 3112 12944 4112
rect 13124 3112 13154 4112
rect 13334 3112 13364 4112
rect 13544 3112 13574 4112
rect 13754 3112 13784 4112
rect 13964 3112 13994 4112
rect 14174 3112 14204 4112
rect 14384 3112 14414 4112
rect 14594 3112 14624 4112
rect 14804 3112 14834 4112
rect 15014 3112 15044 4112
rect 15224 3112 15254 4112
rect 15434 3112 15464 4112
rect 15644 3112 15674 4112
rect 15854 3112 15884 4112
rect 16064 3112 16094 4112
rect 16274 3112 16304 4112
rect 16484 3112 16514 4112
rect 16694 3112 16724 4112
rect 16904 3112 16934 4112
rect 17114 3112 17144 4112
rect 17324 3112 17354 4112
rect 17534 3112 17564 4112
rect 17744 3112 17774 4112
rect 17954 3112 17984 4112
rect 18164 3112 18194 4112
rect 18374 3112 18404 4112
rect 18584 3112 18614 4112
rect 2632 -2586 2662 -1586
rect 2728 -2586 2758 -1586
rect 3370 -2586 3400 -1586
rect 3580 -2586 3610 -1586
rect 3790 -2586 3820 -1586
rect 4000 -2586 4030 -1586
rect 4210 -2586 4240 -1586
rect 4420 -2586 4450 -1586
rect 4630 -2586 4660 -1586
rect 4840 -2586 4870 -1586
rect 5544 -2586 5574 -1586
rect 5754 -2586 5784 -1586
rect 5964 -2586 5994 -1586
rect 6174 -2586 6204 -1586
rect 6384 -2586 6414 -1586
rect 6594 -2586 6624 -1586
rect 6804 -2586 6834 -1586
rect 7014 -2586 7044 -1586
rect 7224 -2586 7254 -1586
rect 7434 -2586 7464 -1586
rect 7644 -2586 7674 -1586
rect 7854 -2586 7884 -1586
rect 8064 -2586 8094 -1586
rect 8274 -2586 8304 -1586
rect 8484 -2586 8514 -1586
rect 8694 -2586 8724 -1586
rect 8904 -2586 8934 -1586
rect 9114 -2586 9144 -1586
rect 5544 -3822 5574 -2822
rect 5754 -3822 5784 -2822
rect 5964 -3822 5994 -2822
rect 6174 -3822 6204 -2822
rect 6384 -3822 6414 -2822
rect 6594 -3822 6624 -2822
rect 6804 -3822 6834 -2822
rect 7014 -3822 7044 -2822
rect 7224 -3822 7254 -2822
rect 7434 -3822 7464 -2822
rect 7644 -3822 7674 -2822
rect 7854 -3822 7884 -2822
rect 8064 -3822 8094 -2822
rect 8274 -3822 8304 -2822
rect 8484 -3822 8514 -2822
rect 8694 -3822 8724 -2822
rect 8904 -3822 8934 -2822
rect 9114 -3822 9144 -2822
<< ndiff >>
rect 10332 13036 10394 13048
rect 10332 12060 10344 13036
rect 10378 12060 10394 13036
rect 10332 12048 10394 12060
rect 10424 13036 10486 13048
rect 10424 12060 10440 13036
rect 10474 12060 10486 13036
rect 10424 12048 10486 12060
rect 10542 13036 10604 13048
rect 10542 12060 10554 13036
rect 10588 12060 10604 13036
rect 10542 12048 10604 12060
rect 10634 13036 10696 13048
rect 10634 12060 10650 13036
rect 10684 12060 10696 13036
rect 10634 12048 10696 12060
rect 10752 13036 10814 13048
rect 10752 12060 10764 13036
rect 10798 12060 10814 13036
rect 10752 12048 10814 12060
rect 10844 13036 10906 13048
rect 10844 12060 10860 13036
rect 10894 12060 10906 13036
rect 10844 12048 10906 12060
rect 10962 13036 11024 13048
rect 10962 12060 10974 13036
rect 11008 12060 11024 13036
rect 10962 12048 11024 12060
rect 11054 13036 11116 13048
rect 11054 12060 11070 13036
rect 11104 12060 11116 13036
rect 11054 12048 11116 12060
rect 11172 13036 11234 13048
rect 11172 12060 11184 13036
rect 11218 12060 11234 13036
rect 11172 12048 11234 12060
rect 11264 13036 11326 13048
rect 11264 12060 11280 13036
rect 11314 12060 11326 13036
rect 11264 12048 11326 12060
rect 11382 13036 11444 13048
rect 11382 12060 11394 13036
rect 11428 12060 11444 13036
rect 11382 12048 11444 12060
rect 11474 13036 11536 13048
rect 11474 12060 11490 13036
rect 11524 12060 11536 13036
rect 11474 12048 11536 12060
rect 11592 13036 11654 13048
rect 11592 12060 11604 13036
rect 11638 12060 11654 13036
rect 11592 12048 11654 12060
rect 11684 13036 11746 13048
rect 11684 12060 11700 13036
rect 11734 12060 11746 13036
rect 11684 12048 11746 12060
rect 11802 13036 11864 13048
rect 11802 12060 11814 13036
rect 11848 12060 11864 13036
rect 11802 12048 11864 12060
rect 11894 13036 11956 13048
rect 11894 12060 11910 13036
rect 11944 12060 11956 13036
rect 11894 12048 11956 12060
rect 12012 13036 12074 13048
rect 12012 12060 12024 13036
rect 12058 12060 12074 13036
rect 12012 12048 12074 12060
rect 12104 13036 12166 13048
rect 12104 12060 12120 13036
rect 12154 12060 12166 13036
rect 12104 12048 12166 12060
rect 12222 13036 12284 13048
rect 12222 12060 12234 13036
rect 12268 12060 12284 13036
rect 12222 12048 12284 12060
rect 12314 13036 12376 13048
rect 12314 12060 12330 13036
rect 12364 12060 12376 13036
rect 12314 12048 12376 12060
rect 12432 13036 12494 13048
rect 12432 12060 12444 13036
rect 12478 12060 12494 13036
rect 12432 12048 12494 12060
rect 12524 13036 12586 13048
rect 12524 12060 12540 13036
rect 12574 12060 12586 13036
rect 12524 12048 12586 12060
rect 12642 13036 12704 13048
rect 12642 12060 12654 13036
rect 12688 12060 12704 13036
rect 12642 12048 12704 12060
rect 12734 13036 12796 13048
rect 12734 12060 12750 13036
rect 12784 12060 12796 13036
rect 12734 12048 12796 12060
rect 12852 13036 12914 13048
rect 12852 12060 12864 13036
rect 12898 12060 12914 13036
rect 12852 12048 12914 12060
rect 12944 13036 13006 13048
rect 12944 12060 12960 13036
rect 12994 12060 13006 13036
rect 12944 12048 13006 12060
rect 13062 13036 13124 13048
rect 13062 12060 13074 13036
rect 13108 12060 13124 13036
rect 13062 12048 13124 12060
rect 13154 13036 13216 13048
rect 13154 12060 13170 13036
rect 13204 12060 13216 13036
rect 13154 12048 13216 12060
rect 13272 13036 13334 13048
rect 13272 12060 13284 13036
rect 13318 12060 13334 13036
rect 13272 12048 13334 12060
rect 13364 13036 13426 13048
rect 13364 12060 13380 13036
rect 13414 12060 13426 13036
rect 13364 12048 13426 12060
rect 13482 13036 13544 13048
rect 13482 12060 13494 13036
rect 13528 12060 13544 13036
rect 13482 12048 13544 12060
rect 13574 13036 13636 13048
rect 13574 12060 13590 13036
rect 13624 12060 13636 13036
rect 13574 12048 13636 12060
rect 13692 13036 13754 13048
rect 13692 12060 13704 13036
rect 13738 12060 13754 13036
rect 13692 12048 13754 12060
rect 13784 13036 13846 13048
rect 13784 12060 13800 13036
rect 13834 12060 13846 13036
rect 13784 12048 13846 12060
rect 13902 13036 13964 13048
rect 13902 12060 13914 13036
rect 13948 12060 13964 13036
rect 13902 12048 13964 12060
rect 13994 13036 14056 13048
rect 13994 12060 14010 13036
rect 14044 12060 14056 13036
rect 13994 12048 14056 12060
rect 14112 13036 14174 13048
rect 14112 12060 14124 13036
rect 14158 12060 14174 13036
rect 14112 12048 14174 12060
rect 14204 13036 14266 13048
rect 14204 12060 14220 13036
rect 14254 12060 14266 13036
rect 14204 12048 14266 12060
rect 14322 13036 14384 13048
rect 14322 12060 14334 13036
rect 14368 12060 14384 13036
rect 14322 12048 14384 12060
rect 14414 13036 14476 13048
rect 14414 12060 14430 13036
rect 14464 12060 14476 13036
rect 14414 12048 14476 12060
rect 14532 13036 14594 13048
rect 14532 12060 14544 13036
rect 14578 12060 14594 13036
rect 14532 12048 14594 12060
rect 14624 13036 14686 13048
rect 14624 12060 14640 13036
rect 14674 12060 14686 13036
rect 14624 12048 14686 12060
rect 14742 13036 14804 13048
rect 14742 12060 14754 13036
rect 14788 12060 14804 13036
rect 14742 12048 14804 12060
rect 14834 13036 14896 13048
rect 14834 12060 14850 13036
rect 14884 12060 14896 13036
rect 14834 12048 14896 12060
rect 14952 13036 15014 13048
rect 14952 12060 14964 13036
rect 14998 12060 15014 13036
rect 14952 12048 15014 12060
rect 15044 13036 15106 13048
rect 15044 12060 15060 13036
rect 15094 12060 15106 13036
rect 15044 12048 15106 12060
rect 15162 13036 15224 13048
rect 15162 12060 15174 13036
rect 15208 12060 15224 13036
rect 15162 12048 15224 12060
rect 15254 13036 15316 13048
rect 15254 12060 15270 13036
rect 15304 12060 15316 13036
rect 15254 12048 15316 12060
rect 15372 13036 15434 13048
rect 15372 12060 15384 13036
rect 15418 12060 15434 13036
rect 15372 12048 15434 12060
rect 15464 13036 15526 13048
rect 15464 12060 15480 13036
rect 15514 12060 15526 13036
rect 15464 12048 15526 12060
rect 15582 13036 15644 13048
rect 15582 12060 15594 13036
rect 15628 12060 15644 13036
rect 15582 12048 15644 12060
rect 15674 13036 15736 13048
rect 15674 12060 15690 13036
rect 15724 12060 15736 13036
rect 15674 12048 15736 12060
rect 15792 13036 15854 13048
rect 15792 12060 15804 13036
rect 15838 12060 15854 13036
rect 15792 12048 15854 12060
rect 15884 13036 15946 13048
rect 15884 12060 15900 13036
rect 15934 12060 15946 13036
rect 15884 12048 15946 12060
rect 16002 13036 16064 13048
rect 16002 12060 16014 13036
rect 16048 12060 16064 13036
rect 16002 12048 16064 12060
rect 16094 13036 16156 13048
rect 16094 12060 16110 13036
rect 16144 12060 16156 13036
rect 16094 12048 16156 12060
rect 16212 13036 16274 13048
rect 16212 12060 16224 13036
rect 16258 12060 16274 13036
rect 16212 12048 16274 12060
rect 16304 13036 16366 13048
rect 16304 12060 16320 13036
rect 16354 12060 16366 13036
rect 16304 12048 16366 12060
rect 16422 13036 16484 13048
rect 16422 12060 16434 13036
rect 16468 12060 16484 13036
rect 16422 12048 16484 12060
rect 16514 13036 16576 13048
rect 16514 12060 16530 13036
rect 16564 12060 16576 13036
rect 16514 12048 16576 12060
rect 16632 13036 16694 13048
rect 16632 12060 16644 13036
rect 16678 12060 16694 13036
rect 16632 12048 16694 12060
rect 16724 13036 16786 13048
rect 16724 12060 16740 13036
rect 16774 12060 16786 13036
rect 16724 12048 16786 12060
rect 16842 13036 16904 13048
rect 16842 12060 16854 13036
rect 16888 12060 16904 13036
rect 16842 12048 16904 12060
rect 16934 13036 16996 13048
rect 16934 12060 16950 13036
rect 16984 12060 16996 13036
rect 16934 12048 16996 12060
rect 17052 13036 17114 13048
rect 17052 12060 17064 13036
rect 17098 12060 17114 13036
rect 17052 12048 17114 12060
rect 17144 13036 17206 13048
rect 17144 12060 17160 13036
rect 17194 12060 17206 13036
rect 17144 12048 17206 12060
rect 17262 13036 17324 13048
rect 17262 12060 17274 13036
rect 17308 12060 17324 13036
rect 17262 12048 17324 12060
rect 17354 13036 17416 13048
rect 17354 12060 17370 13036
rect 17404 12060 17416 13036
rect 17354 12048 17416 12060
rect 17472 13036 17534 13048
rect 17472 12060 17484 13036
rect 17518 12060 17534 13036
rect 17472 12048 17534 12060
rect 17564 13036 17626 13048
rect 17564 12060 17580 13036
rect 17614 12060 17626 13036
rect 17564 12048 17626 12060
rect 17682 13036 17744 13048
rect 17682 12060 17694 13036
rect 17728 12060 17744 13036
rect 17682 12048 17744 12060
rect 17774 13036 17836 13048
rect 17774 12060 17790 13036
rect 17824 12060 17836 13036
rect 17774 12048 17836 12060
rect 17892 13036 17954 13048
rect 17892 12060 17904 13036
rect 17938 12060 17954 13036
rect 17892 12048 17954 12060
rect 17984 13036 18046 13048
rect 17984 12060 18000 13036
rect 18034 12060 18046 13036
rect 17984 12048 18046 12060
rect 18102 13036 18164 13048
rect 18102 12060 18114 13036
rect 18148 12060 18164 13036
rect 18102 12048 18164 12060
rect 18194 13036 18256 13048
rect 18194 12060 18210 13036
rect 18244 12060 18256 13036
rect 18194 12048 18256 12060
rect 18312 13036 18374 13048
rect 18312 12060 18324 13036
rect 18358 12060 18374 13036
rect 18312 12048 18374 12060
rect 18404 13036 18466 13048
rect 18404 12060 18420 13036
rect 18454 12060 18466 13036
rect 18404 12048 18466 12060
rect 18522 13036 18584 13048
rect 18522 12060 18534 13036
rect 18568 12060 18584 13036
rect 18522 12048 18584 12060
rect 18614 13036 18676 13048
rect 18614 12060 18630 13036
rect 18664 12060 18676 13036
rect 18614 12048 18676 12060
rect 10332 11818 10394 11830
rect 10332 10842 10344 11818
rect 10378 10842 10394 11818
rect 10332 10830 10394 10842
rect 10424 11818 10486 11830
rect 10424 10842 10440 11818
rect 10474 10842 10486 11818
rect 10424 10830 10486 10842
rect 10542 11818 10604 11830
rect 10542 10842 10554 11818
rect 10588 10842 10604 11818
rect 10542 10830 10604 10842
rect 10634 11818 10696 11830
rect 10634 10842 10650 11818
rect 10684 10842 10696 11818
rect 10634 10830 10696 10842
rect 10752 11818 10814 11830
rect 10752 10842 10764 11818
rect 10798 10842 10814 11818
rect 10752 10830 10814 10842
rect 10844 11818 10906 11830
rect 10844 10842 10860 11818
rect 10894 10842 10906 11818
rect 10844 10830 10906 10842
rect 10962 11818 11024 11830
rect 10962 10842 10974 11818
rect 11008 10842 11024 11818
rect 10962 10830 11024 10842
rect 11054 11818 11116 11830
rect 11054 10842 11070 11818
rect 11104 10842 11116 11818
rect 11054 10830 11116 10842
rect 11172 11818 11234 11830
rect 11172 10842 11184 11818
rect 11218 10842 11234 11818
rect 11172 10830 11234 10842
rect 11264 11818 11326 11830
rect 11264 10842 11280 11818
rect 11314 10842 11326 11818
rect 11264 10830 11326 10842
rect 11382 11818 11444 11830
rect 11382 10842 11394 11818
rect 11428 10842 11444 11818
rect 11382 10830 11444 10842
rect 11474 11818 11536 11830
rect 11474 10842 11490 11818
rect 11524 10842 11536 11818
rect 11474 10830 11536 10842
rect 11592 11818 11654 11830
rect 11592 10842 11604 11818
rect 11638 10842 11654 11818
rect 11592 10830 11654 10842
rect 11684 11818 11746 11830
rect 11684 10842 11700 11818
rect 11734 10842 11746 11818
rect 11684 10830 11746 10842
rect 11802 11818 11864 11830
rect 11802 10842 11814 11818
rect 11848 10842 11864 11818
rect 11802 10830 11864 10842
rect 11894 11818 11956 11830
rect 11894 10842 11910 11818
rect 11944 10842 11956 11818
rect 11894 10830 11956 10842
rect 12012 11818 12074 11830
rect 12012 10842 12024 11818
rect 12058 10842 12074 11818
rect 12012 10830 12074 10842
rect 12104 11818 12166 11830
rect 12104 10842 12120 11818
rect 12154 10842 12166 11818
rect 12104 10830 12166 10842
rect 12222 11818 12284 11830
rect 12222 10842 12234 11818
rect 12268 10842 12284 11818
rect 12222 10830 12284 10842
rect 12314 11818 12376 11830
rect 12314 10842 12330 11818
rect 12364 10842 12376 11818
rect 12314 10830 12376 10842
rect 12432 11818 12494 11830
rect 12432 10842 12444 11818
rect 12478 10842 12494 11818
rect 12432 10830 12494 10842
rect 12524 11818 12586 11830
rect 12524 10842 12540 11818
rect 12574 10842 12586 11818
rect 12524 10830 12586 10842
rect 12642 11818 12704 11830
rect 12642 10842 12654 11818
rect 12688 10842 12704 11818
rect 12642 10830 12704 10842
rect 12734 11818 12796 11830
rect 12734 10842 12750 11818
rect 12784 10842 12796 11818
rect 12734 10830 12796 10842
rect 12852 11818 12914 11830
rect 12852 10842 12864 11818
rect 12898 10842 12914 11818
rect 12852 10830 12914 10842
rect 12944 11818 13006 11830
rect 12944 10842 12960 11818
rect 12994 10842 13006 11818
rect 12944 10830 13006 10842
rect 13062 11818 13124 11830
rect 13062 10842 13074 11818
rect 13108 10842 13124 11818
rect 13062 10830 13124 10842
rect 13154 11818 13216 11830
rect 13154 10842 13170 11818
rect 13204 10842 13216 11818
rect 13154 10830 13216 10842
rect 13272 11818 13334 11830
rect 13272 10842 13284 11818
rect 13318 10842 13334 11818
rect 13272 10830 13334 10842
rect 13364 11818 13426 11830
rect 13364 10842 13380 11818
rect 13414 10842 13426 11818
rect 13364 10830 13426 10842
rect 13482 11818 13544 11830
rect 13482 10842 13494 11818
rect 13528 10842 13544 11818
rect 13482 10830 13544 10842
rect 13574 11818 13636 11830
rect 13574 10842 13590 11818
rect 13624 10842 13636 11818
rect 13574 10830 13636 10842
rect 13692 11818 13754 11830
rect 13692 10842 13704 11818
rect 13738 10842 13754 11818
rect 13692 10830 13754 10842
rect 13784 11818 13846 11830
rect 13784 10842 13800 11818
rect 13834 10842 13846 11818
rect 13784 10830 13846 10842
rect 13902 11818 13964 11830
rect 13902 10842 13914 11818
rect 13948 10842 13964 11818
rect 13902 10830 13964 10842
rect 13994 11818 14056 11830
rect 13994 10842 14010 11818
rect 14044 10842 14056 11818
rect 13994 10830 14056 10842
rect 14112 11818 14174 11830
rect 14112 10842 14124 11818
rect 14158 10842 14174 11818
rect 14112 10830 14174 10842
rect 14204 11818 14266 11830
rect 14204 10842 14220 11818
rect 14254 10842 14266 11818
rect 14204 10830 14266 10842
rect 14322 11818 14384 11830
rect 14322 10842 14334 11818
rect 14368 10842 14384 11818
rect 14322 10830 14384 10842
rect 14414 11818 14476 11830
rect 14414 10842 14430 11818
rect 14464 10842 14476 11818
rect 14414 10830 14476 10842
rect 14532 11818 14594 11830
rect 14532 10842 14544 11818
rect 14578 10842 14594 11818
rect 14532 10830 14594 10842
rect 14624 11818 14686 11830
rect 14624 10842 14640 11818
rect 14674 10842 14686 11818
rect 14624 10830 14686 10842
rect 14742 11818 14804 11830
rect 14742 10842 14754 11818
rect 14788 10842 14804 11818
rect 14742 10830 14804 10842
rect 14834 11818 14896 11830
rect 14834 10842 14850 11818
rect 14884 10842 14896 11818
rect 14834 10830 14896 10842
rect 14952 11818 15014 11830
rect 14952 10842 14964 11818
rect 14998 10842 15014 11818
rect 14952 10830 15014 10842
rect 15044 11818 15106 11830
rect 15044 10842 15060 11818
rect 15094 10842 15106 11818
rect 15044 10830 15106 10842
rect 15162 11818 15224 11830
rect 15162 10842 15174 11818
rect 15208 10842 15224 11818
rect 15162 10830 15224 10842
rect 15254 11818 15316 11830
rect 15254 10842 15270 11818
rect 15304 10842 15316 11818
rect 15254 10830 15316 10842
rect 15372 11818 15434 11830
rect 15372 10842 15384 11818
rect 15418 10842 15434 11818
rect 15372 10830 15434 10842
rect 15464 11818 15526 11830
rect 15464 10842 15480 11818
rect 15514 10842 15526 11818
rect 15464 10830 15526 10842
rect 15582 11818 15644 11830
rect 15582 10842 15594 11818
rect 15628 10842 15644 11818
rect 15582 10830 15644 10842
rect 15674 11818 15736 11830
rect 15674 10842 15690 11818
rect 15724 10842 15736 11818
rect 15674 10830 15736 10842
rect 15792 11818 15854 11830
rect 15792 10842 15804 11818
rect 15838 10842 15854 11818
rect 15792 10830 15854 10842
rect 15884 11818 15946 11830
rect 15884 10842 15900 11818
rect 15934 10842 15946 11818
rect 15884 10830 15946 10842
rect 16002 11818 16064 11830
rect 16002 10842 16014 11818
rect 16048 10842 16064 11818
rect 16002 10830 16064 10842
rect 16094 11818 16156 11830
rect 16094 10842 16110 11818
rect 16144 10842 16156 11818
rect 16094 10830 16156 10842
rect 16212 11818 16274 11830
rect 16212 10842 16224 11818
rect 16258 10842 16274 11818
rect 16212 10830 16274 10842
rect 16304 11818 16366 11830
rect 16304 10842 16320 11818
rect 16354 10842 16366 11818
rect 16304 10830 16366 10842
rect 16422 11818 16484 11830
rect 16422 10842 16434 11818
rect 16468 10842 16484 11818
rect 16422 10830 16484 10842
rect 16514 11818 16576 11830
rect 16514 10842 16530 11818
rect 16564 10842 16576 11818
rect 16514 10830 16576 10842
rect 16632 11818 16694 11830
rect 16632 10842 16644 11818
rect 16678 10842 16694 11818
rect 16632 10830 16694 10842
rect 16724 11818 16786 11830
rect 16724 10842 16740 11818
rect 16774 10842 16786 11818
rect 16724 10830 16786 10842
rect 16842 11818 16904 11830
rect 16842 10842 16854 11818
rect 16888 10842 16904 11818
rect 16842 10830 16904 10842
rect 16934 11818 16996 11830
rect 16934 10842 16950 11818
rect 16984 10842 16996 11818
rect 16934 10830 16996 10842
rect 17052 11818 17114 11830
rect 17052 10842 17064 11818
rect 17098 10842 17114 11818
rect 17052 10830 17114 10842
rect 17144 11818 17206 11830
rect 17144 10842 17160 11818
rect 17194 10842 17206 11818
rect 17144 10830 17206 10842
rect 17262 11818 17324 11830
rect 17262 10842 17274 11818
rect 17308 10842 17324 11818
rect 17262 10830 17324 10842
rect 17354 11818 17416 11830
rect 17354 10842 17370 11818
rect 17404 10842 17416 11818
rect 17354 10830 17416 10842
rect 17472 11818 17534 11830
rect 17472 10842 17484 11818
rect 17518 10842 17534 11818
rect 17472 10830 17534 10842
rect 17564 11818 17626 11830
rect 17564 10842 17580 11818
rect 17614 10842 17626 11818
rect 17564 10830 17626 10842
rect 17682 11818 17744 11830
rect 17682 10842 17694 11818
rect 17728 10842 17744 11818
rect 17682 10830 17744 10842
rect 17774 11818 17836 11830
rect 17774 10842 17790 11818
rect 17824 10842 17836 11818
rect 17774 10830 17836 10842
rect 17892 11818 17954 11830
rect 17892 10842 17904 11818
rect 17938 10842 17954 11818
rect 17892 10830 17954 10842
rect 17984 11818 18046 11830
rect 17984 10842 18000 11818
rect 18034 10842 18046 11818
rect 17984 10830 18046 10842
rect 18102 11818 18164 11830
rect 18102 10842 18114 11818
rect 18148 10842 18164 11818
rect 18102 10830 18164 10842
rect 18194 11818 18256 11830
rect 18194 10842 18210 11818
rect 18244 10842 18256 11818
rect 18194 10830 18256 10842
rect 18312 11818 18374 11830
rect 18312 10842 18324 11818
rect 18358 10842 18374 11818
rect 18312 10830 18374 10842
rect 18404 11818 18466 11830
rect 18404 10842 18420 11818
rect 18454 10842 18466 11818
rect 18404 10830 18466 10842
rect 18522 11818 18584 11830
rect 18522 10842 18534 11818
rect 18568 10842 18584 11818
rect 18522 10830 18584 10842
rect 18614 11818 18676 11830
rect 18614 10842 18630 11818
rect 18664 10842 18676 11818
rect 18614 10830 18676 10842
rect 5482 6952 5544 6964
rect 5482 5976 5494 6952
rect 5528 5976 5544 6952
rect 5482 5964 5544 5976
rect 5574 6952 5636 6964
rect 5574 5976 5590 6952
rect 5624 5976 5636 6952
rect 5574 5964 5636 5976
rect 5692 6952 5754 6964
rect 5692 5976 5704 6952
rect 5738 5976 5754 6952
rect 5692 5964 5754 5976
rect 5784 6952 5846 6964
rect 5784 5976 5800 6952
rect 5834 5976 5846 6952
rect 5784 5964 5846 5976
rect 5902 6952 5964 6964
rect 5902 5976 5914 6952
rect 5948 5976 5964 6952
rect 5902 5964 5964 5976
rect 5994 6952 6056 6964
rect 5994 5976 6010 6952
rect 6044 5976 6056 6952
rect 5994 5964 6056 5976
rect 6112 6952 6174 6964
rect 6112 5976 6124 6952
rect 6158 5976 6174 6952
rect 6112 5964 6174 5976
rect 6204 6952 6266 6964
rect 6204 5976 6220 6952
rect 6254 5976 6266 6952
rect 6204 5964 6266 5976
rect 6322 6952 6384 6964
rect 6322 5976 6334 6952
rect 6368 5976 6384 6952
rect 6322 5964 6384 5976
rect 6414 6952 6476 6964
rect 6414 5976 6430 6952
rect 6464 5976 6476 6952
rect 6414 5964 6476 5976
rect 6532 6952 6594 6964
rect 6532 5976 6544 6952
rect 6578 5976 6594 6952
rect 6532 5964 6594 5976
rect 6624 6952 6686 6964
rect 6624 5976 6640 6952
rect 6674 5976 6686 6952
rect 6624 5964 6686 5976
rect 6742 6952 6804 6964
rect 6742 5976 6754 6952
rect 6788 5976 6804 6952
rect 6742 5964 6804 5976
rect 6834 6952 6896 6964
rect 6834 5976 6850 6952
rect 6884 5976 6896 6952
rect 6834 5964 6896 5976
rect 6952 6952 7014 6964
rect 6952 5976 6964 6952
rect 6998 5976 7014 6952
rect 6952 5964 7014 5976
rect 7044 6952 7106 6964
rect 7044 5976 7060 6952
rect 7094 5976 7106 6952
rect 7044 5964 7106 5976
rect 7162 6952 7224 6964
rect 7162 5976 7174 6952
rect 7208 5976 7224 6952
rect 7162 5964 7224 5976
rect 7254 6952 7316 6964
rect 7254 5976 7270 6952
rect 7304 5976 7316 6952
rect 7254 5964 7316 5976
rect 7372 6952 7434 6964
rect 7372 5976 7384 6952
rect 7418 5976 7434 6952
rect 7372 5964 7434 5976
rect 7464 6952 7526 6964
rect 7464 5976 7480 6952
rect 7514 5976 7526 6952
rect 7464 5964 7526 5976
rect 7582 6952 7644 6964
rect 7582 5976 7594 6952
rect 7628 5976 7644 6952
rect 7582 5964 7644 5976
rect 7674 6952 7736 6964
rect 7674 5976 7690 6952
rect 7724 5976 7736 6952
rect 7674 5964 7736 5976
rect 7792 6952 7854 6964
rect 7792 5976 7804 6952
rect 7838 5976 7854 6952
rect 7792 5964 7854 5976
rect 7884 6952 7946 6964
rect 7884 5976 7900 6952
rect 7934 5976 7946 6952
rect 7884 5964 7946 5976
rect 8002 6952 8064 6964
rect 8002 5976 8014 6952
rect 8048 5976 8064 6952
rect 8002 5964 8064 5976
rect 8094 6952 8156 6964
rect 8094 5976 8110 6952
rect 8144 5976 8156 6952
rect 8094 5964 8156 5976
rect 8212 6952 8274 6964
rect 8212 5976 8224 6952
rect 8258 5976 8274 6952
rect 8212 5964 8274 5976
rect 8304 6952 8366 6964
rect 8304 5976 8320 6952
rect 8354 5976 8366 6952
rect 8304 5964 8366 5976
rect 8422 6952 8484 6964
rect 8422 5976 8434 6952
rect 8468 5976 8484 6952
rect 8422 5964 8484 5976
rect 8514 6952 8576 6964
rect 8514 5976 8530 6952
rect 8564 5976 8576 6952
rect 8514 5964 8576 5976
rect 8632 6952 8694 6964
rect 8632 5976 8644 6952
rect 8678 5976 8694 6952
rect 8632 5964 8694 5976
rect 8724 6952 8786 6964
rect 8724 5976 8740 6952
rect 8774 5976 8786 6952
rect 8724 5964 8786 5976
rect 8842 6952 8904 6964
rect 8842 5976 8854 6952
rect 8888 5976 8904 6952
rect 8842 5964 8904 5976
rect 8934 6952 8996 6964
rect 8934 5976 8950 6952
rect 8984 5976 8996 6952
rect 8934 5964 8996 5976
rect 9052 6952 9114 6964
rect 9052 5976 9064 6952
rect 9098 5976 9114 6952
rect 9052 5964 9114 5976
rect 9144 6952 9206 6964
rect 9144 5976 9160 6952
rect 9194 5976 9206 6952
rect 9144 5964 9206 5976
rect 2574 5328 2632 5340
rect 2574 4352 2586 5328
rect 2620 4352 2632 5328
rect 2574 4340 2632 4352
rect 2662 5328 2720 5340
rect 2662 4352 2674 5328
rect 2708 4352 2720 5328
rect 3518 5328 3580 5340
rect 2662 4340 2720 4352
rect 3518 4352 3530 5328
rect 3564 4352 3580 5328
rect 3518 4340 3580 4352
rect 3610 5328 3672 5340
rect 3610 4352 3626 5328
rect 3660 4352 3672 5328
rect 3610 4340 3672 4352
rect 3728 5328 3790 5340
rect 3728 4352 3740 5328
rect 3774 4352 3790 5328
rect 3728 4340 3790 4352
rect 3820 5328 3882 5340
rect 3820 4352 3836 5328
rect 3870 4352 3882 5328
rect 3820 4340 3882 4352
rect 3938 5328 4000 5340
rect 3938 4352 3950 5328
rect 3984 4352 4000 5328
rect 3938 4340 4000 4352
rect 4030 5328 4092 5340
rect 4030 4352 4046 5328
rect 4080 4352 4092 5328
rect 4030 4340 4092 4352
rect 4148 5328 4210 5340
rect 4148 4352 4160 5328
rect 4194 4352 4210 5328
rect 4148 4340 4210 4352
rect 4240 5328 4302 5340
rect 4240 4352 4256 5328
rect 4290 4352 4302 5328
rect 4240 4340 4302 4352
rect 2574 -2826 2632 -2814
rect 2574 -3802 2586 -2826
rect 2620 -3802 2632 -2826
rect 2574 -3814 2632 -3802
rect 2662 -2826 2720 -2814
rect 2662 -3802 2674 -2826
rect 2708 -3802 2720 -2826
rect 3518 -2826 3580 -2814
rect 2662 -3814 2720 -3802
rect 3518 -3802 3530 -2826
rect 3564 -3802 3580 -2826
rect 3518 -3814 3580 -3802
rect 3610 -2826 3672 -2814
rect 3610 -3802 3626 -2826
rect 3660 -3802 3672 -2826
rect 3610 -3814 3672 -3802
rect 3728 -2826 3790 -2814
rect 3728 -3802 3740 -2826
rect 3774 -3802 3790 -2826
rect 3728 -3814 3790 -3802
rect 3820 -2826 3882 -2814
rect 3820 -3802 3836 -2826
rect 3870 -3802 3882 -2826
rect 3820 -3814 3882 -3802
rect 3938 -2826 4000 -2814
rect 3938 -3802 3950 -2826
rect 3984 -3802 4000 -2826
rect 3938 -3814 4000 -3802
rect 4030 -2826 4092 -2814
rect 4030 -3802 4046 -2826
rect 4080 -3802 4092 -2826
rect 4030 -3814 4092 -3802
rect 4148 -2826 4210 -2814
rect 4148 -3802 4160 -2826
rect 4194 -3802 4210 -2826
rect 4148 -3814 4210 -3802
rect 4240 -2826 4302 -2814
rect 4240 -3802 4256 -2826
rect 4290 -3802 4302 -2826
rect 4240 -3814 4302 -3802
rect 5482 -5850 5544 -5838
rect 5482 -6826 5494 -5850
rect 5528 -6826 5544 -5850
rect 5482 -6838 5544 -6826
rect 5574 -5850 5636 -5838
rect 5574 -6826 5590 -5850
rect 5624 -6826 5636 -5850
rect 5574 -6838 5636 -6826
rect 5692 -5850 5754 -5838
rect 5692 -6826 5704 -5850
rect 5738 -6826 5754 -5850
rect 5692 -6838 5754 -6826
rect 5784 -5850 5846 -5838
rect 5784 -6826 5800 -5850
rect 5834 -6826 5846 -5850
rect 5784 -6838 5846 -6826
rect 5902 -5850 5964 -5838
rect 5902 -6826 5914 -5850
rect 5948 -6826 5964 -5850
rect 5902 -6838 5964 -6826
rect 5994 -5850 6056 -5838
rect 5994 -6826 6010 -5850
rect 6044 -6826 6056 -5850
rect 5994 -6838 6056 -6826
rect 6112 -5850 6174 -5838
rect 6112 -6826 6124 -5850
rect 6158 -6826 6174 -5850
rect 6112 -6838 6174 -6826
rect 6204 -5850 6266 -5838
rect 6204 -6826 6220 -5850
rect 6254 -6826 6266 -5850
rect 6204 -6838 6266 -6826
rect 6322 -5850 6384 -5838
rect 6322 -6826 6334 -5850
rect 6368 -6826 6384 -5850
rect 6322 -6838 6384 -6826
rect 6414 -5850 6476 -5838
rect 6414 -6826 6430 -5850
rect 6464 -6826 6476 -5850
rect 6414 -6838 6476 -6826
rect 6532 -5850 6594 -5838
rect 6532 -6826 6544 -5850
rect 6578 -6826 6594 -5850
rect 6532 -6838 6594 -6826
rect 6624 -5850 6686 -5838
rect 6624 -6826 6640 -5850
rect 6674 -6826 6686 -5850
rect 6624 -6838 6686 -6826
rect 6742 -5850 6804 -5838
rect 6742 -6826 6754 -5850
rect 6788 -6826 6804 -5850
rect 6742 -6838 6804 -6826
rect 6834 -5850 6896 -5838
rect 6834 -6826 6850 -5850
rect 6884 -6826 6896 -5850
rect 6834 -6838 6896 -6826
rect 6952 -5850 7014 -5838
rect 6952 -6826 6964 -5850
rect 6998 -6826 7014 -5850
rect 6952 -6838 7014 -6826
rect 7044 -5850 7106 -5838
rect 7044 -6826 7060 -5850
rect 7094 -6826 7106 -5850
rect 7044 -6838 7106 -6826
rect 7162 -5850 7224 -5838
rect 7162 -6826 7174 -5850
rect 7208 -6826 7224 -5850
rect 7162 -6838 7224 -6826
rect 7254 -5850 7316 -5838
rect 7254 -6826 7270 -5850
rect 7304 -6826 7316 -5850
rect 7254 -6838 7316 -6826
rect 7372 -5850 7434 -5838
rect 7372 -6826 7384 -5850
rect 7418 -6826 7434 -5850
rect 7372 -6838 7434 -6826
rect 7464 -5850 7526 -5838
rect 7464 -6826 7480 -5850
rect 7514 -6826 7526 -5850
rect 7464 -6838 7526 -6826
rect 7582 -5850 7644 -5838
rect 7582 -6826 7594 -5850
rect 7628 -6826 7644 -5850
rect 7582 -6838 7644 -6826
rect 7674 -5850 7736 -5838
rect 7674 -6826 7690 -5850
rect 7724 -6826 7736 -5850
rect 7674 -6838 7736 -6826
rect 7792 -5850 7854 -5838
rect 7792 -6826 7804 -5850
rect 7838 -6826 7854 -5850
rect 7792 -6838 7854 -6826
rect 7884 -5850 7946 -5838
rect 7884 -6826 7900 -5850
rect 7934 -6826 7946 -5850
rect 7884 -6838 7946 -6826
rect 8002 -5850 8064 -5838
rect 8002 -6826 8014 -5850
rect 8048 -6826 8064 -5850
rect 8002 -6838 8064 -6826
rect 8094 -5850 8156 -5838
rect 8094 -6826 8110 -5850
rect 8144 -6826 8156 -5850
rect 8094 -6838 8156 -6826
rect 8212 -5850 8274 -5838
rect 8212 -6826 8224 -5850
rect 8258 -6826 8274 -5850
rect 8212 -6838 8274 -6826
rect 8304 -5850 8366 -5838
rect 8304 -6826 8320 -5850
rect 8354 -6826 8366 -5850
rect 8304 -6838 8366 -6826
rect 8422 -5850 8484 -5838
rect 8422 -6826 8434 -5850
rect 8468 -6826 8484 -5850
rect 8422 -6838 8484 -6826
rect 8514 -5850 8576 -5838
rect 8514 -6826 8530 -5850
rect 8564 -6826 8576 -5850
rect 8514 -6838 8576 -6826
rect 8632 -5850 8694 -5838
rect 8632 -6826 8644 -5850
rect 8678 -6826 8694 -5850
rect 8632 -6838 8694 -6826
rect 8724 -5850 8786 -5838
rect 8724 -6826 8740 -5850
rect 8774 -6826 8786 -5850
rect 8724 -6838 8786 -6826
rect 8842 -5850 8904 -5838
rect 8842 -6826 8854 -5850
rect 8888 -6826 8904 -5850
rect 8842 -6838 8904 -6826
rect 8934 -5850 8996 -5838
rect 8934 -6826 8950 -5850
rect 8984 -6826 8996 -5850
rect 8934 -6838 8996 -6826
rect 9052 -5850 9114 -5838
rect 9052 -6826 9064 -5850
rect 9098 -6826 9114 -5850
rect 9052 -6838 9114 -6826
rect 9144 -5850 9206 -5838
rect 9144 -6826 9160 -5850
rect 9194 -6826 9206 -5850
rect 9144 -6838 9206 -6826
<< pdiff >>
rect 2570 4100 2632 4112
rect 2570 3124 2582 4100
rect 2616 3124 2632 4100
rect 2570 3112 2632 3124
rect 2662 4100 2728 4112
rect 2662 3124 2678 4100
rect 2712 3124 2728 4100
rect 2662 3112 2728 3124
rect 2758 4100 2820 4112
rect 2758 3124 2774 4100
rect 2808 3124 2820 4100
rect 3308 4100 3370 4112
rect 2758 3112 2820 3124
rect 3308 3124 3320 4100
rect 3354 3124 3370 4100
rect 3308 3112 3370 3124
rect 3400 4100 3462 4112
rect 3400 3124 3416 4100
rect 3450 3124 3462 4100
rect 3400 3112 3462 3124
rect 3518 4100 3580 4112
rect 3518 3124 3530 4100
rect 3564 3124 3580 4100
rect 3518 3112 3580 3124
rect 3610 4100 3672 4112
rect 3610 3124 3626 4100
rect 3660 3124 3672 4100
rect 3610 3112 3672 3124
rect 3728 4100 3790 4112
rect 3728 3124 3740 4100
rect 3774 3124 3790 4100
rect 3728 3112 3790 3124
rect 3820 4100 3882 4112
rect 3820 3124 3836 4100
rect 3870 3124 3882 4100
rect 3820 3112 3882 3124
rect 3938 4100 4000 4112
rect 3938 3124 3950 4100
rect 3984 3124 4000 4100
rect 3938 3112 4000 3124
rect 4030 4100 4092 4112
rect 4030 3124 4046 4100
rect 4080 3124 4092 4100
rect 4030 3112 4092 3124
rect 4148 4100 4210 4112
rect 4148 3124 4160 4100
rect 4194 3124 4210 4100
rect 4148 3112 4210 3124
rect 4240 4100 4302 4112
rect 4240 3124 4256 4100
rect 4290 3124 4302 4100
rect 4240 3112 4302 3124
rect 4358 4100 4420 4112
rect 4358 3124 4370 4100
rect 4404 3124 4420 4100
rect 4358 3112 4420 3124
rect 4450 4100 4512 4112
rect 4450 3124 4466 4100
rect 4500 3124 4512 4100
rect 4450 3112 4512 3124
rect 4568 4100 4630 4112
rect 4568 3124 4580 4100
rect 4614 3124 4630 4100
rect 4568 3112 4630 3124
rect 4660 4100 4722 4112
rect 4660 3124 4676 4100
rect 4710 3124 4722 4100
rect 4660 3112 4722 3124
rect 4778 4100 4840 4112
rect 4778 3124 4790 4100
rect 4824 3124 4840 4100
rect 4778 3112 4840 3124
rect 4870 4100 4932 4112
rect 4870 3124 4886 4100
rect 4920 3124 4932 4100
rect 4870 3112 4932 3124
rect 5482 5336 5544 5348
rect 5482 4360 5494 5336
rect 5528 4360 5544 5336
rect 5482 4348 5544 4360
rect 5574 5336 5636 5348
rect 5574 4360 5590 5336
rect 5624 4360 5636 5336
rect 5574 4348 5636 4360
rect 5692 5336 5754 5348
rect 5692 4360 5704 5336
rect 5738 4360 5754 5336
rect 5692 4348 5754 4360
rect 5784 5336 5846 5348
rect 5784 4360 5800 5336
rect 5834 4360 5846 5336
rect 5784 4348 5846 4360
rect 5902 5336 5964 5348
rect 5902 4360 5914 5336
rect 5948 4360 5964 5336
rect 5902 4348 5964 4360
rect 5994 5336 6056 5348
rect 5994 4360 6010 5336
rect 6044 4360 6056 5336
rect 5994 4348 6056 4360
rect 6112 5336 6174 5348
rect 6112 4360 6124 5336
rect 6158 4360 6174 5336
rect 6112 4348 6174 4360
rect 6204 5336 6266 5348
rect 6204 4360 6220 5336
rect 6254 4360 6266 5336
rect 6204 4348 6266 4360
rect 6322 5336 6384 5348
rect 6322 4360 6334 5336
rect 6368 4360 6384 5336
rect 6322 4348 6384 4360
rect 6414 5336 6476 5348
rect 6414 4360 6430 5336
rect 6464 4360 6476 5336
rect 6414 4348 6476 4360
rect 6532 5336 6594 5348
rect 6532 4360 6544 5336
rect 6578 4360 6594 5336
rect 6532 4348 6594 4360
rect 6624 5336 6686 5348
rect 6624 4360 6640 5336
rect 6674 4360 6686 5336
rect 6624 4348 6686 4360
rect 6742 5336 6804 5348
rect 6742 4360 6754 5336
rect 6788 4360 6804 5336
rect 6742 4348 6804 4360
rect 6834 5336 6896 5348
rect 6834 4360 6850 5336
rect 6884 4360 6896 5336
rect 6834 4348 6896 4360
rect 6952 5336 7014 5348
rect 6952 4360 6964 5336
rect 6998 4360 7014 5336
rect 6952 4348 7014 4360
rect 7044 5336 7106 5348
rect 7044 4360 7060 5336
rect 7094 4360 7106 5336
rect 7044 4348 7106 4360
rect 7162 5336 7224 5348
rect 7162 4360 7174 5336
rect 7208 4360 7224 5336
rect 7162 4348 7224 4360
rect 7254 5336 7316 5348
rect 7254 4360 7270 5336
rect 7304 4360 7316 5336
rect 7254 4348 7316 4360
rect 7372 5336 7434 5348
rect 7372 4360 7384 5336
rect 7418 4360 7434 5336
rect 7372 4348 7434 4360
rect 7464 5336 7526 5348
rect 7464 4360 7480 5336
rect 7514 4360 7526 5336
rect 7464 4348 7526 4360
rect 7582 5336 7644 5348
rect 7582 4360 7594 5336
rect 7628 4360 7644 5336
rect 7582 4348 7644 4360
rect 7674 5336 7736 5348
rect 7674 4360 7690 5336
rect 7724 4360 7736 5336
rect 7674 4348 7736 4360
rect 7792 5336 7854 5348
rect 7792 4360 7804 5336
rect 7838 4360 7854 5336
rect 7792 4348 7854 4360
rect 7884 5336 7946 5348
rect 7884 4360 7900 5336
rect 7934 4360 7946 5336
rect 7884 4348 7946 4360
rect 8002 5336 8064 5348
rect 8002 4360 8014 5336
rect 8048 4360 8064 5336
rect 8002 4348 8064 4360
rect 8094 5336 8156 5348
rect 8094 4360 8110 5336
rect 8144 4360 8156 5336
rect 8094 4348 8156 4360
rect 8212 5336 8274 5348
rect 8212 4360 8224 5336
rect 8258 4360 8274 5336
rect 8212 4348 8274 4360
rect 8304 5336 8366 5348
rect 8304 4360 8320 5336
rect 8354 4360 8366 5336
rect 8304 4348 8366 4360
rect 8422 5336 8484 5348
rect 8422 4360 8434 5336
rect 8468 4360 8484 5336
rect 8422 4348 8484 4360
rect 8514 5336 8576 5348
rect 8514 4360 8530 5336
rect 8564 4360 8576 5336
rect 8514 4348 8576 4360
rect 8632 5336 8694 5348
rect 8632 4360 8644 5336
rect 8678 4360 8694 5336
rect 8632 4348 8694 4360
rect 8724 5336 8786 5348
rect 8724 4360 8740 5336
rect 8774 4360 8786 5336
rect 8724 4348 8786 4360
rect 8842 5336 8904 5348
rect 8842 4360 8854 5336
rect 8888 4360 8904 5336
rect 8842 4348 8904 4360
rect 8934 5336 8996 5348
rect 8934 4360 8950 5336
rect 8984 4360 8996 5336
rect 8934 4348 8996 4360
rect 9052 5336 9114 5348
rect 9052 4360 9064 5336
rect 9098 4360 9114 5336
rect 9052 4348 9114 4360
rect 9144 5336 9206 5348
rect 9144 4360 9160 5336
rect 9194 4360 9206 5336
rect 9144 4348 9206 4360
rect 5482 4100 5544 4112
rect 5482 3124 5494 4100
rect 5528 3124 5544 4100
rect 5482 3112 5544 3124
rect 5574 4100 5636 4112
rect 5574 3124 5590 4100
rect 5624 3124 5636 4100
rect 5574 3112 5636 3124
rect 5692 4100 5754 4112
rect 5692 3124 5704 4100
rect 5738 3124 5754 4100
rect 5692 3112 5754 3124
rect 5784 4100 5846 4112
rect 5784 3124 5800 4100
rect 5834 3124 5846 4100
rect 5784 3112 5846 3124
rect 5902 4100 5964 4112
rect 5902 3124 5914 4100
rect 5948 3124 5964 4100
rect 5902 3112 5964 3124
rect 5994 4100 6056 4112
rect 5994 3124 6010 4100
rect 6044 3124 6056 4100
rect 5994 3112 6056 3124
rect 6112 4100 6174 4112
rect 6112 3124 6124 4100
rect 6158 3124 6174 4100
rect 6112 3112 6174 3124
rect 6204 4100 6266 4112
rect 6204 3124 6220 4100
rect 6254 3124 6266 4100
rect 6204 3112 6266 3124
rect 6322 4100 6384 4112
rect 6322 3124 6334 4100
rect 6368 3124 6384 4100
rect 6322 3112 6384 3124
rect 6414 4100 6476 4112
rect 6414 3124 6430 4100
rect 6464 3124 6476 4100
rect 6414 3112 6476 3124
rect 6532 4100 6594 4112
rect 6532 3124 6544 4100
rect 6578 3124 6594 4100
rect 6532 3112 6594 3124
rect 6624 4100 6686 4112
rect 6624 3124 6640 4100
rect 6674 3124 6686 4100
rect 6624 3112 6686 3124
rect 6742 4100 6804 4112
rect 6742 3124 6754 4100
rect 6788 3124 6804 4100
rect 6742 3112 6804 3124
rect 6834 4100 6896 4112
rect 6834 3124 6850 4100
rect 6884 3124 6896 4100
rect 6834 3112 6896 3124
rect 6952 4100 7014 4112
rect 6952 3124 6964 4100
rect 6998 3124 7014 4100
rect 6952 3112 7014 3124
rect 7044 4100 7106 4112
rect 7044 3124 7060 4100
rect 7094 3124 7106 4100
rect 7044 3112 7106 3124
rect 7162 4100 7224 4112
rect 7162 3124 7174 4100
rect 7208 3124 7224 4100
rect 7162 3112 7224 3124
rect 7254 4100 7316 4112
rect 7254 3124 7270 4100
rect 7304 3124 7316 4100
rect 7254 3112 7316 3124
rect 7372 4100 7434 4112
rect 7372 3124 7384 4100
rect 7418 3124 7434 4100
rect 7372 3112 7434 3124
rect 7464 4100 7526 4112
rect 7464 3124 7480 4100
rect 7514 3124 7526 4100
rect 7464 3112 7526 3124
rect 7582 4100 7644 4112
rect 7582 3124 7594 4100
rect 7628 3124 7644 4100
rect 7582 3112 7644 3124
rect 7674 4100 7736 4112
rect 7674 3124 7690 4100
rect 7724 3124 7736 4100
rect 7674 3112 7736 3124
rect 7792 4100 7854 4112
rect 7792 3124 7804 4100
rect 7838 3124 7854 4100
rect 7792 3112 7854 3124
rect 7884 4100 7946 4112
rect 7884 3124 7900 4100
rect 7934 3124 7946 4100
rect 7884 3112 7946 3124
rect 8002 4100 8064 4112
rect 8002 3124 8014 4100
rect 8048 3124 8064 4100
rect 8002 3112 8064 3124
rect 8094 4100 8156 4112
rect 8094 3124 8110 4100
rect 8144 3124 8156 4100
rect 8094 3112 8156 3124
rect 8212 4100 8274 4112
rect 8212 3124 8224 4100
rect 8258 3124 8274 4100
rect 8212 3112 8274 3124
rect 8304 4100 8366 4112
rect 8304 3124 8320 4100
rect 8354 3124 8366 4100
rect 8304 3112 8366 3124
rect 8422 4100 8484 4112
rect 8422 3124 8434 4100
rect 8468 3124 8484 4100
rect 8422 3112 8484 3124
rect 8514 4100 8576 4112
rect 8514 3124 8530 4100
rect 8564 3124 8576 4100
rect 8514 3112 8576 3124
rect 8632 4100 8694 4112
rect 8632 3124 8644 4100
rect 8678 3124 8694 4100
rect 8632 3112 8694 3124
rect 8724 4100 8786 4112
rect 8724 3124 8740 4100
rect 8774 3124 8786 4100
rect 8724 3112 8786 3124
rect 8842 4100 8904 4112
rect 8842 3124 8854 4100
rect 8888 3124 8904 4100
rect 8842 3112 8904 3124
rect 8934 4100 8996 4112
rect 8934 3124 8950 4100
rect 8984 3124 8996 4100
rect 8934 3112 8996 3124
rect 9052 4100 9114 4112
rect 9052 3124 9064 4100
rect 9098 3124 9114 4100
rect 9052 3112 9114 3124
rect 9144 4100 9206 4112
rect 9144 3124 9160 4100
rect 9194 3124 9206 4100
rect 9144 3112 9206 3124
rect 10332 7808 10394 7820
rect 10332 6832 10344 7808
rect 10378 6832 10394 7808
rect 10332 6820 10394 6832
rect 10424 7808 10486 7820
rect 10424 6832 10440 7808
rect 10474 6832 10486 7808
rect 10424 6820 10486 6832
rect 10542 7808 10604 7820
rect 10542 6832 10554 7808
rect 10588 6832 10604 7808
rect 10542 6820 10604 6832
rect 10634 7808 10696 7820
rect 10634 6832 10650 7808
rect 10684 6832 10696 7808
rect 10634 6820 10696 6832
rect 10752 7808 10814 7820
rect 10752 6832 10764 7808
rect 10798 6832 10814 7808
rect 10752 6820 10814 6832
rect 10844 7808 10906 7820
rect 10844 6832 10860 7808
rect 10894 6832 10906 7808
rect 10844 6820 10906 6832
rect 10962 7808 11024 7820
rect 10962 6832 10974 7808
rect 11008 6832 11024 7808
rect 10962 6820 11024 6832
rect 11054 7808 11116 7820
rect 11054 6832 11070 7808
rect 11104 6832 11116 7808
rect 11054 6820 11116 6832
rect 11172 7808 11234 7820
rect 11172 6832 11184 7808
rect 11218 6832 11234 7808
rect 11172 6820 11234 6832
rect 11264 7808 11326 7820
rect 11264 6832 11280 7808
rect 11314 6832 11326 7808
rect 11264 6820 11326 6832
rect 11382 7808 11444 7820
rect 11382 6832 11394 7808
rect 11428 6832 11444 7808
rect 11382 6820 11444 6832
rect 11474 7808 11536 7820
rect 11474 6832 11490 7808
rect 11524 6832 11536 7808
rect 11474 6820 11536 6832
rect 11592 7808 11654 7820
rect 11592 6832 11604 7808
rect 11638 6832 11654 7808
rect 11592 6820 11654 6832
rect 11684 7808 11746 7820
rect 11684 6832 11700 7808
rect 11734 6832 11746 7808
rect 11684 6820 11746 6832
rect 11802 7808 11864 7820
rect 11802 6832 11814 7808
rect 11848 6832 11864 7808
rect 11802 6820 11864 6832
rect 11894 7808 11956 7820
rect 11894 6832 11910 7808
rect 11944 6832 11956 7808
rect 11894 6820 11956 6832
rect 12012 7808 12074 7820
rect 12012 6832 12024 7808
rect 12058 6832 12074 7808
rect 12012 6820 12074 6832
rect 12104 7808 12166 7820
rect 12104 6832 12120 7808
rect 12154 6832 12166 7808
rect 12104 6820 12166 6832
rect 12222 7808 12284 7820
rect 12222 6832 12234 7808
rect 12268 6832 12284 7808
rect 12222 6820 12284 6832
rect 12314 7808 12376 7820
rect 12314 6832 12330 7808
rect 12364 6832 12376 7808
rect 12314 6820 12376 6832
rect 12432 7808 12494 7820
rect 12432 6832 12444 7808
rect 12478 6832 12494 7808
rect 12432 6820 12494 6832
rect 12524 7808 12586 7820
rect 12524 6832 12540 7808
rect 12574 6832 12586 7808
rect 12524 6820 12586 6832
rect 12642 7808 12704 7820
rect 12642 6832 12654 7808
rect 12688 6832 12704 7808
rect 12642 6820 12704 6832
rect 12734 7808 12796 7820
rect 12734 6832 12750 7808
rect 12784 6832 12796 7808
rect 12734 6820 12796 6832
rect 12852 7808 12914 7820
rect 12852 6832 12864 7808
rect 12898 6832 12914 7808
rect 12852 6820 12914 6832
rect 12944 7808 13006 7820
rect 12944 6832 12960 7808
rect 12994 6832 13006 7808
rect 12944 6820 13006 6832
rect 13062 7808 13124 7820
rect 13062 6832 13074 7808
rect 13108 6832 13124 7808
rect 13062 6820 13124 6832
rect 13154 7808 13216 7820
rect 13154 6832 13170 7808
rect 13204 6832 13216 7808
rect 13154 6820 13216 6832
rect 13272 7808 13334 7820
rect 13272 6832 13284 7808
rect 13318 6832 13334 7808
rect 13272 6820 13334 6832
rect 13364 7808 13426 7820
rect 13364 6832 13380 7808
rect 13414 6832 13426 7808
rect 13364 6820 13426 6832
rect 13482 7808 13544 7820
rect 13482 6832 13494 7808
rect 13528 6832 13544 7808
rect 13482 6820 13544 6832
rect 13574 7808 13636 7820
rect 13574 6832 13590 7808
rect 13624 6832 13636 7808
rect 13574 6820 13636 6832
rect 13692 7808 13754 7820
rect 13692 6832 13704 7808
rect 13738 6832 13754 7808
rect 13692 6820 13754 6832
rect 13784 7808 13846 7820
rect 13784 6832 13800 7808
rect 13834 6832 13846 7808
rect 13784 6820 13846 6832
rect 13902 7808 13964 7820
rect 13902 6832 13914 7808
rect 13948 6832 13964 7808
rect 13902 6820 13964 6832
rect 13994 7808 14056 7820
rect 13994 6832 14010 7808
rect 14044 6832 14056 7808
rect 13994 6820 14056 6832
rect 14112 7808 14174 7820
rect 14112 6832 14124 7808
rect 14158 6832 14174 7808
rect 14112 6820 14174 6832
rect 14204 7808 14266 7820
rect 14204 6832 14220 7808
rect 14254 6832 14266 7808
rect 14204 6820 14266 6832
rect 14322 7808 14384 7820
rect 14322 6832 14334 7808
rect 14368 6832 14384 7808
rect 14322 6820 14384 6832
rect 14414 7808 14476 7820
rect 14414 6832 14430 7808
rect 14464 6832 14476 7808
rect 14414 6820 14476 6832
rect 14532 7808 14594 7820
rect 14532 6832 14544 7808
rect 14578 6832 14594 7808
rect 14532 6820 14594 6832
rect 14624 7808 14686 7820
rect 14624 6832 14640 7808
rect 14674 6832 14686 7808
rect 14624 6820 14686 6832
rect 14742 7808 14804 7820
rect 14742 6832 14754 7808
rect 14788 6832 14804 7808
rect 14742 6820 14804 6832
rect 14834 7808 14896 7820
rect 14834 6832 14850 7808
rect 14884 6832 14896 7808
rect 14834 6820 14896 6832
rect 14952 7808 15014 7820
rect 14952 6832 14964 7808
rect 14998 6832 15014 7808
rect 14952 6820 15014 6832
rect 15044 7808 15106 7820
rect 15044 6832 15060 7808
rect 15094 6832 15106 7808
rect 15044 6820 15106 6832
rect 15162 7808 15224 7820
rect 15162 6832 15174 7808
rect 15208 6832 15224 7808
rect 15162 6820 15224 6832
rect 15254 7808 15316 7820
rect 15254 6832 15270 7808
rect 15304 6832 15316 7808
rect 15254 6820 15316 6832
rect 15372 7808 15434 7820
rect 15372 6832 15384 7808
rect 15418 6832 15434 7808
rect 15372 6820 15434 6832
rect 15464 7808 15526 7820
rect 15464 6832 15480 7808
rect 15514 6832 15526 7808
rect 15464 6820 15526 6832
rect 15582 7808 15644 7820
rect 15582 6832 15594 7808
rect 15628 6832 15644 7808
rect 15582 6820 15644 6832
rect 15674 7808 15736 7820
rect 15674 6832 15690 7808
rect 15724 6832 15736 7808
rect 15674 6820 15736 6832
rect 15792 7808 15854 7820
rect 15792 6832 15804 7808
rect 15838 6832 15854 7808
rect 15792 6820 15854 6832
rect 15884 7808 15946 7820
rect 15884 6832 15900 7808
rect 15934 6832 15946 7808
rect 15884 6820 15946 6832
rect 16002 7808 16064 7820
rect 16002 6832 16014 7808
rect 16048 6832 16064 7808
rect 16002 6820 16064 6832
rect 16094 7808 16156 7820
rect 16094 6832 16110 7808
rect 16144 6832 16156 7808
rect 16094 6820 16156 6832
rect 16212 7808 16274 7820
rect 16212 6832 16224 7808
rect 16258 6832 16274 7808
rect 16212 6820 16274 6832
rect 16304 7808 16366 7820
rect 16304 6832 16320 7808
rect 16354 6832 16366 7808
rect 16304 6820 16366 6832
rect 16422 7808 16484 7820
rect 16422 6832 16434 7808
rect 16468 6832 16484 7808
rect 16422 6820 16484 6832
rect 16514 7808 16576 7820
rect 16514 6832 16530 7808
rect 16564 6832 16576 7808
rect 16514 6820 16576 6832
rect 16632 7808 16694 7820
rect 16632 6832 16644 7808
rect 16678 6832 16694 7808
rect 16632 6820 16694 6832
rect 16724 7808 16786 7820
rect 16724 6832 16740 7808
rect 16774 6832 16786 7808
rect 16724 6820 16786 6832
rect 16842 7808 16904 7820
rect 16842 6832 16854 7808
rect 16888 6832 16904 7808
rect 16842 6820 16904 6832
rect 16934 7808 16996 7820
rect 16934 6832 16950 7808
rect 16984 6832 16996 7808
rect 16934 6820 16996 6832
rect 17052 7808 17114 7820
rect 17052 6832 17064 7808
rect 17098 6832 17114 7808
rect 17052 6820 17114 6832
rect 17144 7808 17206 7820
rect 17144 6832 17160 7808
rect 17194 6832 17206 7808
rect 17144 6820 17206 6832
rect 17262 7808 17324 7820
rect 17262 6832 17274 7808
rect 17308 6832 17324 7808
rect 17262 6820 17324 6832
rect 17354 7808 17416 7820
rect 17354 6832 17370 7808
rect 17404 6832 17416 7808
rect 17354 6820 17416 6832
rect 17472 7808 17534 7820
rect 17472 6832 17484 7808
rect 17518 6832 17534 7808
rect 17472 6820 17534 6832
rect 17564 7808 17626 7820
rect 17564 6832 17580 7808
rect 17614 6832 17626 7808
rect 17564 6820 17626 6832
rect 17682 7808 17744 7820
rect 17682 6832 17694 7808
rect 17728 6832 17744 7808
rect 17682 6820 17744 6832
rect 17774 7808 17836 7820
rect 17774 6832 17790 7808
rect 17824 6832 17836 7808
rect 17774 6820 17836 6832
rect 17892 7808 17954 7820
rect 17892 6832 17904 7808
rect 17938 6832 17954 7808
rect 17892 6820 17954 6832
rect 17984 7808 18046 7820
rect 17984 6832 18000 7808
rect 18034 6832 18046 7808
rect 17984 6820 18046 6832
rect 18102 7808 18164 7820
rect 18102 6832 18114 7808
rect 18148 6832 18164 7808
rect 18102 6820 18164 6832
rect 18194 7808 18256 7820
rect 18194 6832 18210 7808
rect 18244 6832 18256 7808
rect 18194 6820 18256 6832
rect 18312 7808 18374 7820
rect 18312 6832 18324 7808
rect 18358 6832 18374 7808
rect 18312 6820 18374 6832
rect 18404 7808 18466 7820
rect 18404 6832 18420 7808
rect 18454 6832 18466 7808
rect 18404 6820 18466 6832
rect 18522 7808 18584 7820
rect 18522 6832 18534 7808
rect 18568 6832 18584 7808
rect 18522 6820 18584 6832
rect 18614 7808 18676 7820
rect 18614 6832 18630 7808
rect 18664 6832 18676 7808
rect 18614 6820 18676 6832
rect 10332 6572 10394 6584
rect 10332 5596 10344 6572
rect 10378 5596 10394 6572
rect 10332 5584 10394 5596
rect 10424 6572 10486 6584
rect 10424 5596 10440 6572
rect 10474 5596 10486 6572
rect 10424 5584 10486 5596
rect 10542 6572 10604 6584
rect 10542 5596 10554 6572
rect 10588 5596 10604 6572
rect 10542 5584 10604 5596
rect 10634 6572 10696 6584
rect 10634 5596 10650 6572
rect 10684 5596 10696 6572
rect 10634 5584 10696 5596
rect 10752 6572 10814 6584
rect 10752 5596 10764 6572
rect 10798 5596 10814 6572
rect 10752 5584 10814 5596
rect 10844 6572 10906 6584
rect 10844 5596 10860 6572
rect 10894 5596 10906 6572
rect 10844 5584 10906 5596
rect 10962 6572 11024 6584
rect 10962 5596 10974 6572
rect 11008 5596 11024 6572
rect 10962 5584 11024 5596
rect 11054 6572 11116 6584
rect 11054 5596 11070 6572
rect 11104 5596 11116 6572
rect 11054 5584 11116 5596
rect 11172 6572 11234 6584
rect 11172 5596 11184 6572
rect 11218 5596 11234 6572
rect 11172 5584 11234 5596
rect 11264 6572 11326 6584
rect 11264 5596 11280 6572
rect 11314 5596 11326 6572
rect 11264 5584 11326 5596
rect 11382 6572 11444 6584
rect 11382 5596 11394 6572
rect 11428 5596 11444 6572
rect 11382 5584 11444 5596
rect 11474 6572 11536 6584
rect 11474 5596 11490 6572
rect 11524 5596 11536 6572
rect 11474 5584 11536 5596
rect 11592 6572 11654 6584
rect 11592 5596 11604 6572
rect 11638 5596 11654 6572
rect 11592 5584 11654 5596
rect 11684 6572 11746 6584
rect 11684 5596 11700 6572
rect 11734 5596 11746 6572
rect 11684 5584 11746 5596
rect 11802 6572 11864 6584
rect 11802 5596 11814 6572
rect 11848 5596 11864 6572
rect 11802 5584 11864 5596
rect 11894 6572 11956 6584
rect 11894 5596 11910 6572
rect 11944 5596 11956 6572
rect 11894 5584 11956 5596
rect 12012 6572 12074 6584
rect 12012 5596 12024 6572
rect 12058 5596 12074 6572
rect 12012 5584 12074 5596
rect 12104 6572 12166 6584
rect 12104 5596 12120 6572
rect 12154 5596 12166 6572
rect 12104 5584 12166 5596
rect 12222 6572 12284 6584
rect 12222 5596 12234 6572
rect 12268 5596 12284 6572
rect 12222 5584 12284 5596
rect 12314 6572 12376 6584
rect 12314 5596 12330 6572
rect 12364 5596 12376 6572
rect 12314 5584 12376 5596
rect 12432 6572 12494 6584
rect 12432 5596 12444 6572
rect 12478 5596 12494 6572
rect 12432 5584 12494 5596
rect 12524 6572 12586 6584
rect 12524 5596 12540 6572
rect 12574 5596 12586 6572
rect 12524 5584 12586 5596
rect 12642 6572 12704 6584
rect 12642 5596 12654 6572
rect 12688 5596 12704 6572
rect 12642 5584 12704 5596
rect 12734 6572 12796 6584
rect 12734 5596 12750 6572
rect 12784 5596 12796 6572
rect 12734 5584 12796 5596
rect 12852 6572 12914 6584
rect 12852 5596 12864 6572
rect 12898 5596 12914 6572
rect 12852 5584 12914 5596
rect 12944 6572 13006 6584
rect 12944 5596 12960 6572
rect 12994 5596 13006 6572
rect 12944 5584 13006 5596
rect 13062 6572 13124 6584
rect 13062 5596 13074 6572
rect 13108 5596 13124 6572
rect 13062 5584 13124 5596
rect 13154 6572 13216 6584
rect 13154 5596 13170 6572
rect 13204 5596 13216 6572
rect 13154 5584 13216 5596
rect 13272 6572 13334 6584
rect 13272 5596 13284 6572
rect 13318 5596 13334 6572
rect 13272 5584 13334 5596
rect 13364 6572 13426 6584
rect 13364 5596 13380 6572
rect 13414 5596 13426 6572
rect 13364 5584 13426 5596
rect 13482 6572 13544 6584
rect 13482 5596 13494 6572
rect 13528 5596 13544 6572
rect 13482 5584 13544 5596
rect 13574 6572 13636 6584
rect 13574 5596 13590 6572
rect 13624 5596 13636 6572
rect 13574 5584 13636 5596
rect 13692 6572 13754 6584
rect 13692 5596 13704 6572
rect 13738 5596 13754 6572
rect 13692 5584 13754 5596
rect 13784 6572 13846 6584
rect 13784 5596 13800 6572
rect 13834 5596 13846 6572
rect 13784 5584 13846 5596
rect 13902 6572 13964 6584
rect 13902 5596 13914 6572
rect 13948 5596 13964 6572
rect 13902 5584 13964 5596
rect 13994 6572 14056 6584
rect 13994 5596 14010 6572
rect 14044 5596 14056 6572
rect 13994 5584 14056 5596
rect 14112 6572 14174 6584
rect 14112 5596 14124 6572
rect 14158 5596 14174 6572
rect 14112 5584 14174 5596
rect 14204 6572 14266 6584
rect 14204 5596 14220 6572
rect 14254 5596 14266 6572
rect 14204 5584 14266 5596
rect 14322 6572 14384 6584
rect 14322 5596 14334 6572
rect 14368 5596 14384 6572
rect 14322 5584 14384 5596
rect 14414 6572 14476 6584
rect 14414 5596 14430 6572
rect 14464 5596 14476 6572
rect 14414 5584 14476 5596
rect 14532 6572 14594 6584
rect 14532 5596 14544 6572
rect 14578 5596 14594 6572
rect 14532 5584 14594 5596
rect 14624 6572 14686 6584
rect 14624 5596 14640 6572
rect 14674 5596 14686 6572
rect 14624 5584 14686 5596
rect 14742 6572 14804 6584
rect 14742 5596 14754 6572
rect 14788 5596 14804 6572
rect 14742 5584 14804 5596
rect 14834 6572 14896 6584
rect 14834 5596 14850 6572
rect 14884 5596 14896 6572
rect 14834 5584 14896 5596
rect 14952 6572 15014 6584
rect 14952 5596 14964 6572
rect 14998 5596 15014 6572
rect 14952 5584 15014 5596
rect 15044 6572 15106 6584
rect 15044 5596 15060 6572
rect 15094 5596 15106 6572
rect 15044 5584 15106 5596
rect 15162 6572 15224 6584
rect 15162 5596 15174 6572
rect 15208 5596 15224 6572
rect 15162 5584 15224 5596
rect 15254 6572 15316 6584
rect 15254 5596 15270 6572
rect 15304 5596 15316 6572
rect 15254 5584 15316 5596
rect 15372 6572 15434 6584
rect 15372 5596 15384 6572
rect 15418 5596 15434 6572
rect 15372 5584 15434 5596
rect 15464 6572 15526 6584
rect 15464 5596 15480 6572
rect 15514 5596 15526 6572
rect 15464 5584 15526 5596
rect 15582 6572 15644 6584
rect 15582 5596 15594 6572
rect 15628 5596 15644 6572
rect 15582 5584 15644 5596
rect 15674 6572 15736 6584
rect 15674 5596 15690 6572
rect 15724 5596 15736 6572
rect 15674 5584 15736 5596
rect 15792 6572 15854 6584
rect 15792 5596 15804 6572
rect 15838 5596 15854 6572
rect 15792 5584 15854 5596
rect 15884 6572 15946 6584
rect 15884 5596 15900 6572
rect 15934 5596 15946 6572
rect 15884 5584 15946 5596
rect 16002 6572 16064 6584
rect 16002 5596 16014 6572
rect 16048 5596 16064 6572
rect 16002 5584 16064 5596
rect 16094 6572 16156 6584
rect 16094 5596 16110 6572
rect 16144 5596 16156 6572
rect 16094 5584 16156 5596
rect 16212 6572 16274 6584
rect 16212 5596 16224 6572
rect 16258 5596 16274 6572
rect 16212 5584 16274 5596
rect 16304 6572 16366 6584
rect 16304 5596 16320 6572
rect 16354 5596 16366 6572
rect 16304 5584 16366 5596
rect 16422 6572 16484 6584
rect 16422 5596 16434 6572
rect 16468 5596 16484 6572
rect 16422 5584 16484 5596
rect 16514 6572 16576 6584
rect 16514 5596 16530 6572
rect 16564 5596 16576 6572
rect 16514 5584 16576 5596
rect 16632 6572 16694 6584
rect 16632 5596 16644 6572
rect 16678 5596 16694 6572
rect 16632 5584 16694 5596
rect 16724 6572 16786 6584
rect 16724 5596 16740 6572
rect 16774 5596 16786 6572
rect 16724 5584 16786 5596
rect 16842 6572 16904 6584
rect 16842 5596 16854 6572
rect 16888 5596 16904 6572
rect 16842 5584 16904 5596
rect 16934 6572 16996 6584
rect 16934 5596 16950 6572
rect 16984 5596 16996 6572
rect 16934 5584 16996 5596
rect 17052 6572 17114 6584
rect 17052 5596 17064 6572
rect 17098 5596 17114 6572
rect 17052 5584 17114 5596
rect 17144 6572 17206 6584
rect 17144 5596 17160 6572
rect 17194 5596 17206 6572
rect 17144 5584 17206 5596
rect 17262 6572 17324 6584
rect 17262 5596 17274 6572
rect 17308 5596 17324 6572
rect 17262 5584 17324 5596
rect 17354 6572 17416 6584
rect 17354 5596 17370 6572
rect 17404 5596 17416 6572
rect 17354 5584 17416 5596
rect 17472 6572 17534 6584
rect 17472 5596 17484 6572
rect 17518 5596 17534 6572
rect 17472 5584 17534 5596
rect 17564 6572 17626 6584
rect 17564 5596 17580 6572
rect 17614 5596 17626 6572
rect 17564 5584 17626 5596
rect 17682 6572 17744 6584
rect 17682 5596 17694 6572
rect 17728 5596 17744 6572
rect 17682 5584 17744 5596
rect 17774 6572 17836 6584
rect 17774 5596 17790 6572
rect 17824 5596 17836 6572
rect 17774 5584 17836 5596
rect 17892 6572 17954 6584
rect 17892 5596 17904 6572
rect 17938 5596 17954 6572
rect 17892 5584 17954 5596
rect 17984 6572 18046 6584
rect 17984 5596 18000 6572
rect 18034 5596 18046 6572
rect 17984 5584 18046 5596
rect 18102 6572 18164 6584
rect 18102 5596 18114 6572
rect 18148 5596 18164 6572
rect 18102 5584 18164 5596
rect 18194 6572 18256 6584
rect 18194 5596 18210 6572
rect 18244 5596 18256 6572
rect 18194 5584 18256 5596
rect 18312 6572 18374 6584
rect 18312 5596 18324 6572
rect 18358 5596 18374 6572
rect 18312 5584 18374 5596
rect 18404 6572 18466 6584
rect 18404 5596 18420 6572
rect 18454 5596 18466 6572
rect 18404 5584 18466 5596
rect 18522 6572 18584 6584
rect 18522 5596 18534 6572
rect 18568 5596 18584 6572
rect 18522 5584 18584 5596
rect 18614 6572 18676 6584
rect 18614 5596 18630 6572
rect 18664 5596 18676 6572
rect 18614 5584 18676 5596
rect 10332 5336 10394 5348
rect 10332 4360 10344 5336
rect 10378 4360 10394 5336
rect 10332 4348 10394 4360
rect 10424 5336 10486 5348
rect 10424 4360 10440 5336
rect 10474 4360 10486 5336
rect 10424 4348 10486 4360
rect 10542 5336 10604 5348
rect 10542 4360 10554 5336
rect 10588 4360 10604 5336
rect 10542 4348 10604 4360
rect 10634 5336 10696 5348
rect 10634 4360 10650 5336
rect 10684 4360 10696 5336
rect 10634 4348 10696 4360
rect 10752 5336 10814 5348
rect 10752 4360 10764 5336
rect 10798 4360 10814 5336
rect 10752 4348 10814 4360
rect 10844 5336 10906 5348
rect 10844 4360 10860 5336
rect 10894 4360 10906 5336
rect 10844 4348 10906 4360
rect 10962 5336 11024 5348
rect 10962 4360 10974 5336
rect 11008 4360 11024 5336
rect 10962 4348 11024 4360
rect 11054 5336 11116 5348
rect 11054 4360 11070 5336
rect 11104 4360 11116 5336
rect 11054 4348 11116 4360
rect 11172 5336 11234 5348
rect 11172 4360 11184 5336
rect 11218 4360 11234 5336
rect 11172 4348 11234 4360
rect 11264 5336 11326 5348
rect 11264 4360 11280 5336
rect 11314 4360 11326 5336
rect 11264 4348 11326 4360
rect 11382 5336 11444 5348
rect 11382 4360 11394 5336
rect 11428 4360 11444 5336
rect 11382 4348 11444 4360
rect 11474 5336 11536 5348
rect 11474 4360 11490 5336
rect 11524 4360 11536 5336
rect 11474 4348 11536 4360
rect 11592 5336 11654 5348
rect 11592 4360 11604 5336
rect 11638 4360 11654 5336
rect 11592 4348 11654 4360
rect 11684 5336 11746 5348
rect 11684 4360 11700 5336
rect 11734 4360 11746 5336
rect 11684 4348 11746 4360
rect 11802 5336 11864 5348
rect 11802 4360 11814 5336
rect 11848 4360 11864 5336
rect 11802 4348 11864 4360
rect 11894 5336 11956 5348
rect 11894 4360 11910 5336
rect 11944 4360 11956 5336
rect 11894 4348 11956 4360
rect 12012 5336 12074 5348
rect 12012 4360 12024 5336
rect 12058 4360 12074 5336
rect 12012 4348 12074 4360
rect 12104 5336 12166 5348
rect 12104 4360 12120 5336
rect 12154 4360 12166 5336
rect 12104 4348 12166 4360
rect 12222 5336 12284 5348
rect 12222 4360 12234 5336
rect 12268 4360 12284 5336
rect 12222 4348 12284 4360
rect 12314 5336 12376 5348
rect 12314 4360 12330 5336
rect 12364 4360 12376 5336
rect 12314 4348 12376 4360
rect 12432 5336 12494 5348
rect 12432 4360 12444 5336
rect 12478 4360 12494 5336
rect 12432 4348 12494 4360
rect 12524 5336 12586 5348
rect 12524 4360 12540 5336
rect 12574 4360 12586 5336
rect 12524 4348 12586 4360
rect 12642 5336 12704 5348
rect 12642 4360 12654 5336
rect 12688 4360 12704 5336
rect 12642 4348 12704 4360
rect 12734 5336 12796 5348
rect 12734 4360 12750 5336
rect 12784 4360 12796 5336
rect 12734 4348 12796 4360
rect 12852 5336 12914 5348
rect 12852 4360 12864 5336
rect 12898 4360 12914 5336
rect 12852 4348 12914 4360
rect 12944 5336 13006 5348
rect 12944 4360 12960 5336
rect 12994 4360 13006 5336
rect 12944 4348 13006 4360
rect 13062 5336 13124 5348
rect 13062 4360 13074 5336
rect 13108 4360 13124 5336
rect 13062 4348 13124 4360
rect 13154 5336 13216 5348
rect 13154 4360 13170 5336
rect 13204 4360 13216 5336
rect 13154 4348 13216 4360
rect 13272 5336 13334 5348
rect 13272 4360 13284 5336
rect 13318 4360 13334 5336
rect 13272 4348 13334 4360
rect 13364 5336 13426 5348
rect 13364 4360 13380 5336
rect 13414 4360 13426 5336
rect 13364 4348 13426 4360
rect 13482 5336 13544 5348
rect 13482 4360 13494 5336
rect 13528 4360 13544 5336
rect 13482 4348 13544 4360
rect 13574 5336 13636 5348
rect 13574 4360 13590 5336
rect 13624 4360 13636 5336
rect 13574 4348 13636 4360
rect 13692 5336 13754 5348
rect 13692 4360 13704 5336
rect 13738 4360 13754 5336
rect 13692 4348 13754 4360
rect 13784 5336 13846 5348
rect 13784 4360 13800 5336
rect 13834 4360 13846 5336
rect 13784 4348 13846 4360
rect 13902 5336 13964 5348
rect 13902 4360 13914 5336
rect 13948 4360 13964 5336
rect 13902 4348 13964 4360
rect 13994 5336 14056 5348
rect 13994 4360 14010 5336
rect 14044 4360 14056 5336
rect 13994 4348 14056 4360
rect 14112 5336 14174 5348
rect 14112 4360 14124 5336
rect 14158 4360 14174 5336
rect 14112 4348 14174 4360
rect 14204 5336 14266 5348
rect 14204 4360 14220 5336
rect 14254 4360 14266 5336
rect 14204 4348 14266 4360
rect 14322 5336 14384 5348
rect 14322 4360 14334 5336
rect 14368 4360 14384 5336
rect 14322 4348 14384 4360
rect 14414 5336 14476 5348
rect 14414 4360 14430 5336
rect 14464 4360 14476 5336
rect 14414 4348 14476 4360
rect 14532 5336 14594 5348
rect 14532 4360 14544 5336
rect 14578 4360 14594 5336
rect 14532 4348 14594 4360
rect 14624 5336 14686 5348
rect 14624 4360 14640 5336
rect 14674 4360 14686 5336
rect 14624 4348 14686 4360
rect 14742 5336 14804 5348
rect 14742 4360 14754 5336
rect 14788 4360 14804 5336
rect 14742 4348 14804 4360
rect 14834 5336 14896 5348
rect 14834 4360 14850 5336
rect 14884 4360 14896 5336
rect 14834 4348 14896 4360
rect 14952 5336 15014 5348
rect 14952 4360 14964 5336
rect 14998 4360 15014 5336
rect 14952 4348 15014 4360
rect 15044 5336 15106 5348
rect 15044 4360 15060 5336
rect 15094 4360 15106 5336
rect 15044 4348 15106 4360
rect 15162 5336 15224 5348
rect 15162 4360 15174 5336
rect 15208 4360 15224 5336
rect 15162 4348 15224 4360
rect 15254 5336 15316 5348
rect 15254 4360 15270 5336
rect 15304 4360 15316 5336
rect 15254 4348 15316 4360
rect 15372 5336 15434 5348
rect 15372 4360 15384 5336
rect 15418 4360 15434 5336
rect 15372 4348 15434 4360
rect 15464 5336 15526 5348
rect 15464 4360 15480 5336
rect 15514 4360 15526 5336
rect 15464 4348 15526 4360
rect 15582 5336 15644 5348
rect 15582 4360 15594 5336
rect 15628 4360 15644 5336
rect 15582 4348 15644 4360
rect 15674 5336 15736 5348
rect 15674 4360 15690 5336
rect 15724 4360 15736 5336
rect 15674 4348 15736 4360
rect 15792 5336 15854 5348
rect 15792 4360 15804 5336
rect 15838 4360 15854 5336
rect 15792 4348 15854 4360
rect 15884 5336 15946 5348
rect 15884 4360 15900 5336
rect 15934 4360 15946 5336
rect 15884 4348 15946 4360
rect 16002 5336 16064 5348
rect 16002 4360 16014 5336
rect 16048 4360 16064 5336
rect 16002 4348 16064 4360
rect 16094 5336 16156 5348
rect 16094 4360 16110 5336
rect 16144 4360 16156 5336
rect 16094 4348 16156 4360
rect 16212 5336 16274 5348
rect 16212 4360 16224 5336
rect 16258 4360 16274 5336
rect 16212 4348 16274 4360
rect 16304 5336 16366 5348
rect 16304 4360 16320 5336
rect 16354 4360 16366 5336
rect 16304 4348 16366 4360
rect 16422 5336 16484 5348
rect 16422 4360 16434 5336
rect 16468 4360 16484 5336
rect 16422 4348 16484 4360
rect 16514 5336 16576 5348
rect 16514 4360 16530 5336
rect 16564 4360 16576 5336
rect 16514 4348 16576 4360
rect 16632 5336 16694 5348
rect 16632 4360 16644 5336
rect 16678 4360 16694 5336
rect 16632 4348 16694 4360
rect 16724 5336 16786 5348
rect 16724 4360 16740 5336
rect 16774 4360 16786 5336
rect 16724 4348 16786 4360
rect 16842 5336 16904 5348
rect 16842 4360 16854 5336
rect 16888 4360 16904 5336
rect 16842 4348 16904 4360
rect 16934 5336 16996 5348
rect 16934 4360 16950 5336
rect 16984 4360 16996 5336
rect 16934 4348 16996 4360
rect 17052 5336 17114 5348
rect 17052 4360 17064 5336
rect 17098 4360 17114 5336
rect 17052 4348 17114 4360
rect 17144 5336 17206 5348
rect 17144 4360 17160 5336
rect 17194 4360 17206 5336
rect 17144 4348 17206 4360
rect 17262 5336 17324 5348
rect 17262 4360 17274 5336
rect 17308 4360 17324 5336
rect 17262 4348 17324 4360
rect 17354 5336 17416 5348
rect 17354 4360 17370 5336
rect 17404 4360 17416 5336
rect 17354 4348 17416 4360
rect 17472 5336 17534 5348
rect 17472 4360 17484 5336
rect 17518 4360 17534 5336
rect 17472 4348 17534 4360
rect 17564 5336 17626 5348
rect 17564 4360 17580 5336
rect 17614 4360 17626 5336
rect 17564 4348 17626 4360
rect 17682 5336 17744 5348
rect 17682 4360 17694 5336
rect 17728 4360 17744 5336
rect 17682 4348 17744 4360
rect 17774 5336 17836 5348
rect 17774 4360 17790 5336
rect 17824 4360 17836 5336
rect 17774 4348 17836 4360
rect 17892 5336 17954 5348
rect 17892 4360 17904 5336
rect 17938 4360 17954 5336
rect 17892 4348 17954 4360
rect 17984 5336 18046 5348
rect 17984 4360 18000 5336
rect 18034 4360 18046 5336
rect 17984 4348 18046 4360
rect 18102 5336 18164 5348
rect 18102 4360 18114 5336
rect 18148 4360 18164 5336
rect 18102 4348 18164 4360
rect 18194 5336 18256 5348
rect 18194 4360 18210 5336
rect 18244 4360 18256 5336
rect 18194 4348 18256 4360
rect 18312 5336 18374 5348
rect 18312 4360 18324 5336
rect 18358 4360 18374 5336
rect 18312 4348 18374 4360
rect 18404 5336 18466 5348
rect 18404 4360 18420 5336
rect 18454 4360 18466 5336
rect 18404 4348 18466 4360
rect 18522 5336 18584 5348
rect 18522 4360 18534 5336
rect 18568 4360 18584 5336
rect 18522 4348 18584 4360
rect 18614 5336 18676 5348
rect 18614 4360 18630 5336
rect 18664 4360 18676 5336
rect 18614 4348 18676 4360
rect 10332 4100 10394 4112
rect 10332 3124 10344 4100
rect 10378 3124 10394 4100
rect 10332 3112 10394 3124
rect 10424 4100 10486 4112
rect 10424 3124 10440 4100
rect 10474 3124 10486 4100
rect 10424 3112 10486 3124
rect 10542 4100 10604 4112
rect 10542 3124 10554 4100
rect 10588 3124 10604 4100
rect 10542 3112 10604 3124
rect 10634 4100 10696 4112
rect 10634 3124 10650 4100
rect 10684 3124 10696 4100
rect 10634 3112 10696 3124
rect 10752 4100 10814 4112
rect 10752 3124 10764 4100
rect 10798 3124 10814 4100
rect 10752 3112 10814 3124
rect 10844 4100 10906 4112
rect 10844 3124 10860 4100
rect 10894 3124 10906 4100
rect 10844 3112 10906 3124
rect 10962 4100 11024 4112
rect 10962 3124 10974 4100
rect 11008 3124 11024 4100
rect 10962 3112 11024 3124
rect 11054 4100 11116 4112
rect 11054 3124 11070 4100
rect 11104 3124 11116 4100
rect 11054 3112 11116 3124
rect 11172 4100 11234 4112
rect 11172 3124 11184 4100
rect 11218 3124 11234 4100
rect 11172 3112 11234 3124
rect 11264 4100 11326 4112
rect 11264 3124 11280 4100
rect 11314 3124 11326 4100
rect 11264 3112 11326 3124
rect 11382 4100 11444 4112
rect 11382 3124 11394 4100
rect 11428 3124 11444 4100
rect 11382 3112 11444 3124
rect 11474 4100 11536 4112
rect 11474 3124 11490 4100
rect 11524 3124 11536 4100
rect 11474 3112 11536 3124
rect 11592 4100 11654 4112
rect 11592 3124 11604 4100
rect 11638 3124 11654 4100
rect 11592 3112 11654 3124
rect 11684 4100 11746 4112
rect 11684 3124 11700 4100
rect 11734 3124 11746 4100
rect 11684 3112 11746 3124
rect 11802 4100 11864 4112
rect 11802 3124 11814 4100
rect 11848 3124 11864 4100
rect 11802 3112 11864 3124
rect 11894 4100 11956 4112
rect 11894 3124 11910 4100
rect 11944 3124 11956 4100
rect 11894 3112 11956 3124
rect 12012 4100 12074 4112
rect 12012 3124 12024 4100
rect 12058 3124 12074 4100
rect 12012 3112 12074 3124
rect 12104 4100 12166 4112
rect 12104 3124 12120 4100
rect 12154 3124 12166 4100
rect 12104 3112 12166 3124
rect 12222 4100 12284 4112
rect 12222 3124 12234 4100
rect 12268 3124 12284 4100
rect 12222 3112 12284 3124
rect 12314 4100 12376 4112
rect 12314 3124 12330 4100
rect 12364 3124 12376 4100
rect 12314 3112 12376 3124
rect 12432 4100 12494 4112
rect 12432 3124 12444 4100
rect 12478 3124 12494 4100
rect 12432 3112 12494 3124
rect 12524 4100 12586 4112
rect 12524 3124 12540 4100
rect 12574 3124 12586 4100
rect 12524 3112 12586 3124
rect 12642 4100 12704 4112
rect 12642 3124 12654 4100
rect 12688 3124 12704 4100
rect 12642 3112 12704 3124
rect 12734 4100 12796 4112
rect 12734 3124 12750 4100
rect 12784 3124 12796 4100
rect 12734 3112 12796 3124
rect 12852 4100 12914 4112
rect 12852 3124 12864 4100
rect 12898 3124 12914 4100
rect 12852 3112 12914 3124
rect 12944 4100 13006 4112
rect 12944 3124 12960 4100
rect 12994 3124 13006 4100
rect 12944 3112 13006 3124
rect 13062 4100 13124 4112
rect 13062 3124 13074 4100
rect 13108 3124 13124 4100
rect 13062 3112 13124 3124
rect 13154 4100 13216 4112
rect 13154 3124 13170 4100
rect 13204 3124 13216 4100
rect 13154 3112 13216 3124
rect 13272 4100 13334 4112
rect 13272 3124 13284 4100
rect 13318 3124 13334 4100
rect 13272 3112 13334 3124
rect 13364 4100 13426 4112
rect 13364 3124 13380 4100
rect 13414 3124 13426 4100
rect 13364 3112 13426 3124
rect 13482 4100 13544 4112
rect 13482 3124 13494 4100
rect 13528 3124 13544 4100
rect 13482 3112 13544 3124
rect 13574 4100 13636 4112
rect 13574 3124 13590 4100
rect 13624 3124 13636 4100
rect 13574 3112 13636 3124
rect 13692 4100 13754 4112
rect 13692 3124 13704 4100
rect 13738 3124 13754 4100
rect 13692 3112 13754 3124
rect 13784 4100 13846 4112
rect 13784 3124 13800 4100
rect 13834 3124 13846 4100
rect 13784 3112 13846 3124
rect 13902 4100 13964 4112
rect 13902 3124 13914 4100
rect 13948 3124 13964 4100
rect 13902 3112 13964 3124
rect 13994 4100 14056 4112
rect 13994 3124 14010 4100
rect 14044 3124 14056 4100
rect 13994 3112 14056 3124
rect 14112 4100 14174 4112
rect 14112 3124 14124 4100
rect 14158 3124 14174 4100
rect 14112 3112 14174 3124
rect 14204 4100 14266 4112
rect 14204 3124 14220 4100
rect 14254 3124 14266 4100
rect 14204 3112 14266 3124
rect 14322 4100 14384 4112
rect 14322 3124 14334 4100
rect 14368 3124 14384 4100
rect 14322 3112 14384 3124
rect 14414 4100 14476 4112
rect 14414 3124 14430 4100
rect 14464 3124 14476 4100
rect 14414 3112 14476 3124
rect 14532 4100 14594 4112
rect 14532 3124 14544 4100
rect 14578 3124 14594 4100
rect 14532 3112 14594 3124
rect 14624 4100 14686 4112
rect 14624 3124 14640 4100
rect 14674 3124 14686 4100
rect 14624 3112 14686 3124
rect 14742 4100 14804 4112
rect 14742 3124 14754 4100
rect 14788 3124 14804 4100
rect 14742 3112 14804 3124
rect 14834 4100 14896 4112
rect 14834 3124 14850 4100
rect 14884 3124 14896 4100
rect 14834 3112 14896 3124
rect 14952 4100 15014 4112
rect 14952 3124 14964 4100
rect 14998 3124 15014 4100
rect 14952 3112 15014 3124
rect 15044 4100 15106 4112
rect 15044 3124 15060 4100
rect 15094 3124 15106 4100
rect 15044 3112 15106 3124
rect 15162 4100 15224 4112
rect 15162 3124 15174 4100
rect 15208 3124 15224 4100
rect 15162 3112 15224 3124
rect 15254 4100 15316 4112
rect 15254 3124 15270 4100
rect 15304 3124 15316 4100
rect 15254 3112 15316 3124
rect 15372 4100 15434 4112
rect 15372 3124 15384 4100
rect 15418 3124 15434 4100
rect 15372 3112 15434 3124
rect 15464 4100 15526 4112
rect 15464 3124 15480 4100
rect 15514 3124 15526 4100
rect 15464 3112 15526 3124
rect 15582 4100 15644 4112
rect 15582 3124 15594 4100
rect 15628 3124 15644 4100
rect 15582 3112 15644 3124
rect 15674 4100 15736 4112
rect 15674 3124 15690 4100
rect 15724 3124 15736 4100
rect 15674 3112 15736 3124
rect 15792 4100 15854 4112
rect 15792 3124 15804 4100
rect 15838 3124 15854 4100
rect 15792 3112 15854 3124
rect 15884 4100 15946 4112
rect 15884 3124 15900 4100
rect 15934 3124 15946 4100
rect 15884 3112 15946 3124
rect 16002 4100 16064 4112
rect 16002 3124 16014 4100
rect 16048 3124 16064 4100
rect 16002 3112 16064 3124
rect 16094 4100 16156 4112
rect 16094 3124 16110 4100
rect 16144 3124 16156 4100
rect 16094 3112 16156 3124
rect 16212 4100 16274 4112
rect 16212 3124 16224 4100
rect 16258 3124 16274 4100
rect 16212 3112 16274 3124
rect 16304 4100 16366 4112
rect 16304 3124 16320 4100
rect 16354 3124 16366 4100
rect 16304 3112 16366 3124
rect 16422 4100 16484 4112
rect 16422 3124 16434 4100
rect 16468 3124 16484 4100
rect 16422 3112 16484 3124
rect 16514 4100 16576 4112
rect 16514 3124 16530 4100
rect 16564 3124 16576 4100
rect 16514 3112 16576 3124
rect 16632 4100 16694 4112
rect 16632 3124 16644 4100
rect 16678 3124 16694 4100
rect 16632 3112 16694 3124
rect 16724 4100 16786 4112
rect 16724 3124 16740 4100
rect 16774 3124 16786 4100
rect 16724 3112 16786 3124
rect 16842 4100 16904 4112
rect 16842 3124 16854 4100
rect 16888 3124 16904 4100
rect 16842 3112 16904 3124
rect 16934 4100 16996 4112
rect 16934 3124 16950 4100
rect 16984 3124 16996 4100
rect 16934 3112 16996 3124
rect 17052 4100 17114 4112
rect 17052 3124 17064 4100
rect 17098 3124 17114 4100
rect 17052 3112 17114 3124
rect 17144 4100 17206 4112
rect 17144 3124 17160 4100
rect 17194 3124 17206 4100
rect 17144 3112 17206 3124
rect 17262 4100 17324 4112
rect 17262 3124 17274 4100
rect 17308 3124 17324 4100
rect 17262 3112 17324 3124
rect 17354 4100 17416 4112
rect 17354 3124 17370 4100
rect 17404 3124 17416 4100
rect 17354 3112 17416 3124
rect 17472 4100 17534 4112
rect 17472 3124 17484 4100
rect 17518 3124 17534 4100
rect 17472 3112 17534 3124
rect 17564 4100 17626 4112
rect 17564 3124 17580 4100
rect 17614 3124 17626 4100
rect 17564 3112 17626 3124
rect 17682 4100 17744 4112
rect 17682 3124 17694 4100
rect 17728 3124 17744 4100
rect 17682 3112 17744 3124
rect 17774 4100 17836 4112
rect 17774 3124 17790 4100
rect 17824 3124 17836 4100
rect 17774 3112 17836 3124
rect 17892 4100 17954 4112
rect 17892 3124 17904 4100
rect 17938 3124 17954 4100
rect 17892 3112 17954 3124
rect 17984 4100 18046 4112
rect 17984 3124 18000 4100
rect 18034 3124 18046 4100
rect 17984 3112 18046 3124
rect 18102 4100 18164 4112
rect 18102 3124 18114 4100
rect 18148 3124 18164 4100
rect 18102 3112 18164 3124
rect 18194 4100 18256 4112
rect 18194 3124 18210 4100
rect 18244 3124 18256 4100
rect 18194 3112 18256 3124
rect 18312 4100 18374 4112
rect 18312 3124 18324 4100
rect 18358 3124 18374 4100
rect 18312 3112 18374 3124
rect 18404 4100 18466 4112
rect 18404 3124 18420 4100
rect 18454 3124 18466 4100
rect 18404 3112 18466 3124
rect 18522 4100 18584 4112
rect 18522 3124 18534 4100
rect 18568 3124 18584 4100
rect 18522 3112 18584 3124
rect 18614 4100 18676 4112
rect 18614 3124 18630 4100
rect 18664 3124 18676 4100
rect 18614 3112 18676 3124
rect 2570 -1598 2632 -1586
rect 2570 -2574 2582 -1598
rect 2616 -2574 2632 -1598
rect 2570 -2586 2632 -2574
rect 2662 -1598 2728 -1586
rect 2662 -2574 2678 -1598
rect 2712 -2574 2728 -1598
rect 2662 -2586 2728 -2574
rect 2758 -1598 2820 -1586
rect 2758 -2574 2774 -1598
rect 2808 -2574 2820 -1598
rect 3308 -1598 3370 -1586
rect 2758 -2586 2820 -2574
rect 3308 -2574 3320 -1598
rect 3354 -2574 3370 -1598
rect 3308 -2586 3370 -2574
rect 3400 -1598 3462 -1586
rect 3400 -2574 3416 -1598
rect 3450 -2574 3462 -1598
rect 3400 -2586 3462 -2574
rect 3518 -1598 3580 -1586
rect 3518 -2574 3530 -1598
rect 3564 -2574 3580 -1598
rect 3518 -2586 3580 -2574
rect 3610 -1598 3672 -1586
rect 3610 -2574 3626 -1598
rect 3660 -2574 3672 -1598
rect 3610 -2586 3672 -2574
rect 3728 -1598 3790 -1586
rect 3728 -2574 3740 -1598
rect 3774 -2574 3790 -1598
rect 3728 -2586 3790 -2574
rect 3820 -1598 3882 -1586
rect 3820 -2574 3836 -1598
rect 3870 -2574 3882 -1598
rect 3820 -2586 3882 -2574
rect 3938 -1598 4000 -1586
rect 3938 -2574 3950 -1598
rect 3984 -2574 4000 -1598
rect 3938 -2586 4000 -2574
rect 4030 -1598 4092 -1586
rect 4030 -2574 4046 -1598
rect 4080 -2574 4092 -1598
rect 4030 -2586 4092 -2574
rect 4148 -1598 4210 -1586
rect 4148 -2574 4160 -1598
rect 4194 -2574 4210 -1598
rect 4148 -2586 4210 -2574
rect 4240 -1598 4302 -1586
rect 4240 -2574 4256 -1598
rect 4290 -2574 4302 -1598
rect 4240 -2586 4302 -2574
rect 4358 -1598 4420 -1586
rect 4358 -2574 4370 -1598
rect 4404 -2574 4420 -1598
rect 4358 -2586 4420 -2574
rect 4450 -1598 4512 -1586
rect 4450 -2574 4466 -1598
rect 4500 -2574 4512 -1598
rect 4450 -2586 4512 -2574
rect 4568 -1598 4630 -1586
rect 4568 -2574 4580 -1598
rect 4614 -2574 4630 -1598
rect 4568 -2586 4630 -2574
rect 4660 -1598 4722 -1586
rect 4660 -2574 4676 -1598
rect 4710 -2574 4722 -1598
rect 4660 -2586 4722 -2574
rect 4778 -1598 4840 -1586
rect 4778 -2574 4790 -1598
rect 4824 -2574 4840 -1598
rect 4778 -2586 4840 -2574
rect 4870 -1598 4932 -1586
rect 4870 -2574 4886 -1598
rect 4920 -2574 4932 -1598
rect 4870 -2586 4932 -2574
rect 5482 -1598 5544 -1586
rect 5482 -2574 5494 -1598
rect 5528 -2574 5544 -1598
rect 5482 -2586 5544 -2574
rect 5574 -1598 5636 -1586
rect 5574 -2574 5590 -1598
rect 5624 -2574 5636 -1598
rect 5574 -2586 5636 -2574
rect 5692 -1598 5754 -1586
rect 5692 -2574 5704 -1598
rect 5738 -2574 5754 -1598
rect 5692 -2586 5754 -2574
rect 5784 -1598 5846 -1586
rect 5784 -2574 5800 -1598
rect 5834 -2574 5846 -1598
rect 5784 -2586 5846 -2574
rect 5902 -1598 5964 -1586
rect 5902 -2574 5914 -1598
rect 5948 -2574 5964 -1598
rect 5902 -2586 5964 -2574
rect 5994 -1598 6056 -1586
rect 5994 -2574 6010 -1598
rect 6044 -2574 6056 -1598
rect 5994 -2586 6056 -2574
rect 6112 -1598 6174 -1586
rect 6112 -2574 6124 -1598
rect 6158 -2574 6174 -1598
rect 6112 -2586 6174 -2574
rect 6204 -1598 6266 -1586
rect 6204 -2574 6220 -1598
rect 6254 -2574 6266 -1598
rect 6204 -2586 6266 -2574
rect 6322 -1598 6384 -1586
rect 6322 -2574 6334 -1598
rect 6368 -2574 6384 -1598
rect 6322 -2586 6384 -2574
rect 6414 -1598 6476 -1586
rect 6414 -2574 6430 -1598
rect 6464 -2574 6476 -1598
rect 6414 -2586 6476 -2574
rect 6532 -1598 6594 -1586
rect 6532 -2574 6544 -1598
rect 6578 -2574 6594 -1598
rect 6532 -2586 6594 -2574
rect 6624 -1598 6686 -1586
rect 6624 -2574 6640 -1598
rect 6674 -2574 6686 -1598
rect 6624 -2586 6686 -2574
rect 6742 -1598 6804 -1586
rect 6742 -2574 6754 -1598
rect 6788 -2574 6804 -1598
rect 6742 -2586 6804 -2574
rect 6834 -1598 6896 -1586
rect 6834 -2574 6850 -1598
rect 6884 -2574 6896 -1598
rect 6834 -2586 6896 -2574
rect 6952 -1598 7014 -1586
rect 6952 -2574 6964 -1598
rect 6998 -2574 7014 -1598
rect 6952 -2586 7014 -2574
rect 7044 -1598 7106 -1586
rect 7044 -2574 7060 -1598
rect 7094 -2574 7106 -1598
rect 7044 -2586 7106 -2574
rect 7162 -1598 7224 -1586
rect 7162 -2574 7174 -1598
rect 7208 -2574 7224 -1598
rect 7162 -2586 7224 -2574
rect 7254 -1598 7316 -1586
rect 7254 -2574 7270 -1598
rect 7304 -2574 7316 -1598
rect 7254 -2586 7316 -2574
rect 7372 -1598 7434 -1586
rect 7372 -2574 7384 -1598
rect 7418 -2574 7434 -1598
rect 7372 -2586 7434 -2574
rect 7464 -1598 7526 -1586
rect 7464 -2574 7480 -1598
rect 7514 -2574 7526 -1598
rect 7464 -2586 7526 -2574
rect 7582 -1598 7644 -1586
rect 7582 -2574 7594 -1598
rect 7628 -2574 7644 -1598
rect 7582 -2586 7644 -2574
rect 7674 -1598 7736 -1586
rect 7674 -2574 7690 -1598
rect 7724 -2574 7736 -1598
rect 7674 -2586 7736 -2574
rect 7792 -1598 7854 -1586
rect 7792 -2574 7804 -1598
rect 7838 -2574 7854 -1598
rect 7792 -2586 7854 -2574
rect 7884 -1598 7946 -1586
rect 7884 -2574 7900 -1598
rect 7934 -2574 7946 -1598
rect 7884 -2586 7946 -2574
rect 8002 -1598 8064 -1586
rect 8002 -2574 8014 -1598
rect 8048 -2574 8064 -1598
rect 8002 -2586 8064 -2574
rect 8094 -1598 8156 -1586
rect 8094 -2574 8110 -1598
rect 8144 -2574 8156 -1598
rect 8094 -2586 8156 -2574
rect 8212 -1598 8274 -1586
rect 8212 -2574 8224 -1598
rect 8258 -2574 8274 -1598
rect 8212 -2586 8274 -2574
rect 8304 -1598 8366 -1586
rect 8304 -2574 8320 -1598
rect 8354 -2574 8366 -1598
rect 8304 -2586 8366 -2574
rect 8422 -1598 8484 -1586
rect 8422 -2574 8434 -1598
rect 8468 -2574 8484 -1598
rect 8422 -2586 8484 -2574
rect 8514 -1598 8576 -1586
rect 8514 -2574 8530 -1598
rect 8564 -2574 8576 -1598
rect 8514 -2586 8576 -2574
rect 8632 -1598 8694 -1586
rect 8632 -2574 8644 -1598
rect 8678 -2574 8694 -1598
rect 8632 -2586 8694 -2574
rect 8724 -1598 8786 -1586
rect 8724 -2574 8740 -1598
rect 8774 -2574 8786 -1598
rect 8724 -2586 8786 -2574
rect 8842 -1598 8904 -1586
rect 8842 -2574 8854 -1598
rect 8888 -2574 8904 -1598
rect 8842 -2586 8904 -2574
rect 8934 -1598 8996 -1586
rect 8934 -2574 8950 -1598
rect 8984 -2574 8996 -1598
rect 8934 -2586 8996 -2574
rect 9052 -1598 9114 -1586
rect 9052 -2574 9064 -1598
rect 9098 -2574 9114 -1598
rect 9052 -2586 9114 -2574
rect 9144 -1598 9206 -1586
rect 9144 -2574 9160 -1598
rect 9194 -2574 9206 -1598
rect 9144 -2586 9206 -2574
rect 5482 -2834 5544 -2822
rect 5482 -3810 5494 -2834
rect 5528 -3810 5544 -2834
rect 5482 -3822 5544 -3810
rect 5574 -2834 5636 -2822
rect 5574 -3810 5590 -2834
rect 5624 -3810 5636 -2834
rect 5574 -3822 5636 -3810
rect 5692 -2834 5754 -2822
rect 5692 -3810 5704 -2834
rect 5738 -3810 5754 -2834
rect 5692 -3822 5754 -3810
rect 5784 -2834 5846 -2822
rect 5784 -3810 5800 -2834
rect 5834 -3810 5846 -2834
rect 5784 -3822 5846 -3810
rect 5902 -2834 5964 -2822
rect 5902 -3810 5914 -2834
rect 5948 -3810 5964 -2834
rect 5902 -3822 5964 -3810
rect 5994 -2834 6056 -2822
rect 5994 -3810 6010 -2834
rect 6044 -3810 6056 -2834
rect 5994 -3822 6056 -3810
rect 6112 -2834 6174 -2822
rect 6112 -3810 6124 -2834
rect 6158 -3810 6174 -2834
rect 6112 -3822 6174 -3810
rect 6204 -2834 6266 -2822
rect 6204 -3810 6220 -2834
rect 6254 -3810 6266 -2834
rect 6204 -3822 6266 -3810
rect 6322 -2834 6384 -2822
rect 6322 -3810 6334 -2834
rect 6368 -3810 6384 -2834
rect 6322 -3822 6384 -3810
rect 6414 -2834 6476 -2822
rect 6414 -3810 6430 -2834
rect 6464 -3810 6476 -2834
rect 6414 -3822 6476 -3810
rect 6532 -2834 6594 -2822
rect 6532 -3810 6544 -2834
rect 6578 -3810 6594 -2834
rect 6532 -3822 6594 -3810
rect 6624 -2834 6686 -2822
rect 6624 -3810 6640 -2834
rect 6674 -3810 6686 -2834
rect 6624 -3822 6686 -3810
rect 6742 -2834 6804 -2822
rect 6742 -3810 6754 -2834
rect 6788 -3810 6804 -2834
rect 6742 -3822 6804 -3810
rect 6834 -2834 6896 -2822
rect 6834 -3810 6850 -2834
rect 6884 -3810 6896 -2834
rect 6834 -3822 6896 -3810
rect 6952 -2834 7014 -2822
rect 6952 -3810 6964 -2834
rect 6998 -3810 7014 -2834
rect 6952 -3822 7014 -3810
rect 7044 -2834 7106 -2822
rect 7044 -3810 7060 -2834
rect 7094 -3810 7106 -2834
rect 7044 -3822 7106 -3810
rect 7162 -2834 7224 -2822
rect 7162 -3810 7174 -2834
rect 7208 -3810 7224 -2834
rect 7162 -3822 7224 -3810
rect 7254 -2834 7316 -2822
rect 7254 -3810 7270 -2834
rect 7304 -3810 7316 -2834
rect 7254 -3822 7316 -3810
rect 7372 -2834 7434 -2822
rect 7372 -3810 7384 -2834
rect 7418 -3810 7434 -2834
rect 7372 -3822 7434 -3810
rect 7464 -2834 7526 -2822
rect 7464 -3810 7480 -2834
rect 7514 -3810 7526 -2834
rect 7464 -3822 7526 -3810
rect 7582 -2834 7644 -2822
rect 7582 -3810 7594 -2834
rect 7628 -3810 7644 -2834
rect 7582 -3822 7644 -3810
rect 7674 -2834 7736 -2822
rect 7674 -3810 7690 -2834
rect 7724 -3810 7736 -2834
rect 7674 -3822 7736 -3810
rect 7792 -2834 7854 -2822
rect 7792 -3810 7804 -2834
rect 7838 -3810 7854 -2834
rect 7792 -3822 7854 -3810
rect 7884 -2834 7946 -2822
rect 7884 -3810 7900 -2834
rect 7934 -3810 7946 -2834
rect 7884 -3822 7946 -3810
rect 8002 -2834 8064 -2822
rect 8002 -3810 8014 -2834
rect 8048 -3810 8064 -2834
rect 8002 -3822 8064 -3810
rect 8094 -2834 8156 -2822
rect 8094 -3810 8110 -2834
rect 8144 -3810 8156 -2834
rect 8094 -3822 8156 -3810
rect 8212 -2834 8274 -2822
rect 8212 -3810 8224 -2834
rect 8258 -3810 8274 -2834
rect 8212 -3822 8274 -3810
rect 8304 -2834 8366 -2822
rect 8304 -3810 8320 -2834
rect 8354 -3810 8366 -2834
rect 8304 -3822 8366 -3810
rect 8422 -2834 8484 -2822
rect 8422 -3810 8434 -2834
rect 8468 -3810 8484 -2834
rect 8422 -3822 8484 -3810
rect 8514 -2834 8576 -2822
rect 8514 -3810 8530 -2834
rect 8564 -3810 8576 -2834
rect 8514 -3822 8576 -3810
rect 8632 -2834 8694 -2822
rect 8632 -3810 8644 -2834
rect 8678 -3810 8694 -2834
rect 8632 -3822 8694 -3810
rect 8724 -2834 8786 -2822
rect 8724 -3810 8740 -2834
rect 8774 -3810 8786 -2834
rect 8724 -3822 8786 -3810
rect 8842 -2834 8904 -2822
rect 8842 -3810 8854 -2834
rect 8888 -3810 8904 -2834
rect 8842 -3822 8904 -3810
rect 8934 -2834 8996 -2822
rect 8934 -3810 8950 -2834
rect 8984 -3810 8996 -2834
rect 8934 -3822 8996 -3810
rect 9052 -2834 9114 -2822
rect 9052 -3810 9064 -2834
rect 9098 -3810 9114 -2834
rect 9052 -3822 9114 -3810
rect 9144 -2834 9206 -2822
rect 9144 -3810 9160 -2834
rect 9194 -3810 9206 -2834
rect 9144 -3822 9206 -3810
<< ndiffc >>
rect 10344 12060 10378 13036
rect 10440 12060 10474 13036
rect 10554 12060 10588 13036
rect 10650 12060 10684 13036
rect 10764 12060 10798 13036
rect 10860 12060 10894 13036
rect 10974 12060 11008 13036
rect 11070 12060 11104 13036
rect 11184 12060 11218 13036
rect 11280 12060 11314 13036
rect 11394 12060 11428 13036
rect 11490 12060 11524 13036
rect 11604 12060 11638 13036
rect 11700 12060 11734 13036
rect 11814 12060 11848 13036
rect 11910 12060 11944 13036
rect 12024 12060 12058 13036
rect 12120 12060 12154 13036
rect 12234 12060 12268 13036
rect 12330 12060 12364 13036
rect 12444 12060 12478 13036
rect 12540 12060 12574 13036
rect 12654 12060 12688 13036
rect 12750 12060 12784 13036
rect 12864 12060 12898 13036
rect 12960 12060 12994 13036
rect 13074 12060 13108 13036
rect 13170 12060 13204 13036
rect 13284 12060 13318 13036
rect 13380 12060 13414 13036
rect 13494 12060 13528 13036
rect 13590 12060 13624 13036
rect 13704 12060 13738 13036
rect 13800 12060 13834 13036
rect 13914 12060 13948 13036
rect 14010 12060 14044 13036
rect 14124 12060 14158 13036
rect 14220 12060 14254 13036
rect 14334 12060 14368 13036
rect 14430 12060 14464 13036
rect 14544 12060 14578 13036
rect 14640 12060 14674 13036
rect 14754 12060 14788 13036
rect 14850 12060 14884 13036
rect 14964 12060 14998 13036
rect 15060 12060 15094 13036
rect 15174 12060 15208 13036
rect 15270 12060 15304 13036
rect 15384 12060 15418 13036
rect 15480 12060 15514 13036
rect 15594 12060 15628 13036
rect 15690 12060 15724 13036
rect 15804 12060 15838 13036
rect 15900 12060 15934 13036
rect 16014 12060 16048 13036
rect 16110 12060 16144 13036
rect 16224 12060 16258 13036
rect 16320 12060 16354 13036
rect 16434 12060 16468 13036
rect 16530 12060 16564 13036
rect 16644 12060 16678 13036
rect 16740 12060 16774 13036
rect 16854 12060 16888 13036
rect 16950 12060 16984 13036
rect 17064 12060 17098 13036
rect 17160 12060 17194 13036
rect 17274 12060 17308 13036
rect 17370 12060 17404 13036
rect 17484 12060 17518 13036
rect 17580 12060 17614 13036
rect 17694 12060 17728 13036
rect 17790 12060 17824 13036
rect 17904 12060 17938 13036
rect 18000 12060 18034 13036
rect 18114 12060 18148 13036
rect 18210 12060 18244 13036
rect 18324 12060 18358 13036
rect 18420 12060 18454 13036
rect 18534 12060 18568 13036
rect 18630 12060 18664 13036
rect 10344 10842 10378 11818
rect 10440 10842 10474 11818
rect 10554 10842 10588 11818
rect 10650 10842 10684 11818
rect 10764 10842 10798 11818
rect 10860 10842 10894 11818
rect 10974 10842 11008 11818
rect 11070 10842 11104 11818
rect 11184 10842 11218 11818
rect 11280 10842 11314 11818
rect 11394 10842 11428 11818
rect 11490 10842 11524 11818
rect 11604 10842 11638 11818
rect 11700 10842 11734 11818
rect 11814 10842 11848 11818
rect 11910 10842 11944 11818
rect 12024 10842 12058 11818
rect 12120 10842 12154 11818
rect 12234 10842 12268 11818
rect 12330 10842 12364 11818
rect 12444 10842 12478 11818
rect 12540 10842 12574 11818
rect 12654 10842 12688 11818
rect 12750 10842 12784 11818
rect 12864 10842 12898 11818
rect 12960 10842 12994 11818
rect 13074 10842 13108 11818
rect 13170 10842 13204 11818
rect 13284 10842 13318 11818
rect 13380 10842 13414 11818
rect 13494 10842 13528 11818
rect 13590 10842 13624 11818
rect 13704 10842 13738 11818
rect 13800 10842 13834 11818
rect 13914 10842 13948 11818
rect 14010 10842 14044 11818
rect 14124 10842 14158 11818
rect 14220 10842 14254 11818
rect 14334 10842 14368 11818
rect 14430 10842 14464 11818
rect 14544 10842 14578 11818
rect 14640 10842 14674 11818
rect 14754 10842 14788 11818
rect 14850 10842 14884 11818
rect 14964 10842 14998 11818
rect 15060 10842 15094 11818
rect 15174 10842 15208 11818
rect 15270 10842 15304 11818
rect 15384 10842 15418 11818
rect 15480 10842 15514 11818
rect 15594 10842 15628 11818
rect 15690 10842 15724 11818
rect 15804 10842 15838 11818
rect 15900 10842 15934 11818
rect 16014 10842 16048 11818
rect 16110 10842 16144 11818
rect 16224 10842 16258 11818
rect 16320 10842 16354 11818
rect 16434 10842 16468 11818
rect 16530 10842 16564 11818
rect 16644 10842 16678 11818
rect 16740 10842 16774 11818
rect 16854 10842 16888 11818
rect 16950 10842 16984 11818
rect 17064 10842 17098 11818
rect 17160 10842 17194 11818
rect 17274 10842 17308 11818
rect 17370 10842 17404 11818
rect 17484 10842 17518 11818
rect 17580 10842 17614 11818
rect 17694 10842 17728 11818
rect 17790 10842 17824 11818
rect 17904 10842 17938 11818
rect 18000 10842 18034 11818
rect 18114 10842 18148 11818
rect 18210 10842 18244 11818
rect 18324 10842 18358 11818
rect 18420 10842 18454 11818
rect 18534 10842 18568 11818
rect 18630 10842 18664 11818
rect 5494 5976 5528 6952
rect 5590 5976 5624 6952
rect 5704 5976 5738 6952
rect 5800 5976 5834 6952
rect 5914 5976 5948 6952
rect 6010 5976 6044 6952
rect 6124 5976 6158 6952
rect 6220 5976 6254 6952
rect 6334 5976 6368 6952
rect 6430 5976 6464 6952
rect 6544 5976 6578 6952
rect 6640 5976 6674 6952
rect 6754 5976 6788 6952
rect 6850 5976 6884 6952
rect 6964 5976 6998 6952
rect 7060 5976 7094 6952
rect 7174 5976 7208 6952
rect 7270 5976 7304 6952
rect 7384 5976 7418 6952
rect 7480 5976 7514 6952
rect 7594 5976 7628 6952
rect 7690 5976 7724 6952
rect 7804 5976 7838 6952
rect 7900 5976 7934 6952
rect 8014 5976 8048 6952
rect 8110 5976 8144 6952
rect 8224 5976 8258 6952
rect 8320 5976 8354 6952
rect 8434 5976 8468 6952
rect 8530 5976 8564 6952
rect 8644 5976 8678 6952
rect 8740 5976 8774 6952
rect 8854 5976 8888 6952
rect 8950 5976 8984 6952
rect 9064 5976 9098 6952
rect 9160 5976 9194 6952
rect 2586 4352 2620 5328
rect 2674 4352 2708 5328
rect 3530 4352 3564 5328
rect 3626 4352 3660 5328
rect 3740 4352 3774 5328
rect 3836 4352 3870 5328
rect 3950 4352 3984 5328
rect 4046 4352 4080 5328
rect 4160 4352 4194 5328
rect 4256 4352 4290 5328
rect 2586 -3802 2620 -2826
rect 2674 -3802 2708 -2826
rect 3530 -3802 3564 -2826
rect 3626 -3802 3660 -2826
rect 3740 -3802 3774 -2826
rect 3836 -3802 3870 -2826
rect 3950 -3802 3984 -2826
rect 4046 -3802 4080 -2826
rect 4160 -3802 4194 -2826
rect 4256 -3802 4290 -2826
rect 5494 -6826 5528 -5850
rect 5590 -6826 5624 -5850
rect 5704 -6826 5738 -5850
rect 5800 -6826 5834 -5850
rect 5914 -6826 5948 -5850
rect 6010 -6826 6044 -5850
rect 6124 -6826 6158 -5850
rect 6220 -6826 6254 -5850
rect 6334 -6826 6368 -5850
rect 6430 -6826 6464 -5850
rect 6544 -6826 6578 -5850
rect 6640 -6826 6674 -5850
rect 6754 -6826 6788 -5850
rect 6850 -6826 6884 -5850
rect 6964 -6826 6998 -5850
rect 7060 -6826 7094 -5850
rect 7174 -6826 7208 -5850
rect 7270 -6826 7304 -5850
rect 7384 -6826 7418 -5850
rect 7480 -6826 7514 -5850
rect 7594 -6826 7628 -5850
rect 7690 -6826 7724 -5850
rect 7804 -6826 7838 -5850
rect 7900 -6826 7934 -5850
rect 8014 -6826 8048 -5850
rect 8110 -6826 8144 -5850
rect 8224 -6826 8258 -5850
rect 8320 -6826 8354 -5850
rect 8434 -6826 8468 -5850
rect 8530 -6826 8564 -5850
rect 8644 -6826 8678 -5850
rect 8740 -6826 8774 -5850
rect 8854 -6826 8888 -5850
rect 8950 -6826 8984 -5850
rect 9064 -6826 9098 -5850
rect 9160 -6826 9194 -5850
<< pdiffc >>
rect 2582 3124 2616 4100
rect 2678 3124 2712 4100
rect 2774 3124 2808 4100
rect 3320 3124 3354 4100
rect 3416 3124 3450 4100
rect 3530 3124 3564 4100
rect 3626 3124 3660 4100
rect 3740 3124 3774 4100
rect 3836 3124 3870 4100
rect 3950 3124 3984 4100
rect 4046 3124 4080 4100
rect 4160 3124 4194 4100
rect 4256 3124 4290 4100
rect 4370 3124 4404 4100
rect 4466 3124 4500 4100
rect 4580 3124 4614 4100
rect 4676 3124 4710 4100
rect 4790 3124 4824 4100
rect 4886 3124 4920 4100
rect 5494 4360 5528 5336
rect 5590 4360 5624 5336
rect 5704 4360 5738 5336
rect 5800 4360 5834 5336
rect 5914 4360 5948 5336
rect 6010 4360 6044 5336
rect 6124 4360 6158 5336
rect 6220 4360 6254 5336
rect 6334 4360 6368 5336
rect 6430 4360 6464 5336
rect 6544 4360 6578 5336
rect 6640 4360 6674 5336
rect 6754 4360 6788 5336
rect 6850 4360 6884 5336
rect 6964 4360 6998 5336
rect 7060 4360 7094 5336
rect 7174 4360 7208 5336
rect 7270 4360 7304 5336
rect 7384 4360 7418 5336
rect 7480 4360 7514 5336
rect 7594 4360 7628 5336
rect 7690 4360 7724 5336
rect 7804 4360 7838 5336
rect 7900 4360 7934 5336
rect 8014 4360 8048 5336
rect 8110 4360 8144 5336
rect 8224 4360 8258 5336
rect 8320 4360 8354 5336
rect 8434 4360 8468 5336
rect 8530 4360 8564 5336
rect 8644 4360 8678 5336
rect 8740 4360 8774 5336
rect 8854 4360 8888 5336
rect 8950 4360 8984 5336
rect 9064 4360 9098 5336
rect 9160 4360 9194 5336
rect 5494 3124 5528 4100
rect 5590 3124 5624 4100
rect 5704 3124 5738 4100
rect 5800 3124 5834 4100
rect 5914 3124 5948 4100
rect 6010 3124 6044 4100
rect 6124 3124 6158 4100
rect 6220 3124 6254 4100
rect 6334 3124 6368 4100
rect 6430 3124 6464 4100
rect 6544 3124 6578 4100
rect 6640 3124 6674 4100
rect 6754 3124 6788 4100
rect 6850 3124 6884 4100
rect 6964 3124 6998 4100
rect 7060 3124 7094 4100
rect 7174 3124 7208 4100
rect 7270 3124 7304 4100
rect 7384 3124 7418 4100
rect 7480 3124 7514 4100
rect 7594 3124 7628 4100
rect 7690 3124 7724 4100
rect 7804 3124 7838 4100
rect 7900 3124 7934 4100
rect 8014 3124 8048 4100
rect 8110 3124 8144 4100
rect 8224 3124 8258 4100
rect 8320 3124 8354 4100
rect 8434 3124 8468 4100
rect 8530 3124 8564 4100
rect 8644 3124 8678 4100
rect 8740 3124 8774 4100
rect 8854 3124 8888 4100
rect 8950 3124 8984 4100
rect 9064 3124 9098 4100
rect 9160 3124 9194 4100
rect 10344 6832 10378 7808
rect 10440 6832 10474 7808
rect 10554 6832 10588 7808
rect 10650 6832 10684 7808
rect 10764 6832 10798 7808
rect 10860 6832 10894 7808
rect 10974 6832 11008 7808
rect 11070 6832 11104 7808
rect 11184 6832 11218 7808
rect 11280 6832 11314 7808
rect 11394 6832 11428 7808
rect 11490 6832 11524 7808
rect 11604 6832 11638 7808
rect 11700 6832 11734 7808
rect 11814 6832 11848 7808
rect 11910 6832 11944 7808
rect 12024 6832 12058 7808
rect 12120 6832 12154 7808
rect 12234 6832 12268 7808
rect 12330 6832 12364 7808
rect 12444 6832 12478 7808
rect 12540 6832 12574 7808
rect 12654 6832 12688 7808
rect 12750 6832 12784 7808
rect 12864 6832 12898 7808
rect 12960 6832 12994 7808
rect 13074 6832 13108 7808
rect 13170 6832 13204 7808
rect 13284 6832 13318 7808
rect 13380 6832 13414 7808
rect 13494 6832 13528 7808
rect 13590 6832 13624 7808
rect 13704 6832 13738 7808
rect 13800 6832 13834 7808
rect 13914 6832 13948 7808
rect 14010 6832 14044 7808
rect 14124 6832 14158 7808
rect 14220 6832 14254 7808
rect 14334 6832 14368 7808
rect 14430 6832 14464 7808
rect 14544 6832 14578 7808
rect 14640 6832 14674 7808
rect 14754 6832 14788 7808
rect 14850 6832 14884 7808
rect 14964 6832 14998 7808
rect 15060 6832 15094 7808
rect 15174 6832 15208 7808
rect 15270 6832 15304 7808
rect 15384 6832 15418 7808
rect 15480 6832 15514 7808
rect 15594 6832 15628 7808
rect 15690 6832 15724 7808
rect 15804 6832 15838 7808
rect 15900 6832 15934 7808
rect 16014 6832 16048 7808
rect 16110 6832 16144 7808
rect 16224 6832 16258 7808
rect 16320 6832 16354 7808
rect 16434 6832 16468 7808
rect 16530 6832 16564 7808
rect 16644 6832 16678 7808
rect 16740 6832 16774 7808
rect 16854 6832 16888 7808
rect 16950 6832 16984 7808
rect 17064 6832 17098 7808
rect 17160 6832 17194 7808
rect 17274 6832 17308 7808
rect 17370 6832 17404 7808
rect 17484 6832 17518 7808
rect 17580 6832 17614 7808
rect 17694 6832 17728 7808
rect 17790 6832 17824 7808
rect 17904 6832 17938 7808
rect 18000 6832 18034 7808
rect 18114 6832 18148 7808
rect 18210 6832 18244 7808
rect 18324 6832 18358 7808
rect 18420 6832 18454 7808
rect 18534 6832 18568 7808
rect 18630 6832 18664 7808
rect 10344 5596 10378 6572
rect 10440 5596 10474 6572
rect 10554 5596 10588 6572
rect 10650 5596 10684 6572
rect 10764 5596 10798 6572
rect 10860 5596 10894 6572
rect 10974 5596 11008 6572
rect 11070 5596 11104 6572
rect 11184 5596 11218 6572
rect 11280 5596 11314 6572
rect 11394 5596 11428 6572
rect 11490 5596 11524 6572
rect 11604 5596 11638 6572
rect 11700 5596 11734 6572
rect 11814 5596 11848 6572
rect 11910 5596 11944 6572
rect 12024 5596 12058 6572
rect 12120 5596 12154 6572
rect 12234 5596 12268 6572
rect 12330 5596 12364 6572
rect 12444 5596 12478 6572
rect 12540 5596 12574 6572
rect 12654 5596 12688 6572
rect 12750 5596 12784 6572
rect 12864 5596 12898 6572
rect 12960 5596 12994 6572
rect 13074 5596 13108 6572
rect 13170 5596 13204 6572
rect 13284 5596 13318 6572
rect 13380 5596 13414 6572
rect 13494 5596 13528 6572
rect 13590 5596 13624 6572
rect 13704 5596 13738 6572
rect 13800 5596 13834 6572
rect 13914 5596 13948 6572
rect 14010 5596 14044 6572
rect 14124 5596 14158 6572
rect 14220 5596 14254 6572
rect 14334 5596 14368 6572
rect 14430 5596 14464 6572
rect 14544 5596 14578 6572
rect 14640 5596 14674 6572
rect 14754 5596 14788 6572
rect 14850 5596 14884 6572
rect 14964 5596 14998 6572
rect 15060 5596 15094 6572
rect 15174 5596 15208 6572
rect 15270 5596 15304 6572
rect 15384 5596 15418 6572
rect 15480 5596 15514 6572
rect 15594 5596 15628 6572
rect 15690 5596 15724 6572
rect 15804 5596 15838 6572
rect 15900 5596 15934 6572
rect 16014 5596 16048 6572
rect 16110 5596 16144 6572
rect 16224 5596 16258 6572
rect 16320 5596 16354 6572
rect 16434 5596 16468 6572
rect 16530 5596 16564 6572
rect 16644 5596 16678 6572
rect 16740 5596 16774 6572
rect 16854 5596 16888 6572
rect 16950 5596 16984 6572
rect 17064 5596 17098 6572
rect 17160 5596 17194 6572
rect 17274 5596 17308 6572
rect 17370 5596 17404 6572
rect 17484 5596 17518 6572
rect 17580 5596 17614 6572
rect 17694 5596 17728 6572
rect 17790 5596 17824 6572
rect 17904 5596 17938 6572
rect 18000 5596 18034 6572
rect 18114 5596 18148 6572
rect 18210 5596 18244 6572
rect 18324 5596 18358 6572
rect 18420 5596 18454 6572
rect 18534 5596 18568 6572
rect 18630 5596 18664 6572
rect 10344 4360 10378 5336
rect 10440 4360 10474 5336
rect 10554 4360 10588 5336
rect 10650 4360 10684 5336
rect 10764 4360 10798 5336
rect 10860 4360 10894 5336
rect 10974 4360 11008 5336
rect 11070 4360 11104 5336
rect 11184 4360 11218 5336
rect 11280 4360 11314 5336
rect 11394 4360 11428 5336
rect 11490 4360 11524 5336
rect 11604 4360 11638 5336
rect 11700 4360 11734 5336
rect 11814 4360 11848 5336
rect 11910 4360 11944 5336
rect 12024 4360 12058 5336
rect 12120 4360 12154 5336
rect 12234 4360 12268 5336
rect 12330 4360 12364 5336
rect 12444 4360 12478 5336
rect 12540 4360 12574 5336
rect 12654 4360 12688 5336
rect 12750 4360 12784 5336
rect 12864 4360 12898 5336
rect 12960 4360 12994 5336
rect 13074 4360 13108 5336
rect 13170 4360 13204 5336
rect 13284 4360 13318 5336
rect 13380 4360 13414 5336
rect 13494 4360 13528 5336
rect 13590 4360 13624 5336
rect 13704 4360 13738 5336
rect 13800 4360 13834 5336
rect 13914 4360 13948 5336
rect 14010 4360 14044 5336
rect 14124 4360 14158 5336
rect 14220 4360 14254 5336
rect 14334 4360 14368 5336
rect 14430 4360 14464 5336
rect 14544 4360 14578 5336
rect 14640 4360 14674 5336
rect 14754 4360 14788 5336
rect 14850 4360 14884 5336
rect 14964 4360 14998 5336
rect 15060 4360 15094 5336
rect 15174 4360 15208 5336
rect 15270 4360 15304 5336
rect 15384 4360 15418 5336
rect 15480 4360 15514 5336
rect 15594 4360 15628 5336
rect 15690 4360 15724 5336
rect 15804 4360 15838 5336
rect 15900 4360 15934 5336
rect 16014 4360 16048 5336
rect 16110 4360 16144 5336
rect 16224 4360 16258 5336
rect 16320 4360 16354 5336
rect 16434 4360 16468 5336
rect 16530 4360 16564 5336
rect 16644 4360 16678 5336
rect 16740 4360 16774 5336
rect 16854 4360 16888 5336
rect 16950 4360 16984 5336
rect 17064 4360 17098 5336
rect 17160 4360 17194 5336
rect 17274 4360 17308 5336
rect 17370 4360 17404 5336
rect 17484 4360 17518 5336
rect 17580 4360 17614 5336
rect 17694 4360 17728 5336
rect 17790 4360 17824 5336
rect 17904 4360 17938 5336
rect 18000 4360 18034 5336
rect 18114 4360 18148 5336
rect 18210 4360 18244 5336
rect 18324 4360 18358 5336
rect 18420 4360 18454 5336
rect 18534 4360 18568 5336
rect 18630 4360 18664 5336
rect 10344 3124 10378 4100
rect 10440 3124 10474 4100
rect 10554 3124 10588 4100
rect 10650 3124 10684 4100
rect 10764 3124 10798 4100
rect 10860 3124 10894 4100
rect 10974 3124 11008 4100
rect 11070 3124 11104 4100
rect 11184 3124 11218 4100
rect 11280 3124 11314 4100
rect 11394 3124 11428 4100
rect 11490 3124 11524 4100
rect 11604 3124 11638 4100
rect 11700 3124 11734 4100
rect 11814 3124 11848 4100
rect 11910 3124 11944 4100
rect 12024 3124 12058 4100
rect 12120 3124 12154 4100
rect 12234 3124 12268 4100
rect 12330 3124 12364 4100
rect 12444 3124 12478 4100
rect 12540 3124 12574 4100
rect 12654 3124 12688 4100
rect 12750 3124 12784 4100
rect 12864 3124 12898 4100
rect 12960 3124 12994 4100
rect 13074 3124 13108 4100
rect 13170 3124 13204 4100
rect 13284 3124 13318 4100
rect 13380 3124 13414 4100
rect 13494 3124 13528 4100
rect 13590 3124 13624 4100
rect 13704 3124 13738 4100
rect 13800 3124 13834 4100
rect 13914 3124 13948 4100
rect 14010 3124 14044 4100
rect 14124 3124 14158 4100
rect 14220 3124 14254 4100
rect 14334 3124 14368 4100
rect 14430 3124 14464 4100
rect 14544 3124 14578 4100
rect 14640 3124 14674 4100
rect 14754 3124 14788 4100
rect 14850 3124 14884 4100
rect 14964 3124 14998 4100
rect 15060 3124 15094 4100
rect 15174 3124 15208 4100
rect 15270 3124 15304 4100
rect 15384 3124 15418 4100
rect 15480 3124 15514 4100
rect 15594 3124 15628 4100
rect 15690 3124 15724 4100
rect 15804 3124 15838 4100
rect 15900 3124 15934 4100
rect 16014 3124 16048 4100
rect 16110 3124 16144 4100
rect 16224 3124 16258 4100
rect 16320 3124 16354 4100
rect 16434 3124 16468 4100
rect 16530 3124 16564 4100
rect 16644 3124 16678 4100
rect 16740 3124 16774 4100
rect 16854 3124 16888 4100
rect 16950 3124 16984 4100
rect 17064 3124 17098 4100
rect 17160 3124 17194 4100
rect 17274 3124 17308 4100
rect 17370 3124 17404 4100
rect 17484 3124 17518 4100
rect 17580 3124 17614 4100
rect 17694 3124 17728 4100
rect 17790 3124 17824 4100
rect 17904 3124 17938 4100
rect 18000 3124 18034 4100
rect 18114 3124 18148 4100
rect 18210 3124 18244 4100
rect 18324 3124 18358 4100
rect 18420 3124 18454 4100
rect 18534 3124 18568 4100
rect 18630 3124 18664 4100
rect 2582 -2574 2616 -1598
rect 2678 -2574 2712 -1598
rect 2774 -2574 2808 -1598
rect 3320 -2574 3354 -1598
rect 3416 -2574 3450 -1598
rect 3530 -2574 3564 -1598
rect 3626 -2574 3660 -1598
rect 3740 -2574 3774 -1598
rect 3836 -2574 3870 -1598
rect 3950 -2574 3984 -1598
rect 4046 -2574 4080 -1598
rect 4160 -2574 4194 -1598
rect 4256 -2574 4290 -1598
rect 4370 -2574 4404 -1598
rect 4466 -2574 4500 -1598
rect 4580 -2574 4614 -1598
rect 4676 -2574 4710 -1598
rect 4790 -2574 4824 -1598
rect 4886 -2574 4920 -1598
rect 5494 -2574 5528 -1598
rect 5590 -2574 5624 -1598
rect 5704 -2574 5738 -1598
rect 5800 -2574 5834 -1598
rect 5914 -2574 5948 -1598
rect 6010 -2574 6044 -1598
rect 6124 -2574 6158 -1598
rect 6220 -2574 6254 -1598
rect 6334 -2574 6368 -1598
rect 6430 -2574 6464 -1598
rect 6544 -2574 6578 -1598
rect 6640 -2574 6674 -1598
rect 6754 -2574 6788 -1598
rect 6850 -2574 6884 -1598
rect 6964 -2574 6998 -1598
rect 7060 -2574 7094 -1598
rect 7174 -2574 7208 -1598
rect 7270 -2574 7304 -1598
rect 7384 -2574 7418 -1598
rect 7480 -2574 7514 -1598
rect 7594 -2574 7628 -1598
rect 7690 -2574 7724 -1598
rect 7804 -2574 7838 -1598
rect 7900 -2574 7934 -1598
rect 8014 -2574 8048 -1598
rect 8110 -2574 8144 -1598
rect 8224 -2574 8258 -1598
rect 8320 -2574 8354 -1598
rect 8434 -2574 8468 -1598
rect 8530 -2574 8564 -1598
rect 8644 -2574 8678 -1598
rect 8740 -2574 8774 -1598
rect 8854 -2574 8888 -1598
rect 8950 -2574 8984 -1598
rect 9064 -2574 9098 -1598
rect 9160 -2574 9194 -1598
rect 5494 -3810 5528 -2834
rect 5590 -3810 5624 -2834
rect 5704 -3810 5738 -2834
rect 5800 -3810 5834 -2834
rect 5914 -3810 5948 -2834
rect 6010 -3810 6044 -2834
rect 6124 -3810 6158 -2834
rect 6220 -3810 6254 -2834
rect 6334 -3810 6368 -2834
rect 6430 -3810 6464 -2834
rect 6544 -3810 6578 -2834
rect 6640 -3810 6674 -2834
rect 6754 -3810 6788 -2834
rect 6850 -3810 6884 -2834
rect 6964 -3810 6998 -2834
rect 7060 -3810 7094 -2834
rect 7174 -3810 7208 -2834
rect 7270 -3810 7304 -2834
rect 7384 -3810 7418 -2834
rect 7480 -3810 7514 -2834
rect 7594 -3810 7628 -2834
rect 7690 -3810 7724 -2834
rect 7804 -3810 7838 -2834
rect 7900 -3810 7934 -2834
rect 8014 -3810 8048 -2834
rect 8110 -3810 8144 -2834
rect 8224 -3810 8258 -2834
rect 8320 -3810 8354 -2834
rect 8434 -3810 8468 -2834
rect 8530 -3810 8564 -2834
rect 8644 -3810 8678 -2834
rect 8740 -3810 8774 -2834
rect 8854 -3810 8888 -2834
rect 8950 -3810 8984 -2834
rect 9064 -3810 9098 -2834
rect 9160 -3810 9194 -2834
<< psubdiffcont >>
rect 10248 13268 18672 13302
rect 10104 10774 10138 13146
rect 18824 10762 18858 13174
rect 10260 10592 18630 10626
rect 5480 7096 9204 7130
rect 5348 5960 5382 6980
rect 9276 5962 9310 7004
rect 5440 5808 9160 5842
rect 3000 4526 3206 5218
rect 3000 -3692 3206 -3000
rect 5440 -5716 9160 -5682
rect 5348 -6854 5382 -5834
rect 9276 -6878 9310 -5836
rect 5480 -7004 9204 -6970
<< nsubdiffcont >>
rect 10358 7996 18680 8030
rect 5514 5536 9216 5570
rect 2924 3324 3130 4016
rect 5384 3026 5418 5494
rect 9298 3064 9332 5352
rect 10132 3046 10166 7844
rect 18762 3108 18796 7826
rect 5486 2904 9258 2938
rect 10322 2888 18644 2922
rect 5486 -1412 9258 -1378
rect 2924 -2490 3130 -1798
rect 5384 -3968 5418 -1500
rect 9298 -3826 9332 -1538
rect 5514 -4044 9216 -4010
<< poly >>
rect 10376 13120 10492 13136
rect 10376 13086 10392 13120
rect 10476 13086 10492 13120
rect 10376 13070 10492 13086
rect 10796 13120 10912 13136
rect 10796 13086 10812 13120
rect 10896 13086 10912 13120
rect 10394 13048 10424 13070
rect 10604 13048 10634 13074
rect 10796 13070 10912 13086
rect 11216 13120 11332 13136
rect 11216 13086 11232 13120
rect 11316 13086 11332 13120
rect 10814 13048 10844 13070
rect 11024 13048 11054 13074
rect 11216 13070 11332 13086
rect 11636 13120 11752 13136
rect 11636 13086 11652 13120
rect 11736 13086 11752 13120
rect 11234 13048 11264 13070
rect 11444 13048 11474 13074
rect 11636 13070 11752 13086
rect 12056 13120 12172 13136
rect 12056 13086 12072 13120
rect 12156 13086 12172 13120
rect 11654 13048 11684 13070
rect 11864 13048 11894 13074
rect 12056 13070 12172 13086
rect 12476 13120 12592 13136
rect 12476 13086 12492 13120
rect 12576 13086 12592 13120
rect 12074 13048 12104 13070
rect 12284 13048 12314 13074
rect 12476 13070 12592 13086
rect 12896 13120 13012 13136
rect 12896 13086 12912 13120
rect 12996 13086 13012 13120
rect 12494 13048 12524 13070
rect 12704 13048 12734 13074
rect 12896 13070 13012 13086
rect 13316 13120 13432 13136
rect 13316 13086 13332 13120
rect 13416 13086 13432 13120
rect 12914 13048 12944 13070
rect 13124 13048 13154 13074
rect 13316 13070 13432 13086
rect 13736 13120 13852 13136
rect 13736 13086 13752 13120
rect 13836 13086 13852 13120
rect 13334 13048 13364 13070
rect 13544 13048 13574 13074
rect 13736 13070 13852 13086
rect 14156 13120 14272 13136
rect 14156 13086 14172 13120
rect 14256 13086 14272 13120
rect 13754 13048 13784 13070
rect 13964 13048 13994 13074
rect 14156 13070 14272 13086
rect 14576 13120 14692 13136
rect 14576 13086 14592 13120
rect 14676 13086 14692 13120
rect 14174 13048 14204 13070
rect 14384 13048 14414 13074
rect 14576 13070 14692 13086
rect 14996 13120 15112 13136
rect 14996 13086 15012 13120
rect 15096 13086 15112 13120
rect 14594 13048 14624 13070
rect 14804 13048 14834 13074
rect 14996 13070 15112 13086
rect 15416 13120 15532 13136
rect 15416 13086 15432 13120
rect 15516 13086 15532 13120
rect 15014 13048 15044 13070
rect 15224 13048 15254 13074
rect 15416 13070 15532 13086
rect 15836 13120 15952 13136
rect 15836 13086 15852 13120
rect 15936 13086 15952 13120
rect 15434 13048 15464 13070
rect 15644 13048 15674 13074
rect 15836 13070 15952 13086
rect 16256 13120 16372 13136
rect 16256 13086 16272 13120
rect 16356 13086 16372 13120
rect 15854 13048 15884 13070
rect 16064 13048 16094 13074
rect 16256 13070 16372 13086
rect 16676 13120 16792 13136
rect 16676 13086 16692 13120
rect 16776 13086 16792 13120
rect 16274 13048 16304 13070
rect 16484 13048 16514 13074
rect 16676 13070 16792 13086
rect 17096 13120 17212 13136
rect 17096 13086 17112 13120
rect 17196 13086 17212 13120
rect 16694 13048 16724 13070
rect 16904 13048 16934 13074
rect 17096 13070 17212 13086
rect 17516 13120 17632 13136
rect 17516 13086 17532 13120
rect 17616 13086 17632 13120
rect 17114 13048 17144 13070
rect 17324 13048 17354 13074
rect 17516 13070 17632 13086
rect 17936 13120 18052 13136
rect 17936 13086 17952 13120
rect 18036 13086 18052 13120
rect 17534 13048 17564 13070
rect 17744 13048 17774 13074
rect 17936 13070 18052 13086
rect 18356 13120 18472 13136
rect 18356 13086 18372 13120
rect 18456 13086 18472 13120
rect 17954 13048 17984 13070
rect 18164 13048 18194 13074
rect 18356 13070 18472 13086
rect 18374 13048 18404 13070
rect 18584 13048 18614 13074
rect 10394 12022 10424 12048
rect 10604 12026 10634 12048
rect 10586 12010 10652 12026
rect 10814 12022 10844 12048
rect 11024 12026 11054 12048
rect 10586 11868 10602 12010
rect 10636 11868 10652 12010
rect 10394 11830 10424 11856
rect 10586 11852 10652 11868
rect 11006 12010 11072 12026
rect 11234 12022 11264 12048
rect 11444 12026 11474 12048
rect 11006 11868 11022 12010
rect 11056 11868 11072 12010
rect 10604 11830 10634 11852
rect 10814 11830 10844 11856
rect 11006 11852 11072 11868
rect 11426 12010 11492 12026
rect 11654 12022 11684 12048
rect 11864 12026 11894 12048
rect 11426 11868 11442 12010
rect 11476 11868 11492 12010
rect 11024 11830 11054 11852
rect 11234 11830 11264 11856
rect 11426 11852 11492 11868
rect 11846 12010 11912 12026
rect 12074 12022 12104 12048
rect 12284 12026 12314 12048
rect 11846 11868 11862 12010
rect 11896 11868 11912 12010
rect 11444 11830 11474 11852
rect 11654 11830 11684 11856
rect 11846 11852 11912 11868
rect 12266 12010 12332 12026
rect 12494 12022 12524 12048
rect 12704 12026 12734 12048
rect 12266 11868 12282 12010
rect 12316 11868 12332 12010
rect 11864 11830 11894 11852
rect 12074 11830 12104 11856
rect 12266 11852 12332 11868
rect 12686 12010 12752 12026
rect 12914 12022 12944 12048
rect 13124 12026 13154 12048
rect 12686 11868 12702 12010
rect 12736 11868 12752 12010
rect 12284 11830 12314 11852
rect 12494 11830 12524 11856
rect 12686 11852 12752 11868
rect 13106 12010 13172 12026
rect 13334 12022 13364 12048
rect 13544 12026 13574 12048
rect 13106 11868 13122 12010
rect 13156 11868 13172 12010
rect 12704 11830 12734 11852
rect 12914 11830 12944 11856
rect 13106 11852 13172 11868
rect 13526 12010 13592 12026
rect 13754 12022 13784 12048
rect 13964 12026 13994 12048
rect 13526 11868 13542 12010
rect 13576 11868 13592 12010
rect 13124 11830 13154 11852
rect 13334 11830 13364 11856
rect 13526 11852 13592 11868
rect 13946 12010 14012 12026
rect 14174 12022 14204 12048
rect 14384 12026 14414 12048
rect 13946 11868 13962 12010
rect 13996 11868 14012 12010
rect 13544 11830 13574 11852
rect 13754 11830 13784 11856
rect 13946 11852 14012 11868
rect 14366 12010 14432 12026
rect 14594 12022 14624 12048
rect 14804 12026 14834 12048
rect 14366 11868 14382 12010
rect 14416 11868 14432 12010
rect 13964 11830 13994 11852
rect 14174 11830 14204 11856
rect 14366 11852 14432 11868
rect 14786 12010 14852 12026
rect 15014 12022 15044 12048
rect 15224 12026 15254 12048
rect 14786 11868 14802 12010
rect 14836 11868 14852 12010
rect 14384 11830 14414 11852
rect 14594 11830 14624 11856
rect 14786 11852 14852 11868
rect 15206 12010 15272 12026
rect 15434 12022 15464 12048
rect 15644 12026 15674 12048
rect 15206 11868 15222 12010
rect 15256 11868 15272 12010
rect 14804 11830 14834 11852
rect 15014 11830 15044 11856
rect 15206 11852 15272 11868
rect 15626 12010 15692 12026
rect 15854 12022 15884 12048
rect 16064 12026 16094 12048
rect 15626 11868 15642 12010
rect 15676 11868 15692 12010
rect 15224 11830 15254 11852
rect 15434 11830 15464 11856
rect 15626 11852 15692 11868
rect 16046 12010 16112 12026
rect 16274 12022 16304 12048
rect 16484 12026 16514 12048
rect 16046 11868 16062 12010
rect 16096 11868 16112 12010
rect 15644 11830 15674 11852
rect 15854 11830 15884 11856
rect 16046 11852 16112 11868
rect 16466 12010 16532 12026
rect 16694 12022 16724 12048
rect 16904 12026 16934 12048
rect 16466 11868 16482 12010
rect 16516 11868 16532 12010
rect 16064 11830 16094 11852
rect 16274 11830 16304 11856
rect 16466 11852 16532 11868
rect 16886 12010 16952 12026
rect 17114 12022 17144 12048
rect 17324 12026 17354 12048
rect 16886 11868 16902 12010
rect 16936 11868 16952 12010
rect 16484 11830 16514 11852
rect 16694 11830 16724 11856
rect 16886 11852 16952 11868
rect 17306 12010 17372 12026
rect 17534 12022 17564 12048
rect 17744 12026 17774 12048
rect 17306 11868 17322 12010
rect 17356 11868 17372 12010
rect 16904 11830 16934 11852
rect 17114 11830 17144 11856
rect 17306 11852 17372 11868
rect 17726 12010 17792 12026
rect 17954 12022 17984 12048
rect 18164 12026 18194 12048
rect 17726 11868 17742 12010
rect 17776 11868 17792 12010
rect 17324 11830 17354 11852
rect 17534 11830 17564 11856
rect 17726 11852 17792 11868
rect 18146 12010 18212 12026
rect 18374 12022 18404 12048
rect 18584 12026 18614 12048
rect 18146 11868 18162 12010
rect 18196 11868 18212 12010
rect 17744 11830 17774 11852
rect 17954 11830 17984 11856
rect 18146 11852 18212 11868
rect 18566 12010 18632 12026
rect 18566 11868 18582 12010
rect 18616 11868 18632 12010
rect 18164 11830 18194 11852
rect 18374 11830 18404 11856
rect 18566 11852 18632 11868
rect 18584 11830 18614 11852
rect 10394 10808 10424 10830
rect 10376 10792 10492 10808
rect 10604 10804 10634 10830
rect 10814 10808 10844 10830
rect 10376 10758 10392 10792
rect 10476 10758 10492 10792
rect 10376 10742 10492 10758
rect 10796 10792 10912 10808
rect 11024 10804 11054 10830
rect 11234 10808 11264 10830
rect 10796 10758 10812 10792
rect 10896 10758 10912 10792
rect 10796 10742 10912 10758
rect 11216 10792 11332 10808
rect 11444 10804 11474 10830
rect 11654 10808 11684 10830
rect 11216 10758 11232 10792
rect 11316 10758 11332 10792
rect 11216 10742 11332 10758
rect 11636 10792 11752 10808
rect 11864 10804 11894 10830
rect 12074 10808 12104 10830
rect 11636 10758 11652 10792
rect 11736 10758 11752 10792
rect 11636 10742 11752 10758
rect 12056 10792 12172 10808
rect 12284 10804 12314 10830
rect 12494 10808 12524 10830
rect 12056 10758 12072 10792
rect 12156 10758 12172 10792
rect 12056 10742 12172 10758
rect 12476 10792 12592 10808
rect 12704 10804 12734 10830
rect 12914 10808 12944 10830
rect 12476 10758 12492 10792
rect 12576 10758 12592 10792
rect 12476 10742 12592 10758
rect 12896 10792 13012 10808
rect 13124 10804 13154 10830
rect 13334 10808 13364 10830
rect 12896 10758 12912 10792
rect 12996 10758 13012 10792
rect 12896 10742 13012 10758
rect 13316 10792 13432 10808
rect 13544 10804 13574 10830
rect 13754 10808 13784 10830
rect 13316 10758 13332 10792
rect 13416 10758 13432 10792
rect 13316 10742 13432 10758
rect 13736 10792 13852 10808
rect 13964 10804 13994 10830
rect 14174 10808 14204 10830
rect 13736 10758 13752 10792
rect 13836 10758 13852 10792
rect 13736 10742 13852 10758
rect 14156 10792 14272 10808
rect 14384 10804 14414 10830
rect 14594 10808 14624 10830
rect 14156 10758 14172 10792
rect 14256 10758 14272 10792
rect 14156 10742 14272 10758
rect 14576 10792 14692 10808
rect 14804 10804 14834 10830
rect 15014 10808 15044 10830
rect 14576 10758 14592 10792
rect 14676 10758 14692 10792
rect 14576 10742 14692 10758
rect 14996 10792 15112 10808
rect 15224 10804 15254 10830
rect 15434 10808 15464 10830
rect 14996 10758 15012 10792
rect 15096 10758 15112 10792
rect 14996 10742 15112 10758
rect 15416 10792 15532 10808
rect 15644 10804 15674 10830
rect 15854 10808 15884 10830
rect 15416 10758 15432 10792
rect 15516 10758 15532 10792
rect 15416 10742 15532 10758
rect 15836 10792 15952 10808
rect 16064 10804 16094 10830
rect 16274 10808 16304 10830
rect 15836 10758 15852 10792
rect 15936 10758 15952 10792
rect 15836 10742 15952 10758
rect 16256 10792 16372 10808
rect 16484 10804 16514 10830
rect 16694 10808 16724 10830
rect 16256 10758 16272 10792
rect 16356 10758 16372 10792
rect 16256 10742 16372 10758
rect 16676 10792 16792 10808
rect 16904 10804 16934 10830
rect 17114 10808 17144 10830
rect 16676 10758 16692 10792
rect 16776 10758 16792 10792
rect 16676 10742 16792 10758
rect 17096 10792 17212 10808
rect 17324 10804 17354 10830
rect 17534 10808 17564 10830
rect 17096 10758 17112 10792
rect 17196 10758 17212 10792
rect 17096 10742 17212 10758
rect 17516 10792 17632 10808
rect 17744 10804 17774 10830
rect 17954 10808 17984 10830
rect 17516 10758 17532 10792
rect 17616 10758 17632 10792
rect 17516 10742 17632 10758
rect 17936 10792 18052 10808
rect 18164 10804 18194 10830
rect 18374 10808 18404 10830
rect 17936 10758 17952 10792
rect 18036 10758 18052 10792
rect 17936 10742 18052 10758
rect 18356 10792 18472 10808
rect 18584 10804 18614 10830
rect 18356 10758 18372 10792
rect 18456 10758 18472 10792
rect 18356 10742 18472 10758
rect 10376 7901 10492 7918
rect 10376 7866 10392 7901
rect 10426 7900 10492 7901
rect 10476 7866 10492 7900
rect 10376 7850 10492 7866
rect 10796 7901 10912 7918
rect 10796 7866 10812 7901
rect 10846 7900 10912 7901
rect 10896 7866 10912 7900
rect 10796 7850 10912 7866
rect 11216 7901 11332 7918
rect 11216 7866 11232 7901
rect 11266 7900 11332 7901
rect 11316 7866 11332 7900
rect 11216 7850 11332 7866
rect 11636 7901 11752 7918
rect 11636 7866 11652 7901
rect 11686 7900 11752 7901
rect 11736 7866 11752 7900
rect 11636 7850 11752 7866
rect 12056 7901 12172 7918
rect 12056 7866 12072 7901
rect 12106 7900 12172 7901
rect 12156 7866 12172 7900
rect 12056 7850 12172 7866
rect 12476 7901 12592 7918
rect 12476 7866 12492 7901
rect 12526 7900 12592 7901
rect 12576 7866 12592 7900
rect 12476 7850 12592 7866
rect 12896 7901 13012 7918
rect 12896 7866 12912 7901
rect 12946 7900 13012 7901
rect 12996 7866 13012 7900
rect 12896 7850 13012 7866
rect 13316 7901 13432 7918
rect 13316 7866 13332 7901
rect 13366 7900 13432 7901
rect 13416 7866 13432 7900
rect 13316 7850 13432 7866
rect 13736 7901 13852 7918
rect 13736 7866 13752 7901
rect 13786 7900 13852 7901
rect 13836 7866 13852 7900
rect 13736 7850 13852 7866
rect 14156 7901 14272 7918
rect 14156 7866 14172 7901
rect 14206 7900 14272 7901
rect 14256 7866 14272 7900
rect 14156 7850 14272 7866
rect 14576 7901 14692 7918
rect 14576 7866 14592 7901
rect 14626 7900 14692 7901
rect 14676 7866 14692 7900
rect 14576 7850 14692 7866
rect 14996 7901 15112 7918
rect 14996 7866 15012 7901
rect 15046 7900 15112 7901
rect 15096 7866 15112 7900
rect 14996 7850 15112 7866
rect 15416 7901 15532 7918
rect 15416 7866 15432 7901
rect 15466 7900 15532 7901
rect 15516 7866 15532 7900
rect 15416 7850 15532 7866
rect 15836 7901 15952 7918
rect 15836 7866 15852 7901
rect 15886 7900 15952 7901
rect 15936 7866 15952 7900
rect 15836 7850 15952 7866
rect 16256 7901 16372 7918
rect 16256 7866 16272 7901
rect 16306 7900 16372 7901
rect 16356 7866 16372 7900
rect 16256 7850 16372 7866
rect 16676 7901 16792 7918
rect 16676 7866 16692 7901
rect 16726 7900 16792 7901
rect 16776 7866 16792 7900
rect 16676 7850 16792 7866
rect 17096 7901 17212 7918
rect 17096 7866 17112 7901
rect 17146 7900 17212 7901
rect 17196 7866 17212 7900
rect 17096 7850 17212 7866
rect 17516 7901 17632 7918
rect 17516 7866 17532 7901
rect 17566 7900 17632 7901
rect 17616 7866 17632 7900
rect 17516 7850 17632 7866
rect 17936 7901 18052 7918
rect 17936 7866 17952 7901
rect 17986 7900 18052 7901
rect 18036 7866 18052 7900
rect 17936 7850 18052 7866
rect 18356 7901 18472 7918
rect 18356 7866 18372 7901
rect 18406 7900 18472 7901
rect 18456 7866 18472 7900
rect 18356 7850 18472 7866
rect 5736 7044 5852 7062
rect 5736 7010 5752 7044
rect 5836 7010 5852 7044
rect 5736 6994 5852 7010
rect 6156 7044 6272 7062
rect 6156 7002 6172 7044
rect 6256 7010 6272 7044
rect 6206 7002 6272 7010
rect 6156 6994 6272 7002
rect 6576 7044 6692 7062
rect 6576 7002 6592 7044
rect 6676 7010 6692 7044
rect 6626 7002 6692 7010
rect 6576 6994 6692 7002
rect 6996 7044 7112 7062
rect 6996 7002 7012 7044
rect 7096 7010 7112 7044
rect 7046 7002 7112 7010
rect 6996 6994 7112 7002
rect 7416 7044 7532 7062
rect 7416 7002 7432 7044
rect 7516 7010 7532 7044
rect 7466 7002 7532 7010
rect 7416 6994 7532 7002
rect 7836 7044 7952 7062
rect 7836 7002 7852 7044
rect 7936 7010 7952 7044
rect 7886 7002 7952 7010
rect 7836 6994 7952 7002
rect 8256 7044 8372 7062
rect 8256 7002 8272 7044
rect 8356 7010 8372 7044
rect 8306 7002 8372 7010
rect 8256 6994 8372 7002
rect 8676 7044 8792 7062
rect 8676 7002 8692 7044
rect 8776 7010 8792 7044
rect 8726 7002 8792 7010
rect 8676 6994 8792 7002
rect 9096 7044 9212 7062
rect 9096 7002 9112 7044
rect 9196 7010 9212 7044
rect 9146 7002 9212 7010
rect 9096 6994 9212 7002
rect 5544 6964 5574 6990
rect 5754 6964 5784 6994
rect 5964 6964 5994 6990
rect 6156 6986 6222 6994
rect 6174 6964 6204 6986
rect 6384 6964 6414 6990
rect 6576 6986 6642 6994
rect 6594 6964 6624 6986
rect 6804 6964 6834 6990
rect 6996 6986 7062 6994
rect 7014 6964 7044 6986
rect 7224 6964 7254 6990
rect 7416 6986 7482 6994
rect 7434 6964 7464 6986
rect 7644 6964 7674 6990
rect 7836 6986 7902 6994
rect 7854 6964 7884 6986
rect 8064 6964 8094 6990
rect 8256 6986 8322 6994
rect 8274 6964 8304 6986
rect 8484 6964 8514 6990
rect 8676 6986 8742 6994
rect 8694 6964 8724 6986
rect 8904 6964 8934 6990
rect 9096 6986 9162 6994
rect 9114 6964 9144 6986
rect 5544 5938 5574 5964
rect 5754 5938 5784 5964
rect 5964 5938 5994 5964
rect 6174 5938 6204 5964
rect 6384 5942 6414 5964
rect 6366 5938 6432 5942
rect 6594 5938 6624 5964
rect 6804 5942 6834 5964
rect 6786 5938 6852 5942
rect 7014 5938 7044 5964
rect 7224 5942 7254 5964
rect 7206 5938 7272 5942
rect 7434 5938 7464 5964
rect 7644 5942 7674 5964
rect 7626 5938 7692 5942
rect 7854 5938 7884 5964
rect 8064 5942 8094 5964
rect 8046 5938 8112 5942
rect 8274 5938 8304 5964
rect 8484 5942 8514 5964
rect 8466 5938 8532 5942
rect 8694 5938 8724 5964
rect 8904 5942 8934 5964
rect 8886 5938 8952 5942
rect 9114 5938 9144 5964
rect 5526 5921 5642 5938
rect 5526 5886 5542 5921
rect 5576 5920 5642 5921
rect 5626 5886 5642 5920
rect 5526 5870 5642 5886
rect 5946 5921 6062 5938
rect 5946 5886 5962 5921
rect 5996 5920 6062 5921
rect 6046 5886 6062 5920
rect 5946 5870 6062 5886
rect 6366 5926 6482 5938
rect 6366 5886 6382 5926
rect 6416 5920 6482 5926
rect 6466 5886 6482 5920
rect 6366 5870 6482 5886
rect 6786 5926 6902 5938
rect 6786 5886 6802 5926
rect 6836 5920 6902 5926
rect 6886 5886 6902 5920
rect 6786 5870 6902 5886
rect 7206 5926 7322 5938
rect 7206 5886 7222 5926
rect 7256 5920 7322 5926
rect 7306 5886 7322 5920
rect 7206 5870 7322 5886
rect 7626 5926 7742 5938
rect 7626 5886 7642 5926
rect 7676 5920 7742 5926
rect 7726 5886 7742 5920
rect 7626 5870 7742 5886
rect 8046 5926 8162 5938
rect 8046 5886 8062 5926
rect 8096 5920 8162 5926
rect 8146 5886 8162 5920
rect 8046 5870 8162 5886
rect 8466 5926 8582 5938
rect 8466 5886 8482 5926
rect 8516 5920 8582 5926
rect 8566 5886 8582 5920
rect 8466 5870 8582 5886
rect 8886 5926 9002 5938
rect 8886 5886 8902 5926
rect 8936 5920 9002 5926
rect 8986 5886 9002 5920
rect 8886 5870 9002 5886
rect 3772 5421 3888 5438
rect 3772 5386 3788 5421
rect 3822 5420 3888 5421
rect 3872 5386 3888 5420
rect 3772 5370 3888 5386
rect 4192 5421 4308 5438
rect 4192 5386 4208 5421
rect 4242 5420 4308 5421
rect 4292 5386 4308 5420
rect 4192 5370 4308 5386
rect 2632 5340 2662 5366
rect 3580 5340 3610 5366
rect 3790 5340 3820 5370
rect 4000 5340 4030 5366
rect 4210 5340 4240 5370
rect 2632 4318 2662 4340
rect 3580 4318 3610 4340
rect 2614 4302 2680 4318
rect 2614 4159 2630 4302
rect 2664 4159 2680 4302
rect 2614 4143 2680 4159
rect 3562 4302 3628 4318
rect 3790 4314 3820 4340
rect 4000 4318 4030 4340
rect 3562 4159 3578 4302
rect 3612 4159 3628 4302
rect 3562 4143 3628 4159
rect 3982 4302 4048 4318
rect 4210 4314 4240 4340
rect 3982 4159 3998 4302
rect 4032 4159 4048 4302
rect 3982 4143 4048 4159
rect 4402 4193 4518 4210
rect 4402 4158 4418 4193
rect 4452 4192 4518 4193
rect 4502 4158 4518 4192
rect 2632 4112 2662 4143
rect 2728 4112 2758 4138
rect 3370 4112 3400 4138
rect 3580 4112 3610 4143
rect 3790 4112 3820 4138
rect 4000 4112 4030 4143
rect 4402 4142 4518 4158
rect 4822 4193 4938 4210
rect 4822 4158 4838 4193
rect 4872 4192 4938 4193
rect 4922 4158 4938 4192
rect 4822 4142 4938 4158
rect 4210 4112 4240 4138
rect 4420 4112 4450 4142
rect 4630 4112 4660 4138
rect 4840 4112 4870 4142
rect 2632 3086 2662 3112
rect 2728 3082 2758 3112
rect 3370 3082 3400 3112
rect 3580 3086 3610 3112
rect 3790 3082 3820 3112
rect 4000 3086 4030 3112
rect 4210 3082 4240 3112
rect 4420 3086 4450 3112
rect 4630 3082 4660 3112
rect 4840 3086 4870 3112
rect 2710 3066 2826 3082
rect 2710 3032 2726 3066
rect 2810 3032 2826 3066
rect 2710 3016 2826 3032
rect 3352 3065 3468 3082
rect 3352 3030 3368 3065
rect 3402 3064 3468 3065
rect 3452 3030 3468 3064
rect 3352 3014 3468 3030
rect 3772 3065 3888 3082
rect 3772 3030 3788 3065
rect 3822 3064 3888 3065
rect 3872 3030 3888 3064
rect 3772 3014 3888 3030
rect 4192 3065 4308 3082
rect 4192 3030 4208 3065
rect 4242 3064 4308 3065
rect 4292 3030 4308 3064
rect 4192 3014 4308 3030
rect 4612 3065 4728 3082
rect 4612 3030 4628 3065
rect 4662 3064 4728 3065
rect 4712 3030 4728 3064
rect 4612 3014 4728 3030
rect 5526 5429 5642 5446
rect 5526 5394 5542 5429
rect 5576 5428 5642 5429
rect 5626 5394 5642 5428
rect 5526 5378 5642 5394
rect 5946 5429 6062 5446
rect 5946 5394 5962 5429
rect 5996 5428 6062 5429
rect 6046 5394 6062 5428
rect 5946 5378 6062 5394
rect 6366 5429 6482 5446
rect 6366 5394 6382 5429
rect 6416 5428 6482 5429
rect 6466 5394 6482 5428
rect 6366 5378 6482 5394
rect 6786 5429 6902 5446
rect 6786 5394 6802 5429
rect 6836 5428 6902 5429
rect 6886 5394 6902 5428
rect 6786 5378 6902 5394
rect 7206 5429 7322 5446
rect 7206 5394 7222 5429
rect 7256 5428 7322 5429
rect 7306 5394 7322 5428
rect 7206 5378 7322 5394
rect 7626 5429 7742 5446
rect 7626 5394 7642 5429
rect 7676 5428 7742 5429
rect 7726 5394 7742 5428
rect 7626 5378 7742 5394
rect 8046 5429 8162 5446
rect 8046 5394 8062 5429
rect 8096 5428 8162 5429
rect 8146 5394 8162 5428
rect 8046 5378 8162 5394
rect 8466 5429 8582 5446
rect 8466 5394 8482 5429
rect 8516 5428 8582 5429
rect 8566 5394 8582 5428
rect 8466 5378 8582 5394
rect 8886 5429 9002 5446
rect 8886 5394 8902 5429
rect 8936 5428 9002 5429
rect 8986 5394 9002 5428
rect 8886 5378 9002 5394
rect 5544 5348 5574 5378
rect 5754 5348 5784 5374
rect 5964 5348 5994 5378
rect 6174 5348 6204 5374
rect 6384 5348 6414 5378
rect 6594 5348 6624 5374
rect 6804 5348 6834 5378
rect 7014 5348 7044 5374
rect 7224 5348 7254 5378
rect 7434 5348 7464 5374
rect 7644 5348 7674 5378
rect 7854 5348 7884 5374
rect 8064 5348 8094 5378
rect 8274 5348 8304 5374
rect 8484 5348 8514 5378
rect 8694 5348 8724 5374
rect 8904 5348 8934 5378
rect 9114 5348 9144 5374
rect 5544 4322 5574 4348
rect 5754 4317 5784 4348
rect 5964 4322 5994 4348
rect 6174 4317 6204 4348
rect 6384 4322 6414 4348
rect 6594 4317 6624 4348
rect 6804 4322 6834 4348
rect 7014 4317 7044 4348
rect 7224 4322 7254 4348
rect 7434 4317 7464 4348
rect 7644 4322 7674 4348
rect 7854 4317 7884 4348
rect 8064 4322 8094 4348
rect 8274 4317 8304 4348
rect 8484 4322 8514 4348
rect 8694 4317 8724 4348
rect 8904 4322 8934 4348
rect 9114 4317 9144 4348
rect 5736 4301 5802 4317
rect 5736 4159 5752 4301
rect 5786 4159 5802 4301
rect 5736 4143 5802 4159
rect 6156 4301 6222 4317
rect 6156 4159 6172 4301
rect 6206 4159 6222 4301
rect 6156 4143 6222 4159
rect 6576 4301 6642 4317
rect 6576 4159 6592 4301
rect 6626 4159 6642 4301
rect 6576 4143 6642 4159
rect 6996 4301 7062 4317
rect 6996 4159 7012 4301
rect 7046 4159 7062 4301
rect 6996 4143 7062 4159
rect 7416 4301 7482 4317
rect 7416 4159 7432 4301
rect 7466 4159 7482 4301
rect 7416 4143 7482 4159
rect 7836 4301 7902 4317
rect 7836 4159 7852 4301
rect 7886 4159 7902 4301
rect 7836 4143 7902 4159
rect 8256 4301 8322 4317
rect 8256 4159 8272 4301
rect 8306 4159 8322 4301
rect 8256 4143 8322 4159
rect 8676 4301 8742 4317
rect 8676 4159 8692 4301
rect 8726 4159 8742 4301
rect 8676 4143 8742 4159
rect 9096 4301 9162 4317
rect 9096 4159 9112 4301
rect 9146 4159 9162 4301
rect 9096 4143 9162 4159
rect 5544 4112 5574 4138
rect 5754 4112 5784 4143
rect 5964 4112 5994 4138
rect 6174 4112 6204 4143
rect 6384 4112 6414 4138
rect 6594 4112 6624 4143
rect 6804 4112 6834 4138
rect 7014 4112 7044 4143
rect 7224 4112 7254 4138
rect 7434 4112 7464 4143
rect 7644 4112 7674 4138
rect 7854 4112 7884 4143
rect 8064 4112 8094 4138
rect 8274 4112 8304 4143
rect 8484 4112 8514 4138
rect 8694 4112 8724 4143
rect 8904 4112 8934 4138
rect 9114 4112 9144 4143
rect 5544 3082 5574 3112
rect 5754 3086 5784 3112
rect 5964 3082 5994 3112
rect 6174 3086 6204 3112
rect 6384 3082 6414 3112
rect 6594 3086 6624 3112
rect 6804 3082 6834 3112
rect 7014 3086 7044 3112
rect 7224 3082 7254 3112
rect 7434 3086 7464 3112
rect 7644 3082 7674 3112
rect 7854 3086 7884 3112
rect 8064 3082 8094 3112
rect 8274 3086 8304 3112
rect 8484 3082 8514 3112
rect 8694 3086 8724 3112
rect 8904 3082 8934 3112
rect 9114 3086 9144 3112
rect 5526 3065 5642 3082
rect 5526 3030 5542 3065
rect 5576 3064 5642 3065
rect 5626 3030 5642 3064
rect 5526 3014 5642 3030
rect 5946 3065 6062 3082
rect 5946 3030 5962 3065
rect 5996 3064 6062 3065
rect 6046 3030 6062 3064
rect 5946 3014 6062 3030
rect 6366 3065 6482 3082
rect 6366 3030 6382 3065
rect 6416 3064 6482 3065
rect 6466 3030 6482 3064
rect 6366 3014 6482 3030
rect 6786 3065 6902 3082
rect 6786 3030 6802 3065
rect 6836 3064 6902 3065
rect 6886 3030 6902 3064
rect 6786 3014 6902 3030
rect 7206 3065 7322 3082
rect 7206 3030 7222 3065
rect 7256 3064 7322 3065
rect 7306 3030 7322 3064
rect 7206 3014 7322 3030
rect 7626 3065 7742 3082
rect 7626 3030 7642 3065
rect 7676 3064 7742 3065
rect 7726 3030 7742 3064
rect 7626 3014 7742 3030
rect 8046 3065 8162 3082
rect 8046 3030 8062 3065
rect 8096 3064 8162 3065
rect 8146 3030 8162 3064
rect 8046 3014 8162 3030
rect 8466 3065 8582 3082
rect 8466 3030 8482 3065
rect 8516 3064 8582 3065
rect 8566 3030 8582 3064
rect 8466 3014 8582 3030
rect 8886 3065 9002 3082
rect 8886 3030 8902 3065
rect 8936 3064 9002 3065
rect 8986 3030 9002 3064
rect 10394 7820 10424 7850
rect 10604 7820 10634 7846
rect 10814 7820 10844 7850
rect 11024 7820 11054 7846
rect 11234 7820 11264 7850
rect 11444 7820 11474 7846
rect 11654 7820 11684 7850
rect 11864 7820 11894 7846
rect 12074 7820 12104 7850
rect 12284 7820 12314 7846
rect 12494 7820 12524 7850
rect 12704 7820 12734 7846
rect 12914 7820 12944 7850
rect 13124 7820 13154 7846
rect 13334 7820 13364 7850
rect 13544 7820 13574 7846
rect 13754 7820 13784 7850
rect 13964 7820 13994 7846
rect 14174 7820 14204 7850
rect 14384 7820 14414 7846
rect 14594 7820 14624 7850
rect 14804 7820 14834 7846
rect 15014 7820 15044 7850
rect 15224 7820 15254 7846
rect 15434 7820 15464 7850
rect 15644 7820 15674 7846
rect 15854 7820 15884 7850
rect 16064 7820 16094 7846
rect 16274 7820 16304 7850
rect 16484 7820 16514 7846
rect 16694 7820 16724 7850
rect 16904 7820 16934 7846
rect 17114 7820 17144 7850
rect 17324 7820 17354 7846
rect 17534 7820 17564 7850
rect 17744 7820 17774 7846
rect 17954 7820 17984 7850
rect 18164 7820 18194 7846
rect 18374 7820 18404 7850
rect 18584 7820 18614 7846
rect 10394 6794 10424 6820
rect 10604 6789 10634 6820
rect 10814 6794 10844 6820
rect 11024 6789 11054 6820
rect 11234 6794 11264 6820
rect 11444 6789 11474 6820
rect 11654 6794 11684 6820
rect 11864 6789 11894 6820
rect 12074 6794 12104 6820
rect 12284 6789 12314 6820
rect 12494 6794 12524 6820
rect 12704 6789 12734 6820
rect 12914 6794 12944 6820
rect 13124 6789 13154 6820
rect 13334 6794 13364 6820
rect 13544 6789 13574 6820
rect 13754 6794 13784 6820
rect 13964 6789 13994 6820
rect 14174 6794 14204 6820
rect 14384 6789 14414 6820
rect 14594 6794 14624 6820
rect 14804 6789 14834 6820
rect 15014 6794 15044 6820
rect 15224 6789 15254 6820
rect 15434 6794 15464 6820
rect 15644 6789 15674 6820
rect 15854 6794 15884 6820
rect 16064 6789 16094 6820
rect 16274 6794 16304 6820
rect 16484 6789 16514 6820
rect 16694 6794 16724 6820
rect 16904 6789 16934 6820
rect 17114 6794 17144 6820
rect 17324 6789 17354 6820
rect 17534 6794 17564 6820
rect 17744 6789 17774 6820
rect 17954 6794 17984 6820
rect 18164 6789 18194 6820
rect 18374 6794 18404 6820
rect 18584 6789 18614 6820
rect 10586 6773 10652 6789
rect 10586 6631 10602 6773
rect 10636 6631 10652 6773
rect 10586 6615 10652 6631
rect 11006 6773 11072 6789
rect 11006 6631 11022 6773
rect 11056 6631 11072 6773
rect 11006 6615 11072 6631
rect 11426 6773 11492 6789
rect 11426 6631 11442 6773
rect 11476 6631 11492 6773
rect 11426 6615 11492 6631
rect 11846 6773 11912 6789
rect 11846 6631 11862 6773
rect 11896 6631 11912 6773
rect 11846 6615 11912 6631
rect 12266 6773 12332 6789
rect 12266 6631 12282 6773
rect 12316 6631 12332 6773
rect 12266 6615 12332 6631
rect 12686 6773 12752 6789
rect 12686 6631 12702 6773
rect 12736 6631 12752 6773
rect 12686 6615 12752 6631
rect 13106 6773 13172 6789
rect 13106 6631 13122 6773
rect 13156 6631 13172 6773
rect 13106 6615 13172 6631
rect 13526 6773 13592 6789
rect 13526 6631 13542 6773
rect 13576 6631 13592 6773
rect 13526 6615 13592 6631
rect 13946 6773 14012 6789
rect 13946 6631 13962 6773
rect 13996 6631 14012 6773
rect 13946 6615 14012 6631
rect 14366 6773 14432 6789
rect 14366 6631 14382 6773
rect 14416 6631 14432 6773
rect 14366 6615 14432 6631
rect 14786 6773 14852 6789
rect 14786 6631 14802 6773
rect 14836 6631 14852 6773
rect 14786 6615 14852 6631
rect 15206 6773 15272 6789
rect 15206 6631 15222 6773
rect 15256 6631 15272 6773
rect 15206 6615 15272 6631
rect 15626 6773 15692 6789
rect 15626 6631 15642 6773
rect 15676 6631 15692 6773
rect 15626 6615 15692 6631
rect 16046 6773 16112 6789
rect 16046 6631 16062 6773
rect 16096 6631 16112 6773
rect 16046 6615 16112 6631
rect 16466 6773 16532 6789
rect 16466 6631 16482 6773
rect 16516 6631 16532 6773
rect 16466 6615 16532 6631
rect 16886 6773 16952 6789
rect 16886 6631 16902 6773
rect 16936 6631 16952 6773
rect 16886 6615 16952 6631
rect 17306 6773 17372 6789
rect 17306 6631 17322 6773
rect 17356 6631 17372 6773
rect 17306 6615 17372 6631
rect 17726 6773 17792 6789
rect 17726 6631 17742 6773
rect 17776 6631 17792 6773
rect 17726 6615 17792 6631
rect 18146 6773 18212 6789
rect 18146 6631 18162 6773
rect 18196 6631 18212 6773
rect 18146 6615 18212 6631
rect 18566 6773 18632 6789
rect 18566 6631 18582 6773
rect 18616 6631 18632 6773
rect 18566 6615 18632 6631
rect 10394 6584 10424 6610
rect 10604 6584 10634 6615
rect 10814 6584 10844 6610
rect 11024 6584 11054 6615
rect 11234 6584 11264 6610
rect 11444 6584 11474 6615
rect 11654 6584 11684 6610
rect 11864 6584 11894 6615
rect 12074 6584 12104 6610
rect 12284 6584 12314 6615
rect 12494 6584 12524 6610
rect 12704 6584 12734 6615
rect 12914 6584 12944 6610
rect 13124 6584 13154 6615
rect 13334 6584 13364 6610
rect 13544 6584 13574 6615
rect 13754 6584 13784 6610
rect 13964 6584 13994 6615
rect 14174 6584 14204 6610
rect 14384 6584 14414 6615
rect 14594 6584 14624 6610
rect 14804 6584 14834 6615
rect 15014 6584 15044 6610
rect 15224 6584 15254 6615
rect 15434 6584 15464 6610
rect 15644 6584 15674 6615
rect 15854 6584 15884 6610
rect 16064 6584 16094 6615
rect 16274 6584 16304 6610
rect 16484 6584 16514 6615
rect 16694 6584 16724 6610
rect 16904 6584 16934 6615
rect 17114 6584 17144 6610
rect 17324 6584 17354 6615
rect 17534 6584 17564 6610
rect 17744 6584 17774 6615
rect 17954 6584 17984 6610
rect 18164 6584 18194 6615
rect 18374 6584 18404 6610
rect 18584 6584 18614 6615
rect 10394 5553 10424 5584
rect 10604 5558 10634 5584
rect 10814 5553 10844 5584
rect 11024 5558 11054 5584
rect 11234 5553 11264 5584
rect 11444 5558 11474 5584
rect 11654 5553 11684 5584
rect 11864 5558 11894 5584
rect 12074 5553 12104 5584
rect 12284 5558 12314 5584
rect 12494 5553 12524 5584
rect 12704 5558 12734 5584
rect 12914 5553 12944 5584
rect 13124 5558 13154 5584
rect 13334 5553 13364 5584
rect 13544 5558 13574 5584
rect 13754 5553 13784 5584
rect 13964 5558 13994 5584
rect 14174 5553 14204 5584
rect 14384 5558 14414 5584
rect 14594 5553 14624 5584
rect 14804 5558 14834 5584
rect 15014 5553 15044 5584
rect 15224 5558 15254 5584
rect 15434 5553 15464 5584
rect 15644 5558 15674 5584
rect 15854 5553 15884 5584
rect 16064 5558 16094 5584
rect 16274 5553 16304 5584
rect 16484 5558 16514 5584
rect 16694 5553 16724 5584
rect 16904 5558 16934 5584
rect 17114 5553 17144 5584
rect 17324 5558 17354 5584
rect 17534 5553 17564 5584
rect 17744 5558 17774 5584
rect 17954 5553 17984 5584
rect 18164 5558 18194 5584
rect 18374 5553 18404 5584
rect 18584 5558 18614 5584
rect 10376 5537 10442 5553
rect 10376 5395 10392 5537
rect 10426 5395 10442 5537
rect 10376 5379 10442 5395
rect 10796 5537 10862 5553
rect 10796 5395 10812 5537
rect 10846 5395 10862 5537
rect 10796 5379 10862 5395
rect 11216 5537 11282 5553
rect 11216 5395 11232 5537
rect 11266 5395 11282 5537
rect 11216 5379 11282 5395
rect 11636 5537 11702 5553
rect 11636 5395 11652 5537
rect 11686 5395 11702 5537
rect 11636 5379 11702 5395
rect 12056 5537 12122 5553
rect 12056 5395 12072 5537
rect 12106 5395 12122 5537
rect 12056 5379 12122 5395
rect 12476 5537 12542 5553
rect 12476 5395 12492 5537
rect 12526 5395 12542 5537
rect 12476 5379 12542 5395
rect 12896 5537 12962 5553
rect 12896 5395 12912 5537
rect 12946 5395 12962 5537
rect 12896 5379 12962 5395
rect 13316 5537 13382 5553
rect 13316 5395 13332 5537
rect 13366 5395 13382 5537
rect 13316 5379 13382 5395
rect 13736 5537 13802 5553
rect 13736 5395 13752 5537
rect 13786 5395 13802 5537
rect 13736 5379 13802 5395
rect 14156 5537 14222 5553
rect 14156 5395 14172 5537
rect 14206 5395 14222 5537
rect 14156 5379 14222 5395
rect 14576 5537 14642 5553
rect 14576 5395 14592 5537
rect 14626 5395 14642 5537
rect 14576 5379 14642 5395
rect 14996 5537 15062 5553
rect 14996 5395 15012 5537
rect 15046 5395 15062 5537
rect 14996 5379 15062 5395
rect 15416 5537 15482 5553
rect 15416 5395 15432 5537
rect 15466 5395 15482 5537
rect 15416 5379 15482 5395
rect 15836 5537 15902 5553
rect 15836 5395 15852 5537
rect 15886 5395 15902 5537
rect 15836 5379 15902 5395
rect 16256 5537 16322 5553
rect 16256 5395 16272 5537
rect 16306 5395 16322 5537
rect 16256 5379 16322 5395
rect 16676 5537 16742 5553
rect 16676 5395 16692 5537
rect 16726 5395 16742 5537
rect 16676 5379 16742 5395
rect 17096 5537 17162 5553
rect 17096 5395 17112 5537
rect 17146 5395 17162 5537
rect 17096 5379 17162 5395
rect 17516 5537 17582 5553
rect 17516 5395 17532 5537
rect 17566 5395 17582 5537
rect 17516 5379 17582 5395
rect 17936 5537 18002 5553
rect 17936 5395 17952 5537
rect 17986 5395 18002 5537
rect 17936 5379 18002 5395
rect 18356 5537 18422 5553
rect 18356 5395 18372 5537
rect 18406 5395 18422 5537
rect 18356 5379 18422 5395
rect 10394 5348 10424 5379
rect 10604 5348 10634 5374
rect 10814 5348 10844 5379
rect 11024 5348 11054 5374
rect 11234 5348 11264 5379
rect 11444 5348 11474 5374
rect 11654 5348 11684 5379
rect 11864 5348 11894 5374
rect 12074 5348 12104 5379
rect 12284 5348 12314 5374
rect 12494 5348 12524 5379
rect 12704 5348 12734 5374
rect 12914 5348 12944 5379
rect 13124 5348 13154 5374
rect 13334 5348 13364 5379
rect 13544 5348 13574 5374
rect 13754 5348 13784 5379
rect 13964 5348 13994 5374
rect 14174 5348 14204 5379
rect 14384 5348 14414 5374
rect 14594 5348 14624 5379
rect 14804 5348 14834 5374
rect 15014 5348 15044 5379
rect 15224 5348 15254 5374
rect 15434 5348 15464 5379
rect 15644 5348 15674 5374
rect 15854 5348 15884 5379
rect 16064 5348 16094 5374
rect 16274 5348 16304 5379
rect 16484 5348 16514 5374
rect 16694 5348 16724 5379
rect 16904 5348 16934 5374
rect 17114 5348 17144 5379
rect 17324 5348 17354 5374
rect 17534 5348 17564 5379
rect 17744 5348 17774 5374
rect 17954 5348 17984 5379
rect 18164 5348 18194 5374
rect 18374 5348 18404 5379
rect 18584 5348 18614 5374
rect 10394 4322 10424 4348
rect 10604 4317 10634 4348
rect 10814 4322 10844 4348
rect 11024 4317 11054 4348
rect 11234 4322 11264 4348
rect 11444 4317 11474 4348
rect 11654 4322 11684 4348
rect 11864 4317 11894 4348
rect 12074 4322 12104 4348
rect 12284 4317 12314 4348
rect 12494 4322 12524 4348
rect 12704 4317 12734 4348
rect 12914 4322 12944 4348
rect 13124 4317 13154 4348
rect 13334 4322 13364 4348
rect 13544 4317 13574 4348
rect 13754 4322 13784 4348
rect 13964 4317 13994 4348
rect 14174 4322 14204 4348
rect 14384 4317 14414 4348
rect 14594 4322 14624 4348
rect 14804 4317 14834 4348
rect 15014 4322 15044 4348
rect 15224 4317 15254 4348
rect 15434 4322 15464 4348
rect 15644 4317 15674 4348
rect 15854 4322 15884 4348
rect 16064 4317 16094 4348
rect 16274 4322 16304 4348
rect 16484 4317 16514 4348
rect 16694 4322 16724 4348
rect 16904 4317 16934 4348
rect 17114 4322 17144 4348
rect 17324 4317 17354 4348
rect 17534 4322 17564 4348
rect 17744 4317 17774 4348
rect 17954 4322 17984 4348
rect 18164 4317 18194 4348
rect 18374 4322 18404 4348
rect 18584 4317 18614 4348
rect 10586 4301 10652 4317
rect 10586 4159 10602 4301
rect 10636 4159 10652 4301
rect 10586 4143 10652 4159
rect 11006 4301 11072 4317
rect 11006 4159 11022 4301
rect 11056 4159 11072 4301
rect 11006 4143 11072 4159
rect 11426 4301 11492 4317
rect 11426 4159 11442 4301
rect 11476 4159 11492 4301
rect 11426 4143 11492 4159
rect 11846 4301 11912 4317
rect 11846 4159 11862 4301
rect 11896 4159 11912 4301
rect 11846 4143 11912 4159
rect 12266 4301 12332 4317
rect 12266 4159 12282 4301
rect 12316 4159 12332 4301
rect 12266 4143 12332 4159
rect 12686 4301 12752 4317
rect 12686 4159 12702 4301
rect 12736 4159 12752 4301
rect 12686 4143 12752 4159
rect 13106 4301 13172 4317
rect 13106 4159 13122 4301
rect 13156 4159 13172 4301
rect 13106 4143 13172 4159
rect 13526 4301 13592 4317
rect 13526 4159 13542 4301
rect 13576 4159 13592 4301
rect 13526 4143 13592 4159
rect 13946 4301 14012 4317
rect 13946 4159 13962 4301
rect 13996 4159 14012 4301
rect 13946 4143 14012 4159
rect 14366 4301 14432 4317
rect 14366 4159 14382 4301
rect 14416 4159 14432 4301
rect 14366 4143 14432 4159
rect 14786 4301 14852 4317
rect 14786 4159 14802 4301
rect 14836 4159 14852 4301
rect 14786 4143 14852 4159
rect 15206 4301 15272 4317
rect 15206 4159 15222 4301
rect 15256 4159 15272 4301
rect 15206 4143 15272 4159
rect 15626 4301 15692 4317
rect 15626 4159 15642 4301
rect 15676 4159 15692 4301
rect 15626 4143 15692 4159
rect 16046 4301 16112 4317
rect 16046 4159 16062 4301
rect 16096 4159 16112 4301
rect 16046 4143 16112 4159
rect 16466 4301 16532 4317
rect 16466 4159 16482 4301
rect 16516 4159 16532 4301
rect 16466 4143 16532 4159
rect 16886 4301 16952 4317
rect 16886 4159 16902 4301
rect 16936 4159 16952 4301
rect 16886 4143 16952 4159
rect 17306 4301 17372 4317
rect 17306 4159 17322 4301
rect 17356 4159 17372 4301
rect 17306 4143 17372 4159
rect 17726 4301 17792 4317
rect 17726 4159 17742 4301
rect 17776 4159 17792 4301
rect 17726 4143 17792 4159
rect 18146 4301 18212 4317
rect 18146 4159 18162 4301
rect 18196 4159 18212 4301
rect 18146 4143 18212 4159
rect 18566 4301 18632 4317
rect 18566 4159 18582 4301
rect 18616 4159 18632 4301
rect 18566 4143 18632 4159
rect 10394 4112 10424 4138
rect 10604 4112 10634 4143
rect 10814 4112 10844 4138
rect 11024 4112 11054 4143
rect 11234 4112 11264 4138
rect 11444 4112 11474 4143
rect 11654 4112 11684 4138
rect 11864 4112 11894 4143
rect 12074 4112 12104 4138
rect 12284 4112 12314 4143
rect 12494 4112 12524 4138
rect 12704 4112 12734 4143
rect 12914 4112 12944 4138
rect 13124 4112 13154 4143
rect 13334 4112 13364 4138
rect 13544 4112 13574 4143
rect 13754 4112 13784 4138
rect 13964 4112 13994 4143
rect 14174 4112 14204 4138
rect 14384 4112 14414 4143
rect 14594 4112 14624 4138
rect 14804 4112 14834 4143
rect 15014 4112 15044 4138
rect 15224 4112 15254 4143
rect 15434 4112 15464 4138
rect 15644 4112 15674 4143
rect 15854 4112 15884 4138
rect 16064 4112 16094 4143
rect 16274 4112 16304 4138
rect 16484 4112 16514 4143
rect 16694 4112 16724 4138
rect 16904 4112 16934 4143
rect 17114 4112 17144 4138
rect 17324 4112 17354 4143
rect 17534 4112 17564 4138
rect 17744 4112 17774 4143
rect 17954 4112 17984 4138
rect 18164 4112 18194 4143
rect 18374 4112 18404 4138
rect 18584 4112 18614 4143
rect 10394 3082 10424 3112
rect 10604 3086 10634 3112
rect 10814 3082 10844 3112
rect 11024 3086 11054 3112
rect 11234 3082 11264 3112
rect 11444 3086 11474 3112
rect 11654 3082 11684 3112
rect 11864 3086 11894 3112
rect 12074 3082 12104 3112
rect 12284 3086 12314 3112
rect 12494 3082 12524 3112
rect 12704 3086 12734 3112
rect 12914 3082 12944 3112
rect 13124 3086 13154 3112
rect 13334 3082 13364 3112
rect 13544 3086 13574 3112
rect 13754 3082 13784 3112
rect 13964 3086 13994 3112
rect 14174 3082 14204 3112
rect 14384 3086 14414 3112
rect 14594 3082 14624 3112
rect 14804 3086 14834 3112
rect 15014 3082 15044 3112
rect 15224 3086 15254 3112
rect 15434 3082 15464 3112
rect 15644 3086 15674 3112
rect 15854 3082 15884 3112
rect 16064 3086 16094 3112
rect 16274 3082 16304 3112
rect 16484 3086 16514 3112
rect 16694 3082 16724 3112
rect 16904 3086 16934 3112
rect 17114 3082 17144 3112
rect 17324 3086 17354 3112
rect 17534 3082 17564 3112
rect 17744 3086 17774 3112
rect 17954 3082 17984 3112
rect 18164 3086 18194 3112
rect 18374 3082 18404 3112
rect 18584 3086 18614 3112
rect 10376 3065 10492 3082
rect 8886 3014 9002 3030
rect 10376 3030 10392 3065
rect 10426 3064 10492 3065
rect 10476 3030 10492 3064
rect 10376 3014 10492 3030
rect 10796 3065 10912 3082
rect 10796 3030 10812 3065
rect 10846 3064 10912 3065
rect 10896 3030 10912 3064
rect 10796 3014 10912 3030
rect 11216 3065 11332 3082
rect 11216 3030 11232 3065
rect 11266 3064 11332 3065
rect 11316 3030 11332 3064
rect 11216 3014 11332 3030
rect 11636 3065 11752 3082
rect 11636 3030 11652 3065
rect 11686 3064 11752 3065
rect 11736 3030 11752 3064
rect 11636 3014 11752 3030
rect 12056 3065 12172 3082
rect 12056 3030 12072 3065
rect 12106 3064 12172 3065
rect 12156 3030 12172 3064
rect 12056 3014 12172 3030
rect 12476 3065 12592 3082
rect 12476 3030 12492 3065
rect 12526 3064 12592 3065
rect 12576 3030 12592 3064
rect 12476 3014 12592 3030
rect 12896 3065 13012 3082
rect 12896 3030 12912 3065
rect 12946 3064 13012 3065
rect 12996 3030 13012 3064
rect 12896 3014 13012 3030
rect 13316 3065 13432 3082
rect 13316 3030 13332 3065
rect 13366 3064 13432 3065
rect 13416 3030 13432 3064
rect 13316 3014 13432 3030
rect 13736 3065 13852 3082
rect 13736 3030 13752 3065
rect 13786 3064 13852 3065
rect 13836 3030 13852 3064
rect 13736 3014 13852 3030
rect 14156 3065 14272 3082
rect 14156 3030 14172 3065
rect 14206 3064 14272 3065
rect 14256 3030 14272 3064
rect 14156 3014 14272 3030
rect 14576 3065 14692 3082
rect 14576 3030 14592 3065
rect 14626 3064 14692 3065
rect 14676 3030 14692 3064
rect 14576 3014 14692 3030
rect 14996 3065 15112 3082
rect 14996 3030 15012 3065
rect 15046 3064 15112 3065
rect 15096 3030 15112 3064
rect 14996 3014 15112 3030
rect 15416 3065 15532 3082
rect 15416 3030 15432 3065
rect 15466 3064 15532 3065
rect 15516 3030 15532 3064
rect 15416 3014 15532 3030
rect 15836 3065 15952 3082
rect 15836 3030 15852 3065
rect 15886 3064 15952 3065
rect 15936 3030 15952 3064
rect 15836 3014 15952 3030
rect 16256 3065 16372 3082
rect 16256 3030 16272 3065
rect 16306 3064 16372 3065
rect 16356 3030 16372 3064
rect 16256 3014 16372 3030
rect 16676 3065 16792 3082
rect 16676 3030 16692 3065
rect 16726 3064 16792 3065
rect 16776 3030 16792 3064
rect 16676 3014 16792 3030
rect 17096 3065 17212 3082
rect 17096 3030 17112 3065
rect 17146 3064 17212 3065
rect 17196 3030 17212 3064
rect 17096 3014 17212 3030
rect 17516 3065 17632 3082
rect 17516 3030 17532 3065
rect 17566 3064 17632 3065
rect 17616 3030 17632 3064
rect 17516 3014 17632 3030
rect 17936 3065 18052 3082
rect 17936 3030 17952 3065
rect 17986 3064 18052 3065
rect 18036 3030 18052 3064
rect 17936 3014 18052 3030
rect 18356 3065 18472 3082
rect 18356 3030 18372 3065
rect 18406 3064 18472 3065
rect 18456 3030 18472 3064
rect 18356 3014 18472 3030
rect 2710 -1506 2826 -1490
rect 2710 -1540 2726 -1506
rect 2810 -1540 2826 -1506
rect 2710 -1556 2826 -1540
rect 3352 -1504 3468 -1488
rect 3352 -1539 3368 -1504
rect 3452 -1538 3468 -1504
rect 3402 -1539 3468 -1538
rect 3352 -1556 3468 -1539
rect 3772 -1504 3888 -1488
rect 3772 -1539 3788 -1504
rect 3872 -1538 3888 -1504
rect 3822 -1539 3888 -1538
rect 3772 -1556 3888 -1539
rect 4192 -1504 4308 -1488
rect 4192 -1539 4208 -1504
rect 4292 -1538 4308 -1504
rect 4242 -1539 4308 -1538
rect 4192 -1556 4308 -1539
rect 4612 -1504 4728 -1488
rect 4612 -1539 4628 -1504
rect 4712 -1538 4728 -1504
rect 4662 -1539 4728 -1538
rect 4612 -1556 4728 -1539
rect 2632 -1586 2662 -1560
rect 2728 -1586 2758 -1556
rect 3370 -1586 3400 -1556
rect 3580 -1586 3610 -1560
rect 3790 -1586 3820 -1556
rect 4000 -1586 4030 -1560
rect 4210 -1586 4240 -1556
rect 4420 -1586 4450 -1560
rect 4630 -1586 4660 -1556
rect 4840 -1586 4870 -1560
rect 2632 -2617 2662 -2586
rect 2728 -2612 2758 -2586
rect 3370 -2612 3400 -2586
rect 3580 -2617 3610 -2586
rect 3790 -2612 3820 -2586
rect 4000 -2617 4030 -2586
rect 4210 -2612 4240 -2586
rect 4420 -2616 4450 -2586
rect 4630 -2612 4660 -2586
rect 4840 -2616 4870 -2586
rect 2614 -2633 2680 -2617
rect 2614 -2776 2630 -2633
rect 2664 -2776 2680 -2633
rect 2614 -2792 2680 -2776
rect 3562 -2633 3628 -2617
rect 3562 -2776 3578 -2633
rect 3612 -2776 3628 -2633
rect 3562 -2792 3628 -2776
rect 3982 -2633 4048 -2617
rect 3982 -2776 3998 -2633
rect 4032 -2776 4048 -2633
rect 4402 -2632 4518 -2616
rect 4402 -2667 4418 -2632
rect 4502 -2666 4518 -2632
rect 4452 -2667 4518 -2666
rect 4402 -2684 4518 -2667
rect 4822 -2632 4938 -2616
rect 4822 -2667 4838 -2632
rect 4922 -2666 4938 -2632
rect 4872 -2667 4938 -2666
rect 4822 -2684 4938 -2667
rect 2632 -2814 2662 -2792
rect 3580 -2814 3610 -2792
rect 3790 -2814 3820 -2788
rect 3982 -2792 4048 -2776
rect 4000 -2814 4030 -2792
rect 4210 -2814 4240 -2788
rect 2632 -3840 2662 -3814
rect 3580 -3840 3610 -3814
rect 3790 -3844 3820 -3814
rect 4000 -3840 4030 -3814
rect 4210 -3844 4240 -3814
rect 3772 -3860 3888 -3844
rect 3772 -3895 3788 -3860
rect 3872 -3894 3888 -3860
rect 3822 -3895 3888 -3894
rect 3772 -3912 3888 -3895
rect 4192 -3860 4308 -3844
rect 4192 -3895 4208 -3860
rect 4292 -3894 4308 -3860
rect 4242 -3895 4308 -3894
rect 4192 -3912 4308 -3895
rect 5526 -1504 5642 -1488
rect 5526 -1539 5542 -1504
rect 5626 -1538 5642 -1504
rect 5576 -1539 5642 -1538
rect 5526 -1556 5642 -1539
rect 5946 -1504 6062 -1488
rect 5946 -1539 5962 -1504
rect 6046 -1538 6062 -1504
rect 5996 -1539 6062 -1538
rect 5946 -1556 6062 -1539
rect 6366 -1504 6482 -1488
rect 6366 -1539 6382 -1504
rect 6466 -1538 6482 -1504
rect 6416 -1539 6482 -1538
rect 6366 -1556 6482 -1539
rect 6786 -1504 6902 -1488
rect 6786 -1539 6802 -1504
rect 6886 -1538 6902 -1504
rect 6836 -1539 6902 -1538
rect 6786 -1556 6902 -1539
rect 7206 -1504 7322 -1488
rect 7206 -1539 7222 -1504
rect 7306 -1538 7322 -1504
rect 7256 -1539 7322 -1538
rect 7206 -1556 7322 -1539
rect 7626 -1504 7742 -1488
rect 7626 -1539 7642 -1504
rect 7726 -1538 7742 -1504
rect 7676 -1539 7742 -1538
rect 7626 -1556 7742 -1539
rect 8046 -1504 8162 -1488
rect 8046 -1539 8062 -1504
rect 8146 -1538 8162 -1504
rect 8096 -1539 8162 -1538
rect 8046 -1556 8162 -1539
rect 8466 -1504 8582 -1488
rect 8466 -1539 8482 -1504
rect 8566 -1538 8582 -1504
rect 8516 -1539 8582 -1538
rect 8466 -1556 8582 -1539
rect 8886 -1504 9002 -1488
rect 8886 -1539 8902 -1504
rect 8986 -1538 9002 -1504
rect 8936 -1539 9002 -1538
rect 8886 -1556 9002 -1539
rect 5544 -1586 5574 -1556
rect 5754 -1586 5784 -1560
rect 5964 -1586 5994 -1556
rect 6174 -1586 6204 -1560
rect 6384 -1586 6414 -1556
rect 6594 -1586 6624 -1560
rect 6804 -1586 6834 -1556
rect 7014 -1586 7044 -1560
rect 7224 -1586 7254 -1556
rect 7434 -1586 7464 -1560
rect 7644 -1586 7674 -1556
rect 7854 -1586 7884 -1560
rect 8064 -1586 8094 -1556
rect 8274 -1586 8304 -1560
rect 8484 -1586 8514 -1556
rect 8694 -1586 8724 -1560
rect 8904 -1586 8934 -1556
rect 9114 -1586 9144 -1560
rect 5544 -2612 5574 -2586
rect 5754 -2617 5784 -2586
rect 5964 -2612 5994 -2586
rect 6174 -2617 6204 -2586
rect 6384 -2612 6414 -2586
rect 6594 -2617 6624 -2586
rect 6804 -2612 6834 -2586
rect 7014 -2617 7044 -2586
rect 7224 -2612 7254 -2586
rect 7434 -2617 7464 -2586
rect 7644 -2612 7674 -2586
rect 7854 -2617 7884 -2586
rect 8064 -2612 8094 -2586
rect 8274 -2617 8304 -2586
rect 8484 -2612 8514 -2586
rect 8694 -2617 8724 -2586
rect 8904 -2612 8934 -2586
rect 9114 -2617 9144 -2586
rect 5736 -2633 5802 -2617
rect 5736 -2775 5752 -2633
rect 5786 -2775 5802 -2633
rect 5736 -2791 5802 -2775
rect 6156 -2633 6222 -2617
rect 6156 -2775 6172 -2633
rect 6206 -2775 6222 -2633
rect 6156 -2791 6222 -2775
rect 6576 -2633 6642 -2617
rect 6576 -2775 6592 -2633
rect 6626 -2775 6642 -2633
rect 6576 -2791 6642 -2775
rect 6996 -2633 7062 -2617
rect 6996 -2775 7012 -2633
rect 7046 -2775 7062 -2633
rect 6996 -2791 7062 -2775
rect 7416 -2633 7482 -2617
rect 7416 -2775 7432 -2633
rect 7466 -2775 7482 -2633
rect 7416 -2791 7482 -2775
rect 7836 -2633 7902 -2617
rect 7836 -2775 7852 -2633
rect 7886 -2775 7902 -2633
rect 7836 -2791 7902 -2775
rect 8256 -2633 8322 -2617
rect 8256 -2775 8272 -2633
rect 8306 -2775 8322 -2633
rect 8256 -2791 8322 -2775
rect 8676 -2633 8742 -2617
rect 8676 -2775 8692 -2633
rect 8726 -2775 8742 -2633
rect 8676 -2791 8742 -2775
rect 9096 -2633 9162 -2617
rect 9096 -2775 9112 -2633
rect 9146 -2775 9162 -2633
rect 9096 -2791 9162 -2775
rect 5544 -2822 5574 -2796
rect 5754 -2822 5784 -2791
rect 5964 -2822 5994 -2796
rect 6174 -2822 6204 -2791
rect 6384 -2822 6414 -2796
rect 6594 -2822 6624 -2791
rect 6804 -2822 6834 -2796
rect 7014 -2822 7044 -2791
rect 7224 -2822 7254 -2796
rect 7434 -2822 7464 -2791
rect 7644 -2822 7674 -2796
rect 7854 -2822 7884 -2791
rect 8064 -2822 8094 -2796
rect 8274 -2822 8304 -2791
rect 8484 -2822 8514 -2796
rect 8694 -2822 8724 -2791
rect 8904 -2822 8934 -2796
rect 9114 -2822 9144 -2791
rect 5544 -3852 5574 -3822
rect 5754 -3848 5784 -3822
rect 5964 -3852 5994 -3822
rect 6174 -3848 6204 -3822
rect 6384 -3852 6414 -3822
rect 6594 -3848 6624 -3822
rect 6804 -3852 6834 -3822
rect 7014 -3848 7044 -3822
rect 7224 -3852 7254 -3822
rect 7434 -3848 7464 -3822
rect 7644 -3852 7674 -3822
rect 7854 -3848 7884 -3822
rect 8064 -3852 8094 -3822
rect 8274 -3848 8304 -3822
rect 8484 -3852 8514 -3822
rect 8694 -3848 8724 -3822
rect 8904 -3852 8934 -3822
rect 9114 -3848 9144 -3822
rect 5526 -3868 5642 -3852
rect 5526 -3903 5542 -3868
rect 5626 -3902 5642 -3868
rect 5576 -3903 5642 -3902
rect 5526 -3920 5642 -3903
rect 5946 -3868 6062 -3852
rect 5946 -3903 5962 -3868
rect 6046 -3902 6062 -3868
rect 5996 -3903 6062 -3902
rect 5946 -3920 6062 -3903
rect 6366 -3868 6482 -3852
rect 6366 -3903 6382 -3868
rect 6466 -3902 6482 -3868
rect 6416 -3903 6482 -3902
rect 6366 -3920 6482 -3903
rect 6786 -3868 6902 -3852
rect 6786 -3903 6802 -3868
rect 6886 -3902 6902 -3868
rect 6836 -3903 6902 -3902
rect 6786 -3920 6902 -3903
rect 7206 -3868 7322 -3852
rect 7206 -3903 7222 -3868
rect 7306 -3902 7322 -3868
rect 7256 -3903 7322 -3902
rect 7206 -3920 7322 -3903
rect 7626 -3868 7742 -3852
rect 7626 -3903 7642 -3868
rect 7726 -3902 7742 -3868
rect 7676 -3903 7742 -3902
rect 7626 -3920 7742 -3903
rect 8046 -3868 8162 -3852
rect 8046 -3903 8062 -3868
rect 8146 -3902 8162 -3868
rect 8096 -3903 8162 -3902
rect 8046 -3920 8162 -3903
rect 8466 -3868 8582 -3852
rect 8466 -3903 8482 -3868
rect 8566 -3902 8582 -3868
rect 8516 -3903 8582 -3902
rect 8466 -3920 8582 -3903
rect 8886 -3868 9002 -3852
rect 8886 -3903 8902 -3868
rect 8986 -3902 9002 -3868
rect 8936 -3903 9002 -3902
rect 8886 -3920 9002 -3903
rect 5526 -5760 5642 -5744
rect 5526 -5795 5542 -5760
rect 5626 -5794 5642 -5760
rect 5576 -5795 5642 -5794
rect 5526 -5812 5642 -5795
rect 5946 -5760 6062 -5744
rect 5946 -5795 5962 -5760
rect 6046 -5794 6062 -5760
rect 5996 -5795 6062 -5794
rect 5946 -5812 6062 -5795
rect 6366 -5760 6482 -5744
rect 6366 -5800 6382 -5760
rect 6466 -5794 6482 -5760
rect 6416 -5800 6482 -5794
rect 6366 -5812 6482 -5800
rect 6786 -5760 6902 -5744
rect 6786 -5800 6802 -5760
rect 6886 -5794 6902 -5760
rect 6836 -5800 6902 -5794
rect 6786 -5812 6902 -5800
rect 7206 -5760 7322 -5744
rect 7206 -5800 7222 -5760
rect 7306 -5794 7322 -5760
rect 7256 -5800 7322 -5794
rect 7206 -5812 7322 -5800
rect 7626 -5760 7742 -5744
rect 7626 -5800 7642 -5760
rect 7726 -5794 7742 -5760
rect 7676 -5800 7742 -5794
rect 7626 -5812 7742 -5800
rect 8046 -5760 8162 -5744
rect 8046 -5800 8062 -5760
rect 8146 -5794 8162 -5760
rect 8096 -5800 8162 -5794
rect 8046 -5812 8162 -5800
rect 8466 -5760 8582 -5744
rect 8466 -5800 8482 -5760
rect 8566 -5794 8582 -5760
rect 8516 -5800 8582 -5794
rect 8466 -5812 8582 -5800
rect 8886 -5760 9002 -5744
rect 8886 -5800 8902 -5760
rect 8986 -5794 9002 -5760
rect 8936 -5800 9002 -5794
rect 8886 -5812 9002 -5800
rect 5544 -5838 5574 -5812
rect 5754 -5838 5784 -5812
rect 5964 -5838 5994 -5812
rect 6174 -5838 6204 -5812
rect 6366 -5816 6432 -5812
rect 6384 -5838 6414 -5816
rect 6594 -5838 6624 -5812
rect 6786 -5816 6852 -5812
rect 6804 -5838 6834 -5816
rect 7014 -5838 7044 -5812
rect 7206 -5816 7272 -5812
rect 7224 -5838 7254 -5816
rect 7434 -5838 7464 -5812
rect 7626 -5816 7692 -5812
rect 7644 -5838 7674 -5816
rect 7854 -5838 7884 -5812
rect 8046 -5816 8112 -5812
rect 8064 -5838 8094 -5816
rect 8274 -5838 8304 -5812
rect 8466 -5816 8532 -5812
rect 8484 -5838 8514 -5816
rect 8694 -5838 8724 -5812
rect 8886 -5816 8952 -5812
rect 8904 -5838 8934 -5816
rect 9114 -5838 9144 -5812
rect 5544 -6864 5574 -6838
rect 5754 -6868 5784 -6838
rect 5964 -6864 5994 -6838
rect 6174 -6860 6204 -6838
rect 6156 -6868 6222 -6860
rect 6384 -6864 6414 -6838
rect 6594 -6860 6624 -6838
rect 6576 -6868 6642 -6860
rect 6804 -6864 6834 -6838
rect 7014 -6860 7044 -6838
rect 6996 -6868 7062 -6860
rect 7224 -6864 7254 -6838
rect 7434 -6860 7464 -6838
rect 7416 -6868 7482 -6860
rect 7644 -6864 7674 -6838
rect 7854 -6860 7884 -6838
rect 7836 -6868 7902 -6860
rect 8064 -6864 8094 -6838
rect 8274 -6860 8304 -6838
rect 8256 -6868 8322 -6860
rect 8484 -6864 8514 -6838
rect 8694 -6860 8724 -6838
rect 8676 -6868 8742 -6860
rect 8904 -6864 8934 -6838
rect 9114 -6860 9144 -6838
rect 9096 -6868 9162 -6860
rect 5736 -6884 5852 -6868
rect 5736 -6918 5752 -6884
rect 5836 -6918 5852 -6884
rect 5736 -6936 5852 -6918
rect 6156 -6876 6272 -6868
rect 6156 -6918 6172 -6876
rect 6206 -6884 6272 -6876
rect 6256 -6918 6272 -6884
rect 6156 -6936 6272 -6918
rect 6576 -6876 6692 -6868
rect 6576 -6918 6592 -6876
rect 6626 -6884 6692 -6876
rect 6676 -6918 6692 -6884
rect 6576 -6936 6692 -6918
rect 6996 -6876 7112 -6868
rect 6996 -6918 7012 -6876
rect 7046 -6884 7112 -6876
rect 7096 -6918 7112 -6884
rect 6996 -6936 7112 -6918
rect 7416 -6876 7532 -6868
rect 7416 -6918 7432 -6876
rect 7466 -6884 7532 -6876
rect 7516 -6918 7532 -6884
rect 7416 -6936 7532 -6918
rect 7836 -6876 7952 -6868
rect 7836 -6918 7852 -6876
rect 7886 -6884 7952 -6876
rect 7936 -6918 7952 -6884
rect 7836 -6936 7952 -6918
rect 8256 -6876 8372 -6868
rect 8256 -6918 8272 -6876
rect 8306 -6884 8372 -6876
rect 8356 -6918 8372 -6884
rect 8256 -6936 8372 -6918
rect 8676 -6876 8792 -6868
rect 8676 -6918 8692 -6876
rect 8726 -6884 8792 -6876
rect 8776 -6918 8792 -6884
rect 8676 -6936 8792 -6918
rect 9096 -6876 9212 -6868
rect 9096 -6918 9112 -6876
rect 9146 -6884 9212 -6876
rect 9196 -6918 9212 -6884
rect 9096 -6936 9212 -6918
<< polycont >>
rect 10392 13086 10476 13120
rect 10812 13086 10896 13120
rect 11232 13086 11316 13120
rect 11652 13086 11736 13120
rect 12072 13086 12156 13120
rect 12492 13086 12576 13120
rect 12912 13086 12996 13120
rect 13332 13086 13416 13120
rect 13752 13086 13836 13120
rect 14172 13086 14256 13120
rect 14592 13086 14676 13120
rect 15012 13086 15096 13120
rect 15432 13086 15516 13120
rect 15852 13086 15936 13120
rect 16272 13086 16356 13120
rect 16692 13086 16776 13120
rect 17112 13086 17196 13120
rect 17532 13086 17616 13120
rect 17952 13086 18036 13120
rect 18372 13086 18456 13120
rect 10602 11868 10636 12010
rect 11022 11868 11056 12010
rect 11442 11868 11476 12010
rect 11862 11868 11896 12010
rect 12282 11868 12316 12010
rect 12702 11868 12736 12010
rect 13122 11868 13156 12010
rect 13542 11868 13576 12010
rect 13962 11868 13996 12010
rect 14382 11868 14416 12010
rect 14802 11868 14836 12010
rect 15222 11868 15256 12010
rect 15642 11868 15676 12010
rect 16062 11868 16096 12010
rect 16482 11868 16516 12010
rect 16902 11868 16936 12010
rect 17322 11868 17356 12010
rect 17742 11868 17776 12010
rect 18162 11868 18196 12010
rect 18582 11868 18616 12010
rect 10392 10758 10476 10792
rect 10812 10758 10896 10792
rect 11232 10758 11316 10792
rect 11652 10758 11736 10792
rect 12072 10758 12156 10792
rect 12492 10758 12576 10792
rect 12912 10758 12996 10792
rect 13332 10758 13416 10792
rect 13752 10758 13836 10792
rect 14172 10758 14256 10792
rect 14592 10758 14676 10792
rect 15012 10758 15096 10792
rect 15432 10758 15516 10792
rect 15852 10758 15936 10792
rect 16272 10758 16356 10792
rect 16692 10758 16776 10792
rect 17112 10758 17196 10792
rect 17532 10758 17616 10792
rect 17952 10758 18036 10792
rect 18372 10758 18456 10792
rect 10392 7900 10426 7901
rect 10392 7866 10476 7900
rect 10812 7900 10846 7901
rect 10812 7866 10896 7900
rect 11232 7900 11266 7901
rect 11232 7866 11316 7900
rect 11652 7900 11686 7901
rect 11652 7866 11736 7900
rect 12072 7900 12106 7901
rect 12072 7866 12156 7900
rect 12492 7900 12526 7901
rect 12492 7866 12576 7900
rect 12912 7900 12946 7901
rect 12912 7866 12996 7900
rect 13332 7900 13366 7901
rect 13332 7866 13416 7900
rect 13752 7900 13786 7901
rect 13752 7866 13836 7900
rect 14172 7900 14206 7901
rect 14172 7866 14256 7900
rect 14592 7900 14626 7901
rect 14592 7866 14676 7900
rect 15012 7900 15046 7901
rect 15012 7866 15096 7900
rect 15432 7900 15466 7901
rect 15432 7866 15516 7900
rect 15852 7900 15886 7901
rect 15852 7866 15936 7900
rect 16272 7900 16306 7901
rect 16272 7866 16356 7900
rect 16692 7900 16726 7901
rect 16692 7866 16776 7900
rect 17112 7900 17146 7901
rect 17112 7866 17196 7900
rect 17532 7900 17566 7901
rect 17532 7866 17616 7900
rect 17952 7900 17986 7901
rect 17952 7866 18036 7900
rect 18372 7900 18406 7901
rect 18372 7866 18456 7900
rect 5752 7010 5836 7044
rect 6172 7010 6256 7044
rect 6172 7002 6206 7010
rect 6592 7010 6676 7044
rect 6592 7002 6626 7010
rect 7012 7010 7096 7044
rect 7012 7002 7046 7010
rect 7432 7010 7516 7044
rect 7432 7002 7466 7010
rect 7852 7010 7936 7044
rect 7852 7002 7886 7010
rect 8272 7010 8356 7044
rect 8272 7002 8306 7010
rect 8692 7010 8776 7044
rect 8692 7002 8726 7010
rect 9112 7010 9196 7044
rect 9112 7002 9146 7010
rect 5542 5920 5576 5921
rect 5542 5886 5626 5920
rect 5962 5920 5996 5921
rect 5962 5886 6046 5920
rect 6382 5920 6416 5926
rect 6382 5886 6466 5920
rect 6802 5920 6836 5926
rect 6802 5886 6886 5920
rect 7222 5920 7256 5926
rect 7222 5886 7306 5920
rect 7642 5920 7676 5926
rect 7642 5886 7726 5920
rect 8062 5920 8096 5926
rect 8062 5886 8146 5920
rect 8482 5920 8516 5926
rect 8482 5886 8566 5920
rect 8902 5920 8936 5926
rect 8902 5886 8986 5920
rect 3788 5420 3822 5421
rect 3788 5386 3872 5420
rect 4208 5420 4242 5421
rect 4208 5386 4292 5420
rect 2630 4159 2664 4302
rect 3578 4159 3612 4302
rect 3998 4159 4032 4302
rect 4418 4192 4452 4193
rect 4418 4158 4502 4192
rect 4838 4192 4872 4193
rect 4838 4158 4922 4192
rect 2726 3032 2810 3066
rect 3368 3064 3402 3065
rect 3368 3030 3452 3064
rect 3788 3064 3822 3065
rect 3788 3030 3872 3064
rect 4208 3064 4242 3065
rect 4208 3030 4292 3064
rect 4628 3064 4662 3065
rect 4628 3030 4712 3064
rect 5542 5428 5576 5429
rect 5542 5394 5626 5428
rect 5962 5428 5996 5429
rect 5962 5394 6046 5428
rect 6382 5428 6416 5429
rect 6382 5394 6466 5428
rect 6802 5428 6836 5429
rect 6802 5394 6886 5428
rect 7222 5428 7256 5429
rect 7222 5394 7306 5428
rect 7642 5428 7676 5429
rect 7642 5394 7726 5428
rect 8062 5428 8096 5429
rect 8062 5394 8146 5428
rect 8482 5428 8516 5429
rect 8482 5394 8566 5428
rect 8902 5428 8936 5429
rect 8902 5394 8986 5428
rect 5752 4159 5786 4301
rect 6172 4159 6206 4301
rect 6592 4159 6626 4301
rect 7012 4159 7046 4301
rect 7432 4159 7466 4301
rect 7852 4159 7886 4301
rect 8272 4159 8306 4301
rect 8692 4159 8726 4301
rect 9112 4159 9146 4301
rect 5542 3064 5576 3065
rect 5542 3030 5626 3064
rect 5962 3064 5996 3065
rect 5962 3030 6046 3064
rect 6382 3064 6416 3065
rect 6382 3030 6466 3064
rect 6802 3064 6836 3065
rect 6802 3030 6886 3064
rect 7222 3064 7256 3065
rect 7222 3030 7306 3064
rect 7642 3064 7676 3065
rect 7642 3030 7726 3064
rect 8062 3064 8096 3065
rect 8062 3030 8146 3064
rect 8482 3064 8516 3065
rect 8482 3030 8566 3064
rect 8902 3064 8936 3065
rect 8902 3030 8986 3064
rect 10602 6631 10636 6773
rect 11022 6631 11056 6773
rect 11442 6631 11476 6773
rect 11862 6631 11896 6773
rect 12282 6631 12316 6773
rect 12702 6631 12736 6773
rect 13122 6631 13156 6773
rect 13542 6631 13576 6773
rect 13962 6631 13996 6773
rect 14382 6631 14416 6773
rect 14802 6631 14836 6773
rect 15222 6631 15256 6773
rect 15642 6631 15676 6773
rect 16062 6631 16096 6773
rect 16482 6631 16516 6773
rect 16902 6631 16936 6773
rect 17322 6631 17356 6773
rect 17742 6631 17776 6773
rect 18162 6631 18196 6773
rect 18582 6631 18616 6773
rect 10392 5395 10426 5537
rect 10812 5395 10846 5537
rect 11232 5395 11266 5537
rect 11652 5395 11686 5537
rect 12072 5395 12106 5537
rect 12492 5395 12526 5537
rect 12912 5395 12946 5537
rect 13332 5395 13366 5537
rect 13752 5395 13786 5537
rect 14172 5395 14206 5537
rect 14592 5395 14626 5537
rect 15012 5395 15046 5537
rect 15432 5395 15466 5537
rect 15852 5395 15886 5537
rect 16272 5395 16306 5537
rect 16692 5395 16726 5537
rect 17112 5395 17146 5537
rect 17532 5395 17566 5537
rect 17952 5395 17986 5537
rect 18372 5395 18406 5537
rect 10602 4159 10636 4301
rect 11022 4159 11056 4301
rect 11442 4159 11476 4301
rect 11862 4159 11896 4301
rect 12282 4159 12316 4301
rect 12702 4159 12736 4301
rect 13122 4159 13156 4301
rect 13542 4159 13576 4301
rect 13962 4159 13996 4301
rect 14382 4159 14416 4301
rect 14802 4159 14836 4301
rect 15222 4159 15256 4301
rect 15642 4159 15676 4301
rect 16062 4159 16096 4301
rect 16482 4159 16516 4301
rect 16902 4159 16936 4301
rect 17322 4159 17356 4301
rect 17742 4159 17776 4301
rect 18162 4159 18196 4301
rect 18582 4159 18616 4301
rect 10392 3064 10426 3065
rect 10392 3030 10476 3064
rect 10812 3064 10846 3065
rect 10812 3030 10896 3064
rect 11232 3064 11266 3065
rect 11232 3030 11316 3064
rect 11652 3064 11686 3065
rect 11652 3030 11736 3064
rect 12072 3064 12106 3065
rect 12072 3030 12156 3064
rect 12492 3064 12526 3065
rect 12492 3030 12576 3064
rect 12912 3064 12946 3065
rect 12912 3030 12996 3064
rect 13332 3064 13366 3065
rect 13332 3030 13416 3064
rect 13752 3064 13786 3065
rect 13752 3030 13836 3064
rect 14172 3064 14206 3065
rect 14172 3030 14256 3064
rect 14592 3064 14626 3065
rect 14592 3030 14676 3064
rect 15012 3064 15046 3065
rect 15012 3030 15096 3064
rect 15432 3064 15466 3065
rect 15432 3030 15516 3064
rect 15852 3064 15886 3065
rect 15852 3030 15936 3064
rect 16272 3064 16306 3065
rect 16272 3030 16356 3064
rect 16692 3064 16726 3065
rect 16692 3030 16776 3064
rect 17112 3064 17146 3065
rect 17112 3030 17196 3064
rect 17532 3064 17566 3065
rect 17532 3030 17616 3064
rect 17952 3064 17986 3065
rect 17952 3030 18036 3064
rect 18372 3064 18406 3065
rect 18372 3030 18456 3064
rect 2726 -1540 2810 -1506
rect 3368 -1538 3452 -1504
rect 3368 -1539 3402 -1538
rect 3788 -1538 3872 -1504
rect 3788 -1539 3822 -1538
rect 4208 -1538 4292 -1504
rect 4208 -1539 4242 -1538
rect 4628 -1538 4712 -1504
rect 4628 -1539 4662 -1538
rect 2630 -2776 2664 -2633
rect 3578 -2776 3612 -2633
rect 3998 -2776 4032 -2633
rect 4418 -2666 4502 -2632
rect 4418 -2667 4452 -2666
rect 4838 -2666 4922 -2632
rect 4838 -2667 4872 -2666
rect 3788 -3894 3872 -3860
rect 3788 -3895 3822 -3894
rect 4208 -3894 4292 -3860
rect 4208 -3895 4242 -3894
rect 5542 -1538 5626 -1504
rect 5542 -1539 5576 -1538
rect 5962 -1538 6046 -1504
rect 5962 -1539 5996 -1538
rect 6382 -1538 6466 -1504
rect 6382 -1539 6416 -1538
rect 6802 -1538 6886 -1504
rect 6802 -1539 6836 -1538
rect 7222 -1538 7306 -1504
rect 7222 -1539 7256 -1538
rect 7642 -1538 7726 -1504
rect 7642 -1539 7676 -1538
rect 8062 -1538 8146 -1504
rect 8062 -1539 8096 -1538
rect 8482 -1538 8566 -1504
rect 8482 -1539 8516 -1538
rect 8902 -1538 8986 -1504
rect 8902 -1539 8936 -1538
rect 5752 -2775 5786 -2633
rect 6172 -2775 6206 -2633
rect 6592 -2775 6626 -2633
rect 7012 -2775 7046 -2633
rect 7432 -2775 7466 -2633
rect 7852 -2775 7886 -2633
rect 8272 -2775 8306 -2633
rect 8692 -2775 8726 -2633
rect 9112 -2775 9146 -2633
rect 5542 -3902 5626 -3868
rect 5542 -3903 5576 -3902
rect 5962 -3902 6046 -3868
rect 5962 -3903 5996 -3902
rect 6382 -3902 6466 -3868
rect 6382 -3903 6416 -3902
rect 6802 -3902 6886 -3868
rect 6802 -3903 6836 -3902
rect 7222 -3902 7306 -3868
rect 7222 -3903 7256 -3902
rect 7642 -3902 7726 -3868
rect 7642 -3903 7676 -3902
rect 8062 -3902 8146 -3868
rect 8062 -3903 8096 -3902
rect 8482 -3902 8566 -3868
rect 8482 -3903 8516 -3902
rect 8902 -3902 8986 -3868
rect 8902 -3903 8936 -3902
rect 5542 -5794 5626 -5760
rect 5542 -5795 5576 -5794
rect 5962 -5794 6046 -5760
rect 5962 -5795 5996 -5794
rect 6382 -5794 6466 -5760
rect 6382 -5800 6416 -5794
rect 6802 -5794 6886 -5760
rect 6802 -5800 6836 -5794
rect 7222 -5794 7306 -5760
rect 7222 -5800 7256 -5794
rect 7642 -5794 7726 -5760
rect 7642 -5800 7676 -5794
rect 8062 -5794 8146 -5760
rect 8062 -5800 8096 -5794
rect 8482 -5794 8566 -5760
rect 8482 -5800 8516 -5794
rect 8902 -5794 8986 -5760
rect 8902 -5800 8936 -5794
rect 5752 -6918 5836 -6884
rect 6172 -6884 6206 -6876
rect 6172 -6918 6256 -6884
rect 6592 -6884 6626 -6876
rect 6592 -6918 6676 -6884
rect 7012 -6884 7046 -6876
rect 7012 -6918 7096 -6884
rect 7432 -6884 7466 -6876
rect 7432 -6918 7516 -6884
rect 7852 -6884 7886 -6876
rect 7852 -6918 7936 -6884
rect 8272 -6884 8306 -6876
rect 8272 -6918 8356 -6884
rect 8692 -6884 8726 -6876
rect 8692 -6918 8776 -6884
rect 9112 -6884 9146 -6876
rect 9112 -6918 9196 -6884
<< locali >>
rect 10104 13268 10248 13302
rect 18728 13268 18858 13302
rect 10104 13146 10138 13268
rect 18824 13174 18858 13268
rect 10376 13086 10392 13120
rect 10476 13086 10492 13120
rect 10796 13086 10812 13120
rect 10896 13086 10912 13120
rect 11216 13086 11232 13120
rect 11316 13086 11332 13120
rect 11636 13086 11652 13120
rect 11736 13086 11752 13120
rect 12056 13086 12072 13120
rect 12156 13086 12172 13120
rect 12476 13086 12492 13120
rect 12576 13086 12592 13120
rect 12896 13086 12912 13120
rect 12996 13086 13012 13120
rect 13316 13086 13332 13120
rect 13416 13086 13432 13120
rect 13736 13086 13752 13120
rect 13836 13086 13852 13120
rect 14156 13086 14172 13120
rect 14256 13086 14272 13120
rect 14576 13086 14592 13120
rect 14676 13086 14692 13120
rect 14996 13086 15012 13120
rect 15096 13086 15112 13120
rect 15416 13086 15432 13120
rect 15516 13086 15532 13120
rect 15836 13086 15852 13120
rect 15936 13086 15952 13120
rect 16256 13086 16272 13120
rect 16356 13086 16372 13120
rect 16676 13086 16692 13120
rect 16776 13086 16792 13120
rect 17096 13086 17112 13120
rect 17196 13086 17212 13120
rect 17516 13086 17532 13120
rect 17616 13086 17632 13120
rect 17936 13086 17952 13120
rect 18036 13086 18052 13120
rect 18356 13086 18372 13120
rect 18456 13086 18472 13120
rect 10344 13036 10378 13052
rect 10344 12044 10378 12060
rect 10440 13036 10474 13052
rect 10440 12044 10474 12060
rect 10554 13036 10588 13052
rect 10554 12044 10588 12060
rect 10650 13036 10684 13052
rect 10650 12044 10684 12060
rect 10764 13036 10798 13052
rect 10764 12044 10798 12060
rect 10860 13036 10894 13052
rect 10860 12044 10894 12060
rect 10974 13036 11008 13052
rect 10974 12044 11008 12060
rect 11070 13036 11104 13052
rect 11070 12044 11104 12060
rect 11184 13036 11218 13052
rect 11184 12044 11218 12060
rect 11280 13036 11314 13052
rect 11280 12044 11314 12060
rect 11394 13036 11428 13052
rect 11394 12044 11428 12060
rect 11490 13036 11524 13052
rect 11490 12044 11524 12060
rect 11604 13036 11638 13052
rect 11604 12044 11638 12060
rect 11700 13036 11734 13052
rect 11700 12044 11734 12060
rect 11814 13036 11848 13052
rect 11814 12044 11848 12060
rect 11910 13036 11944 13052
rect 11910 12044 11944 12060
rect 12024 13036 12058 13052
rect 12024 12044 12058 12060
rect 12120 13036 12154 13052
rect 12120 12044 12154 12060
rect 12234 13036 12268 13052
rect 12234 12044 12268 12060
rect 12330 13036 12364 13052
rect 12330 12044 12364 12060
rect 12444 13036 12478 13052
rect 12444 12044 12478 12060
rect 12540 13036 12574 13052
rect 12540 12044 12574 12060
rect 12654 13036 12688 13052
rect 12654 12044 12688 12060
rect 12750 13036 12784 13052
rect 12750 12044 12784 12060
rect 12864 13036 12898 13052
rect 12864 12044 12898 12060
rect 12960 13036 12994 13052
rect 12960 12044 12994 12060
rect 13074 13036 13108 13052
rect 13074 12044 13108 12060
rect 13170 13036 13204 13052
rect 13170 12044 13204 12060
rect 13284 13036 13318 13052
rect 13284 12044 13318 12060
rect 13380 13036 13414 13052
rect 13380 12044 13414 12060
rect 13494 13036 13528 13052
rect 13494 12044 13528 12060
rect 13590 13036 13624 13052
rect 13590 12044 13624 12060
rect 13704 13036 13738 13052
rect 13704 12044 13738 12060
rect 13800 13036 13834 13052
rect 13800 12044 13834 12060
rect 13914 13036 13948 13052
rect 13914 12044 13948 12060
rect 14010 13036 14044 13052
rect 14010 12044 14044 12060
rect 14124 13036 14158 13052
rect 14124 12044 14158 12060
rect 14220 13036 14254 13052
rect 14220 12044 14254 12060
rect 14334 13036 14368 13052
rect 14334 12044 14368 12060
rect 14430 13036 14464 13052
rect 14430 12044 14464 12060
rect 14544 13036 14578 13052
rect 14544 12044 14578 12060
rect 14640 13036 14674 13052
rect 14640 12044 14674 12060
rect 14754 13036 14788 13052
rect 14754 12044 14788 12060
rect 14850 13036 14884 13052
rect 14850 12044 14884 12060
rect 14964 13036 14998 13052
rect 14964 12044 14998 12060
rect 15060 13036 15094 13052
rect 15060 12044 15094 12060
rect 15174 13036 15208 13052
rect 15174 12044 15208 12060
rect 15270 13036 15304 13052
rect 15270 12044 15304 12060
rect 15384 13036 15418 13052
rect 15384 12044 15418 12060
rect 15480 13036 15514 13052
rect 15480 12044 15514 12060
rect 15594 13036 15628 13052
rect 15594 12044 15628 12060
rect 15690 13036 15724 13052
rect 15690 12044 15724 12060
rect 15804 13036 15838 13052
rect 15804 12044 15838 12060
rect 15900 13036 15934 13052
rect 15900 12044 15934 12060
rect 16014 13036 16048 13052
rect 16014 12044 16048 12060
rect 16110 13036 16144 13052
rect 16110 12044 16144 12060
rect 16224 13036 16258 13052
rect 16224 12044 16258 12060
rect 16320 13036 16354 13052
rect 16320 12044 16354 12060
rect 16434 13036 16468 13052
rect 16434 12044 16468 12060
rect 16530 13036 16564 13052
rect 16530 12044 16564 12060
rect 16644 13036 16678 13052
rect 16644 12044 16678 12060
rect 16740 13036 16774 13052
rect 16740 12044 16774 12060
rect 16854 13036 16888 13052
rect 16854 12044 16888 12060
rect 16950 13036 16984 13052
rect 16950 12044 16984 12060
rect 17064 13036 17098 13052
rect 17064 12044 17098 12060
rect 17160 13036 17194 13052
rect 17160 12044 17194 12060
rect 17274 13036 17308 13052
rect 17274 12044 17308 12060
rect 17370 13036 17404 13052
rect 17370 12044 17404 12060
rect 17484 13036 17518 13052
rect 17484 12044 17518 12060
rect 17580 13036 17614 13052
rect 17580 12044 17614 12060
rect 17694 13036 17728 13052
rect 17694 12044 17728 12060
rect 17790 13036 17824 13052
rect 17790 12044 17824 12060
rect 17904 13036 17938 13052
rect 17904 12044 17938 12060
rect 18000 13036 18034 13052
rect 18000 12044 18034 12060
rect 18114 13036 18148 13052
rect 18114 12044 18148 12060
rect 18210 13036 18244 13052
rect 18210 12044 18244 12060
rect 18324 13036 18358 13052
rect 18324 12044 18358 12060
rect 18420 13036 18454 13052
rect 18420 12044 18454 12060
rect 18534 13036 18568 13052
rect 18534 12044 18568 12060
rect 18630 13036 18664 13052
rect 18630 12044 18664 12060
rect 10586 11976 10602 12010
rect 10586 11868 10602 11902
rect 10636 11976 10652 12010
rect 11006 11976 11022 12010
rect 10636 11868 10652 11902
rect 11006 11868 11022 11902
rect 11056 11976 11072 12010
rect 11426 11976 11442 12010
rect 11056 11868 11072 11902
rect 11426 11868 11442 11902
rect 11476 11976 11492 12010
rect 11846 11976 11862 12010
rect 11476 11868 11492 11902
rect 11846 11868 11862 11902
rect 11896 11976 11912 12010
rect 12266 11976 12282 12010
rect 11896 11868 11912 11902
rect 12266 11868 12282 11902
rect 12316 11976 12332 12010
rect 12686 11976 12702 12010
rect 12316 11868 12332 11902
rect 12686 11868 12702 11902
rect 12736 11976 12752 12010
rect 13106 11976 13122 12010
rect 12736 11868 12752 11902
rect 13106 11868 13122 11902
rect 13156 11976 13172 12010
rect 13526 11976 13542 12010
rect 13156 11868 13172 11902
rect 13526 11868 13542 11902
rect 13576 11976 13592 12010
rect 13946 11976 13962 12010
rect 13576 11868 13592 11902
rect 13946 11868 13962 11902
rect 13996 11976 14012 12010
rect 14366 11976 14382 12010
rect 13996 11868 14012 11902
rect 14366 11868 14382 11902
rect 14416 11976 14432 12010
rect 14786 11976 14802 12010
rect 14416 11868 14432 11902
rect 14786 11868 14802 11902
rect 14836 11976 14852 12010
rect 15206 11976 15222 12010
rect 14836 11868 14852 11902
rect 15206 11868 15222 11902
rect 15256 11976 15272 12010
rect 15626 11976 15642 12010
rect 15256 11868 15272 11902
rect 15626 11868 15642 11902
rect 15676 11976 15692 12010
rect 16046 11976 16062 12010
rect 15676 11868 15692 11902
rect 16046 11868 16062 11902
rect 16096 11976 16112 12010
rect 16466 11976 16482 12010
rect 16096 11868 16112 11902
rect 16466 11868 16482 11902
rect 16516 11976 16532 12010
rect 16886 11976 16902 12010
rect 16516 11868 16532 11902
rect 16886 11868 16902 11902
rect 16936 11976 16952 12010
rect 17306 11976 17322 12010
rect 16936 11868 16952 11902
rect 17306 11868 17322 11902
rect 17356 11976 17372 12010
rect 17726 11976 17742 12010
rect 17356 11868 17372 11902
rect 17726 11868 17742 11902
rect 17776 11976 17792 12010
rect 18146 11976 18162 12010
rect 17776 11868 17792 11902
rect 18146 11868 18162 11902
rect 18196 11976 18212 12010
rect 18566 11976 18582 12010
rect 18196 11868 18212 11902
rect 18566 11868 18582 11902
rect 18616 11976 18632 12010
rect 18616 11868 18632 11902
rect 10344 11818 10378 11834
rect 10344 10826 10378 10842
rect 10440 11818 10474 11834
rect 10440 10826 10474 10842
rect 10554 11818 10588 11834
rect 10554 10826 10588 10842
rect 10650 11818 10684 11834
rect 10650 10826 10684 10842
rect 10764 11818 10798 11834
rect 10764 10826 10798 10842
rect 10860 11818 10894 11834
rect 10860 10826 10894 10842
rect 10974 11818 11008 11834
rect 10974 10826 11008 10842
rect 11070 11818 11104 11834
rect 11070 10826 11104 10842
rect 11184 11818 11218 11834
rect 11184 10826 11218 10842
rect 11280 11818 11314 11834
rect 11280 10826 11314 10842
rect 11394 11818 11428 11834
rect 11394 10826 11428 10842
rect 11490 11818 11524 11834
rect 11490 10826 11524 10842
rect 11604 11818 11638 11834
rect 11604 10826 11638 10842
rect 11700 11818 11734 11834
rect 11700 10826 11734 10842
rect 11814 11818 11848 11834
rect 11814 10826 11848 10842
rect 11910 11818 11944 11834
rect 11910 10826 11944 10842
rect 12024 11818 12058 11834
rect 12024 10826 12058 10842
rect 12120 11818 12154 11834
rect 12120 10826 12154 10842
rect 12234 11818 12268 11834
rect 12234 10826 12268 10842
rect 12330 11818 12364 11834
rect 12330 10826 12364 10842
rect 12444 11818 12478 11834
rect 12444 10826 12478 10842
rect 12540 11818 12574 11834
rect 12540 10826 12574 10842
rect 12654 11818 12688 11834
rect 12654 10826 12688 10842
rect 12750 11818 12784 11834
rect 12750 10826 12784 10842
rect 12864 11818 12898 11834
rect 12864 10826 12898 10842
rect 12960 11818 12994 11834
rect 12960 10826 12994 10842
rect 13074 11818 13108 11834
rect 13074 10826 13108 10842
rect 13170 11818 13204 11834
rect 13170 10826 13204 10842
rect 13284 11818 13318 11834
rect 13284 10826 13318 10842
rect 13380 11818 13414 11834
rect 13380 10826 13414 10842
rect 13494 11818 13528 11834
rect 13494 10826 13528 10842
rect 13590 11818 13624 11834
rect 13590 10826 13624 10842
rect 13704 11818 13738 11834
rect 13704 10826 13738 10842
rect 13800 11818 13834 11834
rect 13800 10826 13834 10842
rect 13914 11818 13948 11834
rect 13914 10826 13948 10842
rect 14010 11818 14044 11834
rect 14010 10826 14044 10842
rect 14124 11818 14158 11834
rect 14124 10826 14158 10842
rect 14220 11818 14254 11834
rect 14220 10826 14254 10842
rect 14334 11818 14368 11834
rect 14334 10826 14368 10842
rect 14430 11818 14464 11834
rect 14430 10826 14464 10842
rect 14544 11818 14578 11834
rect 14544 10826 14578 10842
rect 14640 11818 14674 11834
rect 14640 10826 14674 10842
rect 14754 11818 14788 11834
rect 14754 10826 14788 10842
rect 14850 11818 14884 11834
rect 14850 10826 14884 10842
rect 14964 11818 14998 11834
rect 14964 10826 14998 10842
rect 15060 11818 15094 11834
rect 15060 10826 15094 10842
rect 15174 11818 15208 11834
rect 15174 10826 15208 10842
rect 15270 11818 15304 11834
rect 15270 10826 15304 10842
rect 15384 11818 15418 11834
rect 15384 10826 15418 10842
rect 15480 11818 15514 11834
rect 15480 10826 15514 10842
rect 15594 11818 15628 11834
rect 15594 10826 15628 10842
rect 15690 11818 15724 11834
rect 15690 10826 15724 10842
rect 15804 11818 15838 11834
rect 15804 10826 15838 10842
rect 15900 11818 15934 11834
rect 15900 10826 15934 10842
rect 16014 11818 16048 11834
rect 16014 10826 16048 10842
rect 16110 11818 16144 11834
rect 16110 10826 16144 10842
rect 16224 11818 16258 11834
rect 16224 10826 16258 10842
rect 16320 11818 16354 11834
rect 16320 10826 16354 10842
rect 16434 11818 16468 11834
rect 16434 10826 16468 10842
rect 16530 11818 16564 11834
rect 16530 10826 16564 10842
rect 16644 11818 16678 11834
rect 16644 10826 16678 10842
rect 16740 11818 16774 11834
rect 16740 10826 16774 10842
rect 16854 11818 16888 11834
rect 16854 10826 16888 10842
rect 16950 11818 16984 11834
rect 16950 10826 16984 10842
rect 17064 11818 17098 11834
rect 17064 10826 17098 10842
rect 17160 11818 17194 11834
rect 17160 10826 17194 10842
rect 17274 11818 17308 11834
rect 17274 10826 17308 10842
rect 17370 11818 17404 11834
rect 17370 10826 17404 10842
rect 17484 11818 17518 11834
rect 17484 10826 17518 10842
rect 17580 11818 17614 11834
rect 17580 10826 17614 10842
rect 17694 11818 17728 11834
rect 17694 10826 17728 10842
rect 17790 11818 17824 11834
rect 17790 10826 17824 10842
rect 17904 11818 17938 11834
rect 17904 10826 17938 10842
rect 18000 11818 18034 11834
rect 18000 10826 18034 10842
rect 18114 11818 18148 11834
rect 18114 10826 18148 10842
rect 18210 11818 18244 11834
rect 18210 10826 18244 10842
rect 18324 11818 18358 11834
rect 18324 10826 18358 10842
rect 18420 11818 18454 11834
rect 18420 10826 18454 10842
rect 18534 11818 18568 11834
rect 18534 10826 18568 10842
rect 18630 11818 18664 11834
rect 18630 10826 18664 10842
rect 10104 10626 10138 10774
rect 10376 10758 10392 10792
rect 10476 10758 10492 10792
rect 10796 10758 10812 10792
rect 10896 10758 10912 10792
rect 11216 10758 11232 10792
rect 11316 10758 11332 10792
rect 11636 10758 11652 10792
rect 11736 10758 11752 10792
rect 12056 10758 12072 10792
rect 12156 10758 12172 10792
rect 12476 10758 12492 10792
rect 12576 10758 12592 10792
rect 12896 10758 12912 10792
rect 12996 10758 13012 10792
rect 13316 10758 13332 10792
rect 13416 10758 13432 10792
rect 13736 10758 13752 10792
rect 13836 10758 13852 10792
rect 14156 10758 14172 10792
rect 14256 10758 14272 10792
rect 14576 10758 14592 10792
rect 14676 10758 14692 10792
rect 14996 10758 15012 10792
rect 15096 10758 15112 10792
rect 15416 10758 15432 10792
rect 15516 10758 15532 10792
rect 15836 10758 15852 10792
rect 15936 10758 15952 10792
rect 16256 10758 16272 10792
rect 16356 10758 16372 10792
rect 16676 10758 16692 10792
rect 16776 10758 16792 10792
rect 17096 10758 17112 10792
rect 17196 10758 17212 10792
rect 17516 10758 17532 10792
rect 17616 10758 17632 10792
rect 17936 10758 17952 10792
rect 18036 10758 18052 10792
rect 18356 10758 18372 10792
rect 18456 10758 18472 10792
rect 18824 10626 18858 10762
rect 10104 10592 10260 10626
rect 18630 10592 18858 10626
rect 10132 7996 10358 8030
rect 18680 7996 18796 8030
rect 10132 7844 10166 7996
rect 10376 7901 10427 7906
rect 10796 7901 10847 7906
rect 11216 7901 11267 7906
rect 11636 7901 11687 7906
rect 12056 7901 12107 7906
rect 12476 7901 12527 7906
rect 12896 7901 12947 7906
rect 13316 7901 13367 7906
rect 13736 7901 13787 7906
rect 14156 7901 14207 7906
rect 14576 7901 14627 7906
rect 14996 7901 15047 7906
rect 15416 7901 15467 7906
rect 15836 7901 15887 7906
rect 16256 7901 16307 7906
rect 16676 7901 16727 7906
rect 17096 7901 17147 7906
rect 17516 7901 17567 7906
rect 17936 7901 17987 7906
rect 18356 7901 18407 7906
rect 10376 7866 10392 7901
rect 10426 7900 10442 7901
rect 10476 7866 10492 7900
rect 10796 7866 10812 7901
rect 10846 7900 10862 7901
rect 10896 7866 10912 7900
rect 11216 7866 11232 7901
rect 11266 7900 11282 7901
rect 11316 7866 11332 7900
rect 11636 7866 11652 7901
rect 11686 7900 11702 7901
rect 11736 7866 11752 7900
rect 12056 7866 12072 7901
rect 12106 7900 12122 7901
rect 12156 7866 12172 7900
rect 12476 7866 12492 7901
rect 12526 7900 12542 7901
rect 12576 7866 12592 7900
rect 12896 7866 12912 7901
rect 12946 7900 12962 7901
rect 12996 7866 13012 7900
rect 13316 7866 13332 7901
rect 13366 7900 13382 7901
rect 13416 7866 13432 7900
rect 13736 7866 13752 7901
rect 13786 7900 13802 7901
rect 13836 7866 13852 7900
rect 14156 7866 14172 7901
rect 14206 7900 14222 7901
rect 14256 7866 14272 7900
rect 14576 7866 14592 7901
rect 14626 7900 14642 7901
rect 14676 7866 14692 7900
rect 14996 7866 15012 7901
rect 15046 7900 15062 7901
rect 15096 7866 15112 7900
rect 15416 7866 15432 7901
rect 15466 7900 15482 7901
rect 15516 7866 15532 7900
rect 15836 7866 15852 7901
rect 15886 7900 15902 7901
rect 15936 7866 15952 7900
rect 16256 7866 16272 7901
rect 16306 7900 16322 7901
rect 16356 7866 16372 7900
rect 16676 7866 16692 7901
rect 16726 7900 16742 7901
rect 16776 7866 16792 7900
rect 17096 7866 17112 7901
rect 17146 7900 17162 7901
rect 17196 7866 17212 7900
rect 17516 7866 17532 7901
rect 17566 7900 17582 7901
rect 17616 7866 17632 7900
rect 17936 7866 17952 7901
rect 17986 7900 18002 7901
rect 18036 7866 18052 7900
rect 18356 7866 18372 7901
rect 18406 7900 18422 7901
rect 18456 7866 18472 7900
rect 10376 7858 10427 7866
rect 10796 7858 10847 7866
rect 11216 7858 11267 7866
rect 11636 7858 11687 7866
rect 12056 7858 12107 7866
rect 12476 7858 12527 7866
rect 12896 7858 12947 7866
rect 13316 7858 13367 7866
rect 13736 7858 13787 7866
rect 14156 7858 14207 7866
rect 14576 7858 14627 7866
rect 14996 7858 15047 7866
rect 15416 7858 15467 7866
rect 15836 7858 15887 7866
rect 16256 7858 16307 7866
rect 16676 7858 16727 7866
rect 17096 7858 17147 7866
rect 17516 7858 17567 7866
rect 17936 7858 17987 7866
rect 18356 7858 18407 7866
rect 5348 7096 5480 7130
rect 9204 7096 9310 7130
rect 5348 6980 5382 7096
rect 5736 7045 5787 7050
rect 6156 7045 6207 7050
rect 6576 7045 6627 7050
rect 6996 7045 7047 7050
rect 7416 7045 7467 7050
rect 7836 7045 7887 7050
rect 8256 7045 8307 7050
rect 8676 7045 8727 7050
rect 9096 7045 9147 7050
rect 5736 7044 5802 7045
rect 6156 7044 6222 7045
rect 6576 7044 6642 7045
rect 6996 7044 7062 7045
rect 7416 7044 7482 7045
rect 7836 7044 7902 7045
rect 8256 7044 8322 7045
rect 8676 7044 8742 7045
rect 9096 7044 9162 7045
rect 5736 7010 5752 7044
rect 5836 7010 5852 7044
rect 5736 7002 5787 7010
rect 6156 7002 6172 7044
rect 6256 7010 6272 7044
rect 6206 7002 6222 7010
rect 6576 7002 6592 7044
rect 6676 7010 6692 7044
rect 6626 7002 6642 7010
rect 6996 7002 7012 7044
rect 7096 7010 7112 7044
rect 7046 7002 7062 7010
rect 7416 7002 7432 7044
rect 7516 7010 7532 7044
rect 7466 7002 7482 7010
rect 7836 7002 7852 7044
rect 7936 7010 7952 7044
rect 7886 7002 7902 7010
rect 8256 7002 8272 7044
rect 8356 7010 8372 7044
rect 8306 7002 8322 7010
rect 8676 7002 8692 7044
rect 8776 7010 8792 7044
rect 8726 7002 8742 7010
rect 9096 7002 9112 7044
rect 9196 7010 9212 7044
rect 9146 7002 9162 7010
rect 9276 7004 9310 7096
rect 5494 6952 5528 6968
rect 5494 5960 5528 5976
rect 5590 6952 5624 6968
rect 5590 5960 5624 5976
rect 5704 6952 5738 6968
rect 5704 5960 5738 5976
rect 5800 6952 5834 6968
rect 5800 5960 5834 5976
rect 5914 6952 5948 6968
rect 5914 5960 5948 5976
rect 6010 6952 6044 6968
rect 6010 5960 6044 5976
rect 6124 6952 6158 6968
rect 6124 5960 6158 5976
rect 6220 6952 6254 6968
rect 6220 5960 6254 5976
rect 6334 6952 6368 6968
rect 6334 5960 6368 5976
rect 6430 6952 6464 6968
rect 6430 5960 6464 5976
rect 6544 6952 6578 6968
rect 6544 5960 6578 5976
rect 6640 6952 6674 6968
rect 6640 5960 6674 5976
rect 6754 6952 6788 6968
rect 6754 5960 6788 5976
rect 6850 6952 6884 6968
rect 6850 5960 6884 5976
rect 6964 6952 6998 6968
rect 6964 5960 6998 5976
rect 7060 6952 7094 6968
rect 7060 5960 7094 5976
rect 7174 6952 7208 6968
rect 7174 5960 7208 5976
rect 7270 6952 7304 6968
rect 7270 5960 7304 5976
rect 7384 6952 7418 6968
rect 7384 5960 7418 5976
rect 7480 6952 7514 6968
rect 7480 5960 7514 5976
rect 7594 6952 7628 6968
rect 7594 5960 7628 5976
rect 7690 6952 7724 6968
rect 7690 5960 7724 5976
rect 7804 6952 7838 6968
rect 7804 5960 7838 5976
rect 7900 6952 7934 6968
rect 7900 5960 7934 5976
rect 8014 6952 8048 6968
rect 8014 5960 8048 5976
rect 8110 6952 8144 6968
rect 8110 5960 8144 5976
rect 8224 6952 8258 6968
rect 8224 5960 8258 5976
rect 8320 6952 8354 6968
rect 8320 5960 8354 5976
rect 8434 6952 8468 6968
rect 8434 5960 8468 5976
rect 8530 6952 8564 6968
rect 8530 5960 8564 5976
rect 8644 6952 8678 6968
rect 8644 5960 8678 5976
rect 8740 6952 8774 6968
rect 8740 5960 8774 5976
rect 8854 6952 8888 6968
rect 8854 5960 8888 5976
rect 8950 6952 8984 6968
rect 8950 5960 8984 5976
rect 9064 6952 9098 6968
rect 9064 5960 9098 5976
rect 9160 6952 9194 6968
rect 9160 5960 9194 5976
rect 5348 5842 5382 5960
rect 5526 5921 5577 5926
rect 5946 5921 5997 5926
rect 5526 5886 5542 5921
rect 5576 5920 5592 5921
rect 5626 5886 5642 5920
rect 5946 5886 5962 5921
rect 5996 5920 6012 5921
rect 6046 5886 6062 5920
rect 6366 5886 6382 5926
rect 6416 5920 6432 5926
rect 6466 5886 6482 5920
rect 6786 5886 6802 5926
rect 6836 5920 6852 5926
rect 6886 5886 6902 5920
rect 7206 5886 7222 5926
rect 7256 5920 7272 5926
rect 7306 5886 7322 5920
rect 7626 5886 7642 5926
rect 7676 5920 7692 5926
rect 7726 5886 7742 5920
rect 8046 5886 8062 5926
rect 8096 5920 8112 5926
rect 8146 5886 8162 5920
rect 8466 5886 8482 5926
rect 8516 5920 8532 5926
rect 8566 5886 8582 5920
rect 8886 5886 8902 5926
rect 8936 5920 8952 5926
rect 8986 5886 9002 5920
rect 5526 5878 5577 5886
rect 5946 5878 5997 5886
rect 6366 5878 6417 5886
rect 6786 5878 6837 5886
rect 7206 5878 7257 5886
rect 7626 5878 7677 5886
rect 8046 5878 8097 5886
rect 8466 5878 8517 5886
rect 8886 5878 8937 5886
rect 9276 5842 9310 5962
rect 5348 5808 5440 5842
rect 9160 5808 9310 5842
rect 5384 5536 5514 5570
rect 9216 5536 9332 5570
rect 2586 5328 2620 5344
rect 2586 4336 2620 4352
rect 2674 5328 2708 5344
rect 3064 5234 3160 5516
rect 5384 5494 5418 5536
rect 3772 5421 3823 5426
rect 4192 5421 4243 5426
rect 3772 5386 3788 5421
rect 3822 5420 3838 5421
rect 3872 5386 3888 5420
rect 4192 5386 4208 5421
rect 4242 5420 4258 5421
rect 4292 5386 4308 5420
rect 3772 5378 3823 5386
rect 4192 5378 4243 5386
rect 3530 5328 3564 5344
rect 3000 5218 3206 5234
rect 3000 4510 3206 4526
rect 2674 4336 2708 4352
rect 3530 4336 3564 4352
rect 3626 5328 3660 5344
rect 3626 4336 3660 4352
rect 3740 5328 3774 5344
rect 3740 4336 3774 4352
rect 3836 5328 3870 5344
rect 3836 4336 3870 4352
rect 3950 5328 3984 5344
rect 3950 4336 3984 4352
rect 4046 5328 4080 5344
rect 4046 4336 4080 4352
rect 4160 5328 4194 5344
rect 4160 4336 4194 4352
rect 4256 5328 4290 5344
rect 4256 4336 4290 4352
rect 2614 4268 2630 4302
rect 2614 4159 2630 4193
rect 2664 4268 2680 4302
rect 3562 4268 3578 4302
rect 2664 4159 2680 4193
rect 3562 4159 3578 4193
rect 3612 4268 3628 4302
rect 3982 4268 3998 4302
rect 3612 4159 3628 4193
rect 3982 4159 3998 4193
rect 4032 4268 4048 4302
rect 4402 4193 4453 4198
rect 4822 4193 4873 4198
rect 4032 4159 4048 4193
rect 4402 4158 4418 4193
rect 4452 4192 4468 4193
rect 4502 4158 4518 4192
rect 4822 4158 4838 4193
rect 4872 4192 4888 4193
rect 4922 4158 4938 4192
rect 4402 4150 4453 4158
rect 4822 4150 4873 4158
rect 2582 4100 2616 4116
rect 2582 3108 2616 3124
rect 2678 4100 2712 4116
rect 2678 3108 2712 3124
rect 2774 4100 2808 4116
rect 3320 4100 3354 4116
rect 2924 4016 3130 4032
rect 2924 3308 3130 3324
rect 2774 3108 2808 3124
rect 2710 3066 2761 3072
rect 2710 3032 2726 3066
rect 2810 3032 2826 3066
rect 2710 3024 2761 3032
rect 3010 2838 3104 3308
rect 3320 3108 3354 3124
rect 3416 4100 3450 4116
rect 3416 3108 3450 3124
rect 3530 4100 3564 4116
rect 3530 3108 3564 3124
rect 3626 4100 3660 4116
rect 3626 3108 3660 3124
rect 3740 4100 3774 4116
rect 3740 3108 3774 3124
rect 3836 4100 3870 4116
rect 3836 3108 3870 3124
rect 3950 4100 3984 4116
rect 3950 3108 3984 3124
rect 4046 4100 4080 4116
rect 4046 3108 4080 3124
rect 4160 4100 4194 4116
rect 4160 3108 4194 3124
rect 4256 4100 4290 4116
rect 4256 3108 4290 3124
rect 4370 4100 4404 4116
rect 4370 3108 4404 3124
rect 4466 4100 4500 4116
rect 4466 3108 4500 3124
rect 4580 4100 4614 4116
rect 4580 3108 4614 3124
rect 4676 4100 4710 4116
rect 4676 3108 4710 3124
rect 4790 4100 4824 4116
rect 4790 3108 4824 3124
rect 4886 4100 4920 4116
rect 4886 3108 4920 3124
rect 3352 3065 3403 3070
rect 3772 3065 3823 3070
rect 4192 3065 4243 3070
rect 4612 3065 4663 3070
rect 3352 3030 3368 3065
rect 3402 3064 3418 3065
rect 3452 3030 3468 3064
rect 3772 3030 3788 3065
rect 3822 3064 3838 3065
rect 3872 3030 3888 3064
rect 4192 3030 4208 3065
rect 4242 3064 4258 3065
rect 4292 3030 4308 3064
rect 4612 3030 4628 3065
rect 4662 3064 4678 3065
rect 4712 3030 4728 3064
rect 3352 3022 3403 3030
rect 3772 3022 3823 3030
rect 4192 3022 4243 3030
rect 4612 3022 4663 3030
rect 5526 5429 5577 5434
rect 5946 5429 5997 5434
rect 6366 5429 6417 5434
rect 6786 5429 6837 5434
rect 7206 5429 7257 5434
rect 7626 5429 7677 5434
rect 8046 5429 8097 5434
rect 8466 5429 8517 5434
rect 8886 5429 8937 5434
rect 5526 5394 5542 5429
rect 5576 5428 5592 5429
rect 5626 5394 5642 5428
rect 5946 5394 5962 5429
rect 5996 5428 6012 5429
rect 6046 5394 6062 5428
rect 6366 5394 6382 5429
rect 6416 5428 6432 5429
rect 6466 5394 6482 5428
rect 6786 5394 6802 5429
rect 6836 5428 6852 5429
rect 6886 5394 6902 5428
rect 7206 5394 7222 5429
rect 7256 5428 7272 5429
rect 7306 5394 7322 5428
rect 7626 5394 7642 5429
rect 7676 5428 7692 5429
rect 7726 5394 7742 5428
rect 8046 5394 8062 5429
rect 8096 5428 8112 5429
rect 8146 5394 8162 5428
rect 8466 5394 8482 5429
rect 8516 5428 8532 5429
rect 8566 5394 8582 5428
rect 8886 5394 8902 5429
rect 8936 5428 8952 5429
rect 8986 5394 9002 5428
rect 5526 5386 5577 5394
rect 5946 5386 5997 5394
rect 6366 5386 6417 5394
rect 6786 5386 6837 5394
rect 7206 5386 7257 5394
rect 7626 5386 7677 5394
rect 8046 5386 8097 5394
rect 8466 5386 8517 5394
rect 8886 5386 8937 5394
rect 9298 5352 9332 5536
rect 5494 5336 5528 5352
rect 5494 4344 5528 4360
rect 5590 5336 5624 5352
rect 5590 4344 5624 4360
rect 5704 5336 5738 5352
rect 5704 4344 5738 4360
rect 5800 5336 5834 5352
rect 5800 4344 5834 4360
rect 5914 5336 5948 5352
rect 5914 4344 5948 4360
rect 6010 5336 6044 5352
rect 6010 4344 6044 4360
rect 6124 5336 6158 5352
rect 6124 4344 6158 4360
rect 6220 5336 6254 5352
rect 6220 4344 6254 4360
rect 6334 5336 6368 5352
rect 6334 4344 6368 4360
rect 6430 5336 6464 5352
rect 6430 4344 6464 4360
rect 6544 5336 6578 5352
rect 6544 4344 6578 4360
rect 6640 5336 6674 5352
rect 6640 4344 6674 4360
rect 6754 5336 6788 5352
rect 6754 4344 6788 4360
rect 6850 5336 6884 5352
rect 6850 4344 6884 4360
rect 6964 5336 6998 5352
rect 6964 4344 6998 4360
rect 7060 5336 7094 5352
rect 7060 4344 7094 4360
rect 7174 5336 7208 5352
rect 7174 4344 7208 4360
rect 7270 5336 7304 5352
rect 7270 4344 7304 4360
rect 7384 5336 7418 5352
rect 7384 4344 7418 4360
rect 7480 5336 7514 5352
rect 7480 4344 7514 4360
rect 7594 5336 7628 5352
rect 7594 4344 7628 4360
rect 7690 5336 7724 5352
rect 7690 4344 7724 4360
rect 7804 5336 7838 5352
rect 7804 4344 7838 4360
rect 7900 5336 7934 5352
rect 7900 4344 7934 4360
rect 8014 5336 8048 5352
rect 8014 4344 8048 4360
rect 8110 5336 8144 5352
rect 8110 4344 8144 4360
rect 8224 5336 8258 5352
rect 8224 4344 8258 4360
rect 8320 5336 8354 5352
rect 8320 4344 8354 4360
rect 8434 5336 8468 5352
rect 8434 4344 8468 4360
rect 8530 5336 8564 5352
rect 8530 4344 8564 4360
rect 8644 5336 8678 5352
rect 8644 4344 8678 4360
rect 8740 5336 8774 5352
rect 8740 4344 8774 4360
rect 8854 5336 8888 5352
rect 8854 4344 8888 4360
rect 8950 5336 8984 5352
rect 8950 4344 8984 4360
rect 9064 5336 9098 5352
rect 9064 4344 9098 4360
rect 9160 5336 9194 5352
rect 9160 4344 9194 4360
rect 5736 4267 5752 4301
rect 5736 4159 5752 4193
rect 5786 4267 5802 4301
rect 6156 4267 6172 4301
rect 5786 4159 5802 4193
rect 6156 4159 6172 4193
rect 6206 4267 6222 4301
rect 6576 4267 6592 4301
rect 6206 4159 6222 4193
rect 6576 4159 6592 4193
rect 6626 4267 6642 4301
rect 6996 4267 7012 4301
rect 6626 4159 6642 4193
rect 6996 4159 7012 4193
rect 7046 4267 7062 4301
rect 7416 4267 7432 4301
rect 7046 4159 7062 4193
rect 7416 4159 7432 4193
rect 7466 4267 7482 4301
rect 7836 4267 7852 4301
rect 7466 4159 7482 4193
rect 7836 4159 7852 4193
rect 7886 4267 7902 4301
rect 8256 4267 8272 4301
rect 7886 4159 7902 4193
rect 8256 4159 8272 4193
rect 8306 4267 8322 4301
rect 8676 4267 8692 4301
rect 8306 4159 8322 4193
rect 8676 4159 8692 4193
rect 8726 4267 8742 4301
rect 9096 4267 9112 4301
rect 8726 4159 8742 4193
rect 9096 4159 9112 4193
rect 9146 4267 9162 4301
rect 9146 4159 9162 4193
rect 5494 4100 5528 4116
rect 5494 3108 5528 3124
rect 5590 4100 5624 4116
rect 5590 3108 5624 3124
rect 5704 4100 5738 4116
rect 5704 3108 5738 3124
rect 5800 4100 5834 4116
rect 5800 3108 5834 3124
rect 5914 4100 5948 4116
rect 5914 3108 5948 3124
rect 6010 4100 6044 4116
rect 6010 3108 6044 3124
rect 6124 4100 6158 4116
rect 6124 3108 6158 3124
rect 6220 4100 6254 4116
rect 6220 3108 6254 3124
rect 6334 4100 6368 4116
rect 6334 3108 6368 3124
rect 6430 4100 6464 4116
rect 6430 3108 6464 3124
rect 6544 4100 6578 4116
rect 6544 3108 6578 3124
rect 6640 4100 6674 4116
rect 6640 3108 6674 3124
rect 6754 4100 6788 4116
rect 6754 3108 6788 3124
rect 6850 4100 6884 4116
rect 6850 3108 6884 3124
rect 6964 4100 6998 4116
rect 6964 3108 6998 3124
rect 7060 4100 7094 4116
rect 7060 3108 7094 3124
rect 7174 4100 7208 4116
rect 7174 3108 7208 3124
rect 7270 4100 7304 4116
rect 7270 3108 7304 3124
rect 7384 4100 7418 4116
rect 7384 3108 7418 3124
rect 7480 4100 7514 4116
rect 7480 3108 7514 3124
rect 7594 4100 7628 4116
rect 7594 3108 7628 3124
rect 7690 4100 7724 4116
rect 7690 3108 7724 3124
rect 7804 4100 7838 4116
rect 7804 3108 7838 3124
rect 7900 4100 7934 4116
rect 7900 3108 7934 3124
rect 8014 4100 8048 4116
rect 8014 3108 8048 3124
rect 8110 4100 8144 4116
rect 8110 3108 8144 3124
rect 8224 4100 8258 4116
rect 8224 3108 8258 3124
rect 8320 4100 8354 4116
rect 8320 3108 8354 3124
rect 8434 4100 8468 4116
rect 8434 3108 8468 3124
rect 8530 4100 8564 4116
rect 8530 3108 8564 3124
rect 8644 4100 8678 4116
rect 8644 3108 8678 3124
rect 8740 4100 8774 4116
rect 8740 3108 8774 3124
rect 8854 4100 8888 4116
rect 8854 3108 8888 3124
rect 8950 4100 8984 4116
rect 8950 3108 8984 3124
rect 9064 4100 9098 4116
rect 9064 3108 9098 3124
rect 9160 4100 9194 4116
rect 9160 3108 9194 3124
rect 5384 2970 5418 3026
rect 5526 3065 5577 3070
rect 5946 3065 5997 3070
rect 6366 3065 6417 3070
rect 6786 3065 6837 3070
rect 7206 3065 7257 3070
rect 7626 3065 7677 3070
rect 8046 3065 8097 3070
rect 8466 3065 8517 3070
rect 8886 3065 8937 3070
rect 5526 3030 5542 3065
rect 5576 3064 5592 3065
rect 5626 3030 5642 3064
rect 5946 3030 5962 3065
rect 5996 3064 6012 3065
rect 6046 3030 6062 3064
rect 6366 3030 6382 3065
rect 6416 3064 6432 3065
rect 6466 3030 6482 3064
rect 6786 3030 6802 3065
rect 6836 3064 6852 3065
rect 6886 3030 6902 3064
rect 7206 3030 7222 3065
rect 7256 3064 7272 3065
rect 7306 3030 7322 3064
rect 7626 3030 7642 3065
rect 7676 3064 7692 3065
rect 7726 3030 7742 3064
rect 8046 3030 8062 3065
rect 8096 3064 8112 3065
rect 8146 3030 8162 3064
rect 8466 3030 8482 3065
rect 8516 3064 8532 3065
rect 8566 3030 8582 3064
rect 8886 3030 8902 3065
rect 8936 3064 8952 3065
rect 8986 3030 9002 3064
rect 5526 3022 5577 3030
rect 5946 3022 5997 3030
rect 6366 3022 6417 3030
rect 6786 3022 6837 3030
rect 7206 3022 7257 3030
rect 7626 3022 7677 3030
rect 8046 3022 8097 3030
rect 8466 3022 8517 3030
rect 8886 3022 8937 3030
rect 9298 2938 9332 3064
rect 5466 2904 5486 2938
rect 9258 2904 9332 2938
rect 18762 7826 18796 7996
rect 10344 7808 10378 7824
rect 10344 6816 10378 6832
rect 10440 7808 10474 7824
rect 10440 6816 10474 6832
rect 10554 7808 10588 7824
rect 10554 6816 10588 6832
rect 10650 7808 10684 7824
rect 10650 6816 10684 6832
rect 10764 7808 10798 7824
rect 10764 6816 10798 6832
rect 10860 7808 10894 7824
rect 10860 6816 10894 6832
rect 10974 7808 11008 7824
rect 10974 6816 11008 6832
rect 11070 7808 11104 7824
rect 11070 6816 11104 6832
rect 11184 7808 11218 7824
rect 11184 6816 11218 6832
rect 11280 7808 11314 7824
rect 11280 6816 11314 6832
rect 11394 7808 11428 7824
rect 11394 6816 11428 6832
rect 11490 7808 11524 7824
rect 11490 6816 11524 6832
rect 11604 7808 11638 7824
rect 11604 6816 11638 6832
rect 11700 7808 11734 7824
rect 11700 6816 11734 6832
rect 11814 7808 11848 7824
rect 11814 6816 11848 6832
rect 11910 7808 11944 7824
rect 11910 6816 11944 6832
rect 12024 7808 12058 7824
rect 12024 6816 12058 6832
rect 12120 7808 12154 7824
rect 12120 6816 12154 6832
rect 12234 7808 12268 7824
rect 12234 6816 12268 6832
rect 12330 7808 12364 7824
rect 12330 6816 12364 6832
rect 12444 7808 12478 7824
rect 12444 6816 12478 6832
rect 12540 7808 12574 7824
rect 12540 6816 12574 6832
rect 12654 7808 12688 7824
rect 12654 6816 12688 6832
rect 12750 7808 12784 7824
rect 12750 6816 12784 6832
rect 12864 7808 12898 7824
rect 12864 6816 12898 6832
rect 12960 7808 12994 7824
rect 12960 6816 12994 6832
rect 13074 7808 13108 7824
rect 13074 6816 13108 6832
rect 13170 7808 13204 7824
rect 13170 6816 13204 6832
rect 13284 7808 13318 7824
rect 13284 6816 13318 6832
rect 13380 7808 13414 7824
rect 13380 6816 13414 6832
rect 13494 7808 13528 7824
rect 13494 6816 13528 6832
rect 13590 7808 13624 7824
rect 13590 6816 13624 6832
rect 13704 7808 13738 7824
rect 13704 6816 13738 6832
rect 13800 7808 13834 7824
rect 13800 6816 13834 6832
rect 13914 7808 13948 7824
rect 13914 6816 13948 6832
rect 14010 7808 14044 7824
rect 14010 6816 14044 6832
rect 14124 7808 14158 7824
rect 14124 6816 14158 6832
rect 14220 7808 14254 7824
rect 14220 6816 14254 6832
rect 14334 7808 14368 7824
rect 14334 6816 14368 6832
rect 14430 7808 14464 7824
rect 14430 6816 14464 6832
rect 14544 7808 14578 7824
rect 14544 6816 14578 6832
rect 14640 7808 14674 7824
rect 14640 6816 14674 6832
rect 14754 7808 14788 7824
rect 14754 6816 14788 6832
rect 14850 7808 14884 7824
rect 14850 6816 14884 6832
rect 14964 7808 14998 7824
rect 14964 6816 14998 6832
rect 15060 7808 15094 7824
rect 15060 6816 15094 6832
rect 15174 7808 15208 7824
rect 15174 6816 15208 6832
rect 15270 7808 15304 7824
rect 15270 6816 15304 6832
rect 15384 7808 15418 7824
rect 15384 6816 15418 6832
rect 15480 7808 15514 7824
rect 15480 6816 15514 6832
rect 15594 7808 15628 7824
rect 15594 6816 15628 6832
rect 15690 7808 15724 7824
rect 15690 6816 15724 6832
rect 15804 7808 15838 7824
rect 15804 6816 15838 6832
rect 15900 7808 15934 7824
rect 15900 6816 15934 6832
rect 16014 7808 16048 7824
rect 16014 6816 16048 6832
rect 16110 7808 16144 7824
rect 16110 6816 16144 6832
rect 16224 7808 16258 7824
rect 16224 6816 16258 6832
rect 16320 7808 16354 7824
rect 16320 6816 16354 6832
rect 16434 7808 16468 7824
rect 16434 6816 16468 6832
rect 16530 7808 16564 7824
rect 16530 6816 16564 6832
rect 16644 7808 16678 7824
rect 16644 6816 16678 6832
rect 16740 7808 16774 7824
rect 16740 6816 16774 6832
rect 16854 7808 16888 7824
rect 16854 6816 16888 6832
rect 16950 7808 16984 7824
rect 16950 6816 16984 6832
rect 17064 7808 17098 7824
rect 17064 6816 17098 6832
rect 17160 7808 17194 7824
rect 17160 6816 17194 6832
rect 17274 7808 17308 7824
rect 17274 6816 17308 6832
rect 17370 7808 17404 7824
rect 17370 6816 17404 6832
rect 17484 7808 17518 7824
rect 17484 6816 17518 6832
rect 17580 7808 17614 7824
rect 17580 6816 17614 6832
rect 17694 7808 17728 7824
rect 17694 6816 17728 6832
rect 17790 7808 17824 7824
rect 17790 6816 17824 6832
rect 17904 7808 17938 7824
rect 17904 6816 17938 6832
rect 18000 7808 18034 7824
rect 18000 6816 18034 6832
rect 18114 7808 18148 7824
rect 18114 6816 18148 6832
rect 18210 7808 18244 7824
rect 18210 6816 18244 6832
rect 18324 7808 18358 7824
rect 18324 6816 18358 6832
rect 18420 7808 18454 7824
rect 18420 6816 18454 6832
rect 18534 7808 18568 7824
rect 18534 6816 18568 6832
rect 18630 7808 18664 7824
rect 18630 6816 18664 6832
rect 10586 6739 10602 6773
rect 10586 6631 10602 6665
rect 10636 6739 10652 6773
rect 11006 6739 11022 6773
rect 10636 6631 10652 6665
rect 11006 6631 11022 6665
rect 11056 6739 11072 6773
rect 11426 6739 11442 6773
rect 11056 6631 11072 6665
rect 11426 6631 11442 6665
rect 11476 6739 11492 6773
rect 11846 6739 11862 6773
rect 11476 6631 11492 6665
rect 11846 6631 11862 6665
rect 11896 6739 11912 6773
rect 12266 6739 12282 6773
rect 11896 6631 11912 6665
rect 12266 6631 12282 6665
rect 12316 6739 12332 6773
rect 12686 6739 12702 6773
rect 12316 6631 12332 6665
rect 12686 6631 12702 6665
rect 12736 6739 12752 6773
rect 13106 6739 13122 6773
rect 12736 6631 12752 6665
rect 13106 6631 13122 6665
rect 13156 6739 13172 6773
rect 13526 6739 13542 6773
rect 13156 6631 13172 6665
rect 13526 6631 13542 6665
rect 13576 6739 13592 6773
rect 13946 6739 13962 6773
rect 13576 6631 13592 6665
rect 13946 6631 13962 6665
rect 13996 6739 14012 6773
rect 14366 6739 14382 6773
rect 13996 6631 14012 6665
rect 14366 6631 14382 6665
rect 14416 6739 14432 6773
rect 14786 6739 14802 6773
rect 14416 6631 14432 6665
rect 14786 6631 14802 6665
rect 14836 6739 14852 6773
rect 15206 6739 15222 6773
rect 14836 6631 14852 6665
rect 15206 6631 15222 6665
rect 15256 6739 15272 6773
rect 15626 6739 15642 6773
rect 15256 6631 15272 6665
rect 15626 6631 15642 6665
rect 15676 6739 15692 6773
rect 16046 6739 16062 6773
rect 15676 6631 15692 6665
rect 16046 6631 16062 6665
rect 16096 6739 16112 6773
rect 16466 6739 16482 6773
rect 16096 6631 16112 6665
rect 16466 6631 16482 6665
rect 16516 6739 16532 6773
rect 16886 6739 16902 6773
rect 16516 6631 16532 6665
rect 16886 6631 16902 6665
rect 16936 6739 16952 6773
rect 17306 6739 17322 6773
rect 16936 6631 16952 6665
rect 17306 6631 17322 6665
rect 17356 6739 17372 6773
rect 17726 6739 17742 6773
rect 17356 6631 17372 6665
rect 17726 6631 17742 6665
rect 17776 6739 17792 6773
rect 18146 6739 18162 6773
rect 17776 6631 17792 6665
rect 18146 6631 18162 6665
rect 18196 6739 18212 6773
rect 18566 6739 18582 6773
rect 18196 6631 18212 6665
rect 18566 6631 18582 6665
rect 18616 6739 18632 6773
rect 18616 6631 18632 6665
rect 10344 6572 10378 6588
rect 10344 5580 10378 5596
rect 10440 6572 10474 6588
rect 10440 5580 10474 5596
rect 10554 6572 10588 6588
rect 10554 5580 10588 5596
rect 10650 6572 10684 6588
rect 10650 5580 10684 5596
rect 10764 6572 10798 6588
rect 10764 5580 10798 5596
rect 10860 6572 10894 6588
rect 10860 5580 10894 5596
rect 10974 6572 11008 6588
rect 10974 5580 11008 5596
rect 11070 6572 11104 6588
rect 11070 5580 11104 5596
rect 11184 6572 11218 6588
rect 11184 5580 11218 5596
rect 11280 6572 11314 6588
rect 11280 5580 11314 5596
rect 11394 6572 11428 6588
rect 11394 5580 11428 5596
rect 11490 6572 11524 6588
rect 11490 5580 11524 5596
rect 11604 6572 11638 6588
rect 11604 5580 11638 5596
rect 11700 6572 11734 6588
rect 11700 5580 11734 5596
rect 11814 6572 11848 6588
rect 11814 5580 11848 5596
rect 11910 6572 11944 6588
rect 11910 5580 11944 5596
rect 12024 6572 12058 6588
rect 12024 5580 12058 5596
rect 12120 6572 12154 6588
rect 12120 5580 12154 5596
rect 12234 6572 12268 6588
rect 12234 5580 12268 5596
rect 12330 6572 12364 6588
rect 12330 5580 12364 5596
rect 12444 6572 12478 6588
rect 12444 5580 12478 5596
rect 12540 6572 12574 6588
rect 12540 5580 12574 5596
rect 12654 6572 12688 6588
rect 12654 5580 12688 5596
rect 12750 6572 12784 6588
rect 12750 5580 12784 5596
rect 12864 6572 12898 6588
rect 12864 5580 12898 5596
rect 12960 6572 12994 6588
rect 12960 5580 12994 5596
rect 13074 6572 13108 6588
rect 13074 5580 13108 5596
rect 13170 6572 13204 6588
rect 13170 5580 13204 5596
rect 13284 6572 13318 6588
rect 13284 5580 13318 5596
rect 13380 6572 13414 6588
rect 13380 5580 13414 5596
rect 13494 6572 13528 6588
rect 13494 5580 13528 5596
rect 13590 6572 13624 6588
rect 13590 5580 13624 5596
rect 13704 6572 13738 6588
rect 13704 5580 13738 5596
rect 13800 6572 13834 6588
rect 13800 5580 13834 5596
rect 13914 6572 13948 6588
rect 13914 5580 13948 5596
rect 14010 6572 14044 6588
rect 14010 5580 14044 5596
rect 14124 6572 14158 6588
rect 14124 5580 14158 5596
rect 14220 6572 14254 6588
rect 14220 5580 14254 5596
rect 14334 6572 14368 6588
rect 14334 5580 14368 5596
rect 14430 6572 14464 6588
rect 14430 5580 14464 5596
rect 14544 6572 14578 6588
rect 14544 5580 14578 5596
rect 14640 6572 14674 6588
rect 14640 5580 14674 5596
rect 14754 6572 14788 6588
rect 14754 5580 14788 5596
rect 14850 6572 14884 6588
rect 14850 5580 14884 5596
rect 14964 6572 14998 6588
rect 14964 5580 14998 5596
rect 15060 6572 15094 6588
rect 15060 5580 15094 5596
rect 15174 6572 15208 6588
rect 15174 5580 15208 5596
rect 15270 6572 15304 6588
rect 15270 5580 15304 5596
rect 15384 6572 15418 6588
rect 15384 5580 15418 5596
rect 15480 6572 15514 6588
rect 15480 5580 15514 5596
rect 15594 6572 15628 6588
rect 15594 5580 15628 5596
rect 15690 6572 15724 6588
rect 15690 5580 15724 5596
rect 15804 6572 15838 6588
rect 15804 5580 15838 5596
rect 15900 6572 15934 6588
rect 15900 5580 15934 5596
rect 16014 6572 16048 6588
rect 16014 5580 16048 5596
rect 16110 6572 16144 6588
rect 16110 5580 16144 5596
rect 16224 6572 16258 6588
rect 16224 5580 16258 5596
rect 16320 6572 16354 6588
rect 16320 5580 16354 5596
rect 16434 6572 16468 6588
rect 16434 5580 16468 5596
rect 16530 6572 16564 6588
rect 16530 5580 16564 5596
rect 16644 6572 16678 6588
rect 16644 5580 16678 5596
rect 16740 6572 16774 6588
rect 16740 5580 16774 5596
rect 16854 6572 16888 6588
rect 16854 5580 16888 5596
rect 16950 6572 16984 6588
rect 16950 5580 16984 5596
rect 17064 6572 17098 6588
rect 17064 5580 17098 5596
rect 17160 6572 17194 6588
rect 17160 5580 17194 5596
rect 17274 6572 17308 6588
rect 17274 5580 17308 5596
rect 17370 6572 17404 6588
rect 17370 5580 17404 5596
rect 17484 6572 17518 6588
rect 17484 5580 17518 5596
rect 17580 6572 17614 6588
rect 17580 5580 17614 5596
rect 17694 6572 17728 6588
rect 17694 5580 17728 5596
rect 17790 6572 17824 6588
rect 17790 5580 17824 5596
rect 17904 6572 17938 6588
rect 17904 5580 17938 5596
rect 18000 6572 18034 6588
rect 18000 5580 18034 5596
rect 18114 6572 18148 6588
rect 18114 5580 18148 5596
rect 18210 6572 18244 6588
rect 18210 5580 18244 5596
rect 18324 6572 18358 6588
rect 18324 5580 18358 5596
rect 18420 6572 18454 6588
rect 18420 5580 18454 5596
rect 18534 6572 18568 6588
rect 18534 5580 18568 5596
rect 18630 6572 18664 6588
rect 18630 5580 18664 5596
rect 10376 5503 10392 5537
rect 10376 5395 10392 5429
rect 10426 5503 10442 5537
rect 10796 5503 10812 5537
rect 10426 5395 10442 5429
rect 10796 5395 10812 5429
rect 10846 5503 10862 5537
rect 11216 5503 11232 5537
rect 10846 5395 10862 5429
rect 11216 5395 11232 5429
rect 11266 5503 11282 5537
rect 11636 5503 11652 5537
rect 11266 5395 11282 5429
rect 11636 5395 11652 5429
rect 11686 5503 11702 5537
rect 12056 5503 12072 5537
rect 11686 5395 11702 5429
rect 12056 5395 12072 5429
rect 12106 5503 12122 5537
rect 12476 5503 12492 5537
rect 12106 5395 12122 5429
rect 12476 5395 12492 5429
rect 12526 5503 12542 5537
rect 12896 5503 12912 5537
rect 12526 5395 12542 5429
rect 12896 5395 12912 5429
rect 12946 5503 12962 5537
rect 13316 5503 13332 5537
rect 12946 5395 12962 5429
rect 13316 5395 13332 5429
rect 13366 5503 13382 5537
rect 13736 5503 13752 5537
rect 13366 5395 13382 5429
rect 13736 5395 13752 5429
rect 13786 5503 13802 5537
rect 14156 5503 14172 5537
rect 13786 5395 13802 5429
rect 14156 5395 14172 5429
rect 14206 5503 14222 5537
rect 14576 5503 14592 5537
rect 14206 5395 14222 5429
rect 14576 5395 14592 5429
rect 14626 5503 14642 5537
rect 14996 5503 15012 5537
rect 14626 5395 14642 5429
rect 14996 5395 15012 5429
rect 15046 5503 15062 5537
rect 15416 5503 15432 5537
rect 15046 5395 15062 5429
rect 15416 5395 15432 5429
rect 15466 5503 15482 5537
rect 15836 5503 15852 5537
rect 15466 5395 15482 5429
rect 15836 5395 15852 5429
rect 15886 5503 15902 5537
rect 16256 5503 16272 5537
rect 15886 5395 15902 5429
rect 16256 5395 16272 5429
rect 16306 5503 16322 5537
rect 16676 5503 16692 5537
rect 16306 5395 16322 5429
rect 16676 5395 16692 5429
rect 16726 5503 16742 5537
rect 17096 5503 17112 5537
rect 16726 5395 16742 5429
rect 17096 5395 17112 5429
rect 17146 5503 17162 5537
rect 17516 5503 17532 5537
rect 17146 5395 17162 5429
rect 17516 5395 17532 5429
rect 17566 5503 17582 5537
rect 17936 5503 17952 5537
rect 17566 5395 17582 5429
rect 17936 5395 17952 5429
rect 17986 5503 18002 5537
rect 18356 5503 18372 5537
rect 17986 5395 18002 5429
rect 18356 5395 18372 5429
rect 18406 5503 18422 5537
rect 18406 5395 18422 5429
rect 10344 5336 10378 5352
rect 10344 4344 10378 4360
rect 10440 5336 10474 5352
rect 10440 4344 10474 4360
rect 10554 5336 10588 5352
rect 10554 4344 10588 4360
rect 10650 5336 10684 5352
rect 10650 4344 10684 4360
rect 10764 5336 10798 5352
rect 10764 4344 10798 4360
rect 10860 5336 10894 5352
rect 10860 4344 10894 4360
rect 10974 5336 11008 5352
rect 10974 4344 11008 4360
rect 11070 5336 11104 5352
rect 11070 4344 11104 4360
rect 11184 5336 11218 5352
rect 11184 4344 11218 4360
rect 11280 5336 11314 5352
rect 11280 4344 11314 4360
rect 11394 5336 11428 5352
rect 11394 4344 11428 4360
rect 11490 5336 11524 5352
rect 11490 4344 11524 4360
rect 11604 5336 11638 5352
rect 11604 4344 11638 4360
rect 11700 5336 11734 5352
rect 11700 4344 11734 4360
rect 11814 5336 11848 5352
rect 11814 4344 11848 4360
rect 11910 5336 11944 5352
rect 11910 4344 11944 4360
rect 12024 5336 12058 5352
rect 12024 4344 12058 4360
rect 12120 5336 12154 5352
rect 12120 4344 12154 4360
rect 12234 5336 12268 5352
rect 12234 4344 12268 4360
rect 12330 5336 12364 5352
rect 12330 4344 12364 4360
rect 12444 5336 12478 5352
rect 12444 4344 12478 4360
rect 12540 5336 12574 5352
rect 12540 4344 12574 4360
rect 12654 5336 12688 5352
rect 12654 4344 12688 4360
rect 12750 5336 12784 5352
rect 12750 4344 12784 4360
rect 12864 5336 12898 5352
rect 12864 4344 12898 4360
rect 12960 5336 12994 5352
rect 12960 4344 12994 4360
rect 13074 5336 13108 5352
rect 13074 4344 13108 4360
rect 13170 5336 13204 5352
rect 13170 4344 13204 4360
rect 13284 5336 13318 5352
rect 13284 4344 13318 4360
rect 13380 5336 13414 5352
rect 13380 4344 13414 4360
rect 13494 5336 13528 5352
rect 13494 4344 13528 4360
rect 13590 5336 13624 5352
rect 13590 4344 13624 4360
rect 13704 5336 13738 5352
rect 13704 4344 13738 4360
rect 13800 5336 13834 5352
rect 13800 4344 13834 4360
rect 13914 5336 13948 5352
rect 13914 4344 13948 4360
rect 14010 5336 14044 5352
rect 14010 4344 14044 4360
rect 14124 5336 14158 5352
rect 14124 4344 14158 4360
rect 14220 5336 14254 5352
rect 14220 4344 14254 4360
rect 14334 5336 14368 5352
rect 14334 4344 14368 4360
rect 14430 5336 14464 5352
rect 14430 4344 14464 4360
rect 14544 5336 14578 5352
rect 14544 4344 14578 4360
rect 14640 5336 14674 5352
rect 14640 4344 14674 4360
rect 14754 5336 14788 5352
rect 14754 4344 14788 4360
rect 14850 5336 14884 5352
rect 14850 4344 14884 4360
rect 14964 5336 14998 5352
rect 14964 4344 14998 4360
rect 15060 5336 15094 5352
rect 15060 4344 15094 4360
rect 15174 5336 15208 5352
rect 15174 4344 15208 4360
rect 15270 5336 15304 5352
rect 15270 4344 15304 4360
rect 15384 5336 15418 5352
rect 15384 4344 15418 4360
rect 15480 5336 15514 5352
rect 15480 4344 15514 4360
rect 15594 5336 15628 5352
rect 15594 4344 15628 4360
rect 15690 5336 15724 5352
rect 15690 4344 15724 4360
rect 15804 5336 15838 5352
rect 15804 4344 15838 4360
rect 15900 5336 15934 5352
rect 15900 4344 15934 4360
rect 16014 5336 16048 5352
rect 16014 4344 16048 4360
rect 16110 5336 16144 5352
rect 16110 4344 16144 4360
rect 16224 5336 16258 5352
rect 16224 4344 16258 4360
rect 16320 5336 16354 5352
rect 16320 4344 16354 4360
rect 16434 5336 16468 5352
rect 16434 4344 16468 4360
rect 16530 5336 16564 5352
rect 16530 4344 16564 4360
rect 16644 5336 16678 5352
rect 16644 4344 16678 4360
rect 16740 5336 16774 5352
rect 16740 4344 16774 4360
rect 16854 5336 16888 5352
rect 16854 4344 16888 4360
rect 16950 5336 16984 5352
rect 16950 4344 16984 4360
rect 17064 5336 17098 5352
rect 17064 4344 17098 4360
rect 17160 5336 17194 5352
rect 17160 4344 17194 4360
rect 17274 5336 17308 5352
rect 17274 4344 17308 4360
rect 17370 5336 17404 5352
rect 17370 4344 17404 4360
rect 17484 5336 17518 5352
rect 17484 4344 17518 4360
rect 17580 5336 17614 5352
rect 17580 4344 17614 4360
rect 17694 5336 17728 5352
rect 17694 4344 17728 4360
rect 17790 5336 17824 5352
rect 17790 4344 17824 4360
rect 17904 5336 17938 5352
rect 17904 4344 17938 4360
rect 18000 5336 18034 5352
rect 18000 4344 18034 4360
rect 18114 5336 18148 5352
rect 18114 4344 18148 4360
rect 18210 5336 18244 5352
rect 18210 4344 18244 4360
rect 18324 5336 18358 5352
rect 18324 4344 18358 4360
rect 18420 5336 18454 5352
rect 18420 4344 18454 4360
rect 18534 5336 18568 5352
rect 18534 4344 18568 4360
rect 18630 5336 18664 5352
rect 18630 4344 18664 4360
rect 10586 4267 10602 4301
rect 10586 4159 10602 4193
rect 10636 4267 10652 4301
rect 11006 4267 11022 4301
rect 10636 4159 10652 4193
rect 11006 4159 11022 4193
rect 11056 4267 11072 4301
rect 11426 4267 11442 4301
rect 11056 4159 11072 4193
rect 11426 4159 11442 4193
rect 11476 4267 11492 4301
rect 11846 4267 11862 4301
rect 11476 4159 11492 4193
rect 11846 4159 11862 4193
rect 11896 4267 11912 4301
rect 12266 4267 12282 4301
rect 11896 4159 11912 4193
rect 12266 4159 12282 4193
rect 12316 4267 12332 4301
rect 12686 4267 12702 4301
rect 12316 4159 12332 4193
rect 12686 4159 12702 4193
rect 12736 4267 12752 4301
rect 13106 4267 13122 4301
rect 12736 4159 12752 4193
rect 13106 4159 13122 4193
rect 13156 4267 13172 4301
rect 13526 4267 13542 4301
rect 13156 4159 13172 4193
rect 13526 4159 13542 4193
rect 13576 4267 13592 4301
rect 13946 4267 13962 4301
rect 13576 4159 13592 4193
rect 13946 4159 13962 4193
rect 13996 4267 14012 4301
rect 14366 4267 14382 4301
rect 13996 4159 14012 4193
rect 14366 4159 14382 4193
rect 14416 4267 14432 4301
rect 14786 4267 14802 4301
rect 14416 4159 14432 4193
rect 14786 4159 14802 4193
rect 14836 4267 14852 4301
rect 15206 4267 15222 4301
rect 14836 4159 14852 4193
rect 15206 4159 15222 4193
rect 15256 4267 15272 4301
rect 15626 4267 15642 4301
rect 15256 4159 15272 4193
rect 15626 4159 15642 4193
rect 15676 4267 15692 4301
rect 16046 4267 16062 4301
rect 15676 4159 15692 4193
rect 16046 4159 16062 4193
rect 16096 4267 16112 4301
rect 16466 4267 16482 4301
rect 16096 4159 16112 4193
rect 16466 4159 16482 4193
rect 16516 4267 16532 4301
rect 16886 4267 16902 4301
rect 16516 4159 16532 4193
rect 16886 4159 16902 4193
rect 16936 4267 16952 4301
rect 17306 4267 17322 4301
rect 16936 4159 16952 4193
rect 17306 4159 17322 4193
rect 17356 4267 17372 4301
rect 17726 4267 17742 4301
rect 17356 4159 17372 4193
rect 17726 4159 17742 4193
rect 17776 4267 17792 4301
rect 18146 4267 18162 4301
rect 17776 4159 17792 4193
rect 18146 4159 18162 4193
rect 18196 4267 18212 4301
rect 18566 4267 18582 4301
rect 18196 4159 18212 4193
rect 18566 4159 18582 4193
rect 18616 4267 18632 4301
rect 18616 4159 18632 4193
rect 10344 4100 10378 4116
rect 10344 3108 10378 3124
rect 10440 4100 10474 4116
rect 10440 3108 10474 3124
rect 10554 4100 10588 4116
rect 10554 3108 10588 3124
rect 10650 4100 10684 4116
rect 10650 3108 10684 3124
rect 10764 4100 10798 4116
rect 10764 3108 10798 3124
rect 10860 4100 10894 4116
rect 10860 3108 10894 3124
rect 10974 4100 11008 4116
rect 10974 3108 11008 3124
rect 11070 4100 11104 4116
rect 11070 3108 11104 3124
rect 11184 4100 11218 4116
rect 11184 3108 11218 3124
rect 11280 4100 11314 4116
rect 11280 3108 11314 3124
rect 11394 4100 11428 4116
rect 11394 3108 11428 3124
rect 11490 4100 11524 4116
rect 11490 3108 11524 3124
rect 11604 4100 11638 4116
rect 11604 3108 11638 3124
rect 11700 4100 11734 4116
rect 11700 3108 11734 3124
rect 11814 4100 11848 4116
rect 11814 3108 11848 3124
rect 11910 4100 11944 4116
rect 11910 3108 11944 3124
rect 12024 4100 12058 4116
rect 12024 3108 12058 3124
rect 12120 4100 12154 4116
rect 12120 3108 12154 3124
rect 12234 4100 12268 4116
rect 12234 3108 12268 3124
rect 12330 4100 12364 4116
rect 12330 3108 12364 3124
rect 12444 4100 12478 4116
rect 12444 3108 12478 3124
rect 12540 4100 12574 4116
rect 12540 3108 12574 3124
rect 12654 4100 12688 4116
rect 12654 3108 12688 3124
rect 12750 4100 12784 4116
rect 12750 3108 12784 3124
rect 12864 4100 12898 4116
rect 12864 3108 12898 3124
rect 12960 4100 12994 4116
rect 12960 3108 12994 3124
rect 13074 4100 13108 4116
rect 13074 3108 13108 3124
rect 13170 4100 13204 4116
rect 13170 3108 13204 3124
rect 13284 4100 13318 4116
rect 13284 3108 13318 3124
rect 13380 4100 13414 4116
rect 13380 3108 13414 3124
rect 13494 4100 13528 4116
rect 13494 3108 13528 3124
rect 13590 4100 13624 4116
rect 13590 3108 13624 3124
rect 13704 4100 13738 4116
rect 13704 3108 13738 3124
rect 13800 4100 13834 4116
rect 13800 3108 13834 3124
rect 13914 4100 13948 4116
rect 13914 3108 13948 3124
rect 14010 4100 14044 4116
rect 14010 3108 14044 3124
rect 14124 4100 14158 4116
rect 14124 3108 14158 3124
rect 14220 4100 14254 4116
rect 14220 3108 14254 3124
rect 14334 4100 14368 4116
rect 14334 3108 14368 3124
rect 14430 4100 14464 4116
rect 14430 3108 14464 3124
rect 14544 4100 14578 4116
rect 14544 3108 14578 3124
rect 14640 4100 14674 4116
rect 14640 3108 14674 3124
rect 14754 4100 14788 4116
rect 14754 3108 14788 3124
rect 14850 4100 14884 4116
rect 14850 3108 14884 3124
rect 14964 4100 14998 4116
rect 14964 3108 14998 3124
rect 15060 4100 15094 4116
rect 15060 3108 15094 3124
rect 15174 4100 15208 4116
rect 15174 3108 15208 3124
rect 15270 4100 15304 4116
rect 15270 3108 15304 3124
rect 15384 4100 15418 4116
rect 15384 3108 15418 3124
rect 15480 4100 15514 4116
rect 15480 3108 15514 3124
rect 15594 4100 15628 4116
rect 15594 3108 15628 3124
rect 15690 4100 15724 4116
rect 15690 3108 15724 3124
rect 15804 4100 15838 4116
rect 15804 3108 15838 3124
rect 15900 4100 15934 4116
rect 15900 3108 15934 3124
rect 16014 4100 16048 4116
rect 16014 3108 16048 3124
rect 16110 4100 16144 4116
rect 16110 3108 16144 3124
rect 16224 4100 16258 4116
rect 16224 3108 16258 3124
rect 16320 4100 16354 4116
rect 16320 3108 16354 3124
rect 16434 4100 16468 4116
rect 16434 3108 16468 3124
rect 16530 4100 16564 4116
rect 16530 3108 16564 3124
rect 16644 4100 16678 4116
rect 16644 3108 16678 3124
rect 16740 4100 16774 4116
rect 16740 3108 16774 3124
rect 16854 4100 16888 4116
rect 16854 3108 16888 3124
rect 16950 4100 16984 4116
rect 16950 3108 16984 3124
rect 17064 4100 17098 4116
rect 17064 3108 17098 3124
rect 17160 4100 17194 4116
rect 17160 3108 17194 3124
rect 17274 4100 17308 4116
rect 17274 3108 17308 3124
rect 17370 4100 17404 4116
rect 17370 3108 17404 3124
rect 17484 4100 17518 4116
rect 17484 3108 17518 3124
rect 17580 4100 17614 4116
rect 17580 3108 17614 3124
rect 17694 4100 17728 4116
rect 17694 3108 17728 3124
rect 17790 4100 17824 4116
rect 17790 3108 17824 3124
rect 17904 4100 17938 4116
rect 17904 3108 17938 3124
rect 18000 4100 18034 4116
rect 18000 3108 18034 3124
rect 18114 4100 18148 4116
rect 18114 3108 18148 3124
rect 18210 4100 18244 4116
rect 18210 3108 18244 3124
rect 18324 4100 18358 4116
rect 18324 3108 18358 3124
rect 18420 4100 18454 4116
rect 18420 3108 18454 3124
rect 18534 4100 18568 4116
rect 18534 3108 18568 3124
rect 18630 4100 18664 4116
rect 18630 3108 18664 3124
rect 10132 2922 10166 3046
rect 10376 3065 10427 3070
rect 10796 3065 10847 3070
rect 11216 3065 11267 3070
rect 11636 3065 11687 3070
rect 12056 3065 12107 3070
rect 12476 3065 12527 3070
rect 12896 3065 12947 3070
rect 13316 3065 13367 3070
rect 13736 3065 13787 3070
rect 14156 3065 14207 3070
rect 14576 3065 14627 3070
rect 14996 3065 15047 3070
rect 15416 3065 15467 3070
rect 15836 3065 15887 3070
rect 16256 3065 16307 3070
rect 16676 3065 16727 3070
rect 17096 3065 17147 3070
rect 17516 3065 17567 3070
rect 17936 3065 17987 3070
rect 18356 3065 18407 3070
rect 10376 3030 10392 3065
rect 10426 3064 10442 3065
rect 10476 3030 10492 3064
rect 10796 3030 10812 3065
rect 10846 3064 10862 3065
rect 10896 3030 10912 3064
rect 11216 3030 11232 3065
rect 11266 3064 11282 3065
rect 11316 3030 11332 3064
rect 11636 3030 11652 3065
rect 11686 3064 11702 3065
rect 11736 3030 11752 3064
rect 12056 3030 12072 3065
rect 12106 3064 12122 3065
rect 12156 3030 12172 3064
rect 12476 3030 12492 3065
rect 12526 3064 12542 3065
rect 12576 3030 12592 3064
rect 12896 3030 12912 3065
rect 12946 3064 12962 3065
rect 12996 3030 13012 3064
rect 13316 3030 13332 3065
rect 13366 3064 13382 3065
rect 13416 3030 13432 3064
rect 13736 3030 13752 3065
rect 13786 3064 13802 3065
rect 13836 3030 13852 3064
rect 14156 3030 14172 3065
rect 14206 3064 14222 3065
rect 14256 3030 14272 3064
rect 14576 3030 14592 3065
rect 14626 3064 14642 3065
rect 14676 3030 14692 3064
rect 14996 3030 15012 3065
rect 15046 3064 15062 3065
rect 15096 3030 15112 3064
rect 15416 3030 15432 3065
rect 15466 3064 15482 3065
rect 15516 3030 15532 3064
rect 15836 3030 15852 3065
rect 15886 3064 15902 3065
rect 15936 3030 15952 3064
rect 16256 3030 16272 3065
rect 16306 3064 16322 3065
rect 16356 3030 16372 3064
rect 16676 3030 16692 3065
rect 16726 3064 16742 3065
rect 16776 3030 16792 3064
rect 17096 3030 17112 3065
rect 17146 3064 17162 3065
rect 17196 3030 17212 3064
rect 17516 3030 17532 3065
rect 17566 3064 17582 3065
rect 17616 3030 17632 3064
rect 17936 3030 17952 3065
rect 17986 3064 18002 3065
rect 18036 3030 18052 3064
rect 18356 3030 18372 3065
rect 18406 3064 18422 3065
rect 18456 3030 18472 3064
rect 10376 3022 10427 3030
rect 10796 3022 10847 3030
rect 11216 3022 11267 3030
rect 11636 3022 11687 3030
rect 12056 3022 12107 3030
rect 12476 3022 12527 3030
rect 12896 3022 12947 3030
rect 13316 3022 13367 3030
rect 13736 3022 13787 3030
rect 14156 3022 14207 3030
rect 14576 3022 14627 3030
rect 14996 3022 15047 3030
rect 15416 3022 15467 3030
rect 15836 3022 15887 3030
rect 16256 3022 16307 3030
rect 16676 3022 16727 3030
rect 17096 3022 17147 3030
rect 17516 3022 17567 3030
rect 17936 3022 17987 3030
rect 18356 3022 18407 3030
rect 10132 2888 10208 2922
rect 18762 2922 18796 3108
rect 10308 2888 10322 2922
rect 18708 2888 18796 2922
rect 2710 -1506 2761 -1498
rect 2710 -1540 2726 -1506
rect 2810 -1540 2826 -1506
rect 2710 -1546 2761 -1540
rect 2582 -1598 2616 -1582
rect 2582 -2590 2616 -2574
rect 2678 -1598 2712 -1582
rect 2678 -2590 2712 -2574
rect 2774 -1598 2808 -1582
rect 3010 -1782 3104 -1312
rect 5466 -1412 5486 -1378
rect 9258 -1412 9332 -1378
rect 3352 -1504 3403 -1496
rect 3772 -1504 3823 -1496
rect 4192 -1504 4243 -1496
rect 4612 -1504 4663 -1496
rect 5384 -1500 5418 -1444
rect 3352 -1539 3368 -1504
rect 3452 -1538 3468 -1504
rect 3402 -1539 3418 -1538
rect 3772 -1539 3788 -1504
rect 3872 -1538 3888 -1504
rect 3822 -1539 3838 -1538
rect 4192 -1539 4208 -1504
rect 4292 -1538 4308 -1504
rect 4242 -1539 4258 -1538
rect 4612 -1539 4628 -1504
rect 4712 -1538 4728 -1504
rect 4662 -1539 4678 -1538
rect 3352 -1544 3403 -1539
rect 3772 -1544 3823 -1539
rect 4192 -1544 4243 -1539
rect 4612 -1544 4663 -1539
rect 3320 -1598 3354 -1582
rect 2924 -1798 3130 -1782
rect 2924 -2506 3130 -2490
rect 2774 -2590 2808 -2574
rect 3320 -2590 3354 -2574
rect 3416 -1598 3450 -1582
rect 3416 -2590 3450 -2574
rect 3530 -1598 3564 -1582
rect 3530 -2590 3564 -2574
rect 3626 -1598 3660 -1582
rect 3626 -2590 3660 -2574
rect 3740 -1598 3774 -1582
rect 3740 -2590 3774 -2574
rect 3836 -1598 3870 -1582
rect 3836 -2590 3870 -2574
rect 3950 -1598 3984 -1582
rect 3950 -2590 3984 -2574
rect 4046 -1598 4080 -1582
rect 4046 -2590 4080 -2574
rect 4160 -1598 4194 -1582
rect 4160 -2590 4194 -2574
rect 4256 -1598 4290 -1582
rect 4256 -2590 4290 -2574
rect 4370 -1598 4404 -1582
rect 4370 -2590 4404 -2574
rect 4466 -1598 4500 -1582
rect 4466 -2590 4500 -2574
rect 4580 -1598 4614 -1582
rect 4580 -2590 4614 -2574
rect 4676 -1598 4710 -1582
rect 4676 -2590 4710 -2574
rect 4790 -1598 4824 -1582
rect 4790 -2590 4824 -2574
rect 4886 -1598 4920 -1582
rect 4886 -2590 4920 -2574
rect 4402 -2632 4453 -2624
rect 4822 -2632 4873 -2624
rect 2614 -2667 2630 -2633
rect 2614 -2776 2630 -2742
rect 2664 -2667 2680 -2633
rect 3562 -2667 3578 -2633
rect 2664 -2776 2680 -2742
rect 3562 -2776 3578 -2742
rect 3612 -2667 3628 -2633
rect 3982 -2667 3998 -2633
rect 3612 -2776 3628 -2742
rect 3982 -2776 3998 -2742
rect 4032 -2667 4048 -2633
rect 4402 -2667 4418 -2632
rect 4502 -2666 4518 -2632
rect 4452 -2667 4468 -2666
rect 4822 -2667 4838 -2632
rect 4922 -2666 4938 -2632
rect 4872 -2667 4888 -2666
rect 4402 -2672 4453 -2667
rect 4822 -2672 4873 -2667
rect 4032 -2776 4048 -2742
rect 2586 -2826 2620 -2810
rect 2586 -3818 2620 -3802
rect 2674 -2826 2708 -2810
rect 3530 -2826 3564 -2810
rect 3000 -3000 3206 -2984
rect 3000 -3708 3206 -3692
rect 2674 -3818 2708 -3802
rect 3064 -3990 3160 -3708
rect 3530 -3818 3564 -3802
rect 3626 -2826 3660 -2810
rect 3626 -3818 3660 -3802
rect 3740 -2826 3774 -2810
rect 3740 -3818 3774 -3802
rect 3836 -2826 3870 -2810
rect 3836 -3818 3870 -3802
rect 3950 -2826 3984 -2810
rect 3950 -3818 3984 -3802
rect 4046 -2826 4080 -2810
rect 4046 -3818 4080 -3802
rect 4160 -2826 4194 -2810
rect 4160 -3818 4194 -3802
rect 4256 -2826 4290 -2810
rect 4256 -3818 4290 -3802
rect 3772 -3860 3823 -3852
rect 4192 -3860 4243 -3852
rect 3772 -3895 3788 -3860
rect 3872 -3894 3888 -3860
rect 3822 -3895 3838 -3894
rect 4192 -3895 4208 -3860
rect 4292 -3894 4308 -3860
rect 4242 -3895 4258 -3894
rect 3772 -3900 3823 -3895
rect 4192 -3900 4243 -3895
rect 5526 -1504 5577 -1496
rect 5946 -1504 5997 -1496
rect 6366 -1504 6417 -1496
rect 6786 -1504 6837 -1496
rect 7206 -1504 7257 -1496
rect 7626 -1504 7677 -1496
rect 8046 -1504 8097 -1496
rect 8466 -1504 8517 -1496
rect 8886 -1504 8937 -1496
rect 5526 -1539 5542 -1504
rect 5626 -1538 5642 -1504
rect 5576 -1539 5592 -1538
rect 5946 -1539 5962 -1504
rect 6046 -1538 6062 -1504
rect 5996 -1539 6012 -1538
rect 6366 -1539 6382 -1504
rect 6466 -1538 6482 -1504
rect 6416 -1539 6432 -1538
rect 6786 -1539 6802 -1504
rect 6886 -1538 6902 -1504
rect 6836 -1539 6852 -1538
rect 7206 -1539 7222 -1504
rect 7306 -1538 7322 -1504
rect 7256 -1539 7272 -1538
rect 7626 -1539 7642 -1504
rect 7726 -1538 7742 -1504
rect 7676 -1539 7692 -1538
rect 8046 -1539 8062 -1504
rect 8146 -1538 8162 -1504
rect 8096 -1539 8112 -1538
rect 8466 -1539 8482 -1504
rect 8566 -1538 8582 -1504
rect 8516 -1539 8532 -1538
rect 8886 -1539 8902 -1504
rect 8986 -1538 9002 -1504
rect 9298 -1538 9332 -1412
rect 8936 -1539 8952 -1538
rect 5526 -1544 5577 -1539
rect 5946 -1544 5997 -1539
rect 6366 -1544 6417 -1539
rect 6786 -1544 6837 -1539
rect 7206 -1544 7257 -1539
rect 7626 -1544 7677 -1539
rect 8046 -1544 8097 -1539
rect 8466 -1544 8517 -1539
rect 8886 -1544 8937 -1539
rect 5494 -1598 5528 -1582
rect 5494 -2590 5528 -2574
rect 5590 -1598 5624 -1582
rect 5590 -2590 5624 -2574
rect 5704 -1598 5738 -1582
rect 5704 -2590 5738 -2574
rect 5800 -1598 5834 -1582
rect 5800 -2590 5834 -2574
rect 5914 -1598 5948 -1582
rect 5914 -2590 5948 -2574
rect 6010 -1598 6044 -1582
rect 6010 -2590 6044 -2574
rect 6124 -1598 6158 -1582
rect 6124 -2590 6158 -2574
rect 6220 -1598 6254 -1582
rect 6220 -2590 6254 -2574
rect 6334 -1598 6368 -1582
rect 6334 -2590 6368 -2574
rect 6430 -1598 6464 -1582
rect 6430 -2590 6464 -2574
rect 6544 -1598 6578 -1582
rect 6544 -2590 6578 -2574
rect 6640 -1598 6674 -1582
rect 6640 -2590 6674 -2574
rect 6754 -1598 6788 -1582
rect 6754 -2590 6788 -2574
rect 6850 -1598 6884 -1582
rect 6850 -2590 6884 -2574
rect 6964 -1598 6998 -1582
rect 6964 -2590 6998 -2574
rect 7060 -1598 7094 -1582
rect 7060 -2590 7094 -2574
rect 7174 -1598 7208 -1582
rect 7174 -2590 7208 -2574
rect 7270 -1598 7304 -1582
rect 7270 -2590 7304 -2574
rect 7384 -1598 7418 -1582
rect 7384 -2590 7418 -2574
rect 7480 -1598 7514 -1582
rect 7480 -2590 7514 -2574
rect 7594 -1598 7628 -1582
rect 7594 -2590 7628 -2574
rect 7690 -1598 7724 -1582
rect 7690 -2590 7724 -2574
rect 7804 -1598 7838 -1582
rect 7804 -2590 7838 -2574
rect 7900 -1598 7934 -1582
rect 7900 -2590 7934 -2574
rect 8014 -1598 8048 -1582
rect 8014 -2590 8048 -2574
rect 8110 -1598 8144 -1582
rect 8110 -2590 8144 -2574
rect 8224 -1598 8258 -1582
rect 8224 -2590 8258 -2574
rect 8320 -1598 8354 -1582
rect 8320 -2590 8354 -2574
rect 8434 -1598 8468 -1582
rect 8434 -2590 8468 -2574
rect 8530 -1598 8564 -1582
rect 8530 -2590 8564 -2574
rect 8644 -1598 8678 -1582
rect 8644 -2590 8678 -2574
rect 8740 -1598 8774 -1582
rect 8740 -2590 8774 -2574
rect 8854 -1598 8888 -1582
rect 8854 -2590 8888 -2574
rect 8950 -1598 8984 -1582
rect 8950 -2590 8984 -2574
rect 9064 -1598 9098 -1582
rect 9064 -2590 9098 -2574
rect 9160 -1598 9194 -1582
rect 9160 -2590 9194 -2574
rect 5736 -2667 5752 -2633
rect 5736 -2775 5752 -2741
rect 5786 -2667 5802 -2633
rect 6156 -2667 6172 -2633
rect 5786 -2775 5802 -2741
rect 6156 -2775 6172 -2741
rect 6206 -2667 6222 -2633
rect 6576 -2667 6592 -2633
rect 6206 -2775 6222 -2741
rect 6576 -2775 6592 -2741
rect 6626 -2667 6642 -2633
rect 6996 -2667 7012 -2633
rect 6626 -2775 6642 -2741
rect 6996 -2775 7012 -2741
rect 7046 -2667 7062 -2633
rect 7416 -2667 7432 -2633
rect 7046 -2775 7062 -2741
rect 7416 -2775 7432 -2741
rect 7466 -2667 7482 -2633
rect 7836 -2667 7852 -2633
rect 7466 -2775 7482 -2741
rect 7836 -2775 7852 -2741
rect 7886 -2667 7902 -2633
rect 8256 -2667 8272 -2633
rect 7886 -2775 7902 -2741
rect 8256 -2775 8272 -2741
rect 8306 -2667 8322 -2633
rect 8676 -2667 8692 -2633
rect 8306 -2775 8322 -2741
rect 8676 -2775 8692 -2741
rect 8726 -2667 8742 -2633
rect 9096 -2667 9112 -2633
rect 8726 -2775 8742 -2741
rect 9096 -2775 9112 -2741
rect 9146 -2667 9162 -2633
rect 9146 -2775 9162 -2741
rect 5494 -2834 5528 -2818
rect 5494 -3826 5528 -3810
rect 5590 -2834 5624 -2818
rect 5590 -3826 5624 -3810
rect 5704 -2834 5738 -2818
rect 5704 -3826 5738 -3810
rect 5800 -2834 5834 -2818
rect 5800 -3826 5834 -3810
rect 5914 -2834 5948 -2818
rect 5914 -3826 5948 -3810
rect 6010 -2834 6044 -2818
rect 6010 -3826 6044 -3810
rect 6124 -2834 6158 -2818
rect 6124 -3826 6158 -3810
rect 6220 -2834 6254 -2818
rect 6220 -3826 6254 -3810
rect 6334 -2834 6368 -2818
rect 6334 -3826 6368 -3810
rect 6430 -2834 6464 -2818
rect 6430 -3826 6464 -3810
rect 6544 -2834 6578 -2818
rect 6544 -3826 6578 -3810
rect 6640 -2834 6674 -2818
rect 6640 -3826 6674 -3810
rect 6754 -2834 6788 -2818
rect 6754 -3826 6788 -3810
rect 6850 -2834 6884 -2818
rect 6850 -3826 6884 -3810
rect 6964 -2834 6998 -2818
rect 6964 -3826 6998 -3810
rect 7060 -2834 7094 -2818
rect 7060 -3826 7094 -3810
rect 7174 -2834 7208 -2818
rect 7174 -3826 7208 -3810
rect 7270 -2834 7304 -2818
rect 7270 -3826 7304 -3810
rect 7384 -2834 7418 -2818
rect 7384 -3826 7418 -3810
rect 7480 -2834 7514 -2818
rect 7480 -3826 7514 -3810
rect 7594 -2834 7628 -2818
rect 7594 -3826 7628 -3810
rect 7690 -2834 7724 -2818
rect 7690 -3826 7724 -3810
rect 7804 -2834 7838 -2818
rect 7804 -3826 7838 -3810
rect 7900 -2834 7934 -2818
rect 7900 -3826 7934 -3810
rect 8014 -2834 8048 -2818
rect 8014 -3826 8048 -3810
rect 8110 -2834 8144 -2818
rect 8110 -3826 8144 -3810
rect 8224 -2834 8258 -2818
rect 8224 -3826 8258 -3810
rect 8320 -2834 8354 -2818
rect 8320 -3826 8354 -3810
rect 8434 -2834 8468 -2818
rect 8434 -3826 8468 -3810
rect 8530 -2834 8564 -2818
rect 8530 -3826 8564 -3810
rect 8644 -2834 8678 -2818
rect 8644 -3826 8678 -3810
rect 8740 -2834 8774 -2818
rect 8740 -3826 8774 -3810
rect 8854 -2834 8888 -2818
rect 8854 -3826 8888 -3810
rect 8950 -2834 8984 -2818
rect 8950 -3826 8984 -3810
rect 9064 -2834 9098 -2818
rect 9064 -3826 9098 -3810
rect 9160 -2834 9194 -2818
rect 9160 -3826 9194 -3810
rect 5526 -3868 5577 -3860
rect 5946 -3868 5997 -3860
rect 6366 -3868 6417 -3860
rect 6786 -3868 6837 -3860
rect 7206 -3868 7257 -3860
rect 7626 -3868 7677 -3860
rect 8046 -3868 8097 -3860
rect 8466 -3868 8517 -3860
rect 8886 -3868 8937 -3860
rect 5526 -3903 5542 -3868
rect 5626 -3902 5642 -3868
rect 5576 -3903 5592 -3902
rect 5946 -3903 5962 -3868
rect 6046 -3902 6062 -3868
rect 5996 -3903 6012 -3902
rect 6366 -3903 6382 -3868
rect 6466 -3902 6482 -3868
rect 6416 -3903 6432 -3902
rect 6786 -3903 6802 -3868
rect 6886 -3902 6902 -3868
rect 6836 -3903 6852 -3902
rect 7206 -3903 7222 -3868
rect 7306 -3902 7322 -3868
rect 7256 -3903 7272 -3902
rect 7626 -3903 7642 -3868
rect 7726 -3902 7742 -3868
rect 7676 -3903 7692 -3902
rect 8046 -3903 8062 -3868
rect 8146 -3902 8162 -3868
rect 8096 -3903 8112 -3902
rect 8466 -3903 8482 -3868
rect 8566 -3902 8582 -3868
rect 8516 -3903 8532 -3902
rect 8886 -3903 8902 -3868
rect 8986 -3902 9002 -3868
rect 8936 -3903 8952 -3902
rect 5526 -3908 5577 -3903
rect 5946 -3908 5997 -3903
rect 6366 -3908 6417 -3903
rect 6786 -3908 6837 -3903
rect 7206 -3908 7257 -3903
rect 7626 -3908 7677 -3903
rect 8046 -3908 8097 -3903
rect 8466 -3908 8517 -3903
rect 8886 -3908 8937 -3903
rect 5384 -4010 5418 -3968
rect 9298 -4010 9332 -3826
rect 5384 -4044 5514 -4010
rect 9216 -4044 9332 -4010
rect 5348 -5716 5440 -5682
rect 9160 -5716 9310 -5682
rect 5348 -5834 5382 -5716
rect 5526 -5760 5577 -5752
rect 5946 -5760 5997 -5752
rect 6366 -5760 6417 -5752
rect 6786 -5760 6837 -5752
rect 7206 -5760 7257 -5752
rect 7626 -5760 7677 -5752
rect 8046 -5760 8097 -5752
rect 8466 -5760 8517 -5752
rect 8886 -5760 8937 -5752
rect 5526 -5795 5542 -5760
rect 5626 -5794 5642 -5760
rect 5576 -5795 5592 -5794
rect 5946 -5795 5962 -5760
rect 6046 -5794 6062 -5760
rect 5996 -5795 6012 -5794
rect 5526 -5800 5577 -5795
rect 5946 -5800 5997 -5795
rect 6366 -5800 6382 -5760
rect 6466 -5794 6482 -5760
rect 6416 -5800 6432 -5794
rect 6786 -5800 6802 -5760
rect 6886 -5794 6902 -5760
rect 6836 -5800 6852 -5794
rect 7206 -5800 7222 -5760
rect 7306 -5794 7322 -5760
rect 7256 -5800 7272 -5794
rect 7626 -5800 7642 -5760
rect 7726 -5794 7742 -5760
rect 7676 -5800 7692 -5794
rect 8046 -5800 8062 -5760
rect 8146 -5794 8162 -5760
rect 8096 -5800 8112 -5794
rect 8466 -5800 8482 -5760
rect 8566 -5794 8582 -5760
rect 8516 -5800 8532 -5794
rect 8886 -5800 8902 -5760
rect 8986 -5794 9002 -5760
rect 8936 -5800 8952 -5794
rect 5494 -5850 5528 -5834
rect 5494 -6842 5528 -6826
rect 5590 -5850 5624 -5834
rect 5590 -6842 5624 -6826
rect 5704 -5850 5738 -5834
rect 5704 -6842 5738 -6826
rect 5800 -5850 5834 -5834
rect 5800 -6842 5834 -6826
rect 5914 -5850 5948 -5834
rect 5914 -6842 5948 -6826
rect 6010 -5850 6044 -5834
rect 6010 -6842 6044 -6826
rect 6124 -5850 6158 -5834
rect 6124 -6842 6158 -6826
rect 6220 -5850 6254 -5834
rect 6220 -6842 6254 -6826
rect 6334 -5850 6368 -5834
rect 6334 -6842 6368 -6826
rect 6430 -5850 6464 -5834
rect 6430 -6842 6464 -6826
rect 6544 -5850 6578 -5834
rect 6544 -6842 6578 -6826
rect 6640 -5850 6674 -5834
rect 6640 -6842 6674 -6826
rect 6754 -5850 6788 -5834
rect 6754 -6842 6788 -6826
rect 6850 -5850 6884 -5834
rect 6850 -6842 6884 -6826
rect 6964 -5850 6998 -5834
rect 6964 -6842 6998 -6826
rect 7060 -5850 7094 -5834
rect 7060 -6842 7094 -6826
rect 7174 -5850 7208 -5834
rect 7174 -6842 7208 -6826
rect 7270 -5850 7304 -5834
rect 7270 -6842 7304 -6826
rect 7384 -5850 7418 -5834
rect 7384 -6842 7418 -6826
rect 7480 -5850 7514 -5834
rect 7480 -6842 7514 -6826
rect 7594 -5850 7628 -5834
rect 7594 -6842 7628 -6826
rect 7690 -5850 7724 -5834
rect 7690 -6842 7724 -6826
rect 7804 -5850 7838 -5834
rect 7804 -6842 7838 -6826
rect 7900 -5850 7934 -5834
rect 7900 -6842 7934 -6826
rect 8014 -5850 8048 -5834
rect 8014 -6842 8048 -6826
rect 8110 -5850 8144 -5834
rect 8110 -6842 8144 -6826
rect 8224 -5850 8258 -5834
rect 8224 -6842 8258 -6826
rect 8320 -5850 8354 -5834
rect 8320 -6842 8354 -6826
rect 8434 -5850 8468 -5834
rect 8434 -6842 8468 -6826
rect 8530 -5850 8564 -5834
rect 8530 -6842 8564 -6826
rect 8644 -5850 8678 -5834
rect 8644 -6842 8678 -6826
rect 8740 -5850 8774 -5834
rect 8740 -6842 8774 -6826
rect 8854 -5850 8888 -5834
rect 8854 -6842 8888 -6826
rect 8950 -5850 8984 -5834
rect 8950 -6842 8984 -6826
rect 9064 -5850 9098 -5834
rect 9064 -6842 9098 -6826
rect 9160 -5850 9194 -5834
rect 9160 -6842 9194 -6826
rect 9276 -5836 9310 -5716
rect 5348 -6970 5382 -6854
rect 5736 -6884 5787 -6876
rect 5736 -6918 5752 -6884
rect 5836 -6918 5852 -6884
rect 6156 -6918 6172 -6876
rect 6206 -6884 6222 -6876
rect 6256 -6918 6272 -6884
rect 6576 -6918 6592 -6876
rect 6626 -6884 6642 -6876
rect 6676 -6918 6692 -6884
rect 6996 -6918 7012 -6876
rect 7046 -6884 7062 -6876
rect 7096 -6918 7112 -6884
rect 7416 -6918 7432 -6876
rect 7466 -6884 7482 -6876
rect 7516 -6918 7532 -6884
rect 7836 -6918 7852 -6876
rect 7886 -6884 7902 -6876
rect 7936 -6918 7952 -6884
rect 8256 -6918 8272 -6876
rect 8306 -6884 8322 -6876
rect 8356 -6918 8372 -6884
rect 8676 -6918 8692 -6876
rect 8726 -6884 8742 -6876
rect 8776 -6918 8792 -6884
rect 9096 -6918 9112 -6876
rect 9146 -6884 9162 -6876
rect 9196 -6918 9212 -6884
rect 5736 -6919 5802 -6918
rect 6156 -6919 6222 -6918
rect 6576 -6919 6642 -6918
rect 6996 -6919 7062 -6918
rect 7416 -6919 7482 -6918
rect 7836 -6919 7902 -6918
rect 8256 -6919 8322 -6918
rect 8676 -6919 8742 -6918
rect 9096 -6919 9162 -6918
rect 5736 -6924 5787 -6919
rect 6156 -6924 6207 -6919
rect 6576 -6924 6627 -6919
rect 6996 -6924 7047 -6919
rect 7416 -6924 7467 -6919
rect 7836 -6924 7887 -6919
rect 8256 -6924 8307 -6919
rect 8676 -6924 8727 -6919
rect 9096 -6924 9147 -6919
rect 9276 -6970 9310 -6878
rect 5348 -7004 5480 -6970
rect 9204 -7004 9310 -6970
<< viali >>
rect 10302 13302 10400 13372
rect 10722 13302 10820 13372
rect 11142 13302 11240 13372
rect 11562 13302 11660 13372
rect 11982 13302 12080 13372
rect 12402 13302 12500 13372
rect 12822 13302 12920 13372
rect 13242 13302 13340 13372
rect 13662 13302 13760 13372
rect 14082 13302 14180 13372
rect 14502 13302 14600 13372
rect 14922 13302 15020 13372
rect 15342 13302 15440 13372
rect 15762 13302 15860 13372
rect 16182 13302 16280 13372
rect 16602 13302 16700 13372
rect 17022 13302 17120 13372
rect 17442 13302 17540 13372
rect 17862 13302 17960 13372
rect 18282 13302 18380 13372
rect 18630 13302 18728 13372
rect 10302 13268 10400 13302
rect 10722 13268 10820 13302
rect 11142 13268 11240 13302
rect 11562 13268 11660 13302
rect 11982 13268 12080 13302
rect 12402 13268 12500 13302
rect 12822 13268 12920 13302
rect 13242 13268 13340 13302
rect 13662 13268 13760 13302
rect 14082 13268 14180 13302
rect 14502 13268 14600 13302
rect 14922 13268 15020 13302
rect 15342 13268 15440 13302
rect 15762 13268 15860 13302
rect 16182 13268 16280 13302
rect 16602 13268 16700 13302
rect 17022 13268 17120 13302
rect 17442 13268 17540 13302
rect 17862 13268 17960 13302
rect 18282 13268 18380 13302
rect 18630 13268 18672 13302
rect 18672 13268 18728 13302
rect 10392 13086 10476 13120
rect 10812 13086 10896 13120
rect 11232 13086 11316 13120
rect 11652 13086 11736 13120
rect 12072 13086 12156 13120
rect 12492 13086 12576 13120
rect 12912 13086 12996 13120
rect 13332 13086 13416 13120
rect 13752 13086 13836 13120
rect 14172 13086 14256 13120
rect 14592 13086 14676 13120
rect 15012 13086 15096 13120
rect 15432 13086 15516 13120
rect 15852 13086 15936 13120
rect 16272 13086 16356 13120
rect 16692 13086 16776 13120
rect 17112 13086 17196 13120
rect 17532 13086 17616 13120
rect 17952 13086 18036 13120
rect 18372 13086 18456 13120
rect 10344 12060 10378 13036
rect 10440 12060 10474 13036
rect 10554 12060 10588 13036
rect 10650 12060 10684 13036
rect 10764 12060 10798 13036
rect 10860 12060 10894 13036
rect 10974 12060 11008 13036
rect 11070 12060 11104 13036
rect 11184 12060 11218 13036
rect 11280 12060 11314 13036
rect 11394 12060 11428 13036
rect 11490 12060 11524 13036
rect 11604 12060 11638 13036
rect 11700 12060 11734 13036
rect 11814 12060 11848 13036
rect 11910 12060 11944 13036
rect 12024 12060 12058 13036
rect 12120 12060 12154 13036
rect 12234 12060 12268 13036
rect 12330 12060 12364 13036
rect 12444 12060 12478 13036
rect 12540 12060 12574 13036
rect 12654 12060 12688 13036
rect 12750 12060 12784 13036
rect 12864 12060 12898 13036
rect 12960 12060 12994 13036
rect 13074 12060 13108 13036
rect 13170 12060 13204 13036
rect 13284 12060 13318 13036
rect 13380 12060 13414 13036
rect 13494 12060 13528 13036
rect 13590 12060 13624 13036
rect 13704 12060 13738 13036
rect 13800 12060 13834 13036
rect 13914 12060 13948 13036
rect 14010 12060 14044 13036
rect 14124 12060 14158 13036
rect 14220 12060 14254 13036
rect 14334 12060 14368 13036
rect 14430 12060 14464 13036
rect 14544 12060 14578 13036
rect 14640 12060 14674 13036
rect 14754 12060 14788 13036
rect 14850 12060 14884 13036
rect 14964 12060 14998 13036
rect 15060 12060 15094 13036
rect 15174 12060 15208 13036
rect 15270 12060 15304 13036
rect 15384 12060 15418 13036
rect 15480 12060 15514 13036
rect 15594 12060 15628 13036
rect 15690 12060 15724 13036
rect 15804 12060 15838 13036
rect 15900 12060 15934 13036
rect 16014 12060 16048 13036
rect 16110 12060 16144 13036
rect 16224 12060 16258 13036
rect 16320 12060 16354 13036
rect 16434 12060 16468 13036
rect 16530 12060 16564 13036
rect 16644 12060 16678 13036
rect 16740 12060 16774 13036
rect 16854 12060 16888 13036
rect 16950 12060 16984 13036
rect 17064 12060 17098 13036
rect 17160 12060 17194 13036
rect 17274 12060 17308 13036
rect 17370 12060 17404 13036
rect 17484 12060 17518 13036
rect 17580 12060 17614 13036
rect 17694 12060 17728 13036
rect 17790 12060 17824 13036
rect 17904 12060 17938 13036
rect 18000 12060 18034 13036
rect 18114 12060 18148 13036
rect 18210 12060 18244 13036
rect 18324 12060 18358 13036
rect 18420 12060 18454 13036
rect 18534 12060 18568 13036
rect 18630 12060 18664 13036
rect 10602 11868 10636 12010
rect 11022 11868 11056 12010
rect 11442 11868 11476 12010
rect 11862 11868 11896 12010
rect 12282 11868 12316 12010
rect 12702 11868 12736 12010
rect 13122 11868 13156 12010
rect 13542 11868 13576 12010
rect 13962 11868 13996 12010
rect 14382 11868 14416 12010
rect 14802 11868 14836 12010
rect 15222 11868 15256 12010
rect 15642 11868 15676 12010
rect 16062 11868 16096 12010
rect 16482 11868 16516 12010
rect 16902 11868 16936 12010
rect 17322 11868 17356 12010
rect 17742 11868 17776 12010
rect 18162 11868 18196 12010
rect 18582 11868 18616 12010
rect 10344 10842 10378 11818
rect 10440 10842 10474 11818
rect 10554 10842 10588 11818
rect 10650 10842 10684 11818
rect 10764 10842 10798 11818
rect 10860 10842 10894 11818
rect 10974 10842 11008 11818
rect 11070 10842 11104 11818
rect 11184 10842 11218 11818
rect 11280 10842 11314 11818
rect 11394 10842 11428 11818
rect 11490 10842 11524 11818
rect 11604 10842 11638 11818
rect 11700 10842 11734 11818
rect 11814 10842 11848 11818
rect 11910 10842 11944 11818
rect 12024 10842 12058 11818
rect 12120 10842 12154 11818
rect 12234 10842 12268 11818
rect 12330 10842 12364 11818
rect 12444 10842 12478 11818
rect 12540 10842 12574 11818
rect 12654 10842 12688 11818
rect 12750 10842 12784 11818
rect 12864 10842 12898 11818
rect 12960 10842 12994 11818
rect 13074 10842 13108 11818
rect 13170 10842 13204 11818
rect 13284 10842 13318 11818
rect 13380 10842 13414 11818
rect 13494 10842 13528 11818
rect 13590 10842 13624 11818
rect 13704 10842 13738 11818
rect 13800 10842 13834 11818
rect 13914 10842 13948 11818
rect 14010 10842 14044 11818
rect 14124 10842 14158 11818
rect 14220 10842 14254 11818
rect 14334 10842 14368 11818
rect 14430 10842 14464 11818
rect 14544 10842 14578 11818
rect 14640 10842 14674 11818
rect 14754 10842 14788 11818
rect 14850 10842 14884 11818
rect 14964 10842 14998 11818
rect 15060 10842 15094 11818
rect 15174 10842 15208 11818
rect 15270 10842 15304 11818
rect 15384 10842 15418 11818
rect 15480 10842 15514 11818
rect 15594 10842 15628 11818
rect 15690 10842 15724 11818
rect 15804 10842 15838 11818
rect 15900 10842 15934 11818
rect 16014 10842 16048 11818
rect 16110 10842 16144 11818
rect 16224 10842 16258 11818
rect 16320 10842 16354 11818
rect 16434 10842 16468 11818
rect 16530 10842 16564 11818
rect 16644 10842 16678 11818
rect 16740 10842 16774 11818
rect 16854 10842 16888 11818
rect 16950 10842 16984 11818
rect 17064 10842 17098 11818
rect 17160 10842 17194 11818
rect 17274 10842 17308 11818
rect 17370 10842 17404 11818
rect 17484 10842 17518 11818
rect 17580 10842 17614 11818
rect 17694 10842 17728 11818
rect 17790 10842 17824 11818
rect 17904 10842 17938 11818
rect 18000 10842 18034 11818
rect 18114 10842 18148 11818
rect 18210 10842 18244 11818
rect 18324 10842 18358 11818
rect 18420 10842 18454 11818
rect 18534 10842 18568 11818
rect 18630 10842 18664 11818
rect 10392 10758 10476 10792
rect 10812 10758 10896 10792
rect 11232 10758 11316 10792
rect 11652 10758 11736 10792
rect 12072 10758 12156 10792
rect 12492 10758 12576 10792
rect 12912 10758 12996 10792
rect 13332 10758 13416 10792
rect 13752 10758 13836 10792
rect 14172 10758 14256 10792
rect 14592 10758 14676 10792
rect 15012 10758 15096 10792
rect 15432 10758 15516 10792
rect 15852 10758 15936 10792
rect 16272 10758 16356 10792
rect 16692 10758 16776 10792
rect 17112 10758 17196 10792
rect 17532 10758 17616 10792
rect 17952 10758 18036 10792
rect 18372 10758 18456 10792
rect 10392 7900 10426 7901
rect 10392 7866 10476 7900
rect 10812 7900 10846 7901
rect 10812 7866 10896 7900
rect 11232 7900 11266 7901
rect 11232 7866 11316 7900
rect 11652 7900 11686 7901
rect 11652 7866 11736 7900
rect 12072 7900 12106 7901
rect 12072 7866 12156 7900
rect 12492 7900 12526 7901
rect 12492 7866 12576 7900
rect 12912 7900 12946 7901
rect 12912 7866 12996 7900
rect 13332 7900 13366 7901
rect 13332 7866 13416 7900
rect 13752 7900 13786 7901
rect 13752 7866 13836 7900
rect 14172 7900 14206 7901
rect 14172 7866 14256 7900
rect 14592 7900 14626 7901
rect 14592 7866 14676 7900
rect 15012 7900 15046 7901
rect 15012 7866 15096 7900
rect 15432 7900 15466 7901
rect 15432 7866 15516 7900
rect 15852 7900 15886 7901
rect 15852 7866 15936 7900
rect 16272 7900 16306 7901
rect 16272 7866 16356 7900
rect 16692 7900 16726 7901
rect 16692 7866 16776 7900
rect 17112 7900 17146 7901
rect 17112 7866 17196 7900
rect 17532 7900 17566 7901
rect 17532 7866 17616 7900
rect 17952 7900 17986 7901
rect 17952 7866 18036 7900
rect 18372 7900 18406 7901
rect 18372 7866 18456 7900
rect 5490 7130 5590 7230
rect 5910 7130 6010 7230
rect 6330 7130 6430 7230
rect 6750 7130 6850 7230
rect 7170 7130 7270 7230
rect 7590 7130 7690 7230
rect 8010 7130 8110 7230
rect 8430 7130 8530 7230
rect 8850 7130 8950 7230
rect 9176 7130 9276 7230
rect 5752 7010 5836 7044
rect 6172 7010 6256 7044
rect 6172 7002 6206 7010
rect 6592 7010 6676 7044
rect 6592 7002 6626 7010
rect 7012 7010 7096 7044
rect 7012 7002 7046 7010
rect 7432 7010 7516 7044
rect 7432 7002 7466 7010
rect 7852 7010 7936 7044
rect 7852 7002 7886 7010
rect 8272 7010 8356 7044
rect 8272 7002 8306 7010
rect 8692 7010 8776 7044
rect 8692 7002 8726 7010
rect 9112 7010 9196 7044
rect 9112 7002 9146 7010
rect 5494 5976 5528 6952
rect 5590 5976 5624 6952
rect 5704 5976 5738 6952
rect 5800 5976 5834 6952
rect 5914 5976 5948 6952
rect 6010 5976 6044 6952
rect 6124 5976 6158 6952
rect 6220 5976 6254 6952
rect 6334 5976 6368 6952
rect 6430 5976 6464 6952
rect 6544 5976 6578 6952
rect 6640 5976 6674 6952
rect 6754 5976 6788 6952
rect 6850 5976 6884 6952
rect 6964 5976 6998 6952
rect 7060 5976 7094 6952
rect 7174 5976 7208 6952
rect 7270 5976 7304 6952
rect 7384 5976 7418 6952
rect 7480 5976 7514 6952
rect 7594 5976 7628 6952
rect 7690 5976 7724 6952
rect 7804 5976 7838 6952
rect 7900 5976 7934 6952
rect 8014 5976 8048 6952
rect 8110 5976 8144 6952
rect 8224 5976 8258 6952
rect 8320 5976 8354 6952
rect 8434 5976 8468 6952
rect 8530 5976 8564 6952
rect 8644 5976 8678 6952
rect 8740 5976 8774 6952
rect 8854 5976 8888 6952
rect 8950 5976 8984 6952
rect 9064 5976 9098 6952
rect 9160 5976 9194 6952
rect 5542 5920 5576 5921
rect 5542 5886 5626 5920
rect 5962 5920 5996 5921
rect 5962 5886 6046 5920
rect 6382 5920 6416 5926
rect 6382 5886 6466 5920
rect 6802 5920 6836 5926
rect 6802 5886 6886 5920
rect 7222 5920 7256 5926
rect 7222 5886 7306 5920
rect 7642 5920 7676 5926
rect 7642 5886 7726 5920
rect 8062 5920 8096 5926
rect 8062 5886 8146 5920
rect 8482 5920 8516 5926
rect 8482 5886 8566 5920
rect 8902 5920 8936 5926
rect 8902 5886 8986 5920
rect 2950 5516 3248 5798
rect 2586 4352 2620 5328
rect 2674 4352 2708 5328
rect 3788 5420 3822 5421
rect 3788 5386 3872 5420
rect 4208 5420 4242 5421
rect 4208 5386 4292 5420
rect 3530 4352 3564 5328
rect 3626 4352 3660 5328
rect 3740 4352 3774 5328
rect 3836 4352 3870 5328
rect 3950 4352 3984 5328
rect 4046 4352 4080 5328
rect 4160 4352 4194 5328
rect 4256 4352 4290 5328
rect 2630 4159 2664 4302
rect 3578 4159 3612 4302
rect 3998 4159 4032 4302
rect 4418 4192 4452 4193
rect 4418 4158 4502 4192
rect 4838 4192 4872 4193
rect 4838 4158 4922 4192
rect 2582 3124 2616 4100
rect 2678 3124 2712 4100
rect 2774 3124 2808 4100
rect 2726 3032 2810 3066
rect 3320 3124 3354 4100
rect 3416 3124 3450 4100
rect 3530 3124 3564 4100
rect 3626 3124 3660 4100
rect 3740 3124 3774 4100
rect 3836 3124 3870 4100
rect 3950 3124 3984 4100
rect 4046 3124 4080 4100
rect 4160 3124 4194 4100
rect 4256 3124 4290 4100
rect 4370 3124 4404 4100
rect 4466 3124 4500 4100
rect 4580 3124 4614 4100
rect 4676 3124 4710 4100
rect 4790 3124 4824 4100
rect 4886 3124 4920 4100
rect 3368 3064 3402 3065
rect 3368 3030 3452 3064
rect 3788 3064 3822 3065
rect 3788 3030 3872 3064
rect 4208 3064 4242 3065
rect 4208 3030 4292 3064
rect 4628 3064 4662 3065
rect 4628 3030 4712 3064
rect 5542 5428 5576 5429
rect 5542 5394 5626 5428
rect 5962 5428 5996 5429
rect 5962 5394 6046 5428
rect 6382 5428 6416 5429
rect 6382 5394 6466 5428
rect 6802 5428 6836 5429
rect 6802 5394 6886 5428
rect 7222 5428 7256 5429
rect 7222 5394 7306 5428
rect 7642 5428 7676 5429
rect 7642 5394 7726 5428
rect 8062 5428 8096 5429
rect 8062 5394 8146 5428
rect 8482 5428 8516 5429
rect 8482 5394 8566 5428
rect 8902 5428 8936 5429
rect 8902 5394 8986 5428
rect 5494 4360 5528 5336
rect 5590 4360 5624 5336
rect 5704 4360 5738 5336
rect 5800 4360 5834 5336
rect 5914 4360 5948 5336
rect 6010 4360 6044 5336
rect 6124 4360 6158 5336
rect 6220 4360 6254 5336
rect 6334 4360 6368 5336
rect 6430 4360 6464 5336
rect 6544 4360 6578 5336
rect 6640 4360 6674 5336
rect 6754 4360 6788 5336
rect 6850 4360 6884 5336
rect 6964 4360 6998 5336
rect 7060 4360 7094 5336
rect 7174 4360 7208 5336
rect 7270 4360 7304 5336
rect 7384 4360 7418 5336
rect 7480 4360 7514 5336
rect 7594 4360 7628 5336
rect 7690 4360 7724 5336
rect 7804 4360 7838 5336
rect 7900 4360 7934 5336
rect 8014 4360 8048 5336
rect 8110 4360 8144 5336
rect 8224 4360 8258 5336
rect 8320 4360 8354 5336
rect 8434 4360 8468 5336
rect 8530 4360 8564 5336
rect 8644 4360 8678 5336
rect 8740 4360 8774 5336
rect 8854 4360 8888 5336
rect 8950 4360 8984 5336
rect 9064 4360 9098 5336
rect 9160 4360 9194 5336
rect 5752 4159 5786 4301
rect 6172 4159 6206 4301
rect 6592 4159 6626 4301
rect 7012 4159 7046 4301
rect 7432 4159 7466 4301
rect 7852 4159 7886 4301
rect 8272 4159 8306 4301
rect 8692 4159 8726 4301
rect 9112 4159 9146 4301
rect 5494 3124 5528 4100
rect 5590 3124 5624 4100
rect 5704 3124 5738 4100
rect 5800 3124 5834 4100
rect 5914 3124 5948 4100
rect 6010 3124 6044 4100
rect 6124 3124 6158 4100
rect 6220 3124 6254 4100
rect 6334 3124 6368 4100
rect 6430 3124 6464 4100
rect 6544 3124 6578 4100
rect 6640 3124 6674 4100
rect 6754 3124 6788 4100
rect 6850 3124 6884 4100
rect 6964 3124 6998 4100
rect 7060 3124 7094 4100
rect 7174 3124 7208 4100
rect 7270 3124 7304 4100
rect 7384 3124 7418 4100
rect 7480 3124 7514 4100
rect 7594 3124 7628 4100
rect 7690 3124 7724 4100
rect 7804 3124 7838 4100
rect 7900 3124 7934 4100
rect 8014 3124 8048 4100
rect 8110 3124 8144 4100
rect 8224 3124 8258 4100
rect 8320 3124 8354 4100
rect 8434 3124 8468 4100
rect 8530 3124 8564 4100
rect 8644 3124 8678 4100
rect 8740 3124 8774 4100
rect 8854 3124 8888 4100
rect 8950 3124 8984 4100
rect 9064 3124 9098 4100
rect 9160 3124 9194 4100
rect 5542 3064 5576 3065
rect 5542 3030 5626 3064
rect 5962 3064 5996 3065
rect 5962 3030 6046 3064
rect 6382 3064 6416 3065
rect 6382 3030 6466 3064
rect 6802 3064 6836 3065
rect 6802 3030 6886 3064
rect 7222 3064 7256 3065
rect 7222 3030 7306 3064
rect 7642 3064 7676 3065
rect 7642 3030 7726 3064
rect 8062 3064 8096 3065
rect 8062 3030 8146 3064
rect 8482 3064 8516 3065
rect 8482 3030 8566 3064
rect 8902 3064 8936 3065
rect 8902 3030 8986 3064
rect 5366 2870 5466 2970
rect 5786 2938 5886 2970
rect 6206 2938 6306 2970
rect 6626 2938 6726 2970
rect 7046 2938 7146 2970
rect 7466 2938 7566 2970
rect 7886 2938 7986 2970
rect 8306 2938 8406 2970
rect 8726 2938 8826 2970
rect 9146 2938 9246 2970
rect 5786 2904 5886 2938
rect 6206 2904 6306 2938
rect 6626 2904 6726 2938
rect 7046 2904 7146 2938
rect 7466 2904 7566 2938
rect 7886 2904 7986 2938
rect 8306 2904 8406 2938
rect 8726 2904 8826 2938
rect 9146 2904 9246 2938
rect 10344 6832 10378 7808
rect 10440 6832 10474 7808
rect 10554 6832 10588 7808
rect 10650 6832 10684 7808
rect 10764 6832 10798 7808
rect 10860 6832 10894 7808
rect 10974 6832 11008 7808
rect 11070 6832 11104 7808
rect 11184 6832 11218 7808
rect 11280 6832 11314 7808
rect 11394 6832 11428 7808
rect 11490 6832 11524 7808
rect 11604 6832 11638 7808
rect 11700 6832 11734 7808
rect 11814 6832 11848 7808
rect 11910 6832 11944 7808
rect 12024 6832 12058 7808
rect 12120 6832 12154 7808
rect 12234 6832 12268 7808
rect 12330 6832 12364 7808
rect 12444 6832 12478 7808
rect 12540 6832 12574 7808
rect 12654 6832 12688 7808
rect 12750 6832 12784 7808
rect 12864 6832 12898 7808
rect 12960 6832 12994 7808
rect 13074 6832 13108 7808
rect 13170 6832 13204 7808
rect 13284 6832 13318 7808
rect 13380 6832 13414 7808
rect 13494 6832 13528 7808
rect 13590 6832 13624 7808
rect 13704 6832 13738 7808
rect 13800 6832 13834 7808
rect 13914 6832 13948 7808
rect 14010 6832 14044 7808
rect 14124 6832 14158 7808
rect 14220 6832 14254 7808
rect 14334 6832 14368 7808
rect 14430 6832 14464 7808
rect 14544 6832 14578 7808
rect 14640 6832 14674 7808
rect 14754 6832 14788 7808
rect 14850 6832 14884 7808
rect 14964 6832 14998 7808
rect 15060 6832 15094 7808
rect 15174 6832 15208 7808
rect 15270 6832 15304 7808
rect 15384 6832 15418 7808
rect 15480 6832 15514 7808
rect 15594 6832 15628 7808
rect 15690 6832 15724 7808
rect 15804 6832 15838 7808
rect 15900 6832 15934 7808
rect 16014 6832 16048 7808
rect 16110 6832 16144 7808
rect 16224 6832 16258 7808
rect 16320 6832 16354 7808
rect 16434 6832 16468 7808
rect 16530 6832 16564 7808
rect 16644 6832 16678 7808
rect 16740 6832 16774 7808
rect 16854 6832 16888 7808
rect 16950 6832 16984 7808
rect 17064 6832 17098 7808
rect 17160 6832 17194 7808
rect 17274 6832 17308 7808
rect 17370 6832 17404 7808
rect 17484 6832 17518 7808
rect 17580 6832 17614 7808
rect 17694 6832 17728 7808
rect 17790 6832 17824 7808
rect 17904 6832 17938 7808
rect 18000 6832 18034 7808
rect 18114 6832 18148 7808
rect 18210 6832 18244 7808
rect 18324 6832 18358 7808
rect 18420 6832 18454 7808
rect 18534 6832 18568 7808
rect 18630 6832 18664 7808
rect 10602 6631 10636 6773
rect 11022 6631 11056 6773
rect 11442 6631 11476 6773
rect 11862 6631 11896 6773
rect 12282 6631 12316 6773
rect 12702 6631 12736 6773
rect 13122 6631 13156 6773
rect 13542 6631 13576 6773
rect 13962 6631 13996 6773
rect 14382 6631 14416 6773
rect 14802 6631 14836 6773
rect 15222 6631 15256 6773
rect 15642 6631 15676 6773
rect 16062 6631 16096 6773
rect 16482 6631 16516 6773
rect 16902 6631 16936 6773
rect 17322 6631 17356 6773
rect 17742 6631 17776 6773
rect 18162 6631 18196 6773
rect 18582 6631 18616 6773
rect 10344 5596 10378 6572
rect 10440 5596 10474 6572
rect 10554 5596 10588 6572
rect 10650 5596 10684 6572
rect 10764 5596 10798 6572
rect 10860 5596 10894 6572
rect 10974 5596 11008 6572
rect 11070 5596 11104 6572
rect 11184 5596 11218 6572
rect 11280 5596 11314 6572
rect 11394 5596 11428 6572
rect 11490 5596 11524 6572
rect 11604 5596 11638 6572
rect 11700 5596 11734 6572
rect 11814 5596 11848 6572
rect 11910 5596 11944 6572
rect 12024 5596 12058 6572
rect 12120 5596 12154 6572
rect 12234 5596 12268 6572
rect 12330 5596 12364 6572
rect 12444 5596 12478 6572
rect 12540 5596 12574 6572
rect 12654 5596 12688 6572
rect 12750 5596 12784 6572
rect 12864 5596 12898 6572
rect 12960 5596 12994 6572
rect 13074 5596 13108 6572
rect 13170 5596 13204 6572
rect 13284 5596 13318 6572
rect 13380 5596 13414 6572
rect 13494 5596 13528 6572
rect 13590 5596 13624 6572
rect 13704 5596 13738 6572
rect 13800 5596 13834 6572
rect 13914 5596 13948 6572
rect 14010 5596 14044 6572
rect 14124 5596 14158 6572
rect 14220 5596 14254 6572
rect 14334 5596 14368 6572
rect 14430 5596 14464 6572
rect 14544 5596 14578 6572
rect 14640 5596 14674 6572
rect 14754 5596 14788 6572
rect 14850 5596 14884 6572
rect 14964 5596 14998 6572
rect 15060 5596 15094 6572
rect 15174 5596 15208 6572
rect 15270 5596 15304 6572
rect 15384 5596 15418 6572
rect 15480 5596 15514 6572
rect 15594 5596 15628 6572
rect 15690 5596 15724 6572
rect 15804 5596 15838 6572
rect 15900 5596 15934 6572
rect 16014 5596 16048 6572
rect 16110 5596 16144 6572
rect 16224 5596 16258 6572
rect 16320 5596 16354 6572
rect 16434 5596 16468 6572
rect 16530 5596 16564 6572
rect 16644 5596 16678 6572
rect 16740 5596 16774 6572
rect 16854 5596 16888 6572
rect 16950 5596 16984 6572
rect 17064 5596 17098 6572
rect 17160 5596 17194 6572
rect 17274 5596 17308 6572
rect 17370 5596 17404 6572
rect 17484 5596 17518 6572
rect 17580 5596 17614 6572
rect 17694 5596 17728 6572
rect 17790 5596 17824 6572
rect 17904 5596 17938 6572
rect 18000 5596 18034 6572
rect 18114 5596 18148 6572
rect 18210 5596 18244 6572
rect 18324 5596 18358 6572
rect 18420 5596 18454 6572
rect 18534 5596 18568 6572
rect 18630 5596 18664 6572
rect 10392 5395 10426 5537
rect 10812 5395 10846 5537
rect 11232 5395 11266 5537
rect 11652 5395 11686 5537
rect 12072 5395 12106 5537
rect 12492 5395 12526 5537
rect 12912 5395 12946 5537
rect 13332 5395 13366 5537
rect 13752 5395 13786 5537
rect 14172 5395 14206 5537
rect 14592 5395 14626 5537
rect 15012 5395 15046 5537
rect 15432 5395 15466 5537
rect 15852 5395 15886 5537
rect 16272 5395 16306 5537
rect 16692 5395 16726 5537
rect 17112 5395 17146 5537
rect 17532 5395 17566 5537
rect 17952 5395 17986 5537
rect 18372 5395 18406 5537
rect 10344 4360 10378 5336
rect 10440 4360 10474 5336
rect 10554 4360 10588 5336
rect 10650 4360 10684 5336
rect 10764 4360 10798 5336
rect 10860 4360 10894 5336
rect 10974 4360 11008 5336
rect 11070 4360 11104 5336
rect 11184 4360 11218 5336
rect 11280 4360 11314 5336
rect 11394 4360 11428 5336
rect 11490 4360 11524 5336
rect 11604 4360 11638 5336
rect 11700 4360 11734 5336
rect 11814 4360 11848 5336
rect 11910 4360 11944 5336
rect 12024 4360 12058 5336
rect 12120 4360 12154 5336
rect 12234 4360 12268 5336
rect 12330 4360 12364 5336
rect 12444 4360 12478 5336
rect 12540 4360 12574 5336
rect 12654 4360 12688 5336
rect 12750 4360 12784 5336
rect 12864 4360 12898 5336
rect 12960 4360 12994 5336
rect 13074 4360 13108 5336
rect 13170 4360 13204 5336
rect 13284 4360 13318 5336
rect 13380 4360 13414 5336
rect 13494 4360 13528 5336
rect 13590 4360 13624 5336
rect 13704 4360 13738 5336
rect 13800 4360 13834 5336
rect 13914 4360 13948 5336
rect 14010 4360 14044 5336
rect 14124 4360 14158 5336
rect 14220 4360 14254 5336
rect 14334 4360 14368 5336
rect 14430 4360 14464 5336
rect 14544 4360 14578 5336
rect 14640 4360 14674 5336
rect 14754 4360 14788 5336
rect 14850 4360 14884 5336
rect 14964 4360 14998 5336
rect 15060 4360 15094 5336
rect 15174 4360 15208 5336
rect 15270 4360 15304 5336
rect 15384 4360 15418 5336
rect 15480 4360 15514 5336
rect 15594 4360 15628 5336
rect 15690 4360 15724 5336
rect 15804 4360 15838 5336
rect 15900 4360 15934 5336
rect 16014 4360 16048 5336
rect 16110 4360 16144 5336
rect 16224 4360 16258 5336
rect 16320 4360 16354 5336
rect 16434 4360 16468 5336
rect 16530 4360 16564 5336
rect 16644 4360 16678 5336
rect 16740 4360 16774 5336
rect 16854 4360 16888 5336
rect 16950 4360 16984 5336
rect 17064 4360 17098 5336
rect 17160 4360 17194 5336
rect 17274 4360 17308 5336
rect 17370 4360 17404 5336
rect 17484 4360 17518 5336
rect 17580 4360 17614 5336
rect 17694 4360 17728 5336
rect 17790 4360 17824 5336
rect 17904 4360 17938 5336
rect 18000 4360 18034 5336
rect 18114 4360 18148 5336
rect 18210 4360 18244 5336
rect 18324 4360 18358 5336
rect 18420 4360 18454 5336
rect 18534 4360 18568 5336
rect 18630 4360 18664 5336
rect 10602 4159 10636 4301
rect 11022 4159 11056 4301
rect 11442 4159 11476 4301
rect 11862 4159 11896 4301
rect 12282 4159 12316 4301
rect 12702 4159 12736 4301
rect 13122 4159 13156 4301
rect 13542 4159 13576 4301
rect 13962 4159 13996 4301
rect 14382 4159 14416 4301
rect 14802 4159 14836 4301
rect 15222 4159 15256 4301
rect 15642 4159 15676 4301
rect 16062 4159 16096 4301
rect 16482 4159 16516 4301
rect 16902 4159 16936 4301
rect 17322 4159 17356 4301
rect 17742 4159 17776 4301
rect 18162 4159 18196 4301
rect 18582 4159 18616 4301
rect 10344 3124 10378 4100
rect 10440 3124 10474 4100
rect 10554 3124 10588 4100
rect 10650 3124 10684 4100
rect 10764 3124 10798 4100
rect 10860 3124 10894 4100
rect 10974 3124 11008 4100
rect 11070 3124 11104 4100
rect 11184 3124 11218 4100
rect 11280 3124 11314 4100
rect 11394 3124 11428 4100
rect 11490 3124 11524 4100
rect 11604 3124 11638 4100
rect 11700 3124 11734 4100
rect 11814 3124 11848 4100
rect 11910 3124 11944 4100
rect 12024 3124 12058 4100
rect 12120 3124 12154 4100
rect 12234 3124 12268 4100
rect 12330 3124 12364 4100
rect 12444 3124 12478 4100
rect 12540 3124 12574 4100
rect 12654 3124 12688 4100
rect 12750 3124 12784 4100
rect 12864 3124 12898 4100
rect 12960 3124 12994 4100
rect 13074 3124 13108 4100
rect 13170 3124 13204 4100
rect 13284 3124 13318 4100
rect 13380 3124 13414 4100
rect 13494 3124 13528 4100
rect 13590 3124 13624 4100
rect 13704 3124 13738 4100
rect 13800 3124 13834 4100
rect 13914 3124 13948 4100
rect 14010 3124 14044 4100
rect 14124 3124 14158 4100
rect 14220 3124 14254 4100
rect 14334 3124 14368 4100
rect 14430 3124 14464 4100
rect 14544 3124 14578 4100
rect 14640 3124 14674 4100
rect 14754 3124 14788 4100
rect 14850 3124 14884 4100
rect 14964 3124 14998 4100
rect 15060 3124 15094 4100
rect 15174 3124 15208 4100
rect 15270 3124 15304 4100
rect 15384 3124 15418 4100
rect 15480 3124 15514 4100
rect 15594 3124 15628 4100
rect 15690 3124 15724 4100
rect 15804 3124 15838 4100
rect 15900 3124 15934 4100
rect 16014 3124 16048 4100
rect 16110 3124 16144 4100
rect 16224 3124 16258 4100
rect 16320 3124 16354 4100
rect 16434 3124 16468 4100
rect 16530 3124 16564 4100
rect 16644 3124 16678 4100
rect 16740 3124 16774 4100
rect 16854 3124 16888 4100
rect 16950 3124 16984 4100
rect 17064 3124 17098 4100
rect 17160 3124 17194 4100
rect 17274 3124 17308 4100
rect 17370 3124 17404 4100
rect 17484 3124 17518 4100
rect 17580 3124 17614 4100
rect 17694 3124 17728 4100
rect 17790 3124 17824 4100
rect 17904 3124 17938 4100
rect 18000 3124 18034 4100
rect 18114 3124 18148 4100
rect 18210 3124 18244 4100
rect 18324 3124 18358 4100
rect 18420 3124 18454 4100
rect 18534 3124 18568 4100
rect 18630 3124 18664 4100
rect 10392 3064 10426 3065
rect 10392 3030 10476 3064
rect 10812 3064 10846 3065
rect 10812 3030 10896 3064
rect 11232 3064 11266 3065
rect 11232 3030 11316 3064
rect 11652 3064 11686 3065
rect 11652 3030 11736 3064
rect 12072 3064 12106 3065
rect 12072 3030 12156 3064
rect 12492 3064 12526 3065
rect 12492 3030 12576 3064
rect 12912 3064 12946 3065
rect 12912 3030 12996 3064
rect 13332 3064 13366 3065
rect 13332 3030 13416 3064
rect 13752 3064 13786 3065
rect 13752 3030 13836 3064
rect 14172 3064 14206 3065
rect 14172 3030 14256 3064
rect 14592 3064 14626 3065
rect 14592 3030 14676 3064
rect 15012 3064 15046 3065
rect 15012 3030 15096 3064
rect 15432 3064 15466 3065
rect 15432 3030 15516 3064
rect 15852 3064 15886 3065
rect 15852 3030 15936 3064
rect 16272 3064 16306 3065
rect 16272 3030 16356 3064
rect 16692 3064 16726 3065
rect 16692 3030 16776 3064
rect 17112 3064 17146 3065
rect 17112 3030 17196 3064
rect 17532 3064 17566 3065
rect 17532 3030 17616 3064
rect 17952 3064 17986 3065
rect 17952 3030 18036 3064
rect 18372 3064 18406 3065
rect 18372 3030 18456 3064
rect 5786 2870 5886 2904
rect 6206 2870 6306 2904
rect 6626 2870 6726 2904
rect 7046 2870 7146 2904
rect 7466 2870 7566 2904
rect 7886 2870 7986 2904
rect 8306 2870 8406 2904
rect 8726 2870 8826 2904
rect 9146 2870 9246 2904
rect 10208 2854 10308 2954
rect 10628 2922 10728 2954
rect 11048 2922 11148 2954
rect 11468 2922 11568 2954
rect 11888 2922 11988 2954
rect 12308 2922 12408 2954
rect 12728 2922 12828 2954
rect 13148 2922 13248 2954
rect 13568 2922 13668 2954
rect 13988 2922 14088 2954
rect 14408 2922 14508 2954
rect 14828 2922 14928 2954
rect 15248 2922 15348 2954
rect 15668 2922 15768 2954
rect 16088 2922 16188 2954
rect 16508 2922 16608 2954
rect 16928 2922 17028 2954
rect 17348 2922 17448 2954
rect 17768 2922 17868 2954
rect 18188 2922 18288 2954
rect 18608 2922 18708 2954
rect 10628 2888 10728 2922
rect 11048 2888 11148 2922
rect 11468 2888 11568 2922
rect 11888 2888 11988 2922
rect 12308 2888 12408 2922
rect 12728 2888 12828 2922
rect 13148 2888 13248 2922
rect 13568 2888 13668 2922
rect 13988 2888 14088 2922
rect 14408 2888 14508 2922
rect 14828 2888 14928 2922
rect 15248 2888 15348 2922
rect 15668 2888 15768 2922
rect 16088 2888 16188 2922
rect 16508 2888 16608 2922
rect 16928 2888 17028 2922
rect 17348 2888 17448 2922
rect 17768 2888 17868 2922
rect 18188 2888 18288 2922
rect 18608 2888 18644 2922
rect 18644 2888 18708 2922
rect 10628 2854 10728 2888
rect 11048 2854 11148 2888
rect 11468 2854 11568 2888
rect 11888 2854 11988 2888
rect 12308 2854 12408 2888
rect 12728 2854 12828 2888
rect 13148 2854 13248 2888
rect 13568 2854 13668 2888
rect 13988 2854 14088 2888
rect 14408 2854 14508 2888
rect 14828 2854 14928 2888
rect 15248 2854 15348 2888
rect 15668 2854 15768 2888
rect 16088 2854 16188 2888
rect 16508 2854 16608 2888
rect 16928 2854 17028 2888
rect 17348 2854 17448 2888
rect 17768 2854 17868 2888
rect 18188 2854 18288 2888
rect 18608 2854 18708 2888
rect 2984 2690 3128 2838
rect 2984 -1312 3128 -1164
rect 2726 -1540 2810 -1506
rect 2582 -2574 2616 -1598
rect 2678 -2574 2712 -1598
rect 2774 -2574 2808 -1598
rect 5366 -1444 5466 -1344
rect 5786 -1378 5886 -1344
rect 6206 -1378 6306 -1344
rect 6626 -1378 6726 -1344
rect 7046 -1378 7146 -1344
rect 7466 -1378 7566 -1344
rect 7886 -1378 7986 -1344
rect 8306 -1378 8406 -1344
rect 8726 -1378 8826 -1344
rect 9146 -1378 9246 -1344
rect 5786 -1412 5886 -1378
rect 6206 -1412 6306 -1378
rect 6626 -1412 6726 -1378
rect 7046 -1412 7146 -1378
rect 7466 -1412 7566 -1378
rect 7886 -1412 7986 -1378
rect 8306 -1412 8406 -1378
rect 8726 -1412 8826 -1378
rect 9146 -1412 9246 -1378
rect 5786 -1444 5886 -1412
rect 6206 -1444 6306 -1412
rect 6626 -1444 6726 -1412
rect 7046 -1444 7146 -1412
rect 7466 -1444 7566 -1412
rect 7886 -1444 7986 -1412
rect 8306 -1444 8406 -1412
rect 8726 -1444 8826 -1412
rect 9146 -1444 9246 -1412
rect 3368 -1538 3452 -1504
rect 3368 -1539 3402 -1538
rect 3788 -1538 3872 -1504
rect 3788 -1539 3822 -1538
rect 4208 -1538 4292 -1504
rect 4208 -1539 4242 -1538
rect 4628 -1538 4712 -1504
rect 4628 -1539 4662 -1538
rect 3320 -2574 3354 -1598
rect 3416 -2574 3450 -1598
rect 3530 -2574 3564 -1598
rect 3626 -2574 3660 -1598
rect 3740 -2574 3774 -1598
rect 3836 -2574 3870 -1598
rect 3950 -2574 3984 -1598
rect 4046 -2574 4080 -1598
rect 4160 -2574 4194 -1598
rect 4256 -2574 4290 -1598
rect 4370 -2574 4404 -1598
rect 4466 -2574 4500 -1598
rect 4580 -2574 4614 -1598
rect 4676 -2574 4710 -1598
rect 4790 -2574 4824 -1598
rect 4886 -2574 4920 -1598
rect 2630 -2776 2664 -2633
rect 3578 -2776 3612 -2633
rect 3998 -2776 4032 -2633
rect 4418 -2666 4502 -2632
rect 4418 -2667 4452 -2666
rect 4838 -2666 4922 -2632
rect 4838 -2667 4872 -2666
rect 2586 -3802 2620 -2826
rect 2674 -3802 2708 -2826
rect 3530 -3802 3564 -2826
rect 3626 -3802 3660 -2826
rect 3740 -3802 3774 -2826
rect 3836 -3802 3870 -2826
rect 3950 -3802 3984 -2826
rect 4046 -3802 4080 -2826
rect 4160 -3802 4194 -2826
rect 4256 -3802 4290 -2826
rect 3788 -3894 3872 -3860
rect 3788 -3895 3822 -3894
rect 4208 -3894 4292 -3860
rect 4208 -3895 4242 -3894
rect 5542 -1538 5626 -1504
rect 5542 -1539 5576 -1538
rect 5962 -1538 6046 -1504
rect 5962 -1539 5996 -1538
rect 6382 -1538 6466 -1504
rect 6382 -1539 6416 -1538
rect 6802 -1538 6886 -1504
rect 6802 -1539 6836 -1538
rect 7222 -1538 7306 -1504
rect 7222 -1539 7256 -1538
rect 7642 -1538 7726 -1504
rect 7642 -1539 7676 -1538
rect 8062 -1538 8146 -1504
rect 8062 -1539 8096 -1538
rect 8482 -1538 8566 -1504
rect 8482 -1539 8516 -1538
rect 8902 -1538 8986 -1504
rect 8902 -1539 8936 -1538
rect 5494 -2574 5528 -1598
rect 5590 -2574 5624 -1598
rect 5704 -2574 5738 -1598
rect 5800 -2574 5834 -1598
rect 5914 -2574 5948 -1598
rect 6010 -2574 6044 -1598
rect 6124 -2574 6158 -1598
rect 6220 -2574 6254 -1598
rect 6334 -2574 6368 -1598
rect 6430 -2574 6464 -1598
rect 6544 -2574 6578 -1598
rect 6640 -2574 6674 -1598
rect 6754 -2574 6788 -1598
rect 6850 -2574 6884 -1598
rect 6964 -2574 6998 -1598
rect 7060 -2574 7094 -1598
rect 7174 -2574 7208 -1598
rect 7270 -2574 7304 -1598
rect 7384 -2574 7418 -1598
rect 7480 -2574 7514 -1598
rect 7594 -2574 7628 -1598
rect 7690 -2574 7724 -1598
rect 7804 -2574 7838 -1598
rect 7900 -2574 7934 -1598
rect 8014 -2574 8048 -1598
rect 8110 -2574 8144 -1598
rect 8224 -2574 8258 -1598
rect 8320 -2574 8354 -1598
rect 8434 -2574 8468 -1598
rect 8530 -2574 8564 -1598
rect 8644 -2574 8678 -1598
rect 8740 -2574 8774 -1598
rect 8854 -2574 8888 -1598
rect 8950 -2574 8984 -1598
rect 9064 -2574 9098 -1598
rect 9160 -2574 9194 -1598
rect 5752 -2775 5786 -2633
rect 6172 -2775 6206 -2633
rect 6592 -2775 6626 -2633
rect 7012 -2775 7046 -2633
rect 7432 -2775 7466 -2633
rect 7852 -2775 7886 -2633
rect 8272 -2775 8306 -2633
rect 8692 -2775 8726 -2633
rect 9112 -2775 9146 -2633
rect 5494 -3810 5528 -2834
rect 5590 -3810 5624 -2834
rect 5704 -3810 5738 -2834
rect 5800 -3810 5834 -2834
rect 5914 -3810 5948 -2834
rect 6010 -3810 6044 -2834
rect 6124 -3810 6158 -2834
rect 6220 -3810 6254 -2834
rect 6334 -3810 6368 -2834
rect 6430 -3810 6464 -2834
rect 6544 -3810 6578 -2834
rect 6640 -3810 6674 -2834
rect 6754 -3810 6788 -2834
rect 6850 -3810 6884 -2834
rect 6964 -3810 6998 -2834
rect 7060 -3810 7094 -2834
rect 7174 -3810 7208 -2834
rect 7270 -3810 7304 -2834
rect 7384 -3810 7418 -2834
rect 7480 -3810 7514 -2834
rect 7594 -3810 7628 -2834
rect 7690 -3810 7724 -2834
rect 7804 -3810 7838 -2834
rect 7900 -3810 7934 -2834
rect 8014 -3810 8048 -2834
rect 8110 -3810 8144 -2834
rect 8224 -3810 8258 -2834
rect 8320 -3810 8354 -2834
rect 8434 -3810 8468 -2834
rect 8530 -3810 8564 -2834
rect 8644 -3810 8678 -2834
rect 8740 -3810 8774 -2834
rect 8854 -3810 8888 -2834
rect 8950 -3810 8984 -2834
rect 9064 -3810 9098 -2834
rect 9160 -3810 9194 -2834
rect 5542 -3902 5626 -3868
rect 5542 -3903 5576 -3902
rect 5962 -3902 6046 -3868
rect 5962 -3903 5996 -3902
rect 6382 -3902 6466 -3868
rect 6382 -3903 6416 -3902
rect 6802 -3902 6886 -3868
rect 6802 -3903 6836 -3902
rect 7222 -3902 7306 -3868
rect 7222 -3903 7256 -3902
rect 7642 -3902 7726 -3868
rect 7642 -3903 7676 -3902
rect 8062 -3902 8146 -3868
rect 8062 -3903 8096 -3902
rect 8482 -3902 8566 -3868
rect 8482 -3903 8516 -3902
rect 8902 -3902 8986 -3868
rect 8902 -3903 8936 -3902
rect 2950 -4272 3248 -3990
rect 5542 -5794 5626 -5760
rect 5542 -5795 5576 -5794
rect 5962 -5794 6046 -5760
rect 5962 -5795 5996 -5794
rect 6382 -5794 6466 -5760
rect 6382 -5800 6416 -5794
rect 6802 -5794 6886 -5760
rect 6802 -5800 6836 -5794
rect 7222 -5794 7306 -5760
rect 7222 -5800 7256 -5794
rect 7642 -5794 7726 -5760
rect 7642 -5800 7676 -5794
rect 8062 -5794 8146 -5760
rect 8062 -5800 8096 -5794
rect 8482 -5794 8566 -5760
rect 8482 -5800 8516 -5794
rect 8902 -5794 8986 -5760
rect 8902 -5800 8936 -5794
rect 5494 -6826 5528 -5850
rect 5590 -6826 5624 -5850
rect 5704 -6826 5738 -5850
rect 5800 -6826 5834 -5850
rect 5914 -6826 5948 -5850
rect 6010 -6826 6044 -5850
rect 6124 -6826 6158 -5850
rect 6220 -6826 6254 -5850
rect 6334 -6826 6368 -5850
rect 6430 -6826 6464 -5850
rect 6544 -6826 6578 -5850
rect 6640 -6826 6674 -5850
rect 6754 -6826 6788 -5850
rect 6850 -6826 6884 -5850
rect 6964 -6826 6998 -5850
rect 7060 -6826 7094 -5850
rect 7174 -6826 7208 -5850
rect 7270 -6826 7304 -5850
rect 7384 -6826 7418 -5850
rect 7480 -6826 7514 -5850
rect 7594 -6826 7628 -5850
rect 7690 -6826 7724 -5850
rect 7804 -6826 7838 -5850
rect 7900 -6826 7934 -5850
rect 8014 -6826 8048 -5850
rect 8110 -6826 8144 -5850
rect 8224 -6826 8258 -5850
rect 8320 -6826 8354 -5850
rect 8434 -6826 8468 -5850
rect 8530 -6826 8564 -5850
rect 8644 -6826 8678 -5850
rect 8740 -6826 8774 -5850
rect 8854 -6826 8888 -5850
rect 8950 -6826 8984 -5850
rect 9064 -6826 9098 -5850
rect 9160 -6826 9194 -5850
rect 5752 -6918 5836 -6884
rect 6172 -6884 6206 -6876
rect 6172 -6918 6256 -6884
rect 6592 -6884 6626 -6876
rect 6592 -6918 6676 -6884
rect 7012 -6884 7046 -6876
rect 7012 -6918 7096 -6884
rect 7432 -6884 7466 -6876
rect 7432 -6918 7516 -6884
rect 7852 -6884 7886 -6876
rect 7852 -6918 7936 -6884
rect 8272 -6884 8306 -6876
rect 8272 -6918 8356 -6884
rect 8692 -6884 8726 -6876
rect 8692 -6918 8776 -6884
rect 9112 -6884 9146 -6876
rect 9112 -6918 9196 -6884
rect 5490 -7104 5590 -7004
rect 5910 -7104 6010 -7004
rect 6330 -7104 6430 -7004
rect 6750 -7104 6850 -7004
rect 7170 -7104 7270 -7004
rect 7590 -7104 7690 -7004
rect 8010 -7104 8110 -7004
rect 8430 -7104 8530 -7004
rect 8850 -7104 8950 -7004
rect 9176 -7104 9276 -7004
<< metal1 >>
rect 10296 13372 10406 13384
rect 10716 13372 10826 13384
rect 11136 13372 11246 13384
rect 11556 13372 11666 13384
rect 11976 13372 12086 13384
rect 12396 13372 12506 13384
rect 12816 13372 12926 13384
rect 13236 13372 13346 13384
rect 13656 13372 13766 13384
rect 14076 13372 14186 13384
rect 14496 13372 14606 13384
rect 14916 13372 15026 13384
rect 15336 13372 15446 13384
rect 15756 13372 15866 13384
rect 16176 13372 16286 13384
rect 16596 13372 16706 13384
rect 17016 13372 17126 13384
rect 17436 13372 17546 13384
rect 17856 13372 17966 13384
rect 18276 13372 18386 13384
rect 18624 13372 18734 13384
rect 10292 13268 10302 13372
rect 10400 13268 10410 13372
rect 10712 13268 10722 13372
rect 10820 13268 10830 13372
rect 11132 13268 11142 13372
rect 11240 13268 11250 13372
rect 11552 13268 11562 13372
rect 11660 13268 11670 13372
rect 11972 13268 11982 13372
rect 12080 13268 12090 13372
rect 12392 13268 12402 13372
rect 12500 13268 12510 13372
rect 12812 13268 12822 13372
rect 12920 13268 12930 13372
rect 13232 13268 13242 13372
rect 13340 13268 13350 13372
rect 13652 13268 13662 13372
rect 13760 13268 13770 13372
rect 14072 13268 14082 13372
rect 14180 13268 14190 13372
rect 14492 13268 14502 13372
rect 14600 13268 14610 13372
rect 14912 13268 14922 13372
rect 15020 13268 15030 13372
rect 15332 13268 15342 13372
rect 15440 13268 15450 13372
rect 15752 13268 15762 13372
rect 15860 13268 15870 13372
rect 16172 13268 16182 13372
rect 16280 13268 16290 13372
rect 16592 13268 16602 13372
rect 16700 13268 16710 13372
rect 17012 13268 17022 13372
rect 17120 13268 17130 13372
rect 17432 13268 17442 13372
rect 17540 13268 17550 13372
rect 17852 13268 17862 13372
rect 17960 13268 17970 13372
rect 18272 13268 18282 13372
rect 18380 13268 18390 13372
rect 18620 13268 18630 13372
rect 18728 13268 18738 13372
rect 10296 13256 10406 13268
rect 10716 13256 10826 13268
rect 11136 13256 11246 13268
rect 11556 13256 11666 13268
rect 11976 13256 12086 13268
rect 12396 13256 12506 13268
rect 12816 13256 12926 13268
rect 13236 13256 13346 13268
rect 13656 13256 13766 13268
rect 14076 13256 14186 13268
rect 14496 13256 14606 13268
rect 14916 13256 15026 13268
rect 15336 13256 15446 13268
rect 15756 13256 15866 13268
rect 16176 13256 16286 13268
rect 16596 13256 16706 13268
rect 17016 13256 17126 13268
rect 17436 13256 17546 13268
rect 17856 13256 17966 13268
rect 18276 13256 18386 13268
rect 18624 13256 18734 13268
rect 9426 13120 18468 13126
rect 9426 13086 10392 13120
rect 10476 13086 10812 13120
rect 10896 13086 11232 13120
rect 11316 13086 11652 13120
rect 11736 13086 12072 13120
rect 12156 13086 12492 13120
rect 12576 13086 12912 13120
rect 12996 13086 13332 13120
rect 13416 13086 13752 13120
rect 13836 13086 14172 13120
rect 14256 13086 14592 13120
rect 14676 13086 15012 13120
rect 15096 13086 15432 13120
rect 15516 13086 15852 13120
rect 15936 13086 16272 13120
rect 16356 13086 16692 13120
rect 16776 13086 17112 13120
rect 17196 13086 17532 13120
rect 17616 13086 17952 13120
rect 18036 13086 18372 13120
rect 18456 13086 18468 13120
rect 9426 13080 18468 13086
rect 9426 12020 9898 13080
rect 10338 13036 10384 13048
rect 10434 13036 10480 13048
rect 10548 13036 10594 13048
rect 10644 13036 10690 13048
rect 10758 13036 10804 13048
rect 10854 13036 10900 13048
rect 10968 13036 11014 13048
rect 11064 13036 11110 13048
rect 11178 13036 11224 13048
rect 11274 13036 11320 13048
rect 11388 13036 11434 13048
rect 11484 13036 11530 13048
rect 11598 13036 11644 13048
rect 11694 13036 11740 13048
rect 11808 13036 11854 13048
rect 11904 13036 11950 13048
rect 12018 13036 12064 13048
rect 12114 13036 12160 13048
rect 12228 13036 12274 13048
rect 12324 13036 12370 13048
rect 12438 13036 12484 13048
rect 12534 13036 12580 13048
rect 12648 13036 12694 13048
rect 12744 13036 12790 13048
rect 12858 13036 12904 13048
rect 12954 13036 13000 13048
rect 13068 13036 13114 13048
rect 13164 13036 13210 13048
rect 13278 13036 13324 13048
rect 13374 13036 13420 13048
rect 13488 13036 13534 13048
rect 13584 13036 13630 13048
rect 13698 13036 13744 13048
rect 13794 13036 13840 13048
rect 13908 13036 13954 13048
rect 14004 13036 14050 13048
rect 14118 13036 14164 13048
rect 14214 13036 14260 13048
rect 14328 13036 14374 13048
rect 14424 13036 14470 13048
rect 14538 13036 14584 13048
rect 14634 13036 14680 13048
rect 14748 13036 14794 13048
rect 14844 13036 14890 13048
rect 14958 13036 15004 13048
rect 15054 13036 15100 13048
rect 15168 13036 15214 13048
rect 15264 13036 15310 13048
rect 15378 13036 15424 13048
rect 15474 13036 15520 13048
rect 15588 13036 15634 13048
rect 15684 13036 15730 13048
rect 15798 13036 15844 13048
rect 15894 13036 15940 13048
rect 16008 13036 16054 13048
rect 16104 13036 16150 13048
rect 16218 13036 16264 13048
rect 16314 13036 16360 13048
rect 16428 13036 16474 13048
rect 16524 13036 16570 13048
rect 16638 13036 16684 13048
rect 16734 13036 16780 13048
rect 16848 13036 16894 13048
rect 16944 13036 16990 13048
rect 17058 13036 17104 13048
rect 17154 13036 17200 13048
rect 17268 13036 17314 13048
rect 17364 13036 17410 13048
rect 17478 13036 17524 13048
rect 17574 13036 17620 13048
rect 17688 13036 17734 13048
rect 17784 13036 17830 13048
rect 17898 13036 17944 13048
rect 17994 13036 18040 13048
rect 18108 13036 18154 13048
rect 18204 13036 18250 13048
rect 18318 13036 18364 13048
rect 18414 13036 18460 13048
rect 18528 13036 18574 13048
rect 18624 13036 18670 13048
rect 10310 12060 10320 13036
rect 10378 12060 10388 13036
rect 10430 12060 10440 13036
rect 10588 12060 10598 13036
rect 10640 12060 10650 13036
rect 10798 12060 10808 13036
rect 10850 12060 10860 13036
rect 11008 12060 11018 13036
rect 11060 12060 11070 13036
rect 11218 12060 11228 13036
rect 11270 12060 11280 13036
rect 11428 12060 11438 13036
rect 11480 12060 11490 13036
rect 11638 12060 11648 13036
rect 11690 12060 11700 13036
rect 11848 12060 11858 13036
rect 11900 12060 11910 13036
rect 12058 12060 12068 13036
rect 12110 12060 12120 13036
rect 12268 12060 12278 13036
rect 12320 12060 12330 13036
rect 12478 12060 12488 13036
rect 12530 12060 12540 13036
rect 12688 12060 12698 13036
rect 12740 12060 12750 13036
rect 12898 12060 12908 13036
rect 12950 12060 12960 13036
rect 13108 12060 13118 13036
rect 13160 12060 13170 13036
rect 13318 12060 13328 13036
rect 13370 12060 13380 13036
rect 13528 12060 13538 13036
rect 13580 12060 13590 13036
rect 13738 12060 13748 13036
rect 13790 12060 13800 13036
rect 13948 12060 13958 13036
rect 14000 12060 14010 13036
rect 14158 12060 14168 13036
rect 14210 12060 14220 13036
rect 14368 12060 14378 13036
rect 14420 12060 14430 13036
rect 14578 12060 14588 13036
rect 14630 12060 14640 13036
rect 14788 12060 14798 13036
rect 14840 12060 14850 13036
rect 14998 12060 15008 13036
rect 15050 12060 15060 13036
rect 15208 12060 15218 13036
rect 15260 12060 15270 13036
rect 15418 12060 15428 13036
rect 15470 12060 15480 13036
rect 15628 12060 15638 13036
rect 15680 12060 15690 13036
rect 15838 12060 15848 13036
rect 15890 12060 15900 13036
rect 16048 12060 16058 13036
rect 16100 12060 16110 13036
rect 16258 12060 16268 13036
rect 16310 12060 16320 13036
rect 16468 12060 16478 13036
rect 16520 12060 16530 13036
rect 16678 12060 16688 13036
rect 16730 12060 16740 13036
rect 16888 12060 16898 13036
rect 16940 12060 16950 13036
rect 17098 12060 17108 13036
rect 17150 12060 17160 13036
rect 17308 12060 17318 13036
rect 17360 12060 17370 13036
rect 17518 12060 17528 13036
rect 17570 12060 17580 13036
rect 17728 12060 17738 13036
rect 17780 12060 17790 13036
rect 17938 12060 17948 13036
rect 17990 12060 18000 13036
rect 18148 12060 18158 13036
rect 18200 12060 18210 13036
rect 18358 12060 18368 13036
rect 18410 12060 18420 13036
rect 18568 12060 18578 13036
rect 18620 12060 18630 13036
rect 18688 12060 18698 13036
rect 10338 12048 10384 12060
rect 10434 12048 10480 12060
rect 10548 12048 10594 12060
rect 10644 12048 10690 12060
rect 10758 12048 10804 12060
rect 10854 12048 10900 12060
rect 10968 12048 11014 12060
rect 11064 12048 11110 12060
rect 11178 12048 11224 12060
rect 11274 12048 11320 12060
rect 11388 12048 11434 12060
rect 11484 12048 11530 12060
rect 11598 12048 11644 12060
rect 11694 12048 11740 12060
rect 11808 12048 11854 12060
rect 11904 12048 11950 12060
rect 12018 12048 12064 12060
rect 12114 12048 12160 12060
rect 12228 12048 12274 12060
rect 12324 12048 12370 12060
rect 12438 12048 12484 12060
rect 12534 12048 12580 12060
rect 12648 12048 12694 12060
rect 12744 12048 12790 12060
rect 12858 12048 12904 12060
rect 12954 12048 13000 12060
rect 13068 12048 13114 12060
rect 13164 12048 13210 12060
rect 13278 12048 13324 12060
rect 13374 12048 13420 12060
rect 13488 12048 13534 12060
rect 13584 12048 13630 12060
rect 13698 12048 13744 12060
rect 13794 12048 13840 12060
rect 13908 12048 13954 12060
rect 14004 12048 14050 12060
rect 14118 12048 14164 12060
rect 14214 12048 14260 12060
rect 14328 12048 14374 12060
rect 14424 12048 14470 12060
rect 14538 12048 14584 12060
rect 14634 12048 14680 12060
rect 14748 12048 14794 12060
rect 14844 12048 14890 12060
rect 14958 12048 15004 12060
rect 15054 12048 15100 12060
rect 15168 12048 15214 12060
rect 15264 12048 15310 12060
rect 15378 12048 15424 12060
rect 15474 12048 15520 12060
rect 15588 12048 15634 12060
rect 15684 12048 15730 12060
rect 15798 12048 15844 12060
rect 15894 12048 15940 12060
rect 16008 12048 16054 12060
rect 16104 12048 16150 12060
rect 16218 12048 16264 12060
rect 16314 12048 16360 12060
rect 16428 12048 16474 12060
rect 16524 12048 16570 12060
rect 16638 12048 16684 12060
rect 16734 12048 16780 12060
rect 16848 12048 16894 12060
rect 16944 12048 16990 12060
rect 17058 12048 17104 12060
rect 17154 12048 17200 12060
rect 17268 12048 17314 12060
rect 17364 12048 17410 12060
rect 17478 12048 17524 12060
rect 17574 12048 17620 12060
rect 17688 12048 17734 12060
rect 17784 12048 17830 12060
rect 17898 12048 17944 12060
rect 17994 12048 18040 12060
rect 18108 12048 18154 12060
rect 18204 12048 18250 12060
rect 18318 12048 18364 12060
rect 18414 12048 18460 12060
rect 18528 12048 18574 12060
rect 18624 12048 18670 12060
rect 9426 12010 18628 12020
rect 9426 11868 10602 12010
rect 10636 11868 11022 12010
rect 11056 11868 11442 12010
rect 11476 11868 11862 12010
rect 11896 11868 12282 12010
rect 12316 11868 12702 12010
rect 12736 11868 13122 12010
rect 13156 11868 13542 12010
rect 13576 11868 13962 12010
rect 13996 11868 14382 12010
rect 14416 11868 14802 12010
rect 14836 11868 15222 12010
rect 15256 11868 15642 12010
rect 15676 11868 16062 12010
rect 16096 11868 16482 12010
rect 16516 11868 16902 12010
rect 16936 11868 17322 12010
rect 17356 11868 17742 12010
rect 17776 11868 18162 12010
rect 18196 11868 18582 12010
rect 18616 11868 18628 12010
rect 9426 11858 18628 11868
rect 9426 10798 9898 11858
rect 10338 11818 10384 11830
rect 10434 11818 10480 11830
rect 10548 11818 10594 11830
rect 10644 11818 10690 11830
rect 10758 11818 10804 11830
rect 10854 11818 10900 11830
rect 10968 11818 11014 11830
rect 11064 11818 11110 11830
rect 11178 11818 11224 11830
rect 11274 11818 11320 11830
rect 11388 11818 11434 11830
rect 11484 11818 11530 11830
rect 11598 11818 11644 11830
rect 11694 11818 11740 11830
rect 11808 11818 11854 11830
rect 11904 11818 11950 11830
rect 12018 11818 12064 11830
rect 12114 11818 12160 11830
rect 12228 11818 12274 11830
rect 12324 11818 12370 11830
rect 12438 11818 12484 11830
rect 12534 11818 12580 11830
rect 12648 11818 12694 11830
rect 12744 11818 12790 11830
rect 12858 11818 12904 11830
rect 12954 11818 13000 11830
rect 13068 11818 13114 11830
rect 13164 11818 13210 11830
rect 13278 11818 13324 11830
rect 13374 11818 13420 11830
rect 13488 11818 13534 11830
rect 13584 11818 13630 11830
rect 13698 11818 13744 11830
rect 13794 11818 13840 11830
rect 13908 11818 13954 11830
rect 14004 11818 14050 11830
rect 14118 11818 14164 11830
rect 14214 11818 14260 11830
rect 14328 11818 14374 11830
rect 14424 11818 14470 11830
rect 14538 11818 14584 11830
rect 14634 11818 14680 11830
rect 14748 11818 14794 11830
rect 14844 11818 14890 11830
rect 14958 11818 15004 11830
rect 15054 11818 15100 11830
rect 15168 11818 15214 11830
rect 15264 11818 15310 11830
rect 15378 11818 15424 11830
rect 15474 11818 15520 11830
rect 15588 11818 15634 11830
rect 15684 11818 15730 11830
rect 15798 11818 15844 11830
rect 15894 11818 15940 11830
rect 16008 11818 16054 11830
rect 16104 11818 16150 11830
rect 16218 11818 16264 11830
rect 16314 11818 16360 11830
rect 16428 11818 16474 11830
rect 16524 11818 16570 11830
rect 16638 11818 16684 11830
rect 16734 11818 16780 11830
rect 16848 11818 16894 11830
rect 16944 11818 16990 11830
rect 17058 11818 17104 11830
rect 17154 11818 17200 11830
rect 17268 11818 17314 11830
rect 17364 11818 17410 11830
rect 17478 11818 17524 11830
rect 17574 11818 17620 11830
rect 17688 11818 17734 11830
rect 17784 11818 17830 11830
rect 17898 11818 17944 11830
rect 17994 11818 18040 11830
rect 18108 11818 18154 11830
rect 18204 11818 18250 11830
rect 18318 11818 18364 11830
rect 18414 11818 18460 11830
rect 18528 11818 18574 11830
rect 18624 11818 18670 11830
rect 10310 10842 10320 11818
rect 10378 10842 10388 11818
rect 10430 10842 10440 11818
rect 10588 10842 10598 11818
rect 10640 10842 10650 11818
rect 10798 10842 10808 11818
rect 10850 10842 10860 11818
rect 11008 10842 11018 11818
rect 11060 10842 11070 11818
rect 11218 10842 11228 11818
rect 11270 10842 11280 11818
rect 11428 10842 11438 11818
rect 11480 10842 11490 11818
rect 11638 10842 11648 11818
rect 11690 10842 11700 11818
rect 11848 10842 11858 11818
rect 11900 10842 11910 11818
rect 12058 10842 12068 11818
rect 12110 10842 12120 11818
rect 12268 10842 12278 11818
rect 12320 10842 12330 11818
rect 12478 10842 12488 11818
rect 12530 10842 12540 11818
rect 12688 10842 12698 11818
rect 12740 10842 12750 11818
rect 12898 10842 12908 11818
rect 12950 10842 12960 11818
rect 13108 10842 13118 11818
rect 13160 10842 13170 11818
rect 13318 10842 13328 11818
rect 13370 10842 13380 11818
rect 13528 10842 13538 11818
rect 13580 10842 13590 11818
rect 13738 10842 13748 11818
rect 13790 10842 13800 11818
rect 13948 10842 13958 11818
rect 14000 10842 14010 11818
rect 14158 10842 14168 11818
rect 14210 10842 14220 11818
rect 14368 10842 14378 11818
rect 14420 10842 14430 11818
rect 14578 10842 14588 11818
rect 14630 10842 14640 11818
rect 14788 10842 14798 11818
rect 14840 10842 14850 11818
rect 14998 10842 15008 11818
rect 15050 10842 15060 11818
rect 15208 10842 15218 11818
rect 15260 10842 15270 11818
rect 15418 10842 15428 11818
rect 15470 10842 15480 11818
rect 15628 10842 15638 11818
rect 15680 10842 15690 11818
rect 15838 10842 15848 11818
rect 15890 10842 15900 11818
rect 16048 10842 16058 11818
rect 16100 10842 16110 11818
rect 16258 10842 16268 11818
rect 16310 10842 16320 11818
rect 16468 10842 16478 11818
rect 16520 10842 16530 11818
rect 16678 10842 16688 11818
rect 16730 10842 16740 11818
rect 16888 10842 16898 11818
rect 16940 10842 16950 11818
rect 17098 10842 17108 11818
rect 17150 10842 17160 11818
rect 17308 10842 17318 11818
rect 17360 10842 17370 11818
rect 17518 10842 17528 11818
rect 17570 10842 17580 11818
rect 17728 10842 17738 11818
rect 17780 10842 17790 11818
rect 17938 10842 17948 11818
rect 17990 10842 18000 11818
rect 18148 10842 18158 11818
rect 18200 10842 18210 11818
rect 18358 10842 18368 11818
rect 18410 10842 18420 11818
rect 18568 10842 18578 11818
rect 18620 10842 18630 11818
rect 18688 10842 18698 11818
rect 10338 10830 10384 10842
rect 10434 10830 10480 10842
rect 10548 10830 10594 10842
rect 10644 10830 10690 10842
rect 10758 10830 10804 10842
rect 10854 10830 10900 10842
rect 10968 10830 11014 10842
rect 11064 10830 11110 10842
rect 11178 10830 11224 10842
rect 11274 10830 11320 10842
rect 11388 10830 11434 10842
rect 11484 10830 11530 10842
rect 11598 10830 11644 10842
rect 11694 10830 11740 10842
rect 11808 10830 11854 10842
rect 11904 10830 11950 10842
rect 12018 10830 12064 10842
rect 12114 10830 12160 10842
rect 12228 10830 12274 10842
rect 12324 10830 12370 10842
rect 12438 10830 12484 10842
rect 12534 10830 12580 10842
rect 12648 10830 12694 10842
rect 12744 10830 12790 10842
rect 12858 10830 12904 10842
rect 12954 10830 13000 10842
rect 13068 10830 13114 10842
rect 13164 10830 13210 10842
rect 13278 10830 13324 10842
rect 13374 10830 13420 10842
rect 13488 10830 13534 10842
rect 13584 10830 13630 10842
rect 13698 10830 13744 10842
rect 13794 10830 13840 10842
rect 13908 10830 13954 10842
rect 14004 10830 14050 10842
rect 14118 10830 14164 10842
rect 14214 10830 14260 10842
rect 14328 10830 14374 10842
rect 14424 10830 14470 10842
rect 14538 10830 14584 10842
rect 14634 10830 14680 10842
rect 14748 10830 14794 10842
rect 14844 10830 14890 10842
rect 14958 10830 15004 10842
rect 15054 10830 15100 10842
rect 15168 10830 15214 10842
rect 15264 10830 15310 10842
rect 15378 10830 15424 10842
rect 15474 10830 15520 10842
rect 15588 10830 15634 10842
rect 15684 10830 15730 10842
rect 15798 10830 15844 10842
rect 15894 10830 15940 10842
rect 16008 10830 16054 10842
rect 16104 10830 16150 10842
rect 16218 10830 16264 10842
rect 16314 10830 16360 10842
rect 16428 10830 16474 10842
rect 16524 10830 16570 10842
rect 16638 10830 16684 10842
rect 16734 10830 16780 10842
rect 16848 10830 16894 10842
rect 16944 10830 16990 10842
rect 17058 10830 17104 10842
rect 17154 10830 17200 10842
rect 17268 10830 17314 10842
rect 17364 10830 17410 10842
rect 17478 10830 17524 10842
rect 17574 10830 17620 10842
rect 17688 10830 17734 10842
rect 17784 10830 17830 10842
rect 17898 10830 17944 10842
rect 17994 10830 18040 10842
rect 18108 10830 18154 10842
rect 18204 10830 18250 10842
rect 18318 10830 18364 10842
rect 18414 10830 18460 10842
rect 18528 10830 18574 10842
rect 18624 10830 18670 10842
rect 9426 10792 18468 10798
rect 9426 10758 10392 10792
rect 10476 10758 10812 10792
rect 10896 10758 11232 10792
rect 11316 10758 11652 10792
rect 11736 10758 12072 10792
rect 12156 10758 12492 10792
rect 12576 10758 12912 10792
rect 12996 10758 13332 10792
rect 13416 10758 13752 10792
rect 13836 10758 14172 10792
rect 14256 10758 14592 10792
rect 14676 10758 15012 10792
rect 15096 10758 15432 10792
rect 15516 10758 15852 10792
rect 15936 10758 16272 10792
rect 16356 10758 16692 10792
rect 16776 10758 17112 10792
rect 17196 10758 17532 10792
rect 17616 10758 17952 10792
rect 18036 10758 18372 10792
rect 18456 10758 18468 10792
rect 9426 10752 18468 10758
rect 9426 7908 9898 10752
rect 9426 7901 18468 7908
rect 9426 7866 10392 7901
rect 10426 7900 10812 7901
rect 10846 7900 11232 7901
rect 11266 7900 11652 7901
rect 11686 7900 12072 7901
rect 12106 7900 12492 7901
rect 12526 7900 12912 7901
rect 12946 7900 13332 7901
rect 13366 7900 13752 7901
rect 13786 7900 14172 7901
rect 14206 7900 14592 7901
rect 14626 7900 15012 7901
rect 15046 7900 15432 7901
rect 15466 7900 15852 7901
rect 15886 7900 16272 7901
rect 16306 7900 16692 7901
rect 16726 7900 17112 7901
rect 17146 7900 17532 7901
rect 17566 7900 17952 7901
rect 17986 7900 18372 7901
rect 18406 7900 18468 7901
rect 10476 7866 10812 7900
rect 10896 7866 11232 7900
rect 11316 7866 11652 7900
rect 11736 7866 12072 7900
rect 12156 7866 12492 7900
rect 12576 7866 12912 7900
rect 12996 7866 13332 7900
rect 13416 7866 13752 7900
rect 13836 7866 14172 7900
rect 14256 7866 14592 7900
rect 14676 7866 15012 7900
rect 15096 7866 15432 7900
rect 15516 7866 15852 7900
rect 15936 7866 16272 7900
rect 16356 7866 16692 7900
rect 16776 7866 17112 7900
rect 17196 7866 17532 7900
rect 17616 7866 17952 7900
rect 18036 7866 18372 7900
rect 18456 7866 18468 7900
rect 9426 7858 18468 7866
rect 5478 7230 5602 7236
rect 5478 7130 5490 7230
rect 5590 7130 5602 7230
rect 5478 7124 5602 7130
rect 5898 7230 6022 7236
rect 5898 7130 5910 7230
rect 6010 7130 6022 7230
rect 5898 7124 6022 7130
rect 6318 7230 6442 7236
rect 6318 7130 6330 7230
rect 6430 7130 6442 7230
rect 6318 7124 6442 7130
rect 6738 7230 6862 7236
rect 6738 7130 6750 7230
rect 6850 7130 6862 7230
rect 6738 7124 6862 7130
rect 7158 7230 7282 7236
rect 7158 7130 7170 7230
rect 7270 7130 7282 7230
rect 7158 7124 7282 7130
rect 7578 7230 7702 7236
rect 7578 7130 7590 7230
rect 7690 7130 7702 7230
rect 7578 7124 7702 7130
rect 7998 7230 8122 7236
rect 7998 7130 8010 7230
rect 8110 7130 8122 7230
rect 7998 7124 8122 7130
rect 8418 7230 8542 7236
rect 8418 7130 8430 7230
rect 8530 7130 8542 7230
rect 8418 7124 8542 7130
rect 8838 7230 8962 7236
rect 8838 7130 8850 7230
rect 8950 7130 8962 7230
rect 8838 7124 8962 7130
rect 9164 7230 9288 7236
rect 9164 7130 9176 7230
rect 9276 7130 9288 7230
rect 9164 7124 9288 7130
rect 5052 7044 9212 7052
rect 5052 7010 5752 7044
rect 5836 7010 6172 7044
rect 6256 7010 6592 7044
rect 6676 7010 7012 7044
rect 7096 7010 7432 7044
rect 7516 7010 7852 7044
rect 7936 7010 8272 7044
rect 8356 7010 8692 7044
rect 8776 7010 9112 7044
rect 9196 7010 9212 7044
rect 5052 7002 6172 7010
rect 6206 7002 6592 7010
rect 6626 7002 7012 7010
rect 7046 7002 7432 7010
rect 7466 7002 7852 7010
rect 7886 7002 8272 7010
rect 8306 7002 8692 7010
rect 8726 7002 9112 7010
rect 9146 7002 9212 7010
rect 5052 6996 9212 7002
rect 5052 5932 5238 6996
rect 5488 6952 5534 6964
rect 5584 6952 5630 6964
rect 5698 6952 5744 6964
rect 5794 6952 5840 6964
rect 5908 6952 5954 6964
rect 6004 6952 6050 6964
rect 6118 6952 6164 6964
rect 6214 6952 6260 6964
rect 6328 6952 6374 6964
rect 6424 6952 6470 6964
rect 6538 6952 6584 6964
rect 6634 6952 6680 6964
rect 6748 6952 6794 6964
rect 6844 6952 6890 6964
rect 6958 6952 7004 6964
rect 7054 6952 7100 6964
rect 7168 6952 7214 6964
rect 7264 6952 7310 6964
rect 7378 6952 7424 6964
rect 7474 6952 7520 6964
rect 7588 6952 7634 6964
rect 7684 6952 7730 6964
rect 7798 6952 7844 6964
rect 7894 6952 7940 6964
rect 8008 6952 8054 6964
rect 8104 6952 8150 6964
rect 8218 6952 8264 6964
rect 8314 6952 8360 6964
rect 8428 6952 8474 6964
rect 8524 6952 8570 6964
rect 8638 6952 8684 6964
rect 8734 6952 8780 6964
rect 8848 6952 8894 6964
rect 8944 6952 8990 6964
rect 9058 6952 9104 6964
rect 9154 6952 9200 6964
rect 5460 5976 5470 6952
rect 5528 5976 5538 6952
rect 5580 5976 5590 6952
rect 5738 5976 5748 6952
rect 5790 5976 5800 6952
rect 5948 5976 5958 6952
rect 6000 5976 6010 6952
rect 6158 5976 6168 6952
rect 6210 5976 6220 6952
rect 6368 5976 6378 6952
rect 6420 5976 6430 6952
rect 6578 5976 6588 6952
rect 6630 5976 6640 6952
rect 6788 5976 6798 6952
rect 6840 5976 6850 6952
rect 6998 5976 7008 6952
rect 7050 5976 7060 6952
rect 7208 5976 7218 6952
rect 7260 5976 7270 6952
rect 7418 5976 7428 6952
rect 7470 5976 7480 6952
rect 7628 5976 7638 6952
rect 7680 5976 7690 6952
rect 7838 5976 7848 6952
rect 7890 5976 7900 6952
rect 8048 5976 8058 6952
rect 8100 5976 8110 6952
rect 8258 5976 8268 6952
rect 8310 5976 8320 6952
rect 8468 5976 8478 6952
rect 8520 5976 8530 6952
rect 8678 5976 8688 6952
rect 8730 5976 8740 6952
rect 8888 5976 8898 6952
rect 8940 5976 8950 6952
rect 9098 5976 9108 6952
rect 9150 5976 9160 6952
rect 9218 5976 9228 6952
rect 9426 6780 9898 7858
rect 10338 7808 10384 7820
rect 10434 7808 10480 7820
rect 10548 7808 10594 7820
rect 10644 7808 10690 7820
rect 10758 7808 10804 7820
rect 10854 7808 10900 7820
rect 10968 7808 11014 7820
rect 11064 7808 11110 7820
rect 11178 7808 11224 7820
rect 11274 7808 11320 7820
rect 11388 7808 11434 7820
rect 11484 7808 11530 7820
rect 11598 7808 11644 7820
rect 11694 7808 11740 7820
rect 11808 7808 11854 7820
rect 11904 7808 11950 7820
rect 12018 7808 12064 7820
rect 12114 7808 12160 7820
rect 12228 7808 12274 7820
rect 12324 7808 12370 7820
rect 12438 7808 12484 7820
rect 12534 7808 12580 7820
rect 12648 7808 12694 7820
rect 12744 7808 12790 7820
rect 12858 7808 12904 7820
rect 12954 7808 13000 7820
rect 13068 7808 13114 7820
rect 13164 7808 13210 7820
rect 13278 7808 13324 7820
rect 13374 7808 13420 7820
rect 13488 7808 13534 7820
rect 13584 7808 13630 7820
rect 13698 7808 13744 7820
rect 13794 7808 13840 7820
rect 13908 7808 13954 7820
rect 14004 7808 14050 7820
rect 14118 7808 14164 7820
rect 14214 7808 14260 7820
rect 14328 7808 14374 7820
rect 14424 7808 14470 7820
rect 14538 7808 14584 7820
rect 14634 7808 14680 7820
rect 14748 7808 14794 7820
rect 14844 7808 14890 7820
rect 14958 7808 15004 7820
rect 15054 7808 15100 7820
rect 15168 7808 15214 7820
rect 15264 7808 15310 7820
rect 15378 7808 15424 7820
rect 15474 7808 15520 7820
rect 15588 7808 15634 7820
rect 15684 7808 15730 7820
rect 15798 7808 15844 7820
rect 15894 7808 15940 7820
rect 16008 7808 16054 7820
rect 16104 7808 16150 7820
rect 16218 7808 16264 7820
rect 16314 7808 16360 7820
rect 16428 7808 16474 7820
rect 16524 7808 16570 7820
rect 16638 7808 16684 7820
rect 16734 7808 16780 7820
rect 16848 7808 16894 7820
rect 16944 7808 16990 7820
rect 17058 7808 17104 7820
rect 17154 7808 17200 7820
rect 17268 7808 17314 7820
rect 17364 7808 17410 7820
rect 17478 7808 17524 7820
rect 17574 7808 17620 7820
rect 17688 7808 17734 7820
rect 17784 7808 17830 7820
rect 17898 7808 17944 7820
rect 17994 7808 18040 7820
rect 18108 7808 18154 7820
rect 18204 7808 18250 7820
rect 18318 7808 18364 7820
rect 18414 7808 18460 7820
rect 18528 7808 18574 7820
rect 18624 7808 18670 7820
rect 10310 6832 10320 7808
rect 10378 6832 10388 7808
rect 10430 6832 10440 7808
rect 10588 6832 10598 7808
rect 10640 6832 10650 7808
rect 10798 6832 10808 7808
rect 10850 6832 10860 7808
rect 11008 6832 11018 7808
rect 11060 6832 11070 7808
rect 11218 6832 11228 7808
rect 11270 6832 11280 7808
rect 11428 6832 11438 7808
rect 11480 6832 11490 7808
rect 11638 6832 11648 7808
rect 11690 6832 11700 7808
rect 11848 6832 11858 7808
rect 11900 6832 11910 7808
rect 12058 6832 12068 7808
rect 12110 6832 12120 7808
rect 12268 6832 12278 7808
rect 12320 6832 12330 7808
rect 12478 6832 12488 7808
rect 12530 6832 12540 7808
rect 12688 6832 12698 7808
rect 12740 6832 12750 7808
rect 12898 6832 12908 7808
rect 12950 6832 12960 7808
rect 13108 6832 13118 7808
rect 13160 6832 13170 7808
rect 13318 6832 13328 7808
rect 13370 6832 13380 7808
rect 13528 6832 13538 7808
rect 13580 6832 13590 7808
rect 13738 6832 13748 7808
rect 13790 6832 13800 7808
rect 13948 6832 13958 7808
rect 14000 6832 14010 7808
rect 14158 6832 14168 7808
rect 14210 6832 14220 7808
rect 14368 6832 14378 7808
rect 14420 6832 14430 7808
rect 14578 6832 14588 7808
rect 14630 6832 14640 7808
rect 14788 6832 14798 7808
rect 14840 6832 14850 7808
rect 14998 6832 15008 7808
rect 15050 6832 15060 7808
rect 15208 6832 15218 7808
rect 15260 6832 15270 7808
rect 15418 6832 15428 7808
rect 15470 6832 15480 7808
rect 15628 6832 15638 7808
rect 15680 6832 15690 7808
rect 15838 6832 15848 7808
rect 15890 6832 15900 7808
rect 16048 6832 16058 7808
rect 16100 6832 16110 7808
rect 16258 6832 16268 7808
rect 16310 6832 16320 7808
rect 16468 6832 16478 7808
rect 16520 6832 16530 7808
rect 16678 6832 16688 7808
rect 16730 6832 16740 7808
rect 16888 6832 16898 7808
rect 16940 6832 16950 7808
rect 17098 6832 17108 7808
rect 17150 6832 17160 7808
rect 17308 6832 17318 7808
rect 17360 6832 17370 7808
rect 17518 6832 17528 7808
rect 17570 6832 17580 7808
rect 17728 6832 17738 7808
rect 17780 6832 17790 7808
rect 17938 6832 17948 7808
rect 17990 6832 18000 7808
rect 18148 6832 18158 7808
rect 18200 6832 18210 7808
rect 18358 6832 18368 7808
rect 18410 6832 18420 7808
rect 18568 6832 18578 7808
rect 18620 6832 18630 7808
rect 18688 6832 18698 7808
rect 10338 6820 10384 6832
rect 10434 6820 10480 6832
rect 10548 6820 10594 6832
rect 10644 6820 10690 6832
rect 10758 6820 10804 6832
rect 10854 6820 10900 6832
rect 10968 6820 11014 6832
rect 11064 6820 11110 6832
rect 11178 6820 11224 6832
rect 11274 6820 11320 6832
rect 11388 6820 11434 6832
rect 11484 6820 11530 6832
rect 11598 6820 11644 6832
rect 11694 6820 11740 6832
rect 11808 6820 11854 6832
rect 11904 6820 11950 6832
rect 12018 6820 12064 6832
rect 12114 6820 12160 6832
rect 12228 6820 12274 6832
rect 12324 6820 12370 6832
rect 12438 6820 12484 6832
rect 12534 6820 12580 6832
rect 12648 6820 12694 6832
rect 12744 6820 12790 6832
rect 12858 6820 12904 6832
rect 12954 6820 13000 6832
rect 13068 6820 13114 6832
rect 13164 6820 13210 6832
rect 13278 6820 13324 6832
rect 13374 6820 13420 6832
rect 13488 6820 13534 6832
rect 13584 6820 13630 6832
rect 13698 6820 13744 6832
rect 13794 6820 13840 6832
rect 13908 6820 13954 6832
rect 14004 6820 14050 6832
rect 14118 6820 14164 6832
rect 14214 6820 14260 6832
rect 14328 6820 14374 6832
rect 14424 6820 14470 6832
rect 14538 6820 14584 6832
rect 14634 6820 14680 6832
rect 14748 6820 14794 6832
rect 14844 6820 14890 6832
rect 14958 6820 15004 6832
rect 15054 6820 15100 6832
rect 15168 6820 15214 6832
rect 15264 6820 15310 6832
rect 15378 6820 15424 6832
rect 15474 6820 15520 6832
rect 15588 6820 15634 6832
rect 15684 6820 15730 6832
rect 15798 6820 15844 6832
rect 15894 6820 15940 6832
rect 16008 6820 16054 6832
rect 16104 6820 16150 6832
rect 16218 6820 16264 6832
rect 16314 6820 16360 6832
rect 16428 6820 16474 6832
rect 16524 6820 16570 6832
rect 16638 6820 16684 6832
rect 16734 6820 16780 6832
rect 16848 6820 16894 6832
rect 16944 6820 16990 6832
rect 17058 6820 17104 6832
rect 17154 6820 17200 6832
rect 17268 6820 17314 6832
rect 17364 6820 17410 6832
rect 17478 6820 17524 6832
rect 17574 6820 17620 6832
rect 17688 6820 17734 6832
rect 17784 6820 17830 6832
rect 17898 6820 17944 6832
rect 17994 6820 18040 6832
rect 18108 6820 18154 6832
rect 18204 6820 18250 6832
rect 18318 6820 18364 6832
rect 18414 6820 18460 6832
rect 18528 6820 18574 6832
rect 18624 6820 18670 6832
rect 9426 6773 18628 6780
rect 9426 6631 10602 6773
rect 10636 6631 11022 6773
rect 11056 6631 11442 6773
rect 11476 6631 11862 6773
rect 11896 6631 12282 6773
rect 12316 6631 12702 6773
rect 12736 6631 13122 6773
rect 13156 6631 13542 6773
rect 13576 6631 13962 6773
rect 13996 6631 14382 6773
rect 14416 6631 14802 6773
rect 14836 6631 15222 6773
rect 15256 6631 15642 6773
rect 15676 6631 16062 6773
rect 16096 6631 16482 6773
rect 16516 6631 16902 6773
rect 16936 6631 17322 6773
rect 17356 6631 17742 6773
rect 17776 6631 18162 6773
rect 18196 6631 18582 6773
rect 18616 6631 18628 6773
rect 9426 6624 18628 6631
rect 9426 5996 9898 6624
rect 10338 6572 10384 6584
rect 10434 6572 10480 6584
rect 10548 6572 10594 6584
rect 10644 6572 10690 6584
rect 10758 6572 10804 6584
rect 10854 6572 10900 6584
rect 10968 6572 11014 6584
rect 11064 6572 11110 6584
rect 11178 6572 11224 6584
rect 11274 6572 11320 6584
rect 11388 6572 11434 6584
rect 11484 6572 11530 6584
rect 11598 6572 11644 6584
rect 11694 6572 11740 6584
rect 11808 6572 11854 6584
rect 11904 6572 11950 6584
rect 12018 6572 12064 6584
rect 12114 6572 12160 6584
rect 12228 6572 12274 6584
rect 12324 6572 12370 6584
rect 12438 6572 12484 6584
rect 12534 6572 12580 6584
rect 12648 6572 12694 6584
rect 12744 6572 12790 6584
rect 12858 6572 12904 6584
rect 12954 6572 13000 6584
rect 13068 6572 13114 6584
rect 13164 6572 13210 6584
rect 13278 6572 13324 6584
rect 13374 6572 13420 6584
rect 13488 6572 13534 6584
rect 13584 6572 13630 6584
rect 13698 6572 13744 6584
rect 13794 6572 13840 6584
rect 13908 6572 13954 6584
rect 14004 6572 14050 6584
rect 14118 6572 14164 6584
rect 14214 6572 14260 6584
rect 14328 6572 14374 6584
rect 14424 6572 14470 6584
rect 14538 6572 14584 6584
rect 14634 6572 14680 6584
rect 14748 6572 14794 6584
rect 14844 6572 14890 6584
rect 14958 6572 15004 6584
rect 15054 6572 15100 6584
rect 15168 6572 15214 6584
rect 15264 6572 15310 6584
rect 15378 6572 15424 6584
rect 15474 6572 15520 6584
rect 15588 6572 15634 6584
rect 15684 6572 15730 6584
rect 15798 6572 15844 6584
rect 15894 6572 15940 6584
rect 16008 6572 16054 6584
rect 16104 6572 16150 6584
rect 16218 6572 16264 6584
rect 16314 6572 16360 6584
rect 16428 6572 16474 6584
rect 16524 6572 16570 6584
rect 16638 6572 16684 6584
rect 16734 6572 16780 6584
rect 16848 6572 16894 6584
rect 16944 6572 16990 6584
rect 17058 6572 17104 6584
rect 17154 6572 17200 6584
rect 17268 6572 17314 6584
rect 17364 6572 17410 6584
rect 17478 6572 17524 6584
rect 17574 6572 17620 6584
rect 17688 6572 17734 6584
rect 17784 6572 17830 6584
rect 17898 6572 17944 6584
rect 17994 6572 18040 6584
rect 18108 6572 18154 6584
rect 18204 6572 18250 6584
rect 18318 6572 18364 6584
rect 18414 6572 18460 6584
rect 18528 6572 18574 6584
rect 18624 6572 18670 6584
rect 5488 5964 5534 5976
rect 5584 5964 5630 5976
rect 5698 5964 5744 5976
rect 5794 5964 5840 5976
rect 5908 5964 5954 5976
rect 6004 5964 6050 5976
rect 6118 5964 6164 5976
rect 6214 5964 6260 5976
rect 6328 5964 6374 5976
rect 6424 5964 6470 5976
rect 6538 5964 6584 5976
rect 6634 5964 6680 5976
rect 6748 5964 6794 5976
rect 6844 5964 6890 5976
rect 6958 5964 7004 5976
rect 7054 5964 7100 5976
rect 7168 5964 7214 5976
rect 7264 5964 7310 5976
rect 7378 5964 7424 5976
rect 7474 5964 7520 5976
rect 7588 5964 7634 5976
rect 7684 5964 7730 5976
rect 7798 5964 7844 5976
rect 7894 5964 7940 5976
rect 8008 5964 8054 5976
rect 8104 5964 8150 5976
rect 8218 5964 8264 5976
rect 8314 5964 8360 5976
rect 8428 5964 8474 5976
rect 8524 5964 8570 5976
rect 8638 5964 8684 5976
rect 8734 5964 8780 5976
rect 8848 5964 8894 5976
rect 8944 5964 8990 5976
rect 9058 5964 9104 5976
rect 9154 5964 9200 5976
rect 5052 5926 9098 5932
rect 5052 5921 6382 5926
rect 5052 5886 5542 5921
rect 5576 5920 5962 5921
rect 5996 5920 6382 5921
rect 6416 5920 6802 5926
rect 6836 5920 7222 5926
rect 7256 5920 7642 5926
rect 7676 5920 8062 5926
rect 8096 5920 8482 5926
rect 8516 5920 8902 5926
rect 8936 5920 9098 5926
rect 5626 5886 5962 5920
rect 6046 5886 6382 5920
rect 6466 5886 6802 5920
rect 6886 5886 7222 5920
rect 7306 5886 7642 5920
rect 7726 5886 8062 5920
rect 8146 5886 8482 5920
rect 8566 5886 8902 5920
rect 8986 5886 9098 5920
rect 5052 5872 9098 5886
rect 2938 5798 3260 5804
rect 2938 5516 2950 5798
rect 3248 5516 3260 5798
rect 2938 5510 3260 5516
rect 5052 5436 5238 5872
rect 5052 5429 9098 5436
rect 2784 5421 4304 5428
rect 2784 5386 3788 5421
rect 3822 5420 4208 5421
rect 4242 5420 4304 5421
rect 3872 5386 4208 5420
rect 4292 5386 4304 5420
rect 2784 5372 4304 5386
rect 5052 5394 5542 5429
rect 5576 5428 5962 5429
rect 5996 5428 6382 5429
rect 6416 5428 6802 5429
rect 6836 5428 7222 5429
rect 7256 5428 7642 5429
rect 7676 5428 8062 5429
rect 8096 5428 8482 5429
rect 8516 5428 8902 5429
rect 8936 5428 9098 5429
rect 5626 5394 5962 5428
rect 6046 5394 6382 5428
rect 6466 5394 6802 5428
rect 6886 5394 7222 5428
rect 7306 5394 7642 5428
rect 7726 5394 8062 5428
rect 8146 5394 8482 5428
rect 8566 5394 8902 5428
rect 8986 5394 9098 5428
rect 5052 5386 9098 5394
rect 2580 5328 2626 5340
rect 2668 5328 2714 5340
rect 2556 4352 2566 5328
rect 2620 4352 2630 5328
rect 2664 4352 2674 5328
rect 2728 4352 2738 5328
rect 2784 4404 2898 5372
rect 3524 5328 3570 5340
rect 3620 5328 3666 5340
rect 3734 5328 3780 5340
rect 3830 5328 3876 5340
rect 3944 5328 3990 5340
rect 4040 5328 4086 5340
rect 4154 5328 4200 5340
rect 4250 5328 4296 5340
rect 2580 4340 2626 4352
rect 2668 4340 2714 4352
rect 2618 4302 2676 4308
rect 2618 4250 2630 4302
rect 2228 4202 2630 4250
rect 2228 3072 2322 4202
rect 2618 4159 2630 4202
rect 2664 4159 2676 4302
rect 2784 4256 2794 4404
rect 2936 4274 2946 4404
rect 3500 4352 3510 5328
rect 3564 4352 3574 5328
rect 3616 4352 3626 5328
rect 3774 4352 3784 5328
rect 3826 4352 3836 5328
rect 3984 4352 3994 5328
rect 4036 4352 4046 5328
rect 4194 4352 4204 5328
rect 4246 4352 4256 5328
rect 4310 4352 4320 5328
rect 4716 4500 4726 4764
rect 5008 4736 5018 4764
rect 5052 4736 5238 5386
rect 9316 5378 9326 5996
rect 9936 5544 9946 5996
rect 10310 5596 10320 6572
rect 10378 5596 10388 6572
rect 10430 5596 10440 6572
rect 10588 5596 10598 6572
rect 10640 5596 10650 6572
rect 10798 5596 10808 6572
rect 10850 5596 10860 6572
rect 11008 5596 11018 6572
rect 11060 5596 11070 6572
rect 11218 5596 11228 6572
rect 11270 5596 11280 6572
rect 11428 5596 11438 6572
rect 11480 5596 11490 6572
rect 11638 5596 11648 6572
rect 11690 5596 11700 6572
rect 11848 5596 11858 6572
rect 11900 5596 11910 6572
rect 12058 5596 12068 6572
rect 12110 5596 12120 6572
rect 12268 5596 12278 6572
rect 12320 5596 12330 6572
rect 12478 5596 12488 6572
rect 12530 5596 12540 6572
rect 12688 5596 12698 6572
rect 12740 5596 12750 6572
rect 12898 5596 12908 6572
rect 12950 5596 12960 6572
rect 13108 5596 13118 6572
rect 13160 5596 13170 6572
rect 13318 5596 13328 6572
rect 13370 5596 13380 6572
rect 13528 5596 13538 6572
rect 13580 5596 13590 6572
rect 13738 5596 13748 6572
rect 13790 5596 13800 6572
rect 13948 5596 13958 6572
rect 14000 5596 14010 6572
rect 14158 5596 14168 6572
rect 14210 5596 14220 6572
rect 14368 5596 14378 6572
rect 14420 5596 14430 6572
rect 14578 5596 14588 6572
rect 14630 5596 14640 6572
rect 14788 5596 14798 6572
rect 14840 5596 14850 6572
rect 14998 5596 15008 6572
rect 15050 5596 15060 6572
rect 15208 5596 15218 6572
rect 15260 5596 15270 6572
rect 15418 5596 15428 6572
rect 15470 5596 15480 6572
rect 15628 5596 15638 6572
rect 15680 5596 15690 6572
rect 15838 5596 15848 6572
rect 15890 5596 15900 6572
rect 16048 5596 16058 6572
rect 16100 5596 16110 6572
rect 16258 5596 16268 6572
rect 16310 5596 16320 6572
rect 16468 5596 16478 6572
rect 16520 5596 16530 6572
rect 16678 5596 16688 6572
rect 16730 5596 16740 6572
rect 16888 5596 16898 6572
rect 16940 5596 16950 6572
rect 17098 5596 17108 6572
rect 17150 5596 17160 6572
rect 17308 5596 17318 6572
rect 17360 5596 17370 6572
rect 17518 5596 17528 6572
rect 17570 5596 17580 6572
rect 17728 5596 17738 6572
rect 17780 5596 17790 6572
rect 17938 5596 17948 6572
rect 17990 5596 18000 6572
rect 18148 5596 18158 6572
rect 18200 5596 18210 6572
rect 18358 5596 18368 6572
rect 18410 5596 18420 6572
rect 18568 5596 18578 6572
rect 18620 5596 18630 6572
rect 18688 5596 18698 6572
rect 10338 5584 10384 5596
rect 10434 5584 10480 5596
rect 10548 5584 10594 5596
rect 10644 5584 10690 5596
rect 10758 5584 10804 5596
rect 10854 5584 10900 5596
rect 10968 5584 11014 5596
rect 11064 5584 11110 5596
rect 11178 5584 11224 5596
rect 11274 5584 11320 5596
rect 11388 5584 11434 5596
rect 11484 5584 11530 5596
rect 11598 5584 11644 5596
rect 11694 5584 11740 5596
rect 11808 5584 11854 5596
rect 11904 5584 11950 5596
rect 12018 5584 12064 5596
rect 12114 5584 12160 5596
rect 12228 5584 12274 5596
rect 12324 5584 12370 5596
rect 12438 5584 12484 5596
rect 12534 5584 12580 5596
rect 12648 5584 12694 5596
rect 12744 5584 12790 5596
rect 12858 5584 12904 5596
rect 12954 5584 13000 5596
rect 13068 5584 13114 5596
rect 13164 5584 13210 5596
rect 13278 5584 13324 5596
rect 13374 5584 13420 5596
rect 13488 5584 13534 5596
rect 13584 5584 13630 5596
rect 13698 5584 13744 5596
rect 13794 5584 13840 5596
rect 13908 5584 13954 5596
rect 14004 5584 14050 5596
rect 14118 5584 14164 5596
rect 14214 5584 14260 5596
rect 14328 5584 14374 5596
rect 14424 5584 14470 5596
rect 14538 5584 14584 5596
rect 14634 5584 14680 5596
rect 14748 5584 14794 5596
rect 14844 5584 14890 5596
rect 14958 5584 15004 5596
rect 15054 5584 15100 5596
rect 15168 5584 15214 5596
rect 15264 5584 15310 5596
rect 15378 5584 15424 5596
rect 15474 5584 15520 5596
rect 15588 5584 15634 5596
rect 15684 5584 15730 5596
rect 15798 5584 15844 5596
rect 15894 5584 15940 5596
rect 16008 5584 16054 5596
rect 16104 5584 16150 5596
rect 16218 5584 16264 5596
rect 16314 5584 16360 5596
rect 16428 5584 16474 5596
rect 16524 5584 16570 5596
rect 16638 5584 16684 5596
rect 16734 5584 16780 5596
rect 16848 5584 16894 5596
rect 16944 5584 16990 5596
rect 17058 5584 17104 5596
rect 17154 5584 17200 5596
rect 17268 5584 17314 5596
rect 17364 5584 17410 5596
rect 17478 5584 17524 5596
rect 17574 5584 17620 5596
rect 17688 5584 17734 5596
rect 17784 5584 17830 5596
rect 17898 5584 17944 5596
rect 17994 5584 18040 5596
rect 18108 5584 18154 5596
rect 18204 5584 18250 5596
rect 18318 5584 18364 5596
rect 18414 5584 18460 5596
rect 18528 5584 18574 5596
rect 18624 5584 18670 5596
rect 9936 5537 18418 5544
rect 9936 5395 10392 5537
rect 10426 5395 10812 5537
rect 10846 5395 11232 5537
rect 11266 5395 11652 5537
rect 11686 5395 12072 5537
rect 12106 5395 12492 5537
rect 12526 5395 12912 5537
rect 12946 5395 13332 5537
rect 13366 5395 13752 5537
rect 13786 5395 14172 5537
rect 14206 5395 14592 5537
rect 14626 5395 15012 5537
rect 15046 5395 15432 5537
rect 15466 5395 15852 5537
rect 15886 5395 16272 5537
rect 16306 5395 16692 5537
rect 16726 5395 17112 5537
rect 17146 5395 17532 5537
rect 17566 5395 17952 5537
rect 17986 5395 18372 5537
rect 18406 5395 18418 5537
rect 9936 5388 18418 5395
rect 9936 5378 9946 5388
rect 5488 5336 5534 5348
rect 5584 5336 5630 5348
rect 5698 5336 5744 5348
rect 5794 5336 5840 5348
rect 5908 5336 5954 5348
rect 6004 5336 6050 5348
rect 6118 5336 6164 5348
rect 6214 5336 6260 5348
rect 6328 5336 6374 5348
rect 6424 5336 6470 5348
rect 6538 5336 6584 5348
rect 6634 5336 6680 5348
rect 6748 5336 6794 5348
rect 6844 5336 6890 5348
rect 6958 5336 7004 5348
rect 7054 5336 7100 5348
rect 7168 5336 7214 5348
rect 7264 5336 7310 5348
rect 7378 5336 7424 5348
rect 7474 5336 7520 5348
rect 7588 5336 7634 5348
rect 7684 5336 7730 5348
rect 7798 5336 7844 5348
rect 7894 5336 7940 5348
rect 8008 5336 8054 5348
rect 8104 5336 8150 5348
rect 8218 5336 8264 5348
rect 8314 5336 8360 5348
rect 8428 5336 8474 5348
rect 8524 5336 8570 5348
rect 8638 5336 8684 5348
rect 8734 5336 8780 5348
rect 8848 5336 8894 5348
rect 8944 5336 8990 5348
rect 9058 5336 9104 5348
rect 9154 5336 9200 5348
rect 5008 4520 5238 4736
rect 5008 4500 5018 4520
rect 3524 4340 3570 4352
rect 3620 4340 3666 4352
rect 3734 4340 3780 4352
rect 3830 4340 3876 4352
rect 3944 4340 3990 4352
rect 4040 4340 4086 4352
rect 4154 4340 4200 4352
rect 4250 4340 4296 4352
rect 3566 4302 3624 4308
rect 3566 4274 3578 4302
rect 2936 4256 3578 4274
rect 2784 4196 3578 4256
rect 2618 4152 2676 4159
rect 2576 4100 2622 4112
rect 2672 4100 2718 4112
rect 2768 4100 2814 4112
rect 2534 3124 2544 4100
rect 2616 3124 2626 4100
rect 2658 3124 2668 4100
rect 2722 3124 2732 4100
rect 2764 3124 2774 4100
rect 2846 3124 2856 4100
rect 2576 3112 2622 3124
rect 2672 3112 2718 3124
rect 2768 3112 2814 3124
rect 2996 3072 3110 4196
rect 3566 4159 3578 4196
rect 3612 4274 3624 4302
rect 3986 4302 4044 4308
rect 3986 4274 3998 4302
rect 3612 4196 3998 4274
rect 3612 4159 3624 4196
rect 3566 4153 3624 4159
rect 3986 4159 3998 4196
rect 4032 4262 4044 4302
rect 5052 4302 5238 4520
rect 5460 4360 5470 5336
rect 5528 4360 5538 5336
rect 5580 4360 5590 5336
rect 5738 4360 5748 5336
rect 5790 4360 5800 5336
rect 5948 4360 5958 5336
rect 6000 4360 6010 5336
rect 6158 4360 6168 5336
rect 6210 4360 6220 5336
rect 6368 4360 6378 5336
rect 6420 4360 6430 5336
rect 6578 4360 6588 5336
rect 6630 4360 6640 5336
rect 6788 4360 6798 5336
rect 6840 4360 6850 5336
rect 6998 4360 7008 5336
rect 7050 4360 7060 5336
rect 7208 4360 7218 5336
rect 7260 4360 7270 5336
rect 7418 4360 7428 5336
rect 7470 4360 7480 5336
rect 7628 4360 7638 5336
rect 7680 4360 7690 5336
rect 7838 4360 7848 5336
rect 7890 4360 7900 5336
rect 8048 4360 8058 5336
rect 8100 4360 8110 5336
rect 8258 4360 8268 5336
rect 8310 4360 8320 5336
rect 8468 4360 8478 5336
rect 8520 4360 8530 5336
rect 8678 4360 8688 5336
rect 8730 4360 8740 5336
rect 8888 4360 8898 5336
rect 8940 4360 8950 5336
rect 9098 4360 9108 5336
rect 9150 4360 9160 5336
rect 9218 4360 9228 5336
rect 5488 4348 5534 4360
rect 5584 4348 5630 4360
rect 5698 4348 5744 4360
rect 5794 4348 5840 4360
rect 5908 4348 5954 4360
rect 6004 4348 6050 4360
rect 6118 4348 6164 4360
rect 6214 4348 6260 4360
rect 6328 4348 6374 4360
rect 6424 4348 6470 4360
rect 6538 4348 6584 4360
rect 6634 4348 6680 4360
rect 6748 4348 6794 4360
rect 6844 4348 6890 4360
rect 6958 4348 7004 4360
rect 7054 4348 7100 4360
rect 7168 4348 7214 4360
rect 7264 4348 7310 4360
rect 7378 4348 7424 4360
rect 7474 4348 7520 4360
rect 7588 4348 7634 4360
rect 7684 4348 7730 4360
rect 7798 4348 7844 4360
rect 7894 4348 7940 4360
rect 8008 4348 8054 4360
rect 8104 4348 8150 4360
rect 8218 4348 8264 4360
rect 8314 4348 8360 4360
rect 8428 4348 8474 4360
rect 8524 4348 8570 4360
rect 8638 4348 8684 4360
rect 8734 4348 8780 4360
rect 8848 4348 8894 4360
rect 8944 4348 8990 4360
rect 9058 4348 9104 4360
rect 9154 4348 9200 4360
rect 9426 4308 9898 5378
rect 10338 5336 10384 5348
rect 10434 5336 10480 5348
rect 10548 5336 10594 5348
rect 10644 5336 10690 5348
rect 10758 5336 10804 5348
rect 10854 5336 10900 5348
rect 10968 5336 11014 5348
rect 11064 5336 11110 5348
rect 11178 5336 11224 5348
rect 11274 5336 11320 5348
rect 11388 5336 11434 5348
rect 11484 5336 11530 5348
rect 11598 5336 11644 5348
rect 11694 5336 11740 5348
rect 11808 5336 11854 5348
rect 11904 5336 11950 5348
rect 12018 5336 12064 5348
rect 12114 5336 12160 5348
rect 12228 5336 12274 5348
rect 12324 5336 12370 5348
rect 12438 5336 12484 5348
rect 12534 5336 12580 5348
rect 12648 5336 12694 5348
rect 12744 5336 12790 5348
rect 12858 5336 12904 5348
rect 12954 5336 13000 5348
rect 13068 5336 13114 5348
rect 13164 5336 13210 5348
rect 13278 5336 13324 5348
rect 13374 5336 13420 5348
rect 13488 5336 13534 5348
rect 13584 5336 13630 5348
rect 13698 5336 13744 5348
rect 13794 5336 13840 5348
rect 13908 5336 13954 5348
rect 14004 5336 14050 5348
rect 14118 5336 14164 5348
rect 14214 5336 14260 5348
rect 14328 5336 14374 5348
rect 14424 5336 14470 5348
rect 14538 5336 14584 5348
rect 14634 5336 14680 5348
rect 14748 5336 14794 5348
rect 14844 5336 14890 5348
rect 14958 5336 15004 5348
rect 15054 5336 15100 5348
rect 15168 5336 15214 5348
rect 15264 5336 15310 5348
rect 15378 5336 15424 5348
rect 15474 5336 15520 5348
rect 15588 5336 15634 5348
rect 15684 5336 15730 5348
rect 15798 5336 15844 5348
rect 15894 5336 15940 5348
rect 16008 5336 16054 5348
rect 16104 5336 16150 5348
rect 16218 5336 16264 5348
rect 16314 5336 16360 5348
rect 16428 5336 16474 5348
rect 16524 5336 16570 5348
rect 16638 5336 16684 5348
rect 16734 5336 16780 5348
rect 16848 5336 16894 5348
rect 16944 5336 16990 5348
rect 17058 5336 17104 5348
rect 17154 5336 17200 5348
rect 17268 5336 17314 5348
rect 17364 5336 17410 5348
rect 17478 5336 17524 5348
rect 17574 5336 17620 5348
rect 17688 5336 17734 5348
rect 17784 5336 17830 5348
rect 17898 5336 17944 5348
rect 17994 5336 18040 5348
rect 18108 5336 18154 5348
rect 18204 5336 18250 5348
rect 18318 5336 18364 5348
rect 18414 5336 18460 5348
rect 18528 5336 18574 5348
rect 18624 5336 18670 5348
rect 10310 4360 10320 5336
rect 10378 4360 10388 5336
rect 10430 4360 10440 5336
rect 10588 4360 10598 5336
rect 10640 4360 10650 5336
rect 10798 4360 10808 5336
rect 10850 4360 10860 5336
rect 11008 4360 11018 5336
rect 11060 4360 11070 5336
rect 11218 4360 11228 5336
rect 11270 4360 11280 5336
rect 11428 4360 11438 5336
rect 11480 4360 11490 5336
rect 11638 4360 11648 5336
rect 11690 4360 11700 5336
rect 11848 4360 11858 5336
rect 11900 4360 11910 5336
rect 12058 4360 12068 5336
rect 12110 4360 12120 5336
rect 12268 4360 12278 5336
rect 12320 4360 12330 5336
rect 12478 4360 12488 5336
rect 12530 4360 12540 5336
rect 12688 4360 12698 5336
rect 12740 4360 12750 5336
rect 12898 4360 12908 5336
rect 12950 4360 12960 5336
rect 13108 4360 13118 5336
rect 13160 4360 13170 5336
rect 13318 4360 13328 5336
rect 13370 4360 13380 5336
rect 13528 4360 13538 5336
rect 13580 4360 13590 5336
rect 13738 4360 13748 5336
rect 13790 4360 13800 5336
rect 13948 4360 13958 5336
rect 14000 4360 14010 5336
rect 14158 4360 14168 5336
rect 14210 4360 14220 5336
rect 14368 4360 14378 5336
rect 14420 4360 14430 5336
rect 14578 4360 14588 5336
rect 14630 4360 14640 5336
rect 14788 4360 14798 5336
rect 14840 4360 14850 5336
rect 14998 4360 15008 5336
rect 15050 4360 15060 5336
rect 15208 4360 15218 5336
rect 15260 4360 15270 5336
rect 15418 4360 15428 5336
rect 15470 4360 15480 5336
rect 15628 4360 15638 5336
rect 15680 4360 15690 5336
rect 15838 4360 15848 5336
rect 15890 4360 15900 5336
rect 16048 4360 16058 5336
rect 16100 4360 16110 5336
rect 16258 4360 16268 5336
rect 16310 4360 16320 5336
rect 16468 4360 16478 5336
rect 16520 4360 16530 5336
rect 16678 4360 16688 5336
rect 16730 4360 16740 5336
rect 16888 4360 16898 5336
rect 16940 4360 16950 5336
rect 17098 4360 17108 5336
rect 17150 4360 17160 5336
rect 17308 4360 17318 5336
rect 17360 4360 17370 5336
rect 17518 4360 17528 5336
rect 17570 4360 17580 5336
rect 17728 4360 17738 5336
rect 17780 4360 17790 5336
rect 17938 4360 17948 5336
rect 17990 4360 18000 5336
rect 18148 4360 18158 5336
rect 18200 4360 18210 5336
rect 18358 4360 18368 5336
rect 18410 4360 18420 5336
rect 18568 4360 18578 5336
rect 18620 4360 18630 5336
rect 18688 4360 18698 5336
rect 10338 4348 10384 4360
rect 10434 4348 10480 4360
rect 10548 4348 10594 4360
rect 10644 4348 10690 4360
rect 10758 4348 10804 4360
rect 10854 4348 10900 4360
rect 10968 4348 11014 4360
rect 11064 4348 11110 4360
rect 11178 4348 11224 4360
rect 11274 4348 11320 4360
rect 11388 4348 11434 4360
rect 11484 4348 11530 4360
rect 11598 4348 11644 4360
rect 11694 4348 11740 4360
rect 11808 4348 11854 4360
rect 11904 4348 11950 4360
rect 12018 4348 12064 4360
rect 12114 4348 12160 4360
rect 12228 4348 12274 4360
rect 12324 4348 12370 4360
rect 12438 4348 12484 4360
rect 12534 4348 12580 4360
rect 12648 4348 12694 4360
rect 12744 4348 12790 4360
rect 12858 4348 12904 4360
rect 12954 4348 13000 4360
rect 13068 4348 13114 4360
rect 13164 4348 13210 4360
rect 13278 4348 13324 4360
rect 13374 4348 13420 4360
rect 13488 4348 13534 4360
rect 13584 4348 13630 4360
rect 13698 4348 13744 4360
rect 13794 4348 13840 4360
rect 13908 4348 13954 4360
rect 14004 4348 14050 4360
rect 14118 4348 14164 4360
rect 14214 4348 14260 4360
rect 14328 4348 14374 4360
rect 14424 4348 14470 4360
rect 14538 4348 14584 4360
rect 14634 4348 14680 4360
rect 14748 4348 14794 4360
rect 14844 4348 14890 4360
rect 14958 4348 15004 4360
rect 15054 4348 15100 4360
rect 15168 4348 15214 4360
rect 15264 4348 15310 4360
rect 15378 4348 15424 4360
rect 15474 4348 15520 4360
rect 15588 4348 15634 4360
rect 15684 4348 15730 4360
rect 15798 4348 15844 4360
rect 15894 4348 15940 4360
rect 16008 4348 16054 4360
rect 16104 4348 16150 4360
rect 16218 4348 16264 4360
rect 16314 4348 16360 4360
rect 16428 4348 16474 4360
rect 16524 4348 16570 4360
rect 16638 4348 16684 4360
rect 16734 4348 16780 4360
rect 16848 4348 16894 4360
rect 16944 4348 16990 4360
rect 17058 4348 17104 4360
rect 17154 4348 17200 4360
rect 17268 4348 17314 4360
rect 17364 4348 17410 4360
rect 17478 4348 17524 4360
rect 17574 4348 17620 4360
rect 17688 4348 17734 4360
rect 17784 4348 17830 4360
rect 17898 4348 17944 4360
rect 17994 4348 18040 4360
rect 18108 4348 18154 4360
rect 18204 4348 18250 4360
rect 18318 4348 18364 4360
rect 18414 4348 18460 4360
rect 18528 4348 18574 4360
rect 18624 4348 18670 4360
rect 5740 4302 5798 4307
rect 6160 4302 6218 4307
rect 6580 4302 6638 4307
rect 7000 4302 7058 4307
rect 7420 4302 7478 4307
rect 7840 4302 7898 4307
rect 8260 4302 8318 4307
rect 8680 4302 8738 4307
rect 9100 4302 9158 4307
rect 5052 4301 9158 4302
rect 4032 4200 4038 4262
rect 4032 4193 4934 4200
rect 4032 4159 4418 4193
rect 4452 4192 4838 4193
rect 4872 4192 4934 4193
rect 3986 4158 4418 4159
rect 4502 4158 4838 4192
rect 4922 4158 4934 4192
rect 3986 4153 4934 4158
rect 4036 4150 4934 4153
rect 5052 4159 5752 4301
rect 5786 4159 6172 4301
rect 6206 4159 6592 4301
rect 6626 4159 7012 4301
rect 7046 4159 7432 4301
rect 7466 4159 7852 4301
rect 7886 4159 8272 4301
rect 8306 4159 8692 4301
rect 8726 4159 9112 4301
rect 9146 4159 9158 4301
rect 5052 4152 9158 4159
rect 9426 4301 18628 4308
rect 9426 4159 10602 4301
rect 10636 4159 11022 4301
rect 11056 4159 11442 4301
rect 11476 4159 11862 4301
rect 11896 4159 12282 4301
rect 12316 4159 12702 4301
rect 12736 4159 13122 4301
rect 13156 4159 13542 4301
rect 13576 4159 13962 4301
rect 13996 4159 14382 4301
rect 14416 4159 14802 4301
rect 14836 4159 15222 4301
rect 15256 4159 15642 4301
rect 15676 4159 16062 4301
rect 16096 4159 16482 4301
rect 16516 4159 16902 4301
rect 16936 4159 17322 4301
rect 17356 4159 17742 4301
rect 17776 4159 18162 4301
rect 18196 4159 18582 4301
rect 18616 4159 18628 4301
rect 9426 4152 18628 4159
rect 3314 4100 3360 4112
rect 3410 4100 3456 4112
rect 3524 4100 3570 4112
rect 3620 4100 3666 4112
rect 3734 4100 3780 4112
rect 3830 4100 3876 4112
rect 3944 4100 3990 4112
rect 4040 4100 4086 4112
rect 4154 4100 4200 4112
rect 4250 4100 4296 4112
rect 4364 4100 4410 4112
rect 4460 4100 4506 4112
rect 4574 4100 4620 4112
rect 4670 4100 4716 4112
rect 4784 4100 4830 4112
rect 4880 4100 4926 4112
rect 3286 3124 3296 4100
rect 3354 3124 3364 4100
rect 3406 3124 3416 4100
rect 3564 3124 3574 4100
rect 3616 3124 3626 4100
rect 3774 3124 3784 4100
rect 3826 3124 3836 4100
rect 3984 3124 3994 4100
rect 4036 3124 4046 4100
rect 4194 3124 4204 4100
rect 4246 3124 4256 4100
rect 4404 3124 4414 4100
rect 4456 3124 4466 4100
rect 4614 3124 4624 4100
rect 4666 3124 4676 4100
rect 4824 3124 4834 4100
rect 4876 3124 4886 4100
rect 4944 3124 4954 4100
rect 3314 3112 3360 3124
rect 3410 3112 3456 3124
rect 3524 3112 3570 3124
rect 3620 3112 3666 3124
rect 3734 3112 3780 3124
rect 3830 3112 3876 3124
rect 3944 3112 3990 3124
rect 4040 3112 4086 3124
rect 4154 3112 4200 3124
rect 4250 3112 4296 3124
rect 4364 3112 4410 3124
rect 4460 3112 4506 3124
rect 4574 3112 4620 3124
rect 4670 3112 4716 3124
rect 4784 3112 4830 3124
rect 4880 3112 4926 3124
rect 5052 3072 5238 4152
rect 5488 4100 5534 4112
rect 5584 4100 5630 4112
rect 5698 4100 5744 4112
rect 5794 4100 5840 4112
rect 5908 4100 5954 4112
rect 6004 4100 6050 4112
rect 6118 4100 6164 4112
rect 6214 4100 6260 4112
rect 6328 4100 6374 4112
rect 6424 4100 6470 4112
rect 6538 4100 6584 4112
rect 6634 4100 6680 4112
rect 6748 4100 6794 4112
rect 6844 4100 6890 4112
rect 6958 4100 7004 4112
rect 7054 4100 7100 4112
rect 7168 4100 7214 4112
rect 7264 4100 7310 4112
rect 7378 4100 7424 4112
rect 7474 4100 7520 4112
rect 7588 4100 7634 4112
rect 7684 4100 7730 4112
rect 7798 4100 7844 4112
rect 7894 4100 7940 4112
rect 8008 4100 8054 4112
rect 8104 4100 8150 4112
rect 8218 4100 8264 4112
rect 8314 4100 8360 4112
rect 8428 4100 8474 4112
rect 8524 4100 8570 4112
rect 8638 4100 8684 4112
rect 8734 4100 8780 4112
rect 8848 4100 8894 4112
rect 8944 4100 8990 4112
rect 9058 4100 9104 4112
rect 9154 4100 9200 4112
rect 5460 3124 5470 4100
rect 5528 3124 5538 4100
rect 5580 3124 5590 4100
rect 5738 3124 5748 4100
rect 5790 3124 5800 4100
rect 5948 3124 5958 4100
rect 6000 3124 6010 4100
rect 6158 3124 6168 4100
rect 6210 3124 6220 4100
rect 6368 3124 6378 4100
rect 6420 3124 6430 4100
rect 6578 3124 6588 4100
rect 6630 3124 6640 4100
rect 6788 3124 6798 4100
rect 6840 3124 6850 4100
rect 6998 3124 7008 4100
rect 7050 3124 7060 4100
rect 7208 3124 7218 4100
rect 7260 3124 7270 4100
rect 7418 3124 7428 4100
rect 7470 3124 7480 4100
rect 7628 3124 7638 4100
rect 7680 3124 7690 4100
rect 7838 3124 7848 4100
rect 7890 3124 7900 4100
rect 8048 3124 8058 4100
rect 8100 3124 8110 4100
rect 8258 3124 8268 4100
rect 8310 3124 8320 4100
rect 8468 3124 8478 4100
rect 8520 3124 8530 4100
rect 8678 3124 8688 4100
rect 8730 3124 8740 4100
rect 8888 3124 8898 4100
rect 8940 3124 8950 4100
rect 9098 3124 9108 4100
rect 9150 3124 9160 4100
rect 9218 3124 9228 4100
rect 5488 3112 5534 3124
rect 5584 3112 5630 3124
rect 5698 3112 5744 3124
rect 5794 3112 5840 3124
rect 5908 3112 5954 3124
rect 6004 3112 6050 3124
rect 6118 3112 6164 3124
rect 6214 3112 6260 3124
rect 6328 3112 6374 3124
rect 6424 3112 6470 3124
rect 6538 3112 6584 3124
rect 6634 3112 6680 3124
rect 6748 3112 6794 3124
rect 6844 3112 6890 3124
rect 6958 3112 7004 3124
rect 7054 3112 7100 3124
rect 7168 3112 7214 3124
rect 7264 3112 7310 3124
rect 7378 3112 7424 3124
rect 7474 3112 7520 3124
rect 7588 3112 7634 3124
rect 7684 3112 7730 3124
rect 7798 3112 7844 3124
rect 7894 3112 7940 3124
rect 8008 3112 8054 3124
rect 8104 3112 8150 3124
rect 8218 3112 8264 3124
rect 8314 3112 8360 3124
rect 8428 3112 8474 3124
rect 8524 3112 8570 3124
rect 8638 3112 8684 3124
rect 8734 3112 8780 3124
rect 8848 3112 8894 3124
rect 8944 3112 8990 3124
rect 9058 3112 9104 3124
rect 9154 3112 9200 3124
rect 9426 3072 9898 4152
rect 10338 4100 10384 4112
rect 10434 4100 10480 4112
rect 10548 4100 10594 4112
rect 10644 4100 10690 4112
rect 10758 4100 10804 4112
rect 10854 4100 10900 4112
rect 10968 4100 11014 4112
rect 11064 4100 11110 4112
rect 11178 4100 11224 4112
rect 11274 4100 11320 4112
rect 11388 4100 11434 4112
rect 11484 4100 11530 4112
rect 11598 4100 11644 4112
rect 11694 4100 11740 4112
rect 11808 4100 11854 4112
rect 11904 4100 11950 4112
rect 12018 4100 12064 4112
rect 12114 4100 12160 4112
rect 12228 4100 12274 4112
rect 12324 4100 12370 4112
rect 12438 4100 12484 4112
rect 12534 4100 12580 4112
rect 12648 4100 12694 4112
rect 12744 4100 12790 4112
rect 12858 4100 12904 4112
rect 12954 4100 13000 4112
rect 13068 4100 13114 4112
rect 13164 4100 13210 4112
rect 13278 4100 13324 4112
rect 13374 4100 13420 4112
rect 13488 4100 13534 4112
rect 13584 4100 13630 4112
rect 13698 4100 13744 4112
rect 13794 4100 13840 4112
rect 13908 4100 13954 4112
rect 14004 4100 14050 4112
rect 14118 4100 14164 4112
rect 14214 4100 14260 4112
rect 14328 4100 14374 4112
rect 14424 4100 14470 4112
rect 14538 4100 14584 4112
rect 14634 4100 14680 4112
rect 14748 4100 14794 4112
rect 14844 4100 14890 4112
rect 14958 4100 15004 4112
rect 15054 4100 15100 4112
rect 15168 4100 15214 4112
rect 15264 4100 15310 4112
rect 15378 4100 15424 4112
rect 15474 4100 15520 4112
rect 15588 4100 15634 4112
rect 15684 4100 15730 4112
rect 15798 4100 15844 4112
rect 15894 4100 15940 4112
rect 16008 4100 16054 4112
rect 16104 4100 16150 4112
rect 16218 4100 16264 4112
rect 16314 4100 16360 4112
rect 16428 4100 16474 4112
rect 16524 4100 16570 4112
rect 16638 4100 16684 4112
rect 16734 4100 16780 4112
rect 16848 4100 16894 4112
rect 16944 4100 16990 4112
rect 17058 4100 17104 4112
rect 17154 4100 17200 4112
rect 17268 4100 17314 4112
rect 17364 4100 17410 4112
rect 17478 4100 17524 4112
rect 17574 4100 17620 4112
rect 17688 4100 17734 4112
rect 17784 4100 17830 4112
rect 17898 4100 17944 4112
rect 17994 4100 18040 4112
rect 18108 4100 18154 4112
rect 18204 4100 18250 4112
rect 18318 4100 18364 4112
rect 18414 4100 18460 4112
rect 18528 4100 18574 4112
rect 18624 4100 18670 4112
rect 10310 3124 10320 4100
rect 10378 3124 10388 4100
rect 10430 3124 10440 4100
rect 10588 3124 10598 4100
rect 10640 3124 10650 4100
rect 10798 3124 10808 4100
rect 10850 3124 10860 4100
rect 11008 3124 11018 4100
rect 11060 3124 11070 4100
rect 11218 3124 11228 4100
rect 11270 3124 11280 4100
rect 11428 3124 11438 4100
rect 11480 3124 11490 4100
rect 11638 3124 11648 4100
rect 11690 3124 11700 4100
rect 11848 3124 11858 4100
rect 11900 3124 11910 4100
rect 12058 3124 12068 4100
rect 12110 3124 12120 4100
rect 12268 3124 12278 4100
rect 12320 3124 12330 4100
rect 12478 3124 12488 4100
rect 12530 3124 12540 4100
rect 12688 3124 12698 4100
rect 12740 3124 12750 4100
rect 12898 3124 12908 4100
rect 12950 3124 12960 4100
rect 13108 3124 13118 4100
rect 13160 3124 13170 4100
rect 13318 3124 13328 4100
rect 13370 3124 13380 4100
rect 13528 3124 13538 4100
rect 13580 3124 13590 4100
rect 13738 3124 13748 4100
rect 13790 3124 13800 4100
rect 13948 3124 13958 4100
rect 14000 3124 14010 4100
rect 14158 3124 14168 4100
rect 14210 3124 14220 4100
rect 14368 3124 14378 4100
rect 14420 3124 14430 4100
rect 14578 3124 14588 4100
rect 14630 3124 14640 4100
rect 14788 3124 14798 4100
rect 14840 3124 14850 4100
rect 14998 3124 15008 4100
rect 15050 3124 15060 4100
rect 15208 3124 15218 4100
rect 15260 3124 15270 4100
rect 15418 3124 15428 4100
rect 15470 3124 15480 4100
rect 15628 3124 15638 4100
rect 15680 3124 15690 4100
rect 15838 3124 15848 4100
rect 15890 3124 15900 4100
rect 16048 3124 16058 4100
rect 16100 3124 16110 4100
rect 16258 3124 16268 4100
rect 16310 3124 16320 4100
rect 16468 3124 16478 4100
rect 16520 3124 16530 4100
rect 16678 3124 16688 4100
rect 16730 3124 16740 4100
rect 16888 3124 16898 4100
rect 16940 3124 16950 4100
rect 17098 3124 17108 4100
rect 17150 3124 17160 4100
rect 17308 3124 17318 4100
rect 17360 3124 17370 4100
rect 17518 3124 17528 4100
rect 17570 3124 17580 4100
rect 17728 3124 17738 4100
rect 17780 3124 17790 4100
rect 17938 3124 17948 4100
rect 17990 3124 18000 4100
rect 18148 3124 18158 4100
rect 18200 3124 18210 4100
rect 18358 3124 18368 4100
rect 18410 3124 18420 4100
rect 18568 3124 18578 4100
rect 18620 3124 18630 4100
rect 18688 3124 18698 4100
rect 10338 3112 10384 3124
rect 10434 3112 10480 3124
rect 10548 3112 10594 3124
rect 10644 3112 10690 3124
rect 10758 3112 10804 3124
rect 10854 3112 10900 3124
rect 10968 3112 11014 3124
rect 11064 3112 11110 3124
rect 11178 3112 11224 3124
rect 11274 3112 11320 3124
rect 11388 3112 11434 3124
rect 11484 3112 11530 3124
rect 11598 3112 11644 3124
rect 11694 3112 11740 3124
rect 11808 3112 11854 3124
rect 11904 3112 11950 3124
rect 12018 3112 12064 3124
rect 12114 3112 12160 3124
rect 12228 3112 12274 3124
rect 12324 3112 12370 3124
rect 12438 3112 12484 3124
rect 12534 3112 12580 3124
rect 12648 3112 12694 3124
rect 12744 3112 12790 3124
rect 12858 3112 12904 3124
rect 12954 3112 13000 3124
rect 13068 3112 13114 3124
rect 13164 3112 13210 3124
rect 13278 3112 13324 3124
rect 13374 3112 13420 3124
rect 13488 3112 13534 3124
rect 13584 3112 13630 3124
rect 13698 3112 13744 3124
rect 13794 3112 13840 3124
rect 13908 3112 13954 3124
rect 14004 3112 14050 3124
rect 14118 3112 14164 3124
rect 14214 3112 14260 3124
rect 14328 3112 14374 3124
rect 14424 3112 14470 3124
rect 14538 3112 14584 3124
rect 14634 3112 14680 3124
rect 14748 3112 14794 3124
rect 14844 3112 14890 3124
rect 14958 3112 15004 3124
rect 15054 3112 15100 3124
rect 15168 3112 15214 3124
rect 15264 3112 15310 3124
rect 15378 3112 15424 3124
rect 15474 3112 15520 3124
rect 15588 3112 15634 3124
rect 15684 3112 15730 3124
rect 15798 3112 15844 3124
rect 15894 3112 15940 3124
rect 16008 3112 16054 3124
rect 16104 3112 16150 3124
rect 16218 3112 16264 3124
rect 16314 3112 16360 3124
rect 16428 3112 16474 3124
rect 16524 3112 16570 3124
rect 16638 3112 16684 3124
rect 16734 3112 16780 3124
rect 16848 3112 16894 3124
rect 16944 3112 16990 3124
rect 17058 3112 17104 3124
rect 17154 3112 17200 3124
rect 17268 3112 17314 3124
rect 17364 3112 17410 3124
rect 17478 3112 17524 3124
rect 17574 3112 17620 3124
rect 17688 3112 17734 3124
rect 17784 3112 17830 3124
rect 17898 3112 17944 3124
rect 17994 3112 18040 3124
rect 18108 3112 18154 3124
rect 18204 3112 18250 3124
rect 18318 3112 18364 3124
rect 18414 3112 18460 3124
rect 18528 3112 18574 3124
rect 18624 3112 18670 3124
rect 2228 3066 2822 3072
rect 2228 3032 2726 3066
rect 2810 3032 2822 3066
rect 2228 3026 2822 3032
rect 2996 3070 3150 3072
rect 3356 3070 3414 3071
rect 3776 3070 3834 3071
rect 4196 3070 4254 3071
rect 4616 3070 4674 3071
rect 2996 3065 4724 3070
rect 2996 3030 3368 3065
rect 3402 3064 3788 3065
rect 3822 3064 4208 3065
rect 4242 3064 4628 3065
rect 4662 3064 4724 3065
rect 3452 3030 3788 3064
rect 3872 3030 4208 3064
rect 4292 3030 4628 3064
rect 4712 3030 4724 3064
rect 2228 3024 2768 3026
rect 2996 3024 4724 3030
rect 5052 3065 8998 3072
rect 5052 3030 5542 3065
rect 5576 3064 5962 3065
rect 5996 3064 6382 3065
rect 6416 3064 6802 3065
rect 6836 3064 7222 3065
rect 7256 3064 7642 3065
rect 7676 3064 8062 3065
rect 8096 3064 8482 3065
rect 8516 3064 8902 3065
rect 8936 3064 8998 3065
rect 5626 3030 5962 3064
rect 6046 3030 6382 3064
rect 6466 3030 6802 3064
rect 6886 3030 7222 3064
rect 7306 3030 7642 3064
rect 7726 3030 8062 3064
rect 8146 3030 8482 3064
rect 8566 3030 8902 3064
rect 8986 3030 8998 3064
rect 186 2220 196 2482
rect 524 2220 534 2482
rect 304 2122 416 2220
rect 2228 2122 2322 3024
rect 3352 3022 3410 3024
rect 3772 3022 3830 3024
rect 4192 3022 4250 3024
rect 4612 3022 4670 3024
rect 5052 3022 8998 3030
rect 9426 3065 18468 3072
rect 9426 3030 10392 3065
rect 10426 3064 10812 3065
rect 10846 3064 11232 3065
rect 11266 3064 11652 3065
rect 11686 3064 12072 3065
rect 12106 3064 12492 3065
rect 12526 3064 12912 3065
rect 12946 3064 13332 3065
rect 13366 3064 13752 3065
rect 13786 3064 14172 3065
rect 14206 3064 14592 3065
rect 14626 3064 15012 3065
rect 15046 3064 15432 3065
rect 15466 3064 15852 3065
rect 15886 3064 16272 3065
rect 16306 3064 16692 3065
rect 16726 3064 17112 3065
rect 17146 3064 17532 3065
rect 17566 3064 17952 3065
rect 17986 3064 18372 3065
rect 18406 3064 18468 3065
rect 10476 3030 10812 3064
rect 10896 3030 11232 3064
rect 11316 3030 11652 3064
rect 11736 3030 12072 3064
rect 12156 3030 12492 3064
rect 12576 3030 12912 3064
rect 12996 3030 13332 3064
rect 13416 3030 13752 3064
rect 13836 3030 14172 3064
rect 14256 3030 14592 3064
rect 14676 3030 15012 3064
rect 15096 3030 15432 3064
rect 15516 3030 15852 3064
rect 15936 3030 16272 3064
rect 16356 3030 16692 3064
rect 16776 3030 17112 3064
rect 17196 3030 17532 3064
rect 17616 3030 17952 3064
rect 18036 3030 18372 3064
rect 18456 3030 18468 3064
rect 9426 3022 18468 3030
rect 2978 2838 3134 2850
rect 2974 2690 2984 2838
rect 3128 2690 3138 2838
rect 2978 2678 3134 2690
rect 304 2044 2322 2122
rect -958 1486 -16 1544
rect -958 48 -886 1486
rect -198 1400 -188 1458
rect -114 1400 -104 1458
rect 304 1446 416 2044
rect 90 1406 416 1446
rect 4376 1286 4386 1534
rect 4630 1286 4640 1534
rect -528 68 -192 126
rect -958 2 -712 48
rect -36 -14 -26 40
rect 36 -14 46 40
rect 124 10 416 50
rect 304 -518 416 10
rect 4416 -468 4600 1286
rect 5054 222 5238 3022
rect 5354 2970 5478 2976
rect 5354 2870 5366 2970
rect 5466 2870 5478 2970
rect 5354 2864 5478 2870
rect 5774 2970 5898 2976
rect 5774 2870 5786 2970
rect 5886 2870 5898 2970
rect 5774 2864 5898 2870
rect 6194 2970 6318 2976
rect 6194 2870 6206 2970
rect 6306 2870 6318 2970
rect 6194 2864 6318 2870
rect 6614 2970 6738 2976
rect 6614 2870 6626 2970
rect 6726 2870 6738 2970
rect 6614 2864 6738 2870
rect 7034 2970 7158 2976
rect 7034 2870 7046 2970
rect 7146 2870 7158 2970
rect 7034 2864 7158 2870
rect 7454 2970 7578 2976
rect 7454 2870 7466 2970
rect 7566 2870 7578 2970
rect 7454 2864 7578 2870
rect 7874 2970 7998 2976
rect 7874 2870 7886 2970
rect 7986 2870 7998 2970
rect 7874 2864 7998 2870
rect 8294 2970 8418 2976
rect 8294 2870 8306 2970
rect 8406 2870 8418 2970
rect 8294 2864 8418 2870
rect 8714 2970 8838 2976
rect 8714 2870 8726 2970
rect 8826 2870 8838 2970
rect 8714 2864 8838 2870
rect 9134 2970 9258 2976
rect 9134 2870 9146 2970
rect 9246 2870 9258 2970
rect 9134 2864 9258 2870
rect 10196 2954 10320 2960
rect 10196 2854 10208 2954
rect 10308 2854 10320 2954
rect 10196 2848 10320 2854
rect 10616 2954 10740 2960
rect 10616 2854 10628 2954
rect 10728 2854 10740 2954
rect 10616 2848 10740 2854
rect 11036 2954 11160 2960
rect 11036 2854 11048 2954
rect 11148 2854 11160 2954
rect 11036 2848 11160 2854
rect 11456 2954 11580 2960
rect 11456 2854 11468 2954
rect 11568 2854 11580 2954
rect 11456 2848 11580 2854
rect 11876 2954 12000 2960
rect 11876 2854 11888 2954
rect 11988 2854 12000 2954
rect 11876 2848 12000 2854
rect 12296 2954 12420 2960
rect 12296 2854 12308 2954
rect 12408 2854 12420 2954
rect 12296 2848 12420 2854
rect 12716 2954 12840 2960
rect 12716 2854 12728 2954
rect 12828 2854 12840 2954
rect 12716 2848 12840 2854
rect 13136 2954 13260 2960
rect 13136 2854 13148 2954
rect 13248 2854 13260 2954
rect 13136 2848 13260 2854
rect 13556 2954 13680 2960
rect 13556 2854 13568 2954
rect 13668 2854 13680 2954
rect 13556 2848 13680 2854
rect 13976 2954 14100 2960
rect 13976 2854 13988 2954
rect 14088 2854 14100 2954
rect 13976 2848 14100 2854
rect 14396 2954 14520 2960
rect 14396 2854 14408 2954
rect 14508 2854 14520 2954
rect 14396 2848 14520 2854
rect 14816 2954 14940 2960
rect 14816 2854 14828 2954
rect 14928 2854 14940 2954
rect 14816 2848 14940 2854
rect 15236 2954 15360 2960
rect 15236 2854 15248 2954
rect 15348 2854 15360 2954
rect 15236 2848 15360 2854
rect 15656 2954 15780 2960
rect 15656 2854 15668 2954
rect 15768 2854 15780 2954
rect 15656 2848 15780 2854
rect 16076 2954 16200 2960
rect 16076 2854 16088 2954
rect 16188 2854 16200 2954
rect 16076 2848 16200 2854
rect 16496 2954 16620 2960
rect 16496 2854 16508 2954
rect 16608 2854 16620 2954
rect 16496 2848 16620 2854
rect 16916 2954 17040 2960
rect 16916 2854 16928 2954
rect 17028 2854 17040 2954
rect 16916 2848 17040 2854
rect 17336 2954 17460 2960
rect 17336 2854 17348 2954
rect 17448 2854 17460 2954
rect 17336 2848 17460 2854
rect 17756 2954 17880 2960
rect 17756 2854 17768 2954
rect 17868 2854 17880 2954
rect 17756 2848 17880 2854
rect 18176 2954 18300 2960
rect 18176 2854 18188 2954
rect 18288 2854 18300 2954
rect 18176 2848 18300 2854
rect 18596 2954 18720 2960
rect 18596 2854 18608 2954
rect 18708 2854 18720 2954
rect 18596 2848 18720 2854
rect 5010 -26 5020 222
rect 5264 -26 5274 222
rect 304 -596 2322 -518
rect 304 -694 416 -596
rect 186 -956 196 -694
rect 524 -956 534 -694
rect 2228 -1498 2322 -596
rect 4416 -636 5238 -468
rect 2978 -1164 3134 -1152
rect 2974 -1312 2984 -1164
rect 3128 -1312 3138 -1164
rect 2978 -1324 3134 -1312
rect 5052 -1496 5238 -636
rect 5354 -1344 5478 -1338
rect 5354 -1444 5366 -1344
rect 5466 -1444 5478 -1344
rect 5354 -1450 5478 -1444
rect 5774 -1344 5898 -1338
rect 5774 -1444 5786 -1344
rect 5886 -1444 5898 -1344
rect 5774 -1450 5898 -1444
rect 6194 -1344 6318 -1338
rect 6194 -1444 6206 -1344
rect 6306 -1444 6318 -1344
rect 6194 -1450 6318 -1444
rect 6614 -1344 6738 -1338
rect 6614 -1444 6626 -1344
rect 6726 -1444 6738 -1344
rect 6614 -1450 6738 -1444
rect 7034 -1344 7158 -1338
rect 7034 -1444 7046 -1344
rect 7146 -1444 7158 -1344
rect 7034 -1450 7158 -1444
rect 7454 -1344 7578 -1338
rect 7454 -1444 7466 -1344
rect 7566 -1444 7578 -1344
rect 7454 -1450 7578 -1444
rect 7874 -1344 7998 -1338
rect 7874 -1444 7886 -1344
rect 7986 -1444 7998 -1344
rect 7874 -1450 7998 -1444
rect 8294 -1344 8418 -1338
rect 8294 -1444 8306 -1344
rect 8406 -1444 8418 -1344
rect 8294 -1450 8418 -1444
rect 8714 -1344 8838 -1338
rect 8714 -1444 8726 -1344
rect 8826 -1444 8838 -1344
rect 8714 -1450 8838 -1444
rect 9134 -1344 9258 -1338
rect 9134 -1444 9146 -1344
rect 9246 -1444 9258 -1344
rect 9134 -1450 9258 -1444
rect 3352 -1498 3410 -1496
rect 3772 -1498 3830 -1496
rect 4192 -1498 4250 -1496
rect 4612 -1498 4670 -1496
rect 2228 -1500 2768 -1498
rect 2228 -1506 2822 -1500
rect 2228 -1540 2726 -1506
rect 2810 -1540 2822 -1506
rect 2228 -1546 2822 -1540
rect 2996 -1504 4724 -1498
rect 2996 -1539 3368 -1504
rect 3452 -1538 3788 -1504
rect 3872 -1538 4208 -1504
rect 4292 -1538 4628 -1504
rect 4712 -1538 4724 -1504
rect 3402 -1539 3788 -1538
rect 3822 -1539 4208 -1538
rect 4242 -1539 4628 -1538
rect 4662 -1539 4724 -1538
rect 2996 -1544 4724 -1539
rect 5052 -1504 8998 -1496
rect 5052 -1539 5542 -1504
rect 5626 -1538 5962 -1504
rect 6046 -1538 6382 -1504
rect 6466 -1538 6802 -1504
rect 6886 -1538 7222 -1504
rect 7306 -1538 7642 -1504
rect 7726 -1538 8062 -1504
rect 8146 -1538 8482 -1504
rect 8566 -1538 8902 -1504
rect 8986 -1538 8998 -1504
rect 5576 -1539 5962 -1538
rect 5996 -1539 6382 -1538
rect 6416 -1539 6802 -1538
rect 6836 -1539 7222 -1538
rect 7256 -1539 7642 -1538
rect 7676 -1539 8062 -1538
rect 8096 -1539 8482 -1538
rect 8516 -1539 8902 -1538
rect 8936 -1539 8998 -1538
rect 2996 -1546 3150 -1544
rect 3356 -1545 3414 -1544
rect 3776 -1545 3834 -1544
rect 4196 -1545 4254 -1544
rect 4616 -1545 4674 -1544
rect 5052 -1546 8998 -1539
rect 2228 -2676 2322 -1546
rect 2576 -1598 2622 -1586
rect 2672 -1598 2718 -1586
rect 2768 -1598 2814 -1586
rect 2534 -2574 2544 -1598
rect 2616 -2574 2626 -1598
rect 2658 -2574 2668 -1598
rect 2722 -2574 2732 -1598
rect 2764 -2574 2774 -1598
rect 2846 -2574 2856 -1598
rect 2576 -2586 2622 -2574
rect 2672 -2586 2718 -2574
rect 2768 -2586 2814 -2574
rect 2618 -2633 2676 -2626
rect 2618 -2676 2630 -2633
rect 2228 -2724 2630 -2676
rect 2618 -2776 2630 -2724
rect 2664 -2776 2676 -2633
rect 2996 -2670 3110 -1546
rect 3314 -1598 3360 -1586
rect 3410 -1598 3456 -1586
rect 3524 -1598 3570 -1586
rect 3620 -1598 3666 -1586
rect 3734 -1598 3780 -1586
rect 3830 -1598 3876 -1586
rect 3944 -1598 3990 -1586
rect 4040 -1598 4086 -1586
rect 4154 -1598 4200 -1586
rect 4250 -1598 4296 -1586
rect 4364 -1598 4410 -1586
rect 4460 -1598 4506 -1586
rect 4574 -1598 4620 -1586
rect 4670 -1598 4716 -1586
rect 4784 -1598 4830 -1586
rect 4880 -1598 4926 -1586
rect 3286 -2574 3296 -1598
rect 3354 -2574 3364 -1598
rect 3406 -2574 3416 -1598
rect 3564 -2574 3574 -1598
rect 3616 -2574 3626 -1598
rect 3774 -2574 3784 -1598
rect 3826 -2574 3836 -1598
rect 3984 -2574 3994 -1598
rect 4036 -2574 4046 -1598
rect 4194 -2574 4204 -1598
rect 4246 -2574 4256 -1598
rect 4404 -2574 4414 -1598
rect 4456 -2574 4466 -1598
rect 4614 -2574 4624 -1598
rect 4666 -2574 4676 -1598
rect 4824 -2574 4834 -1598
rect 4876 -2574 4886 -1598
rect 4944 -2574 4954 -1598
rect 3314 -2586 3360 -2574
rect 3410 -2586 3456 -2574
rect 3524 -2586 3570 -2574
rect 3620 -2586 3666 -2574
rect 3734 -2586 3780 -2574
rect 3830 -2586 3876 -2574
rect 3944 -2586 3990 -2574
rect 4040 -2586 4086 -2574
rect 4154 -2586 4200 -2574
rect 4250 -2586 4296 -2574
rect 4364 -2586 4410 -2574
rect 4460 -2586 4506 -2574
rect 4574 -2586 4620 -2574
rect 4670 -2586 4716 -2574
rect 4784 -2586 4830 -2574
rect 4880 -2586 4926 -2574
rect 4036 -2627 4934 -2624
rect 3566 -2633 3624 -2627
rect 3566 -2670 3578 -2633
rect 2618 -2782 2676 -2776
rect 2784 -2730 3578 -2670
rect 2580 -2826 2626 -2814
rect 2668 -2826 2714 -2814
rect 2556 -3802 2566 -2826
rect 2620 -3802 2630 -2826
rect 2664 -3802 2674 -2826
rect 2728 -3802 2738 -2826
rect 2784 -2878 2794 -2730
rect 2936 -2748 3578 -2730
rect 2936 -2878 2946 -2748
rect 3566 -2776 3578 -2748
rect 3612 -2670 3624 -2633
rect 3986 -2632 4934 -2627
rect 3986 -2633 4418 -2632
rect 3986 -2670 3998 -2633
rect 3612 -2748 3998 -2670
rect 3612 -2776 3624 -2748
rect 3566 -2782 3624 -2776
rect 3986 -2776 3998 -2748
rect 4032 -2667 4418 -2633
rect 4502 -2666 4838 -2632
rect 4922 -2666 4934 -2632
rect 4452 -2667 4838 -2666
rect 4872 -2667 4934 -2666
rect 4032 -2674 4934 -2667
rect 5052 -2626 5238 -1546
rect 5488 -1598 5534 -1586
rect 5584 -1598 5630 -1586
rect 5698 -1598 5744 -1586
rect 5794 -1598 5840 -1586
rect 5908 -1598 5954 -1586
rect 6004 -1598 6050 -1586
rect 6118 -1598 6164 -1586
rect 6214 -1598 6260 -1586
rect 6328 -1598 6374 -1586
rect 6424 -1598 6470 -1586
rect 6538 -1598 6584 -1586
rect 6634 -1598 6680 -1586
rect 6748 -1598 6794 -1586
rect 6844 -1598 6890 -1586
rect 6958 -1598 7004 -1586
rect 7054 -1598 7100 -1586
rect 7168 -1598 7214 -1586
rect 7264 -1598 7310 -1586
rect 7378 -1598 7424 -1586
rect 7474 -1598 7520 -1586
rect 7588 -1598 7634 -1586
rect 7684 -1598 7730 -1586
rect 7798 -1598 7844 -1586
rect 7894 -1598 7940 -1586
rect 8008 -1598 8054 -1586
rect 8104 -1598 8150 -1586
rect 8218 -1598 8264 -1586
rect 8314 -1598 8360 -1586
rect 8428 -1598 8474 -1586
rect 8524 -1598 8570 -1586
rect 8638 -1598 8684 -1586
rect 8734 -1598 8780 -1586
rect 8848 -1598 8894 -1586
rect 8944 -1598 8990 -1586
rect 9058 -1598 9104 -1586
rect 9154 -1598 9200 -1586
rect 5460 -2574 5470 -1598
rect 5528 -2574 5538 -1598
rect 5580 -2574 5590 -1598
rect 5738 -2574 5748 -1598
rect 5790 -2574 5800 -1598
rect 5948 -2574 5958 -1598
rect 6000 -2574 6010 -1598
rect 6158 -2574 6168 -1598
rect 6210 -2574 6220 -1598
rect 6368 -2574 6378 -1598
rect 6420 -2574 6430 -1598
rect 6578 -2574 6588 -1598
rect 6630 -2574 6640 -1598
rect 6788 -2574 6798 -1598
rect 6840 -2574 6850 -1598
rect 6998 -2574 7008 -1598
rect 7050 -2574 7060 -1598
rect 7208 -2574 7218 -1598
rect 7260 -2574 7270 -1598
rect 7418 -2574 7428 -1598
rect 7470 -2574 7480 -1598
rect 7628 -2574 7638 -1598
rect 7680 -2574 7690 -1598
rect 7838 -2574 7848 -1598
rect 7890 -2574 7900 -1598
rect 8048 -2574 8058 -1598
rect 8100 -2574 8110 -1598
rect 8258 -2574 8268 -1598
rect 8310 -2574 8320 -1598
rect 8468 -2574 8478 -1598
rect 8520 -2574 8530 -1598
rect 8678 -2574 8688 -1598
rect 8730 -2574 8740 -1598
rect 8888 -2574 8898 -1598
rect 8940 -2574 8950 -1598
rect 9098 -2574 9108 -1598
rect 9150 -2574 9160 -1598
rect 9218 -2574 9228 -1598
rect 5488 -2586 5534 -2574
rect 5584 -2586 5630 -2574
rect 5698 -2586 5744 -2574
rect 5794 -2586 5840 -2574
rect 5908 -2586 5954 -2574
rect 6004 -2586 6050 -2574
rect 6118 -2586 6164 -2574
rect 6214 -2586 6260 -2574
rect 6328 -2586 6374 -2574
rect 6424 -2586 6470 -2574
rect 6538 -2586 6584 -2574
rect 6634 -2586 6680 -2574
rect 6748 -2586 6794 -2574
rect 6844 -2586 6890 -2574
rect 6958 -2586 7004 -2574
rect 7054 -2586 7100 -2574
rect 7168 -2586 7214 -2574
rect 7264 -2586 7310 -2574
rect 7378 -2586 7424 -2574
rect 7474 -2586 7520 -2574
rect 7588 -2586 7634 -2574
rect 7684 -2586 7730 -2574
rect 7798 -2586 7844 -2574
rect 7894 -2586 7940 -2574
rect 8008 -2586 8054 -2574
rect 8104 -2586 8150 -2574
rect 8218 -2586 8264 -2574
rect 8314 -2586 8360 -2574
rect 8428 -2586 8474 -2574
rect 8524 -2586 8570 -2574
rect 8638 -2586 8684 -2574
rect 8734 -2586 8780 -2574
rect 8848 -2586 8894 -2574
rect 8944 -2586 8990 -2574
rect 9058 -2586 9104 -2574
rect 9154 -2586 9200 -2574
rect 5052 -2633 9158 -2626
rect 4032 -2736 4038 -2674
rect 4032 -2776 4044 -2736
rect 3986 -2782 4044 -2776
rect 5052 -2775 5752 -2633
rect 5786 -2775 6172 -2633
rect 6206 -2775 6592 -2633
rect 6626 -2775 7012 -2633
rect 7046 -2775 7432 -2633
rect 7466 -2775 7852 -2633
rect 7886 -2775 8272 -2633
rect 8306 -2775 8692 -2633
rect 8726 -2775 9112 -2633
rect 9146 -2775 9158 -2633
rect 5052 -2776 9158 -2775
rect 3524 -2826 3570 -2814
rect 3620 -2826 3666 -2814
rect 3734 -2826 3780 -2814
rect 3830 -2826 3876 -2814
rect 3944 -2826 3990 -2814
rect 4040 -2826 4086 -2814
rect 4154 -2826 4200 -2814
rect 4250 -2826 4296 -2814
rect 2580 -3814 2626 -3802
rect 2668 -3814 2714 -3802
rect 2784 -3846 2898 -2878
rect 3500 -3802 3510 -2826
rect 3564 -3802 3574 -2826
rect 3616 -3802 3626 -2826
rect 3774 -3802 3784 -2826
rect 3826 -3802 3836 -2826
rect 3984 -3802 3994 -2826
rect 4036 -3802 4046 -2826
rect 4194 -3802 4204 -2826
rect 4246 -3802 4256 -2826
rect 4310 -3802 4320 -2826
rect 4716 -3238 4726 -2974
rect 5008 -2994 5018 -2974
rect 5052 -2994 5238 -2776
rect 5740 -2781 5798 -2776
rect 6160 -2781 6218 -2776
rect 6580 -2781 6638 -2776
rect 7000 -2781 7058 -2776
rect 7420 -2781 7478 -2776
rect 7840 -2781 7898 -2776
rect 8260 -2781 8318 -2776
rect 8680 -2781 8738 -2776
rect 9100 -2781 9158 -2776
rect 5488 -2834 5534 -2822
rect 5584 -2834 5630 -2822
rect 5698 -2834 5744 -2822
rect 5794 -2834 5840 -2822
rect 5908 -2834 5954 -2822
rect 6004 -2834 6050 -2822
rect 6118 -2834 6164 -2822
rect 6214 -2834 6260 -2822
rect 6328 -2834 6374 -2822
rect 6424 -2834 6470 -2822
rect 6538 -2834 6584 -2822
rect 6634 -2834 6680 -2822
rect 6748 -2834 6794 -2822
rect 6844 -2834 6890 -2822
rect 6958 -2834 7004 -2822
rect 7054 -2834 7100 -2822
rect 7168 -2834 7214 -2822
rect 7264 -2834 7310 -2822
rect 7378 -2834 7424 -2822
rect 7474 -2834 7520 -2822
rect 7588 -2834 7634 -2822
rect 7684 -2834 7730 -2822
rect 7798 -2834 7844 -2822
rect 7894 -2834 7940 -2822
rect 8008 -2834 8054 -2822
rect 8104 -2834 8150 -2822
rect 8218 -2834 8264 -2822
rect 8314 -2834 8360 -2822
rect 8428 -2834 8474 -2822
rect 8524 -2834 8570 -2822
rect 8638 -2834 8684 -2822
rect 8734 -2834 8780 -2822
rect 8848 -2834 8894 -2822
rect 8944 -2834 8990 -2822
rect 9058 -2834 9104 -2822
rect 9154 -2834 9200 -2822
rect 5008 -3210 5238 -2994
rect 5008 -3238 5018 -3210
rect 3524 -3814 3570 -3802
rect 3620 -3814 3666 -3802
rect 3734 -3814 3780 -3802
rect 3830 -3814 3876 -3802
rect 3944 -3814 3990 -3802
rect 4040 -3814 4086 -3802
rect 4154 -3814 4200 -3802
rect 4250 -3814 4296 -3802
rect 2784 -3860 4304 -3846
rect 2784 -3895 3788 -3860
rect 3872 -3894 4208 -3860
rect 4292 -3894 4304 -3860
rect 3822 -3895 4208 -3894
rect 4242 -3895 4304 -3894
rect 2784 -3902 4304 -3895
rect 5052 -3860 5238 -3210
rect 5460 -3810 5470 -2834
rect 5528 -3810 5538 -2834
rect 5580 -3810 5590 -2834
rect 5738 -3810 5748 -2834
rect 5790 -3810 5800 -2834
rect 5948 -3810 5958 -2834
rect 6000 -3810 6010 -2834
rect 6158 -3810 6168 -2834
rect 6210 -3810 6220 -2834
rect 6368 -3810 6378 -2834
rect 6420 -3810 6430 -2834
rect 6578 -3810 6588 -2834
rect 6630 -3810 6640 -2834
rect 6788 -3810 6798 -2834
rect 6840 -3810 6850 -2834
rect 6998 -3810 7008 -2834
rect 7050 -3810 7060 -2834
rect 7208 -3810 7218 -2834
rect 7260 -3810 7270 -2834
rect 7418 -3810 7428 -2834
rect 7470 -3810 7480 -2834
rect 7628 -3810 7638 -2834
rect 7680 -3810 7690 -2834
rect 7838 -3810 7848 -2834
rect 7890 -3810 7900 -2834
rect 8048 -3810 8058 -2834
rect 8100 -3810 8110 -2834
rect 8258 -3810 8268 -2834
rect 8310 -3810 8320 -2834
rect 8468 -3810 8478 -2834
rect 8520 -3810 8530 -2834
rect 8678 -3810 8688 -2834
rect 8730 -3810 8740 -2834
rect 8888 -3810 8898 -2834
rect 8940 -3810 8950 -2834
rect 9098 -3810 9108 -2834
rect 9150 -3810 9160 -2834
rect 9218 -3810 9228 -2834
rect 5488 -3822 5534 -3810
rect 5584 -3822 5630 -3810
rect 5698 -3822 5744 -3810
rect 5794 -3822 5840 -3810
rect 5908 -3822 5954 -3810
rect 6004 -3822 6050 -3810
rect 6118 -3822 6164 -3810
rect 6214 -3822 6260 -3810
rect 6328 -3822 6374 -3810
rect 6424 -3822 6470 -3810
rect 6538 -3822 6584 -3810
rect 6634 -3822 6680 -3810
rect 6748 -3822 6794 -3810
rect 6844 -3822 6890 -3810
rect 6958 -3822 7004 -3810
rect 7054 -3822 7100 -3810
rect 7168 -3822 7214 -3810
rect 7264 -3822 7310 -3810
rect 7378 -3822 7424 -3810
rect 7474 -3822 7520 -3810
rect 7588 -3822 7634 -3810
rect 7684 -3822 7730 -3810
rect 7798 -3822 7844 -3810
rect 7894 -3822 7940 -3810
rect 8008 -3822 8054 -3810
rect 8104 -3822 8150 -3810
rect 8218 -3822 8264 -3810
rect 8314 -3822 8360 -3810
rect 8428 -3822 8474 -3810
rect 8524 -3822 8570 -3810
rect 8638 -3822 8684 -3810
rect 8734 -3822 8780 -3810
rect 8848 -3822 8894 -3810
rect 8944 -3822 8990 -3810
rect 9058 -3822 9104 -3810
rect 9154 -3822 9200 -3810
rect 5052 -3868 9098 -3860
rect 5052 -3903 5542 -3868
rect 5626 -3902 5962 -3868
rect 6046 -3902 6382 -3868
rect 6466 -3902 6802 -3868
rect 6886 -3902 7222 -3868
rect 7306 -3902 7642 -3868
rect 7726 -3902 8062 -3868
rect 8146 -3902 8482 -3868
rect 8566 -3902 8902 -3868
rect 8986 -3902 9098 -3868
rect 5576 -3903 5962 -3902
rect 5996 -3903 6382 -3902
rect 6416 -3903 6802 -3902
rect 6836 -3903 7222 -3902
rect 7256 -3903 7642 -3902
rect 7676 -3903 8062 -3902
rect 8096 -3903 8482 -3902
rect 8516 -3903 8902 -3902
rect 8936 -3903 9098 -3902
rect 5052 -3910 9098 -3903
rect 2938 -3990 3260 -3984
rect 2938 -4272 2950 -3990
rect 3248 -4272 3260 -3990
rect 2938 -4278 3260 -4272
rect 5052 -5746 5238 -3910
rect 5052 -5760 9098 -5746
rect 5052 -5795 5542 -5760
rect 5626 -5794 5962 -5760
rect 6046 -5794 6382 -5760
rect 6466 -5794 6802 -5760
rect 6886 -5794 7222 -5760
rect 7306 -5794 7642 -5760
rect 7726 -5794 8062 -5760
rect 8146 -5794 8482 -5760
rect 8566 -5794 8902 -5760
rect 8986 -5794 9098 -5760
rect 5576 -5795 5962 -5794
rect 5996 -5795 6382 -5794
rect 5052 -5800 6382 -5795
rect 6416 -5800 6802 -5794
rect 6836 -5800 7222 -5794
rect 7256 -5800 7642 -5794
rect 7676 -5800 8062 -5794
rect 8096 -5800 8482 -5794
rect 8516 -5800 8902 -5794
rect 8936 -5800 9098 -5794
rect 5052 -5806 9098 -5800
rect 5052 -6870 5238 -5806
rect 5488 -5850 5534 -5838
rect 5584 -5850 5630 -5838
rect 5698 -5850 5744 -5838
rect 5794 -5850 5840 -5838
rect 5908 -5850 5954 -5838
rect 6004 -5850 6050 -5838
rect 6118 -5850 6164 -5838
rect 6214 -5850 6260 -5838
rect 6328 -5850 6374 -5838
rect 6424 -5850 6470 -5838
rect 6538 -5850 6584 -5838
rect 6634 -5850 6680 -5838
rect 6748 -5850 6794 -5838
rect 6844 -5850 6890 -5838
rect 6958 -5850 7004 -5838
rect 7054 -5850 7100 -5838
rect 7168 -5850 7214 -5838
rect 7264 -5850 7310 -5838
rect 7378 -5850 7424 -5838
rect 7474 -5850 7520 -5838
rect 7588 -5850 7634 -5838
rect 7684 -5850 7730 -5838
rect 7798 -5850 7844 -5838
rect 7894 -5850 7940 -5838
rect 8008 -5850 8054 -5838
rect 8104 -5850 8150 -5838
rect 8218 -5850 8264 -5838
rect 8314 -5850 8360 -5838
rect 8428 -5850 8474 -5838
rect 8524 -5850 8570 -5838
rect 8638 -5850 8684 -5838
rect 8734 -5850 8780 -5838
rect 8848 -5850 8894 -5838
rect 8944 -5850 8990 -5838
rect 9058 -5850 9104 -5838
rect 9154 -5850 9200 -5838
rect 5460 -6826 5470 -5850
rect 5528 -6826 5538 -5850
rect 5580 -6826 5590 -5850
rect 5738 -6826 5748 -5850
rect 5790 -6826 5800 -5850
rect 5948 -6826 5958 -5850
rect 6000 -6826 6010 -5850
rect 6158 -6826 6168 -5850
rect 6210 -6826 6220 -5850
rect 6368 -6826 6378 -5850
rect 6420 -6826 6430 -5850
rect 6578 -6826 6588 -5850
rect 6630 -6826 6640 -5850
rect 6788 -6826 6798 -5850
rect 6840 -6826 6850 -5850
rect 6998 -6826 7008 -5850
rect 7050 -6826 7060 -5850
rect 7208 -6826 7218 -5850
rect 7260 -6826 7270 -5850
rect 7418 -6826 7428 -5850
rect 7470 -6826 7480 -5850
rect 7628 -6826 7638 -5850
rect 7680 -6826 7690 -5850
rect 7838 -6826 7848 -5850
rect 7890 -6826 7900 -5850
rect 8048 -6826 8058 -5850
rect 8100 -6826 8110 -5850
rect 8258 -6826 8268 -5850
rect 8310 -6826 8320 -5850
rect 8468 -6826 8478 -5850
rect 8520 -6826 8530 -5850
rect 8678 -6826 8688 -5850
rect 8730 -6826 8740 -5850
rect 8888 -6826 8898 -5850
rect 8940 -6826 8950 -5850
rect 9098 -6826 9108 -5850
rect 9150 -6826 9160 -5850
rect 9218 -6826 9228 -5850
rect 5488 -6838 5534 -6826
rect 5584 -6838 5630 -6826
rect 5698 -6838 5744 -6826
rect 5794 -6838 5840 -6826
rect 5908 -6838 5954 -6826
rect 6004 -6838 6050 -6826
rect 6118 -6838 6164 -6826
rect 6214 -6838 6260 -6826
rect 6328 -6838 6374 -6826
rect 6424 -6838 6470 -6826
rect 6538 -6838 6584 -6826
rect 6634 -6838 6680 -6826
rect 6748 -6838 6794 -6826
rect 6844 -6838 6890 -6826
rect 6958 -6838 7004 -6826
rect 7054 -6838 7100 -6826
rect 7168 -6838 7214 -6826
rect 7264 -6838 7310 -6826
rect 7378 -6838 7424 -6826
rect 7474 -6838 7520 -6826
rect 7588 -6838 7634 -6826
rect 7684 -6838 7730 -6826
rect 7798 -6838 7844 -6826
rect 7894 -6838 7940 -6826
rect 8008 -6838 8054 -6826
rect 8104 -6838 8150 -6826
rect 8218 -6838 8264 -6826
rect 8314 -6838 8360 -6826
rect 8428 -6838 8474 -6826
rect 8524 -6838 8570 -6826
rect 8638 -6838 8684 -6826
rect 8734 -6838 8780 -6826
rect 8848 -6838 8894 -6826
rect 8944 -6838 8990 -6826
rect 9058 -6838 9104 -6826
rect 9154 -6838 9200 -6826
rect 5052 -6876 9212 -6870
rect 5052 -6884 6172 -6876
rect 6206 -6884 6592 -6876
rect 6626 -6884 7012 -6876
rect 7046 -6884 7432 -6876
rect 7466 -6884 7852 -6876
rect 7886 -6884 8272 -6876
rect 8306 -6884 8692 -6876
rect 8726 -6884 9112 -6876
rect 9146 -6884 9212 -6876
rect 5052 -6918 5752 -6884
rect 5836 -6918 6172 -6884
rect 6256 -6918 6592 -6884
rect 6676 -6918 7012 -6884
rect 7096 -6918 7432 -6884
rect 7516 -6918 7852 -6884
rect 7936 -6918 8272 -6884
rect 8356 -6918 8692 -6884
rect 8776 -6918 9112 -6884
rect 9196 -6918 9212 -6884
rect 5052 -6926 9212 -6918
rect 5478 -7004 5602 -6998
rect 5478 -7104 5490 -7004
rect 5590 -7104 5602 -7004
rect 5478 -7110 5602 -7104
rect 5898 -7004 6022 -6998
rect 5898 -7104 5910 -7004
rect 6010 -7104 6022 -7004
rect 5898 -7110 6022 -7104
rect 6318 -7004 6442 -6998
rect 6318 -7104 6330 -7004
rect 6430 -7104 6442 -7004
rect 6318 -7110 6442 -7104
rect 6738 -7004 6862 -6998
rect 6738 -7104 6750 -7004
rect 6850 -7104 6862 -7004
rect 6738 -7110 6862 -7104
rect 7158 -7004 7282 -6998
rect 7158 -7104 7170 -7004
rect 7270 -7104 7282 -7004
rect 7158 -7110 7282 -7104
rect 7578 -7004 7702 -6998
rect 7578 -7104 7590 -7004
rect 7690 -7104 7702 -7004
rect 7578 -7110 7702 -7104
rect 7998 -7004 8122 -6998
rect 7998 -7104 8010 -7004
rect 8110 -7104 8122 -7004
rect 7998 -7110 8122 -7104
rect 8418 -7004 8542 -6998
rect 8418 -7104 8430 -7004
rect 8530 -7104 8542 -7004
rect 8418 -7110 8542 -7104
rect 8838 -7004 8962 -6998
rect 8838 -7104 8850 -7004
rect 8950 -7104 8962 -7004
rect 8838 -7110 8962 -7104
rect 9164 -7004 9288 -6998
rect 9164 -7104 9176 -7004
rect 9276 -7104 9288 -7004
rect 9164 -7110 9288 -7104
<< via1 >>
rect 10302 13268 10400 13372
rect 10722 13268 10820 13372
rect 11142 13268 11240 13372
rect 11562 13268 11660 13372
rect 11982 13268 12080 13372
rect 12402 13268 12500 13372
rect 12822 13268 12920 13372
rect 13242 13268 13340 13372
rect 13662 13268 13760 13372
rect 14082 13268 14180 13372
rect 14502 13268 14600 13372
rect 14922 13268 15020 13372
rect 15342 13268 15440 13372
rect 15762 13268 15860 13372
rect 16182 13268 16280 13372
rect 16602 13268 16700 13372
rect 17022 13268 17120 13372
rect 17442 13268 17540 13372
rect 17862 13268 17960 13372
rect 18282 13268 18380 13372
rect 18630 13268 18728 13372
rect 10320 12060 10344 13036
rect 10344 12060 10378 13036
rect 10440 12060 10474 13036
rect 10474 12060 10554 13036
rect 10554 12060 10588 13036
rect 10650 12060 10684 13036
rect 10684 12060 10764 13036
rect 10764 12060 10798 13036
rect 10860 12060 10894 13036
rect 10894 12060 10974 13036
rect 10974 12060 11008 13036
rect 11070 12060 11104 13036
rect 11104 12060 11184 13036
rect 11184 12060 11218 13036
rect 11280 12060 11314 13036
rect 11314 12060 11394 13036
rect 11394 12060 11428 13036
rect 11490 12060 11524 13036
rect 11524 12060 11604 13036
rect 11604 12060 11638 13036
rect 11700 12060 11734 13036
rect 11734 12060 11814 13036
rect 11814 12060 11848 13036
rect 11910 12060 11944 13036
rect 11944 12060 12024 13036
rect 12024 12060 12058 13036
rect 12120 12060 12154 13036
rect 12154 12060 12234 13036
rect 12234 12060 12268 13036
rect 12330 12060 12364 13036
rect 12364 12060 12444 13036
rect 12444 12060 12478 13036
rect 12540 12060 12574 13036
rect 12574 12060 12654 13036
rect 12654 12060 12688 13036
rect 12750 12060 12784 13036
rect 12784 12060 12864 13036
rect 12864 12060 12898 13036
rect 12960 12060 12994 13036
rect 12994 12060 13074 13036
rect 13074 12060 13108 13036
rect 13170 12060 13204 13036
rect 13204 12060 13284 13036
rect 13284 12060 13318 13036
rect 13380 12060 13414 13036
rect 13414 12060 13494 13036
rect 13494 12060 13528 13036
rect 13590 12060 13624 13036
rect 13624 12060 13704 13036
rect 13704 12060 13738 13036
rect 13800 12060 13834 13036
rect 13834 12060 13914 13036
rect 13914 12060 13948 13036
rect 14010 12060 14044 13036
rect 14044 12060 14124 13036
rect 14124 12060 14158 13036
rect 14220 12060 14254 13036
rect 14254 12060 14334 13036
rect 14334 12060 14368 13036
rect 14430 12060 14464 13036
rect 14464 12060 14544 13036
rect 14544 12060 14578 13036
rect 14640 12060 14674 13036
rect 14674 12060 14754 13036
rect 14754 12060 14788 13036
rect 14850 12060 14884 13036
rect 14884 12060 14964 13036
rect 14964 12060 14998 13036
rect 15060 12060 15094 13036
rect 15094 12060 15174 13036
rect 15174 12060 15208 13036
rect 15270 12060 15304 13036
rect 15304 12060 15384 13036
rect 15384 12060 15418 13036
rect 15480 12060 15514 13036
rect 15514 12060 15594 13036
rect 15594 12060 15628 13036
rect 15690 12060 15724 13036
rect 15724 12060 15804 13036
rect 15804 12060 15838 13036
rect 15900 12060 15934 13036
rect 15934 12060 16014 13036
rect 16014 12060 16048 13036
rect 16110 12060 16144 13036
rect 16144 12060 16224 13036
rect 16224 12060 16258 13036
rect 16320 12060 16354 13036
rect 16354 12060 16434 13036
rect 16434 12060 16468 13036
rect 16530 12060 16564 13036
rect 16564 12060 16644 13036
rect 16644 12060 16678 13036
rect 16740 12060 16774 13036
rect 16774 12060 16854 13036
rect 16854 12060 16888 13036
rect 16950 12060 16984 13036
rect 16984 12060 17064 13036
rect 17064 12060 17098 13036
rect 17160 12060 17194 13036
rect 17194 12060 17274 13036
rect 17274 12060 17308 13036
rect 17370 12060 17404 13036
rect 17404 12060 17484 13036
rect 17484 12060 17518 13036
rect 17580 12060 17614 13036
rect 17614 12060 17694 13036
rect 17694 12060 17728 13036
rect 17790 12060 17824 13036
rect 17824 12060 17904 13036
rect 17904 12060 17938 13036
rect 18000 12060 18034 13036
rect 18034 12060 18114 13036
rect 18114 12060 18148 13036
rect 18210 12060 18244 13036
rect 18244 12060 18324 13036
rect 18324 12060 18358 13036
rect 18420 12060 18454 13036
rect 18454 12060 18534 13036
rect 18534 12060 18568 13036
rect 18630 12060 18664 13036
rect 18664 12060 18688 13036
rect 10320 10842 10344 11818
rect 10344 10842 10378 11818
rect 10440 10842 10474 11818
rect 10474 10842 10554 11818
rect 10554 10842 10588 11818
rect 10650 10842 10684 11818
rect 10684 10842 10764 11818
rect 10764 10842 10798 11818
rect 10860 10842 10894 11818
rect 10894 10842 10974 11818
rect 10974 10842 11008 11818
rect 11070 10842 11104 11818
rect 11104 10842 11184 11818
rect 11184 10842 11218 11818
rect 11280 10842 11314 11818
rect 11314 10842 11394 11818
rect 11394 10842 11428 11818
rect 11490 10842 11524 11818
rect 11524 10842 11604 11818
rect 11604 10842 11638 11818
rect 11700 10842 11734 11818
rect 11734 10842 11814 11818
rect 11814 10842 11848 11818
rect 11910 10842 11944 11818
rect 11944 10842 12024 11818
rect 12024 10842 12058 11818
rect 12120 10842 12154 11818
rect 12154 10842 12234 11818
rect 12234 10842 12268 11818
rect 12330 10842 12364 11818
rect 12364 10842 12444 11818
rect 12444 10842 12478 11818
rect 12540 10842 12574 11818
rect 12574 10842 12654 11818
rect 12654 10842 12688 11818
rect 12750 10842 12784 11818
rect 12784 10842 12864 11818
rect 12864 10842 12898 11818
rect 12960 10842 12994 11818
rect 12994 10842 13074 11818
rect 13074 10842 13108 11818
rect 13170 10842 13204 11818
rect 13204 10842 13284 11818
rect 13284 10842 13318 11818
rect 13380 10842 13414 11818
rect 13414 10842 13494 11818
rect 13494 10842 13528 11818
rect 13590 10842 13624 11818
rect 13624 10842 13704 11818
rect 13704 10842 13738 11818
rect 13800 10842 13834 11818
rect 13834 10842 13914 11818
rect 13914 10842 13948 11818
rect 14010 10842 14044 11818
rect 14044 10842 14124 11818
rect 14124 10842 14158 11818
rect 14220 10842 14254 11818
rect 14254 10842 14334 11818
rect 14334 10842 14368 11818
rect 14430 10842 14464 11818
rect 14464 10842 14544 11818
rect 14544 10842 14578 11818
rect 14640 10842 14674 11818
rect 14674 10842 14754 11818
rect 14754 10842 14788 11818
rect 14850 10842 14884 11818
rect 14884 10842 14964 11818
rect 14964 10842 14998 11818
rect 15060 10842 15094 11818
rect 15094 10842 15174 11818
rect 15174 10842 15208 11818
rect 15270 10842 15304 11818
rect 15304 10842 15384 11818
rect 15384 10842 15418 11818
rect 15480 10842 15514 11818
rect 15514 10842 15594 11818
rect 15594 10842 15628 11818
rect 15690 10842 15724 11818
rect 15724 10842 15804 11818
rect 15804 10842 15838 11818
rect 15900 10842 15934 11818
rect 15934 10842 16014 11818
rect 16014 10842 16048 11818
rect 16110 10842 16144 11818
rect 16144 10842 16224 11818
rect 16224 10842 16258 11818
rect 16320 10842 16354 11818
rect 16354 10842 16434 11818
rect 16434 10842 16468 11818
rect 16530 10842 16564 11818
rect 16564 10842 16644 11818
rect 16644 10842 16678 11818
rect 16740 10842 16774 11818
rect 16774 10842 16854 11818
rect 16854 10842 16888 11818
rect 16950 10842 16984 11818
rect 16984 10842 17064 11818
rect 17064 10842 17098 11818
rect 17160 10842 17194 11818
rect 17194 10842 17274 11818
rect 17274 10842 17308 11818
rect 17370 10842 17404 11818
rect 17404 10842 17484 11818
rect 17484 10842 17518 11818
rect 17580 10842 17614 11818
rect 17614 10842 17694 11818
rect 17694 10842 17728 11818
rect 17790 10842 17824 11818
rect 17824 10842 17904 11818
rect 17904 10842 17938 11818
rect 18000 10842 18034 11818
rect 18034 10842 18114 11818
rect 18114 10842 18148 11818
rect 18210 10842 18244 11818
rect 18244 10842 18324 11818
rect 18324 10842 18358 11818
rect 18420 10842 18454 11818
rect 18454 10842 18534 11818
rect 18534 10842 18568 11818
rect 18630 10842 18664 11818
rect 18664 10842 18688 11818
rect 5490 7130 5590 7230
rect 5910 7130 6010 7230
rect 6330 7130 6430 7230
rect 6750 7130 6850 7230
rect 7170 7130 7270 7230
rect 7590 7130 7690 7230
rect 8010 7130 8110 7230
rect 8430 7130 8530 7230
rect 8850 7130 8950 7230
rect 9176 7130 9276 7230
rect 5470 5976 5494 6952
rect 5494 5976 5528 6952
rect 5590 5976 5624 6952
rect 5624 5976 5704 6952
rect 5704 5976 5738 6952
rect 5800 5976 5834 6952
rect 5834 5976 5914 6952
rect 5914 5976 5948 6952
rect 6010 5976 6044 6952
rect 6044 5976 6124 6952
rect 6124 5976 6158 6952
rect 6220 5976 6254 6952
rect 6254 5976 6334 6952
rect 6334 5976 6368 6952
rect 6430 5976 6464 6952
rect 6464 5976 6544 6952
rect 6544 5976 6578 6952
rect 6640 5976 6674 6952
rect 6674 5976 6754 6952
rect 6754 5976 6788 6952
rect 6850 5976 6884 6952
rect 6884 5976 6964 6952
rect 6964 5976 6998 6952
rect 7060 5976 7094 6952
rect 7094 5976 7174 6952
rect 7174 5976 7208 6952
rect 7270 5976 7304 6952
rect 7304 5976 7384 6952
rect 7384 5976 7418 6952
rect 7480 5976 7514 6952
rect 7514 5976 7594 6952
rect 7594 5976 7628 6952
rect 7690 5976 7724 6952
rect 7724 5976 7804 6952
rect 7804 5976 7838 6952
rect 7900 5976 7934 6952
rect 7934 5976 8014 6952
rect 8014 5976 8048 6952
rect 8110 5976 8144 6952
rect 8144 5976 8224 6952
rect 8224 5976 8258 6952
rect 8320 5976 8354 6952
rect 8354 5976 8434 6952
rect 8434 5976 8468 6952
rect 8530 5976 8564 6952
rect 8564 5976 8644 6952
rect 8644 5976 8678 6952
rect 8740 5976 8774 6952
rect 8774 5976 8854 6952
rect 8854 5976 8888 6952
rect 8950 5976 8984 6952
rect 8984 5976 9064 6952
rect 9064 5976 9098 6952
rect 9160 5976 9194 6952
rect 9194 5976 9218 6952
rect 10320 6832 10344 7808
rect 10344 6832 10378 7808
rect 10440 6832 10474 7808
rect 10474 6832 10554 7808
rect 10554 6832 10588 7808
rect 10650 6832 10684 7808
rect 10684 6832 10764 7808
rect 10764 6832 10798 7808
rect 10860 6832 10894 7808
rect 10894 6832 10974 7808
rect 10974 6832 11008 7808
rect 11070 6832 11104 7808
rect 11104 6832 11184 7808
rect 11184 6832 11218 7808
rect 11280 6832 11314 7808
rect 11314 6832 11394 7808
rect 11394 6832 11428 7808
rect 11490 6832 11524 7808
rect 11524 6832 11604 7808
rect 11604 6832 11638 7808
rect 11700 6832 11734 7808
rect 11734 6832 11814 7808
rect 11814 6832 11848 7808
rect 11910 6832 11944 7808
rect 11944 6832 12024 7808
rect 12024 6832 12058 7808
rect 12120 6832 12154 7808
rect 12154 6832 12234 7808
rect 12234 6832 12268 7808
rect 12330 6832 12364 7808
rect 12364 6832 12444 7808
rect 12444 6832 12478 7808
rect 12540 6832 12574 7808
rect 12574 6832 12654 7808
rect 12654 6832 12688 7808
rect 12750 6832 12784 7808
rect 12784 6832 12864 7808
rect 12864 6832 12898 7808
rect 12960 6832 12994 7808
rect 12994 6832 13074 7808
rect 13074 6832 13108 7808
rect 13170 6832 13204 7808
rect 13204 6832 13284 7808
rect 13284 6832 13318 7808
rect 13380 6832 13414 7808
rect 13414 6832 13494 7808
rect 13494 6832 13528 7808
rect 13590 6832 13624 7808
rect 13624 6832 13704 7808
rect 13704 6832 13738 7808
rect 13800 6832 13834 7808
rect 13834 6832 13914 7808
rect 13914 6832 13948 7808
rect 14010 6832 14044 7808
rect 14044 6832 14124 7808
rect 14124 6832 14158 7808
rect 14220 6832 14254 7808
rect 14254 6832 14334 7808
rect 14334 6832 14368 7808
rect 14430 6832 14464 7808
rect 14464 6832 14544 7808
rect 14544 6832 14578 7808
rect 14640 6832 14674 7808
rect 14674 6832 14754 7808
rect 14754 6832 14788 7808
rect 14850 6832 14884 7808
rect 14884 6832 14964 7808
rect 14964 6832 14998 7808
rect 15060 6832 15094 7808
rect 15094 6832 15174 7808
rect 15174 6832 15208 7808
rect 15270 6832 15304 7808
rect 15304 6832 15384 7808
rect 15384 6832 15418 7808
rect 15480 6832 15514 7808
rect 15514 6832 15594 7808
rect 15594 6832 15628 7808
rect 15690 6832 15724 7808
rect 15724 6832 15804 7808
rect 15804 6832 15838 7808
rect 15900 6832 15934 7808
rect 15934 6832 16014 7808
rect 16014 6832 16048 7808
rect 16110 6832 16144 7808
rect 16144 6832 16224 7808
rect 16224 6832 16258 7808
rect 16320 6832 16354 7808
rect 16354 6832 16434 7808
rect 16434 6832 16468 7808
rect 16530 6832 16564 7808
rect 16564 6832 16644 7808
rect 16644 6832 16678 7808
rect 16740 6832 16774 7808
rect 16774 6832 16854 7808
rect 16854 6832 16888 7808
rect 16950 6832 16984 7808
rect 16984 6832 17064 7808
rect 17064 6832 17098 7808
rect 17160 6832 17194 7808
rect 17194 6832 17274 7808
rect 17274 6832 17308 7808
rect 17370 6832 17404 7808
rect 17404 6832 17484 7808
rect 17484 6832 17518 7808
rect 17580 6832 17614 7808
rect 17614 6832 17694 7808
rect 17694 6832 17728 7808
rect 17790 6832 17824 7808
rect 17824 6832 17904 7808
rect 17904 6832 17938 7808
rect 18000 6832 18034 7808
rect 18034 6832 18114 7808
rect 18114 6832 18148 7808
rect 18210 6832 18244 7808
rect 18244 6832 18324 7808
rect 18324 6832 18358 7808
rect 18420 6832 18454 7808
rect 18454 6832 18534 7808
rect 18534 6832 18568 7808
rect 18630 6832 18664 7808
rect 18664 6832 18688 7808
rect 2950 5516 3248 5798
rect 2566 4352 2586 5328
rect 2586 4352 2620 5328
rect 2674 4352 2708 5328
rect 2708 4352 2728 5328
rect 2794 4256 2936 4404
rect 3510 4352 3530 5328
rect 3530 4352 3564 5328
rect 3626 4352 3660 5328
rect 3660 4352 3740 5328
rect 3740 4352 3774 5328
rect 3836 4352 3870 5328
rect 3870 4352 3950 5328
rect 3950 4352 3984 5328
rect 4046 4352 4080 5328
rect 4080 4352 4160 5328
rect 4160 4352 4194 5328
rect 4256 4352 4290 5328
rect 4290 4352 4310 5328
rect 4726 4500 5008 4764
rect 9326 5378 9936 5996
rect 10320 5596 10344 6572
rect 10344 5596 10378 6572
rect 10440 5596 10474 6572
rect 10474 5596 10554 6572
rect 10554 5596 10588 6572
rect 10650 5596 10684 6572
rect 10684 5596 10764 6572
rect 10764 5596 10798 6572
rect 10860 5596 10894 6572
rect 10894 5596 10974 6572
rect 10974 5596 11008 6572
rect 11070 5596 11104 6572
rect 11104 5596 11184 6572
rect 11184 5596 11218 6572
rect 11280 5596 11314 6572
rect 11314 5596 11394 6572
rect 11394 5596 11428 6572
rect 11490 5596 11524 6572
rect 11524 5596 11604 6572
rect 11604 5596 11638 6572
rect 11700 5596 11734 6572
rect 11734 5596 11814 6572
rect 11814 5596 11848 6572
rect 11910 5596 11944 6572
rect 11944 5596 12024 6572
rect 12024 5596 12058 6572
rect 12120 5596 12154 6572
rect 12154 5596 12234 6572
rect 12234 5596 12268 6572
rect 12330 5596 12364 6572
rect 12364 5596 12444 6572
rect 12444 5596 12478 6572
rect 12540 5596 12574 6572
rect 12574 5596 12654 6572
rect 12654 5596 12688 6572
rect 12750 5596 12784 6572
rect 12784 5596 12864 6572
rect 12864 5596 12898 6572
rect 12960 5596 12994 6572
rect 12994 5596 13074 6572
rect 13074 5596 13108 6572
rect 13170 5596 13204 6572
rect 13204 5596 13284 6572
rect 13284 5596 13318 6572
rect 13380 5596 13414 6572
rect 13414 5596 13494 6572
rect 13494 5596 13528 6572
rect 13590 5596 13624 6572
rect 13624 5596 13704 6572
rect 13704 5596 13738 6572
rect 13800 5596 13834 6572
rect 13834 5596 13914 6572
rect 13914 5596 13948 6572
rect 14010 5596 14044 6572
rect 14044 5596 14124 6572
rect 14124 5596 14158 6572
rect 14220 5596 14254 6572
rect 14254 5596 14334 6572
rect 14334 5596 14368 6572
rect 14430 5596 14464 6572
rect 14464 5596 14544 6572
rect 14544 5596 14578 6572
rect 14640 5596 14674 6572
rect 14674 5596 14754 6572
rect 14754 5596 14788 6572
rect 14850 5596 14884 6572
rect 14884 5596 14964 6572
rect 14964 5596 14998 6572
rect 15060 5596 15094 6572
rect 15094 5596 15174 6572
rect 15174 5596 15208 6572
rect 15270 5596 15304 6572
rect 15304 5596 15384 6572
rect 15384 5596 15418 6572
rect 15480 5596 15514 6572
rect 15514 5596 15594 6572
rect 15594 5596 15628 6572
rect 15690 5596 15724 6572
rect 15724 5596 15804 6572
rect 15804 5596 15838 6572
rect 15900 5596 15934 6572
rect 15934 5596 16014 6572
rect 16014 5596 16048 6572
rect 16110 5596 16144 6572
rect 16144 5596 16224 6572
rect 16224 5596 16258 6572
rect 16320 5596 16354 6572
rect 16354 5596 16434 6572
rect 16434 5596 16468 6572
rect 16530 5596 16564 6572
rect 16564 5596 16644 6572
rect 16644 5596 16678 6572
rect 16740 5596 16774 6572
rect 16774 5596 16854 6572
rect 16854 5596 16888 6572
rect 16950 5596 16984 6572
rect 16984 5596 17064 6572
rect 17064 5596 17098 6572
rect 17160 5596 17194 6572
rect 17194 5596 17274 6572
rect 17274 5596 17308 6572
rect 17370 5596 17404 6572
rect 17404 5596 17484 6572
rect 17484 5596 17518 6572
rect 17580 5596 17614 6572
rect 17614 5596 17694 6572
rect 17694 5596 17728 6572
rect 17790 5596 17824 6572
rect 17824 5596 17904 6572
rect 17904 5596 17938 6572
rect 18000 5596 18034 6572
rect 18034 5596 18114 6572
rect 18114 5596 18148 6572
rect 18210 5596 18244 6572
rect 18244 5596 18324 6572
rect 18324 5596 18358 6572
rect 18420 5596 18454 6572
rect 18454 5596 18534 6572
rect 18534 5596 18568 6572
rect 18630 5596 18664 6572
rect 18664 5596 18688 6572
rect 2544 3124 2582 4100
rect 2582 3124 2616 4100
rect 2668 3124 2678 4100
rect 2678 3124 2712 4100
rect 2712 3124 2722 4100
rect 2774 3124 2808 4100
rect 2808 3124 2846 4100
rect 5470 4360 5494 5336
rect 5494 4360 5528 5336
rect 5590 4360 5624 5336
rect 5624 4360 5704 5336
rect 5704 4360 5738 5336
rect 5800 4360 5834 5336
rect 5834 4360 5914 5336
rect 5914 4360 5948 5336
rect 6010 4360 6044 5336
rect 6044 4360 6124 5336
rect 6124 4360 6158 5336
rect 6220 4360 6254 5336
rect 6254 4360 6334 5336
rect 6334 4360 6368 5336
rect 6430 4360 6464 5336
rect 6464 4360 6544 5336
rect 6544 4360 6578 5336
rect 6640 4360 6674 5336
rect 6674 4360 6754 5336
rect 6754 4360 6788 5336
rect 6850 4360 6884 5336
rect 6884 4360 6964 5336
rect 6964 4360 6998 5336
rect 7060 4360 7094 5336
rect 7094 4360 7174 5336
rect 7174 4360 7208 5336
rect 7270 4360 7304 5336
rect 7304 4360 7384 5336
rect 7384 4360 7418 5336
rect 7480 4360 7514 5336
rect 7514 4360 7594 5336
rect 7594 4360 7628 5336
rect 7690 4360 7724 5336
rect 7724 4360 7804 5336
rect 7804 4360 7838 5336
rect 7900 4360 7934 5336
rect 7934 4360 8014 5336
rect 8014 4360 8048 5336
rect 8110 4360 8144 5336
rect 8144 4360 8224 5336
rect 8224 4360 8258 5336
rect 8320 4360 8354 5336
rect 8354 4360 8434 5336
rect 8434 4360 8468 5336
rect 8530 4360 8564 5336
rect 8564 4360 8644 5336
rect 8644 4360 8678 5336
rect 8740 4360 8774 5336
rect 8774 4360 8854 5336
rect 8854 4360 8888 5336
rect 8950 4360 8984 5336
rect 8984 4360 9064 5336
rect 9064 4360 9098 5336
rect 9160 4360 9194 5336
rect 9194 4360 9218 5336
rect 10320 4360 10344 5336
rect 10344 4360 10378 5336
rect 10440 4360 10474 5336
rect 10474 4360 10554 5336
rect 10554 4360 10588 5336
rect 10650 4360 10684 5336
rect 10684 4360 10764 5336
rect 10764 4360 10798 5336
rect 10860 4360 10894 5336
rect 10894 4360 10974 5336
rect 10974 4360 11008 5336
rect 11070 4360 11104 5336
rect 11104 4360 11184 5336
rect 11184 4360 11218 5336
rect 11280 4360 11314 5336
rect 11314 4360 11394 5336
rect 11394 4360 11428 5336
rect 11490 4360 11524 5336
rect 11524 4360 11604 5336
rect 11604 4360 11638 5336
rect 11700 4360 11734 5336
rect 11734 4360 11814 5336
rect 11814 4360 11848 5336
rect 11910 4360 11944 5336
rect 11944 4360 12024 5336
rect 12024 4360 12058 5336
rect 12120 4360 12154 5336
rect 12154 4360 12234 5336
rect 12234 4360 12268 5336
rect 12330 4360 12364 5336
rect 12364 4360 12444 5336
rect 12444 4360 12478 5336
rect 12540 4360 12574 5336
rect 12574 4360 12654 5336
rect 12654 4360 12688 5336
rect 12750 4360 12784 5336
rect 12784 4360 12864 5336
rect 12864 4360 12898 5336
rect 12960 4360 12994 5336
rect 12994 4360 13074 5336
rect 13074 4360 13108 5336
rect 13170 4360 13204 5336
rect 13204 4360 13284 5336
rect 13284 4360 13318 5336
rect 13380 4360 13414 5336
rect 13414 4360 13494 5336
rect 13494 4360 13528 5336
rect 13590 4360 13624 5336
rect 13624 4360 13704 5336
rect 13704 4360 13738 5336
rect 13800 4360 13834 5336
rect 13834 4360 13914 5336
rect 13914 4360 13948 5336
rect 14010 4360 14044 5336
rect 14044 4360 14124 5336
rect 14124 4360 14158 5336
rect 14220 4360 14254 5336
rect 14254 4360 14334 5336
rect 14334 4360 14368 5336
rect 14430 4360 14464 5336
rect 14464 4360 14544 5336
rect 14544 4360 14578 5336
rect 14640 4360 14674 5336
rect 14674 4360 14754 5336
rect 14754 4360 14788 5336
rect 14850 4360 14884 5336
rect 14884 4360 14964 5336
rect 14964 4360 14998 5336
rect 15060 4360 15094 5336
rect 15094 4360 15174 5336
rect 15174 4360 15208 5336
rect 15270 4360 15304 5336
rect 15304 4360 15384 5336
rect 15384 4360 15418 5336
rect 15480 4360 15514 5336
rect 15514 4360 15594 5336
rect 15594 4360 15628 5336
rect 15690 4360 15724 5336
rect 15724 4360 15804 5336
rect 15804 4360 15838 5336
rect 15900 4360 15934 5336
rect 15934 4360 16014 5336
rect 16014 4360 16048 5336
rect 16110 4360 16144 5336
rect 16144 4360 16224 5336
rect 16224 4360 16258 5336
rect 16320 4360 16354 5336
rect 16354 4360 16434 5336
rect 16434 4360 16468 5336
rect 16530 4360 16564 5336
rect 16564 4360 16644 5336
rect 16644 4360 16678 5336
rect 16740 4360 16774 5336
rect 16774 4360 16854 5336
rect 16854 4360 16888 5336
rect 16950 4360 16984 5336
rect 16984 4360 17064 5336
rect 17064 4360 17098 5336
rect 17160 4360 17194 5336
rect 17194 4360 17274 5336
rect 17274 4360 17308 5336
rect 17370 4360 17404 5336
rect 17404 4360 17484 5336
rect 17484 4360 17518 5336
rect 17580 4360 17614 5336
rect 17614 4360 17694 5336
rect 17694 4360 17728 5336
rect 17790 4360 17824 5336
rect 17824 4360 17904 5336
rect 17904 4360 17938 5336
rect 18000 4360 18034 5336
rect 18034 4360 18114 5336
rect 18114 4360 18148 5336
rect 18210 4360 18244 5336
rect 18244 4360 18324 5336
rect 18324 4360 18358 5336
rect 18420 4360 18454 5336
rect 18454 4360 18534 5336
rect 18534 4360 18568 5336
rect 18630 4360 18664 5336
rect 18664 4360 18688 5336
rect 3296 3124 3320 4100
rect 3320 3124 3354 4100
rect 3416 3124 3450 4100
rect 3450 3124 3530 4100
rect 3530 3124 3564 4100
rect 3626 3124 3660 4100
rect 3660 3124 3740 4100
rect 3740 3124 3774 4100
rect 3836 3124 3870 4100
rect 3870 3124 3950 4100
rect 3950 3124 3984 4100
rect 4046 3124 4080 4100
rect 4080 3124 4160 4100
rect 4160 3124 4194 4100
rect 4256 3124 4290 4100
rect 4290 3124 4370 4100
rect 4370 3124 4404 4100
rect 4466 3124 4500 4100
rect 4500 3124 4580 4100
rect 4580 3124 4614 4100
rect 4676 3124 4710 4100
rect 4710 3124 4790 4100
rect 4790 3124 4824 4100
rect 4886 3124 4920 4100
rect 4920 3124 4944 4100
rect 5470 3124 5494 4100
rect 5494 3124 5528 4100
rect 5590 3124 5624 4100
rect 5624 3124 5704 4100
rect 5704 3124 5738 4100
rect 5800 3124 5834 4100
rect 5834 3124 5914 4100
rect 5914 3124 5948 4100
rect 6010 3124 6044 4100
rect 6044 3124 6124 4100
rect 6124 3124 6158 4100
rect 6220 3124 6254 4100
rect 6254 3124 6334 4100
rect 6334 3124 6368 4100
rect 6430 3124 6464 4100
rect 6464 3124 6544 4100
rect 6544 3124 6578 4100
rect 6640 3124 6674 4100
rect 6674 3124 6754 4100
rect 6754 3124 6788 4100
rect 6850 3124 6884 4100
rect 6884 3124 6964 4100
rect 6964 3124 6998 4100
rect 7060 3124 7094 4100
rect 7094 3124 7174 4100
rect 7174 3124 7208 4100
rect 7270 3124 7304 4100
rect 7304 3124 7384 4100
rect 7384 3124 7418 4100
rect 7480 3124 7514 4100
rect 7514 3124 7594 4100
rect 7594 3124 7628 4100
rect 7690 3124 7724 4100
rect 7724 3124 7804 4100
rect 7804 3124 7838 4100
rect 7900 3124 7934 4100
rect 7934 3124 8014 4100
rect 8014 3124 8048 4100
rect 8110 3124 8144 4100
rect 8144 3124 8224 4100
rect 8224 3124 8258 4100
rect 8320 3124 8354 4100
rect 8354 3124 8434 4100
rect 8434 3124 8468 4100
rect 8530 3124 8564 4100
rect 8564 3124 8644 4100
rect 8644 3124 8678 4100
rect 8740 3124 8774 4100
rect 8774 3124 8854 4100
rect 8854 3124 8888 4100
rect 8950 3124 8984 4100
rect 8984 3124 9064 4100
rect 9064 3124 9098 4100
rect 9160 3124 9194 4100
rect 9194 3124 9218 4100
rect 10320 3124 10344 4100
rect 10344 3124 10378 4100
rect 10440 3124 10474 4100
rect 10474 3124 10554 4100
rect 10554 3124 10588 4100
rect 10650 3124 10684 4100
rect 10684 3124 10764 4100
rect 10764 3124 10798 4100
rect 10860 3124 10894 4100
rect 10894 3124 10974 4100
rect 10974 3124 11008 4100
rect 11070 3124 11104 4100
rect 11104 3124 11184 4100
rect 11184 3124 11218 4100
rect 11280 3124 11314 4100
rect 11314 3124 11394 4100
rect 11394 3124 11428 4100
rect 11490 3124 11524 4100
rect 11524 3124 11604 4100
rect 11604 3124 11638 4100
rect 11700 3124 11734 4100
rect 11734 3124 11814 4100
rect 11814 3124 11848 4100
rect 11910 3124 11944 4100
rect 11944 3124 12024 4100
rect 12024 3124 12058 4100
rect 12120 3124 12154 4100
rect 12154 3124 12234 4100
rect 12234 3124 12268 4100
rect 12330 3124 12364 4100
rect 12364 3124 12444 4100
rect 12444 3124 12478 4100
rect 12540 3124 12574 4100
rect 12574 3124 12654 4100
rect 12654 3124 12688 4100
rect 12750 3124 12784 4100
rect 12784 3124 12864 4100
rect 12864 3124 12898 4100
rect 12960 3124 12994 4100
rect 12994 3124 13074 4100
rect 13074 3124 13108 4100
rect 13170 3124 13204 4100
rect 13204 3124 13284 4100
rect 13284 3124 13318 4100
rect 13380 3124 13414 4100
rect 13414 3124 13494 4100
rect 13494 3124 13528 4100
rect 13590 3124 13624 4100
rect 13624 3124 13704 4100
rect 13704 3124 13738 4100
rect 13800 3124 13834 4100
rect 13834 3124 13914 4100
rect 13914 3124 13948 4100
rect 14010 3124 14044 4100
rect 14044 3124 14124 4100
rect 14124 3124 14158 4100
rect 14220 3124 14254 4100
rect 14254 3124 14334 4100
rect 14334 3124 14368 4100
rect 14430 3124 14464 4100
rect 14464 3124 14544 4100
rect 14544 3124 14578 4100
rect 14640 3124 14674 4100
rect 14674 3124 14754 4100
rect 14754 3124 14788 4100
rect 14850 3124 14884 4100
rect 14884 3124 14964 4100
rect 14964 3124 14998 4100
rect 15060 3124 15094 4100
rect 15094 3124 15174 4100
rect 15174 3124 15208 4100
rect 15270 3124 15304 4100
rect 15304 3124 15384 4100
rect 15384 3124 15418 4100
rect 15480 3124 15514 4100
rect 15514 3124 15594 4100
rect 15594 3124 15628 4100
rect 15690 3124 15724 4100
rect 15724 3124 15804 4100
rect 15804 3124 15838 4100
rect 15900 3124 15934 4100
rect 15934 3124 16014 4100
rect 16014 3124 16048 4100
rect 16110 3124 16144 4100
rect 16144 3124 16224 4100
rect 16224 3124 16258 4100
rect 16320 3124 16354 4100
rect 16354 3124 16434 4100
rect 16434 3124 16468 4100
rect 16530 3124 16564 4100
rect 16564 3124 16644 4100
rect 16644 3124 16678 4100
rect 16740 3124 16774 4100
rect 16774 3124 16854 4100
rect 16854 3124 16888 4100
rect 16950 3124 16984 4100
rect 16984 3124 17064 4100
rect 17064 3124 17098 4100
rect 17160 3124 17194 4100
rect 17194 3124 17274 4100
rect 17274 3124 17308 4100
rect 17370 3124 17404 4100
rect 17404 3124 17484 4100
rect 17484 3124 17518 4100
rect 17580 3124 17614 4100
rect 17614 3124 17694 4100
rect 17694 3124 17728 4100
rect 17790 3124 17824 4100
rect 17824 3124 17904 4100
rect 17904 3124 17938 4100
rect 18000 3124 18034 4100
rect 18034 3124 18114 4100
rect 18114 3124 18148 4100
rect 18210 3124 18244 4100
rect 18244 3124 18324 4100
rect 18324 3124 18358 4100
rect 18420 3124 18454 4100
rect 18454 3124 18534 4100
rect 18534 3124 18568 4100
rect 18630 3124 18664 4100
rect 18664 3124 18688 4100
rect 196 2220 524 2482
rect 2984 2690 3128 2838
rect -188 1400 -114 1458
rect 4386 1286 4630 1534
rect -26 -14 36 40
rect 5366 2870 5466 2970
rect 5786 2870 5886 2970
rect 6206 2870 6306 2970
rect 6626 2870 6726 2970
rect 7046 2870 7146 2970
rect 7466 2870 7566 2970
rect 7886 2870 7986 2970
rect 8306 2870 8406 2970
rect 8726 2870 8826 2970
rect 9146 2870 9246 2970
rect 10208 2854 10308 2954
rect 10628 2854 10728 2954
rect 11048 2854 11148 2954
rect 11468 2854 11568 2954
rect 11888 2854 11988 2954
rect 12308 2854 12408 2954
rect 12728 2854 12828 2954
rect 13148 2854 13248 2954
rect 13568 2854 13668 2954
rect 13988 2854 14088 2954
rect 14408 2854 14508 2954
rect 14828 2854 14928 2954
rect 15248 2854 15348 2954
rect 15668 2854 15768 2954
rect 16088 2854 16188 2954
rect 16508 2854 16608 2954
rect 16928 2854 17028 2954
rect 17348 2854 17448 2954
rect 17768 2854 17868 2954
rect 18188 2854 18288 2954
rect 18608 2854 18708 2954
rect 5020 -26 5264 222
rect 196 -956 524 -694
rect 2984 -1312 3128 -1164
rect 5366 -1444 5466 -1344
rect 5786 -1444 5886 -1344
rect 6206 -1444 6306 -1344
rect 6626 -1444 6726 -1344
rect 7046 -1444 7146 -1344
rect 7466 -1444 7566 -1344
rect 7886 -1444 7986 -1344
rect 8306 -1444 8406 -1344
rect 8726 -1444 8826 -1344
rect 9146 -1444 9246 -1344
rect 2544 -2574 2582 -1598
rect 2582 -2574 2616 -1598
rect 2668 -2574 2678 -1598
rect 2678 -2574 2712 -1598
rect 2712 -2574 2722 -1598
rect 2774 -2574 2808 -1598
rect 2808 -2574 2846 -1598
rect 3296 -2574 3320 -1598
rect 3320 -2574 3354 -1598
rect 3416 -2574 3450 -1598
rect 3450 -2574 3530 -1598
rect 3530 -2574 3564 -1598
rect 3626 -2574 3660 -1598
rect 3660 -2574 3740 -1598
rect 3740 -2574 3774 -1598
rect 3836 -2574 3870 -1598
rect 3870 -2574 3950 -1598
rect 3950 -2574 3984 -1598
rect 4046 -2574 4080 -1598
rect 4080 -2574 4160 -1598
rect 4160 -2574 4194 -1598
rect 4256 -2574 4290 -1598
rect 4290 -2574 4370 -1598
rect 4370 -2574 4404 -1598
rect 4466 -2574 4500 -1598
rect 4500 -2574 4580 -1598
rect 4580 -2574 4614 -1598
rect 4676 -2574 4710 -1598
rect 4710 -2574 4790 -1598
rect 4790 -2574 4824 -1598
rect 4886 -2574 4920 -1598
rect 4920 -2574 4944 -1598
rect 2566 -3802 2586 -2826
rect 2586 -3802 2620 -2826
rect 2674 -3802 2708 -2826
rect 2708 -3802 2728 -2826
rect 2794 -2878 2936 -2730
rect 5470 -2574 5494 -1598
rect 5494 -2574 5528 -1598
rect 5590 -2574 5624 -1598
rect 5624 -2574 5704 -1598
rect 5704 -2574 5738 -1598
rect 5800 -2574 5834 -1598
rect 5834 -2574 5914 -1598
rect 5914 -2574 5948 -1598
rect 6010 -2574 6044 -1598
rect 6044 -2574 6124 -1598
rect 6124 -2574 6158 -1598
rect 6220 -2574 6254 -1598
rect 6254 -2574 6334 -1598
rect 6334 -2574 6368 -1598
rect 6430 -2574 6464 -1598
rect 6464 -2574 6544 -1598
rect 6544 -2574 6578 -1598
rect 6640 -2574 6674 -1598
rect 6674 -2574 6754 -1598
rect 6754 -2574 6788 -1598
rect 6850 -2574 6884 -1598
rect 6884 -2574 6964 -1598
rect 6964 -2574 6998 -1598
rect 7060 -2574 7094 -1598
rect 7094 -2574 7174 -1598
rect 7174 -2574 7208 -1598
rect 7270 -2574 7304 -1598
rect 7304 -2574 7384 -1598
rect 7384 -2574 7418 -1598
rect 7480 -2574 7514 -1598
rect 7514 -2574 7594 -1598
rect 7594 -2574 7628 -1598
rect 7690 -2574 7724 -1598
rect 7724 -2574 7804 -1598
rect 7804 -2574 7838 -1598
rect 7900 -2574 7934 -1598
rect 7934 -2574 8014 -1598
rect 8014 -2574 8048 -1598
rect 8110 -2574 8144 -1598
rect 8144 -2574 8224 -1598
rect 8224 -2574 8258 -1598
rect 8320 -2574 8354 -1598
rect 8354 -2574 8434 -1598
rect 8434 -2574 8468 -1598
rect 8530 -2574 8564 -1598
rect 8564 -2574 8644 -1598
rect 8644 -2574 8678 -1598
rect 8740 -2574 8774 -1598
rect 8774 -2574 8854 -1598
rect 8854 -2574 8888 -1598
rect 8950 -2574 8984 -1598
rect 8984 -2574 9064 -1598
rect 9064 -2574 9098 -1598
rect 9160 -2574 9194 -1598
rect 9194 -2574 9218 -1598
rect 3510 -3802 3530 -2826
rect 3530 -3802 3564 -2826
rect 3626 -3802 3660 -2826
rect 3660 -3802 3740 -2826
rect 3740 -3802 3774 -2826
rect 3836 -3802 3870 -2826
rect 3870 -3802 3950 -2826
rect 3950 -3802 3984 -2826
rect 4046 -3802 4080 -2826
rect 4080 -3802 4160 -2826
rect 4160 -3802 4194 -2826
rect 4256 -3802 4290 -2826
rect 4290 -3802 4310 -2826
rect 4726 -3238 5008 -2974
rect 5470 -3810 5494 -2834
rect 5494 -3810 5528 -2834
rect 5590 -3810 5624 -2834
rect 5624 -3810 5704 -2834
rect 5704 -3810 5738 -2834
rect 5800 -3810 5834 -2834
rect 5834 -3810 5914 -2834
rect 5914 -3810 5948 -2834
rect 6010 -3810 6044 -2834
rect 6044 -3810 6124 -2834
rect 6124 -3810 6158 -2834
rect 6220 -3810 6254 -2834
rect 6254 -3810 6334 -2834
rect 6334 -3810 6368 -2834
rect 6430 -3810 6464 -2834
rect 6464 -3810 6544 -2834
rect 6544 -3810 6578 -2834
rect 6640 -3810 6674 -2834
rect 6674 -3810 6754 -2834
rect 6754 -3810 6788 -2834
rect 6850 -3810 6884 -2834
rect 6884 -3810 6964 -2834
rect 6964 -3810 6998 -2834
rect 7060 -3810 7094 -2834
rect 7094 -3810 7174 -2834
rect 7174 -3810 7208 -2834
rect 7270 -3810 7304 -2834
rect 7304 -3810 7384 -2834
rect 7384 -3810 7418 -2834
rect 7480 -3810 7514 -2834
rect 7514 -3810 7594 -2834
rect 7594 -3810 7628 -2834
rect 7690 -3810 7724 -2834
rect 7724 -3810 7804 -2834
rect 7804 -3810 7838 -2834
rect 7900 -3810 7934 -2834
rect 7934 -3810 8014 -2834
rect 8014 -3810 8048 -2834
rect 8110 -3810 8144 -2834
rect 8144 -3810 8224 -2834
rect 8224 -3810 8258 -2834
rect 8320 -3810 8354 -2834
rect 8354 -3810 8434 -2834
rect 8434 -3810 8468 -2834
rect 8530 -3810 8564 -2834
rect 8564 -3810 8644 -2834
rect 8644 -3810 8678 -2834
rect 8740 -3810 8774 -2834
rect 8774 -3810 8854 -2834
rect 8854 -3810 8888 -2834
rect 8950 -3810 8984 -2834
rect 8984 -3810 9064 -2834
rect 9064 -3810 9098 -2834
rect 9160 -3810 9194 -2834
rect 9194 -3810 9218 -2834
rect 2950 -4272 3248 -3990
rect 5470 -6826 5494 -5850
rect 5494 -6826 5528 -5850
rect 5590 -6826 5624 -5850
rect 5624 -6826 5704 -5850
rect 5704 -6826 5738 -5850
rect 5800 -6826 5834 -5850
rect 5834 -6826 5914 -5850
rect 5914 -6826 5948 -5850
rect 6010 -6826 6044 -5850
rect 6044 -6826 6124 -5850
rect 6124 -6826 6158 -5850
rect 6220 -6826 6254 -5850
rect 6254 -6826 6334 -5850
rect 6334 -6826 6368 -5850
rect 6430 -6826 6464 -5850
rect 6464 -6826 6544 -5850
rect 6544 -6826 6578 -5850
rect 6640 -6826 6674 -5850
rect 6674 -6826 6754 -5850
rect 6754 -6826 6788 -5850
rect 6850 -6826 6884 -5850
rect 6884 -6826 6964 -5850
rect 6964 -6826 6998 -5850
rect 7060 -6826 7094 -5850
rect 7094 -6826 7174 -5850
rect 7174 -6826 7208 -5850
rect 7270 -6826 7304 -5850
rect 7304 -6826 7384 -5850
rect 7384 -6826 7418 -5850
rect 7480 -6826 7514 -5850
rect 7514 -6826 7594 -5850
rect 7594 -6826 7628 -5850
rect 7690 -6826 7724 -5850
rect 7724 -6826 7804 -5850
rect 7804 -6826 7838 -5850
rect 7900 -6826 7934 -5850
rect 7934 -6826 8014 -5850
rect 8014 -6826 8048 -5850
rect 8110 -6826 8144 -5850
rect 8144 -6826 8224 -5850
rect 8224 -6826 8258 -5850
rect 8320 -6826 8354 -5850
rect 8354 -6826 8434 -5850
rect 8434 -6826 8468 -5850
rect 8530 -6826 8564 -5850
rect 8564 -6826 8644 -5850
rect 8644 -6826 8678 -5850
rect 8740 -6826 8774 -5850
rect 8774 -6826 8854 -5850
rect 8854 -6826 8888 -5850
rect 8950 -6826 8984 -5850
rect 8984 -6826 9064 -5850
rect 9064 -6826 9098 -5850
rect 9160 -6826 9194 -5850
rect 9194 -6826 9218 -5850
rect 5490 -7104 5590 -7004
rect 5910 -7104 6010 -7004
rect 6330 -7104 6430 -7004
rect 6750 -7104 6850 -7004
rect 7170 -7104 7270 -7004
rect 7590 -7104 7690 -7004
rect 8010 -7104 8110 -7004
rect 8430 -7104 8530 -7004
rect 8850 -7104 8950 -7004
rect 9176 -7104 9276 -7004
<< metal2 >>
rect 10130 13618 10428 13628
rect 10130 13326 10302 13336
rect 10400 13326 10428 13336
rect 10580 13618 10878 13628
rect 10580 13326 10722 13336
rect 10302 13258 10400 13268
rect 10650 13268 10722 13326
rect 10820 13326 10878 13336
rect 11000 13618 11298 13628
rect 11000 13326 11142 13336
rect 10650 13258 10820 13268
rect 11070 13268 11142 13326
rect 11240 13326 11298 13336
rect 11420 13618 11718 13628
rect 11420 13326 11562 13336
rect 11070 13258 11240 13268
rect 11490 13268 11562 13326
rect 11660 13326 11718 13336
rect 11840 13618 12138 13628
rect 11840 13326 11982 13336
rect 11490 13258 11660 13268
rect 11910 13268 11982 13326
rect 12080 13326 12138 13336
rect 12260 13618 12558 13628
rect 12260 13326 12402 13336
rect 11910 13258 12080 13268
rect 12330 13268 12402 13326
rect 12500 13326 12558 13336
rect 12680 13618 12978 13628
rect 12680 13326 12822 13336
rect 12330 13258 12500 13268
rect 12750 13268 12822 13326
rect 12920 13326 12978 13336
rect 13100 13618 13398 13628
rect 13100 13326 13242 13336
rect 12750 13258 12920 13268
rect 13170 13268 13242 13326
rect 13340 13326 13398 13336
rect 13520 13618 13818 13628
rect 13520 13326 13662 13336
rect 13170 13258 13340 13268
rect 13590 13268 13662 13326
rect 13760 13326 13818 13336
rect 13940 13618 14238 13628
rect 13940 13326 14082 13336
rect 13590 13258 13760 13268
rect 14010 13268 14082 13326
rect 14180 13326 14238 13336
rect 14360 13618 14658 13628
rect 14360 13326 14502 13336
rect 14010 13258 14180 13268
rect 14430 13268 14502 13326
rect 14600 13326 14658 13336
rect 14780 13618 15078 13628
rect 14780 13326 14922 13336
rect 14430 13258 14600 13268
rect 14850 13268 14922 13326
rect 15020 13326 15078 13336
rect 15200 13618 15498 13628
rect 15200 13326 15342 13336
rect 14850 13258 15020 13268
rect 15270 13268 15342 13326
rect 15440 13326 15498 13336
rect 15620 13618 15918 13628
rect 15620 13326 15762 13336
rect 15270 13258 15440 13268
rect 15690 13268 15762 13326
rect 15860 13326 15918 13336
rect 16040 13618 16338 13628
rect 16040 13326 16182 13336
rect 15690 13258 15860 13268
rect 16110 13268 16182 13326
rect 16280 13326 16338 13336
rect 16460 13618 16758 13628
rect 16460 13326 16602 13336
rect 16110 13258 16280 13268
rect 16530 13268 16602 13326
rect 16700 13326 16758 13336
rect 16880 13618 17178 13628
rect 16880 13326 17022 13336
rect 16530 13258 16700 13268
rect 16950 13268 17022 13326
rect 17120 13326 17178 13336
rect 17300 13618 17598 13628
rect 17300 13326 17442 13336
rect 16950 13258 17120 13268
rect 17370 13268 17442 13326
rect 17540 13326 17598 13336
rect 17720 13618 18018 13628
rect 17720 13326 17862 13336
rect 17370 13258 17540 13268
rect 17790 13268 17862 13326
rect 17960 13326 18018 13336
rect 18140 13618 18438 13628
rect 18140 13326 18282 13336
rect 17790 13258 17960 13268
rect 18210 13268 18282 13326
rect 18380 13326 18438 13336
rect 18560 13618 18858 13628
rect 18560 13326 18630 13336
rect 18210 13258 18380 13268
rect 18728 13326 18858 13336
rect 18630 13258 18728 13268
rect 10320 13036 10378 13258
rect 10320 11818 10378 12060
rect 10320 10832 10378 10842
rect 10440 13036 10588 13046
rect 10440 11818 10588 12060
rect 10440 10704 10588 10842
rect 10650 13036 10798 13258
rect 10650 11818 10798 12060
rect 10650 10832 10798 10842
rect 10860 13036 11008 13046
rect 10860 11818 11008 12060
rect 10860 10704 11008 10842
rect 11070 13036 11218 13258
rect 11070 11818 11218 12060
rect 11070 10832 11218 10842
rect 11280 13036 11428 13046
rect 11280 11818 11428 12060
rect 11280 10704 11428 10842
rect 11490 13036 11638 13258
rect 11490 11818 11638 12060
rect 11490 10832 11638 10842
rect 11700 13036 11848 13046
rect 11700 11818 11848 12060
rect 11700 10704 11848 10842
rect 11910 13036 12058 13258
rect 11910 11818 12058 12060
rect 11910 10832 12058 10842
rect 12120 13036 12268 13046
rect 12120 11818 12268 12060
rect 12120 10704 12268 10842
rect 12330 13036 12478 13258
rect 12330 11818 12478 12060
rect 12330 10832 12478 10842
rect 12540 13036 12688 13046
rect 12540 11818 12688 12060
rect 12540 10704 12688 10842
rect 12750 13036 12898 13258
rect 12750 11818 12898 12060
rect 12750 10832 12898 10842
rect 12960 13036 13108 13046
rect 12960 11818 13108 12060
rect 12960 10704 13108 10842
rect 13170 13036 13318 13258
rect 13170 11818 13318 12060
rect 13170 10832 13318 10842
rect 13380 13036 13528 13046
rect 13380 11818 13528 12060
rect 13380 10704 13528 10842
rect 13590 13036 13738 13258
rect 13590 11818 13738 12060
rect 13590 10832 13738 10842
rect 13800 13036 13948 13046
rect 13800 11818 13948 12060
rect 13800 10704 13948 10842
rect 14010 13036 14158 13258
rect 14010 11818 14158 12060
rect 14010 10832 14158 10842
rect 14220 13036 14368 13046
rect 14220 11818 14368 12060
rect 14220 10704 14368 10842
rect 14430 13036 14578 13258
rect 14430 11818 14578 12060
rect 14430 10832 14578 10842
rect 14640 13036 14788 13046
rect 14640 11818 14788 12060
rect 14640 10704 14788 10842
rect 14850 13036 14998 13258
rect 14850 11818 14998 12060
rect 14850 10832 14998 10842
rect 15060 13036 15208 13046
rect 15060 11818 15208 12060
rect 15060 10704 15208 10842
rect 15270 13036 15418 13258
rect 15270 11818 15418 12060
rect 15270 10832 15418 10842
rect 15480 13036 15628 13046
rect 15480 11818 15628 12060
rect 15480 10704 15628 10842
rect 15690 13036 15838 13258
rect 15690 11818 15838 12060
rect 15690 10832 15838 10842
rect 15900 13036 16048 13046
rect 15900 11818 16048 12060
rect 15900 10704 16048 10842
rect 16110 13036 16258 13258
rect 16110 11818 16258 12060
rect 16110 10832 16258 10842
rect 16320 13036 16468 13046
rect 16320 11818 16468 12060
rect 16320 10704 16468 10842
rect 16530 13036 16678 13258
rect 16530 11818 16678 12060
rect 16530 10832 16678 10842
rect 16740 13036 16888 13046
rect 16740 11818 16888 12060
rect 16740 10704 16888 10842
rect 16950 13036 17098 13258
rect 16950 11818 17098 12060
rect 16950 10832 17098 10842
rect 17160 13036 17308 13046
rect 17160 11818 17308 12060
rect 17160 10704 17308 10842
rect 17370 13036 17518 13258
rect 17370 11818 17518 12060
rect 17370 10832 17518 10842
rect 17580 13036 17728 13046
rect 17580 11818 17728 12060
rect 17580 10704 17728 10842
rect 17790 13036 17938 13258
rect 17790 11818 17938 12060
rect 17790 10832 17938 10842
rect 18000 13036 18148 13046
rect 18000 11818 18148 12060
rect 18000 10704 18148 10842
rect 18210 13036 18358 13258
rect 18210 11818 18358 12060
rect 18210 10832 18358 10842
rect 18420 13036 18568 13046
rect 18420 11818 18568 12060
rect 18420 10704 18568 10842
rect 18630 13036 18688 13258
rect 18630 11818 18688 12060
rect 18630 10832 18688 10842
rect 10440 8006 18568 10704
rect 10320 7808 10378 7818
rect 5292 7440 5590 7450
rect 5292 7148 5490 7158
rect 5470 7130 5490 7148
rect 5712 7440 6010 7450
rect 5712 7148 5910 7158
rect 5470 7120 5590 7130
rect 5800 7130 5910 7148
rect 6132 7440 6430 7450
rect 6132 7148 6330 7158
rect 5800 7124 6010 7130
rect 6220 7130 6330 7148
rect 6552 7440 6850 7450
rect 6552 7148 6750 7158
rect 6220 7124 6430 7130
rect 6640 7130 6750 7148
rect 6972 7440 7270 7450
rect 6972 7148 7170 7158
rect 6640 7124 6850 7130
rect 7060 7130 7170 7148
rect 7392 7440 7690 7450
rect 7392 7148 7590 7158
rect 7060 7124 7270 7130
rect 7480 7130 7590 7148
rect 7812 7440 8110 7450
rect 7812 7148 8010 7158
rect 7480 7124 7690 7130
rect 7900 7130 8010 7148
rect 8232 7440 8530 7450
rect 8232 7148 8430 7158
rect 7900 7124 8110 7130
rect 8320 7130 8430 7148
rect 8652 7440 8950 7450
rect 8652 7148 8850 7158
rect 8320 7124 8530 7130
rect 8740 7130 8850 7148
rect 9072 7440 9370 7450
rect 9072 7148 9176 7158
rect 8740 7124 8950 7130
rect 9160 7130 9176 7148
rect 9276 7148 9370 7158
rect 5470 6952 5528 7120
rect 5470 5966 5528 5976
rect 5590 6952 5738 6962
rect 5590 5850 5738 5976
rect 5800 6952 5948 7124
rect 5800 5966 5948 5976
rect 6010 6952 6158 6962
rect 6010 5850 6158 5976
rect 6220 6952 6368 7124
rect 6220 5966 6368 5976
rect 6430 6952 6578 6962
rect 6430 5850 6578 5976
rect 6640 6952 6788 7124
rect 6640 5966 6788 5976
rect 6850 6952 6998 6962
rect 6850 5850 6998 5976
rect 7060 6952 7208 7124
rect 7060 5966 7208 5976
rect 7270 6952 7418 6962
rect 7270 5850 7418 5976
rect 7480 6952 7628 7124
rect 7480 5966 7628 5976
rect 7690 6952 7838 6962
rect 7690 5850 7838 5976
rect 7900 6952 8048 7124
rect 7900 5966 8048 5976
rect 8110 6952 8258 6962
rect 8110 5850 8258 5976
rect 8320 6952 8468 7124
rect 8320 5966 8468 5976
rect 8530 6952 8678 6962
rect 8530 5850 8678 5976
rect 8740 6952 8888 7124
rect 9160 7120 9276 7130
rect 8740 5966 8888 5976
rect 8950 6952 9098 6962
rect 8950 5850 9098 5976
rect 9160 6952 9218 7120
rect 10320 6572 10378 6832
rect 9160 5966 9218 5976
rect 9326 5996 9936 6006
rect 2490 5798 2788 5808
rect 2490 5506 2788 5516
rect 2950 5798 3248 5808
rect 2950 5506 3248 5516
rect 3350 5798 3648 5808
rect 3350 5506 3648 5516
rect 3770 5798 4068 5808
rect 3770 5506 4068 5516
rect 4190 5798 4488 5808
rect 4190 5506 4488 5516
rect 2566 5328 2620 5506
rect 2566 4342 2620 4352
rect 2668 5328 2728 5338
rect 2668 4352 2674 5328
rect 3510 5328 3564 5506
rect 2668 4342 2728 4352
rect 2794 4404 2936 4414
rect 2668 4272 2794 4342
rect 2544 4100 2616 4110
rect 2544 3012 2616 3124
rect 2668 4100 2722 4272
rect 3510 4342 3564 4352
rect 3626 5328 3774 5338
rect 3626 4288 3774 4352
rect 3836 5328 3984 5506
rect 3836 4342 3984 4352
rect 4046 5328 4194 5338
rect 4046 4288 4194 4352
rect 4256 5328 4310 5506
rect 4350 5504 4404 5506
rect 5590 5470 9326 5850
rect 5470 5336 5528 5346
rect 4726 4764 5008 4774
rect 4726 4490 5008 4500
rect 4256 4342 4310 4352
rect 4790 4288 4944 4490
rect 2794 4246 2936 4256
rect 3296 4168 4944 4288
rect 2668 3114 2722 3124
rect 2774 4100 2846 4110
rect 2774 3012 2846 3124
rect 3296 4100 3354 4168
rect 3296 3114 3354 3124
rect 3416 4100 3564 4110
rect 2492 3002 2886 3012
rect 3416 2970 3564 3124
rect 3626 4100 3774 4168
rect 3626 3114 3774 3124
rect 3836 4100 3984 4110
rect 3836 2970 3984 3124
rect 4046 4100 4194 4168
rect 4046 3114 4194 3124
rect 4256 4100 4404 4110
rect 4256 2970 4404 3124
rect 4466 4100 4614 4168
rect 4466 3114 4614 3124
rect 4676 4100 4824 4110
rect 4676 2970 4824 3124
rect 4886 4100 4944 4168
rect 4886 3114 4944 3124
rect 5470 4100 5528 4360
rect 5470 2980 5528 3124
rect 5590 5336 5738 5470
rect 5590 4100 5738 4360
rect 5590 3114 5738 3124
rect 5800 5336 5948 5346
rect 5800 4100 5948 4360
rect 5800 2980 5948 3124
rect 6010 5336 6158 5470
rect 6010 4100 6158 4360
rect 6010 3114 6158 3124
rect 6220 5336 6368 5346
rect 6220 4100 6368 4360
rect 5366 2970 5528 2980
rect 5786 2970 5948 2980
rect 6220 2976 6368 3124
rect 6430 5336 6578 5470
rect 6430 4100 6578 4360
rect 6430 3114 6578 3124
rect 6640 5336 6788 5346
rect 6640 4100 6788 4360
rect 6640 2976 6788 3124
rect 6850 5336 6998 5470
rect 6850 4100 6998 4360
rect 6850 3114 6998 3124
rect 7060 5336 7208 5346
rect 7060 4100 7208 4360
rect 7060 2976 7208 3124
rect 7270 5336 7418 5470
rect 7270 4100 7418 4360
rect 7270 3114 7418 3124
rect 7480 5336 7628 5346
rect 7480 4100 7628 4360
rect 7480 2976 7628 3124
rect 7690 5336 7838 5470
rect 7690 4100 7838 4360
rect 7690 3114 7838 3124
rect 7900 5336 8048 5346
rect 7900 4100 8048 4360
rect 7900 2976 8048 3124
rect 8110 5336 8258 5470
rect 8110 4100 8258 4360
rect 8110 3114 8258 3124
rect 8320 5336 8468 5346
rect 8320 4100 8468 4360
rect 8320 2976 8468 3124
rect 8530 5336 8678 5470
rect 8530 4100 8678 4360
rect 8530 3114 8678 3124
rect 8740 5336 8888 5346
rect 8740 4100 8888 4360
rect 8740 2976 8888 3124
rect 8950 5336 9098 5470
rect 9326 5368 9936 5378
rect 8950 4100 9098 4360
rect 8950 3114 9098 3124
rect 9160 5336 9218 5346
rect 9160 4100 9218 4360
rect 9160 2976 9218 3124
rect 10320 5336 10378 5596
rect 10320 4100 10378 4360
rect 6206 2970 6368 2976
rect 6626 2970 6788 2976
rect 7046 2970 7208 2976
rect 7466 2970 7628 2976
rect 7886 2970 8048 2976
rect 8306 2970 8468 2976
rect 8726 2970 8888 2976
rect 9146 2970 9258 2976
rect 10320 2970 10378 3124
rect 10440 7808 10588 8006
rect 10440 6572 10588 6832
rect 10440 5336 10588 5596
rect 10440 4100 10588 4360
rect 10440 3114 10588 3124
rect 10650 7808 10798 7818
rect 10650 6572 10798 6832
rect 10650 5336 10798 5596
rect 10650 4100 10798 4360
rect 10650 2970 10798 3124
rect 10860 7808 11008 8006
rect 10860 6572 11008 6832
rect 10860 5336 11008 5596
rect 10860 4100 11008 4360
rect 10860 3114 11008 3124
rect 11070 7808 11218 7818
rect 11070 6572 11218 6832
rect 11070 5336 11218 5596
rect 11070 4100 11218 4360
rect 11070 2970 11218 3124
rect 11280 7808 11428 8006
rect 11280 6572 11428 6832
rect 11280 5336 11428 5596
rect 11280 4100 11428 4360
rect 11280 3114 11428 3124
rect 11490 7808 11638 7818
rect 11490 6572 11638 6832
rect 11490 5336 11638 5596
rect 11490 4100 11638 4360
rect 11490 2970 11638 3124
rect 11700 7808 11848 8006
rect 11700 6572 11848 6832
rect 11700 5336 11848 5596
rect 11700 4100 11848 4360
rect 11700 3114 11848 3124
rect 11910 7808 12058 7818
rect 11910 6572 12058 6832
rect 11910 5336 12058 5596
rect 11910 4100 12058 4360
rect 11910 2970 12058 3124
rect 12120 7808 12268 8006
rect 12120 6572 12268 6832
rect 12120 5336 12268 5596
rect 12120 4100 12268 4360
rect 12120 3114 12268 3124
rect 12330 7808 12478 7818
rect 12330 6572 12478 6832
rect 12330 5336 12478 5596
rect 12330 4100 12478 4360
rect 12330 2970 12478 3124
rect 12540 7808 12688 8006
rect 12540 6572 12688 6832
rect 12540 5336 12688 5596
rect 12540 4100 12688 4360
rect 12540 3114 12688 3124
rect 12750 7808 12898 7818
rect 12750 6572 12898 6832
rect 12750 5336 12898 5596
rect 12750 4100 12898 4360
rect 12750 2970 12898 3124
rect 12960 7808 13108 8006
rect 12960 6572 13108 6832
rect 12960 5336 13108 5596
rect 12960 4100 13108 4360
rect 12960 3114 13108 3124
rect 13170 7808 13318 7818
rect 13170 6572 13318 6832
rect 13170 5336 13318 5596
rect 13170 4100 13318 4360
rect 13170 2970 13318 3124
rect 13380 7808 13528 8006
rect 13380 6572 13528 6832
rect 13380 5336 13528 5596
rect 13380 4100 13528 4360
rect 13380 3114 13528 3124
rect 13590 7808 13738 7818
rect 13590 6572 13738 6832
rect 13590 5336 13738 5596
rect 13590 4100 13738 4360
rect 13590 2970 13738 3124
rect 13800 7808 13948 8006
rect 13800 6572 13948 6832
rect 13800 5336 13948 5596
rect 13800 4100 13948 4360
rect 13800 3114 13948 3124
rect 14010 7808 14158 7818
rect 14010 6572 14158 6832
rect 14010 5336 14158 5596
rect 14010 4100 14158 4360
rect 14010 2970 14158 3124
rect 14220 7808 14368 8006
rect 14220 6572 14368 6832
rect 14220 5336 14368 5596
rect 14220 4100 14368 4360
rect 14220 3114 14368 3124
rect 14430 7808 14578 7818
rect 14430 6572 14578 6832
rect 14430 5336 14578 5596
rect 14430 4100 14578 4360
rect 14430 2970 14578 3124
rect 14640 7808 14788 8006
rect 14640 6572 14788 6832
rect 14640 5336 14788 5596
rect 14640 4100 14788 4360
rect 14640 3114 14788 3124
rect 14850 7808 14998 7818
rect 14850 6572 14998 6832
rect 14850 5336 14998 5596
rect 14850 4100 14998 4360
rect 14850 2970 14998 3124
rect 15060 7808 15208 8006
rect 15060 6572 15208 6832
rect 15060 5336 15208 5596
rect 15060 4100 15208 4360
rect 15060 3114 15208 3124
rect 15270 7808 15418 7818
rect 15270 6572 15418 6832
rect 15270 5336 15418 5596
rect 15270 4100 15418 4360
rect 15270 2970 15418 3124
rect 15480 7808 15628 8006
rect 15480 6572 15628 6832
rect 15480 5336 15628 5596
rect 15480 4100 15628 4360
rect 15480 3114 15628 3124
rect 15690 7808 15838 7818
rect 15690 6572 15838 6832
rect 15690 5336 15838 5596
rect 15690 4100 15838 4360
rect 15690 2970 15838 3124
rect 15900 7808 16048 8006
rect 15900 6572 16048 6832
rect 15900 5336 16048 5596
rect 15900 4100 16048 4360
rect 15900 3114 16048 3124
rect 16110 7808 16258 7818
rect 16110 6572 16258 6832
rect 16110 5336 16258 5596
rect 16110 4100 16258 4360
rect 16110 2970 16258 3124
rect 16320 7808 16468 8006
rect 16320 6572 16468 6832
rect 16320 5336 16468 5596
rect 16320 4100 16468 4360
rect 16320 3114 16468 3124
rect 16530 7808 16678 7818
rect 16530 6572 16678 6832
rect 16530 5336 16678 5596
rect 16530 4100 16678 4360
rect 16530 2970 16678 3124
rect 16740 7808 16888 8006
rect 16740 6572 16888 6832
rect 16740 5336 16888 5596
rect 16740 4100 16888 4360
rect 16740 3114 16888 3124
rect 16950 7808 17098 7818
rect 16950 6572 17098 6832
rect 16950 5336 17098 5596
rect 16950 4100 17098 4360
rect 16950 2970 17098 3124
rect 17160 7808 17308 8006
rect 17160 6572 17308 6832
rect 17160 5336 17308 5596
rect 17160 4100 17308 4360
rect 17160 3114 17308 3124
rect 17370 7808 17518 7818
rect 17370 6572 17518 6832
rect 17370 5336 17518 5596
rect 17370 4100 17518 4360
rect 17370 2970 17518 3124
rect 17580 7808 17728 8006
rect 17580 6572 17728 6832
rect 17580 5336 17728 5596
rect 17580 4100 17728 4360
rect 17580 3114 17728 3124
rect 17790 7808 17938 7818
rect 17790 6572 17938 6832
rect 17790 5336 17938 5596
rect 17790 4100 17938 4360
rect 17790 2970 17938 3124
rect 18000 7808 18148 8006
rect 18000 6572 18148 6832
rect 18000 5336 18148 5596
rect 18000 4100 18148 4360
rect 18000 3114 18148 3124
rect 18210 7808 18358 7818
rect 18210 6572 18358 6832
rect 18210 5336 18358 5596
rect 18210 4100 18358 4360
rect 18210 2970 18358 3124
rect 18420 7808 18568 8006
rect 18420 6572 18568 6832
rect 18420 5336 18568 5596
rect 18420 4100 18568 4360
rect 18420 3114 18568 3124
rect 18630 7808 18688 7818
rect 18630 6572 18688 6832
rect 18630 5336 18688 5596
rect 18630 4100 18688 4360
rect 18630 2970 18688 3124
rect 3338 2960 3636 2970
rect 2492 2828 2886 2838
rect 2984 2838 3128 2848
rect 2984 2680 3128 2690
rect 3338 2668 3636 2678
rect 3758 2960 4056 2970
rect 3758 2668 4056 2678
rect 4178 2960 4476 2970
rect 4178 2668 4476 2678
rect 4598 2960 4896 2970
rect 4598 2668 4896 2678
rect 5298 2960 5366 2970
rect 5466 2960 5596 2970
rect 5298 2668 5596 2678
rect 5728 2960 5786 2970
rect 5886 2960 6026 2970
rect 5728 2668 6026 2678
rect 6148 2960 6206 2970
rect 6306 2960 6446 2970
rect 6148 2668 6446 2678
rect 6568 2960 6626 2970
rect 6726 2960 6866 2970
rect 6568 2668 6866 2678
rect 6988 2960 7046 2970
rect 7146 2960 7286 2970
rect 6988 2668 7286 2678
rect 7408 2960 7466 2970
rect 7566 2960 7706 2970
rect 7408 2668 7706 2678
rect 7828 2960 7886 2970
rect 7986 2960 8126 2970
rect 7828 2668 8126 2678
rect 8248 2960 8306 2970
rect 8406 2960 8546 2970
rect 8248 2668 8546 2678
rect 8668 2960 8726 2970
rect 8826 2960 8966 2970
rect 8668 2668 8966 2678
rect 9088 2960 9146 2970
rect 9246 2960 9386 2970
rect 9088 2668 9386 2678
rect 10128 2960 10426 2970
rect 10128 2668 10426 2678
rect 10578 2960 10876 2970
rect 10578 2668 10876 2678
rect 10998 2960 11296 2970
rect 10998 2668 11296 2678
rect 11418 2960 11716 2970
rect 11418 2668 11716 2678
rect 11838 2960 12136 2970
rect 11838 2668 12136 2678
rect 12258 2960 12556 2970
rect 12258 2668 12556 2678
rect 12678 2960 12976 2970
rect 12678 2668 12976 2678
rect 13098 2960 13396 2970
rect 13098 2668 13396 2678
rect 13518 2960 13816 2970
rect 13518 2668 13816 2678
rect 13938 2960 14236 2970
rect 13938 2668 14236 2678
rect 14358 2960 14656 2970
rect 14358 2668 14656 2678
rect 14778 2960 15076 2970
rect 14778 2668 15076 2678
rect 15198 2960 15496 2970
rect 15198 2668 15496 2678
rect 15618 2960 15916 2970
rect 15618 2668 15916 2678
rect 16038 2960 16336 2970
rect 16038 2668 16336 2678
rect 16458 2960 16756 2970
rect 16458 2668 16756 2678
rect 16878 2960 17176 2970
rect 16878 2668 17176 2678
rect 17298 2960 17596 2970
rect 17298 2668 17596 2678
rect 17718 2960 18016 2970
rect 17718 2668 18016 2678
rect 18138 2960 18436 2970
rect 18138 2668 18436 2678
rect 18558 2960 18856 2970
rect 18558 2668 18856 2678
rect 196 2482 524 2492
rect 196 2210 524 2220
rect 4386 1534 4630 1544
rect -188 1458 4386 1468
rect -114 1400 4386 1458
rect -188 1390 4386 1400
rect 4386 1276 4630 1286
rect 5020 222 5264 232
rect -26 40 5020 52
rect 36 -14 5020 40
rect -26 -26 5020 -14
rect 5020 -36 5264 -26
rect 196 -694 524 -684
rect 196 -966 524 -956
rect 3338 -1152 3636 -1142
rect 2984 -1164 3128 -1154
rect 2492 -1312 2886 -1302
rect 2984 -1322 3128 -1312
rect 3338 -1444 3636 -1434
rect 3758 -1152 4056 -1142
rect 3758 -1444 4056 -1434
rect 4178 -1152 4476 -1142
rect 4178 -1444 4476 -1434
rect 4598 -1152 4896 -1142
rect 4598 -1444 4896 -1434
rect 5298 -1152 5596 -1142
rect 5298 -1444 5366 -1434
rect 5466 -1444 5596 -1434
rect 5728 -1152 6026 -1142
rect 5728 -1444 5786 -1434
rect 5886 -1444 6026 -1434
rect 6148 -1152 6446 -1142
rect 6148 -1444 6206 -1434
rect 6306 -1444 6446 -1434
rect 6568 -1152 6866 -1142
rect 6568 -1444 6626 -1434
rect 6726 -1444 6866 -1434
rect 6988 -1152 7286 -1142
rect 6988 -1444 7046 -1434
rect 7146 -1444 7286 -1434
rect 7408 -1152 7706 -1142
rect 7408 -1444 7466 -1434
rect 7566 -1444 7706 -1434
rect 7828 -1152 8126 -1142
rect 7828 -1444 7886 -1434
rect 7986 -1444 8126 -1434
rect 8248 -1152 8546 -1142
rect 8248 -1444 8306 -1434
rect 8406 -1444 8546 -1434
rect 8668 -1152 8966 -1142
rect 8668 -1444 8726 -1434
rect 8826 -1444 8966 -1434
rect 9088 -1152 9386 -1142
rect 9088 -1444 9146 -1434
rect 9246 -1444 9386 -1434
rect 2492 -1486 2886 -1476
rect 2544 -1598 2616 -1486
rect 2544 -2584 2616 -2574
rect 2668 -1598 2722 -1588
rect 2668 -2746 2722 -2574
rect 2774 -1598 2846 -1486
rect 2774 -2584 2846 -2574
rect 3296 -1598 3354 -1588
rect 3296 -2642 3354 -2574
rect 3416 -1598 3564 -1444
rect 3416 -2584 3564 -2574
rect 3626 -1598 3774 -1588
rect 3626 -2642 3774 -2574
rect 3836 -1598 3984 -1444
rect 3836 -2584 3984 -2574
rect 4046 -1598 4194 -1588
rect 4046 -2642 4194 -2574
rect 4256 -1598 4404 -1444
rect 4256 -2584 4404 -2574
rect 4466 -1598 4614 -1588
rect 4466 -2642 4614 -2574
rect 4676 -1598 4824 -1444
rect 5366 -1454 5528 -1444
rect 5786 -1454 5948 -1444
rect 6206 -1450 6368 -1444
rect 6626 -1450 6788 -1444
rect 7046 -1450 7208 -1444
rect 7466 -1450 7628 -1444
rect 7886 -1450 8048 -1444
rect 8306 -1450 8468 -1444
rect 8726 -1450 8888 -1444
rect 9146 -1450 9258 -1444
rect 4676 -2584 4824 -2574
rect 4886 -1598 4944 -1588
rect 4886 -2642 4944 -2574
rect 2794 -2730 2936 -2720
rect 2668 -2816 2794 -2746
rect 2566 -2826 2620 -2816
rect 2566 -3980 2620 -3802
rect 2668 -2826 2728 -2816
rect 2668 -3802 2674 -2826
rect 3296 -2762 4944 -2642
rect 2794 -2888 2936 -2878
rect 3510 -2826 3564 -2816
rect 2668 -3812 2728 -3802
rect 3510 -3980 3564 -3802
rect 3626 -2826 3774 -2762
rect 3626 -3812 3774 -3802
rect 3836 -2826 3984 -2816
rect 3836 -3980 3984 -3802
rect 4046 -2826 4194 -2762
rect 4046 -3812 4194 -3802
rect 4256 -2826 4310 -2816
rect 4790 -2964 4944 -2762
rect 5470 -1598 5528 -1454
rect 5470 -2834 5528 -2574
rect 4726 -2974 5008 -2964
rect 4726 -3248 5008 -3238
rect 4256 -3980 4310 -3802
rect 5470 -3820 5528 -3810
rect 5590 -1598 5738 -1588
rect 5590 -2834 5738 -2574
rect 5590 -3944 5738 -3810
rect 5800 -1598 5948 -1454
rect 5800 -2834 5948 -2574
rect 5800 -3820 5948 -3810
rect 6010 -1598 6158 -1588
rect 6010 -2834 6158 -2574
rect 6010 -3944 6158 -3810
rect 6220 -1598 6368 -1450
rect 6220 -2834 6368 -2574
rect 6220 -3820 6368 -3810
rect 6430 -1598 6578 -1588
rect 6430 -2834 6578 -2574
rect 6430 -3944 6578 -3810
rect 6640 -1598 6788 -1450
rect 6640 -2834 6788 -2574
rect 6640 -3820 6788 -3810
rect 6850 -1598 6998 -1588
rect 6850 -2834 6998 -2574
rect 6850 -3944 6998 -3810
rect 7060 -1598 7208 -1450
rect 7060 -2834 7208 -2574
rect 7060 -3820 7208 -3810
rect 7270 -1598 7418 -1588
rect 7270 -2834 7418 -2574
rect 7270 -3944 7418 -3810
rect 7480 -1598 7628 -1450
rect 7480 -2834 7628 -2574
rect 7480 -3820 7628 -3810
rect 7690 -1598 7838 -1588
rect 7690 -2834 7838 -2574
rect 7690 -3944 7838 -3810
rect 7900 -1598 8048 -1450
rect 7900 -2834 8048 -2574
rect 7900 -3820 8048 -3810
rect 8110 -1598 8258 -1588
rect 8110 -2834 8258 -2574
rect 8110 -3944 8258 -3810
rect 8320 -1598 8468 -1450
rect 8320 -2834 8468 -2574
rect 8320 -3820 8468 -3810
rect 8530 -1598 8678 -1588
rect 8530 -2834 8678 -2574
rect 8530 -3944 8678 -3810
rect 8740 -1598 8888 -1450
rect 8740 -2834 8888 -2574
rect 8740 -3820 8888 -3810
rect 8950 -1598 9098 -1588
rect 8950 -2834 9098 -2574
rect 8950 -3944 9098 -3810
rect 9160 -1598 9218 -1450
rect 9160 -2834 9218 -2574
rect 9160 -3820 9218 -3810
rect 4350 -3980 4404 -3978
rect 2490 -3990 2788 -3980
rect 2490 -4282 2788 -4272
rect 2950 -3990 3248 -3980
rect 2950 -4282 3248 -4272
rect 3350 -3990 3648 -3980
rect 3350 -4282 3648 -4272
rect 3770 -3990 4068 -3980
rect 3770 -4282 4068 -4272
rect 4190 -3990 4488 -3980
rect 4190 -4282 4488 -4272
rect 5590 -5724 9314 -3944
rect 5470 -5850 5528 -5840
rect 5470 -6994 5528 -6826
rect 5590 -5850 5738 -5724
rect 5590 -6836 5738 -6826
rect 5800 -5850 5948 -5840
rect 5470 -7004 5590 -6994
rect 5470 -7022 5490 -7004
rect 5292 -7032 5490 -7022
rect 5800 -6998 5948 -6826
rect 6010 -5850 6158 -5724
rect 6010 -6836 6158 -6826
rect 6220 -5850 6368 -5840
rect 6220 -6998 6368 -6826
rect 6430 -5850 6578 -5724
rect 6430 -6836 6578 -6826
rect 6640 -5850 6788 -5840
rect 6640 -6998 6788 -6826
rect 6850 -5850 6998 -5724
rect 6850 -6836 6998 -6826
rect 7060 -5850 7208 -5840
rect 7060 -6998 7208 -6826
rect 7270 -5850 7418 -5724
rect 7270 -6836 7418 -6826
rect 7480 -5850 7628 -5840
rect 7480 -6998 7628 -6826
rect 7690 -5850 7838 -5724
rect 7690 -6836 7838 -6826
rect 7900 -5850 8048 -5840
rect 7900 -6998 8048 -6826
rect 8110 -5850 8258 -5724
rect 8110 -6836 8258 -6826
rect 8320 -5850 8468 -5840
rect 8320 -6998 8468 -6826
rect 8530 -5850 8678 -5724
rect 8530 -6836 8678 -6826
rect 8740 -5850 8888 -5840
rect 8740 -6998 8888 -6826
rect 8950 -5850 9098 -5724
rect 8950 -6836 9098 -6826
rect 9160 -5850 9218 -5840
rect 9160 -6994 9218 -6826
rect 5800 -7004 6010 -6998
rect 5800 -7022 5910 -7004
rect 5292 -7324 5590 -7314
rect 5712 -7032 5910 -7022
rect 6220 -7004 6430 -6998
rect 6220 -7022 6330 -7004
rect 5712 -7324 6010 -7314
rect 6132 -7032 6330 -7022
rect 6640 -7004 6850 -6998
rect 6640 -7022 6750 -7004
rect 6132 -7324 6430 -7314
rect 6552 -7032 6750 -7022
rect 7060 -7004 7270 -6998
rect 7060 -7022 7170 -7004
rect 6552 -7324 6850 -7314
rect 6972 -7032 7170 -7022
rect 7480 -7004 7690 -6998
rect 7480 -7022 7590 -7004
rect 6972 -7324 7270 -7314
rect 7392 -7032 7590 -7022
rect 7900 -7004 8110 -6998
rect 7900 -7022 8010 -7004
rect 7392 -7324 7690 -7314
rect 7812 -7032 8010 -7022
rect 8320 -7004 8530 -6998
rect 8320 -7022 8430 -7004
rect 7812 -7324 8110 -7314
rect 8232 -7032 8430 -7022
rect 8740 -7004 8950 -6998
rect 8740 -7022 8850 -7004
rect 8232 -7324 8530 -7314
rect 8652 -7032 8850 -7022
rect 9160 -7004 9276 -6994
rect 9160 -7022 9176 -7004
rect 8652 -7324 8950 -7314
rect 9072 -7032 9176 -7022
rect 9276 -7032 9370 -7022
rect 9072 -7324 9370 -7314
<< via2 >>
rect 10130 13372 10428 13618
rect 10130 13336 10302 13372
rect 10302 13336 10400 13372
rect 10400 13336 10428 13372
rect 10580 13372 10878 13618
rect 10580 13336 10722 13372
rect 10722 13336 10820 13372
rect 10820 13336 10878 13372
rect 11000 13372 11298 13618
rect 11000 13336 11142 13372
rect 11142 13336 11240 13372
rect 11240 13336 11298 13372
rect 11420 13372 11718 13618
rect 11420 13336 11562 13372
rect 11562 13336 11660 13372
rect 11660 13336 11718 13372
rect 11840 13372 12138 13618
rect 11840 13336 11982 13372
rect 11982 13336 12080 13372
rect 12080 13336 12138 13372
rect 12260 13372 12558 13618
rect 12260 13336 12402 13372
rect 12402 13336 12500 13372
rect 12500 13336 12558 13372
rect 12680 13372 12978 13618
rect 12680 13336 12822 13372
rect 12822 13336 12920 13372
rect 12920 13336 12978 13372
rect 13100 13372 13398 13618
rect 13100 13336 13242 13372
rect 13242 13336 13340 13372
rect 13340 13336 13398 13372
rect 13520 13372 13818 13618
rect 13520 13336 13662 13372
rect 13662 13336 13760 13372
rect 13760 13336 13818 13372
rect 13940 13372 14238 13618
rect 13940 13336 14082 13372
rect 14082 13336 14180 13372
rect 14180 13336 14238 13372
rect 14360 13372 14658 13618
rect 14360 13336 14502 13372
rect 14502 13336 14600 13372
rect 14600 13336 14658 13372
rect 14780 13372 15078 13618
rect 14780 13336 14922 13372
rect 14922 13336 15020 13372
rect 15020 13336 15078 13372
rect 15200 13372 15498 13618
rect 15200 13336 15342 13372
rect 15342 13336 15440 13372
rect 15440 13336 15498 13372
rect 15620 13372 15918 13618
rect 15620 13336 15762 13372
rect 15762 13336 15860 13372
rect 15860 13336 15918 13372
rect 16040 13372 16338 13618
rect 16040 13336 16182 13372
rect 16182 13336 16280 13372
rect 16280 13336 16338 13372
rect 16460 13372 16758 13618
rect 16460 13336 16602 13372
rect 16602 13336 16700 13372
rect 16700 13336 16758 13372
rect 16880 13372 17178 13618
rect 16880 13336 17022 13372
rect 17022 13336 17120 13372
rect 17120 13336 17178 13372
rect 17300 13372 17598 13618
rect 17300 13336 17442 13372
rect 17442 13336 17540 13372
rect 17540 13336 17598 13372
rect 17720 13372 18018 13618
rect 17720 13336 17862 13372
rect 17862 13336 17960 13372
rect 17960 13336 18018 13372
rect 18140 13372 18438 13618
rect 18140 13336 18282 13372
rect 18282 13336 18380 13372
rect 18380 13336 18438 13372
rect 18560 13372 18858 13618
rect 18560 13336 18630 13372
rect 18630 13336 18728 13372
rect 18728 13336 18858 13372
rect 5292 7230 5590 7440
rect 5292 7158 5490 7230
rect 5490 7158 5590 7230
rect 5712 7230 6010 7440
rect 5712 7158 5910 7230
rect 5910 7158 6010 7230
rect 6132 7230 6430 7440
rect 6132 7158 6330 7230
rect 6330 7158 6430 7230
rect 6552 7230 6850 7440
rect 6552 7158 6750 7230
rect 6750 7158 6850 7230
rect 6972 7230 7270 7440
rect 6972 7158 7170 7230
rect 7170 7158 7270 7230
rect 7392 7230 7690 7440
rect 7392 7158 7590 7230
rect 7590 7158 7690 7230
rect 7812 7230 8110 7440
rect 7812 7158 8010 7230
rect 8010 7158 8110 7230
rect 8232 7230 8530 7440
rect 8232 7158 8430 7230
rect 8430 7158 8530 7230
rect 8652 7230 8950 7440
rect 8652 7158 8850 7230
rect 8850 7158 8950 7230
rect 9072 7230 9370 7440
rect 9072 7158 9176 7230
rect 9176 7158 9276 7230
rect 9276 7158 9370 7230
rect 2490 5516 2788 5798
rect 2950 5516 3248 5798
rect 3350 5516 3648 5798
rect 3770 5516 4068 5798
rect 4190 5516 4488 5798
rect 2492 2838 2886 3002
rect 2984 2690 3128 2838
rect 3338 2678 3636 2960
rect 3758 2678 4056 2960
rect 4178 2678 4476 2960
rect 4598 2678 4896 2960
rect 5298 2870 5366 2960
rect 5366 2870 5466 2960
rect 5466 2870 5596 2960
rect 5298 2678 5596 2870
rect 5728 2870 5786 2960
rect 5786 2870 5886 2960
rect 5886 2870 6026 2960
rect 5728 2678 6026 2870
rect 6148 2870 6206 2960
rect 6206 2870 6306 2960
rect 6306 2870 6446 2960
rect 6148 2678 6446 2870
rect 6568 2870 6626 2960
rect 6626 2870 6726 2960
rect 6726 2870 6866 2960
rect 6568 2678 6866 2870
rect 6988 2870 7046 2960
rect 7046 2870 7146 2960
rect 7146 2870 7286 2960
rect 6988 2678 7286 2870
rect 7408 2870 7466 2960
rect 7466 2870 7566 2960
rect 7566 2870 7706 2960
rect 7408 2678 7706 2870
rect 7828 2870 7886 2960
rect 7886 2870 7986 2960
rect 7986 2870 8126 2960
rect 7828 2678 8126 2870
rect 8248 2870 8306 2960
rect 8306 2870 8406 2960
rect 8406 2870 8546 2960
rect 8248 2678 8546 2870
rect 8668 2870 8726 2960
rect 8726 2870 8826 2960
rect 8826 2870 8966 2960
rect 8668 2678 8966 2870
rect 9088 2870 9146 2960
rect 9146 2870 9246 2960
rect 9246 2870 9386 2960
rect 9088 2678 9386 2870
rect 10128 2954 10426 2960
rect 10128 2854 10208 2954
rect 10208 2854 10308 2954
rect 10308 2854 10426 2954
rect 10128 2678 10426 2854
rect 10578 2954 10876 2960
rect 10578 2854 10628 2954
rect 10628 2854 10728 2954
rect 10728 2854 10876 2954
rect 10578 2678 10876 2854
rect 10998 2954 11296 2960
rect 10998 2854 11048 2954
rect 11048 2854 11148 2954
rect 11148 2854 11296 2954
rect 10998 2678 11296 2854
rect 11418 2954 11716 2960
rect 11418 2854 11468 2954
rect 11468 2854 11568 2954
rect 11568 2854 11716 2954
rect 11418 2678 11716 2854
rect 11838 2954 12136 2960
rect 11838 2854 11888 2954
rect 11888 2854 11988 2954
rect 11988 2854 12136 2954
rect 11838 2678 12136 2854
rect 12258 2954 12556 2960
rect 12258 2854 12308 2954
rect 12308 2854 12408 2954
rect 12408 2854 12556 2954
rect 12258 2678 12556 2854
rect 12678 2954 12976 2960
rect 12678 2854 12728 2954
rect 12728 2854 12828 2954
rect 12828 2854 12976 2954
rect 12678 2678 12976 2854
rect 13098 2954 13396 2960
rect 13098 2854 13148 2954
rect 13148 2854 13248 2954
rect 13248 2854 13396 2954
rect 13098 2678 13396 2854
rect 13518 2954 13816 2960
rect 13518 2854 13568 2954
rect 13568 2854 13668 2954
rect 13668 2854 13816 2954
rect 13518 2678 13816 2854
rect 13938 2954 14236 2960
rect 13938 2854 13988 2954
rect 13988 2854 14088 2954
rect 14088 2854 14236 2954
rect 13938 2678 14236 2854
rect 14358 2954 14656 2960
rect 14358 2854 14408 2954
rect 14408 2854 14508 2954
rect 14508 2854 14656 2954
rect 14358 2678 14656 2854
rect 14778 2954 15076 2960
rect 14778 2854 14828 2954
rect 14828 2854 14928 2954
rect 14928 2854 15076 2954
rect 14778 2678 15076 2854
rect 15198 2954 15496 2960
rect 15198 2854 15248 2954
rect 15248 2854 15348 2954
rect 15348 2854 15496 2954
rect 15198 2678 15496 2854
rect 15618 2954 15916 2960
rect 15618 2854 15668 2954
rect 15668 2854 15768 2954
rect 15768 2854 15916 2954
rect 15618 2678 15916 2854
rect 16038 2954 16336 2960
rect 16038 2854 16088 2954
rect 16088 2854 16188 2954
rect 16188 2854 16336 2954
rect 16038 2678 16336 2854
rect 16458 2954 16756 2960
rect 16458 2854 16508 2954
rect 16508 2854 16608 2954
rect 16608 2854 16756 2954
rect 16458 2678 16756 2854
rect 16878 2954 17176 2960
rect 16878 2854 16928 2954
rect 16928 2854 17028 2954
rect 17028 2854 17176 2954
rect 16878 2678 17176 2854
rect 17298 2954 17596 2960
rect 17298 2854 17348 2954
rect 17348 2854 17448 2954
rect 17448 2854 17596 2954
rect 17298 2678 17596 2854
rect 17718 2954 18016 2960
rect 17718 2854 17768 2954
rect 17768 2854 17868 2954
rect 17868 2854 18016 2954
rect 17718 2678 18016 2854
rect 18138 2954 18436 2960
rect 18138 2854 18188 2954
rect 18188 2854 18288 2954
rect 18288 2854 18436 2954
rect 18138 2678 18436 2854
rect 18558 2954 18856 2960
rect 18558 2854 18608 2954
rect 18608 2854 18708 2954
rect 18708 2854 18856 2954
rect 18558 2678 18856 2854
rect 196 2220 524 2482
rect 196 -956 524 -694
rect 2492 -1476 2886 -1312
rect 2984 -1312 3128 -1164
rect 3338 -1434 3636 -1152
rect 3758 -1434 4056 -1152
rect 4178 -1434 4476 -1152
rect 4598 -1434 4896 -1152
rect 5298 -1344 5596 -1152
rect 5298 -1434 5366 -1344
rect 5366 -1434 5466 -1344
rect 5466 -1434 5596 -1344
rect 5728 -1344 6026 -1152
rect 5728 -1434 5786 -1344
rect 5786 -1434 5886 -1344
rect 5886 -1434 6026 -1344
rect 6148 -1344 6446 -1152
rect 6148 -1434 6206 -1344
rect 6206 -1434 6306 -1344
rect 6306 -1434 6446 -1344
rect 6568 -1344 6866 -1152
rect 6568 -1434 6626 -1344
rect 6626 -1434 6726 -1344
rect 6726 -1434 6866 -1344
rect 6988 -1344 7286 -1152
rect 6988 -1434 7046 -1344
rect 7046 -1434 7146 -1344
rect 7146 -1434 7286 -1344
rect 7408 -1344 7706 -1152
rect 7408 -1434 7466 -1344
rect 7466 -1434 7566 -1344
rect 7566 -1434 7706 -1344
rect 7828 -1344 8126 -1152
rect 7828 -1434 7886 -1344
rect 7886 -1434 7986 -1344
rect 7986 -1434 8126 -1344
rect 8248 -1344 8546 -1152
rect 8248 -1434 8306 -1344
rect 8306 -1434 8406 -1344
rect 8406 -1434 8546 -1344
rect 8668 -1344 8966 -1152
rect 8668 -1434 8726 -1344
rect 8726 -1434 8826 -1344
rect 8826 -1434 8966 -1344
rect 9088 -1344 9386 -1152
rect 9088 -1434 9146 -1344
rect 9146 -1434 9246 -1344
rect 9246 -1434 9386 -1344
rect 2490 -4272 2788 -3990
rect 2950 -4272 3248 -3990
rect 3350 -4272 3648 -3990
rect 3770 -4272 4068 -3990
rect 4190 -4272 4488 -3990
rect 5292 -7104 5490 -7032
rect 5490 -7104 5590 -7032
rect 5292 -7314 5590 -7104
rect 5712 -7104 5910 -7032
rect 5910 -7104 6010 -7032
rect 5712 -7314 6010 -7104
rect 6132 -7104 6330 -7032
rect 6330 -7104 6430 -7032
rect 6132 -7314 6430 -7104
rect 6552 -7104 6750 -7032
rect 6750 -7104 6850 -7032
rect 6552 -7314 6850 -7104
rect 6972 -7104 7170 -7032
rect 7170 -7104 7270 -7032
rect 6972 -7314 7270 -7104
rect 7392 -7104 7590 -7032
rect 7590 -7104 7690 -7032
rect 7392 -7314 7690 -7104
rect 7812 -7104 8010 -7032
rect 8010 -7104 8110 -7032
rect 7812 -7314 8110 -7104
rect 8232 -7104 8430 -7032
rect 8430 -7104 8530 -7032
rect 8232 -7314 8530 -7104
rect 8652 -7104 8850 -7032
rect 8850 -7104 8950 -7032
rect 8652 -7314 8950 -7104
rect 9072 -7104 9176 -7032
rect 9176 -7104 9276 -7032
rect 9276 -7104 9370 -7032
rect 9072 -7314 9370 -7104
<< metal3 >>
rect -14714 6676 612 18022
rect 10120 13618 10438 13623
rect 10120 13336 10130 13618
rect 10428 13336 10438 13618
rect 10120 13331 10438 13336
rect 10570 13618 10888 13623
rect 10570 13336 10580 13618
rect 10878 13336 10888 13618
rect 10570 13331 10888 13336
rect 10990 13618 11308 13623
rect 10990 13336 11000 13618
rect 11298 13336 11308 13618
rect 10990 13331 11308 13336
rect 11410 13618 11728 13623
rect 11410 13336 11420 13618
rect 11718 13336 11728 13618
rect 11410 13331 11728 13336
rect 11830 13618 12148 13623
rect 11830 13336 11840 13618
rect 12138 13336 12148 13618
rect 11830 13331 12148 13336
rect 12250 13618 12568 13623
rect 12250 13336 12260 13618
rect 12558 13336 12568 13618
rect 12250 13331 12568 13336
rect 12670 13618 12988 13623
rect 12670 13336 12680 13618
rect 12978 13336 12988 13618
rect 12670 13331 12988 13336
rect 13090 13618 13408 13623
rect 13090 13336 13100 13618
rect 13398 13336 13408 13618
rect 13090 13331 13408 13336
rect 13510 13618 13828 13623
rect 13510 13336 13520 13618
rect 13818 13336 13828 13618
rect 13510 13331 13828 13336
rect 13930 13618 14248 13623
rect 13930 13336 13940 13618
rect 14238 13336 14248 13618
rect 13930 13331 14248 13336
rect 14350 13618 14668 13623
rect 14350 13336 14360 13618
rect 14658 13336 14668 13618
rect 14350 13331 14668 13336
rect 14770 13618 15088 13623
rect 14770 13336 14780 13618
rect 15078 13336 15088 13618
rect 14770 13331 15088 13336
rect 15190 13618 15508 13623
rect 15190 13336 15200 13618
rect 15498 13336 15508 13618
rect 15190 13331 15508 13336
rect 15610 13618 15928 13623
rect 15610 13336 15620 13618
rect 15918 13336 15928 13618
rect 15610 13331 15928 13336
rect 16030 13618 16348 13623
rect 16030 13336 16040 13618
rect 16338 13336 16348 13618
rect 16030 13331 16348 13336
rect 16450 13618 16768 13623
rect 16450 13336 16460 13618
rect 16758 13336 16768 13618
rect 16450 13331 16768 13336
rect 16870 13618 17188 13623
rect 16870 13336 16880 13618
rect 17178 13336 17188 13618
rect 16870 13331 17188 13336
rect 17290 13618 17608 13623
rect 17290 13336 17300 13618
rect 17598 13336 17608 13618
rect 17290 13331 17608 13336
rect 17710 13618 18028 13623
rect 17710 13336 17720 13618
rect 18018 13336 18028 13618
rect 17710 13331 18028 13336
rect 18130 13618 18448 13623
rect 18130 13336 18140 13618
rect 18438 13336 18448 13618
rect 18130 13331 18448 13336
rect 18550 13618 18868 13623
rect 18550 13336 18560 13618
rect 18858 13336 18868 13618
rect 18550 13331 18868 13336
rect 2450 12788 4460 12846
rect 5276 12788 9352 12916
rect 2450 12506 3154 12788
rect 3452 12506 3574 12788
rect 3872 12506 3994 12788
rect 4292 12506 4414 12788
rect 4712 12506 4722 12788
rect 4824 12506 4834 12788
rect 5132 12506 5142 12788
rect 5244 12506 5254 12788
rect 5552 12506 5674 12788
rect 5972 12506 6094 12788
rect 6392 12506 6514 12788
rect 6812 12506 6934 12788
rect 7232 12506 7354 12788
rect 7652 12506 7774 12788
rect 8072 12506 8194 12788
rect 8492 12506 8614 12788
rect 8912 12506 9352 12788
rect 2450 12368 4460 12506
rect 5276 12368 9352 12506
rect 2450 12086 3154 12368
rect 3452 12086 3574 12368
rect 3872 12086 3994 12368
rect 4292 12086 4414 12368
rect 4712 12086 4722 12368
rect 4824 12086 4834 12368
rect 5132 12086 5142 12368
rect 5244 12086 5254 12368
rect 5552 12086 5674 12368
rect 5972 12086 6094 12368
rect 6392 12086 6514 12368
rect 6812 12086 6934 12368
rect 7232 12086 7354 12368
rect 7652 12086 7774 12368
rect 8072 12086 8194 12368
rect 8492 12086 8614 12368
rect 8912 12086 9352 12368
rect 2450 6676 4460 12086
rect 5276 7445 9352 12086
rect 5276 7440 9380 7445
rect 5276 7158 5292 7440
rect 5590 7158 5712 7440
rect 6010 7158 6132 7440
rect 6430 7158 6552 7440
rect 6850 7158 6972 7440
rect 7270 7158 7392 7440
rect 7690 7158 7812 7440
rect 8110 7158 8232 7440
rect 8530 7158 8652 7440
rect 8950 7158 9072 7440
rect 9370 7158 9380 7440
rect 5276 7153 9380 7158
rect 5276 6894 9352 7153
rect -14714 6314 4460 6676
rect -14714 2722 612 6314
rect 2450 5812 4460 6314
rect 2450 5798 4494 5812
rect 2450 5516 2490 5798
rect 2788 5516 2950 5798
rect 3248 5516 3350 5798
rect 3648 5516 3770 5798
rect 4068 5516 4190 5798
rect 4488 5516 4494 5798
rect 2450 5504 4494 5516
rect 2450 5260 4460 5504
rect 2482 3002 2896 3007
rect 2482 2838 2492 3002
rect 2886 2838 2896 3002
rect 3328 2960 3646 2965
rect 2482 2833 2896 2838
rect 2974 2838 3138 2843
rect 2974 2690 2984 2838
rect 3128 2690 3138 2838
rect 2974 2685 3138 2690
rect 3328 2678 3338 2960
rect 3636 2678 3646 2960
rect 3328 2673 3646 2678
rect 3748 2960 4066 2965
rect 3748 2678 3758 2960
rect 4056 2678 4066 2960
rect 3748 2673 4066 2678
rect 4168 2960 4486 2965
rect 4168 2678 4178 2960
rect 4476 2678 4486 2960
rect 4168 2673 4486 2678
rect 4588 2960 4906 2965
rect 4588 2678 4598 2960
rect 4896 2678 4906 2960
rect 4588 2673 4906 2678
rect 5288 2960 5606 2965
rect 5288 2678 5298 2960
rect 5596 2678 5606 2960
rect 5288 2673 5606 2678
rect 5718 2960 6036 2965
rect 5718 2678 5728 2960
rect 6026 2678 6036 2960
rect 5718 2673 6036 2678
rect 6138 2960 6456 2965
rect 6138 2678 6148 2960
rect 6446 2678 6456 2960
rect 6138 2673 6456 2678
rect 6558 2960 6876 2965
rect 6558 2678 6568 2960
rect 6866 2678 6876 2960
rect 6558 2673 6876 2678
rect 6978 2960 7296 2965
rect 6978 2678 6988 2960
rect 7286 2678 7296 2960
rect 6978 2673 7296 2678
rect 7398 2960 7716 2965
rect 7398 2678 7408 2960
rect 7706 2678 7716 2960
rect 7398 2673 7716 2678
rect 7818 2960 8136 2965
rect 7818 2678 7828 2960
rect 8126 2678 8136 2960
rect 7818 2673 8136 2678
rect 8238 2960 8556 2965
rect 8238 2678 8248 2960
rect 8546 2678 8556 2960
rect 8238 2673 8556 2678
rect 8658 2960 8976 2965
rect 8658 2678 8668 2960
rect 8966 2678 8976 2960
rect 8658 2673 8976 2678
rect 9078 2960 9396 2965
rect 9078 2678 9088 2960
rect 9386 2678 9396 2960
rect 9078 2673 9396 2678
rect 10118 2960 10436 2965
rect 10118 2678 10128 2960
rect 10426 2678 10436 2960
rect 10118 2673 10436 2678
rect 10568 2960 10886 2965
rect 10568 2678 10578 2960
rect 10876 2678 10886 2960
rect 10568 2673 10886 2678
rect 10988 2960 11306 2965
rect 10988 2678 10998 2960
rect 11296 2678 11306 2960
rect 10988 2673 11306 2678
rect 11408 2960 11726 2965
rect 11408 2678 11418 2960
rect 11716 2678 11726 2960
rect 11408 2673 11726 2678
rect 11828 2960 12146 2965
rect 11828 2678 11838 2960
rect 12136 2678 12146 2960
rect 11828 2673 12146 2678
rect 12248 2960 12566 2965
rect 12248 2678 12258 2960
rect 12556 2678 12566 2960
rect 12248 2673 12566 2678
rect 12668 2960 12986 2965
rect 12668 2678 12678 2960
rect 12976 2678 12986 2960
rect 12668 2673 12986 2678
rect 13088 2960 13406 2965
rect 13088 2678 13098 2960
rect 13396 2678 13406 2960
rect 13088 2673 13406 2678
rect 13508 2960 13826 2965
rect 13508 2678 13518 2960
rect 13816 2678 13826 2960
rect 13508 2673 13826 2678
rect 13928 2960 14246 2965
rect 13928 2678 13938 2960
rect 14236 2678 14246 2960
rect 13928 2673 14246 2678
rect 14348 2960 14666 2965
rect 14348 2678 14358 2960
rect 14656 2678 14666 2960
rect 14348 2673 14666 2678
rect 14768 2960 15086 2965
rect 14768 2678 14778 2960
rect 15076 2678 15086 2960
rect 14768 2673 15086 2678
rect 15188 2960 15506 2965
rect 15188 2678 15198 2960
rect 15496 2678 15506 2960
rect 15188 2673 15506 2678
rect 15608 2960 15926 2965
rect 15608 2678 15618 2960
rect 15916 2678 15926 2960
rect 15608 2673 15926 2678
rect 16028 2960 16346 2965
rect 16028 2678 16038 2960
rect 16336 2678 16346 2960
rect 16028 2673 16346 2678
rect 16448 2960 16766 2965
rect 16448 2678 16458 2960
rect 16756 2678 16766 2960
rect 16448 2673 16766 2678
rect 16868 2960 17186 2965
rect 16868 2678 16878 2960
rect 17176 2678 17186 2960
rect 16868 2673 17186 2678
rect 17288 2960 17606 2965
rect 17288 2678 17298 2960
rect 17596 2678 17606 2960
rect 17288 2673 17606 2678
rect 17708 2960 18026 2965
rect 17708 2678 17718 2960
rect 18016 2678 18026 2960
rect 17708 2673 18026 2678
rect 18128 2960 18446 2965
rect 18128 2678 18138 2960
rect 18436 2678 18446 2960
rect 18128 2673 18446 2678
rect 18548 2960 18866 2965
rect 18548 2678 18558 2960
rect 18856 2678 18866 2960
rect 18548 2673 18866 2678
rect 186 2482 534 2487
rect 186 2220 196 2482
rect 524 2220 534 2482
rect 186 2215 534 2220
rect -184 726 -80 800
rect -18 798 90 802
rect -18 728 102 798
rect -18 724 90 728
rect 186 -694 534 -689
rect 186 -956 196 -694
rect 524 -956 534 -694
rect 186 -961 534 -956
rect 3328 -1152 3646 -1147
rect 2974 -1164 3138 -1159
rect -14714 -4788 612 -1196
rect 2482 -1312 2896 -1307
rect 2482 -1476 2492 -1312
rect 2886 -1476 2896 -1312
rect 2974 -1312 2984 -1164
rect 3128 -1312 3138 -1164
rect 2974 -1317 3138 -1312
rect 3328 -1434 3338 -1152
rect 3636 -1434 3646 -1152
rect 3328 -1439 3646 -1434
rect 3748 -1152 4066 -1147
rect 3748 -1434 3758 -1152
rect 4056 -1434 4066 -1152
rect 3748 -1439 4066 -1434
rect 4168 -1152 4486 -1147
rect 4168 -1434 4178 -1152
rect 4476 -1434 4486 -1152
rect 4168 -1439 4486 -1434
rect 4588 -1152 4906 -1147
rect 4588 -1434 4598 -1152
rect 4896 -1434 4906 -1152
rect 4588 -1439 4906 -1434
rect 5288 -1152 5606 -1147
rect 5288 -1434 5298 -1152
rect 5596 -1434 5606 -1152
rect 5288 -1439 5606 -1434
rect 5718 -1152 6036 -1147
rect 5718 -1434 5728 -1152
rect 6026 -1434 6036 -1152
rect 5718 -1439 6036 -1434
rect 6138 -1152 6456 -1147
rect 6138 -1434 6148 -1152
rect 6446 -1434 6456 -1152
rect 6138 -1439 6456 -1434
rect 6558 -1152 6876 -1147
rect 6558 -1434 6568 -1152
rect 6866 -1434 6876 -1152
rect 6558 -1439 6876 -1434
rect 6978 -1152 7296 -1147
rect 6978 -1434 6988 -1152
rect 7286 -1434 7296 -1152
rect 6978 -1439 7296 -1434
rect 7398 -1152 7716 -1147
rect 7398 -1434 7408 -1152
rect 7706 -1434 7716 -1152
rect 7398 -1439 7716 -1434
rect 7818 -1152 8136 -1147
rect 7818 -1434 7828 -1152
rect 8126 -1434 8136 -1152
rect 7818 -1439 8136 -1434
rect 8238 -1152 8556 -1147
rect 8238 -1434 8248 -1152
rect 8546 -1434 8556 -1152
rect 8238 -1439 8556 -1434
rect 8658 -1152 8976 -1147
rect 8658 -1434 8668 -1152
rect 8966 -1434 8976 -1152
rect 8658 -1439 8976 -1434
rect 9078 -1152 9396 -1147
rect 9078 -1434 9088 -1152
rect 9386 -1434 9396 -1152
rect 9078 -1439 9396 -1434
rect 2482 -1481 2896 -1476
rect 2450 -3978 4460 -3734
rect 2450 -3990 4494 -3978
rect 2450 -4272 2490 -3990
rect 2788 -4272 2950 -3990
rect 3248 -4272 3350 -3990
rect 3648 -4272 3770 -3990
rect 4068 -4272 4190 -3990
rect 4488 -4272 4494 -3990
rect 2450 -4286 4494 -4272
rect 2450 -4788 4460 -4286
rect -14714 -5150 4460 -4788
rect -14714 -16496 612 -5150
rect 2450 -10560 4460 -5150
rect 5276 -7027 9352 -6768
rect 5276 -7032 9380 -7027
rect 5276 -7314 5292 -7032
rect 5590 -7314 5712 -7032
rect 6010 -7314 6132 -7032
rect 6430 -7314 6552 -7032
rect 6850 -7314 6972 -7032
rect 7270 -7314 7392 -7032
rect 7690 -7314 7812 -7032
rect 8110 -7314 8232 -7032
rect 8530 -7314 8652 -7032
rect 8950 -7314 9072 -7032
rect 9370 -7314 9380 -7032
rect 5276 -7319 9380 -7314
rect 5276 -10560 9352 -7319
rect 2450 -10842 3154 -10560
rect 3452 -10842 3574 -10560
rect 3872 -10842 3994 -10560
rect 4292 -10842 4414 -10560
rect 4712 -10842 4722 -10560
rect 4824 -10842 4834 -10560
rect 5132 -10842 5142 -10560
rect 5244 -10842 5254 -10560
rect 5552 -10842 5674 -10560
rect 5972 -10842 6094 -10560
rect 6392 -10842 6514 -10560
rect 6812 -10842 6934 -10560
rect 7232 -10842 7354 -10560
rect 7652 -10842 7774 -10560
rect 8072 -10842 8194 -10560
rect 8492 -10842 8614 -10560
rect 8912 -10842 9352 -10560
rect 2450 -10980 4460 -10842
rect 5276 -10980 9352 -10842
rect 2450 -11262 3154 -10980
rect 3452 -11262 3574 -10980
rect 3872 -11262 3994 -10980
rect 4292 -11262 4414 -10980
rect 4712 -11262 4722 -10980
rect 4824 -11262 4834 -10980
rect 5132 -11262 5142 -10980
rect 5244 -11262 5254 -10980
rect 5552 -11262 5674 -10980
rect 5972 -11262 6094 -10980
rect 6392 -11262 6514 -10980
rect 6812 -11262 6934 -10980
rect 7232 -11262 7354 -10980
rect 7652 -11262 7774 -10980
rect 8072 -11262 8194 -10980
rect 8492 -11262 8614 -10980
rect 8912 -11262 9352 -10980
rect 2450 -11320 4460 -11262
rect 5276 -11390 9352 -11262
<< via3 >>
rect 10130 13336 10428 13618
rect 10580 13336 10878 13618
rect 11000 13336 11298 13618
rect 11420 13336 11718 13618
rect 11840 13336 12138 13618
rect 12260 13336 12558 13618
rect 12680 13336 12978 13618
rect 13100 13336 13398 13618
rect 13520 13336 13818 13618
rect 13940 13336 14238 13618
rect 14360 13336 14658 13618
rect 14780 13336 15078 13618
rect 15200 13336 15498 13618
rect 15620 13336 15918 13618
rect 16040 13336 16338 13618
rect 16460 13336 16758 13618
rect 16880 13336 17178 13618
rect 17300 13336 17598 13618
rect 17720 13336 18018 13618
rect 18140 13336 18438 13618
rect 18560 13336 18858 13618
rect 3154 12506 3452 12788
rect 3574 12506 3872 12788
rect 3994 12506 4292 12788
rect 4414 12506 4712 12788
rect 4834 12506 5132 12788
rect 5254 12506 5552 12788
rect 5674 12506 5972 12788
rect 6094 12506 6392 12788
rect 6514 12506 6812 12788
rect 6934 12506 7232 12788
rect 7354 12506 7652 12788
rect 7774 12506 8072 12788
rect 8194 12506 8492 12788
rect 8614 12506 8912 12788
rect 3154 12086 3452 12368
rect 3574 12086 3872 12368
rect 3994 12086 4292 12368
rect 4414 12086 4712 12368
rect 4834 12086 5132 12368
rect 5254 12086 5552 12368
rect 5674 12086 5972 12368
rect 6094 12086 6392 12368
rect 6514 12086 6812 12368
rect 6934 12086 7232 12368
rect 7354 12086 7652 12368
rect 7774 12086 8072 12368
rect 8194 12086 8492 12368
rect 8614 12086 8912 12368
rect 2492 2838 2886 3002
rect 2984 2690 3128 2838
rect 3338 2678 3636 2960
rect 3758 2678 4056 2960
rect 4178 2678 4476 2960
rect 4598 2678 4896 2960
rect 5298 2678 5596 2960
rect 5728 2678 6026 2960
rect 6148 2678 6446 2960
rect 6568 2678 6866 2960
rect 6988 2678 7286 2960
rect 7408 2678 7706 2960
rect 7828 2678 8126 2960
rect 8248 2678 8546 2960
rect 8668 2678 8966 2960
rect 9088 2678 9386 2960
rect 10128 2678 10426 2960
rect 10578 2678 10876 2960
rect 10998 2678 11296 2960
rect 11418 2678 11716 2960
rect 11838 2678 12136 2960
rect 12258 2678 12556 2960
rect 12678 2678 12976 2960
rect 13098 2678 13396 2960
rect 13518 2678 13816 2960
rect 13938 2678 14236 2960
rect 14358 2678 14656 2960
rect 14778 2678 15076 2960
rect 15198 2678 15496 2960
rect 15618 2678 15916 2960
rect 16038 2678 16336 2960
rect 16458 2678 16756 2960
rect 16878 2678 17176 2960
rect 17298 2678 17596 2960
rect 17718 2678 18016 2960
rect 18138 2678 18436 2960
rect 18558 2678 18856 2960
rect 196 2220 524 2482
rect 196 -956 524 -694
rect 2492 -1476 2886 -1312
rect 2984 -1312 3128 -1164
rect 3338 -1434 3636 -1152
rect 3758 -1434 4056 -1152
rect 4178 -1434 4476 -1152
rect 4598 -1434 4896 -1152
rect 5298 -1434 5596 -1152
rect 5728 -1434 6026 -1152
rect 6148 -1434 6446 -1152
rect 6568 -1434 6866 -1152
rect 6988 -1434 7286 -1152
rect 7408 -1434 7706 -1152
rect 7828 -1434 8126 -1152
rect 8248 -1434 8546 -1152
rect 8668 -1434 8966 -1152
rect 9088 -1434 9386 -1152
rect 3154 -10842 3452 -10560
rect 3574 -10842 3872 -10560
rect 3994 -10842 4292 -10560
rect 4414 -10842 4712 -10560
rect 4834 -10842 5132 -10560
rect 5254 -10842 5552 -10560
rect 5674 -10842 5972 -10560
rect 6094 -10842 6392 -10560
rect 6514 -10842 6812 -10560
rect 6934 -10842 7232 -10560
rect 7354 -10842 7652 -10560
rect 7774 -10842 8072 -10560
rect 8194 -10842 8492 -10560
rect 8614 -10842 8912 -10560
rect 3154 -11262 3452 -10980
rect 3574 -11262 3872 -10980
rect 3994 -11262 4292 -10980
rect 4414 -11262 4712 -10980
rect 4834 -11262 5132 -10980
rect 5254 -11262 5552 -10980
rect 5674 -11262 5972 -10980
rect 6094 -11262 6392 -10980
rect 6514 -11262 6812 -10980
rect 6934 -11262 7232 -10980
rect 7354 -11262 7652 -10980
rect 7774 -11262 8072 -10980
rect 8194 -11262 8492 -10980
rect 8614 -11262 8912 -10980
<< mimcap >>
rect -14613 17882 -11063 17922
rect -14613 14412 -14573 17882
rect -11103 14412 -11063 17882
rect -14613 14372 -11063 14412
rect -10744 17882 -7194 17922
rect -10744 14412 -10704 17882
rect -7234 14412 -7194 17882
rect -10744 14372 -7194 14412
rect -6875 17882 -3325 17922
rect -6875 14412 -6835 17882
rect -3365 14412 -3325 17882
rect -6875 14372 -3325 14412
rect -3006 17882 544 17922
rect -3006 14412 -2966 17882
rect 504 14412 544 17882
rect -3006 14372 544 14412
rect -14613 14032 -11063 14072
rect -14613 10562 -14573 14032
rect -11103 10562 -11063 14032
rect -14613 10522 -11063 10562
rect -10744 14032 -7194 14072
rect -10744 10562 -10704 14032
rect -7234 10562 -7194 14032
rect -10744 10522 -7194 10562
rect -6875 14032 -3325 14072
rect -6875 10562 -6835 14032
rect -3365 10562 -3325 14032
rect -6875 10522 -3325 10562
rect -3006 14032 544 14072
rect -3006 10562 -2966 14032
rect 504 10562 544 14032
rect -3006 10522 544 10562
rect -14613 10182 -11063 10222
rect -14613 6712 -14573 10182
rect -11103 6712 -11063 10182
rect -14613 6672 -11063 6712
rect -10744 10182 -7194 10222
rect -10744 6712 -10704 10182
rect -7234 6712 -7194 10182
rect -10744 6672 -7194 6712
rect -6875 10182 -3325 10222
rect -6875 6712 -6835 10182
rect -3365 6712 -3325 10182
rect -6875 6672 -3325 6712
rect -3006 10182 544 10222
rect -3006 6712 -2966 10182
rect 504 6712 544 10182
rect -3006 6672 544 6712
rect -14613 6332 -11063 6372
rect -14613 2862 -14573 6332
rect -11103 2862 -11063 6332
rect -14613 2822 -11063 2862
rect -10744 6332 -7194 6372
rect -10744 2862 -10704 6332
rect -7234 2862 -7194 6332
rect -10744 2822 -7194 2862
rect -6875 6332 -3325 6372
rect -6875 2862 -6835 6332
rect -3365 2862 -3325 6332
rect -6875 2822 -3325 2862
rect -3006 6332 544 6372
rect -3006 2862 -2966 6332
rect 504 2862 544 6332
rect -3006 2822 544 2862
rect -14613 -1336 -11063 -1296
rect -14613 -4806 -14573 -1336
rect -11103 -4806 -11063 -1336
rect -14613 -4846 -11063 -4806
rect -10744 -1336 -7194 -1296
rect -10744 -4806 -10704 -1336
rect -7234 -4806 -7194 -1336
rect -10744 -4846 -7194 -4806
rect -6875 -1336 -3325 -1296
rect -6875 -4806 -6835 -1336
rect -3365 -4806 -3325 -1336
rect -6875 -4846 -3325 -4806
rect -3006 -1336 544 -1296
rect -3006 -4806 -2966 -1336
rect 504 -4806 544 -1336
rect -3006 -4846 544 -4806
rect -14613 -5186 -11063 -5146
rect -14613 -8656 -14573 -5186
rect -11103 -8656 -11063 -5186
rect -14613 -8696 -11063 -8656
rect -10744 -5186 -7194 -5146
rect -10744 -8656 -10704 -5186
rect -7234 -8656 -7194 -5186
rect -10744 -8696 -7194 -8656
rect -6875 -5186 -3325 -5146
rect -6875 -8656 -6835 -5186
rect -3365 -8656 -3325 -5186
rect -6875 -8696 -3325 -8656
rect -3006 -5186 544 -5146
rect -3006 -8656 -2966 -5186
rect 504 -8656 544 -5186
rect -3006 -8696 544 -8656
rect -14613 -9036 -11063 -8996
rect -14613 -12506 -14573 -9036
rect -11103 -12506 -11063 -9036
rect -14613 -12546 -11063 -12506
rect -10744 -9036 -7194 -8996
rect -10744 -12506 -10704 -9036
rect -7234 -12506 -7194 -9036
rect -10744 -12546 -7194 -12506
rect -6875 -9036 -3325 -8996
rect -6875 -12506 -6835 -9036
rect -3365 -12506 -3325 -9036
rect -6875 -12546 -3325 -12506
rect -3006 -9036 544 -8996
rect -3006 -12506 -2966 -9036
rect 504 -12506 544 -9036
rect -3006 -12546 544 -12506
rect -14613 -12886 -11063 -12846
rect -14613 -16356 -14573 -12886
rect -11103 -16356 -11063 -12886
rect -14613 -16396 -11063 -16356
rect -10744 -12886 -7194 -12846
rect -10744 -16356 -10704 -12886
rect -7234 -16356 -7194 -12886
rect -10744 -16396 -7194 -16356
rect -6875 -12886 -3325 -12846
rect -6875 -16356 -6835 -12886
rect -3365 -16356 -3325 -12886
rect -6875 -16396 -3325 -16356
rect -3006 -12886 544 -12846
rect -3006 -16356 -2966 -12886
rect 504 -16356 544 -12886
rect -3006 -16396 544 -16356
<< mimcapcontact >>
rect -14573 14412 -11103 17882
rect -10704 14412 -7234 17882
rect -6835 14412 -3365 17882
rect -2966 14412 504 17882
rect -14573 10562 -11103 14032
rect -10704 10562 -7234 14032
rect -6835 10562 -3365 14032
rect -2966 10562 504 14032
rect -14573 6712 -11103 10182
rect -10704 6712 -7234 10182
rect -6835 6712 -3365 10182
rect -2966 6712 504 10182
rect -14573 2862 -11103 6332
rect -10704 2862 -7234 6332
rect -6835 2862 -3365 6332
rect -2966 2862 504 6332
rect -14573 -4806 -11103 -1336
rect -10704 -4806 -7234 -1336
rect -6835 -4806 -3365 -1336
rect -2966 -4806 504 -1336
rect -14573 -8656 -11103 -5186
rect -10704 -8656 -7234 -5186
rect -6835 -8656 -3365 -5186
rect -2966 -8656 504 -5186
rect -14573 -12506 -11103 -9036
rect -10704 -12506 -7234 -9036
rect -6835 -12506 -3365 -9036
rect -2966 -12506 504 -9036
rect -14573 -16356 -11103 -12886
rect -10704 -16356 -7234 -12886
rect -6835 -16356 -3365 -12886
rect -2966 -16356 504 -12886
<< metal4 >>
rect -12890 18022 -12786 18072
rect -9021 18022 -8917 18072
rect -5152 18022 -5048 18072
rect -1283 18022 -1179 18072
rect -14714 17882 612 18022
rect -14714 14412 -14573 17882
rect -11103 14412 -10704 17882
rect -7234 14412 -6835 17882
rect -3365 14412 -2966 17882
rect 504 14412 612 17882
rect -14714 14032 612 14412
rect 9376 14200 19390 14210
rect -14714 10562 -14573 14032
rect -11103 10562 -10704 14032
rect -7234 10562 -6835 14032
rect -3365 10562 -2966 14032
rect 504 10562 612 14032
rect 2800 13618 19390 14200
rect 2800 13542 10130 13618
rect 2774 13336 10130 13542
rect 10428 13336 10580 13618
rect 10878 13336 11000 13618
rect 11298 13336 11420 13618
rect 11718 13336 11840 13618
rect 12138 13336 12260 13618
rect 12558 13336 12680 13618
rect 12978 13336 13100 13618
rect 13398 13336 13520 13618
rect 13818 13336 13940 13618
rect 14238 13336 14360 13618
rect 14658 13336 14780 13618
rect 15078 13336 15200 13618
rect 15498 13336 15620 13618
rect 15918 13336 16040 13618
rect 16338 13336 16460 13618
rect 16758 13336 16880 13618
rect 17178 13336 17300 13618
rect 17598 13336 17720 13618
rect 18018 13336 18140 13618
rect 18438 13336 18560 13618
rect 18858 13336 19390 13618
rect 2774 12788 19390 13336
rect 2774 12716 3154 12788
rect -14714 10182 612 10562
rect -14714 6712 -14573 10182
rect -11103 6712 -10704 10182
rect -7234 6712 -6835 10182
rect -3365 6712 -2966 10182
rect 504 6712 612 10182
rect 2772 12506 3154 12716
rect 3452 12506 3574 12788
rect 3872 12506 3994 12788
rect 4292 12506 4414 12788
rect 4712 12506 4834 12788
rect 5132 12506 5254 12788
rect 5552 12506 5674 12788
rect 5972 12506 6094 12788
rect 6392 12506 6514 12788
rect 6812 12506 6934 12788
rect 7232 12506 7354 12788
rect 7652 12506 7774 12788
rect 8072 12506 8194 12788
rect 8492 12506 8614 12788
rect 8912 12506 19390 12788
rect 2772 12368 19390 12506
rect 2772 12086 3154 12368
rect 3452 12086 3574 12368
rect 3872 12086 3994 12368
rect 4292 12086 4414 12368
rect 4712 12086 4834 12368
rect 5132 12086 5254 12368
rect 5552 12086 5674 12368
rect 5972 12086 6094 12368
rect 6392 12086 6514 12368
rect 6812 12086 6934 12368
rect 7232 12086 7354 12368
rect 7652 12086 7774 12368
rect 8072 12086 8194 12368
rect 8492 12086 8614 12368
rect 8912 12086 19390 12368
rect 2772 11900 19390 12086
rect 2772 7716 3130 11900
rect -14714 6332 612 6712
rect -14714 2862 -14573 6332
rect -11103 2862 -10704 6332
rect -7234 2862 -6835 6332
rect -3365 2862 -2966 6332
rect 504 2862 612 6332
rect -14714 2722 612 2862
rect 858 7460 3130 7716
rect 274 2483 446 2722
rect 858 2650 1098 7460
rect 195 2482 525 2483
rect 195 2220 196 2482
rect 524 2220 525 2482
rect 195 2219 525 2220
rect 856 2122 1098 2650
rect 2080 3002 19064 3024
rect 2080 2838 2492 3002
rect 2886 2960 19064 3002
rect 2886 2838 3338 2960
rect 2080 2690 2984 2838
rect 3128 2690 3338 2838
rect 2080 2678 3338 2690
rect 3636 2678 3758 2960
rect 4056 2678 4178 2960
rect 4476 2678 4598 2960
rect 4896 2678 5298 2960
rect 5596 2678 5728 2960
rect 6026 2678 6148 2960
rect 6446 2678 6568 2960
rect 6866 2678 6988 2960
rect 7286 2678 7408 2960
rect 7706 2678 7828 2960
rect 8126 2678 8248 2960
rect 8546 2678 8668 2960
rect 8966 2678 9088 2960
rect 9386 2678 10128 2960
rect 10426 2678 10578 2960
rect 10876 2678 10998 2960
rect 11296 2678 11418 2960
rect 11716 2678 11838 2960
rect 12136 2678 12258 2960
rect 12556 2678 12678 2960
rect 12976 2678 13098 2960
rect 13396 2678 13518 2960
rect 13816 2678 13938 2960
rect 14236 2678 14358 2960
rect 14656 2678 14778 2960
rect 15076 2678 15198 2960
rect 15496 2678 15618 2960
rect 15916 2678 16038 2960
rect 16336 2678 16458 2960
rect 16756 2678 16878 2960
rect 17176 2678 17298 2960
rect 17596 2678 17718 2960
rect 18016 2678 18138 2960
rect 18436 2678 18558 2960
rect 18856 2678 19064 2960
rect -182 2016 1108 2122
rect 2080 1428 19064 2678
rect -1172 254 19064 1428
rect -708 -490 -538 -326
rect -708 -594 1098 -490
rect 195 -694 525 -693
rect 195 -956 196 -694
rect 524 -956 525 -694
rect 195 -957 525 -956
rect 274 -1196 446 -957
rect -14714 -1336 612 -1196
rect -14714 -4806 -14573 -1336
rect -11103 -4806 -10704 -1336
rect -7234 -4806 -6835 -1336
rect -3365 -4806 -2966 -1336
rect 504 -4806 612 -1336
rect -14714 -5186 612 -4806
rect -14714 -8656 -14573 -5186
rect -11103 -8656 -10704 -5186
rect -7234 -8656 -6835 -5186
rect -3365 -8656 -2966 -5186
rect 504 -8656 612 -5186
rect 858 -5934 1098 -594
rect 2080 -1152 19064 254
rect 2080 -1164 3338 -1152
rect 2080 -1312 2984 -1164
rect 3128 -1312 3338 -1164
rect 2080 -1476 2492 -1312
rect 2886 -1434 3338 -1312
rect 3636 -1434 3758 -1152
rect 4056 -1434 4178 -1152
rect 4476 -1434 4598 -1152
rect 4896 -1434 5298 -1152
rect 5596 -1434 5728 -1152
rect 6026 -1434 6148 -1152
rect 6446 -1434 6568 -1152
rect 6866 -1434 6988 -1152
rect 7286 -1434 7408 -1152
rect 7706 -1434 7828 -1152
rect 8126 -1434 8248 -1152
rect 8546 -1434 8668 -1152
rect 8966 -1434 9088 -1152
rect 9386 -1434 19064 -1152
rect 2886 -1476 19064 -1434
rect 2080 -1498 19064 -1476
rect 858 -6190 3130 -5934
rect -14714 -9036 612 -8656
rect -14714 -12506 -14573 -9036
rect -11103 -12506 -10704 -9036
rect -7234 -12506 -6835 -9036
rect -3365 -12506 -2966 -9036
rect 504 -12506 612 -9036
rect 2772 -10464 3130 -6190
rect 2772 -10560 9446 -10464
rect 2772 -10842 3154 -10560
rect 3452 -10842 3574 -10560
rect 3872 -10842 3994 -10560
rect 4292 -10842 4414 -10560
rect 4712 -10842 4834 -10560
rect 5132 -10842 5254 -10560
rect 5552 -10842 5674 -10560
rect 5972 -10842 6094 -10560
rect 6392 -10842 6514 -10560
rect 6812 -10842 6934 -10560
rect 7232 -10842 7354 -10560
rect 7652 -10842 7774 -10560
rect 8072 -10842 8194 -10560
rect 8492 -10842 8614 -10560
rect 8912 -10842 9446 -10560
rect 2772 -10980 9446 -10842
rect 2772 -11262 3154 -10980
rect 3452 -11262 3574 -10980
rect 3872 -11262 3994 -10980
rect 4292 -11262 4414 -10980
rect 4712 -11262 4834 -10980
rect 5132 -11262 5254 -10980
rect 5552 -11262 5674 -10980
rect 5972 -11262 6094 -10980
rect 6392 -11262 6514 -10980
rect 6812 -11262 6934 -10980
rect 7232 -11262 7354 -10980
rect 7652 -11262 7774 -10980
rect 8072 -11262 8194 -10980
rect 8492 -11262 8614 -10980
rect 8912 -11262 9446 -10980
rect 2772 -12016 9446 -11262
rect -14714 -12886 612 -12506
rect -14714 -16356 -14573 -12886
rect -11103 -16356 -10704 -12886
rect -7234 -16356 -6835 -12886
rect -3365 -16356 -2966 -12886
rect 504 -16356 612 -12886
rect -14714 -16496 612 -16356
use nand  nand_0 ~/magic/class_d_audio_amplifier/nand
timestamp 1628437904
transform 1 0 106 0 1 -1138
box -512 542 18 1882
use nand  nand_1
timestamp 1628437904
transform 1 0 106 0 -1 2664
box -512 542 18 1882
use inverter  inverter_0 ~/magic/class_d_audio_amplifier/inverter
timestamp 1628437795
transform 1 0 -238 0 1 -2230
box -622 1804 -274 2934
<< labels >>
flabel metal4 11848 246 11848 246 0 FreeSans 8000 0 0 0 vdd
port 0 nsew
flabel metal2 8334 -4172 8334 -4172 0 FreeSans 8000 0 0 0 vn
port 3 nsew
flabel metal1 2824 4476 2824 4476 0 FreeSans 8000 0 0 0 vp1
flabel metal1 2814 -3050 2814 -3050 0 FreeSans 8000 0 0 0 vn1
flabel metal1 5174 5910 5174 5910 0 FreeSans 1600 0 0 0 vp2
flabel metal1 -914 144 -914 144 0 FreeSans 8000 0 0 0 vin
port 1 nsew
flabel metal1 9632 7278 9632 7278 0 FreeSans 8000 0 0 0 vp3
flabel metal2 17426 8700 17426 8700 0 FreeSans 8000 0 0 0 vp
port 2 nsew
flabel metal1 5128 -5754 5128 -5754 0 FreeSans 8000 0 0 0 vn2
<< end >>
