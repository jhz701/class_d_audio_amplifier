.subckt integrator_input in out
.param R1=10k CF=20p
.model int_fb int(in_offset=0 gain=2e6 out_lower_limit=-100 out_upper_limit=100 limit_range=1e-9 out_ic=0.9)

aint in out int_fb
.ends
