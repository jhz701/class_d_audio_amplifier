* NGSPICE file created from output_driver_post.ext - technology: sky130A

.subckt output_driver_post vdd1 vp_p out_p vss vp_n vn_p out_n vn_n vdd2
X0 out_n.t1761 vn_p.t0 vdd2.t1499 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1 out_n.t1760 vn_p.t1 vdd2.t1498 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2 vdd2.t1497 vn_p.t2 out_n.t1759 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3 out_n.t1758 vn_p.t3 vdd2.t1496 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4 vdd1.t1499 vp_p.t0 out_p.t946 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5 vdd1.t1498 vp_p.t1 out_p.t1090 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6 out_n.t1757 vn_p.t4 vdd2.t1495 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7 out_p.t1094 vp_p.t2 vdd1.t1497 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8 vdd2.t1494 vn_p.t5 out_n.t1756 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9 out_n.t1755 vn_p.t6 vdd2.t1493 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10 vdd2.t1492 vn_p.t7 out_n.t1754 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X11 out_n.t1753 vn_p.t8 vdd2.t1491 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X12 vss.t561 vp_n.t0 out_p.t1777 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 vdd2.t1490 vn_p.t9 out_n.t1752 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14 vss.t258 vn_n.t0 out_n.t258 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X15 out_n.t1751 vn_p.t10 vdd2.t1489 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X16 out_n.t1750 vn_p.t11 vdd2.t1488 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X17 out_n.t1749 vn_p.t12 vdd2.t1487 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 out_n.t1748 vn_p.t13 vdd2.t1486 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 vdd2.t1485 vn_p.t14 out_n.t1747 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X20 out_n.t1746 vn_p.t15 vdd2.t1484 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X21 out_p.t1778 vp_n.t1 vss.t560 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X22 vdd2.t1483 vn_p.t16 out_n.t1745 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X23 vdd2.t1482 vn_p.t17 out_n.t1744 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X24 out_n.t259 vn_n.t1 vss.t259 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X25 vdd2.t1481 vn_p.t18 out_n.t1743 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X26 out_p.t606 vp_p.t3 vdd1.t1496 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X27 vdd1.t1495 vp_p.t4 out_p.t607 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X28 vdd2.t1480 vn_p.t19 out_n.t1742 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X29 out_p.t608 vp_p.t5 vdd1.t1494 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X30 vdd1.t1493 vp_p.t6 out_p.t598 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X31 out_n.t1741 vn_p.t20 vdd2.t1479 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X32 out_p.t599 vp_p.t7 vdd1.t1492 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X33 out_p.t610 vp_p.t8 vdd1.t1491 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X34 vdd2.t1478 vn_p.t21 out_n.t1740 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X35 out_p.t600 vp_p.t9 vdd1.t1490 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X36 vdd1.t1489 vp_p.t10 out_p.t588 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X37 vdd2.t1477 vn_p.t22 out_n.t1739 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X38 vdd1.t1488 vp_p.t11 out_p.t601 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X39 out_p.t589 vp_p.t12 vdd1.t1487 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X40 out_p.t602 vp_p.t13 vdd1.t1486 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X41 vdd1.t1485 vp_p.t14 out_p.t590 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X42 out_n.t260 vn_n.t2 vss.t260 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X43 vdd2.t1476 vn_p.t23 out_n.t1738 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X44 out_n.t1737 vn_p.t24 vdd2.t1475 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X45 out_n.t1736 vn_p.t25 vdd2.t1474 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X46 vdd2.t1473 vn_p.t26 out_n.t1735 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X47 vdd1.t1484 vp_p.t15 out_p.t580 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X48 vdd1.t1483 vp_p.t16 out_p.t591 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X49 vdd2.t1472 vn_p.t27 out_n.t1734 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X50 vss.t261 vn_n.t3 out_n.t261 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X51 out_p.t581 vp_p.t17 vdd1.t1482 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X52 out_p.t592 vp_p.t18 vdd1.t1481 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X53 out_p.t582 vp_p.t19 vdd1.t1480 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X54 out_n.t49 vn_n.t4 vss.t49 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X55 out_p.t573 vp_p.t20 vdd1.t1479 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X56 out_p.t583 vp_p.t21 vdd1.t1478 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X57 vss.t559 vp_n.t2 out_p.t1779 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X58 vdd1.t1477 vp_p.t22 out_p.t574 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X59 vdd1.t1476 vp_p.t23 out_p.t575 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X60 vdd1.t1475 vp_p.t24 out_p.t565 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X61 vss.t50 vn_n.t5 out_n.t50 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X62 out_n.t1733 vn_p.t28 vdd2.t1471 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X63 out_n.t1732 vn_p.t29 vdd2.t1470 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X64 out_p.t84 vp_n.t3 vss.t558 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X65 out_n.t1731 vn_p.t30 vdd2.t1469 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X66 vdd1.t1474 vp_p.t25 out_p.t566 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X67 out_n.t1730 vn_p.t31 vdd2.t1468 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X68 vdd2.t1467 vn_p.t32 out_n.t1729 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X69 out_p.t567 vp_p.t26 vdd1.t1473 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X70 vdd1.t1472 vp_p.t27 out_p.t556 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X71 out_n.t1728 vn_p.t33 vdd2.t1466 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X72 out_n.t1727 vn_p.t34 vdd2.t1465 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X73 out_n.t1726 vn_p.t35 vdd2.t1464 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X74 vdd2.t1463 vn_p.t36 out_n.t1725 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X75 vdd1.t1471 vp_p.t28 out_p.t568 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X76 vdd1.t1470 vp_p.t29 out_p.t557 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X77 vss.t557 vp_n.t4 out_p.t144 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X78 out_p.t569 vp_p.t30 vdd1.t1469 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X79 vdd2.t1462 vn_p.t37 out_n.t1724 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X80 vss.t556 vp_n.t5 out_p.t145 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X81 vdd2.t1461 vn_p.t38 out_n.t1723 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X82 out_n.t1722 vn_p.t39 vdd2.t1460 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X83 vdd2.t1459 vn_p.t40 out_n.t1721 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X84 vdd1.t1468 vp_p.t31 out_p.t558 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X85 vdd1.t1467 vp_p.t32 out_p.t548 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X86 out_n.t1720 vn_p.t41 vdd2.t1458 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X87 vdd2.t1457 vn_p.t42 out_n.t1719 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X88 vdd2.t1456 vn_p.t43 out_n.t1718 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X89 out_p.t146 vp_n.t6 vss.t555 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X90 out_n.t51 vn_n.t6 vss.t51 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X91 vdd1.t1466 vp_p.t33 out_p.t559 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X92 vdd2.t1455 vn_p.t44 out_n.t1717 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X93 vdd2.t1454 vn_p.t45 out_n.t1716 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X94 out_n.t1715 vn_p.t46 vdd2.t1453 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X95 vss.t554 vp_n.t7 out_p.t147 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X96 out_p.t148 vp_n.t8 vss.t553 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X97 vdd2.t1452 vn_p.t47 out_n.t1714 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X98 out_n.t1713 vn_p.t48 vdd2.t1451 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X99 out_p.t549 vp_p.t34 vdd1.t1465 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X100 vdd1.t1464 vp_p.t35 out_p.t560 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X101 out_p.t550 vp_p.t36 vdd1.t1463 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X102 out_p.t539 vp_p.t37 vdd1.t1462 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X103 out_n.t1712 vn_p.t49 vdd2.t1450 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X104 out_n.t1711 vn_p.t50 vdd2.t1449 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X105 vdd2.t1448 vn_p.t51 out_n.t1710 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X106 vdd1.t1461 vp_p.t38 out_p.t551 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X107 vdd2.t1447 vn_p.t52 out_n.t1709 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X108 vdd1.t1460 vp_p.t39 out_p.t540 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X109 vdd1.t1459 vp_p.t40 out_p.t552 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X110 vdd1.t1458 vp_p.t41 out_p.t541 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X111 out_p.t531 vp_p.t42 vdd1.t1457 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X112 vdd1.t1456 vp_p.t43 out_p.t542 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X113 vss.t52 vn_n.t7 out_n.t52 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X114 vdd2.t1446 vn_p.t53 out_n.t1708 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X115 out_n.t1707 vn_p.t54 vdd2.t1445 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X116 vdd2.t1444 vn_p.t55 out_n.t1706 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X117 out_p.t532 vp_p.t44 vdd1.t1455 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X118 out_n.t1705 vn_p.t56 vdd2.t1443 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X119 out_p.t543 vp_p.t45 vdd1.t1454 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X120 vss.t116 vn_n.t8 out_n.t116 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X121 out_n.t1704 vn_p.t57 vdd2.t1442 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X122 vdd1.t1453 vp_p.t46 out_p.t533 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X123 out_p.t522 vp_p.t47 vdd1.t1452 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X124 out_p.t534 vp_p.t48 vdd1.t1451 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X125 vdd2.t1441 vn_p.t58 out_n.t1703 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X126 out_n.t1702 vn_p.t59 vdd2.t1440 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X127 out_n.t1701 vn_p.t60 vdd2.t1439 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X128 vdd2.t1438 vn_p.t61 out_n.t1700 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X129 out_n.t1699 vn_p.t62 vdd2.t1437 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X130 vdd1.t1450 vp_p.t49 out_p.t523 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X131 out_p.t535 vp_p.t50 vdd1.t1449 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X132 out_n.t1698 vn_p.t63 vdd2.t1436 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X133 vdd1.t1448 vp_p.t51 out_p.t524 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X134 vdd1.t1447 vp_p.t52 out_p.t514 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X135 vdd2.t1435 vn_p.t64 out_n.t1697 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X136 out_p.t525 vp_p.t53 vdd1.t1446 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X137 out_p.t515 vp_p.t54 vdd1.t1445 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X138 out_p.t526 vp_p.t55 vdd1.t1444 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X139 out_n.t1696 vn_p.t65 vdd2.t1434 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X140 vss.t552 vp_n.t9 out_p.t149 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X141 vdd1.t1443 vp_p.t56 out_p.t516 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X142 vdd2.t1433 vn_p.t66 out_n.t1695 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X143 out_p.t505 vp_p.t57 vdd1.t1442 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X144 out_p.t517 vp_p.t58 vdd1.t1441 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X145 out_p.t506 vp_p.t59 vdd1.t1440 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X146 vdd2.t1432 vn_p.t67 out_n.t1694 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X147 out_p.t518 vp_p.t60 vdd1.t1439 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X148 vss.t551 vp_n.t10 out_p.t150 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X149 vdd1.t1438 vp_p.t61 out_p.t507 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X150 vdd1.t1437 vp_p.t62 out_p.t497 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X151 out_p.t151 vp_n.t11 vss.t550 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X152 out_p.t508 vp_p.t63 vdd1.t1436 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X153 out_n.t117 vn_n.t9 vss.t117 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X154 out_n.t1693 vn_p.t68 vdd2.t1431 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X155 vss.t118 vn_n.t10 out_n.t118 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X156 out_n.t1692 vn_p.t69 vdd2.t1430 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X157 vdd2.t1429 vn_p.t70 out_n.t1691 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X158 out_n.t119 vn_n.t11 vss.t119 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X159 out_p.t498 vp_p.t64 vdd1.t1435 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X160 vdd2.t1428 vn_p.t71 out_n.t1690 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X161 out_p.t509 vp_p.t65 vdd1.t1434 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X162 vdd2.t1427 vn_p.t72 out_n.t1689 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X163 vdd1.t1433 vp_p.t66 out_p.t499 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X164 out_n.t1688 vn_p.t73 vdd2.t1426 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X165 vdd2.t1425 vn_p.t74 out_n.t1687 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X166 vdd2.t1424 vn_p.t75 out_n.t1686 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X167 out_n.t1685 vn_p.t76 vdd2.t1423 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X168 vss.t549 vp_n.t12 out_p.t152 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X169 vss.t77 vn_n.t12 out_n.t77 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X170 out_p.t488 vp_p.t67 vdd1.t1432 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X171 out_n.t1684 vn_p.t77 vdd2.t1422 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X172 out_p.t153 vp_n.t13 vss.t548 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X173 out_n.t1683 vn_p.t78 vdd2.t1421 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X174 vdd1.t1431 vp_p.t68 out_p.t500 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X175 vdd2.t1420 vn_p.t79 out_n.t1682 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X176 vdd1.t1430 vp_p.t69 out_p.t489 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X177 vdd1.t1429 vp_p.t70 out_p.t501 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X178 vdd1.t1428 vp_p.t71 out_p.t490 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X179 out_p.t480 vp_p.t72 vdd1.t1427 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X180 vdd1.t1426 vp_p.t73 out_p.t491 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X181 vdd2.t1419 vn_p.t80 out_n.t1681 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X182 vdd2.t1418 vn_p.t81 out_n.t1680 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X183 out_n.t1679 vn_p.t82 vdd2.t1417 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X184 out_p.t481 vp_p.t74 vdd1.t1425 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X185 out_p.t492 vp_p.t75 vdd1.t1424 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X186 vdd1.t1423 vp_p.t76 out_p.t482 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X187 out_p.t471 vp_p.t77 vdd1.t1422 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X188 out_p.t483 vp_p.t78 vdd1.t1421 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X189 out_n.t1678 vn_p.t83 vdd2.t1416 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X190 vdd2.t1415 vn_p.t84 out_n.t1677 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X191 out_n.t1676 vn_p.t85 vdd2.t1414 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X192 vdd1.t1420 vp_p.t79 out_p.t472 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X193 vdd2.t1413 vn_p.t86 out_n.t1675 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X194 out_n.t1674 vn_p.t87 vdd2.t1412 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X195 out_p.t154 vp_n.t14 vss.t547 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X196 vdd1.t1419 vp_p.t80 out_p.t484 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X197 vdd1.t1418 vp_p.t81 out_p.t473 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X198 vdd2.t1411 vn_p.t88 out_n.t1673 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X199 vdd2.t1410 vn_p.t89 out_n.t1672 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X200 vdd1.t1417 vp_p.t82 out_p.t463 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X201 vdd2.t1409 vn_p.t90 out_n.t1671 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X202 vdd2.t1408 vn_p.t91 out_n.t1670 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X203 out_p.t474 vp_p.t83 vdd1.t1416 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X204 out_p.t464 vp_p.t84 vdd1.t1415 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X205 vdd1.t1414 vp_p.t85 out_p.t475 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X206 out_p.t465 vp_p.t86 vdd1.t1413 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X207 out_n.t1669 vn_p.t92 vdd2.t1407 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X208 vdd2.t1406 vn_p.t93 out_n.t1668 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X209 out_p.t454 vp_p.t87 vdd1.t1412 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X210 vdd2.t1405 vn_p.t94 out_n.t1667 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X211 vdd1.t1411 vp_p.t88 out_p.t466 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X212 out_p.t455 vp_p.t89 vdd1.t1410 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X213 vdd1.t1409 vp_p.t90 out_p.t467 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X214 vdd1.t1408 vp_p.t91 out_p.t456 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X215 out_n.t78 vn_n.t13 vss.t78 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X216 vdd2.t1404 vn_p.t95 out_n.t1666 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X217 out_p.t155 vp_n.t15 vss.t546 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X218 out_p.t446 vp_p.t92 vdd1.t1407 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X219 out_n.t1665 vn_p.t96 vdd2.t1403 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X220 vss.t79 vn_n.t14 out_n.t79 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X221 vdd2.t1402 vn_p.t97 out_n.t1664 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X222 out_p.t457 vp_p.t93 vdd1.t1406 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X223 vdd1.t1405 vp_p.t94 out_p.t447 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X224 out_p.t458 vp_p.t95 vdd1.t1404 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X225 vdd2.t1401 vn_p.t98 out_n.t1663 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X226 vss.t545 vp_n.t16 out_p.t156 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X227 out_n.t1662 vn_p.t99 vdd2.t1400 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X228 out_n.t1661 vn_p.t100 vdd2.t1399 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X229 out_n.t1660 vn_p.t101 vdd2.t1398 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X230 vss.t544 vp_n.t17 out_p.t157 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X231 vdd2.t1397 vn_p.t102 out_n.t1659 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X232 out_n.t1658 vn_p.t103 vdd2.t1396 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X233 vss.t80 vn_n.t15 out_n.t80 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X234 out_n.t1657 vn_p.t104 vdd2.t1395 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X235 out_n.t1656 vn_p.t105 vdd2.t1394 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X236 out_p.t448 vp_p.t96 vdd1.t1403 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X237 vdd1.t1402 vp_p.t97 out_p.t437 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X238 vdd1.t1401 vp_p.t98 out_p.t449 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X239 out_n.t1655 vn_p.t106 vdd2.t1393 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X240 out_p.t438 vp_p.t99 vdd1.t1400 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X241 out_n.t1654 vn_p.t107 vdd2.t1392 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X242 out_p.t158 vp_n.t18 vss.t543 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X243 vss.t204 vn_n.t16 out_n.t204 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X244 vss.t542 vp_n.t19 out_p.t159 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X245 vdd1.t1399 vp_p.t100 out_p.t450 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X246 vdd2.t1391 vn_p.t108 out_n.t1653 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X247 out_p.t160 vp_n.t20 vss.t541 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X248 vdd2.t1390 vn_p.t109 out_n.t1652 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X249 vdd2.t1389 vn_p.t110 out_n.t1651 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X250 vdd2.t1388 vn_p.t111 out_n.t1650 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X251 out_n.t1649 vn_p.t112 vdd2.t1387 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X252 out_p.t161 vp_n.t21 vss.t540 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X253 vdd2.t1386 vn_p.t113 out_n.t1648 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X254 out_p.t162 vp_n.t22 vss.t539 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X255 vdd2.t1385 vn_p.t114 out_n.t1647 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X256 out_n.t205 vn_n.t17 vss.t205 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X257 out_p.t439 vp_p.t101 vdd1.t1398 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X258 vdd1.t1397 vp_p.t102 out_p.t429 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X259 out_p.t440 vp_p.t103 vdd1.t1396 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X260 vdd2.t1384 vn_p.t115 out_n.t1646 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X261 vdd1.t1395 vp_p.t104 out_p.t430 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X262 vdd1.t1394 vp_p.t105 out_p.t441 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X263 out_p.t431 vp_p.t106 vdd1.t1393 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X264 out_n.t206 vn_n.t18 vss.t206 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X265 vdd2.t1383 vn_p.t116 out_n.t1645 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X266 vdd1.t1392 vp_p.t107 out_p.t419 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X267 vdd1.t1391 vp_p.t108 out_p.t432 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X268 out_p.t420 vp_p.t109 vdd1.t1390 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X269 vdd1.t1389 vp_p.t110 out_p.t433 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X270 vss.t207 vn_n.t19 out_n.t207 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X271 vdd2.t1382 vn_p.t117 out_n.t1644 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X272 out_p.t421 vp_p.t111 vdd1.t1388 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X273 vdd1.t1387 vp_p.t112 out_p.t409 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X274 vdd1.t1386 vp_p.t113 out_p.t422 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X275 out_p.t410 vp_p.t114 vdd1.t1385 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X276 out_p.t423 vp_p.t115 vdd1.t1384 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X277 out_n.t1643 vn_p.t118 vdd2.t1381 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X278 vdd2.t1380 vn_p.t119 out_n.t1642 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X279 out_n.t1641 vn_p.t120 vdd2.t1379 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X280 out_p.t411 vp_p.t116 vdd1.t1383 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X281 out_n.t1640 vn_p.t121 vdd2.t1378 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X282 vdd2.t1377 vn_p.t122 out_n.t1639 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X283 vss.t538 vp_n.t23 out_p.t163 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X284 out_p.t399 vp_p.t117 vdd1.t1382 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X285 out_n.t1638 vn_p.t123 vdd2.t1376 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X286 vss.t40 vn_n.t20 out_n.t40 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X287 vdd1.t1381 vp_p.t118 out_p.t412 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X288 out_n.t1637 vn_p.t124 vdd2.t1375 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X289 out_p.t400 vp_p.t119 vdd1.t1380 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X290 vdd1.t1379 vp_p.t120 out_p.t413 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X291 out_p.t401 vp_p.t121 vdd1.t1378 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X292 vdd2.t1374 vn_p.t125 out_n.t1636 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X293 vdd2.t1373 vn_p.t126 out_n.t1635 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X294 out_p.t389 vp_p.t122 vdd1.t1377 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X295 out_n.t1634 vn_p.t127 vdd2.t1372 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X296 out_p.t402 vp_p.t123 vdd1.t1376 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X297 vdd2.t1371 vn_p.t128 out_n.t1633 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X298 vdd2.t1370 vn_p.t129 out_n.t1632 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X299 out_n.t1631 vn_p.t130 vdd2.t1369 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X300 vdd1.t1375 vp_p.t124 out_p.t390 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X301 out_n.t1630 vn_p.t131 vdd2.t1368 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X302 vdd1.t1374 vp_p.t125 out_p.t403 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X303 vdd2.t1367 vn_p.t132 out_n.t1629 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X304 out_p.t164 vp_n.t24 vss.t537 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X305 out_n.t1628 vn_p.t133 vdd2.t1366 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X306 vdd2.t1365 vn_p.t134 out_n.t1627 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X307 out_n.t41 vn_n.t21 vss.t41 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X308 vdd2.t1364 vn_p.t135 out_n.t1626 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X309 out_n.t1625 vn_p.t136 vdd2.t1363 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X310 out_p.t391 vp_p.t126 vdd1.t1373 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X311 out_p.t378 vp_p.t127 vdd1.t1372 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X312 out_n.t1624 vn_p.t137 vdd2.t1362 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X313 vdd2.t1361 vn_p.t138 out_n.t1623 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X314 vdd2.t1360 vn_p.t139 out_n.t1622 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X315 vdd1.t1371 vp_p.t128 out_p.t392 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X316 out_p.t379 vp_p.t129 vdd1.t1370 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X317 out_p.t165 vp_n.t25 vss.t536 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X318 out_n.t1621 vn_p.t140 vdd2.t1359 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X319 out_p.t393 vp_p.t130 vdd1.t1369 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X320 out_n.t1620 vn_p.t141 vdd2.t1358 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X321 out_n.t1619 vn_p.t142 vdd2.t1357 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X322 vss.t535 vp_n.t26 out_p.t166 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X323 out_n.t42 vn_n.t22 vss.t42 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X324 out_n.t1618 vn_p.t143 vdd2.t1356 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X325 out_p.t380 vp_p.t131 vdd1.t1368 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X326 vss.t43 vn_n.t23 out_n.t43 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X327 vss.t534 vp_n.t27 out_p.t167 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X328 out_n.t1617 vn_p.t144 vdd2.t1355 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X329 vdd2.t1354 vn_p.t145 out_n.t1616 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X330 vdd1.t1367 vp_p.t132 out_p.t368 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X331 out_n.t1615 vn_p.t146 vdd2.t1353 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X332 vdd1.t1366 vp_p.t133 out_p.t381 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X333 out_p.t369 vp_p.t134 vdd1.t1365 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X334 out_p.t382 vp_p.t135 vdd1.t1364 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X335 out_p.t370 vp_p.t136 vdd1.t1363 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X336 vdd1.t1362 vp_p.t137 out_p.t357 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X337 vss.t533 vp_n.t28 out_p.t168 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X338 out_p.t371 vp_p.t138 vdd1.t1361 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X339 out_p.t358 vp_p.t139 vdd1.t1360 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X340 vss.t170 vn_n.t24 out_n.t170 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X341 out_n.t1614 vn_p.t147 vdd2.t1352 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X342 vdd1.t1359 vp_p.t140 out_p.t372 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X343 vdd1.t1358 vp_p.t141 out_p.t359 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X344 vdd2.t1351 vn_p.t148 out_n.t1613 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X345 vdd1.t1357 vp_p.t142 out_p.t347 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X346 out_p.t360 vp_p.t143 vdd1.t1356 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X347 out_p.t348 vp_p.t144 vdd1.t1355 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X348 out_n.t1612 vn_p.t149 vdd2.t1350 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X349 vdd1.t1354 vp_p.t145 out_p.t361 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X350 out_p.t349 vp_p.t146 vdd1.t1353 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X351 vdd1.t1352 vp_p.t147 out_p.t336 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X352 out_n.t1611 vn_p.t150 vdd2.t1349 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X353 out_p.t169 vp_n.t29 vss.t532 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X354 vdd1.t1351 vp_p.t148 out_p.t350 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X355 out_p.t337 vp_p.t149 vdd1.t1350 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X356 out_n.t171 vn_n.t25 vss.t171 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X357 out_n.t172 vn_n.t26 vss.t172 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X358 vdd2.t1348 vn_p.t151 out_n.t1610 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X359 vss.t173 vn_n.t27 out_n.t173 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X360 out_p.t351 vp_p.t150 vdd1.t1349 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X361 out_p.t338 vp_p.t151 vdd1.t1348 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X362 vdd2.t1347 vn_p.t152 out_n.t1609 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X363 vdd2.t1346 vn_p.t153 out_n.t1608 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X364 vdd2.t1345 vn_p.t154 out_n.t1607 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X365 vdd2.t1344 vn_p.t155 out_n.t1606 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X366 out_n.t1605 vn_p.t156 vdd2.t1343 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X367 vdd2.t1342 vn_p.t157 out_n.t1604 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X368 vdd2.t1341 vn_p.t158 out_n.t1603 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X369 out_n.t36 vn_n.t28 vss.t36 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X370 vdd2.t1340 vn_p.t159 out_n.t1602 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X371 out_n.t1601 vn_p.t160 vdd2.t1339 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X372 vdd1.t1347 vp_p.t152 out_p.t326 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X373 out_p.t956 vp_p.t153 vdd1.t1346 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X374 vss.t531 vp_n.t30 out_p.t170 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X375 out_n.t1600 vn_p.t161 vdd2.t1338 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X376 vdd2.t1337 vn_p.t162 out_n.t1599 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X377 vdd1.t1345 vp_p.t154 out_p.t339 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X378 vdd2.t1336 vn_p.t163 out_n.t1598 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X379 out_n.t1597 vn_p.t164 vdd2.t1335 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X380 out_n.t1596 vn_p.t165 vdd2.t1334 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X381 out_n.t1595 vn_p.t166 vdd2.t1333 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X382 vdd1.t1344 vp_p.t155 out_p.t327 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X383 vdd2.t1332 vn_p.t167 out_n.t1594 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X384 out_p.t340 vp_p.t156 vdd1.t1343 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X385 out_p.t328 vp_p.t157 vdd1.t1342 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X386 vdd1.t1341 vp_p.t158 out_p.t315 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X387 vss.t37 vn_n.t29 out_n.t37 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X388 vdd1.t1340 vp_p.t159 out_p.t329 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X389 out_p.t316 vp_p.t160 vdd1.t1339 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X390 out_n.t1593 vn_p.t168 vdd2.t1331 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X391 vdd2.t1330 vn_p.t169 out_n.t1592 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X392 vdd1.t1338 vp_p.t161 out_p.t330 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X393 out_n.t1591 vn_p.t170 vdd2.t1329 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X394 vdd2.t1328 vn_p.t171 out_n.t1590 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X395 out_n.t1589 vn_p.t172 vdd2.t1327 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X396 out_p.t317 vp_p.t162 vdd1.t1337 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X397 out_n.t1588 vn_p.t173 vdd2.t1326 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X398 vdd2.t1325 vn_p.t174 out_n.t1587 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X399 out_n.t1586 vn_p.t175 vdd2.t1324 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X400 out_p.t305 vp_p.t163 vdd1.t1336 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X401 out_p.t171 vp_n.t31 vss.t530 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X402 vdd2.t1323 vn_p.t176 out_n.t1585 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X403 out_p.t318 vp_p.t164 vdd1.t1335 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X404 vdd1.t1334 vp_p.t165 out_p.t306 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X405 out_p.t319 vp_p.t166 vdd1.t1333 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X406 out_p.t307 vp_p.t167 vdd1.t1332 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X407 vdd1.t1331 vp_p.t168 out_p.t294 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X408 vdd1.t1330 vp_p.t169 out_p.t308 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X409 vdd1.t1329 vp_p.t170 out_p.t295 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X410 out_p.t309 vp_p.t171 vdd1.t1328 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X411 out_n.t1584 vn_p.t177 vdd2.t1322 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X412 out_p.t172 vp_n.t32 vss.t529 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X413 out_n.t38 vn_n.t30 vss.t38 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X414 vss.t39 vn_n.t31 out_n.t39 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X415 vdd2.t1321 vn_p.t178 out_n.t1583 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X416 out_n.t140 vn_n.t32 vss.t140 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X417 vdd2.t1320 vn_p.t179 out_n.t1582 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X418 out_p.t296 vp_p.t172 vdd1.t1327 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X419 out_p.t285 vp_p.t173 vdd1.t1326 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X420 out_p.t957 vp_p.t174 vdd1.t1325 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X421 vss.t528 vp_n.t33 out_p.t173 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X422 vdd1.t1324 vp_p.t175 out_p.t286 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X423 out_p.t287 vp_p.t176 vdd1.t1323 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X424 out_p.t276 vp_p.t177 vdd1.t1322 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X425 out_p.t174 vp_n.t34 vss.t527 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X426 out_p.t288 vp_p.t178 vdd1.t1321 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X427 out_n.t1581 vn_p.t180 vdd2.t1319 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X428 vdd2.t1318 vn_p.t181 out_n.t1580 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X429 vdd2.t1317 vn_p.t182 out_n.t1579 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X430 out_n.t1578 vn_p.t183 vdd2.t1316 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X431 vdd2.t1315 vn_p.t184 out_n.t1577 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X432 vdd1.t1320 vp_p.t179 out_p.t277 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X433 out_n.t1576 vn_p.t185 vdd2.t1314 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X434 out_n.t1575 vn_p.t186 vdd2.t1313 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X435 vdd2.t1312 vn_p.t187 out_n.t1574 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X436 out_p.t278 vp_p.t180 vdd1.t1319 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X437 out_n.t1573 vn_p.t188 vdd2.t1311 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X438 out_p.t175 vp_n.t35 vss.t526 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X439 vdd2.t1310 vn_p.t189 out_n.t1572 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X440 vdd2.t1309 vn_p.t190 out_n.t1571 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X441 vss.t141 vn_n.t33 out_n.t141 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X442 out_n.t1570 vn_p.t191 vdd2.t1308 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X443 vss.t142 vn_n.t34 out_n.t142 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X444 vdd2.t1307 vn_p.t192 out_n.t1569 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X445 out_p.t176 vp_n.t36 vss.t525 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X446 out_n.t1568 vn_p.t193 vdd2.t1306 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X447 out_n.t1567 vn_p.t194 vdd2.t1305 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X448 out_n.t1566 vn_p.t195 vdd2.t1304 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X449 out_p.t279 vp_p.t181 vdd1.t1318 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X450 vdd2.t1303 vn_p.t196 out_n.t1565 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X451 out_n.t1564 vn_p.t197 vdd2.t1302 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X452 out_n.t1563 vn_p.t198 vdd2.t1301 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X453 vdd1.t1317 vp_p.t182 out_p.t925 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X454 out_n.t143 vn_n.t35 vss.t143 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X455 vdd2.t1300 vn_p.t199 out_n.t1562 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X456 vdd1.t1316 vp_p.t183 out_p.t926 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X457 out_p.t927 vp_p.t184 vdd1.t1315 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X458 vdd1.t1314 vp_p.t185 out_p.t915 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X459 out_n.t125 vn_n.t36 vss.t125 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X460 out_p.t931 vp_p.t186 vdd1.t1313 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X461 out_p.t916 vp_p.t187 vdd1.t1312 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X462 out_p.t917 vp_p.t188 vdd1.t1311 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X463 vdd1.t1310 vp_p.t189 out_p.t932 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X464 vdd2.t1299 vn_p.t200 out_n.t1561 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X465 out_n.t1560 vn_p.t201 vdd2.t1298 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X466 out_p.t905 vp_p.t190 vdd1.t1309 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X467 out_p.t921 vp_p.t191 vdd1.t1308 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X468 vdd1.t1307 vp_p.t192 out_p.t906 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X469 vdd2.t1297 vn_p.t202 out_n.t1559 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X470 vdd1.t1306 vp_p.t193 out_p.t907 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X471 vdd1.t1305 vp_p.t194 out_p.t922 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X472 out_n.t126 vn_n.t37 vss.t126 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X473 vss.t127 vn_n.t38 out_n.t127 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X474 out_n.t1558 vn_p.t203 vdd2.t1296 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X475 vdd1.t1304 vp_p.t195 out_p.t895 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X476 vdd2.t1295 vn_p.t204 out_n.t1557 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X477 out_n.t1556 vn_p.t205 vdd2.t1294 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X478 out_p.t911 vp_p.t196 vdd1.t1303 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X479 vdd1.t1302 vp_p.t197 out_p.t896 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X480 out_p.t897 vp_p.t198 vdd1.t1301 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X481 vdd2.t1293 vn_p.t206 out_n.t1555 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X482 out_p.t912 vp_p.t199 vdd1.t1300 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X483 out_p.t885 vp_p.t200 vdd1.t1299 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X484 out_p.t901 vp_p.t201 vdd1.t1298 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X485 vdd1.t1297 vp_p.t202 out_p.t886 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X486 out_n.t1554 vn_p.t207 vdd2.t1292 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X487 vss.t128 vn_n.t39 out_n.t128 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X488 vss.t524 vp_n.t37 out_p.t177 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X489 vdd1.t1296 vp_p.t203 out_p.t887 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X490 vdd1.t1295 vp_p.t204 out_p.t902 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X491 out_n.t1553 vn_p.t208 vdd2.t1291 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X492 vdd1.t1294 vp_p.t205 out_p.t875 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X493 out_p.t891 vp_p.t206 vdd1.t1293 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X494 out_n.t1552 vn_p.t209 vdd2.t1290 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X495 out_n.t1551 vn_p.t210 vdd2.t1289 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X496 out_p.t178 vp_n.t38 vss.t523 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X497 vdd1.t1292 vp_p.t207 out_p.t876 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X498 out_n.t1550 vn_p.t211 vdd2.t1288 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X499 vdd1.t1291 vp_p.t208 out_p.t877 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X500 out_n.t1549 vn_p.t212 vdd2.t1287 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X501 out_p.t892 vp_p.t209 vdd1.t1290 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X502 vdd1.t1289 vp_p.t210 out_p.t865 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X503 out_n.t1548 vn_p.t213 vdd2.t1286 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X504 vdd2.t1285 vn_p.t214 out_n.t1547 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X505 out_n.t1546 vn_p.t215 vdd2.t1284 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X506 out_n.t1545 vn_p.t216 vdd2.t1283 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X507 vdd1.t1288 vp_p.t211 out_p.t881 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X508 vdd2.t1282 vn_p.t217 out_n.t1544 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X509 vss.t596 vn_n.t40 out_n.t1796 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X510 out_n.t1797 vn_n.t41 vss.t597 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X511 out_n.t1543 vn_p.t218 vdd2.t1281 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X512 out_p.t179 vp_n.t39 vss.t522 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X513 vdd2.t1280 vn_p.t219 out_n.t1542 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X514 vdd2.t1279 vn_p.t220 out_n.t1541 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X515 out_n.t1540 vn_p.t221 vdd2.t1278 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X516 vdd2.t1277 vn_p.t222 out_n.t1539 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X517 vdd2.t1276 vn_p.t223 out_n.t1538 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X518 vss.t598 vn_n.t42 out_n.t1798 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X519 out_n.t1799 vn_n.t43 vss.t599 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X520 vdd2.t1275 vn_p.t224 out_n.t1537 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X521 vss.t521 vp_n.t40 out_p.t180 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X522 vdd2.t1274 vn_p.t225 out_n.t1536 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X523 out_p.t866 vp_p.t212 vdd1.t1287 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X524 out_p.t867 vp_p.t213 vdd1.t1286 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X525 vdd1.t1285 vp_p.t214 out_p.t882 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X526 vdd2.t1273 vn_p.t226 out_n.t1535 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X527 out_p.t855 vp_p.t215 vdd1.t1284 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X528 out_p.t871 vp_p.t216 vdd1.t1283 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X529 vdd1.t1282 vp_p.t217 out_p.t856 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X530 vdd1.t1281 vp_p.t218 out_p.t857 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X531 out_p.t872 vp_p.t219 vdd1.t1280 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X532 out_n.t185 vn_n.t44 vss.t185 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X533 vdd1.t1279 vp_p.t220 out_p.t845 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X534 out_n.t1534 vn_p.t227 vdd2.t1272 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X535 out_n.t1533 vn_p.t228 vdd2.t1271 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X536 vdd1.t1278 vp_p.t221 out_p.t861 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X537 vdd1.t1277 vp_p.t222 out_p.t846 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X538 out_p.t847 vp_p.t223 vdd1.t1276 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X539 out_n.t1532 vn_p.t229 vdd2.t1270 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X540 out_n.t1531 vn_p.t230 vdd2.t1269 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X541 out_p.t862 vp_p.t224 vdd1.t1275 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X542 vdd1.t1274 vp_p.t225 out_p.t835 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X543 vdd2.t1268 vn_p.t231 out_n.t1530 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X544 out_n.t1529 vn_p.t232 vdd2.t1267 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X545 out_p.t851 vp_p.t226 vdd1.t1273 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X546 vss.t186 vn_n.t45 out_n.t186 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X547 out_p.t836 vp_p.t227 vdd1.t1272 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X548 out_p.t837 vp_p.t228 vdd1.t1271 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X549 out_p.t852 vp_p.t229 vdd1.t1270 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X550 out_p.t825 vp_p.t230 vdd1.t1269 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X551 vss.t187 vn_n.t46 out_n.t187 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X552 out_n.t1528 vn_p.t233 vdd2.t1266 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X553 out_n.t1527 vn_p.t234 vdd2.t1265 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X554 vdd1.t1268 vp_p.t231 out_p.t841 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X555 vdd1.t1267 vp_p.t232 out_p.t826 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X556 vdd2.t1264 vn_p.t235 out_n.t1526 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X557 vdd1.t1266 vp_p.t233 out_p.t827 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X558 out_n.t1525 vn_p.t236 vdd2.t1263 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X559 out_p.t181 vp_n.t41 vss.t520 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X560 vdd1.t1265 vp_p.t234 out_p.t842 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X561 out_p.t815 vp_p.t235 vdd1.t1264 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X562 out_p.t831 vp_p.t236 vdd1.t1263 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X563 vdd2.t1262 vn_p.t237 out_n.t1524 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X564 out_n.t1523 vn_p.t238 vdd2.t1261 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X565 out_n.t1522 vn_p.t239 vdd2.t1260 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X566 vdd2.t1259 vn_p.t240 out_n.t1521 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X567 vss.t519 vp_n.t42 out_p.t182 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X568 vdd1.t1262 vp_p.t237 out_p.t816 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X569 vdd2.t1258 vn_p.t241 out_n.t1520 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X570 out_p.t183 vp_n.t43 vss.t518 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X571 vdd1.t1261 vp_p.t238 out_p.t817 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X572 vdd2.t1257 vn_p.t242 out_n.t1519 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X573 out_p.t832 vp_p.t239 vdd1.t1260 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X574 out_p.t805 vp_p.t240 vdd1.t1259 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X575 out_n.t188 vn_n.t47 vss.t188 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X576 out_p.t184 vp_n.t44 vss.t517 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X577 vdd1.t1258 vp_p.t241 out_p.t821 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X578 vdd2.t1256 vn_p.t243 out_n.t1518 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X579 out_p.t185 vp_n.t45 vss.t516 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X580 out_n.t1517 vn_p.t244 vdd2.t1255 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X581 out_n.t13 vn_n.t48 vss.t13 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X582 vss.t14 vn_n.t49 out_n.t14 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X583 out_p.t186 vp_n.t46 vss.t515 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X584 vdd2.t1254 vn_p.t245 out_n.t1516 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X585 out_p.t806 vp_p.t242 vdd1.t1257 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X586 out_n.t15 vn_n.t50 vss.t15 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X587 vss.t16 vn_n.t51 out_n.t16 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X588 vdd2.t1253 vn_p.t246 out_n.t1515 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X589 vss.t514 vp_n.t47 out_p.t187 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X590 vss.t513 vp_n.t48 out_p.t188 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X591 out_n.t1514 vn_p.t247 vdd2.t1252 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X592 vdd2.t1251 vn_p.t248 out_n.t1513 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X593 out_p.t807 vp_p.t243 vdd1.t1256 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X594 out_n.t1512 vn_p.t249 vdd2.t1250 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X595 vss.t238 vn_n.t52 out_n.t238 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X596 vss.t512 vp_n.t49 out_p.t189 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X597 vss.t239 vn_n.t53 out_n.t239 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X598 vdd2.t1249 vn_p.t250 out_n.t1511 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X599 out_p.t822 vp_p.t244 vdd1.t1255 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X600 out_p.t795 vp_p.t245 vdd1.t1254 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X601 vdd1.t1253 vp_p.t246 out_p.t811 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X602 out_n.t1510 vn_p.t251 vdd2.t1248 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X603 out_p.t796 vp_p.t247 vdd1.t1252 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X604 out_p.t797 vp_p.t248 vdd1.t1251 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X605 vdd1.t1250 vp_p.t249 out_p.t812 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X606 vdd1.t1249 vp_p.t250 out_p.t785 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X607 out_p.t801 vp_p.t251 vdd1.t1248 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X608 vdd2.t1247 vn_p.t252 out_n.t1509 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X609 vdd2.t1246 vn_p.t253 out_n.t1508 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X610 out_n.t1507 vn_p.t254 vdd2.t1245 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X611 out_p.t786 vp_p.t252 vdd1.t1247 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X612 vdd1.t1246 vp_p.t253 out_p.t787 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X613 out_p.t802 vp_p.t254 vdd1.t1245 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X614 out_p.t775 vp_p.t255 vdd1.t1244 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X615 out_n.t240 vn_n.t54 vss.t240 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X616 vss.t241 vn_n.t55 out_n.t241 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X617 vdd2.t1244 vn_p.t255 out_n.t1506 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X618 vdd2.t1243 vn_p.t256 out_n.t1505 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X619 out_n.t155 vn_n.t56 vss.t155 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X620 out_p.t791 vp_p.t256 vdd1.t1243 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X621 vdd1.t1242 vp_p.t257 out_p.t776 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X622 vdd2.t1242 vn_p.t257 out_n.t1504 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X623 out_n.t1503 vn_p.t258 vdd2.t1241 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X624 out_p.t777 vp_p.t258 vdd1.t1241 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X625 vdd2.t1240 vn_p.t259 out_n.t1502 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X626 vdd1.t1240 vp_p.t259 out_p.t792 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X627 vdd1.t1239 vp_p.t260 out_p.t765 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X628 vdd2.t1239 vn_p.t260 out_n.t1501 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X629 out_p.t781 vp_p.t261 vdd1.t1238 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X630 vdd2.t1238 vn_p.t261 out_n.t1500 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X631 out_p.t766 vp_p.t262 vdd1.t1237 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X632 out_p.t767 vp_p.t263 vdd1.t1236 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X633 out_p.t782 vp_p.t264 vdd1.t1235 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X634 vdd1.t1234 vp_p.t265 out_p.t755 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X635 vdd1.t1233 vp_p.t266 out_p.t771 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X636 vdd2.t1237 vn_p.t262 out_n.t1499 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X637 out_p.t190 vp_n.t50 vss.t511 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X638 out_p.t756 vp_p.t267 vdd1.t1232 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X639 vss.t510 vp_n.t51 out_p.t191 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X640 vdd1.t1231 vp_p.t268 out_p.t757 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X641 vss.t156 vn_n.t57 out_n.t156 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X642 out_n.t1498 vn_p.t263 vdd2.t1236 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X643 vdd1.t1230 vp_p.t269 out_p.t772 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X644 out_n.t157 vn_n.t58 vss.t157 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X645 out_p.t745 vp_p.t270 vdd1.t1229 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X646 out_p.t761 vp_p.t271 vdd1.t1228 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X647 vss.t509 vp_n.t52 out_p.t192 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X648 vdd1.t1227 vp_p.t272 out_p.t746 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X649 out_n.t1497 vn_p.t264 vdd2.t1235 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X650 out_n.t1496 vn_p.t265 vdd2.t1234 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X651 vdd2.t1233 vn_p.t266 out_n.t1495 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X652 vdd2.t1232 vn_p.t267 out_n.t1494 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X653 out_n.t1493 vn_p.t268 vdd2.t1231 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X654 out_p.t193 vp_n.t53 vss.t508 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X655 out_n.t1492 vn_p.t269 vdd2.t1230 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X656 vdd1.t1226 vp_p.t273 out_p.t747 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X657 vss.t158 vn_n.t59 out_n.t158 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X658 out_n.t1491 vn_p.t270 vdd2.t1229 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X659 vdd1.t1225 vp_p.t274 out_p.t762 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X660 out_p.t735 vp_p.t275 vdd1.t1224 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X661 out_p.t194 vp_n.t54 vss.t507 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X662 vdd1.t1223 vp_p.t276 out_p.t751 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X663 out_p.t195 vp_n.t55 vss.t506 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X664 vdd2.t1228 vn_p.t271 out_n.t1490 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X665 out_n.t1489 vn_p.t272 vdd2.t1227 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X666 vdd1.t1222 vp_p.t277 out_p.t736 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X667 out_n.t1488 vn_p.t273 vdd2.t1226 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X668 vdd2.t1225 vn_p.t274 out_n.t1487 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X669 vdd1.t1221 vp_p.t278 out_p.t737 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X670 vdd2.t1224 vn_p.t275 out_n.t1486 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X671 vdd2.t1223 vn_p.t276 out_n.t1485 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X672 out_p.t752 vp_p.t279 vdd1.t1220 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X673 out_n.t233 vn_n.t60 vss.t233 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X674 vdd2.t1222 vn_p.t277 out_n.t1484 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X675 out_p.t725 vp_p.t280 vdd1.t1219 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X676 out_p.t741 vp_p.t281 vdd1.t1218 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X677 out_p.t726 vp_p.t282 vdd1.t1217 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X678 vdd1.t1216 vp_p.t283 out_p.t727 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X679 out_p.t742 vp_p.t284 vdd1.t1215 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X680 out_n.t1483 vn_p.t278 vdd2.t1221 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X681 vdd1.t1214 vp_p.t285 out_p.t715 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X682 vdd1.t1213 vp_p.t286 out_p.t731 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X683 vdd2.t1220 vn_p.t279 out_n.t1482 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X684 out_p.t716 vp_p.t287 vdd1.t1212 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X685 vdd1.t1211 vp_p.t288 out_p.t717 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X686 out_p.t732 vp_p.t289 vdd1.t1210 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X687 out_n.t1481 vn_p.t280 vdd2.t1219 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X688 vdd2.t1218 vn_p.t281 out_n.t1480 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X689 vdd1.t1209 vp_p.t290 out_p.t705 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X690 vss.t234 vn_n.t61 out_n.t234 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X691 out_n.t235 vn_n.t62 vss.t235 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X692 out_p.t721 vp_p.t291 vdd1.t1208 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X693 vss.t505 vp_n.t56 out_p.t196 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X694 vdd1.t1207 vp_p.t292 out_p.t706 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X695 out_n.t1479 vn_p.t282 vdd2.t1217 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X696 vdd2.t1216 vn_p.t283 out_n.t1478 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X697 out_n.t1477 vn_p.t284 vdd2.t1215 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X698 out_n.t1476 vn_p.t285 vdd2.t1214 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X699 vdd2.t1213 vn_p.t286 out_n.t1475 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X700 vdd1.t1206 vp_p.t293 out_p.t707 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X701 vdd1.t1205 vp_p.t294 out_p.t722 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X702 out_p.t694 vp_p.t295 vdd1.t1204 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X703 vdd1.t1203 vp_p.t296 out_p.t711 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X704 vdd1.t1202 vp_p.t297 out_p.t695 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X705 vss.t236 vn_n.t63 out_n.t236 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X706 out_p.t696 vp_p.t298 vdd1.t1201 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X707 vss.t237 vn_n.t64 out_n.t237 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X708 vdd1.t1200 vp_p.t299 out_p.t712 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X709 vdd1.t1199 vp_p.t300 out_p.t683 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X710 out_n.t1474 vn_p.t287 vdd2.t1212 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X711 out_p.t700 vp_p.t301 vdd1.t1198 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X712 out_n.t1473 vn_p.t288 vdd2.t1211 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X713 vdd2.t1210 vn_p.t289 out_n.t1472 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X714 vdd2.t1209 vn_p.t290 out_n.t1471 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X715 out_n.t1470 vn_p.t291 vdd2.t1208 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X716 out_n.t1469 vn_p.t292 vdd2.t1207 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X717 vdd2.t1206 vn_p.t293 out_n.t1468 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X718 vdd2.t1205 vn_p.t294 out_n.t1467 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X719 out_n.t1466 vn_p.t295 vdd2.t1204 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X720 out_p.t125 vp_n.t57 vss.t504 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X721 out_n.t218 vn_n.t65 vss.t218 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X722 out_p.t684 vp_p.t302 vdd1.t1197 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X723 vdd2.t1203 vn_p.t296 out_n.t1465 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X724 out_n.t1464 vn_p.t297 vdd2.t1202 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X725 vdd1.t1196 vp_p.t303 out_p.t685 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X726 out_p.t701 vp_p.t304 vdd1.t1195 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X727 vdd1.t1194 vp_p.t305 out_p.t673 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X728 vdd1.t1193 vp_p.t306 out_p.t689 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X729 out_n.t1463 vn_p.t298 vdd2.t1201 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X730 out_n.t1462 vn_p.t299 vdd2.t1200 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X731 vdd2.t1199 vn_p.t300 out_n.t1461 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X732 vss.t503 vp_n.t58 out_p.t126 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X733 out_p.t127 vp_n.t59 vss.t502 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X734 vss.t501 vp_n.t60 out_p.t128 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X735 vdd2.t1198 vn_p.t301 out_n.t1460 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X736 vdd2.t1197 vn_p.t302 out_n.t1459 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X737 out_p.t674 vp_p.t307 vdd1.t1192 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X738 vdd2.t1196 vn_p.t303 out_n.t1458 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X739 out_n.t1457 vn_p.t304 vdd2.t1195 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X740 vss.t219 vn_n.t66 out_n.t219 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X741 vdd1.t1191 vp_p.t308 out_p.t675 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X742 out_p.t690 vp_p.t309 vdd1.t1190 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X743 vdd1.t1189 vp_p.t310 out_p.t663 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X744 vdd1.t1188 vp_p.t311 out_p.t678 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X745 vdd1.t1187 vp_p.t312 out_p.t664 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X746 out_n.t1456 vn_p.t305 vdd2.t1194 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X747 vdd1.t1186 vp_p.t313 out_p.t665 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X748 out_p.t679 vp_p.t314 vdd1.t1185 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X749 vdd1.t1184 vp_p.t315 out_p.t651 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X750 out_n.t1455 vn_p.t306 vdd2.t1193 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X751 vdd2.t1192 vn_p.t307 out_n.t1454 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X752 out_n.t1453 vn_p.t308 vdd2.t1191 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X753 out_p.t129 vp_n.t61 vss.t500 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X754 out_p.t668 vp_p.t316 vdd1.t1183 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X755 out_p.t652 vp_p.t317 vdd1.t1182 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X756 out_p.t653 vp_p.t318 vdd1.t1181 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X757 vdd1.t1180 vp_p.t319 out_p.t669 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X758 out_p.t640 vp_p.t320 vdd1.t1179 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X759 vdd2.t1190 vn_p.t309 out_n.t1452 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X760 out_n.t1451 vn_p.t310 vdd2.t1189 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X761 out_n.t1450 vn_p.t311 vdd2.t1188 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X762 vdd1.t1178 vp_p.t321 out_p.t657 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X763 out_p.t641 vp_p.t322 vdd1.t1177 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X764 out_n.t1449 vn_p.t312 vdd2.t1187 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X765 vdd1.t1176 vp_p.t323 out_p.t642 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X766 out_n.t1448 vn_p.t313 vdd2.t1186 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X767 vdd1.t1175 vp_p.t324 out_p.t658 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X768 vdd2.t1185 vn_p.t314 out_n.t1447 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X769 vdd2.t1184 vn_p.t315 out_n.t1446 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X770 out_p.t130 vp_n.t62 vss.t499 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X771 vdd1.t1174 vp_p.t325 out_p.t628 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X772 vdd1.t1173 vp_p.t326 out_p.t646 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X773 out_n.t1445 vn_p.t316 vdd2.t1183 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X774 out_p.t629 vp_p.t327 vdd1.t1172 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X775 out_p.t630 vp_p.t328 vdd1.t1171 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X776 vdd2.t1182 vn_p.t317 out_n.t1444 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X777 out_n.t220 vn_n.t67 vss.t220 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X778 out_n.t1443 vn_p.t318 vdd2.t1181 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X779 out_n.t1442 vn_p.t319 vdd2.t1180 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X780 vdd2.t1179 vn_p.t320 out_n.t1441 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X781 vdd1.t1170 vp_p.t329 out_p.t648 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X782 out_p.t616 vp_p.t330 vdd1.t1169 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X783 vdd2.t1178 vn_p.t321 out_n.t1440 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X784 vdd1.t1168 vp_p.t331 out_p.t633 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X785 vdd1.t1167 vp_p.t332 out_p.t634 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X786 vss.t498 vp_n.t63 out_p.t131 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X787 vdd2.t1177 vn_p.t322 out_n.t1439 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X788 vdd1.t1166 vp_p.t333 out_p.t617 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X789 vdd2.t1176 vn_p.t323 out_n.t1438 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X790 vdd2.t1175 vn_p.t324 out_n.t1437 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X791 vdd2.t1174 vn_p.t325 out_n.t1436 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X792 out_n.t221 vn_n.t68 vss.t221 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X793 out_n.t1435 vn_p.t326 vdd2.t1173 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X794 vdd2.t1172 vn_p.t327 out_n.t1434 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X795 out_p.t649 vp_p.t334 vdd1.t1165 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X796 vss.t222 vn_n.t69 out_n.t222 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X797 out_n.t1433 vn_p.t328 vdd2.t1171 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X798 vdd2.t1170 vn_p.t329 out_n.t1432 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X799 vdd1.t1164 vp_p.t335 out_p.t618 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X800 out_n.t1431 vn_p.t330 vdd2.t1169 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X801 out_p.t619 vp_p.t336 vdd1.t1163 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X802 vdd1.t1162 vp_p.t337 out_p.t635 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X803 vdd1.t1161 vp_p.t338 out_p.t621 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X804 out_n.t1430 vn_p.t331 vdd2.t1168 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X805 out_p.t622 vp_p.t339 vdd1.t1160 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X806 out_n.t1429 vn_p.t332 vdd2.t1167 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X807 out_n.t1428 vn_p.t333 vdd2.t1166 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X808 vdd2.t1165 vn_p.t334 out_n.t1427 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X809 vdd1.t1159 vp_p.t340 out_p.t636 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X810 out_p.t623 vp_p.t341 vdd1.t1158 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X811 out_n.t1426 vn_p.t335 vdd2.t1164 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X812 vss.t497 vp_n.t64 out_p.t132 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X813 vss.t72 vn_n.t70 out_n.t72 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X814 out_p.t133 vp_n.t65 vss.t496 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X815 out_p.t624 vp_p.t342 vdd1.t1157 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X816 out_n.t1425 vn_p.t336 vdd2.t1163 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X817 vdd1.t1156 vp_p.t343 out_p.t942 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X818 vdd2.t1162 vn_p.t337 out_n.t1424 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X819 out_n.t1423 vn_p.t338 vdd2.t1161 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X820 out_p.t943 vp_p.t344 vdd1.t1155 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X821 vdd2.t1160 vn_p.t339 out_n.t1422 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X822 vdd1.t1154 vp_p.t345 out_p.t944 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X823 out_p.t945 vp_p.t346 vdd1.t1153 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X824 vdd2.t1159 vn_p.t340 out_n.t1421 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X825 out_p.t947 vp_p.t347 vdd1.t1152 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X826 vdd1.t1151 vp_p.t348 out_p.t948 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X827 out_p.t949 vp_p.t349 vdd1.t1150 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X828 vdd2.t1158 vn_p.t341 out_n.t1420 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X829 vdd2.t1157 vn_p.t342 out_n.t1419 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X830 vdd1.t1149 vp_p.t350 out_p.t267 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X831 vdd1.t1148 vp_p.t351 out_p.t1027 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X832 out_p.t638 vp_p.t352 vdd1.t1147 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X833 vdd1.t1146 vp_p.t353 out_p.t1091 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X834 out_p.t134 vp_n.t66 vss.t495 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X835 out_p.t1086 vp_p.t354 vdd1.t1145 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X836 out_p.t1082 vp_p.t355 vdd1.t1144 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X837 vdd1.t1143 vp_p.t356 out_p.t1088 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X838 vdd2.t1156 vn_p.t343 out_n.t1418 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X839 out_n.t73 vn_n.t71 vss.t73 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X840 out_n.t74 vn_n.t72 vss.t74 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X841 vdd1.t1142 vp_p.t357 out_p.t1085 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X842 vss.t75 vn_n.t73 out_n.t75 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X843 vdd2.t1155 vn_p.t344 out_n.t1417 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X844 vss.t494 vp_n.t67 out_p.t135 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X845 out_p.t1093 vp_p.t358 vdd1.t1141 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X846 out_p.t1092 vp_p.t359 vdd1.t1140 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X847 vdd2.t1154 vn_p.t345 out_n.t1416 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X848 out_n.t1415 vn_p.t346 vdd2.t1153 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X849 out_n.t1414 vn_p.t347 vdd2.t1152 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X850 vdd2.t1151 vn_p.t348 out_n.t1413 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X851 vdd1.t1139 vp_p.t360 out_p.t1089 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X852 vdd2.t1150 vn_p.t349 out_n.t1412 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X853 out_n.t1411 vn_p.t350 vdd2.t1149 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X854 out_n.t1410 vn_p.t351 vdd2.t1148 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X855 vdd2.t1147 vn_p.t352 out_n.t1409 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X856 out_n.t1408 vn_p.t353 vdd2.t1146 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X857 out_p.t1081 vp_p.t361 vdd1.t1138 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X858 out_n.t1407 vn_p.t354 vdd2.t1145 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X859 out_n.t1406 vn_p.t355 vdd2.t1144 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X860 vdd1.t1137 vp_p.t362 out_p.t1080 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X861 out_p.t136 vp_n.t68 vss.t493 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X862 vdd2.t1143 vn_p.t356 out_n.t1405 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X863 vdd2.t1142 vn_p.t357 out_n.t1404 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X864 out_n.t1403 vn_p.t358 vdd2.t1141 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X865 vdd2.t1140 vn_p.t359 out_n.t1402 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X866 out_n.t1401 vn_p.t360 vdd2.t1139 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X867 out_p.t1079 vp_p.t363 vdd1.t1136 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X868 out_n.t1400 vn_p.t361 vdd2.t1138 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X869 vdd2.t1137 vn_p.t362 out_n.t1399 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X870 vdd1.t1135 vp_p.t364 out_p.t1078 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X871 out_p.t1077 vp_p.t365 vdd1.t1134 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X872 vdd1.t1133 vp_p.t366 out_p.t1076 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X873 vdd1.t1132 vp_p.t367 out_p.t1075 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X874 out_n.t1398 vn_p.t363 vdd2.t1136 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X875 out_p.t1074 vp_p.t368 vdd1.t1131 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X876 out_p.t1073 vp_p.t369 vdd1.t1130 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X877 vdd1.t1129 vp_p.t370 out_p.t1072 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X878 vdd2.t1135 vn_p.t364 out_n.t1397 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X879 out_n.t76 vn_n.t74 vss.t76 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X880 out_p.t1068 vp_p.t371 vdd1.t1128 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X881 out_n.t159 vn_n.t75 vss.t159 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X882 vdd2.t1134 vn_p.t365 out_n.t1396 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X883 vdd1.t1127 vp_p.t372 out_p.t1071 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X884 out_n.t1395 vn_p.t366 vdd2.t1133 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X885 out_p.t1070 vp_p.t373 vdd1.t1126 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X886 vdd2.t1132 vn_p.t367 out_n.t1394 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X887 out_p.t1069 vp_p.t374 vdd1.t1125 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X888 vdd1.t1124 vp_p.t375 out_p.t1067 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X889 vdd2.t1131 vn_p.t368 out_n.t1393 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X890 out_p.t1066 vp_p.t376 vdd1.t1123 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X891 vss.t492 vp_n.t69 out_p.t137 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X892 vdd1.t1122 vp_p.t377 out_p.t1065 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X893 out_p.t138 vp_n.t70 vss.t491 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X894 vdd1.t1121 vp_p.t378 out_p.t1064 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X895 vdd1.t1120 vp_p.t379 out_p.t1063 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X896 vss.t160 vn_n.t76 out_n.t160 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X897 out_n.t161 vn_n.t77 vss.t161 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X898 vdd2.t1130 vn_p.t369 out_n.t1392 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X899 out_p.t1062 vp_p.t380 vdd1.t1119 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X900 vdd1.t1118 vp_p.t381 out_p.t1061 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X901 out_p.t1060 vp_p.t382 vdd1.t1117 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X902 out_p.t1059 vp_p.t383 vdd1.t1116 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X903 out_p.t1058 vp_p.t384 vdd1.t1115 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X904 vdd1.t1114 vp_p.t385 out_p.t1057 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X905 vdd2.t1129 vn_p.t370 out_n.t1391 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X906 vss.t490 vp_n.t71 out_p.t139 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X907 vss.t489 vp_n.t72 out_p.t140 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X908 vss.t162 vn_n.t78 out_n.t162 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X909 out_p.t1056 vp_p.t386 vdd1.t1113 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X910 out_n.t1390 vn_p.t371 vdd2.t1128 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X911 vdd1.t1112 vp_p.t387 out_p.t1055 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X912 out_n.t1389 vn_p.t372 vdd2.t1127 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X913 vdd2.t1126 vn_p.t373 out_n.t1388 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X914 vss.t163 vn_n.t79 out_n.t163 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X915 out_n.t1387 vn_p.t374 vdd2.t1125 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X916 out_p.t1054 vp_p.t388 vdd1.t1111 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X917 vdd1.t1110 vp_p.t389 out_p.t1053 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X918 out_n.t1386 vn_p.t375 vdd2.t1124 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X919 vdd2.t1123 vn_p.t376 out_n.t1385 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X920 vss.t488 vp_n.t73 out_p.t141 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X921 vdd1.t1109 vp_p.t390 out_p.t1052 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X922 out_n.t1384 vn_p.t377 vdd2.t1122 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X923 out_p.t1051 vp_p.t391 vdd1.t1108 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X924 out_n.t1383 vn_p.t378 vdd2.t1121 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X925 vdd2.t1120 vn_p.t379 out_n.t1382 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X926 out_n.t1381 vn_p.t380 vdd2.t1119 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X927 out_n.t1380 vn_p.t381 vdd2.t1118 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X928 vdd1.t1107 vp_p.t392 out_p.t1050 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X929 vdd2.t1117 vn_p.t382 out_n.t1379 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X930 vdd2.t1116 vn_p.t383 out_n.t1378 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X931 vss.t487 vp_n.t74 out_p.t142 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X932 out_n.t228 vn_n.t80 vss.t228 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X933 vdd2.t1115 vn_p.t384 out_n.t1377 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X934 out_p.t143 vp_n.t75 vss.t486 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X935 vdd2.t1114 vn_p.t385 out_n.t1376 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X936 vss.t485 vp_n.t76 out_p.t0 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X937 vdd2.t1113 vn_p.t386 out_n.t1375 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X938 out_n.t1374 vn_p.t387 vdd2.t1112 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X939 out_n.t1373 vn_p.t388 vdd2.t1111 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X940 vdd2.t1110 vn_p.t389 out_n.t1372 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X941 out_n.t229 vn_n.t81 vss.t229 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X942 out_n.t1371 vn_p.t390 vdd2.t1109 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X943 vdd2.t1108 vn_p.t391 out_n.t1370 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X944 vss.t230 vn_n.t82 out_n.t230 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X945 out_n.t231 vn_n.t83 vss.t231 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X946 vdd1.t1106 vp_p.t393 out_p.t1049 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X947 vdd1.t1105 vp_p.t394 out_p.t1048 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X948 out_p.t1047 vp_p.t395 vdd1.t1104 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X949 vdd1.t1103 vp_p.t396 out_p.t1046 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X950 out_n.t1369 vn_p.t392 vdd2.t1107 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X951 out_p.t1045 vp_p.t397 vdd1.t1102 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X952 out_p.t1044 vp_p.t398 vdd1.t1101 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X953 out_p.t1043 vp_p.t399 vdd1.t1100 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X954 out_p.t1042 vp_p.t400 vdd1.t1099 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X955 vdd2.t1106 vn_p.t393 out_n.t1368 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X956 vdd1.t1098 vp_p.t401 out_p.t1041 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X957 vdd2.t1105 vn_p.t394 out_n.t1367 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X958 vdd1.t1097 vp_p.t402 out_p.t1040 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X959 out_p.t1039 vp_p.t403 vdd1.t1096 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X960 out_n.t1366 vn_p.t395 vdd2.t1104 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X961 vdd1.t1095 vp_p.t404 out_p.t1038 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X962 vdd1.t1094 vp_p.t405 out_p.t1037 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X963 vdd2.t1103 vn_p.t396 out_n.t1365 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X964 out_n.t1364 vn_p.t397 vdd2.t1102 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X965 out_n.t1363 vn_p.t398 vdd2.t1101 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X966 out_p.t1032 vp_p.t406 vdd1.t1093 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X967 vdd2.t1100 vn_p.t399 out_n.t1362 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X968 out_p.t1 vp_n.t77 vss.t484 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X969 out_p.t1036 vp_p.t407 vdd1.t1092 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X970 out_p.t1035 vp_p.t408 vdd1.t1091 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X971 out_n.t1361 vn_p.t400 vdd2.t1099 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X972 vdd2.t1098 vn_p.t401 out_n.t1360 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X973 out_n.t232 vn_n.t84 vss.t232 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X974 out_p.t1034 vp_p.t409 vdd1.t1090 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X975 out_n.t1359 vn_p.t402 vdd2.t1097 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X976 out_p.t1033 vp_p.t410 vdd1.t1089 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X977 vdd1.t1088 vp_p.t411 out_p.t605 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X978 vdd1.t1087 vp_p.t412 out_p.t597 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X979 out_n.t1358 vn_p.t403 vdd2.t1096 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X980 vdd1.t1086 vp_p.t413 out_p.t587 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X981 vdd1.t1085 vp_p.t414 out_p.t612 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X982 out_p.t579 vp_p.t415 vdd1.t1084 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X983 vdd2.t1095 vn_p.t404 out_n.t1357 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X984 out_n.t1356 vn_p.t405 vdd2.t1094 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X985 out_p.t2 vp_n.t78 vss.t483 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X986 out_p.t572 vp_p.t416 vdd1.t1083 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X987 out_p.t614 vp_p.t417 vdd1.t1082 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X988 vdd1.t1081 vp_p.t418 out_p.t564 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X989 vdd1.t1080 vp_p.t419 out_p.t586 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X990 vdd2.t1093 vn_p.t406 out_n.t1355 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X991 vdd2.t1092 vn_p.t407 out_n.t1354 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X992 out_p.t3 vp_n.t79 vss.t482 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X993 vdd2.t1091 vn_p.t408 out_n.t1353 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X994 vdd2.t1090 vn_p.t409 out_n.t1352 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X995 out_n.t1351 vn_p.t410 vdd2.t1089 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X996 vdd2.t1088 vn_p.t411 out_n.t1350 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X997 out_n.t1349 vn_p.t412 vdd2.t1087 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X998 out_p.t585 vp_p.t420 vdd1.t1079 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X999 vdd1.t1078 vp_p.t421 out_p.t595 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1000 vdd2.t1086 vn_p.t413 out_n.t1348 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1001 out_n.t1347 vn_p.t414 vdd2.t1085 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1002 out_p.t555 vp_p.t422 vdd1.t1077 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1003 vdd2.t1084 vn_p.t415 out_n.t1346 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1004 out_n.t89 vn_n.t85 vss.t89 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1005 out_n.t1345 vn_p.t416 vdd2.t1083 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1006 vdd2.t1082 vn_p.t417 out_n.t1344 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1007 out_p.t596 vp_p.t423 vdd1.t1076 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1008 vdd2.t1081 vn_p.t418 out_n.t1343 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1009 vdd2.t1080 vn_p.t419 out_n.t1342 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1010 out_n.t1341 vn_p.t420 vdd2.t1079 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1011 out_n.t1340 vn_p.t421 vdd2.t1078 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1012 out_n.t90 vn_n.t86 vss.t90 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1013 vdd2.t1077 vn_p.t422 out_n.t1339 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1014 out_p.t4 vp_n.t80 vss.t481 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1015 out_p.t5 vp_n.t81 vss.t480 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1016 out_n.t1338 vn_p.t423 vdd2.t1076 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1017 vss.t479 vp_n.t82 out_p.t6 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1018 vss.t91 vn_n.t87 out_n.t91 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1019 vdd2.t1075 vn_p.t424 out_n.t1337 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1020 out_n.t1336 vn_p.t425 vdd2.t1074 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1021 vss.t92 vn_n.t88 out_n.t92 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1022 out_n.t1335 vn_p.t426 vdd2.t1073 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1023 vdd2.t1072 vn_p.t427 out_n.t1334 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1024 out_p.t547 vp_p.t424 vdd1.t1075 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1025 out_p.t538 vp_p.t425 vdd1.t1074 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1026 vdd2.t1071 vn_p.t428 out_n.t1333 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1027 out_n.t1332 vn_p.t429 vdd2.t1070 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1028 vdd1.t1073 vp_p.t426 out_p.t530 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1029 out_p.t571 vp_p.t427 vdd1.t1072 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1030 out_n.t1331 vn_p.t430 vdd2.t1069 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1031 vdd1.t1071 vp_p.t428 out_p.t521 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1032 vdd1.t1070 vp_p.t429 out_p.t563 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1033 vdd1.t1069 vp_p.t430 out_p.t513 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1034 vdd1.t1068 vp_p.t431 out_p.t554 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1035 vdd2.t1068 vn_p.t431 out_n.t1330 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1036 out_p.t504 vp_p.t432 vdd1.t1067 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1037 out_n.t1329 vn_p.t432 vdd2.t1067 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1038 out_p.t546 vp_p.t433 vdd1.t1066 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1039 out_p.t496 vp_p.t434 vdd1.t1065 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1040 vdd1.t1064 vp_p.t435 out_p.t537 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1041 out_n.t1328 vn_p.t433 vdd2.t1066 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1042 vdd1.t1063 vp_p.t436 out_p.t487 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1043 out_n.t93 vn_n.t89 vss.t93 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1044 out_n.t1327 vn_p.t434 vdd2.t1065 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1045 out_p.t529 vp_p.t437 vdd1.t1062 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1046 vdd2.t1064 vn_p.t435 out_n.t1326 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1047 out_n.t1325 vn_p.t436 vdd2.t1063 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1048 out_n.t135 vn_n.t90 vss.t135 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1049 vdd2.t1062 vn_p.t437 out_n.t1324 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1050 vdd1.t1061 vp_p.t438 out_p.t479 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1051 vdd1.t1060 vp_p.t439 out_p.t520 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1052 vdd2.t1061 vn_p.t438 out_n.t1323 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1053 vdd1.t1059 vp_p.t440 out_p.t470 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1054 vdd1.t1058 vp_p.t441 out_p.t512 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1055 vdd2.t1060 vn_p.t439 out_n.t1322 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1056 out_n.t1321 vn_p.t440 vdd2.t1059 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1057 vdd2.t1058 vn_p.t441 out_n.t1320 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1058 vdd2.t1057 vn_p.t442 out_n.t1319 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1059 out_p.t462 vp_p.t442 vdd1.t1057 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1060 vdd2.t1056 vn_p.t443 out_n.t1318 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1061 out_p.t503 vp_p.t443 vdd1.t1056 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1062 out_p.t453 vp_p.t444 vdd1.t1055 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1063 vdd2.t1055 vn_p.t444 out_n.t1317 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1064 vss.t478 vp_n.t83 out_p.t7 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1065 out_p.t8 vp_n.t84 vss.t477 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1066 out_p.t495 vp_p.t445 vdd1.t1054 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1067 vss.t476 vp_n.t85 out_p.t9 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1068 vdd2.t1054 vn_p.t445 out_n.t1316 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1069 vdd1.t1053 vp_p.t446 out_p.t445 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1070 vdd1.t1052 vp_p.t447 out_p.t486 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1071 out_p.t436 vp_p.t448 vdd1.t1051 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1072 out_n.t1315 vn_p.t446 vdd2.t1053 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1073 out_n.t1314 vn_p.t447 vdd2.t1052 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1074 out_n.t1313 vn_p.t448 vdd2.t1051 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1075 vdd2.t1050 vn_p.t449 out_n.t1312 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1076 vss.t136 vn_n.t91 out_n.t136 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1077 vdd1.t1050 vp_p.t449 out_p.t478 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1078 vdd2.t1049 vn_p.t450 out_n.t1311 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1079 out_n.t1310 vn_p.t451 vdd2.t1048 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1080 out_n.t1309 vn_p.t452 vdd2.t1047 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1081 vss.t475 vp_n.t86 out_p.t10 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1082 out_n.t1308 vn_p.t453 vdd2.t1046 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1083 out_n.t1307 vn_p.t454 vdd2.t1045 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1084 vdd1.t1049 vp_p.t450 out_p.t428 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1085 vdd2.t1044 vn_p.t455 out_n.t1306 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1086 out_n.t137 vn_n.t92 vss.t137 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1087 out_n.t1305 vn_p.t456 vdd2.t1043 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1088 out_n.t1304 vn_p.t457 vdd2.t1042 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1089 out_p.t11 vp_n.t87 vss.t474 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1090 vss.t138 vn_n.t93 out_n.t138 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1091 vdd1.t1048 vp_p.t451 out_p.t469 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1092 vdd2.t1041 vn_p.t458 out_n.t1303 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1093 vdd2.t1040 vn_p.t459 out_n.t1302 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1094 vdd1.t1047 vp_p.t452 out_p.t418 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1095 vdd2.t1039 vn_p.t460 out_n.t1301 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1096 out_n.t1300 vn_p.t461 vdd2.t1038 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1097 out_p.t461 vp_p.t453 vdd1.t1046 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1098 vdd2.t1037 vn_p.t462 out_n.t1299 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1099 vdd1.t1045 vp_p.t454 out_p.t408 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1100 out_p.t452 vp_p.t455 vdd1.t1044 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1101 vdd2.t1036 vn_p.t463 out_n.t1298 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1102 out_n.t139 vn_n.t94 vss.t139 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1103 out_p.t398 vp_p.t456 vdd1.t1043 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1104 vdd1.t1042 vp_p.t457 out_p.t444 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1105 vdd2.t1035 vn_p.t464 out_n.t1297 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1106 vdd1.t1041 vp_p.t458 out_p.t388 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1107 out_p.t435 vp_p.t459 vdd1.t1040 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1108 vdd1.t1039 vp_p.t460 out_p.t377 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1109 out_p.t427 vp_p.t461 vdd1.t1038 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1110 out_p.t367 vp_p.t462 vdd1.t1037 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1111 out_p.t417 vp_p.t463 vdd1.t1036 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1112 vdd2.t1034 vn_p.t465 out_n.t1296 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1113 out_n.t1295 vn_p.t466 vdd2.t1033 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1114 vss.t473 vp_n.t88 out_p.t12 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1115 vdd1.t1035 vp_p.t464 out_p.t356 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1116 vdd2.t1032 vn_p.t467 out_n.t1294 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1117 out_p.t384 vp_p.t465 vdd1.t1034 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1118 vdd1.t1033 vp_p.t466 out_p.t407 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1119 vdd1.t1032 vp_p.t467 out_p.t346 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1120 out_n.t1293 vn_p.t468 vdd2.t1031 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1121 vdd2.t1030 vn_p.t469 out_n.t1292 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1122 out_n.t174 vn_n.t95 vss.t174 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1123 out_n.t1291 vn_p.t470 vdd2.t1029 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1124 vdd1.t1031 vp_p.t468 out_p.t397 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1125 out_n.t1290 vn_p.t471 vdd2.t1028 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1126 vdd1.t1030 vp_p.t469 out_p.t335 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1127 out_p.t363 vp_p.t470 vdd1.t1029 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1128 out_n.t1289 vn_p.t472 vdd2.t1027 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1129 out_p.t387 vp_p.t471 vdd1.t1028 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1130 vdd1.t1027 vp_p.t472 out_p.t325 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1131 out_p.t376 vp_p.t473 vdd1.t1026 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1132 vdd1.t1025 vp_p.t474 out_p.t314 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1133 vdd1.t1024 vp_p.t475 out_p.t342 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1134 out_p.t366 vp_p.t476 vdd1.t1023 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1135 vdd2.t1026 vn_p.t473 out_n.t1288 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1136 vss.t175 vn_n.t96 out_n.t175 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1137 vss.t472 vp_n.t89 out_p.t13 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1138 vdd1.t1022 vp_p.t477 out_p.t304 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1139 out_n.t1287 vn_p.t474 vdd2.t1025 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1140 out_p.t355 vp_p.t478 vdd1.t1021 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1141 out_n.t1286 vn_p.t475 vdd2.t1024 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1142 out_p.t14 vp_n.t90 vss.t471 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1143 out_n.t1285 vn_p.t476 vdd2.t1023 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1144 out_p.t293 vp_p.t479 vdd1.t1020 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1145 vdd1.t1019 vp_p.t480 out_p.t292 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1146 vdd2.t1022 vn_p.t477 out_n.t1284 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1147 vdd2.t1021 vn_p.t478 out_n.t1283 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1148 out_n.t1282 vn_p.t479 vdd2.t1020 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1149 out_p.t321 vp_p.t481 vdd1.t1018 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1150 vdd2.t1019 vn_p.t480 out_n.t1281 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1151 out_n.t176 vn_n.t97 vss.t176 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1152 out_n.t1280 vn_p.t481 vdd2.t1018 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1153 out_p.t345 vp_p.t482 vdd1.t1017 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1154 vdd2.t1017 vn_p.t482 out_n.t1279 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1155 vss.t470 vp_n.t91 out_p.t15 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1156 out_p.t284 vp_p.t483 vdd1.t1016 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1157 out_p.t334 vp_p.t484 vdd1.t1015 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1158 out_p.t275 vp_p.t485 vdd1.t1014 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1159 vdd1.t1013 vp_p.t486 out_p.t274 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1160 vdd2.t1016 vn_p.t483 out_n.t1278 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1161 vss.t469 vp_n.t92 out_p.t16 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1162 out_n.t177 vn_n.t98 vss.t177 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1163 out_n.t1277 vn_p.t484 vdd2.t1015 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1164 out_n.t1276 vn_p.t485 vdd2.t1014 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1165 vss.t468 vp_n.t93 out_p.t17 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1166 out_n.t1275 vn_p.t486 vdd2.t1013 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1167 out_n.t1274 vn_p.t487 vdd2.t1012 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1168 vdd2.t1011 vn_p.t488 out_n.t1273 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1169 out_p.t300 vp_p.t487 vdd1.t1012 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1170 vdd2.t1010 vn_p.t489 out_n.t1272 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1171 out_p.t324 vp_p.t488 vdd1.t1011 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1172 vdd1.t1010 vp_p.t489 out_p.t934 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1173 out_p.t935 vp_p.t490 vdd1.t1009 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1174 out_p.t936 vp_p.t491 vdd1.t1008 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1175 vdd1.t1007 vp_p.t492 out_p.t924 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1176 vdd1.t1006 vp_p.t493 out_p.t940 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1177 vdd1.t1005 vp_p.t494 out_p.t939 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1178 out_p.t928 vp_p.t495 vdd1.t1004 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1179 vss.t178 vn_n.t99 out_n.t178 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1180 vdd1.t1003 vp_p.t496 out_p.t914 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1181 vdd1.t1002 vp_p.t497 out_p.t918 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1182 out_p.t904 vp_p.t498 vdd1.t1001 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1183 vss.t100 vn_n.t100 out_n.t100 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1184 vdd1.t1000 vp_p.t499 out_p.t908 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1185 vdd1.t999 vp_p.t500 out_p.t894 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1186 out_n.t1271 vn_p.t490 vdd2.t1009 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1187 out_p.t898 vp_p.t501 vdd1.t998 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1188 out_n.t1270 vn_p.t491 vdd2.t1008 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1189 vdd2.t1007 vn_p.t492 out_n.t1269 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1190 vdd1.t997 vp_p.t502 out_p.t884 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1191 out_p.t18 vp_n.t94 vss.t467 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1192 out_p.t888 vp_p.t503 vdd1.t996 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1193 out_n.t1268 vn_p.t493 vdd2.t1006 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1194 out_n.t101 vn_n.t101 vss.t101 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1195 vdd2.t1005 vn_p.t494 out_n.t1267 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1196 vss.t102 vn_n.t102 out_n.t102 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1197 out_p.t874 vp_p.t504 vdd1.t995 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1198 vdd1.t994 vp_p.t505 out_p.t878 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1199 out_p.t864 vp_p.t506 vdd1.t993 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1200 vdd1.t992 vp_p.t507 out_p.t868 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1201 vdd2.t1004 vn_p.t495 out_n.t1266 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1202 vdd1.t991 vp_p.t508 out_p.t854 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1203 vdd2.t1003 vn_p.t496 out_n.t1265 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1204 out_p.t858 vp_p.t509 vdd1.t990 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1205 vdd2.t1002 vn_p.t497 out_n.t1264 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1206 out_n.t1263 vn_p.t498 vdd2.t1001 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1207 out_n.t103 vn_n.t103 vss.t103 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1208 vdd1.t989 vp_p.t510 out_p.t844 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1209 vdd2.t1000 vn_p.t499 out_n.t1262 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1210 vss.t466 vp_n.t95 out_p.t1780 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1211 vdd2.t999 vn_p.t500 out_n.t1261 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1212 out_p.t848 vp_p.t511 vdd1.t988 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1213 out_n.t1260 vn_p.t501 vdd2.t998 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1214 vdd2.t997 vn_p.t502 out_n.t1259 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1215 vss.t104 vn_n.t104 out_n.t104 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1216 out_n.t1258 vn_p.t503 vdd2.t996 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1217 out_n.t1257 vn_p.t504 vdd2.t995 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1218 vdd1.t987 vp_p.t512 out_p.t834 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1219 vdd1.t986 vp_p.t513 out_p.t838 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1220 out_p.t824 vp_p.t514 vdd1.t985 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1221 out_p.t828 vp_p.t515 vdd1.t984 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1222 vdd2.t994 vn_p.t505 out_n.t1256 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1223 vdd2.t993 vn_p.t506 out_n.t1255 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1224 vss.t465 vp_n.t96 out_p.t1781 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1225 out_n.t1254 vn_p.t507 vdd2.t992 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1226 out_p.t1782 vp_n.t97 vss.t464 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1227 out_n.t1253 vn_p.t508 vdd2.t991 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1228 vss.t105 vn_n.t105 out_n.t105 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1229 vdd2.t990 vn_p.t509 out_n.t1252 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1230 vdd1.t983 vp_p.t516 out_p.t814 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1231 vdd1.t982 vp_p.t517 out_p.t818 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1232 out_p.t804 vp_p.t518 vdd1.t981 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1233 vdd2.t989 vn_p.t510 out_n.t1251 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1234 out_n.t1250 vn_p.t511 vdd2.t988 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1235 out_p.t808 vp_p.t519 vdd1.t980 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1236 out_p.t794 vp_p.t520 vdd1.t979 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1237 out_p.t798 vp_p.t521 vdd1.t978 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1238 out_p.t784 vp_p.t522 vdd1.t977 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1239 out_p.t788 vp_p.t523 vdd1.t976 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1240 vdd1.t975 vp_p.t524 out_p.t774 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1241 out_n.t1249 vn_p.t512 vdd2.t987 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1242 vss.t463 vp_n.t98 out_p.t1783 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1243 vdd1.t974 vp_p.t525 out_p.t778 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1244 vdd1.t973 vp_p.t526 out_p.t764 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1245 out_p.t768 vp_p.t527 vdd1.t972 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1246 out_p.t754 vp_p.t528 vdd1.t971 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1247 vdd2.t986 vn_p.t513 out_n.t1248 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1248 vdd2.t985 vn_p.t514 out_n.t1247 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1249 out_p.t1784 vp_n.t99 vss.t462 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1250 vdd1.t970 vp_p.t529 out_p.t758 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1251 out_p.t744 vp_p.t530 vdd1.t969 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1252 vdd2.t984 vn_p.t515 out_n.t1246 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1253 vdd1.t968 vp_p.t531 out_p.t748 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1254 vss.t461 vp_n.t100 out_p.t1785 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1255 vdd1.t967 vp_p.t532 out_p.t734 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1256 out_p.t738 vp_p.t533 vdd1.t966 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1257 out_p.t724 vp_p.t534 vdd1.t965 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1258 out_n.t106 vn_n.t106 vss.t106 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1259 vss.t107 vn_n.t107 out_n.t107 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1260 vdd2.t983 vn_p.t516 out_n.t1245 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1261 out_n.t108 vn_n.t108 vss.t108 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1262 vdd1.t964 vp_p.t535 out_p.t728 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1263 vdd2.t982 vn_p.t517 out_n.t1244 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1264 out_n.t1243 vn_p.t518 vdd2.t981 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1265 out_n.t1242 vn_p.t519 vdd2.t980 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1266 out_n.t1241 vn_p.t520 vdd2.t979 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1267 vdd2.t978 vn_p.t521 out_n.t1240 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1268 vdd1.t963 vp_p.t536 out_p.t714 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1269 vdd2.t977 vn_p.t522 out_n.t1239 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1270 out_n.t1238 vn_p.t523 vdd2.t976 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1271 out_p.t1786 vp_n.t101 vss.t460 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1272 out_p.t718 vp_p.t537 vdd1.t962 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1273 vdd2.t975 vn_p.t524 out_n.t1237 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1274 out_n.t1236 vn_p.t525 vdd2.t974 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1275 vdd2.t973 vn_p.t526 out_n.t1235 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1276 out_n.t1234 vn_p.t527 vdd2.t972 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1277 vss.t109 vn_n.t109 out_n.t109 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1278 out_n.t1233 vn_p.t528 vdd2.t971 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1279 out_n.t1232 vn_p.t529 vdd2.t970 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1280 vdd1.t961 vp_p.t538 out_p.t704 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1281 out_n.t1231 vn_p.t530 vdd2.t969 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1282 vdd2.t968 vn_p.t531 out_n.t1230 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1283 out_p.t708 vp_p.t539 vdd1.t960 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1284 vdd2.t967 vn_p.t532 out_n.t1229 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1285 out_n.t1228 vn_p.t533 vdd2.t966 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1286 out_p.t693 vp_p.t540 vdd1.t959 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1287 out_n.t1227 vn_p.t534 vdd2.t965 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1288 out_p.t697 vp_p.t541 vdd1.t958 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1289 out_n.t1226 vn_p.t535 vdd2.t964 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1290 vdd1.t957 vp_p.t542 out_p.t682 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1291 out_n.t120 vn_n.t110 vss.t120 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1292 vdd2.t963 vn_p.t536 out_n.t1225 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1293 vdd1.t956 vp_p.t543 out_p.t686 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1294 out_p.t672 vp_p.t544 vdd1.t955 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1295 vdd1.t954 vp_p.t545 out_p.t662 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1296 out_n.t1224 vn_p.t537 vdd2.t962 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1297 vdd2.t961 vn_p.t538 out_n.t1223 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1298 vss.t459 vp_n.t102 out_p.t1787 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1299 vdd2.t960 vn_p.t539 out_n.t1222 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1300 vdd1.t953 vp_p.t546 out_p.t650 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1301 out_p.t654 vp_p.t547 vdd1.t952 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1302 vdd2.t959 vn_p.t540 out_n.t1221 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1303 vdd1.t951 vp_p.t548 out_p.t639 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1304 out_p.t643 vp_p.t549 vdd1.t950 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1305 out_n.t1220 vn_p.t541 vdd2.t958 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1306 out_p.t627 vp_p.t550 vdd1.t949 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1307 vdd2.t957 vn_p.t542 out_n.t1219 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1308 vdd2.t956 vn_p.t543 out_n.t1218 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1309 vdd1.t948 vp_p.t551 out_p.t659 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1310 vdd1.t947 vp_p.t552 out_p.t644 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1311 vdd1.t946 vp_p.t553 out_p.t631 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1312 out_p.t615 vp_p.t554 vdd1.t945 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1313 vdd2.t955 vn_p.t544 out_n.t1217 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1314 out_p.t1788 vp_n.t103 vss.t458 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1315 out_p.t1789 vp_n.t104 vss.t457 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1316 out_p.t632 vp_p.t555 vdd1.t944 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1317 vdd1.t943 vp_p.t556 out_p.t620 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1318 vss.t121 vn_n.t111 out_n.t121 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1319 vdd2.t954 vn_p.t545 out_n.t1216 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1320 vss.t456 vp_n.t105 out_p.t1790 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1321 vdd1.t942 vp_p.t557 out_p.t625 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1322 out_p.t626 vp_p.t558 vdd1.t941 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1323 vss.t122 vn_n.t112 out_n.t122 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1324 out_n.t1215 vn_p.t546 vdd2.t953 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1325 out_n.t1214 vn_p.t547 vdd2.t952 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1326 out_p.t958 vp_p.t559 vdd1.t940 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1327 vdd1.t939 vp_p.t560 out_p.t955 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1328 out_n.t1213 vn_p.t548 vdd2.t951 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1329 vdd2.t950 vn_p.t549 out_n.t1212 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1330 out_n.t1211 vn_p.t550 vdd2.t949 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1331 vdd1.t938 vp_p.t561 out_p.t959 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1332 out_n.t1210 vn_p.t551 vdd2.t948 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1333 out_n.t1209 vn_p.t552 vdd2.t947 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1334 out_n.t1208 vn_p.t553 vdd2.t946 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1335 out_n.t1207 vn_p.t554 vdd2.t945 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1336 out_n.t1206 vn_p.t555 vdd2.t944 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1337 out_n.t1205 vn_p.t556 vdd2.t943 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1338 out_n.t1204 vn_p.t557 vdd2.t942 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1339 vdd2.t941 vn_p.t558 out_n.t1203 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1340 out_n.t1202 vn_p.t559 vdd2.t940 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1341 vss.t455 vp_n.t106 out_p.t1791 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1342 vdd2.t939 vn_p.t560 out_n.t1201 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1343 vdd2.t938 vn_p.t561 out_n.t1200 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1344 vdd2.t937 vn_p.t562 out_n.t1199 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1345 out_n.t1198 vn_p.t563 vdd2.t936 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1346 out_n.t123 vn_n.t113 vss.t123 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1347 out_n.t1197 vn_p.t564 vdd2.t935 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1348 vdd2.t934 vn_p.t565 out_n.t1196 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1349 vdd2.t933 vn_p.t566 out_n.t1195 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1350 vdd2.t932 vn_p.t567 out_n.t1194 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1351 vdd1.t937 vp_p.t562 out_p.t1031 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1352 vdd1.t936 vp_p.t563 out_p.t1029 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1353 vdd2.t931 vn_p.t568 out_n.t1193 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1354 vdd2.t930 vn_p.t569 out_n.t1192 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1355 vdd1.t935 vp_p.t564 out_p.t967 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1356 out_p.t1018 vp_p.t565 vdd1.t934 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1357 out_n.t1191 vn_p.t570 vdd2.t929 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1358 vdd2.t928 vn_p.t571 out_n.t1190 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1359 vdd1.t933 vp_p.t566 out_p.t1012 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1360 vss.t124 vn_n.t114 out_n.t124 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1361 out_n.t223 vn_n.t115 vss.t223 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1362 out_p.t1006 vp_p.t567 vdd1.t932 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1363 out_n.t224 vn_n.t116 vss.t224 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1364 out_n.t1189 vn_p.t572 vdd2.t927 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1365 vdd1.t931 vp_p.t568 out_p.t1000 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1366 out_n.t1188 vn_p.t573 vdd2.t926 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1367 out_p.t993 vp_p.t569 vdd1.t930 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1368 vdd1.t929 vp_p.t570 out_p.t987 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1369 out_p.t981 vp_p.t571 vdd1.t928 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1370 vdd1.t927 vp_p.t572 out_p.t975 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1371 vdd1.t926 vp_p.t573 out_p.t969 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1372 out_n.t1187 vn_p.t574 vdd2.t925 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1373 vdd2.t924 vn_p.t575 out_n.t1186 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1374 out_n.t1185 vn_p.t576 vdd2.t923 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1375 vdd1.t925 vp_p.t574 out_p.t1030 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1376 vdd1.t924 vp_p.t575 out_p.t1087 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1377 vss.t225 vn_n.t117 out_n.t225 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1378 vdd1.t923 vp_p.t576 out_p.t1084 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1379 out_p.t609 vp_p.t577 vdd1.t922 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1380 out_p.t1028 vp_p.t578 vdd1.t921 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1381 out_p.t584 vp_p.t579 vdd1.t920 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1382 vss.t454 vp_n.t107 out_p.t1792 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1383 out_n.t1184 vn_p.t577 vdd2.t922 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1384 out_p.t594 vp_p.t580 vdd1.t919 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1385 out_n.t1183 vn_p.t578 vdd2.t921 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1386 vdd1.t918 vp_p.t581 out_p.t604 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1387 vdd1.t917 vp_p.t582 out_p.t953 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1388 vdd2.t920 vn_p.t579 out_n.t1182 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1389 vdd1.t916 vp_p.t583 out_p.t954 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1390 vdd1.t915 vp_p.t584 out_p.t298 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1391 out_p.t289 vp_p.t585 vdd1.t914 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1392 out_n.t1181 vn_p.t580 vdd2.t919 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1393 out_p.t1793 vp_n.t108 vss.t453 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1394 out_p.t313 vp_p.t586 vdd1.t913 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1395 vdd2.t918 vn_p.t581 out_n.t1180 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1396 out_n.t1179 vn_p.t582 vdd2.t917 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1397 vdd1.t912 vp_p.t587 out_p.t282 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1398 vdd2.t916 vn_p.t583 out_n.t1178 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1399 vdd1.t911 vp_p.t588 out_p.t303 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1400 vdd2.t915 vn_p.t584 out_n.t1177 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1401 out_p.t670 vp_p.t589 vdd1.t910 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1402 vdd2.t914 vn_p.t585 out_n.t1176 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1403 vdd2.t913 vn_p.t586 out_n.t1175 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1404 out_n.t1174 vn_p.t587 vdd2.t912 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1405 out_p.t961 vp_p.t590 vdd1.t909 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1406 vdd2.t911 vn_p.t588 out_n.t1173 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1407 vdd2.t910 vn_p.t589 out_n.t1172 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1408 out_n.t1171 vn_p.t590 vdd2.t909 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1409 out_n.t226 vn_n.t118 vss.t226 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1410 vdd2.t908 vn_p.t591 out_n.t1170 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1411 out_p.t952 vp_p.t591 vdd1.t908 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1412 vdd2.t907 vn_p.t592 out_n.t1169 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1413 out_p.t1794 vp_n.t109 vss.t452 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1414 out_n.t1168 vn_p.t593 vdd2.t906 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1415 vdd2.t905 vn_p.t594 out_n.t1167 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1416 vss.t451 vp_n.t110 out_p.t1795 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1417 out_n.t1166 vn_p.t595 vdd2.t904 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1418 vdd2.t903 vn_p.t596 out_n.t1165 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1419 out_n.t1164 vn_p.t597 vdd2.t902 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1420 out_n.t1163 vn_p.t598 vdd2.t901 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1421 vss.t227 vn_n.t119 out_n.t227 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1422 out_n.t1162 vn_p.t599 vdd2.t900 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1423 out_p.t960 vp_p.t592 vdd1.t907 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1424 out_p.t1083 vp_p.t593 vdd1.t906 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1425 out_p.t1021 vp_p.t594 vdd1.t905 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1426 out_p.t1019 vp_p.t595 vdd1.t904 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1427 vdd1.t903 vp_p.t596 out_p.t1013 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1428 vdd1.t902 vp_p.t597 out_p.t1007 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1429 out_n.t1161 vn_p.t600 vdd2.t899 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1430 out_p.t1001 vp_p.t598 vdd1.t901 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1431 out_p.t994 vp_p.t599 vdd1.t900 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1432 vss.t213 vn_n.t120 out_n.t213 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1433 out_n.t1160 vn_p.t601 vdd2.t898 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1434 vdd1.t899 vp_p.t600 out_p.t988 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1435 vdd1.t898 vp_p.t601 out_p.t982 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1436 vdd1.t897 vp_p.t602 out_p.t976 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1437 vdd2.t897 vn_p.t602 out_n.t1159 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1438 out_p.t970 vp_p.t603 vdd1.t896 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1439 out_n.t1158 vn_p.t603 vdd2.t896 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1440 vdd2.t895 vn_p.t604 out_n.t1157 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1441 vdd2.t894 vn_p.t605 out_n.t1156 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1442 vdd1.t895 vp_p.t604 out_p.t963 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1443 vdd1.t894 vp_p.t605 out_p.t1024 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1444 out_n.t1155 vn_p.t606 vdd2.t893 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1445 out_p.t1015 vp_p.t606 vdd1.t893 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1446 out_p.t1009 vp_p.t607 vdd1.t892 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1447 out_n.t214 vn_n.t121 vss.t214 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1448 out_p.t1003 vp_p.t608 vdd1.t891 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1449 vdd1.t890 vp_p.t609 out_p.t997 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1450 vdd2.t892 vn_p.t607 out_n.t1154 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1451 vss.t450 vp_n.t111 out_p.t1796 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1452 vdd1.t889 vp_p.t610 out_p.t990 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1453 vdd1.t888 vp_p.t611 out_p.t984 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1454 vdd1.t887 vp_p.t612 out_p.t978 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1455 vdd1.t886 vp_p.t613 out_p.t972 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1456 out_n.t215 vn_n.t122 vss.t215 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1457 vdd2.t891 vn_p.t608 out_n.t1153 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1458 vdd1.t885 vp_p.t614 out_p.t965 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1459 vdd1.t884 vp_p.t615 out_p.t1026 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1460 out_p.t611 vp_p.t616 vdd1.t883 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1461 out_n.t1152 vn_p.t609 vdd2.t890 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1462 vdd2.t889 vn_p.t610 out_n.t1151 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1463 out_n.t1150 vn_p.t611 vdd2.t888 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1464 vdd2.t887 vn_p.t612 out_n.t1149 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1465 vdd1.t882 vp_p.t617 out_p.t613 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1466 vdd2.t886 vn_p.t613 out_n.t1148 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1467 vss.t449 vp_n.t112 out_p.t1797 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1468 vdd1.t881 vp_p.t618 out_p.t603 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1469 vdd1.t880 vp_p.t619 out_p.t593 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1470 out_p.t576 vp_p.t620 vdd1.t879 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1471 out_p.t577 vp_p.t621 vdd1.t878 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1472 vss.t448 vp_n.t113 out_p.t1798 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1473 vss.t216 vn_n.t123 out_n.t216 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1474 out_n.t217 vn_n.t124 vss.t217 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1475 out_n.t1147 vn_p.t614 vdd2.t885 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1476 vdd1.t877 vp_p.t622 out_p.t578 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1477 out_n.t1146 vn_p.t615 vdd2.t884 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1478 out_p.t570 vp_p.t623 vdd1.t876 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1479 vdd1.t875 vp_p.t624 out_p.t561 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1480 vdd2.t883 vn_p.t616 out_n.t1145 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1481 out_n.t1144 vn_p.t617 vdd2.t882 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1482 vdd2.t881 vn_p.t618 out_n.t1143 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1483 out_p.t1799 vp_n.t114 vss.t447 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1484 out_n.t1142 vn_p.t619 vdd2.t880 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1485 vss.t446 vp_n.t115 out_p.t1757 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1486 vdd1.t874 vp_p.t625 out_p.t562 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1487 vss.t199 vn_n.t125 out_n.t199 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1488 vss.t445 vp_n.t116 out_p.t1758 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1489 vss.t444 vp_n.t117 out_p.t1759 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1490 out_n.t1141 vn_p.t620 vdd2.t879 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1491 out_p.t1760 vp_n.t118 vss.t443 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1492 out_n.t1140 vn_p.t621 vdd2.t878 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1493 vdd2.t877 vn_p.t622 out_n.t1139 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1494 out_p.t553 vp_p.t626 vdd1.t873 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1495 vdd2.t876 vn_p.t623 out_n.t1138 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1496 out_p.t544 vp_p.t627 vdd1.t872 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1497 vdd2.t875 vn_p.t624 out_n.t1137 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1498 out_n.t1136 vn_p.t625 vdd2.t874 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1499 vdd1.t871 vp_p.t628 out_p.t545 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1500 vdd2.t873 vn_p.t626 out_n.t1135 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1501 out_n.t1134 vn_p.t627 vdd2.t872 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1502 vdd1.t870 vp_p.t629 out_p.t536 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1503 vdd1.t869 vp_p.t630 out_p.t527 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1504 out_p.t528 vp_p.t631 vdd1.t868 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1505 out_n.t1133 vn_p.t628 vdd2.t871 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1506 out_p.t519 vp_p.t632 vdd1.t867 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1507 vdd1.t866 vp_p.t633 out_p.t510 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1508 out_p.t511 vp_p.t634 vdd1.t865 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1509 out_n.t200 vn_n.t126 vss.t200 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1510 out_p.t502 vp_p.t635 vdd1.t864 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1511 out_p.t493 vp_p.t636 vdd1.t863 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1512 out_p.t494 vp_p.t637 vdd1.t862 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1513 vdd2.t870 vn_p.t629 out_n.t1132 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1514 out_p.t485 vp_p.t638 vdd1.t861 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1515 out_n.t201 vn_n.t127 vss.t201 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1516 vdd2.t869 vn_p.t630 out_n.t1131 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1517 vdd1.t860 vp_p.t639 out_p.t476 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1518 out_p.t477 vp_p.t640 vdd1.t859 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1519 vdd1.t858 vp_p.t641 out_p.t468 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1520 out_p.t459 vp_p.t642 vdd1.t857 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1521 out_n.t1130 vn_p.t631 vdd2.t868 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1522 vdd2.t867 vn_p.t632 out_n.t1129 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1523 out_n.t1128 vn_p.t633 vdd2.t866 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1524 vdd1.t856 vp_p.t643 out_p.t460 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1525 vdd2.t865 vn_p.t634 out_n.t1127 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1526 out_p.t451 vp_p.t644 vdd1.t855 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1527 out_p.t442 vp_p.t645 vdd1.t854 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1528 out_p.t443 vp_p.t646 vdd1.t853 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1529 out_p.t434 vp_p.t647 vdd1.t852 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1530 out_p.t424 vp_p.t648 vdd1.t851 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1531 out_n.t1126 vn_p.t635 vdd2.t864 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1532 vdd2.t863 vn_p.t636 out_n.t1125 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1533 out_p.t425 vp_p.t649 vdd1.t850 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1534 out_n.t1124 vn_p.t637 vdd2.t862 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1535 vdd1.t849 vp_p.t650 out_p.t414 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1536 vdd1.t848 vp_p.t651 out_p.t426 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1537 vss.t442 vp_n.t119 out_p.t1761 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1538 vdd1.t847 vp_p.t652 out_p.t415 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1539 out_p.t1762 vp_n.t120 vss.t441 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1540 vdd2.t861 vn_p.t638 out_n.t1123 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1541 vss.t202 vn_n.t128 out_n.t202 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1542 out_n.t203 vn_n.t129 vss.t203 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1543 out_n.t1122 vn_p.t639 vdd2.t860 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1544 vss.t189 vn_n.t130 out_n.t189 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1545 out_p.t404 vp_p.t653 vdd1.t846 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1546 vdd2.t859 vn_p.t640 out_n.t1121 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1547 out_n.t1120 vn_p.t641 vdd2.t858 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1548 out_p.t416 vp_p.t654 vdd1.t845 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1549 out_n.t1119 vn_p.t642 vdd2.t857 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1550 vdd1.t844 vp_p.t655 out_p.t405 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1551 vdd2.t856 vn_p.t643 out_n.t1118 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1552 out_n.t1117 vn_p.t644 vdd2.t855 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1553 out_n.t1116 vn_p.t645 vdd2.t854 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1554 vdd2.t853 vn_p.t646 out_n.t1115 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1555 out_n.t190 vn_n.t131 vss.t190 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1556 vdd2.t852 vn_p.t647 out_n.t1114 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1557 vss.t440 vp_n.t121 out_p.t1763 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1558 out_p.t1764 vp_n.t122 vss.t439 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1559 out_p.t394 vp_p.t656 vdd1.t843 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1560 vdd2.t851 vn_p.t648 out_n.t1113 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1561 vdd2.t850 vn_p.t649 out_n.t1112 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1562 vdd2.t849 vn_p.t650 out_n.t1111 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1563 vss.t438 vp_n.t123 out_p.t1765 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1564 out_n.t1110 vn_p.t651 vdd2.t848 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1565 out_p.t406 vp_p.t657 vdd1.t842 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1566 out_p.t395 vp_p.t658 vdd1.t841 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1567 vdd2.t847 vn_p.t652 out_n.t1109 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1568 vdd1.t840 vp_p.t659 out_p.t383 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1569 out_p.t396 vp_p.t660 vdd1.t839 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1570 out_p.t385 vp_p.t661 vdd1.t838 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1571 out_n.t1108 vn_p.t653 vdd2.t846 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1572 vdd2.t845 vn_p.t654 out_n.t1107 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1573 vdd1.t837 vp_p.t662 out_p.t373 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1574 vss.t191 vn_n.t132 out_n.t191 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1575 out_p.t386 vp_p.t663 vdd1.t836 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1576 out_p.t374 vp_p.t664 vdd1.t835 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1577 vdd1.t834 vp_p.t665 out_p.t362 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1578 vdd1.t833 vp_p.t666 out_p.t375 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1579 out_n.t1106 vn_p.t655 vdd2.t844 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1580 vdd1.t832 vp_p.t667 out_p.t364 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1581 out_p.t352 vp_p.t668 vdd1.t831 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1582 vdd1.t830 vp_p.t669 out_p.t365 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1583 out_n.t1105 vn_p.t656 vdd2.t843 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1584 vdd2.t842 vn_p.t657 out_n.t1104 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1585 vdd2.t841 vn_p.t658 out_n.t1103 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1586 out_p.t1766 vp_n.t124 vss.t437 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1587 out_p.t353 vp_p.t670 vdd1.t829 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1588 vdd1.t828 vp_p.t671 out_p.t341 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1589 out_n.t1102 vn_p.t659 vdd2.t840 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1590 vdd1.t827 vp_p.t672 out_p.t354 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1591 out_n.t1101 vn_p.t660 vdd2.t839 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1592 out_p.t343 vp_p.t673 vdd1.t826 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1593 out_n.t1100 vn_p.t661 vdd2.t838 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1594 out_n.t1099 vn_p.t662 vdd2.t837 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1595 vdd2.t836 vn_p.t663 out_n.t1098 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1596 out_p.t331 vp_p.t674 vdd1.t825 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1597 out_n.t1097 vn_p.t664 vdd2.t835 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1598 out_n.t1096 vn_p.t665 vdd2.t834 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1599 out_p.t344 vp_p.t675 vdd1.t824 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1600 vdd1.t823 vp_p.t676 out_p.t332 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1601 out_p.t320 vp_p.t677 vdd1.t822 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1602 vdd1.t821 vp_p.t678 out_p.t333 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1603 out_n.t1095 vn_p.t666 vdd2.t833 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1604 vdd1.t820 vp_p.t679 out_p.t322 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1605 out_p.t310 vp_p.t680 vdd1.t819 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1606 vdd2.t832 vn_p.t667 out_n.t1094 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1607 out_n.t192 vn_n.t133 vss.t192 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1608 vdd1.t818 vp_p.t681 out_p.t323 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1609 out_n.t1093 vn_p.t668 vdd2.t831 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1610 out_p.t297 vp_p.t682 vdd1.t817 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1611 out_p.t311 vp_p.t683 vdd1.t816 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1612 vdd2.t830 vn_p.t669 out_n.t1092 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1613 out_n.t1091 vn_p.t670 vdd2.t829 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1614 out_p.t299 vp_p.t684 vdd1.t815 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1615 vdd2.t828 vn_p.t671 out_n.t1090 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1616 vdd2.t827 vn_p.t672 out_n.t1089 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1617 vdd2.t826 vn_p.t673 out_n.t1088 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1618 vss.t436 vp_n.t125 out_p.t1767 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1619 vdd2.t825 vn_p.t674 out_n.t1087 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1620 out_n.t193 vn_n.t134 vss.t193 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1621 vdd2.t824 vn_p.t675 out_n.t1086 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1622 vdd2.t823 vn_p.t676 out_n.t1085 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1623 vdd1.t814 vp_p.t685 out_p.t312 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1624 vdd2.t822 vn_p.t677 out_n.t1084 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1625 out_p.t301 vp_p.t686 vdd1.t813 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1626 vdd1.t812 vp_p.t687 out_p.t290 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1627 vdd2.t821 vn_p.t678 out_n.t1083 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1628 out_p.t1768 vp_n.t126 vss.t435 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1629 vss.t434 vp_n.t127 out_p.t1769 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1630 out_n.t194 vn_n.t135 vss.t194 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1631 out_n.t1082 vn_p.t679 vdd2.t820 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1632 out_p.t1770 vp_n.t128 vss.t433 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1633 vdd1.t811 vp_p.t688 out_p.t302 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1634 vdd2.t819 vn_p.t680 out_n.t1081 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1635 out_n.t1080 vn_p.t681 vdd2.t818 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1636 out_p.t291 vp_p.t689 vdd1.t810 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1637 out_n.t1079 vn_p.t682 vdd2.t817 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1638 vdd2.t816 vn_p.t683 out_n.t1078 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1639 out_n.t1077 vn_p.t684 vdd2.t815 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1640 out_n.t1076 vn_p.t685 vdd2.t814 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1641 out_p.t1771 vp_n.t129 vss.t432 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1642 vdd2.t813 vn_p.t686 out_n.t1075 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1643 out_n.t1074 vn_p.t687 vdd2.t812 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1644 out_p.t1772 vp_n.t130 vss.t431 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1645 out_n.t1073 vn_p.t688 vdd2.t811 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1646 out_p.t280 vp_p.t690 vdd1.t809 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1647 vdd2.t810 vn_p.t689 out_n.t1072 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1648 vdd1.t808 vp_p.t691 out_p.t281 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1649 vdd1.t807 vp_p.t692 out_p.t283 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1650 out_n.t1071 vn_p.t690 vdd2.t809 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1651 vdd1.t806 vp_p.t693 out_p.t937 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1652 vdd1.t805 vp_p.t694 out_p.t938 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1653 out_n.t195 vn_n.t136 vss.t195 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1654 vss.t196 vn_n.t137 out_n.t196 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1655 vdd2.t808 vn_p.t691 out_n.t1070 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1656 out_n.t1069 vn_p.t692 vdd2.t807 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1657 vdd1.t804 vp_p.t695 out_p.t930 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1658 out_n.t1068 vn_p.t693 vdd2.t806 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1659 out_p.t929 vp_p.t696 vdd1.t803 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1660 vdd1.t802 vp_p.t697 out_p.t920 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1661 out_p.t941 vp_p.t698 vdd1.t801 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1662 vdd1.t800 vp_p.t699 out_p.t919 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1663 out_p.t910 vp_p.t700 vdd1.t799 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1664 vdd1.t798 vp_p.t701 out_p.t909 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1665 out_p.t900 vp_p.t702 vdd1.t797 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1666 out_p.t933 vp_p.t703 vdd1.t796 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1667 out_n.t1067 vn_p.t694 vdd2.t805 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1668 out_n.t1066 vn_p.t695 vdd2.t804 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1669 vdd2.t803 vn_p.t696 out_n.t1065 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1670 out_p.t899 vp_p.t704 vdd1.t795 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1671 vdd2.t802 vn_p.t697 out_n.t1064 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1672 vss.t430 vp_n.t131 out_p.t1773 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1673 vdd1.t794 vp_p.t705 out_p.t890 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1674 out_p.t923 vp_p.t706 vdd1.t793 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1675 vdd1.t792 vp_p.t707 out_p.t889 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1676 vdd2.t801 vn_p.t698 out_n.t1063 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1677 out_n.t197 vn_n.t138 vss.t197 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1678 vdd1.t791 vp_p.t708 out_p.t880 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1679 vdd2.t800 vn_p.t699 out_n.t1062 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1680 vdd1.t790 vp_p.t709 out_p.t913 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1681 out_n.t1061 vn_p.t700 vdd2.t799 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1682 out_p.t879 vp_p.t710 vdd1.t789 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1683 vdd1.t788 vp_p.t711 out_p.t870 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1684 vdd2.t798 vn_p.t701 out_n.t1060 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1685 out_p.t903 vp_p.t712 vdd1.t787 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1686 vdd1.t786 vp_p.t713 out_p.t869 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1687 out_n.t1059 vn_p.t702 vdd2.t797 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1688 out_p.t1774 vp_n.t132 vss.t429 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1689 out_n.t1058 vn_p.t703 vdd2.t796 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1690 vdd2.t795 vn_p.t704 out_n.t1057 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1691 out_n.t1056 vn_p.t705 vdd2.t794 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1692 vss.t198 vn_n.t139 out_n.t198 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1693 vdd2.t793 vn_p.t706 out_n.t1055 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1694 out_n.t1054 vn_p.t707 vdd2.t792 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1695 vdd2.t791 vn_p.t708 out_n.t1053 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1696 vdd2.t790 vn_p.t709 out_n.t1052 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1697 out_n.t1051 vn_p.t710 vdd2.t789 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1698 vdd1.t785 vp_p.t714 out_p.t860 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1699 out_n.t1050 vn_p.t711 vdd2.t788 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1700 out_n.t1049 vn_p.t712 vdd2.t787 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1701 out_p.t893 vp_p.t715 vdd1.t784 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1702 vdd2.t786 vn_p.t713 out_n.t1048 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1703 out_p.t859 vp_p.t716 vdd1.t783 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1704 out_p.t850 vp_p.t717 vdd1.t782 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1705 vdd1.t781 vp_p.t718 out_p.t883 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1706 vdd2.t785 vn_p.t714 out_n.t1047 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1707 out_n.t1046 vn_p.t715 vdd2.t784 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1708 out_p.t849 vp_p.t719 vdd1.t780 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1709 out_n.t208 vn_n.t140 vss.t208 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1710 vdd2.t783 vn_p.t716 out_n.t1045 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1711 vdd2.t782 vn_p.t717 out_n.t1044 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1712 vss.t428 vp_n.t133 out_p.t1775 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1713 vdd2.t781 vn_p.t718 out_n.t1043 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1714 out_n.t1042 vn_p.t719 vdd2.t780 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1715 out_p.t840 vp_p.t720 vdd1.t779 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1716 out_p.t873 vp_p.t721 vdd1.t778 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1717 vdd1.t777 vp_p.t722 out_p.t839 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1718 vdd2.t779 vn_p.t720 out_n.t1041 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1719 out_p.t830 vp_p.t723 vdd1.t776 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1720 vdd2.t778 vn_p.t721 out_n.t1040 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1721 out_p.t863 vp_p.t724 vdd1.t775 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1722 out_p.t829 vp_p.t725 vdd1.t774 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1723 out_n.t209 vn_n.t141 vss.t209 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1724 vdd2.t777 vn_p.t722 out_n.t1039 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1725 vdd1.t773 vp_p.t726 out_p.t820 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1726 vss.t210 vn_n.t142 out_n.t210 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1727 out_n.t1038 vn_p.t723 vdd2.t776 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1728 vdd2.t775 vn_p.t724 out_n.t1037 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1729 vdd1.t772 vp_p.t727 out_p.t853 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1730 out_p.t1776 vp_n.t134 vss.t427 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1731 out_p.t819 vp_p.t728 vdd1.t771 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1732 out_p.t810 vp_p.t729 vdd1.t770 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1733 vdd1.t769 vp_p.t730 out_p.t843 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1734 vdd1.t768 vp_p.t731 out_p.t809 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1735 vdd1.t767 vp_p.t732 out_p.t800 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1736 vdd2.t774 vn_p.t725 out_n.t1036 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1737 vss.t426 vp_n.t135 out_p.t217 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1738 vdd1.t766 vp_p.t733 out_p.t833 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1739 out_p.t799 vp_p.t734 vdd1.t765 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1740 vss.t211 vn_n.t143 out_n.t211 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1741 out_n.t1035 vn_p.t726 vdd2.t773 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1742 out_n.t212 vn_n.t144 vss.t212 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1743 out_p.t790 vp_p.t735 vdd1.t764 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1744 out_p.t823 vp_p.t736 vdd1.t763 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1745 vdd1.t762 vp_p.t737 out_p.t789 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1746 out_n.t1034 vn_p.t727 vdd2.t772 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1747 out_n.t1033 vn_p.t728 vdd2.t771 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1748 out_n.t1032 vn_p.t729 vdd2.t770 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1749 out_n.t1031 vn_p.t730 vdd2.t769 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1750 vdd2.t768 vn_p.t731 out_n.t1030 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1751 out_n.t1029 vn_p.t732 vdd2.t767 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1752 out_n.t1028 vn_p.t733 vdd2.t766 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1753 out_n.t1027 vn_p.t734 vdd2.t765 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1754 out_p.t780 vp_p.t738 vdd1.t761 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1755 vdd2.t764 vn_p.t735 out_n.t1026 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1756 vdd2.t763 vn_p.t736 out_n.t1025 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1757 out_n.t1024 vn_p.t737 vdd2.t762 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1758 vss.t425 vp_n.t136 out_p.t218 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1759 vdd1.t760 vp_p.t739 out_p.t813 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1760 vdd2.t761 vn_p.t738 out_n.t1023 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1761 out_n.t1022 vn_p.t739 vdd2.t760 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1762 out_n.t1021 vn_p.t740 vdd2.t759 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1763 vdd2.t758 vn_p.t741 out_n.t1020 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1764 out_p.t779 vp_p.t740 vdd1.t759 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1765 out_p.t770 vp_p.t741 vdd1.t758 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1766 out_n.t44 vn_n.t145 vss.t44 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1767 vdd1.t757 vp_p.t742 out_p.t803 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1768 vdd1.t756 vp_p.t743 out_p.t769 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1769 out_p.t760 vp_p.t744 vdd1.t755 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1770 out_n.t1019 vn_p.t742 vdd2.t757 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1771 vdd1.t754 vp_p.t745 out_p.t793 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1772 out_n.t1018 vn_p.t743 vdd2.t756 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1773 vdd2.t755 vn_p.t744 out_n.t1017 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1774 out_p.t759 vp_p.t746 vdd1.t753 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1775 out_p.t750 vp_p.t747 vdd1.t752 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1776 vdd2.t754 vn_p.t745 out_n.t1016 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1777 out_n.t1015 vn_p.t746 vdd2.t753 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1778 vdd1.t751 vp_p.t748 out_p.t783 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1779 out_p.t749 vp_p.t749 vdd1.t750 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1780 out_p.t740 vp_p.t750 vdd1.t749 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1781 out_n.t1014 vn_p.t747 vdd2.t752 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1782 out_p.t219 vp_n.t137 vss.t424 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1783 out_n.t1013 vn_p.t748 vdd2.t751 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1784 vdd2.t750 vn_p.t749 out_n.t1012 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1785 out_p.t773 vp_p.t751 vdd1.t748 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1786 vdd1.t747 vp_p.t752 out_p.t739 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1787 out_p.t730 vp_p.t753 vdd1.t746 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1788 vdd1.t745 vp_p.t754 out_p.t763 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1789 vdd1.t744 vp_p.t755 out_p.t729 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1790 vdd1.t743 vp_p.t756 out_p.t720 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1791 out_p.t753 vp_p.t757 vdd1.t742 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1792 out_n.t1011 vn_p.t750 vdd2.t749 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1793 vdd2.t748 vn_p.t751 out_n.t1010 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1794 out_p.t220 vp_n.t138 vss.t423 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1795 out_p.t719 vp_p.t758 vdd1.t741 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1796 vss.t45 vn_n.t146 out_n.t45 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1797 out_n.t46 vn_n.t147 vss.t46 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1798 vss.t422 vp_n.t139 out_p.t221 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1799 out_p.t710 vp_p.t759 vdd1.t740 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1800 out_p.t743 vp_p.t760 vdd1.t739 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1801 vss.t47 vn_n.t148 out_n.t47 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1802 out_p.t709 vp_p.t761 vdd1.t738 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1803 out_p.t699 vp_p.t762 vdd1.t737 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1804 out_n.t1009 vn_p.t752 vdd2.t747 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1805 vss.t421 vp_n.t140 out_p.t222 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1806 vss.t420 vp_n.t141 out_p.t223 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1807 vdd1.t736 vp_p.t763 out_p.t733 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1808 out_p.t698 vp_p.t764 vdd1.t735 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1809 vdd2.t746 vn_p.t753 out_n.t1008 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1810 out_n.t1007 vn_p.t754 vdd2.t745 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1811 out_p.t224 vp_n.t142 vss.t419 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1812 out_p.t688 vp_p.t765 vdd1.t734 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1813 out_p.t723 vp_p.t766 vdd1.t733 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1814 vdd2.t744 vn_p.t755 out_n.t1006 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1815 out_n.t1005 vn_p.t756 vdd2.t743 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1816 out_n.t1004 vn_p.t757 vdd2.t742 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1817 vdd2.t741 vn_p.t758 out_n.t1003 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1818 out_n.t1002 vn_p.t759 vdd2.t740 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1819 vdd1.t732 vp_p.t767 out_p.t687 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1820 out_p.t677 vp_p.t768 vdd1.t731 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1821 vdd2.t739 vn_p.t760 out_n.t1001 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1822 out_n.t1000 vn_p.t761 vdd2.t738 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1823 vdd2.t737 vn_p.t762 out_n.t999 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1824 out_p.t225 vp_n.t143 vss.t418 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1825 out_n.t998 vn_p.t763 vdd2.t736 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1826 out_n.t997 vn_p.t764 vdd2.t735 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1827 out_n.t48 vn_n.t149 vss.t48 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1828 out_n.t996 vn_p.t765 vdd2.t734 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1829 vdd2.t733 vn_p.t766 out_n.t995 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1830 out_p.t226 vp_n.t144 vss.t417 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1831 out_n.t247 vn_n.t150 vss.t247 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1832 out_p.t227 vp_n.t145 vss.t416 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1833 vss.t248 vn_n.t151 out_n.t248 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1834 vdd2.t732 vn_p.t767 out_n.t994 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1835 vdd2.t731 vn_p.t768 out_n.t993 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1836 out_n.t992 vn_p.t769 vdd2.t730 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1837 vdd2.t729 vn_p.t770 out_n.t991 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1838 out_n.t990 vn_p.t771 vdd2.t728 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1839 vdd2.t727 vn_p.t772 out_n.t989 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1840 out_n.t988 vn_p.t773 vdd2.t726 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1841 vdd1.t730 vp_p.t769 out_p.t713 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1842 vss.t249 vn_n.t152 out_n.t249 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1843 out_p.t702 vp_p.t770 vdd1.t729 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1844 out_p.t676 vp_p.t771 vdd1.t728 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1845 out_p.t667 vp_p.t772 vdd1.t727 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1846 out_p.t703 vp_p.t773 vdd1.t726 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1847 out_p.t691 vp_p.t774 vdd1.t725 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1848 vdd1.t724 vp_p.t775 out_p.t666 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1849 vdd1.t723 vp_p.t776 out_p.t656 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1850 out_p.t692 vp_p.t777 vdd1.t722 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1851 out_n.t987 vn_p.t774 vdd2.t725 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1852 vdd1.t721 vp_p.t778 out_p.t680 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1853 out_n.t986 vn_p.t775 vdd2.t724 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1854 out_n.t985 vn_p.t776 vdd2.t723 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1855 vdd1.t720 vp_p.t779 out_p.t655 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1856 vdd1.t719 vp_p.t780 out_p.t645 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1857 vdd2.t722 vn_p.t777 out_n.t984 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1858 out_n.t983 vn_p.t778 vdd2.t721 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1859 out_n.t250 vn_n.t153 vss.t250 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1860 out_p.t681 vp_p.t781 vdd1.t718 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1861 vdd2.t720 vn_p.t779 out_n.t982 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1862 out_n.t981 vn_p.t780 vdd2.t719 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1863 out_p.t671 vp_p.t782 vdd1.t717 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1864 vdd2.t718 vn_p.t781 out_n.t980 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1865 out_n.t979 vn_p.t782 vdd2.t717 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1866 out_p.t660 vp_p.t783 vdd1.t716 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1867 vdd1.t715 vp_p.t784 out_p.t647 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1868 out_p.t661 vp_p.t785 vdd1.t714 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1869 vdd2.t716 vn_p.t783 out_n.t978 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1870 vdd1.t713 vp_p.t786 out_p.t637 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1871 out_p.t950 vp_p.t787 vdd1.t712 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1872 vdd1.t711 vp_p.t788 out_p.t951 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1873 vss.t415 vp_n.t146 out_p.t228 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1874 out_p.t229 vp_n.t147 vss.t414 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1875 out_p.t962 vp_p.t789 vdd1.t710 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1876 vdd2.t715 vn_p.t784 out_n.t977 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1877 out_n.t976 vn_p.t785 vdd2.t714 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1878 vdd1.t709 vp_p.t790 out_p.t991 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1879 vdd2.t713 vn_p.t786 out_n.t975 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1880 vdd2.t712 vn_p.t787 out_n.t974 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1881 vdd2.t711 vn_p.t788 out_n.t973 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1882 vdd2.t710 vn_p.t789 out_n.t972 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1883 out_p.t998 vp_p.t791 vdd1.t708 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1884 vdd1.t707 vp_p.t792 out_p.t1004 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1885 vdd1.t706 vp_p.t793 out_p.t1010 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1886 vdd2.t709 vn_p.t790 out_n.t971 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1887 out_p.t1016 vp_p.t794 vdd1.t705 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1888 out_p.t1023 vp_p.t795 vdd1.t704 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1889 vdd2.t708 vn_p.t791 out_n.t970 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1890 vss.t413 vp_n.t148 out_p.t230 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1891 vdd2.t707 vn_p.t792 out_n.t969 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1892 vdd1.t703 vp_p.t796 out_p.t262 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1893 out_n.t968 vn_p.t793 vdd2.t706 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1894 vdd1.t702 vp_p.t797 out_p.t985 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1895 out_n.t967 vn_p.t794 vdd2.t705 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1896 vdd2.t704 vn_p.t795 out_n.t966 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1897 out_n.t251 vn_n.t154 vss.t251 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1898 vss.t150 vn_n.t155 out_n.t150 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1899 vdd2.t703 vn_p.t796 out_n.t965 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1900 out_p.t231 vp_n.t149 vss.t412 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1901 out_n.t964 vn_p.t797 vdd2.t702 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1902 out_n.t963 vn_p.t798 vdd2.t701 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1903 vdd2.t700 vn_p.t799 out_n.t962 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1904 out_n.t961 vn_p.t800 vdd2.t699 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1905 out_n.t960 vn_p.t801 vdd2.t698 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1906 vdd1.t701 vp_p.t798 out_p.t1017 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1907 out_n.t959 vn_p.t802 vdd2.t697 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1908 out_n.t958 vn_p.t803 vdd2.t696 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1909 vss.t411 vp_n.t150 out_p.t232 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1910 out_n.t151 vn_n.t156 vss.t151 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1911 vss.t152 vn_n.t157 out_n.t152 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1912 out_p.t1022 vp_p.t799 vdd1.t700 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1913 out_p.t1025 vp_p.t800 vdd1.t699 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1914 out_n.t957 vn_p.t804 vdd2.t695 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1915 out_p.t995 vp_p.t801 vdd1.t698 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1916 vss.t153 vn_n.t158 out_n.t153 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1917 vdd1.t697 vp_p.t802 out_p.t966 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1918 vdd1.t696 vp_p.t803 out_p.t973 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1919 vdd2.t694 vn_p.t805 out_n.t956 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1920 vdd1.t695 vp_p.t804 out_p.t979 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1921 vdd1.t694 vp_p.t805 out_p.t1014 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1922 out_n.t154 vn_n.t159 vss.t154 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1923 out_p.t992 vp_p.t806 vdd1.t693 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1924 vdd2.t693 vn_p.t806 out_n.t955 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1925 vdd2.t692 vn_p.t807 out_n.t954 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1926 vdd1.t692 vp_p.t807 out_p.t996 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1927 out_n.t953 vn_p.t808 vdd2.t691 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1928 out_p.t999 vp_p.t808 vdd1.t691 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1929 vdd1.t690 vp_p.t809 out_p.t1002 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1930 vdd2.t690 vn_p.t809 out_n.t952 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1931 vdd2.t689 vn_p.t810 out_n.t951 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1932 out_p.t1005 vp_p.t810 vdd1.t689 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1933 out_p.t1008 vp_p.t811 vdd1.t688 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1934 vdd1.t687 vp_p.t812 out_p.t1011 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1935 vdd2.t688 vn_p.t811 out_n.t950 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1936 vdd1.t686 vp_p.t813 out_p.t989 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1937 out_n.t164 vn_n.t160 vss.t164 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1938 vdd2.t687 vn_p.t812 out_n.t949 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1939 vdd1.t685 vp_p.t814 out_p.t968 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1940 out_p.t971 vp_p.t815 vdd1.t684 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1941 out_n.t948 vn_p.t813 vdd2.t686 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1942 vdd2.t685 vn_p.t814 out_n.t947 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1943 out_p.t233 vp_n.t151 vss.t410 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1944 out_p.t974 vp_p.t816 vdd1.t683 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1945 out_p.t977 vp_p.t817 vdd1.t682 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1946 out_n.t946 vn_p.t815 vdd2.t684 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1947 vdd2.t683 vn_p.t816 out_n.t945 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1948 vss.t409 vp_n.t152 out_p.t234 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1949 vdd1.t681 vp_p.t818 out_p.t980 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1950 out_p.t235 vp_n.t153 vss.t408 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1951 out_n.t944 vn_p.t817 vdd2.t682 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1952 vdd1.t680 vp_p.t819 out_p.t983 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1953 out_p.t986 vp_p.t820 vdd1.t679 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1954 out_p.t236 vp_n.t154 vss.t407 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1955 vdd2.t681 vn_p.t818 out_n.t943 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1956 vss.t165 vn_n.t161 out_n.t165 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1957 out_n.t942 vn_p.t819 vdd2.t680 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1958 out_n.t941 vn_p.t820 vdd2.t679 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1959 vdd1.t678 vp_p.t821 out_p.t964 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1960 vdd1.t677 vp_p.t822 out_p.t266 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1961 out_n.t940 vn_p.t821 vdd2.t678 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1962 out_p.t197 vp_n.t155 vss.t406 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1963 out_n.t939 vn_p.t822 vdd2.t677 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1964 vdd2.t676 vn_p.t823 out_n.t938 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1965 vdd1.t676 vp_p.t823 out_p.t273 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1966 vdd2.t675 vn_p.t824 out_n.t937 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1967 out_p.t268 vp_p.t824 vdd1.t675 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1968 out_p.t270 vp_p.t825 vdd1.t674 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1969 out_n.t166 vn_n.t162 vss.t166 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1970 vdd2.t674 vn_p.t825 out_n.t936 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1971 out_n.t935 vn_p.t826 vdd2.t673 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1972 vdd2.t672 vn_p.t827 out_n.t934 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1973 vss.t405 vp_n.t156 out_p.t198 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1974 out_p.t199 vp_n.t157 vss.t404 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1975 vdd2.t671 vn_p.t828 out_n.t933 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1976 out_n.t932 vn_p.t829 vdd2.t670 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1977 out_p.t257 vp_p.t826 vdd1.t673 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1978 vdd2.t669 vn_p.t830 out_n.t931 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1979 vdd2.t668 vn_p.t831 out_n.t930 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1980 out_n.t167 vn_n.t163 vss.t167 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1981 vss.t403 vp_n.t158 out_p.t200 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1982 out_p.t269 vp_p.t827 vdd1.t672 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1983 out_n.t929 vn_p.t832 vdd2.t667 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1984 vdd2.t666 vn_p.t833 out_n.t928 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1985 vdd2.t665 vn_p.t834 out_n.t927 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1986 out_n.t926 vn_p.t835 vdd2.t664 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1987 out_p.t1020 vp_p.t828 vdd1.t671 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1988 vdd2.t663 vn_p.t836 out_n.t925 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1989 vdd1.t670 vp_p.t829 out_p.t259 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1990 out_p.t263 vp_p.t830 vdd1.t669 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1991 vdd1.t668 vp_p.t831 out_p.t260 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1992 out_p.t271 vp_p.t832 vdd1.t667 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1993 out_p.t272 vp_p.t833 vdd1.t666 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1994 out_p.t261 vp_p.t834 vdd1.t665 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1995 out_p.t264 vp_p.t835 vdd1.t664 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1996 vdd1.t663 vp_p.t836 out_p.t265 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1997 vdd1.t662 vp_p.t837 out_p.t258 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1998 out_p.t1756 vp_p.t838 vdd1.t661 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1999 vss.t168 vn_n.t164 out_n.t168 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2000 out_n.t169 vn_n.t165 vss.t169 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2001 out_n.t924 vn_p.t837 vdd2.t662 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2002 out_p.t201 vp_n.t159 vss.t402 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2003 vdd1.t660 vp_p.t839 out_p.t1755 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2004 out_n.t923 vn_p.t838 vdd2.t661 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2005 out_n.t922 vn_p.t839 vdd2.t660 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2006 vdd2.t659 vn_p.t840 out_n.t921 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2007 vdd1.t659 vp_p.t840 out_p.t1754 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2008 out_n.t920 vn_p.t841 vdd2.t658 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2009 out_p.t1753 vp_p.t841 vdd1.t658 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2010 out_p.t1752 vp_p.t842 vdd1.t657 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2011 vdd1.t656 vp_p.t843 out_p.t1751 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2012 vdd1.t655 vp_p.t844 out_p.t1750 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2013 out_n.t919 vn_p.t842 vdd2.t657 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2014 out_n.t918 vn_p.t843 vdd2.t656 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2015 out_p.t1749 vp_p.t845 vdd1.t654 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2016 vdd1.t653 vp_p.t846 out_p.t1748 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2017 vdd2.t655 vn_p.t844 out_n.t917 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2018 out_n.t916 vn_p.t845 vdd2.t654 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2019 vdd1.t652 vp_p.t847 out_p.t1747 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2020 vdd1.t651 vp_p.t848 out_p.t1746 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2021 vdd1.t650 vp_p.t849 out_p.t1745 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2022 vss.t66 vn_n.t166 out_n.t66 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2023 vdd2.t653 vn_p.t846 out_n.t915 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2024 vdd2.t652 vn_p.t847 out_n.t914 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2025 out_p.t1744 vp_p.t850 vdd1.t649 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2026 out_p.t1743 vp_p.t851 vdd1.t648 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2027 out_n.t67 vn_n.t167 vss.t67 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2028 vss.t401 vp_n.t160 out_p.t202 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2029 vdd2.t651 vn_p.t848 out_n.t913 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2030 vdd2.t650 vn_p.t849 out_n.t912 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2031 out_n.t911 vn_p.t850 vdd2.t649 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2032 out_n.t910 vn_p.t851 vdd2.t648 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2033 vdd1.t647 vp_p.t852 out_p.t1742 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2034 vdd2.t647 vn_p.t852 out_n.t909 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2035 vdd2.t646 vn_p.t853 out_n.t908 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2036 vdd1.t646 vp_p.t853 out_p.t1741 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2037 out_p.t1740 vp_p.t854 vdd1.t645 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2038 out_p.t203 vp_n.t161 vss.t400 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2039 vss.t399 vp_n.t162 out_p.t204 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2040 out_n.t907 vn_p.t854 vdd2.t645 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2041 vdd1.t644 vp_p.t855 out_p.t1739 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2042 out_n.t906 vn_p.t855 vdd2.t644 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2043 vdd2.t643 vn_p.t856 out_n.t905 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2044 vdd2.t642 vn_p.t857 out_n.t904 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2045 vdd1.t643 vp_p.t856 out_p.t1738 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2046 vdd2.t641 vn_p.t858 out_n.t903 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2047 out_n.t902 vn_p.t859 vdd2.t640 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2048 out_n.t901 vn_p.t860 vdd2.t639 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2049 out_n.t900 vn_p.t861 vdd2.t638 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2050 vdd2.t637 vn_p.t862 out_n.t899 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2051 vss.t68 vn_n.t168 out_n.t68 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2052 vdd1.t642 vp_p.t857 out_p.t1737 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2053 vdd1.t641 vp_p.t858 out_p.t1736 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2054 out_p.t1735 vp_p.t859 vdd1.t640 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2055 out_p.t1734 vp_p.t860 vdd1.t639 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2056 out_p.t1733 vp_p.t861 vdd1.t638 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2057 vdd1.t637 vp_p.t862 out_p.t1732 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2058 vdd1.t636 vp_p.t863 out_p.t1731 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2059 out_n.t898 vn_p.t863 vdd2.t636 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2060 vdd2.t635 vn_p.t864 out_n.t897 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2061 out_p.t1730 vp_p.t864 vdd1.t635 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2062 out_p.t1729 vp_p.t865 vdd1.t634 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2063 out_n.t896 vn_p.t865 vdd2.t634 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2064 vdd1.t633 vp_p.t866 out_p.t1728 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2065 vdd1.t632 vp_p.t867 out_p.t1727 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2066 vdd2.t633 vn_p.t866 out_n.t895 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2067 out_n.t894 vn_p.t867 vdd2.t632 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2068 out_p.t1726 vp_p.t868 vdd1.t631 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2069 vdd1.t630 vp_p.t869 out_p.t1725 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2070 out_p.t1724 vp_p.t870 vdd1.t629 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2071 out_n.t893 vn_p.t868 vdd2.t631 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2072 vss.t398 vp_n.t163 out_p.t205 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2073 out_p.t1723 vp_p.t871 vdd1.t628 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2074 vdd2.t630 vn_p.t869 out_n.t892 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2075 out_p.t1722 vp_p.t872 vdd1.t627 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2076 vdd2.t629 vn_p.t870 out_n.t891 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2077 vdd1.t626 vp_p.t873 out_p.t1721 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2078 out_n.t69 vn_n.t169 vss.t69 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2079 vss.t70 vn_n.t170 out_n.t70 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2080 vdd1.t625 vp_p.t874 out_p.t1720 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2081 out_p.t1719 vp_p.t875 vdd1.t624 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2082 out_n.t71 vn_n.t171 vss.t71 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2083 vdd1.t623 vp_p.t876 out_p.t1718 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2084 vdd1.t622 vp_p.t877 out_p.t1717 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2085 vdd2.t628 vn_p.t871 out_n.t890 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2086 out_p.t1716 vp_p.t878 vdd1.t621 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2087 vdd2.t627 vn_p.t872 out_n.t889 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2088 out_n.t888 vn_p.t873 vdd2.t626 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2089 out_n.t887 vn_p.t874 vdd2.t625 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2090 vdd2.t624 vn_p.t875 out_n.t886 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2091 out_n.t885 vn_p.t876 vdd2.t623 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2092 vdd1.t620 vp_p.t879 out_p.t1715 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2093 vdd2.t622 vn_p.t877 out_n.t884 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2094 out_p.t206 vp_n.t164 vss.t397 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2095 out_p.t1714 vp_p.t880 vdd1.t619 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2096 out_n.t883 vn_p.t878 vdd2.t621 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2097 out_p.t1713 vp_p.t881 vdd1.t618 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2098 vdd1.t617 vp_p.t882 out_p.t1712 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2099 vdd1.t616 vp_p.t883 out_p.t1711 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2100 vdd1.t615 vp_p.t884 out_p.t1710 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2101 vdd2.t620 vn_p.t879 out_n.t882 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2102 out_n.t881 vn_p.t880 vdd2.t619 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2103 out_n.t880 vn_p.t881 vdd2.t618 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2104 vss.t396 vp_n.t165 out_p.t207 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2105 out_p.t1709 vp_p.t885 vdd1.t614 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2106 vdd2.t617 vn_p.t882 out_n.t879 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2107 vdd2.t616 vn_p.t883 out_n.t878 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2108 out_p.t208 vp_n.t166 vss.t395 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2109 vss.t394 vp_n.t167 out_p.t209 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2110 out_n.t877 vn_p.t884 vdd2.t615 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2111 vdd1.t613 vp_p.t886 out_p.t1708 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2112 out_n.t876 vn_p.t885 vdd2.t614 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2113 vdd2.t613 vn_p.t886 out_n.t875 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2114 out_n.t874 vn_p.t887 vdd2.t612 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2115 vdd1.t612 vp_p.t887 out_p.t1707 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2116 vss.t393 vp_n.t168 out_p.t210 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2117 vdd2.t611 vn_p.t888 out_n.t873 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2118 vdd1.t611 vp_p.t888 out_p.t1706 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2119 vdd1.t610 vp_p.t889 out_p.t1705 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2120 out_p.t1704 vp_p.t890 vdd1.t609 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2121 out_p.t1703 vp_p.t891 vdd1.t608 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2122 out_p.t1702 vp_p.t892 vdd1.t607 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2123 out_p.t1701 vp_p.t893 vdd1.t606 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2124 out_p.t1700 vp_p.t894 vdd1.t605 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2125 vdd2.t610 vn_p.t889 out_n.t872 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2126 out_n.t871 vn_p.t890 vdd2.t609 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2127 out_n.t870 vn_p.t891 vdd2.t608 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2128 out_p.t211 vp_n.t169 vss.t392 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2129 out_p.t1699 vp_p.t895 vdd1.t604 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2130 vdd2.t607 vn_p.t892 out_n.t869 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2131 vdd1.t603 vp_p.t896 out_p.t1698 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2132 vdd1.t602 vp_p.t897 out_p.t1697 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2133 vdd1.t601 vp_p.t898 out_p.t1696 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2134 out_p.t1695 vp_p.t899 vdd1.t600 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2135 vdd1.t599 vp_p.t900 out_p.t1694 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2136 vdd1.t598 vp_p.t901 out_p.t1693 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2137 vdd1.t597 vp_p.t902 out_p.t1692 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2138 out_p.t212 vp_n.t170 vss.t391 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2139 out_n.t0 vn_n.t172 vss.t0 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2140 vss.t1 vn_n.t173 out_n.t1 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2141 out_n.t868 vn_p.t893 vdd2.t606 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2142 vdd2.t605 vn_p.t894 out_n.t867 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2143 out_p.t213 vp_n.t171 vss.t390 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2144 vdd1.t596 vp_p.t903 out_p.t1691 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2145 vdd1.t595 vp_p.t904 out_p.t1690 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2146 vdd2.t604 vn_p.t895 out_n.t866 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2147 vdd1.t594 vp_p.t905 out_p.t1689 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2148 out_p.t1688 vp_p.t906 vdd1.t593 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2149 vdd2.t603 vn_p.t896 out_n.t865 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2150 out_n.t864 vn_p.t897 vdd2.t602 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2151 out_n.t863 vn_p.t898 vdd2.t601 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2152 out_n.t862 vn_p.t899 vdd2.t600 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2153 out_n.t861 vn_p.t900 vdd2.t599 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2154 out_n.t860 vn_p.t901 vdd2.t598 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2155 vss.t389 vp_n.t172 out_p.t214 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2156 vdd1.t592 vp_p.t907 out_p.t1687 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2157 out_n.t859 vn_p.t902 vdd2.t597 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2158 vdd1.t591 vp_p.t908 out_p.t1686 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2159 out_n.t858 vn_p.t903 vdd2.t596 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2160 out_n.t857 vn_p.t904 vdd2.t595 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2161 vss.t388 vp_n.t173 out_p.t215 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2162 vss.t2 vn_n.t174 out_n.t2 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2163 vdd2.t594 vn_p.t905 out_n.t856 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2164 out_p.t1685 vp_p.t909 vdd1.t590 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2165 vdd2.t593 vn_p.t906 out_n.t855 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2166 out_n.t3 vn_n.t175 vss.t3 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2167 vdd2.t592 vn_p.t907 out_n.t854 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2168 out_n.t853 vn_p.t908 vdd2.t591 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2169 vdd2.t590 vn_p.t909 out_n.t852 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2170 vdd2.t589 vn_p.t910 out_n.t851 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2171 out_p.t1684 vp_p.t910 vdd1.t589 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2172 vdd2.t588 vn_p.t911 out_n.t850 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2173 vdd2.t587 vn_p.t912 out_n.t849 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2174 vdd1.t588 vp_p.t911 out_p.t1683 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2175 out_p.t1682 vp_p.t912 vdd1.t587 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2176 vdd2.t586 vn_p.t913 out_n.t848 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2177 vss.t4 vn_n.t176 out_n.t4 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2178 out_n.t5 vn_n.t177 vss.t5 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2179 vdd2.t585 vn_p.t914 out_n.t847 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2180 vdd1.t586 vp_p.t913 out_p.t1681 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2181 out_p.t1680 vp_p.t914 vdd1.t585 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2182 vdd1.t584 vp_p.t915 out_p.t1679 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2183 out_n.t846 vn_p.t915 vdd2.t584 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2184 vdd2.t583 vn_p.t916 out_n.t845 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2185 out_n.t844 vn_p.t917 vdd2.t582 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2186 out_p.t1678 vp_p.t916 vdd1.t583 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2187 vdd2.t581 vn_p.t918 out_n.t843 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2188 out_p.t1677 vp_p.t917 vdd1.t582 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2189 vdd1.t581 vp_p.t918 out_p.t1676 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2190 out_p.t1675 vp_p.t919 vdd1.t580 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2191 vss.t570 vn_n.t178 out_n.t1770 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2192 out_n.t842 vn_p.t919 vdd2.t580 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2193 vdd1.t579 vp_p.t920 out_p.t1674 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2194 vdd1.t578 vp_p.t921 out_p.t1673 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2195 out_n.t841 vn_p.t920 vdd2.t579 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2196 vdd1.t577 vp_p.t922 out_p.t1672 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2197 vdd1.t576 vp_p.t923 out_p.t1671 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2198 vdd1.t575 vp_p.t924 out_p.t1670 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2199 out_p.t216 vp_n.t174 vss.t387 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2200 out_p.t1669 vp_p.t925 vdd1.t574 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2201 out_n.t840 vn_p.t921 vdd2.t578 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2202 vdd2.t577 vn_p.t922 out_n.t839 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2203 vss.t571 vn_n.t179 out_n.t1771 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2204 out_n.t1772 vn_n.t180 vss.t572 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2205 vss.t386 vp_n.t175 out_p.t64 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2206 vdd1.t573 vp_p.t926 out_p.t1668 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2207 out_p.t1667 vp_p.t927 vdd1.t572 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2208 out_n.t838 vn_p.t923 vdd2.t576 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2209 out_p.t1666 vp_p.t928 vdd1.t571 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2210 out_p.t1665 vp_p.t929 vdd1.t570 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2211 vdd1.t569 vp_p.t930 out_p.t1664 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2212 out_n.t837 vn_p.t924 vdd2.t575 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2213 vdd2.t574 vn_p.t925 out_n.t836 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2214 out_n.t835 vn_p.t926 vdd2.t573 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2215 vdd2.t572 vn_p.t927 out_n.t834 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2216 vdd1.t568 vp_p.t931 out_p.t1663 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2217 vdd2.t571 vn_p.t928 out_n.t833 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2218 out_n.t832 vn_p.t929 vdd2.t570 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2219 out_p.t1662 vp_p.t932 vdd1.t567 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2220 vdd2.t569 vn_p.t930 out_n.t831 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2221 out_n.t830 vn_p.t931 vdd2.t568 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2222 vdd2.t567 vn_p.t932 out_n.t829 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2223 vdd2.t566 vn_p.t933 out_n.t828 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2224 out_n.t827 vn_p.t934 vdd2.t565 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2225 vdd2.t564 vn_p.t935 out_n.t826 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2226 out_n.t1773 vn_n.t181 vss.t573 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2227 vss.t385 vp_n.t176 out_p.t65 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2228 vdd2.t563 vn_p.t936 out_n.t825 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2229 vdd2.t562 vn_p.t937 out_n.t824 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2230 vdd1.t566 vp_p.t933 out_p.t1661 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2231 out_n.t823 vn_p.t938 vdd2.t561 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2232 out_p.t66 vp_n.t177 vss.t384 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2233 out_n.t822 vn_p.t939 vdd2.t560 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2234 out_n.t821 vn_p.t940 vdd2.t559 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2235 vdd2.t558 vn_p.t941 out_n.t820 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2236 vss.t574 vn_n.t182 out_n.t1774 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2237 out_n.t1775 vn_n.t183 vss.t575 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2238 out_n.t819 vn_p.t942 vdd2.t557 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2239 vdd1.t565 vp_p.t934 out_p.t1660 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2240 out_p.t1659 vp_p.t935 vdd1.t564 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2241 vdd1.t563 vp_p.t936 out_p.t1658 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2242 vdd1.t562 vp_p.t937 out_p.t1657 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2243 out_n.t818 vn_p.t943 vdd2.t556 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2244 vdd2.t555 vn_p.t944 out_n.t817 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2245 out_p.t1656 vp_p.t938 vdd1.t561 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2246 out_p.t1655 vp_p.t939 vdd1.t560 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2247 out_p.t1654 vp_p.t940 vdd1.t559 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2248 vdd1.t558 vp_p.t941 out_p.t1653 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2249 out_n.t816 vn_p.t945 vdd2.t554 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2250 out_p.t1652 vp_p.t942 vdd1.t557 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2251 vss.t129 vn_n.t184 out_n.t129 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2252 out_n.t815 vn_p.t946 vdd2.t553 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2253 vdd1.t556 vp_p.t943 out_p.t1651 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2254 vdd2.t552 vn_p.t947 out_n.t814 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2255 vdd2.t551 vn_p.t948 out_n.t813 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2256 out_p.t1650 vp_p.t944 vdd1.t555 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2257 vdd2.t550 vn_p.t949 out_n.t812 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2258 vdd1.t554 vp_p.t945 out_p.t1649 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2259 out_n.t811 vn_p.t950 vdd2.t549 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2260 out_p.t1648 vp_p.t946 vdd1.t553 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2261 vss.t383 vp_n.t178 out_p.t67 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2262 vdd1.t552 vp_p.t947 out_p.t1647 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2263 out_n.t130 vn_n.t185 vss.t130 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2264 out_n.t131 vn_n.t186 vss.t131 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2265 out_p.t1646 vp_p.t948 vdd1.t551 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2266 out_p.t1645 vp_p.t949 vdd1.t550 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2267 vdd1.t549 vp_p.t950 out_p.t1644 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2268 vss.t132 vn_n.t187 out_n.t132 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2269 out_n.t810 vn_p.t951 vdd2.t548 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2270 out_p.t1643 vp_p.t951 vdd1.t548 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2271 out_p.t1642 vp_p.t952 vdd1.t547 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2272 out_p.t1641 vp_p.t953 vdd1.t546 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2273 vdd1.t545 vp_p.t954 out_p.t1640 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2274 out_n.t133 vn_n.t188 vss.t133 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2275 vdd2.t547 vn_p.t952 out_n.t809 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2276 vss.t382 vp_n.t179 out_p.t68 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2277 vdd1.t544 vp_p.t955 out_p.t1639 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2278 vdd2.t546 vn_p.t953 out_n.t808 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2279 out_p.t69 vp_n.t180 vss.t381 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2280 vdd1.t543 vp_p.t956 out_p.t1638 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2281 out_p.t1637 vp_p.t957 vdd1.t542 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2282 vdd2.t545 vn_p.t954 out_n.t807 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2283 out_n.t806 vn_p.t955 vdd2.t544 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2284 vdd2.t543 vn_p.t956 out_n.t805 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2285 vdd2.t542 vn_p.t957 out_n.t804 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2286 vdd1.t541 vp_p.t958 out_p.t1636 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2287 vdd2.t541 vn_p.t958 out_n.t803 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2288 out_n.t802 vn_p.t959 vdd2.t540 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2289 vss.t380 vp_n.t181 out_p.t70 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2290 vdd1.t540 vp_p.t959 out_p.t1635 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2291 vdd2.t539 vn_p.t960 out_n.t801 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2292 out_p.t1634 vp_p.t960 vdd1.t539 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2293 out_n.t800 vn_p.t961 vdd2.t538 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2294 vdd2.t537 vn_p.t962 out_n.t799 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2295 vdd1.t538 vp_p.t961 out_p.t1633 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2296 out_n.t798 vn_p.t963 vdd2.t536 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2297 vdd2.t535 vn_p.t964 out_n.t797 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2298 out_n.t796 vn_p.t965 vdd2.t534 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2299 vss.t134 vn_n.t189 out_n.t134 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2300 out_n.t795 vn_p.t966 vdd2.t533 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2301 out_n.t794 vn_p.t967 vdd2.t532 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2302 vss.t379 vp_n.t182 out_p.t71 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2303 out_p.t72 vp_n.t183 vss.t378 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2304 vss.t24 vn_n.t190 out_n.t24 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2305 out_n.t793 vn_p.t968 vdd2.t531 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2306 out_n.t792 vn_p.t969 vdd2.t530 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2307 vdd2.t529 vn_p.t970 out_n.t791 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2308 vss.t377 vp_n.t184 out_p.t73 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2309 out_n.t790 vn_p.t971 vdd2.t528 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2310 out_n.t789 vn_p.t972 vdd2.t527 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2311 out_n.t25 vn_n.t191 vss.t25 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2312 vss.t26 vn_n.t192 out_n.t26 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2313 vdd2.t526 vn_p.t973 out_n.t788 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2314 out_p.t1632 vp_p.t962 vdd1.t537 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2315 vdd1.t536 vp_p.t963 out_p.t1631 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2316 out_p.t1630 vp_p.t964 vdd1.t535 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2317 out_p.t1629 vp_p.t965 vdd1.t534 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2318 vdd2.t525 vn_p.t974 out_n.t787 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2319 out_n.t786 vn_p.t975 vdd2.t524 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2320 out_p.t1628 vp_p.t966 vdd1.t533 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2321 vdd1.t532 vp_p.t967 out_p.t1627 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2322 vdd1.t531 vp_p.t968 out_p.t1626 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2323 out_n.t785 vn_p.t976 vdd2.t523 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2324 vdd1.t530 vp_p.t969 out_p.t1625 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2325 vdd1.t529 vp_p.t970 out_p.t1624 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2326 out_p.t1623 vp_p.t971 vdd1.t528 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2327 vdd1.t527 vp_p.t972 out_p.t1622 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2328 out_p.t1621 vp_p.t973 vdd1.t526 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2329 vdd1.t525 vp_p.t974 out_p.t1620 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2330 vdd2.t522 vn_p.t977 out_n.t784 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2331 out_n.t27 vn_n.t193 vss.t27 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2332 out_n.t783 vn_p.t978 vdd2.t521 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2333 vdd2.t520 vn_p.t979 out_n.t782 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2334 out_n.t28 vn_n.t194 vss.t28 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2335 out_p.t1619 vp_p.t975 vdd1.t524 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2336 vdd1.t523 vp_p.t976 out_p.t1618 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2337 out_p.t1617 vp_p.t977 vdd1.t522 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2338 out_n.t781 vn_p.t980 vdd2.t519 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2339 out_n.t780 vn_p.t981 vdd2.t518 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2340 out_p.t1616 vp_p.t978 vdd1.t521 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2341 vdd1.t520 vp_p.t979 out_p.t1615 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2342 vss.t29 vn_n.t195 out_n.t29 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2343 vdd2.t517 vn_p.t982 out_n.t779 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2344 out_p.t1614 vp_p.t980 vdd1.t519 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2345 vdd2.t516 vn_p.t983 out_n.t778 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2346 out_n.t777 vn_p.t984 vdd2.t515 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2347 vdd1.t518 vp_p.t981 out_p.t1613 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2348 vdd2.t514 vn_p.t985 out_n.t776 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2349 vdd2.t513 vn_p.t986 out_n.t775 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2350 vdd1.t517 vp_p.t982 out_p.t1612 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2351 vdd1.t516 vp_p.t983 out_p.t1611 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2352 out_p.t1610 vp_p.t984 vdd1.t515 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2353 vdd1.t514 vp_p.t985 out_p.t1609 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2354 out_p.t1608 vp_p.t986 vdd1.t513 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2355 out_n.t774 vn_p.t987 vdd2.t512 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2356 out_p.t74 vp_n.t185 vss.t376 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2357 vss.t375 vp_n.t186 out_p.t75 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2358 vdd1.t512 vp_p.t987 out_p.t1607 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2359 out_n.t773 vn_p.t988 vdd2.t511 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2360 vdd2.t510 vn_p.t989 out_n.t772 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2361 out_p.t1606 vp_p.t988 vdd1.t511 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2362 out_n.t771 vn_p.t990 vdd2.t509 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2363 out_n.t770 vn_p.t991 vdd2.t508 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2364 out_p.t1605 vp_p.t989 vdd1.t510 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2365 vdd1.t509 vp_p.t990 out_p.t1604 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2366 out_p.t1603 vp_p.t991 vdd1.t508 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2367 vss.t144 vn_n.t196 out_n.t144 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2368 vdd2.t507 vn_p.t992 out_n.t769 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2369 out_n.t768 vn_p.t993 vdd2.t506 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2370 vss.t145 vn_n.t197 out_n.t145 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2371 out_p.t1602 vp_p.t992 vdd1.t507 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2372 out_p.t1601 vp_p.t993 vdd1.t506 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2373 out_n.t767 vn_p.t994 vdd2.t505 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2374 out_n.t766 vn_p.t995 vdd2.t504 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2375 vdd2.t503 vn_p.t996 out_n.t765 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2376 out_n.t764 vn_p.t997 vdd2.t502 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2377 vdd2.t501 vn_p.t998 out_n.t763 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2378 out_n.t762 vn_p.t999 vdd2.t500 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2379 out_p.t76 vp_n.t187 vss.t374 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2380 vss.t373 vp_n.t188 out_p.t77 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2381 out_n.t146 vn_n.t198 vss.t146 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2382 out_n.t147 vn_n.t199 vss.t147 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2383 vdd2.t499 vn_p.t1000 out_n.t761 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2384 out_n.t760 vn_p.t1001 vdd2.t498 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2385 out_p.t1600 vp_p.t994 vdd1.t505 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2386 out_p.t78 vp_n.t189 vss.t372 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2387 vdd2.t497 vn_p.t1002 out_n.t759 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2388 out_p.t1599 vp_p.t995 vdd1.t504 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2389 vdd2.t496 vn_p.t1003 out_n.t758 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2390 out_n.t757 vn_p.t1004 vdd2.t495 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2391 out_p.t1598 vp_p.t996 vdd1.t503 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2392 vdd1.t502 vp_p.t997 out_p.t1597 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2393 vdd1.t501 vp_p.t998 out_p.t1596 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2394 vdd1.t500 vp_p.t999 out_p.t1595 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2395 out_n.t756 vn_p.t1005 vdd2.t494 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2396 vdd1.t499 vp_p.t1000 out_p.t1594 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2397 out_n.t755 vn_p.t1006 vdd2.t493 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2398 vdd2.t492 vn_p.t1007 out_n.t754 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2399 vdd1.t498 vp_p.t1001 out_p.t1593 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2400 vdd1.t497 vp_p.t1002 out_p.t1592 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2401 out_p.t1591 vp_p.t1003 vdd1.t496 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2402 out_p.t1590 vp_p.t1004 vdd1.t495 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2403 vdd2.t491 vn_p.t1008 out_n.t753 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2404 out_p.t1589 vp_p.t1005 vdd1.t494 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2405 out_n.t752 vn_p.t1009 vdd2.t490 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2406 vdd2.t489 vn_p.t1010 out_n.t751 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2407 vss.t148 vn_n.t200 out_n.t148 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2408 vdd2.t488 vn_p.t1011 out_n.t750 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2409 vdd1.t493 vp_p.t1006 out_p.t1588 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2410 vss.t149 vn_n.t201 out_n.t149 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2411 out_n.t749 vn_p.t1012 vdd2.t487 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2412 vdd1.t492 vp_p.t1007 out_p.t1587 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2413 vdd1.t491 vp_p.t1008 out_p.t1586 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2414 out_n.t748 vn_p.t1013 vdd2.t486 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2415 vdd1.t490 vp_p.t1009 out_p.t1585 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2416 out_p.t1584 vp_p.t1010 vdd1.t489 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2417 vdd1.t488 vp_p.t1011 out_p.t1583 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2418 vdd2.t485 vn_p.t1014 out_n.t747 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2419 vdd1.t487 vp_p.t1012 out_p.t1582 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2420 out_p.t1581 vp_p.t1013 vdd1.t486 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2421 out_n.t746 vn_p.t1015 vdd2.t484 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2422 vdd2.t483 vn_p.t1016 out_n.t745 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2423 out_n.t744 vn_p.t1017 vdd2.t482 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2424 out_p.t1580 vp_p.t1014 vdd1.t485 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2425 out_n.t743 vn_p.t1018 vdd2.t481 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2426 out_n.t742 vn_p.t1019 vdd2.t480 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2427 vdd1.t484 vp_p.t1015 out_p.t1579 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2428 out_n.t741 vn_p.t1020 vdd2.t479 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2429 out_p.t1578 vp_p.t1016 vdd1.t483 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2430 vss.t371 vp_n.t190 out_p.t79 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2431 vdd1.t482 vp_p.t1017 out_p.t1577 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2432 out_n.t740 vn_p.t1021 vdd2.t478 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2433 out_p.t80 vp_n.t191 vss.t370 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2434 out_p.t1576 vp_p.t1018 vdd1.t481 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2435 vss.t110 vn_n.t202 out_n.t110 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2436 out_n.t111 vn_n.t203 vss.t111 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2437 vss.t369 vp_n.t192 out_p.t81 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2438 vdd1.t480 vp_p.t1019 out_p.t1575 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2439 vdd1.t479 vp_p.t1020 out_p.t1574 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2440 out_p.t1573 vp_p.t1021 vdd1.t478 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2441 vdd2.t477 vn_p.t1022 out_n.t739 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2442 vss.t368 vp_n.t193 out_p.t82 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2443 vdd1.t477 vp_p.t1022 out_p.t1572 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2444 out_n.t738 vn_p.t1023 vdd2.t476 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2445 out_n.t112 vn_n.t204 vss.t112 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2446 out_n.t737 vn_p.t1024 vdd2.t475 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2447 vdd2.t474 vn_p.t1025 out_n.t736 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2448 out_n.t113 vn_n.t205 vss.t113 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2449 vdd2.t473 vn_p.t1026 out_n.t735 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2450 vdd2.t472 vn_p.t1027 out_n.t734 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2451 vss.t367 vp_n.t194 out_p.t83 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2452 vdd1.t476 vp_p.t1023 out_p.t1571 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2453 vdd1.t475 vp_p.t1024 out_p.t1570 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2454 vdd2.t471 vn_p.t1028 out_n.t733 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2455 out_p.t1569 vp_p.t1025 vdd1.t474 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2456 vss.t114 vn_n.t206 out_n.t114 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2457 vdd2.t470 vn_p.t1029 out_n.t732 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2458 out_p.t237 vp_n.t195 vss.t366 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2459 out_n.t115 vn_n.t207 vss.t115 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2460 vss.t365 vp_n.t196 out_p.t238 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2461 out_p.t239 vp_n.t197 vss.t364 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2462 vdd1.t473 vp_p.t1026 out_p.t1568 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2463 out_n.t731 vn_p.t1030 vdd2.t469 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2464 out_n.t730 vn_p.t1031 vdd2.t468 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2465 vdd2.t467 vn_p.t1032 out_n.t729 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2466 out_p.t1567 vp_p.t1027 vdd1.t472 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2467 out_n.t728 vn_p.t1033 vdd2.t466 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2468 vdd1.t471 vp_p.t1028 out_p.t1566 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2469 out_p.t1565 vp_p.t1029 vdd1.t470 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2470 vdd1.t469 vp_p.t1030 out_p.t1564 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2471 out_n.t727 vn_p.t1034 vdd2.t465 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2472 vss.t582 vn_n.t208 out_n.t1782 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2473 out_p.t1563 vp_p.t1031 vdd1.t468 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2474 out_p.t1562 vp_p.t1032 vdd1.t467 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2475 out_n.t726 vn_p.t1035 vdd2.t464 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2476 vdd1.t466 vp_p.t1033 out_p.t1561 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2477 vss.t363 vp_n.t198 out_p.t240 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2478 out_p.t1560 vp_p.t1034 vdd1.t465 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2479 out_p.t1559 vp_p.t1035 vdd1.t464 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2480 vss.t583 vn_n.t209 out_n.t1783 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2481 out_n.t725 vn_p.t1036 vdd2.t463 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2482 vdd1.t463 vp_p.t1036 out_p.t1558 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2483 out_n.t724 vn_p.t1037 vdd2.t462 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2484 vdd1.t462 vp_p.t1037 out_p.t1557 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2485 out_p.t1556 vp_p.t1038 vdd1.t461 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2486 vdd1.t460 vp_p.t1039 out_p.t1555 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2487 out_p.t1554 vp_p.t1040 vdd1.t459 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2488 vdd2.t461 vn_p.t1038 out_n.t723 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2489 out_p.t1553 vp_p.t1041 vdd1.t458 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2490 vdd2.t460 vn_p.t1039 out_n.t722 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2491 out_n.t721 vn_p.t1040 vdd2.t459 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2492 vdd2.t458 vn_p.t1041 out_n.t720 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2493 out_n.t719 vn_p.t1042 vdd2.t457 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2494 vss.t362 vp_n.t199 out_p.t241 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2495 out_p.t1552 vp_p.t1042 vdd1.t457 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2496 vdd2.t456 vn_p.t1043 out_n.t718 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2497 out_p.t1551 vp_p.t1043 vdd1.t456 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2498 vdd1.t455 vp_p.t1044 out_p.t1550 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2499 vdd1.t454 vp_p.t1045 out_p.t1549 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2500 out_p.t1548 vp_p.t1046 vdd1.t453 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2501 out_p.t1547 vp_p.t1047 vdd1.t452 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2502 vdd2.t455 vn_p.t1044 out_n.t717 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2503 vdd1.t451 vp_p.t1048 out_p.t1546 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2504 vdd1.t450 vp_p.t1049 out_p.t1545 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2505 out_p.t1544 vp_p.t1050 vdd1.t449 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2506 out_p.t1543 vp_p.t1051 vdd1.t448 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2507 vdd1.t447 vp_p.t1052 out_p.t1542 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2508 out_p.t1541 vp_p.t1053 vdd1.t446 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2509 out_p.t1540 vp_p.t1054 vdd1.t445 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2510 out_n.t716 vn_p.t1045 vdd2.t454 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2511 out_n.t1784 vn_n.t210 vss.t584 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2512 vss.t585 vn_n.t211 out_n.t1785 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2513 vdd2.t453 vn_p.t1046 out_n.t715 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2514 out_p.t242 vp_n.t200 vss.t361 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2515 out_p.t1539 vp_p.t1055 vdd1.t444 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2516 vdd2.t452 vn_p.t1047 out_n.t714 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2517 vdd1.t443 vp_p.t1056 out_p.t1538 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2518 out_n.t713 vn_p.t1048 vdd2.t451 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2519 vdd2.t450 vn_p.t1049 out_n.t712 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2520 out_n.t711 vn_p.t1050 vdd2.t449 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2521 vdd2.t448 vn_p.t1051 out_n.t710 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2522 vss.t586 vn_n.t212 out_n.t1786 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2523 out_n.t709 vn_p.t1052 vdd2.t447 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2524 vdd2.t446 vn_p.t1053 out_n.t708 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2525 out_p.t1537 vp_p.t1057 vdd1.t442 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2526 out_p.t1536 vp_p.t1058 vdd1.t441 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2527 out_p.t1535 vp_p.t1059 vdd1.t440 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2528 vdd1.t439 vp_p.t1060 out_p.t1534 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2529 vss.t360 vp_n.t201 out_p.t243 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2530 vdd2.t445 vn_p.t1054 out_n.t707 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2531 out_p.t244 vp_n.t202 vss.t359 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2532 out_n.t706 vn_p.t1055 vdd2.t444 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2533 vss.t358 vp_n.t203 out_p.t245 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2534 vdd2.t443 vn_p.t1056 out_n.t705 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2535 vdd2.t442 vn_p.t1057 out_n.t704 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2536 out_n.t703 vn_p.t1058 vdd2.t441 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2537 out_p.t1533 vp_p.t1061 vdd1.t438 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2538 out_n.t1787 vn_n.t213 vss.t587 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2539 vss.t94 vn_n.t214 out_n.t94 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2540 vdd2.t440 vn_p.t1059 out_n.t702 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2541 out_p.t1532 vp_p.t1062 vdd1.t437 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2542 vdd2.t439 vn_p.t1060 out_n.t701 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2543 out_n.t700 vn_p.t1061 vdd2.t438 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2544 out_p.t1531 vp_p.t1063 vdd1.t436 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2545 vdd1.t435 vp_p.t1064 out_p.t1530 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2546 vdd1.t434 vp_p.t1065 out_p.t1529 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2547 out_p.t1528 vp_p.t1066 vdd1.t433 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2548 vdd1.t432 vp_p.t1067 out_p.t1527 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2549 out_n.t95 vn_n.t215 vss.t95 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2550 out_p.t1526 vp_p.t1068 vdd1.t431 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2551 out_p.t1525 vp_p.t1069 vdd1.t430 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2552 vdd1.t429 vp_p.t1070 out_p.t1524 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2553 out_p.t1523 vp_p.t1071 vdd1.t428 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2554 vss.t357 vp_n.t204 out_p.t246 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2555 vdd1.t427 vp_p.t1072 out_p.t1522 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2556 vdd1.t426 vp_p.t1073 out_p.t1521 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2557 out_n.t96 vn_n.t216 vss.t96 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2558 vdd2.t437 vn_p.t1062 out_n.t699 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2559 out_p.t1520 vp_p.t1074 vdd1.t425 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2560 out_p.t1519 vp_p.t1075 vdd1.t424 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2561 out_n.t698 vn_p.t1063 vdd2.t436 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2562 vdd2.t435 vn_p.t1064 out_n.t697 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2563 vdd1.t423 vp_p.t1076 out_p.t1518 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2564 out_p.t247 vp_n.t205 vss.t356 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2565 out_p.t1517 vp_p.t1077 vdd1.t422 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2566 vdd1.t421 vp_p.t1078 out_p.t1516 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2567 vdd2.t434 vn_p.t1065 out_n.t696 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2568 vss.t97 vn_n.t217 out_n.t97 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2569 vss.t98 vn_n.t218 out_n.t98 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2570 out_n.t695 vn_p.t1066 vdd2.t433 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2571 out_n.t99 vn_n.t219 vss.t99 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2572 out_p.t1515 vp_p.t1079 vdd1.t420 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2573 out_p.t1514 vp_p.t1080 vdd1.t419 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2574 out_n.t694 vn_p.t1067 vdd2.t432 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2575 vdd1.t418 vp_p.t1081 out_p.t1513 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2576 out_n.t693 vn_p.t1068 vdd2.t431 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2577 vdd2.t430 vn_p.t1069 out_n.t692 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2578 out_p.t1512 vp_p.t1082 vdd1.t417 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2579 out_n.t691 vn_p.t1070 vdd2.t429 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2580 out_n.t690 vn_p.t1071 vdd2.t428 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2581 out_n.t689 vn_p.t1072 vdd2.t427 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2582 vdd2.t426 vn_p.t1073 out_n.t688 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2583 vdd1.t416 vp_p.t1083 out_p.t1511 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2584 vss.t179 vn_n.t220 out_n.t179 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2585 out_p.t1510 vp_p.t1084 vdd1.t415 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2586 out_n.t687 vn_p.t1074 vdd2.t425 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2587 vss.t355 vp_n.t206 out_p.t248 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2588 vdd2.t424 vn_p.t1075 out_n.t686 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2589 vdd1.t414 vp_p.t1085 out_p.t1509 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2590 out_n.t685 vn_p.t1076 vdd2.t423 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2591 vdd2.t422 vn_p.t1077 out_n.t684 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2592 vdd1.t413 vp_p.t1086 out_p.t1508 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2593 out_n.t180 vn_n.t221 vss.t180 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2594 vdd2.t421 vn_p.t1078 out_n.t683 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2595 vdd2.t420 vn_p.t1079 out_n.t682 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2596 out_p.t1507 vp_p.t1087 vdd1.t412 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2597 out_p.t1506 vp_p.t1088 vdd1.t411 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2598 out_n.t681 vn_p.t1080 vdd2.t419 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2599 out_p.t249 vp_n.t207 vss.t354 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2600 vdd1.t410 vp_p.t1089 out_p.t1505 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2601 vdd2.t418 vn_p.t1081 out_n.t680 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2602 vss.t353 vp_n.t208 out_p.t250 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2603 out_n.t679 vn_p.t1082 vdd2.t417 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2604 out_p.t251 vp_n.t209 vss.t352 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2605 vdd2.t416 vn_p.t1083 out_n.t678 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2606 out_n.t677 vn_p.t1084 vdd2.t415 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2607 vdd2.t414 vn_p.t1085 out_n.t676 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2608 vss.t181 vn_n.t222 out_n.t181 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2609 out_n.t182 vn_n.t223 vss.t182 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2610 vdd1.t409 vp_p.t1090 out_p.t1504 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2611 vdd1.t408 vp_p.t1091 out_p.t1503 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2612 out_p.t1502 vp_p.t1092 vdd1.t407 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2613 out_n.t675 vn_p.t1086 vdd2.t413 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2614 out_p.t252 vp_n.t210 vss.t351 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2615 vdd2.t412 vn_p.t1087 out_n.t674 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2616 out_p.t1501 vp_p.t1093 vdd1.t406 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2617 out_p.t1500 vp_p.t1094 vdd1.t405 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2618 out_p.t1499 vp_p.t1095 vdd1.t404 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2619 vdd1.t403 vp_p.t1096 out_p.t1498 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2620 vdd1.t402 vp_p.t1097 out_p.t1497 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2621 out_p.t1496 vp_p.t1098 vdd1.t401 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2622 vdd1.t400 vp_p.t1099 out_p.t1495 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2623 vdd1.t399 vp_p.t1100 out_p.t1494 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2624 out_p.t1493 vp_p.t1101 vdd1.t398 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2625 vss.t350 vp_n.t211 out_p.t253 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2626 out_p.t254 vp_n.t212 vss.t349 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2627 vdd1.t397 vp_p.t1102 out_p.t1492 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2628 out_n.t673 vn_p.t1088 vdd2.t411 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2629 out_n.t672 vn_p.t1089 vdd2.t410 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2630 out_p.t1491 vp_p.t1103 vdd1.t396 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2631 out_p.t1490 vp_p.t1104 vdd1.t395 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2632 vdd1.t394 vp_p.t1105 out_p.t1489 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2633 out_n.t671 vn_p.t1090 vdd2.t409 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2634 vss.t348 vp_n.t213 out_p.t255 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2635 out_p.t1488 vp_p.t1106 vdd1.t393 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2636 out_p.t1487 vp_p.t1107 vdd1.t392 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2637 out_n.t670 vn_p.t1091 vdd2.t408 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2638 vdd2.t407 vn_p.t1092 out_n.t669 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2639 out_n.t183 vn_n.t224 vss.t183 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2640 out_n.t668 vn_p.t1093 vdd2.t406 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2641 out_n.t667 vn_p.t1094 vdd2.t405 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2642 vdd1.t391 vp_p.t1108 out_p.t1486 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2643 vdd2.t404 vn_p.t1095 out_n.t666 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2644 out_n.t665 vn_p.t1096 vdd2.t403 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2645 out_n.t664 vn_p.t1097 vdd2.t402 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2646 vdd2.t401 vn_p.t1098 out_n.t663 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2647 vdd2.t400 vn_p.t1099 out_n.t662 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2648 out_n.t661 vn_p.t1100 vdd2.t399 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2649 vdd2.t398 vn_p.t1101 out_n.t660 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2650 out_n.t659 vn_p.t1102 vdd2.t397 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2651 out_p.t256 vp_n.t214 vss.t347 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2652 vdd2.t396 vn_p.t1103 out_n.t658 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2653 out_p.t1485 vp_p.t1109 vdd1.t390 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2654 out_n.t657 vn_p.t1104 vdd2.t395 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2655 out_n.t184 vn_n.t225 vss.t184 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2656 vdd2.t394 vn_p.t1105 out_n.t656 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2657 out_n.t655 vn_p.t1106 vdd2.t393 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2658 out_n.t60 vn_n.t226 vss.t60 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2659 out_p.t19 vp_n.t215 vss.t346 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2660 vdd2.t392 vn_p.t1107 out_n.t654 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2661 vdd1.t389 vp_p.t1110 out_p.t1484 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2662 vdd2.t391 vn_p.t1108 out_n.t653 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2663 out_p.t1483 vp_p.t1111 vdd1.t388 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2664 out_p.t1482 vp_p.t1112 vdd1.t387 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2665 out_n.t652 vn_p.t1109 vdd2.t390 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2666 vdd2.t389 vn_p.t1110 out_n.t651 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2667 vdd2.t388 vn_p.t1111 out_n.t650 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2668 vss.t61 vn_n.t227 out_n.t61 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2669 out_n.t649 vn_p.t1112 vdd2.t387 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2670 vdd1.t386 vp_p.t1113 out_p.t1481 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2671 vss.t62 vn_n.t228 out_n.t62 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2672 vdd1.t385 vp_p.t1114 out_p.t1480 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2673 out_p.t1479 vp_p.t1115 vdd1.t384 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2674 vdd1.t383 vp_p.t1116 out_p.t1478 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2675 out_n.t648 vn_p.t1113 vdd2.t386 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2676 vdd2.t385 vn_p.t1114 out_n.t647 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2677 out_p.t1477 vp_p.t1117 vdd1.t382 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2678 out_n.t646 vn_p.t1115 vdd2.t384 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2679 out_p.t1476 vp_p.t1118 vdd1.t381 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2680 vdd1.t380 vp_p.t1119 out_p.t1475 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2681 vdd2.t383 vn_p.t1116 out_n.t645 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2682 out_n.t644 vn_p.t1117 vdd2.t382 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2683 vdd1.t379 vp_p.t1120 out_p.t1474 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2684 out_p.t1473 vp_p.t1121 vdd1.t378 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2685 out_n.t643 vn_p.t1118 vdd2.t381 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2686 vdd1.t377 vp_p.t1122 out_p.t1472 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2687 vdd2.t380 vn_p.t1119 out_n.t642 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2688 out_n.t641 vn_p.t1120 vdd2.t379 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2689 vdd1.t376 vp_p.t1123 out_p.t1471 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2690 out_p.t1470 vp_p.t1124 vdd1.t375 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2691 vdd1.t374 vp_p.t1125 out_p.t1469 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2692 out_p.t1468 vp_p.t1126 vdd1.t373 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2693 out_p.t20 vp_n.t216 vss.t345 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2694 out_p.t1467 vp_p.t1127 vdd1.t372 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2695 out_p.t1466 vp_p.t1128 vdd1.t371 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2696 out_p.t1465 vp_p.t1129 vdd1.t370 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2697 vdd1.t369 vp_p.t1130 out_p.t1464 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2698 vdd2.t378 vn_p.t1121 out_n.t640 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2699 out_n.t63 vn_n.t229 vss.t63 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2700 out_n.t639 vn_p.t1122 vdd2.t377 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2701 vss.t344 vp_n.t217 out_p.t21 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2702 out_n.t638 vn_p.t1123 vdd2.t376 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2703 out_p.t1463 vp_p.t1131 vdd1.t368 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2704 vdd1.t367 vp_p.t1132 out_p.t1462 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2705 vdd2.t375 vn_p.t1124 out_n.t637 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2706 out_n.t64 vn_n.t230 vss.t64 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2707 vdd2.t374 vn_p.t1125 out_n.t636 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2708 out_p.t22 vp_n.t218 vss.t343 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2709 vdd1.t366 vp_p.t1133 out_p.t1461 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2710 vdd1.t365 vp_p.t1134 out_p.t1460 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2711 vdd2.t373 vn_p.t1126 out_n.t635 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2712 out_n.t634 vn_p.t1127 vdd2.t372 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2713 vdd2.t371 vn_p.t1128 out_n.t633 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2714 vdd1.t364 vp_p.t1135 out_p.t1459 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2715 vdd2.t370 vn_p.t1129 out_n.t632 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2716 vdd2.t369 vn_p.t1130 out_n.t631 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2717 vdd2.t368 vn_p.t1131 out_n.t630 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2718 vdd2.t367 vn_p.t1132 out_n.t629 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2719 vdd1.t363 vp_p.t1136 out_p.t1458 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2720 out_n.t628 vn_p.t1133 vdd2.t366 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2721 vdd2.t365 vn_p.t1134 out_n.t627 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2722 out_n.t626 vn_p.t1135 vdd2.t364 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2723 vdd2.t363 vn_p.t1136 out_n.t625 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2724 vss.t342 vp_n.t219 out_p.t23 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2725 out_p.t24 vp_n.t220 vss.t341 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2726 out_n.t624 vn_p.t1137 vdd2.t362 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2727 out_n.t623 vn_p.t1138 vdd2.t361 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2728 out_n.t622 vn_p.t1139 vdd2.t360 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2729 vdd2.t359 vn_p.t1140 out_n.t621 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2730 vss.t65 vn_n.t231 out_n.t65 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2731 out_n.t620 vn_p.t1141 vdd2.t358 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2732 out_n.t619 vn_p.t1142 vdd2.t357 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2733 vss.t340 vp_n.t221 out_p.t25 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2734 out_n.t618 vn_p.t1143 vdd2.t356 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2735 out_p.t1457 vp_p.t1137 vdd1.t362 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2736 out_n.t30 vn_n.t232 vss.t30 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2737 out_n.t617 vn_p.t1144 vdd2.t355 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2738 vdd1.t361 vp_p.t1138 out_p.t1456 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2739 out_p.t1455 vp_p.t1139 vdd1.t360 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2740 out_p.t1454 vp_p.t1140 vdd1.t359 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2741 vss.t31 vn_n.t233 out_n.t31 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2742 vdd1.t358 vp_p.t1141 out_p.t1453 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2743 vdd1.t357 vp_p.t1142 out_p.t1452 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2744 vdd2.t354 vn_p.t1145 out_n.t616 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2745 vdd1.t356 vp_p.t1143 out_p.t1451 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2746 out_p.t1450 vp_p.t1144 vdd1.t355 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2747 vdd2.t353 vn_p.t1146 out_n.t615 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2748 out_p.t1449 vp_p.t1145 vdd1.t354 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2749 vdd2.t352 vn_p.t1147 out_n.t614 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2750 vdd1.t353 vp_p.t1146 out_p.t1448 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2751 out_n.t613 vn_p.t1148 vdd2.t351 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2752 vdd2.t350 vn_p.t1149 out_n.t612 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2753 vdd1.t352 vp_p.t1147 out_p.t1447 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2754 out_n.t32 vn_n.t234 vss.t32 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2755 out_p.t1446 vp_p.t1148 vdd1.t351 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2756 vdd1.t350 vp_p.t1149 out_p.t1445 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2757 out_p.t1444 vp_p.t1150 vdd1.t349 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2758 out_p.t1443 vp_p.t1151 vdd1.t348 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2759 out_n.t33 vn_n.t235 vss.t33 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2760 vdd2.t349 vn_p.t1150 out_n.t611 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2761 vss.t339 vp_n.t222 out_p.t26 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2762 out_p.t1442 vp_p.t1152 vdd1.t347 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2763 vdd2.t348 vn_p.t1151 out_n.t610 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2764 vdd1.t346 vp_p.t1153 out_p.t1441 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2765 vdd1.t345 vp_p.t1154 out_p.t1440 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2766 out_p.t1439 vp_p.t1155 vdd1.t344 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2767 out_n.t609 vn_p.t1152 vdd2.t347 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2768 vdd1.t343 vp_p.t1156 out_p.t1438 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2769 out_n.t608 vn_p.t1153 vdd2.t346 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2770 vdd2.t345 vn_p.t1154 out_n.t607 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2771 vdd1.t342 vp_p.t1157 out_p.t1437 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2772 vdd1.t341 vp_p.t1158 out_p.t1436 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2773 out_p.t1435 vp_p.t1159 vdd1.t340 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2774 out_n.t606 vn_p.t1155 vdd2.t344 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2775 vdd2.t343 vn_p.t1156 out_n.t605 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2776 out_p.t27 vp_n.t223 vss.t338 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2777 out_p.t1434 vp_p.t1160 vdd1.t339 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2778 vdd2.t342 vn_p.t1157 out_n.t604 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2779 vss.t337 vp_n.t224 out_p.t28 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2780 vdd1.t338 vp_p.t1161 out_p.t1433 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2781 out_p.t29 vp_n.t225 vss.t336 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2782 out_n.t603 vn_p.t1158 vdd2.t341 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2783 out_p.t1432 vp_p.t1162 vdd1.t337 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2784 out_p.t1431 vp_p.t1163 vdd1.t336 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2785 out_n.t602 vn_p.t1159 vdd2.t340 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2786 out_n.t601 vn_p.t1160 vdd2.t339 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2787 out_p.t1430 vp_p.t1164 vdd1.t335 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2788 vdd2.t338 vn_p.t1161 out_n.t600 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2789 vss.t34 vn_n.t236 out_n.t34 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2790 out_n.t599 vn_p.t1162 vdd2.t337 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2791 out_n.t598 vn_p.t1163 vdd2.t336 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2792 out_p.t1429 vp_p.t1165 vdd1.t334 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2793 out_n.t597 vn_p.t1164 vdd2.t335 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2794 out_p.t30 vp_n.t226 vss.t335 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2795 vdd2.t334 vn_p.t1165 out_n.t596 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2796 vss.t334 vp_n.t227 out_p.t31 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2797 vss.t333 vp_n.t228 out_p.t32 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2798 vdd2.t333 vn_p.t1166 out_n.t595 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2799 vdd2.t332 vn_p.t1167 out_n.t594 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2800 out_n.t593 vn_p.t1168 vdd2.t331 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2801 out_n.t35 vn_n.t237 vss.t35 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2802 vdd2.t330 vn_p.t1169 out_n.t592 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2803 out_p.t1428 vp_p.t1166 vdd1.t333 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2804 out_n.t1776 vn_n.t238 vss.t576 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2805 out_p.t1427 vp_p.t1167 vdd1.t332 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2806 vdd1.t331 vp_p.t1168 out_p.t1426 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2807 out_p.t1425 vp_p.t1169 vdd1.t330 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2808 vdd2.t329 vn_p.t1170 out_n.t591 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2809 vdd1.t329 vp_p.t1170 out_p.t1424 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2810 vdd1.t328 vp_p.t1171 out_p.t1423 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2811 out_p.t1422 vp_p.t1172 vdd1.t327 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2812 vdd1.t326 vp_p.t1173 out_p.t1421 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2813 out_p.t1420 vp_p.t1174 vdd1.t325 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2814 vdd1.t324 vp_p.t1175 out_p.t1419 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2815 out_p.t33 vp_n.t229 vss.t332 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2816 vdd1.t323 vp_p.t1176 out_p.t1418 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2817 out_p.t1417 vp_p.t1177 vdd1.t322 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2818 out_n.t590 vn_p.t1171 vdd2.t328 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2819 out_n.t589 vn_p.t1172 vdd2.t327 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2820 vdd2.t326 vn_p.t1173 out_n.t588 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2821 out_p.t1416 vp_p.t1178 vdd1.t321 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2822 vdd1.t320 vp_p.t1179 out_p.t1415 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2823 vdd1.t319 vp_p.t1180 out_p.t1414 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2824 vdd2.t325 vn_p.t1174 out_n.t587 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2825 out_p.t1413 vp_p.t1181 vdd1.t318 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2826 out_n.t586 vn_p.t1175 vdd2.t324 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2827 vss.t577 vn_n.t239 out_n.t1777 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2828 out_p.t1412 vp_p.t1182 vdd1.t317 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2829 vdd1.t316 vp_p.t1183 out_p.t1411 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2830 out_p.t1410 vp_p.t1184 vdd1.t315 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2831 vdd1.t314 vp_p.t1185 out_p.t1409 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2832 vss.t578 vn_n.t240 out_n.t1778 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2833 vdd1.t313 vp_p.t1186 out_p.t1408 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2834 out_p.t1407 vp_p.t1187 vdd1.t312 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2835 out_n.t585 vn_p.t1176 vdd2.t323 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2836 vdd1.t311 vp_p.t1188 out_p.t1406 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2837 vdd2.t322 vn_p.t1177 out_n.t584 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2838 out_n.t583 vn_p.t1178 vdd2.t321 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2839 out_p.t1405 vp_p.t1189 vdd1.t310 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2840 vdd2.t320 vn_p.t1179 out_n.t582 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2841 out_n.t581 vn_p.t1180 vdd2.t319 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2842 out_p.t1404 vp_p.t1190 vdd1.t309 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2843 vdd1.t308 vp_p.t1191 out_p.t1403 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2844 out_n.t580 vn_p.t1181 vdd2.t318 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2845 out_n.t579 vn_p.t1182 vdd2.t317 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2846 vss.t331 vp_n.t230 out_p.t34 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2847 out_p.t35 vp_n.t231 vss.t330 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2848 out_p.t1402 vp_p.t1192 vdd1.t307 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2849 vdd1.t306 vp_p.t1193 out_p.t1401 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2850 vss.t329 vp_n.t232 out_p.t36 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2851 out_n.t1779 vn_n.t241 vss.t579 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2852 vdd2.t316 vn_p.t1183 out_n.t578 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2853 vdd1.t305 vp_p.t1194 out_p.t1400 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2854 vss.t580 vn_n.t242 out_n.t1780 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2855 out_p.t1399 vp_p.t1195 vdd1.t304 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2856 vdd2.t315 vn_p.t1184 out_n.t577 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2857 vdd1.t303 vp_p.t1196 out_p.t1398 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2858 vdd2.t314 vn_p.t1185 out_n.t576 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2859 vdd2.t313 vn_p.t1186 out_n.t575 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2860 out_n.t574 vn_p.t1187 vdd2.t312 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2861 vdd2.t311 vn_p.t1188 out_n.t573 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2862 out_n.t572 vn_p.t1189 vdd2.t310 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2863 out_p.t37 vp_n.t233 vss.t328 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2864 out_n.t1781 vn_n.t243 vss.t581 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2865 vdd2.t309 vn_p.t1190 out_n.t571 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2866 vdd2.t308 vn_p.t1191 out_n.t570 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2867 vdd1.t302 vp_p.t1197 out_p.t1397 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2868 vss.t327 vp_n.t234 out_p.t38 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2869 out_p.t105 vp_n.t235 vss.t326 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2870 out_p.t106 vp_n.t236 vss.t325 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2871 vdd2.t307 vn_p.t1192 out_n.t569 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2872 out_p.t1396 vp_p.t1198 vdd1.t301 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2873 vss.t252 vn_n.t244 out_n.t252 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2874 vdd1.t300 vp_p.t1199 out_p.t1395 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2875 vdd2.t306 vn_p.t1193 out_n.t568 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2876 out_n.t567 vn_p.t1194 vdd2.t305 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2877 out_n.t566 vn_p.t1195 vdd2.t304 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2878 out_n.t565 vn_p.t1196 vdd2.t303 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2879 vdd1.t299 vp_p.t1200 out_p.t1394 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2880 vdd1.t298 vp_p.t1201 out_p.t1393 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2881 out_p.t1392 vp_p.t1202 vdd1.t297 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2882 vdd1.t296 vp_p.t1203 out_p.t1391 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2883 out_p.t1390 vp_p.t1204 vdd1.t295 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2884 out_p.t1389 vp_p.t1205 vdd1.t294 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2885 out_p.t1388 vp_p.t1206 vdd1.t293 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2886 vdd2.t302 vn_p.t1197 out_n.t564 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2887 out_p.t1387 vp_p.t1207 vdd1.t292 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2888 out_p.t1386 vp_p.t1208 vdd1.t291 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2889 vdd1.t290 vp_p.t1209 out_p.t1385 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2890 vdd1.t289 vp_p.t1210 out_p.t1384 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2891 vss.t253 vn_n.t245 out_n.t253 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2892 vdd2.t301 vn_p.t1198 out_n.t563 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2893 out_n.t562 vn_p.t1199 vdd2.t300 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2894 out_n.t561 vn_p.t1200 vdd2.t299 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2895 vdd1.t288 vp_p.t1211 out_p.t1383 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2896 vdd2.t298 vn_p.t1201 out_n.t560 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2897 out_n.t559 vn_p.t1202 vdd2.t297 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2898 vdd2.t296 vn_p.t1203 out_n.t558 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2899 out_n.t557 vn_p.t1204 vdd2.t295 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2900 out_p.t1382 vp_p.t1212 vdd1.t287 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2901 vdd2.t294 vn_p.t1205 out_n.t556 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2902 out_n.t555 vn_p.t1206 vdd2.t293 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2903 out_p.t1381 vp_p.t1213 vdd1.t286 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2904 out_p.t1380 vp_p.t1214 vdd1.t285 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2905 out_p.t1379 vp_p.t1215 vdd1.t284 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2906 vdd1.t283 vp_p.t1216 out_p.t1378 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2907 vdd2.t292 vn_p.t1207 out_n.t554 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2908 out_n.t553 vn_p.t1208 vdd2.t291 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2909 vdd1.t282 vp_p.t1217 out_p.t1377 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2910 out_n.t254 vn_n.t246 vss.t254 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2911 out_p.t1376 vp_p.t1218 vdd1.t281 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2912 vdd2.t290 vn_p.t1209 out_n.t552 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2913 out_p.t107 vp_n.t237 vss.t324 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2914 vdd1.t280 vp_p.t1219 out_p.t1375 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2915 vss.t323 vp_n.t238 out_p.t108 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2916 vdd1.t279 vp_p.t1220 out_p.t1374 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2917 out_p.t109 vp_n.t239 vss.t322 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2918 vdd2.t289 vn_p.t1210 out_n.t551 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2919 vdd2.t288 vn_p.t1211 out_n.t550 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2920 out_n.t549 vn_p.t1212 vdd2.t287 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2921 out_n.t548 vn_p.t1213 vdd2.t286 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2922 out_n.t255 vn_n.t247 vss.t255 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2923 vss.t256 vn_n.t248 out_n.t256 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2924 vdd2.t285 vn_p.t1214 out_n.t547 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2925 vdd1.t278 vp_p.t1221 out_p.t1373 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2926 out_p.t1372 vp_p.t1222 vdd1.t277 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2927 out_n.t546 vn_p.t1215 vdd2.t284 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2928 vdd2.t283 vn_p.t1216 out_n.t545 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2929 out_p.t110 vp_n.t240 vss.t321 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2930 out_n.t544 vn_p.t1217 vdd2.t282 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2931 vss.t257 vn_n.t249 out_n.t257 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2932 out_n.t543 vn_p.t1218 vdd2.t281 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2933 vdd2.t280 vn_p.t1219 out_n.t542 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2934 out_p.t111 vp_n.t241 vss.t320 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2935 out_p.t1371 vp_p.t1223 vdd1.t276 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2936 vdd1.t275 vp_p.t1224 out_p.t1370 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2937 vdd2.t279 vn_p.t1220 out_n.t541 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2938 out_n.t540 vn_p.t1221 vdd2.t278 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2939 out_n.t539 vn_p.t1222 vdd2.t277 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2940 vss.t319 vp_n.t242 out_p.t112 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2941 vdd2.t276 vn_p.t1223 out_n.t538 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2942 out_p.t113 vp_n.t243 vss.t318 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2943 out_n.t537 vn_p.t1224 vdd2.t275 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2944 vss.t317 vp_n.t244 out_p.t114 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2945 out_n.t536 vn_p.t1225 vdd2.t274 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2946 out_n.t535 vn_p.t1226 vdd2.t273 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2947 out_p.t1369 vp_p.t1225 vdd1.t274 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2948 out_n.t534 vn_p.t1227 vdd2.t272 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2949 vdd1.t273 vp_p.t1226 out_p.t1368 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2950 out_p.t1367 vp_p.t1227 vdd1.t272 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2951 out_n.t53 vn_n.t250 vss.t53 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2952 vdd2.t271 vn_p.t1228 out_n.t533 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2953 out_n.t532 vn_p.t1229 vdd2.t270 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2954 vdd1.t271 vp_p.t1228 out_p.t1366 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2955 vdd1.t270 vp_p.t1229 out_p.t1365 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2956 out_p.t1364 vp_p.t1230 vdd1.t269 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2957 out_p.t1363 vp_p.t1231 vdd1.t268 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2958 vdd1.t267 vp_p.t1232 out_p.t1362 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2959 vdd1.t266 vp_p.t1233 out_p.t1361 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2960 vdd1.t265 vp_p.t1234 out_p.t1360 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2961 vdd2.t269 vn_p.t1230 out_n.t531 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2962 vdd1.t264 vp_p.t1235 out_p.t1359 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2963 out_p.t1358 vp_p.t1236 vdd1.t263 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2964 out_p.t115 vp_n.t245 vss.t316 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2965 vdd1.t262 vp_p.t1237 out_p.t1357 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2966 vdd1.t261 vp_p.t1238 out_p.t1356 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2967 vdd2.t268 vn_p.t1231 out_n.t530 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2968 out_n.t529 vn_p.t1232 vdd2.t267 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2969 out_p.t1355 vp_p.t1239 vdd1.t260 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2970 vdd2.t266 vn_p.t1233 out_n.t528 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2971 vdd1.t259 vp_p.t1240 out_p.t1354 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2972 vdd2.t265 vn_p.t1234 out_n.t527 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2973 out_p.t1353 vp_p.t1241 vdd1.t258 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2974 vdd2.t264 vn_p.t1235 out_n.t526 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2975 out_p.t116 vp_n.t246 vss.t315 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2976 out_n.t525 vn_p.t1236 vdd2.t263 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2977 vdd2.t262 vn_p.t1237 out_n.t524 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2978 vdd2.t261 vn_p.t1238 out_n.t523 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2979 out_p.t1352 vp_p.t1242 vdd1.t257 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2980 vdd1.t256 vp_p.t1243 out_p.t1351 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2981 vdd1.t255 vp_p.t1244 out_p.t1350 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2982 vdd2.t260 vn_p.t1239 out_n.t522 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2983 out_p.t1349 vp_p.t1245 vdd1.t254 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2984 out_n.t521 vn_p.t1240 vdd2.t259 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2985 vss.t54 vn_n.t251 out_n.t54 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2986 vdd2.t258 vn_p.t1241 out_n.t520 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2987 vdd1.t253 vp_p.t1246 out_p.t1348 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2988 vss.t55 vn_n.t252 out_n.t55 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2989 out_p.t1347 vp_p.t1247 vdd1.t252 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2990 out_p.t1346 vp_p.t1248 vdd1.t251 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2991 out_n.t519 vn_p.t1242 vdd2.t257 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2992 out_n.t518 vn_p.t1243 vdd2.t256 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2993 vss.t314 vp_n.t247 out_p.t117 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2994 out_n.t517 vn_p.t1244 vdd2.t255 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2995 vdd2.t254 vn_p.t1245 out_n.t516 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2996 vdd1.t250 vp_p.t1249 out_p.t1345 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2997 out_n.t515 vn_p.t1246 vdd2.t253 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2998 out_n.t514 vn_p.t1247 vdd2.t252 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2999 out_n.t513 vn_p.t1248 vdd2.t251 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3000 out_n.t512 vn_p.t1249 vdd2.t250 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3001 vss.t56 vn_n.t253 out_n.t56 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3002 vdd2.t249 vn_p.t1250 out_n.t511 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3003 out_n.t510 vn_p.t1251 vdd2.t248 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3004 out_p.t1344 vp_p.t1250 vdd1.t249 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3005 vdd2.t247 vn_p.t1252 out_n.t509 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3006 vdd1.t248 vp_p.t1251 out_p.t1343 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3007 vdd1.t247 vp_p.t1252 out_p.t1342 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3008 vdd2.t246 vn_p.t1253 out_n.t508 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3009 out_n.t507 vn_p.t1254 vdd2.t245 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3010 vdd1.t246 vp_p.t1253 out_p.t1341 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3011 vdd1.t245 vp_p.t1254 out_p.t1340 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3012 vdd2.t244 vn_p.t1255 out_n.t506 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3013 out_p.t1339 vp_p.t1255 vdd1.t244 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3014 vdd1.t243 vp_p.t1256 out_p.t1338 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3015 out_p.t1337 vp_p.t1257 vdd1.t242 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3016 vdd2.t243 vn_p.t1256 out_n.t505 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3017 out_n.t504 vn_p.t1257 vdd2.t242 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3018 vdd2.t241 vn_p.t1258 out_n.t503 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3019 out_n.t502 vn_p.t1259 vdd2.t240 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3020 vdd2.t239 vn_p.t1260 out_n.t501 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3021 out_n.t500 vn_p.t1261 vdd2.t238 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3022 out_p.t118 vp_n.t248 vss.t313 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3023 vdd2.t237 vn_p.t1262 out_n.t499 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3024 out_p.t119 vp_n.t249 vss.t312 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3025 vdd2.t236 vn_p.t1263 out_n.t498 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3026 vdd1.t241 vp_p.t1258 out_p.t1336 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3027 out_p.t1335 vp_p.t1259 vdd1.t240 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3028 out_n.t497 vn_p.t1264 vdd2.t235 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3029 vdd1.t239 vp_p.t1260 out_p.t1334 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3030 vss.t57 vn_n.t254 out_n.t57 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3031 out_n.t58 vn_n.t255 vss.t58 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3032 out_p.t1333 vp_p.t1261 vdd1.t238 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3033 vdd1.t237 vp_p.t1262 out_p.t1332 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3034 vdd1.t236 vp_p.t1263 out_p.t1331 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3035 out_p.t1330 vp_p.t1264 vdd1.t235 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3036 out_n.t496 vn_p.t1265 vdd2.t234 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3037 out_n.t495 vn_p.t1266 vdd2.t233 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3038 out_p.t1329 vp_p.t1265 vdd1.t234 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3039 vdd1.t233 vp_p.t1266 out_p.t1328 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3040 out_n.t494 vn_p.t1267 vdd2.t232 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3041 vss.t311 vp_n.t250 out_p.t120 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3042 vdd1.t232 vp_p.t1267 out_p.t1327 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3043 vdd1.t231 vp_p.t1268 out_p.t1326 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3044 out_p.t1325 vp_p.t1269 vdd1.t230 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3045 out_p.t1324 vp_p.t1270 vdd1.t229 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3046 vdd1.t228 vp_p.t1271 out_p.t1323 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3047 out_p.t121 vp_n.t251 vss.t310 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3048 out_p.t1322 vp_p.t1272 vdd1.t227 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3049 vdd1.t226 vp_p.t1273 out_p.t1321 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3050 out_n.t493 vn_p.t1268 vdd2.t231 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3051 vss.t59 vn_n.t256 out_n.t59 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3052 out_n.t492 vn_p.t1269 vdd2.t230 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3053 vss.t309 vp_n.t252 out_p.t122 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3054 vdd1.t225 vp_p.t1274 out_p.t1320 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3055 out_p.t1319 vp_p.t1275 vdd1.t224 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3056 out_n.t491 vn_p.t1270 vdd2.t229 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3057 vdd2.t228 vn_p.t1271 out_n.t490 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3058 vdd2.t227 vn_p.t1272 out_n.t489 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3059 vdd1.t223 vp_p.t1276 out_p.t1318 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3060 vdd2.t226 vn_p.t1273 out_n.t488 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3061 out_n.t487 vn_p.t1274 vdd2.t225 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3062 vdd2.t224 vn_p.t1275 out_n.t486 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3063 out_n.t485 vn_p.t1276 vdd2.t223 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3064 vdd2.t222 vn_p.t1277 out_n.t484 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3065 vdd1.t222 vp_p.t1277 out_p.t1317 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3066 out_p.t123 vp_n.t253 vss.t308 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3067 out_n.t483 vn_p.t1278 vdd2.t221 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3068 vdd2.t220 vn_p.t1279 out_n.t482 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3069 vdd2.t219 vn_p.t1280 out_n.t481 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3070 out_n.t17 vn_n.t257 vss.t17 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3071 out_n.t480 vn_p.t1281 vdd2.t218 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3072 out_n.t479 vn_p.t1282 vdd2.t217 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3073 out_n.t478 vn_p.t1283 vdd2.t216 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3074 vdd2.t215 vn_p.t1284 out_n.t477 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3075 out_n.t476 vn_p.t1285 vdd2.t214 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3076 vdd2.t213 vn_p.t1286 out_n.t475 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3077 vdd1.t221 vp_p.t1278 out_p.t1316 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3078 vdd2.t212 vn_p.t1287 out_n.t474 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3079 out_p.t1315 vp_p.t1279 vdd1.t220 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3080 out_p.t1314 vp_p.t1280 vdd1.t219 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3081 vdd1.t218 vp_p.t1281 out_p.t1313 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3082 out_n.t473 vn_p.t1288 vdd2.t211 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3083 vdd2.t210 vn_p.t1289 out_n.t472 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3084 out_n.t471 vn_p.t1290 vdd2.t209 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3085 out_p.t1312 vp_p.t1282 vdd1.t217 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3086 vdd1.t216 vp_p.t1283 out_p.t1311 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3087 vss.t18 vn_n.t258 out_n.t18 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3088 out_n.t470 vn_p.t1291 vdd2.t208 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3089 vss.t19 vn_n.t259 out_n.t19 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3090 vss.t307 vp_n.t254 out_p.t124 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3091 out_n.t469 vn_p.t1292 vdd2.t207 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3092 vdd2.t206 vn_p.t1293 out_n.t468 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3093 out_n.t467 vn_p.t1294 vdd2.t205 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3094 out_p.t1310 vp_p.t1284 vdd1.t215 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3095 out_p.t1309 vp_p.t1285 vdd1.t214 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3096 out_p.t1308 vp_p.t1286 vdd1.t213 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3097 out_p.t1307 vp_p.t1287 vdd1.t212 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3098 vdd1.t211 vp_p.t1288 out_p.t1306 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3099 out_n.t466 vn_p.t1295 vdd2.t204 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3100 vdd1.t210 vp_p.t1289 out_p.t1305 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3101 vdd1.t209 vp_p.t1290 out_p.t1304 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3102 vss.t20 vn_n.t260 out_n.t20 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3103 out_n.t465 vn_p.t1296 vdd2.t203 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3104 vdd1.t208 vp_p.t1291 out_p.t1303 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3105 vdd1.t207 vp_p.t1292 out_p.t1302 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3106 out_n.t21 vn_n.t261 vss.t21 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3107 vdd2.t202 vn_p.t1297 out_n.t464 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3108 vdd1.t206 vp_p.t1293 out_p.t1301 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3109 vss.t22 vn_n.t262 out_n.t22 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3110 out_n.t463 vn_p.t1298 vdd2.t201 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3111 vdd1.t205 vp_p.t1294 out_p.t1300 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3112 out_p.t1299 vp_p.t1295 vdd1.t204 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3113 vdd1.t203 vp_p.t1296 out_p.t1298 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3114 out_p.t1297 vp_p.t1297 vdd1.t202 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3115 out_n.t462 vn_p.t1299 vdd2.t200 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3116 out_p.t85 vp_n.t255 vss.t306 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3117 vss.t305 vp_n.t256 out_p.t86 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3118 out_p.t1296 vp_p.t1298 vdd1.t201 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3119 vss.t304 vp_n.t257 out_p.t87 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3120 vdd1.t200 vp_p.t1299 out_p.t1295 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3121 vdd2.t199 vn_p.t1300 out_n.t461 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3122 vdd1.t199 vp_p.t1300 out_p.t1294 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3123 out_p.t1293 vp_p.t1301 vdd1.t198 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3124 out_n.t23 vn_n.t263 vss.t23 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3125 vdd2.t198 vn_p.t1301 out_n.t460 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3126 out_n.t459 vn_p.t1302 vdd2.t197 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3127 out_p.t1292 vp_p.t1302 vdd1.t197 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3128 out_p.t1291 vp_p.t1303 vdd1.t196 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3129 vdd1.t195 vp_p.t1304 out_p.t1290 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3130 vdd1.t194 vp_p.t1305 out_p.t1289 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3131 vdd2.t196 vn_p.t1303 out_n.t458 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3132 out_n.t457 vn_p.t1304 vdd2.t195 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3133 vdd2.t194 vn_p.t1305 out_n.t456 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3134 vdd2.t193 vn_p.t1306 out_n.t455 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3135 vdd2.t192 vn_p.t1307 out_n.t454 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3136 out_n.t453 vn_p.t1308 vdd2.t191 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3137 vss.t303 vp_n.t258 out_p.t88 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3138 vss.t6 vn_n.t264 out_n.t6 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3139 out_n.t452 vn_p.t1309 vdd2.t190 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3140 out_n.t451 vn_p.t1310 vdd2.t189 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3141 out_n.t450 vn_p.t1311 vdd2.t188 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3142 vdd1.t193 vp_p.t1306 out_p.t1288 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3143 vdd2.t187 vn_p.t1312 out_n.t449 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3144 out_n.t448 vn_p.t1313 vdd2.t186 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3145 vdd2.t185 vn_p.t1314 out_n.t447 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3146 vss.t302 vp_n.t259 out_p.t89 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3147 out_n.t446 vn_p.t1315 vdd2.t184 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3148 vdd2.t183 vn_p.t1316 out_n.t445 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3149 out_p.t1287 vp_p.t1307 vdd1.t192 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3150 vdd2.t182 vn_p.t1317 out_n.t444 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3151 out_n.t443 vn_p.t1318 vdd2.t181 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3152 out_p.t1286 vp_p.t1308 vdd1.t191 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3153 vss.t7 vn_n.t265 out_n.t7 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3154 vdd1.t190 vp_p.t1309 out_p.t1285 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3155 vdd1.t189 vp_p.t1310 out_p.t1284 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3156 vdd1.t188 vp_p.t1311 out_p.t1283 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3157 out_p.t1282 vp_p.t1312 vdd1.t187 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3158 out_p.t1281 vp_p.t1313 vdd1.t186 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3159 vdd1.t185 vp_p.t1314 out_p.t1280 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3160 vdd2.t180 vn_p.t1319 out_n.t442 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3161 out_p.t1279 vp_p.t1315 vdd1.t184 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3162 out_p.t1278 vp_p.t1316 vdd1.t183 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3163 out_n.t441 vn_p.t1320 vdd2.t179 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3164 out_p.t1277 vp_p.t1317 vdd1.t182 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3165 out_n.t440 vn_p.t1321 vdd2.t178 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3166 vdd1.t181 vp_p.t1318 out_p.t1276 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3167 out_p.t1275 vp_p.t1319 vdd1.t180 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3168 out_p.t1274 vp_p.t1320 vdd1.t179 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3169 vdd2.t177 vn_p.t1322 out_n.t439 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3170 vdd2.t176 vn_p.t1323 out_n.t438 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3171 out_n.t437 vn_p.t1324 vdd2.t175 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3172 vdd2.t174 vn_p.t1325 out_n.t436 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3173 vdd1.t178 vp_p.t1321 out_p.t1273 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3174 out_p.t1272 vp_p.t1322 vdd1.t177 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3175 vdd1.t176 vp_p.t1323 out_p.t1271 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3176 vdd1.t175 vp_p.t1324 out_p.t1270 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3177 out_p.t90 vp_n.t260 vss.t301 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3178 out_p.t1269 vp_p.t1325 vdd1.t174 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3179 out_p.t1268 vp_p.t1326 vdd1.t173 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3180 out_n.t8 vn_n.t266 vss.t8 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3181 vss.t9 vn_n.t267 out_n.t9 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3182 out_n.t435 vn_p.t1326 vdd2.t173 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3183 out_p.t1267 vp_p.t1327 vdd1.t172 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3184 out_p.t1266 vp_p.t1328 vdd1.t171 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3185 out_p.t1265 vp_p.t1329 vdd1.t170 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3186 out_n.t10 vn_n.t268 vss.t10 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3187 vdd1.t169 vp_p.t1330 out_p.t1264 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3188 vdd2.t172 vn_p.t1327 out_n.t434 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3189 vss.t300 vp_n.t261 out_p.t91 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3190 vdd1.t168 vp_p.t1331 out_p.t1263 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3191 out_p.t1262 vp_p.t1332 vdd1.t167 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3192 out_n.t433 vn_p.t1328 vdd2.t171 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3193 vdd2.t170 vn_p.t1329 out_n.t432 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3194 out_p.t92 vp_n.t262 vss.t299 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3195 vdd1.t166 vp_p.t1333 out_p.t1261 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3196 vdd1.t165 vp_p.t1334 out_p.t1260 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3197 out_n.t431 vn_p.t1330 vdd2.t169 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3198 out_p.t93 vp_n.t263 vss.t298 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3199 out_n.t430 vn_p.t1331 vdd2.t168 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3200 vdd2.t167 vn_p.t1332 out_n.t429 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3201 vdd2.t166 vn_p.t1333 out_n.t428 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3202 out_p.t1259 vp_p.t1335 vdd1.t164 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3203 vdd2.t165 vn_p.t1334 out_n.t427 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3204 out_n.t426 vn_p.t1335 vdd2.t164 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3205 vdd2.t163 vn_p.t1336 out_n.t425 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3206 out_n.t424 vn_p.t1337 vdd2.t162 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3207 vss.t11 vn_n.t269 out_n.t11 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3208 out_n.t423 vn_p.t1338 vdd2.t161 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3209 vdd2.t160 vn_p.t1339 out_n.t422 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3210 out_p.t1258 vp_p.t1336 vdd1.t163 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3211 vdd2.t159 vn_p.t1340 out_n.t421 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3212 vss.t12 vn_n.t270 out_n.t12 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3213 out_n.t420 vn_p.t1341 vdd2.t158 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3214 out_p.t94 vp_n.t264 vss.t297 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3215 out_p.t95 vp_n.t265 vss.t296 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3216 vss.t81 vn_n.t271 out_n.t81 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3217 vdd2.t157 vn_p.t1342 out_n.t419 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3218 out_n.t418 vn_p.t1343 vdd2.t156 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3219 vss.t295 vp_n.t266 out_p.t96 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3220 out_n.t82 vn_n.t272 vss.t82 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3221 out_n.t417 vn_p.t1344 vdd2.t155 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3222 out_n.t416 vn_p.t1345 vdd2.t154 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3223 vdd2.t153 vn_p.t1346 out_n.t415 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3224 vdd2.t152 vn_p.t1347 out_n.t414 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3225 out_n.t413 vn_p.t1348 vdd2.t151 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3226 vdd2.t150 vn_p.t1349 out_n.t412 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3227 out_n.t411 vn_p.t1350 vdd2.t149 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3228 out_n.t83 vn_n.t273 vss.t83 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3229 vdd2.t148 vn_p.t1351 out_n.t410 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3230 out_p.t1257 vp_p.t1337 vdd1.t162 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3231 out_p.t1256 vp_p.t1338 vdd1.t161 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3232 out_p.t1255 vp_p.t1339 vdd1.t160 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3233 out_p.t1254 vp_p.t1340 vdd1.t159 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3234 out_n.t409 vn_p.t1352 vdd2.t147 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3235 vdd2.t146 vn_p.t1353 out_n.t408 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3236 vdd1.t158 vp_p.t1341 out_p.t1253 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3237 out_p.t1252 vp_p.t1342 vdd1.t157 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3238 vdd2.t145 vn_p.t1354 out_n.t407 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3239 vdd1.t156 vp_p.t1343 out_p.t1251 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3240 vdd1.t155 vp_p.t1344 out_p.t1250 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3241 vdd2.t144 vn_p.t1355 out_n.t406 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3242 vdd1.t154 vp_p.t1345 out_p.t1249 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3243 vdd2.t143 vn_p.t1356 out_n.t405 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3244 vdd1.t153 vp_p.t1346 out_p.t1248 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3245 vss.t84 vn_n.t274 out_n.t84 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3246 out_n.t404 vn_p.t1357 vdd2.t142 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3247 vdd2.t141 vn_p.t1358 out_n.t403 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3248 out_p.t1247 vp_p.t1347 vdd1.t152 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3249 vdd2.t140 vn_p.t1359 out_n.t402 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3250 out_n.t401 vn_p.t1360 vdd2.t139 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3251 vdd2.t138 vn_p.t1361 out_n.t400 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3252 out_p.t1246 vp_p.t1348 vdd1.t151 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3253 vss.t85 vn_n.t275 out_n.t85 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3254 out_n.t399 vn_p.t1362 vdd2.t137 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3255 vdd1.t150 vp_p.t1349 out_p.t1245 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3256 out_p.t1244 vp_p.t1350 vdd1.t149 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3257 out_p.t1243 vp_p.t1351 vdd1.t148 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3258 out_n.t398 vn_p.t1363 vdd2.t136 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3259 vdd1.t147 vp_p.t1352 out_p.t1242 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3260 vdd1.t146 vp_p.t1353 out_p.t1241 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3261 vdd1.t145 vp_p.t1354 out_p.t1240 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3262 out_n.t397 vn_p.t1364 vdd2.t135 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3263 vdd2.t134 vn_p.t1365 out_n.t396 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3264 out_p.t97 vp_n.t267 vss.t294 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3265 out_p.t1239 vp_p.t1355 vdd1.t144 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3266 out_n.t395 vn_p.t1366 vdd2.t133 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3267 vdd1.t143 vp_p.t1356 out_p.t1238 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3268 out_p.t1237 vp_p.t1357 vdd1.t142 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3269 out_n.t394 vn_p.t1367 vdd2.t132 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3270 out_p.t1236 vp_p.t1358 vdd1.t141 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3271 out_p.t1235 vp_p.t1359 vdd1.t140 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3272 vdd1.t139 vp_p.t1360 out_p.t1234 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3273 out_n.t393 vn_p.t1368 vdd2.t131 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3274 vss.t293 vp_n.t268 out_p.t98 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3275 vdd1.t138 vp_p.t1361 out_p.t1233 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3276 out_n.t392 vn_p.t1369 vdd2.t130 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3277 out_p.t99 vp_n.t269 vss.t292 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3278 out_p.t1232 vp_p.t1362 vdd1.t137 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3279 vss.t291 vp_n.t270 out_p.t100 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3280 out_n.t391 vn_p.t1370 vdd2.t129 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3281 vdd1.t136 vp_p.t1363 out_p.t1231 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3282 vdd2.t128 vn_p.t1371 out_n.t390 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3283 vdd2.t127 vn_p.t1372 out_n.t389 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3284 out_n.t86 vn_n.t276 vss.t86 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3285 vdd1.t135 vp_p.t1364 out_p.t1230 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3286 out_n.t388 vn_p.t1373 vdd2.t126 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3287 out_n.t387 vn_p.t1374 vdd2.t125 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3288 vdd2.t124 vn_p.t1375 out_n.t386 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3289 out_n.t385 vn_p.t1376 vdd2.t123 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3290 out_p.t101 vp_n.t271 vss.t290 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3291 vdd2.t122 vn_p.t1377 out_n.t384 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3292 vdd1.t134 vp_p.t1365 out_p.t1229 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3293 vdd2.t121 vn_p.t1378 out_n.t383 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3294 vdd2.t120 vn_p.t1379 out_n.t382 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3295 out_n.t87 vn_n.t277 vss.t87 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3296 vdd2.t119 vn_p.t1380 out_n.t381 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3297 vdd2.t118 vn_p.t1381 out_n.t380 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3298 vss.t289 vp_n.t272 out_p.t102 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3299 vss.t88 vn_n.t278 out_n.t88 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3300 out_p.t103 vp_n.t273 vss.t288 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3301 vdd2.t117 vn_p.t1382 out_n.t379 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3302 vdd1.t133 vp_p.t1366 out_p.t1228 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3303 out_p.t1227 vp_p.t1367 vdd1.t132 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3304 vdd1.t131 vp_p.t1368 out_p.t1226 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3305 vdd1.t130 vp_p.t1369 out_p.t1225 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3306 out_n.t378 vn_p.t1383 vdd2.t116 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3307 out_n.t1762 vn_n.t279 vss.t562 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3308 out_p.t1224 vp_p.t1370 vdd1.t129 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3309 vss.t563 vn_n.t280 out_n.t1763 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3310 vdd2.t115 vn_p.t1384 out_n.t377 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3311 out_n.t376 vn_p.t1385 vdd2.t114 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3312 vdd1.t128 vp_p.t1371 out_p.t1223 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3313 out_n.t375 vn_p.t1386 vdd2.t113 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3314 out_p.t1222 vp_p.t1372 vdd1.t127 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3315 vdd1.t126 vp_p.t1373 out_p.t1221 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3316 out_p.t1220 vp_p.t1374 vdd1.t125 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3317 vdd1.t124 vp_p.t1375 out_p.t1219 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3318 out_p.t1218 vp_p.t1376 vdd1.t123 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3319 out_n.t374 vn_p.t1387 vdd2.t112 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3320 vdd2.t111 vn_p.t1388 out_n.t373 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3321 vss.t287 vp_n.t274 out_p.t104 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3322 vdd1.t122 vp_p.t1377 out_p.t1217 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3323 out_n.t372 vn_p.t1389 vdd2.t110 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3324 vdd1.t121 vp_p.t1378 out_p.t1216 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3325 out_p.t1215 vp_p.t1379 vdd1.t120 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3326 vdd2.t109 vn_p.t1390 out_n.t371 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3327 out_n.t370 vn_p.t1391 vdd2.t108 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3328 vdd1.t119 vp_p.t1380 out_p.t1214 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3329 vdd1.t118 vp_p.t1381 out_p.t1213 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3330 vss.t564 vn_n.t281 out_n.t1764 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3331 vdd2.t107 vn_p.t1392 out_n.t369 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3332 out_n.t368 vn_p.t1393 vdd2.t106 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3333 vdd1.t117 vp_p.t1382 out_p.t1212 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3334 vdd2.t105 vn_p.t1394 out_n.t367 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3335 out_p.t1211 vp_p.t1383 vdd1.t116 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3336 vdd1.t115 vp_p.t1384 out_p.t1210 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3337 out_p.t1209 vp_p.t1385 vdd1.t114 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3338 out_p.t1208 vp_p.t1386 vdd1.t113 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3339 vdd1.t112 vp_p.t1387 out_p.t1207 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3340 vdd2.t104 vn_p.t1395 out_n.t366 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3341 out_n.t365 vn_p.t1396 vdd2.t103 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3342 out_p.t1206 vp_p.t1388 vdd1.t111 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3343 vdd1.t110 vp_p.t1389 out_p.t1205 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3344 vdd1.t109 vp_p.t1390 out_p.t1204 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3345 out_n.t1765 vn_n.t282 vss.t565 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3346 out_p.t44 vp_n.t275 vss.t286 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3347 out_n.t364 vn_p.t1397 vdd2.t102 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3348 vdd2.t101 vn_p.t1398 out_n.t363 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3349 vdd1.t108 vp_p.t1391 out_p.t1203 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3350 vdd2.t100 vn_p.t1399 out_n.t362 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3351 out_p.t45 vp_n.t276 vss.t285 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3352 vdd2.t99 vn_p.t1400 out_n.t361 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3353 out_n.t360 vn_p.t1401 vdd2.t98 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3354 vdd2.t97 vn_p.t1402 out_n.t359 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3355 vdd1.t107 vp_p.t1392 out_p.t1202 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3356 out_p.t1201 vp_p.t1393 vdd1.t106 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3357 out_p.t1200 vp_p.t1394 vdd1.t105 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3358 vss.t566 vn_n.t283 out_n.t1766 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3359 out_n.t358 vn_p.t1403 vdd2.t96 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3360 vss.t284 vp_n.t277 out_p.t46 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3361 out_p.t47 vp_n.t278 vss.t283 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3362 out_p.t1199 vp_p.t1395 vdd1.t104 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3363 out_p.t1198 vp_p.t1396 vdd1.t103 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3364 out_n.t357 vn_p.t1404 vdd2.t95 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3365 out_n.t356 vn_p.t1405 vdd2.t94 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3366 vss.t567 vn_n.t284 out_n.t1767 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3367 vss.t282 vp_n.t279 out_p.t48 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3368 vdd2.t93 vn_p.t1406 out_n.t355 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3369 vdd2.t92 vn_p.t1407 out_n.t354 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3370 out_n.t353 vn_p.t1408 vdd2.t91 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3371 vdd2.t90 vn_p.t1409 out_n.t352 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3372 out_n.t351 vn_p.t1410 vdd2.t89 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3373 vss.t281 vp_n.t280 out_p.t49 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3374 vdd2.t88 vn_p.t1411 out_n.t350 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3375 out_n.t349 vn_p.t1412 vdd2.t87 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3376 out_p.t1197 vp_p.t1397 vdd1.t102 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3377 vdd1.t101 vp_p.t1398 out_p.t1196 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3378 out_p.t1195 vp_p.t1399 vdd1.t100 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3379 vdd1.t99 vp_p.t1400 out_p.t1194 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3380 vdd2.t86 vn_p.t1413 out_n.t348 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3381 out_p.t1193 vp_p.t1401 vdd1.t98 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3382 out_p.t1192 vp_p.t1402 vdd1.t97 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3383 vdd1.t96 vp_p.t1403 out_p.t1191 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3384 out_p.t1190 vp_p.t1404 vdd1.t95 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3385 out_p.t1189 vp_p.t1405 vdd1.t94 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3386 vdd1.t93 vp_p.t1406 out_p.t1188 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3387 vdd1.t92 vp_p.t1407 out_p.t1187 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3388 out_n.t1768 vn_n.t285 vss.t568 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3389 vdd2.t85 vn_p.t1414 out_n.t347 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3390 vdd1.t91 vp_p.t1408 out_p.t1186 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3391 out_p.t50 vp_n.t281 vss.t280 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3392 vdd1.t90 vp_p.t1409 out_p.t1185 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3393 vdd1.t89 vp_p.t1410 out_p.t1184 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3394 vdd2.t84 vn_p.t1415 out_n.t346 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3395 vdd2.t83 vn_p.t1416 out_n.t345 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3396 out_n.t344 vn_p.t1417 vdd2.t82 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3397 out_p.t1183 vp_p.t1411 vdd1.t88 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3398 vdd2.t81 vn_p.t1418 out_n.t343 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3399 out_p.t1182 vp_p.t1412 vdd1.t87 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3400 vdd2.t80 vn_p.t1419 out_n.t342 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3401 out_n.t341 vn_p.t1420 vdd2.t79 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3402 vdd1.t86 vp_p.t1413 out_p.t1181 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3403 vdd1.t85 vp_p.t1414 out_p.t1180 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3404 vss.t569 vn_n.t286 out_n.t1769 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3405 out_n.t340 vn_p.t1421 vdd2.t78 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3406 vdd1.t84 vp_p.t1415 out_p.t1179 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3407 vdd1.t83 vp_p.t1416 out_p.t1178 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3408 out_p.t1177 vp_p.t1417 vdd1.t82 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3409 vdd1.t81 vp_p.t1418 out_p.t1176 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3410 vdd1.t80 vp_p.t1419 out_p.t1175 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3411 out_p.t1174 vp_p.t1420 vdd1.t79 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3412 out_n.t1788 vn_n.t287 vss.t588 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3413 vss.t589 vn_n.t288 out_n.t1789 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3414 out_p.t1173 vp_p.t1421 vdd1.t78 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3415 vss.t279 vp_n.t282 out_p.t51 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3416 out_n.t339 vn_p.t1422 vdd2.t77 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3417 vdd2.t76 vn_p.t1423 out_n.t338 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3418 out_n.t337 vn_p.t1424 vdd2.t75 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3419 out_n.t336 vn_p.t1425 vdd2.t74 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3420 vdd1.t77 vp_p.t1422 out_p.t1172 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3421 out_p.t1171 vp_p.t1423 vdd1.t76 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3422 vdd2.t73 vn_p.t1426 out_n.t335 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3423 out_n.t334 vn_p.t1427 vdd2.t72 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3424 vss.t278 vp_n.t283 out_p.t52 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3425 vdd2.t71 vn_p.t1428 out_n.t333 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3426 vdd1.t75 vp_p.t1424 out_p.t1170 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3427 vdd2.t70 vn_p.t1429 out_n.t332 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3428 out_n.t331 vn_p.t1430 vdd2.t69 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3429 out_n.t330 vn_p.t1431 vdd2.t68 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3430 out_n.t329 vn_p.t1432 vdd2.t67 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3431 vss.t277 vp_n.t284 out_p.t53 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3432 out_n.t328 vn_p.t1433 vdd2.t66 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3433 out_p.t54 vp_n.t285 vss.t276 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3434 vdd2.t65 vn_p.t1434 out_n.t327 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3435 out_n.t1790 vn_n.t289 vss.t590 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3436 vdd2.t64 vn_p.t1435 out_n.t326 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3437 out_p.t1169 vp_p.t1425 vdd1.t74 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3438 out_p.t1168 vp_p.t1426 vdd1.t73 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3439 vdd1.t72 vp_p.t1427 out_p.t1167 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3440 out_p.t1166 vp_p.t1428 vdd1.t71 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3441 vdd1.t70 vp_p.t1429 out_p.t1165 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3442 vdd1.t69 vp_p.t1430 out_p.t1164 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3443 out_n.t325 vn_p.t1436 vdd2.t63 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3444 out_p.t1163 vp_p.t1431 vdd1.t68 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3445 vdd1.t67 vp_p.t1432 out_p.t1162 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3446 out_p.t1161 vp_p.t1433 vdd1.t66 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3447 vdd2.t62 vn_p.t1437 out_n.t324 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3448 out_p.t1160 vp_p.t1434 vdd1.t65 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3449 vdd1.t64 vp_p.t1435 out_p.t1159 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3450 out_p.t1158 vp_p.t1436 vdd1.t63 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3451 out_p.t1157 vp_p.t1437 vdd1.t62 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3452 out_p.t1156 vp_p.t1438 vdd1.t61 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3453 vdd1.t60 vp_p.t1439 out_p.t1155 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3454 vss.t275 vp_n.t286 out_p.t55 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3455 out_p.t1154 vp_p.t1440 vdd1.t59 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3456 out_p.t1153 vp_p.t1441 vdd1.t58 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3457 out_n.t323 vn_p.t1438 vdd2.t61 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3458 vdd2.t60 vn_p.t1439 out_n.t322 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3459 out_n.t321 vn_p.t1440 vdd2.t59 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3460 out_p.t1152 vp_p.t1442 vdd1.t57 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3461 out_n.t320 vn_p.t1441 vdd2.t58 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3462 vdd1.t56 vp_p.t1443 out_p.t1151 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3463 vdd1.t55 vp_p.t1444 out_p.t1150 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3464 vss.t274 vp_n.t287 out_p.t56 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3465 vss.t591 vn_n.t290 out_n.t1791 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3466 out_n.t1792 vn_n.t291 vss.t592 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3467 out_p.t1149 vp_p.t1445 vdd1.t54 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3468 vss.t593 vn_n.t292 out_n.t1793 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3469 out_p.t1148 vp_p.t1446 vdd1.t53 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3470 out_p.t1147 vp_p.t1447 vdd1.t52 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3471 vdd1.t51 vp_p.t1448 out_p.t1146 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3472 out_n.t319 vn_p.t1442 vdd2.t57 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3473 vdd2.t56 vn_p.t1443 out_n.t318 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3474 out_n.t317 vn_p.t1444 vdd2.t55 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3475 out_p.t1145 vp_p.t1449 vdd1.t50 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3476 vdd2.t54 vn_p.t1445 out_n.t316 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3477 vdd1.t49 vp_p.t1450 out_p.t1144 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3478 out_n.t315 vn_p.t1446 vdd2.t53 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3479 vdd2.t52 vn_p.t1447 out_n.t314 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3480 out_n.t313 vn_p.t1448 vdd2.t51 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3481 vdd2.t50 vn_p.t1449 out_n.t312 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3482 vdd1.t48 vp_p.t1451 out_p.t1143 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3483 out_n.t311 vn_p.t1450 vdd2.t49 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3484 out_p.t57 vp_n.t288 vss.t273 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3485 out_p.t1142 vp_p.t1452 vdd1.t47 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3486 vdd2.t48 vn_p.t1451 out_n.t310 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3487 vdd2.t47 vn_p.t1452 out_n.t309 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3488 vdd2.t46 vn_p.t1453 out_n.t308 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3489 vdd1.t46 vp_p.t1453 out_p.t1141 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3490 vdd1.t45 vp_p.t1454 out_p.t1140 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3491 out_p.t1139 vp_p.t1455 vdd1.t44 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3492 out_n.t307 vn_p.t1454 vdd2.t45 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3493 out_p.t1138 vp_p.t1456 vdd1.t43 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3494 out_n.t306 vn_p.t1455 vdd2.t44 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3495 vdd2.t43 vn_p.t1456 out_n.t305 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3496 out_p.t58 vp_n.t289 vss.t272 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3497 out_p.t1137 vp_p.t1457 vdd1.t42 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3498 vdd1.t41 vp_p.t1458 out_p.t1136 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3499 vdd1.t40 vp_p.t1459 out_p.t1135 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3500 vss.t594 vn_n.t293 out_n.t1794 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3501 vdd2.t42 vn_p.t1457 out_n.t304 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3502 vss.t271 vp_n.t290 out_p.t59 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3503 vdd1.t39 vp_p.t1460 out_p.t1134 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3504 out_n.t303 vn_p.t1458 vdd2.t41 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3505 vdd2.t40 vn_p.t1459 out_n.t302 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3506 vss.t270 vp_n.t291 out_p.t60 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3507 out_n.t301 vn_p.t1460 vdd2.t39 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3508 out_p.t1133 vp_p.t1461 vdd1.t38 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3509 vdd1.t37 vp_p.t1462 out_p.t1132 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3510 out_p.t1131 vp_p.t1463 vdd1.t36 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3511 out_p.t1130 vp_p.t1464 vdd1.t35 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3512 out_p.t1129 vp_p.t1465 vdd1.t34 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3513 out_n.t300 vn_p.t1461 vdd2.t38 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3514 out_n.t299 vn_p.t1462 vdd2.t37 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3515 vdd1.t33 vp_p.t1466 out_p.t1128 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3516 vdd1.t32 vp_p.t1467 out_p.t1127 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3517 vdd1.t31 vp_p.t1468 out_p.t1126 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3518 out_n.t298 vn_p.t1463 vdd2.t36 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3519 out_p.t61 vp_n.t292 vss.t269 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3520 out_p.t62 vp_n.t293 vss.t268 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3521 out_p.t1125 vp_p.t1469 vdd1.t30 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3522 vdd1.t29 vp_p.t1470 out_p.t1124 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3523 vdd1.t28 vp_p.t1471 out_p.t1123 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3524 out_n.t1795 vn_n.t294 vss.t595 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3525 vdd2.t35 vn_p.t1464 out_n.t297 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3526 out_n.t296 vn_p.t1465 vdd2.t34 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3527 vss.t267 vp_n.t294 out_p.t63 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3528 vdd1.t27 vp_p.t1472 out_p.t1122 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3529 vdd2.t33 vn_p.t1466 out_n.t295 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3530 vdd2.t32 vn_p.t1467 out_n.t294 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3531 out_n.t293 vn_p.t1468 vdd2.t31 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3532 out_p.t1121 vp_p.t1473 vdd1.t26 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3533 vdd2.t30 vn_p.t1469 out_n.t292 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3534 vdd1.t25 vp_p.t1474 out_p.t1120 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3535 vdd2.t29 vn_p.t1470 out_n.t291 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3536 vdd2.t28 vn_p.t1471 out_n.t290 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3537 vdd2.t27 vn_p.t1472 out_n.t289 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3538 vdd2.t26 vn_p.t1473 out_n.t288 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3539 vdd2.t25 vn_p.t1474 out_n.t287 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3540 vdd2.t24 vn_p.t1475 out_n.t286 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3541 out_p.t1119 vp_p.t1475 vdd1.t24 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3542 vdd2.t23 vn_p.t1476 out_n.t285 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3543 vss.t266 vp_n.t295 out_p.t39 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3544 out_n.t242 vn_n.t295 vss.t242 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3545 out_n.t284 vn_p.t1477 vdd2.t22 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3546 out_n.t283 vn_p.t1478 vdd2.t21 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3547 vdd2.t20 vn_p.t1479 out_n.t282 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3548 vss.t243 vn_n.t296 out_n.t243 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3549 out_n.t281 vn_p.t1480 vdd2.t19 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3550 out_n.t280 vn_p.t1481 vdd2.t18 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3551 vdd2.t17 vn_p.t1482 out_n.t279 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3552 out_n.t278 vn_p.t1483 vdd2.t16 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3553 out_n.t277 vn_p.t1484 vdd2.t15 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3554 vdd1.t23 vp_p.t1476 out_p.t1118 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3555 out_p.t1117 vp_p.t1477 vdd1.t22 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3556 out_n.t276 vn_p.t1485 vdd2.t14 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3557 vdd1.t21 vp_p.t1478 out_p.t1116 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3558 out_n.t275 vn_p.t1486 vdd2.t13 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3559 vdd1.t20 vp_p.t1479 out_p.t1115 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3560 out_n.t274 vn_p.t1487 vdd2.t12 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3561 vdd1.t19 vp_p.t1480 out_p.t1114 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3562 out_n.t244 vn_n.t297 vss.t244 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3563 vss.t245 vn_n.t298 out_n.t245 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3564 vdd2.t11 vn_p.t1488 out_n.t273 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3565 out_n.t272 vn_p.t1489 vdd2.t10 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3566 out_p.t1113 vp_p.t1481 vdd1.t18 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3567 vdd2.t9 vn_p.t1490 out_n.t271 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3568 out_n.t270 vn_p.t1491 vdd2.t8 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3569 out_n.t269 vn_p.t1492 vdd2.t7 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3570 out_p.t1112 vp_p.t1482 vdd1.t17 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3571 out_p.t40 vp_n.t296 vss.t265 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3572 vdd2.t6 vn_p.t1493 out_n.t268 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3573 vdd1.t16 vp_p.t1483 out_p.t1111 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3574 vdd1.t15 vp_p.t1484 out_p.t1110 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3575 vdd1.t14 vp_p.t1485 out_p.t1109 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3576 out_n.t246 vn_n.t299 vss.t246 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3577 vdd2.t5 vn_p.t1494 out_n.t267 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3578 vdd1.t13 vp_p.t1486 out_p.t1108 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3579 out_p.t1107 vp_p.t1487 vdd1.t12 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3580 vdd2.t4 vn_p.t1495 out_n.t266 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3581 vdd1.t11 vp_p.t1488 out_p.t1106 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3582 out_p.t1105 vp_p.t1489 vdd1.t10 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3583 out_p.t41 vp_n.t297 vss.t264 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3584 out_p.t1104 vp_p.t1490 vdd1.t9 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3585 out_p.t1103 vp_p.t1491 vdd1.t8 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3586 vdd2.t3 vn_p.t1496 out_n.t265 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3587 vdd2.t2 vn_p.t1497 out_n.t264 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3588 vdd1.t7 vp_p.t1492 out_p.t1102 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3589 out_n.t263 vn_p.t1498 vdd2.t1 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3590 vss.t263 vp_n.t298 out_p.t42 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3591 vdd1.t6 vp_p.t1493 out_p.t1101 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3592 out_p.t1100 vp_p.t1494 vdd1.t5 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3593 vdd1.t4 vp_p.t1495 out_p.t1099 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3594 out_p.t1098 vp_p.t1496 vdd1.t3 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3595 vdd2.t0 vn_p.t1499 out_n.t262 vdd2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3596 out_p.t43 vp_n.t299 vss.t262 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3597 vdd1.t2 vp_p.t1497 out_p.t1097 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3598 out_p.t1096 vp_p.t1498 vdd1.t1 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3599 vdd1.t0 vp_p.t1499 out_p.t1095 vdd1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
C0 vdd1 vp_p 620.90fF
C1 vdd2 vn_p 620.90fF
C2 vdd1 out_p 4414.79fF
C3 vp_n out_p 102.35fF
C4 out_p vp_p 548.19fF
C5 vdd2 out_n 4414.79fF
C6 vn_p out_n 548.19fF
C7 out_n vn_n 102.36fF
R0 vn_p.n668 vn_p.t330 756.008
R1 vn_p.n668 vn_p.t99 756.008
R2 vn_p.n666 vn_p.t1483 756.008
R3 vn_p.n666 vn_p.t1242 756.008
R4 vn_p.n664 vn_p.t529 756.008
R5 vn_p.n664 vn_p.t287 756.008
R6 vn_p.n662 vn_p.t193 756.008
R7 vn_p.n662 vn_p.t1442 756.008
R8 vn_p.n660 vn_p.t1383 756.008
R9 vn_p.n660 vn_p.t1137 756.008
R10 vn_p.n658 vn_p.t1033 756.008
R11 vn_p.n658 vn_p.t797 756.008
R12 vn_p.n656 vn_p.t687 756.008
R13 vn_p.n656 vn_p.t454 756.008
R14 vn_p.n654 vn_p.t1225 756.008
R15 vn_p.n654 vn_p.t994 756.008
R16 vn_p.n652 vn_p.t884 756.008
R17 vn_p.n652 vn_p.t642 756.008
R18 vn_p.n650 vn_p.t574 756.008
R19 vn_p.n650 vn_p.t331 756.008
R20 vn_p.n648 vn_p.t232 756.008
R21 vn_p.n648 vn_p.t1485 756.008
R22 vn_p.n646 vn_p.t776 756.008
R23 vn_p.n646 vn_p.t530 756.008
R24 vn_p.n644 vn_p.t432 756.008
R25 vn_p.n644 vn_p.t195 756.008
R26 vn_p.n642 vn_p.t83 756.008
R27 vn_p.n642 vn_p.t1345 756.008
R28 vn_p.n640 vn_p.t1268 756.008
R29 vn_p.n640 vn_p.t1034 756.008
R30 vn_p.n638 vn_p.t921 756.008
R31 vn_p.n638 vn_p.t688 756.008
R32 vn_p.n636 vn_p.t1009 756.008
R33 vn_p.n636 vn_p.t771 756.008
R34 vn_p.n634 vn_p.t655 756.008
R35 vn_p.n634 vn_p.t425 756.008
R36 vn_p.n632 vn_p.t305 756.008
R37 vn_p.n632 vn_p.t77 756.008
R38 vn_p.n630 vn_p.t1498 756.008
R39 vn_p.n630 vn_p.t1264 756.008
R40 vn_p.n628 vn_p.t1153 756.008
R41 vn_p.n628 vn_p.t915 756.008
R42 vn_p.n626 vn_p.t207 756.008
R43 vn_p.n626 vn_p.t1458 756.008
R44 vn_p.n624 vn_p.t1363 756.008
R45 vn_p.n624 vn_p.t1113 756.008
R46 vn_p.n622 vn_p.t400 756.008
R47 vn_p.n622 vn_p.t170 756.008
R48 vn_p.n620 vn_p.t700 756.008
R49 vn_p.n620 vn_p.t468 756.008
R50 vn_p.n618 vn_p.t346 756.008
R51 vn_p.n618 vn_p.t118 756.008
R52 vn_p.n616 vn_p.t897 756.008
R53 vn_p.n616 vn_p.t656 756.008
R54 vn_p.n614 vn_p.t548 756.008
R55 vn_p.n614 vn_p.t306 756.008
R56 vn_p.n612 vn_p.t1091 756.008
R57 vn_p.n612 vn_p.t863 756.008
R58 vn_p.n610 vn_p.t1401 756.008
R59 vn_p.n610 vn_p.t1155 756.008
R60 vn_p.n608 vn_p.t447 756.008
R61 vn_p.n608 vn_p.t208 756.008
R62 vn_p.n606 vn_p.t101 756.008
R63 vn_p.n606 vn_p.t1364 756.008
R64 vn_p.n604 vn_p.t1244 756.008
R65 vn_p.n604 vn_p.t1015 756.008
R66 vn_p.n602 vn_p.t288 756.008
R67 vn_p.n602 vn_p.t59 756.008
R68 vn_p.n600 vn_p.t595 756.008
R69 vn_p.n600 vn_p.t351 756.008
R70 vn_p.n598 vn_p.t1138 756.008
R71 vn_p.n598 vn_p.t898 756.008
R72 vn_p.n596 vn_p.t800 756.008
R73 vn_p.n596 vn_p.t553 756.008
R74 vn_p.n594 vn_p.t453 756.008
R75 vn_p.n594 vn_p.t213 756.008
R76 vn_p.n592 vn_p.t995 756.008
R77 vn_p.n592 vn_p.t757 756.008
R78 vn_p.n590 vn_p.t1288 756.008
R79 vn_p.n590 vn_p.t1050 756.008
R80 vn_p.n588 vn_p.t980 756.008
R81 vn_p.n588 vn_p.t743 756.008
R82 vn_p.n586 vn_p.t631 756.008
R83 vn_p.n586 vn_p.t392 756.008
R84 vn_p.n584 vn_p.t1175 756.008
R85 vn_p.n584 vn_p.t943 756.008
R86 vn_p.n582 vn_p.t838 756.008
R87 vn_p.n582 vn_p.t599 756.008
R88 vn_p.n580 vn_p.t1127 756.008
R89 vn_p.n580 vn_p.t890 756.008
R90 vn_p.n578 vn_p.t180 756.008
R91 vn_p.n578 vn_p.t1436 756.008
R92 vn_p.n576 vn_p.t1330 756.008
R93 vn_p.n576 vn_p.t1086 756.008
R94 vn_p.n574 vn_p.t372 756.008
R95 vn_p.n574 vn_p.t144 756.008
R96 vn_p.n572 vn_p.t31 756.008
R97 vn_p.n572 vn_p.t1292 756.008
R98 vn_p.n570 vn_p.t1212 756.008
R99 vn_p.n570 vn_p.t984 756.008
R100 vn_p.n568 vn_p.t873 756.008
R101 vn_p.n568 vn_p.t633 756.008
R102 vn_p.n566 vn_p.t519 756.008
R103 vn_p.n566 vn_p.t284 756.008
R104 vn_p.n564 vn_p.t1068 756.008
R105 vn_p.n564 vn_p.t839 756.008
R106 vn_p.n562 vn_p.t730 756.008
R107 vn_p.n562 vn_p.t490 756.008
R108 vn_p.n560 vn_p.t420 756.008
R109 vn_p.n560 vn_p.t183 756.008
R110 vn_p.n558 vn_p.t73 756.008
R111 vn_p.n558 vn_p.t1331 756.008
R112 vn_p.n556 vn_p.t1217 756.008
R113 vn_p.n556 vn_p.t990 756.008
R114 vn_p.n554 vn_p.t265 756.008
R115 vn_p.n554 vn_p.t34 756.008
R116 vn_p.n552 vn_p.t1422 756.008
R117 vn_p.n552 vn_p.t1180 756.008
R118 vn_p.n550 vn_p.t1109 756.008
R119 vn_p.n550 vn_p.t876 756.008
R120 vn_p.n548 vn_p.t769 756.008
R121 vn_p.n548 vn_p.t523 756.008
R122 vn_p.n546 vn_p.t1313 756.008
R123 vn_p.n546 vn_p.t1071 756.008
R124 vn_p.n544 vn_p.t969 756.008
R125 vn_p.n544 vn_p.t733 756.008
R126 vn_p.n542 vn_p.t620 756.008
R127 vn_p.n542 vn_p.t378 756.008
R128 vn_p.n540 vn_p.t955 756.008
R129 vn_p.n540 vn_p.t719 756.008
R130 vn_p.n538 vn_p.t609 756.008
R131 vn_p.n538 vn_p.t366 756.008
R132 vn_p.n536 vn_p.t1152 756.008
R133 vn_p.n536 vn_p.t917 756.008
R134 vn_p.n534 vn_p.t813 756.008
R135 vn_p.n534 vn_p.t573 756.008
R136 vn_p.n532 vn_p.t471 756.008
R137 vn_p.n532 vn_p.t228 756.008
R138 vn_p.n530 vn_p.t156 756.008
R139 vn_p.n530 vn_p.t1417 756.008
R140 vn_p.n528 vn_p.t1304 756.008
R141 vn_p.n528 vn_p.t1063 756.008
R142 vn_p.n526 vn_p.t347 756.008
R143 vn_p.n526 vn_p.t120 756.008
R144 vn_p.n524 vn_p.t3 756.008
R145 vn_p.n524 vn_p.t1266 756.008
R146 vn_p.n522 vn_p.t550 756.008
R147 vn_p.n522 vn_p.t308 756.008
R148 vn_p.n521 vn_p.t850 756.008
R149 vn_p.n521 vn_p.t611 756.008
R150 vn_p.n519 vn_p.t671 756.008
R151 vn_p.n519 vn_p.t1235 756.008
R152 vn_p.n517 vn_p.t1211 756.008
R153 vn_p.n517 vn_p.t283 756.008
R154 vn_p.n515 vn_p.t872 756.008
R155 vn_p.n515 vn_p.t1439 756.008
R156 vn_p.n513 vn_p.t1165 756.008
R157 vn_p.n513 vn_p.t242 756.008
R158 vn_p.n511 vn_p.t219 756.008
R159 vn_p.n511 vn_p.t790 756.008
R160 vn_p.n509 vn_p.t1377 756.008
R161 vn_p.n509 vn_p.t444 756.008
R162 vn_p.n507 vn_p.t418 756.008
R163 vn_p.n507 vn_p.t989 756.008
R164 vn_p.n505 vn_p.t72 756.008
R165 vn_p.n505 vn_p.t636 756.008
R166 vn_p.n503 vn_p.t1256 756.008
R167 vn_p.n503 vn_p.t322 756.008
R168 vn_p.n501 vn_p.t911 756.008
R169 vn_p.n501 vn_p.t1474 756.008
R170 vn_p.n499 vn_p.t566 756.008
R171 vn_p.n499 vn_p.t1134 756.008
R172 vn_p.n497 vn_p.t1108 756.008
R173 vn_p.n497 vn_p.t187 756.008
R174 vn_p.n495 vn_p.t767 756.008
R175 vn_p.n495 vn_p.t1334 756.008
R176 vn_p.n493 vn_p.t463 756.008
R177 vn_p.n493 vn_p.t1028 756.008
R178 vn_p.n491 vn_p.t114 756.008
R179 vn_p.n491 vn_p.t677 756.008
R180 vn_p.n489 vn_p.t1263 756.008
R181 vn_p.n489 vn_p.t327 756.008
R182 vn_p.n487 vn_p.t1347 756.008
R183 vn_p.n487 vn_p.t415 756.008
R184 vn_p.n485 vn_p.t1002 756.008
R185 vn_p.n485 vn_p.t70 756.008
R186 vn_p.n483 vn_p.t689 756.008
R187 vn_p.n483 vn_p.t1252 756.008
R188 vn_p.n481 vn_p.t337 756.008
R189 vn_p.n481 vn_p.t907 756.008
R190 vn_p.n479 vn_p.t886 756.008
R191 vn_p.n479 vn_p.t1451 756.008
R192 vn_p.n477 vn_p.t538 756.008
R193 vn_p.n477 vn_p.t1105 756.008
R194 vn_p.n475 vn_p.t200 756.008
R195 vn_p.n475 vn_p.t766 756.008
R196 vn_p.n473 vn_p.t1390 756.008
R197 vn_p.n473 vn_p.t459 756.008
R198 vn_p.n471 vn_p.t1039 756.008
R199 vn_p.n471 vn_p.t111 756.008
R200 vn_p.n469 vn_p.t86 756.008
R201 vn_p.n469 vn_p.t648 756.008
R202 vn_p.n467 vn_p.t1231 756.008
R203 vn_p.n467 vn_p.t300 756.008
R204 vn_p.n465 vn_p.t889 756.008
R205 vn_p.n465 vn_p.t1456 756.008
R206 vn_p.n463 vn_p.t581 756.008
R207 vn_p.n463 vn_p.t1147 756.008
R208 vn_p.n461 vn_p.t237 756.008
R209 vn_p.n461 vn_p.t807 756.008
R210 vn_p.n459 vn_p.t784 756.008
R211 vn_p.n459 vn_p.t1354 756.008
R212 vn_p.n457 vn_p.t439 756.008
R213 vn_p.n457 vn_p.t1007 756.008
R214 vn_p.n455 vn_p.t983 756.008
R215 vn_p.n455 vn_p.t51 756.008
R216 vn_p.n453 vn_p.t1275 756.008
R217 vn_p.n453 vn_p.t342 756.008
R218 vn_p.n451 vn_p.t930 756.008
R219 vn_p.n451 vn_p.t1495 756.008
R220 vn_p.n449 vn_p.t1471 756.008
R221 vn_p.n449 vn_p.t543 756.008
R222 vn_p.n447 vn_p.t1129 756.008
R223 vn_p.n447 vn_p.t204 756.008
R224 vn_p.n445 vn_p.t182 756.008
R225 vn_p.n445 vn_p.t749 756.008
R226 vn_p.n443 vn_p.t480 756.008
R227 vn_p.n443 vn_p.t1044 756.008
R228 vn_p.n441 vn_p.t171 756.008
R229 vn_p.n441 vn_p.t736 756.008
R230 vn_p.n439 vn_p.t1319 756.008
R231 vn_p.n439 vn_p.t383 756.008
R232 vn_p.n437 vn_p.t974 756.008
R233 vn_p.n437 vn_p.t43 756.008
R234 vn_p.n435 vn_p.t19 756.008
R235 vn_p.n435 vn_p.t589 756.008
R236 vn_p.n433 vn_p.t309 756.008
R237 vn_p.n433 vn_p.t883 756.008
R238 vn_p.n431 vn_p.t864 756.008
R239 vn_p.n431 vn_p.t1426 756.008
R240 vn_p.n429 vn_p.t510 756.008
R241 vn_p.n429 vn_p.t1079 756.008
R242 vn_p.n427 vn_p.t176 756.008
R243 vn_p.n427 vn_p.t741 756.008
R244 vn_p.n425 vn_p.t718 756.008
R245 vn_p.n425 vn_p.t1286 756.008
R246 vn_p.n423 vn_p.t1016 756.008
R247 vn_p.n423 vn_p.t81 756.008
R248 vn_p.n421 vn_p.t61 756.008
R249 vn_p.n421 vn_p.t624 756.008
R250 vn_p.n419 vn_p.t1203 756.008
R251 vn_p.n419 vn_p.t276 756.008
R252 vn_p.n417 vn_p.t257 756.008
R253 vn_p.n417 vn_p.t833 756.008
R254 vn_p.n415 vn_p.t1415 756.008
R255 vn_p.n415 vn_p.t488 756.008
R256 vn_p.n413 vn_p.t214 756.008
R257 vn_p.n413 vn_p.t779 756.008
R258 vn_p.n411 vn_p.t758 756.008
R259 vn_p.n411 vn_p.t1325 756.008
R260 vn_p.n409 vn_p.t408 756.008
R261 vn_p.n409 vn_p.t979 756.008
R262 vn_p.n407 vn_p.t957 756.008
R263 vn_p.n407 vn_p.t26 756.008
R264 vn_p.n405 vn_p.t612 756.008
R265 vn_p.n405 vn_p.t1173 756.008
R266 vn_p.n403 vn_p.t293 756.008
R267 vn_p.n403 vn_p.t870 756.008
R268 vn_p.n401 vn_p.t1449 756.008
R269 vn_p.n401 vn_p.t515 756.008
R270 vn_p.n399 vn_p.t1099 756.008
R271 vn_p.n399 vn_p.t179 756.008
R272 vn_p.n397 vn_p.t158 756.008
R273 vn_p.n397 vn_p.t724 756.008
R274 vn_p.n395 vn_p.t1306 756.008
R275 vn_p.n395 vn_p.t369 756.008
R276 vn_p.n393 vn_p.t145 756.008
R277 vn_p.n393 vn_p.t709 756.008
R278 vn_p.n391 vn_p.t1293 756.008
R279 vn_p.n391 vn_p.t357 756.008
R280 vn_p.n389 vn_p.t948 756.008
R281 vn_p.n389 vn_p.t17 756.008
R282 vn_p.n387 vn_p.t1490 756.008
R283 vn_p.n387 vn_p.t561 756.008
R284 vn_p.n385 vn_p.t1146 756.008
R285 vn_p.n385 vn_p.t222 756.008
R286 vn_p.n383 vn_p.t840 756.008
R287 vn_p.n383 vn_p.t1409 756.008
R288 vn_p.n381 vn_p.t492 756.008
R289 vn_p.n381 vn_p.t1057 756.008
R290 vn_p.n379 vn_p.t1038 756.008
R291 vn_p.n379 vn_p.t109 756.008
R292 vn_p.n377 vn_p.t696 756.008
R293 vn_p.n377 vn_p.t1260 756.008
R294 vn_p.n375 vn_p.t340 756.008
R295 vn_p.n375 vn_p.t912 756.008
R296 vn_p.n373 vn_p.t36 756.008
R297 vn_p.n373 vn_p.t605 756.008
R298 vn_p.n372 vn_p.t1179 756.008
R299 vn_p.n372 vn_p.t253 756.008
R300 vn_p.n370 vn_p.t662 756.008
R301 vn_p.n370 vn_p.t1226 756.008
R302 vn_p.n368 vn_p.t313 756.008
R303 vn_p.n368 vn_p.t885 756.008
R304 vn_p.n366 vn_p.t868 756.008
R305 vn_p.n366 vn_p.t1431 756.008
R306 vn_p.n364 vn_p.t512 756.008
R307 vn_p.n364 vn_p.t1080 756.008
R308 vn_p.n362 vn_p.t211 756.008
R309 vn_p.n362 vn_p.t778 756.008
R310 vn_p.n360 vn_p.t1368 756.008
R311 vn_p.n360 vn_p.t433 756.008
R312 vn_p.n358 vn_p.t1021 756.008
R313 vn_p.n358 vn_p.t85 756.008
R314 vn_p.n356 vn_p.t65 756.008
R315 vn_p.n356 vn_p.t628 756.008
R316 vn_p.n354 vn_p.t1208 756.008
R317 vn_p.n354 vn_p.t278 756.008
R318 vn_p.n352 vn_p.t902 756.008
R319 vn_p.n352 vn_p.t1463 756.008
R320 vn_p.n350 vn_p.t556 756.008
R321 vn_p.n350 vn_p.t1122 756.008
R322 vn_p.n348 vn_p.t1097 756.008
R323 vn_p.n348 vn_p.t177 756.008
R324 vn_p.n346 vn_p.t761 756.008
R325 vn_p.n346 vn_p.t1326 756.008
R326 vn_p.n344 vn_p.t414 756.008
R327 vn_p.n344 vn_p.t981 756.008
R328 vn_p.n342 vn_p.t106 756.008
R329 vn_p.n342 vn_p.t666 756.008
R330 vn_p.n340 vn_p.t1251 756.008
R331 vn_p.n340 vn_p.t318 756.008
R332 vn_p.n338 vn_p.t1337 756.008
R333 vn_p.n338 vn_p.t402 756.008
R334 vn_p.n336 vn_p.t993 756.008
R335 vn_p.n336 vn_p.t60 756.008
R336 vn_p.n334 vn_p.t639 756.008
R337 vn_p.n334 vn_p.t1202 756.008
R338 vn_p.n332 vn_p.t328 756.008
R339 vn_p.n332 vn_p.t899 756.008
R340 vn_p.n330 vn_p.t1481 756.008
R341 vn_p.n330 vn_p.t552 756.008
R342 vn_p.n328 vn_p.t527 756.008
R343 vn_p.n328 vn_p.t1093 756.008
R344 vn_p.n326 vn_p.t191 756.008
R345 vn_p.n326 vn_p.t756 756.008
R346 vn_p.n324 vn_p.t737 756.008
R347 vn_p.n324 vn_p.t1302 756.008
R348 vn_p.n322 vn_p.t1031 756.008
R349 vn_p.n322 vn_p.t103 756.008
R350 vn_p.n320 vn_p.t685 756.008
R351 vn_p.n320 vn_p.t1247 756.008
R352 vn_p.n318 vn_p.t1222 756.008
R353 vn_p.n318 vn_p.t291 756.008
R354 vn_p.n316 vn_p.t881 756.008
R355 vn_p.n316 vn_p.t1448 756.008
R356 vn_p.n314 vn_p.t1427 756.008
R357 vn_p.n314 vn_p.t498 756.008
R358 vn_p.n312 vn_p.t230 756.008
R359 vn_p.n312 vn_p.t802 756.008
R360 vn_p.n310 vn_p.t774 756.008
R361 vn_p.n310 vn_p.t1341 756.008
R362 vn_p.n308 vn_p.t430 756.008
R363 vn_p.n308 vn_p.t999 756.008
R364 vn_p.n306 vn_p.t82 756.008
R365 vn_p.n306 vn_p.t645 756.008
R366 vn_p.n304 vn_p.t625 756.008
R367 vn_p.n304 vn_p.t1189 756.008
R368 vn_p.n302 vn_p.t920 756.008
R369 vn_p.n302 vn_p.t1486 756.008
R370 vn_p.n300 vn_p.t1462 756.008
R371 vn_p.n300 vn_p.t534 756.008
R372 vn_p.n298 vn_p.t1118 756.008
R373 vn_p.n298 vn_p.t198 756.008
R374 vn_p.n296 vn_p.t780 756.008
R375 vn_p.n296 vn_p.t1350 756.008
R376 vn_p.n294 vn_p.t1324 756.008
R377 vn_p.n294 vn_p.t388 756.008
R378 vn_p.n292 vn_p.t124 756.008
R379 vn_p.n292 vn_p.t690 756.008
R380 vn_p.n290 vn_p.t1310 756.008
R381 vn_p.n290 vn_p.t374 756.008
R382 vn_p.n288 vn_p.t967 756.008
R383 vn_p.n288 vn_p.t33 756.008
R384 vn_p.n286 vn_p.t11 756.008
R385 vn_p.n286 vn_p.t580 756.008
R386 vn_p.n284 vn_p.t1162 756.008
R387 vn_p.n284 vn_p.t236 756.008
R388 vn_p.n282 vn_p.t1455 756.008
R389 vn_p.n282 vn_p.t520 756.008
R390 vn_p.n280 vn_p.t504 756.008
R391 vn_p.n280 vn_p.t1070 756.008
R392 vn_p.n278 vn_p.t166 756.008
R393 vn_p.n278 vn_p.t732 756.008
R394 vn_p.n276 vn_p.t710 756.008
R395 vn_p.n276 vn_p.t1274 756.008
R396 vn_p.n274 vn_p.t358 756.008
R397 vn_p.n274 vn_p.t929 756.008
R398 vn_p.n272 vn_p.t50 756.008
R399 vn_p.n272 vn_p.t617 756.008
R400 vn_p.n270 vn_p.t1196 756.008
R401 vn_p.n270 vn_p.t268 756.008
R402 vn_p.n268 vn_p.t860 756.008
R403 vn_p.n268 vn_p.t1424 756.008
R404 vn_p.n266 vn_p.t1410 756.008
R405 vn_p.n266 vn_p.t479 756.008
R406 vn_p.n264 vn_p.t1055 756.008
R407 vn_p.n264 vn_p.t131 756.008
R408 vn_p.n262 vn_p.t748 756.008
R409 vn_p.n262 vn_p.t1315 756.008
R410 vn_p.n260 vn_p.t398 756.008
R411 vn_p.n260 vn_p.t971 756.008
R412 vn_p.n258 vn_p.t56 756.008
R413 vn_p.n258 vn_p.t621 756.008
R414 vn_p.n256 vn_p.t603 756.008
R415 vn_p.n256 vn_p.t1168 756.008
R416 vn_p.n254 vn_p.t254 756.008
R417 vn_p.n254 vn_p.t829 756.008
R418 vn_p.n252 vn_p.t1441 756.008
R419 vn_p.n252 vn_p.t507 756.008
R420 vn_p.n250 vn_p.t1090 756.008
R421 vn_p.n250 vn_p.t172 756.008
R422 vn_p.n248 vn_p.t149 756.008
R423 vn_p.n248 vn_p.t715 756.008
R424 vn_p.n246 vn_p.t1298 756.008
R425 vn_p.n246 vn_p.t363 756.008
R426 vn_p.n244 vn_p.t951 756.008
R427 vn_p.n244 vn_p.t20 756.008
R428 vn_p.n242 vn_p.t1285 756.008
R429 vn_p.n242 vn_p.t350 756.008
R430 vn_p.n240 vn_p.t940 756.008
R431 vn_p.n240 vn_p.t4 756.008
R432 vn_p.n238 vn_p.t1480 756.008
R433 vn_p.n238 vn_p.t551 756.008
R434 vn_p.n236 vn_p.t1141 756.008
R435 vn_p.n236 vn_p.t212 756.008
R436 vn_p.n234 vn_p.t801 756.008
R437 vn_p.n234 vn_p.t1369 756.008
R438 vn_p.n232 vn_p.t487 756.008
R439 vn_p.n232 vn_p.t1048 756.008
R440 vn_p.n230 vn_p.t142 756.008
R441 vn_p.n230 vn_p.t703 756.008
R442 vn_p.n228 vn_p.t684 756.008
R443 vn_p.n228 vn_p.t1246 756.008
R444 vn_p.n226 vn_p.t333 756.008
R445 vn_p.n226 vn_p.t903 756.008
R446 vn_p.n224 vn_p.t880 756.008
R447 vn_p.n224 vn_p.t1446 756.008
R448 vn_p.n223 vn_p.t1172 756.008
R449 vn_p.n223 vn_p.t247 756.008
R450 vn_p.n221 vn_p.t302 756.008
R451 vn_p.n221 vn_p.t74 756.008
R452 vn_p.n219 vn_p.t857 756.008
R453 vn_p.n219 vn_p.t616 756.008
R454 vn_p.n217 vn_p.t505 756.008
R455 vn_p.n217 vn_p.t267 756.008
R456 vn_p.n215 vn_p.t810 756.008
R457 vn_p.n215 vn_p.t568 756.008
R458 vn_p.n213 vn_p.t1358 756.008
R459 vn_p.n213 vn_p.t1110 756.008
R460 vn_p.n211 vn_p.t1010 756.008
R461 vn_p.n211 vn_p.t770 756.008
R462 vn_p.n209 vn_p.t55 756.008
R463 vn_p.n209 vn_p.t1314 756.008
R464 vn_p.n207 vn_p.t1197 756.008
R465 vn_p.n207 vn_p.t970 756.008
R466 vn_p.n205 vn_p.t894 756.008
R467 vn_p.n205 vn_p.t652 756.008
R468 vn_p.n203 vn_p.t544 756.008
R469 vn_p.n203 vn_p.t303 756.008
R470 vn_p.n201 vn_p.t206 756.008
R471 vn_p.n201 vn_p.t1457 756.008
R472 vn_p.n199 vn_p.t751 756.008
R473 vn_p.n199 vn_p.t506 756.008
R474 vn_p.n197 vn_p.t399 756.008
R475 vn_p.n197 vn_p.t169 756.008
R476 vn_p.n195 vn_p.t95 756.008
R477 vn_p.n195 vn_p.t1359 756.008
R478 vn_p.n193 vn_p.t1239 756.008
R479 vn_p.n193 vn_p.t1011 756.008
R480 vn_p.n191 vn_p.t896 756.008
R481 vn_p.n191 vn_p.t658 756.008
R482 vn_p.n189 vn_p.t982 756.008
R483 vn_p.n189 vn_p.t745 756.008
R484 vn_p.n187 vn_p.t632 756.008
R485 vn_p.n187 vn_p.t393 756.008
R486 vn_p.n185 vn_p.t320 756.008
R487 vn_p.n185 vn_p.t88 756.008
R488 vn_p.n183 vn_p.t1470 756.008
R489 vn_p.n183 vn_p.t1233 756.008
R490 vn_p.n181 vn_p.t516 756.008
R491 vn_p.n181 vn_p.t279 756.008
R492 vn_p.n179 vn_p.t181 756.008
R493 vn_p.n179 vn_p.t1437 756.008
R494 vn_p.n177 vn_p.t1332 756.008
R495 vn_p.n177 vn_p.t1087 756.008
R496 vn_p.n175 vn_p.t1025 756.008
R497 vn_p.n175 vn_p.t787 756.008
R498 vn_p.n173 vn_p.t674 756.008
R499 vn_p.n173 vn_p.t442 756.008
R500 vn_p.n171 vn_p.t1214 756.008
R501 vn_p.n171 vn_p.t986 756.008
R502 vn_p.n169 vn_p.t875 756.008
R503 vn_p.n169 vn_p.t634 756.008
R504 vn_p.n167 vn_p.t521 756.008
R505 vn_p.n167 vn_p.t286 756.008
R506 vn_p.n165 vn_p.t223 756.008
R507 vn_p.n165 vn_p.t1472 756.008
R508 vn_p.n163 vn_p.t1379 756.008
R509 vn_p.n163 vn_p.t1131 756.008
R510 vn_p.n161 vn_p.t422 756.008
R511 vn_p.n161 vn_p.t184 756.008
R512 vn_p.n159 vn_p.t75 756.008
R513 vn_p.n159 vn_p.t1333 756.008
R514 vn_p.n157 vn_p.t618 756.008
R515 vn_p.n157 vn_p.t376 756.008
R516 vn_p.n155 vn_p.t913 756.008
R517 vn_p.n155 vn_p.t676 756.008
R518 vn_p.n153 vn_p.t569 756.008
R519 vn_p.n153 vn_p.t324 756.008
R520 vn_p.n151 vn_p.t1111 756.008
R521 vn_p.n151 vn_p.t877 756.008
R522 vn_p.n149 vn_p.t772 756.008
R523 vn_p.n149 vn_p.t522 756.008
R524 vn_p.n147 vn_p.t1316 756.008
R525 vn_p.n147 vn_p.t1073 756.008
R526 vn_p.n145 vn_p.t115 756.008
R527 vn_p.n145 vn_p.t1381 756.008
R528 vn_p.n143 vn_p.t1301 756.008
R529 vn_p.n143 vn_p.t1060 756.008
R530 vn_p.n141 vn_p.t956 756.008
R531 vn_p.n141 vn_p.t720 756.008
R532 vn_p.n139 vn_p.t610 756.008
R533 vn_p.n139 vn_p.t367 756.008
R534 vn_p.n137 vn_p.t1154 756.008
R535 vn_p.n137 vn_p.t918 756.008
R536 vn_p.n135 vn_p.t1447 756.008
R537 vn_p.n135 vn_p.t1205 756.008
R538 vn_p.n133 vn_p.t497 756.008
R539 vn_p.n133 vn_p.t259 756.008
R540 vn_p.n131 vn_p.t157 756.008
R541 vn_p.n131 vn_p.t1418 756.008
R542 vn_p.n129 vn_p.t1305 756.008
R543 vn_p.n129 vn_p.t1064 756.008
R544 vn_p.n127 vn_p.t348 756.008
R545 vn_p.n127 vn_p.t122 756.008
R546 vn_p.n125 vn_p.t646 756.008
R547 vn_p.n125 vn_p.t411 756.008
R548 vn_p.n123 vn_p.t1188 756.008
R549 vn_p.n123 vn_p.t958 756.008
R550 vn_p.n121 vn_p.t852 756.008
R551 vn_p.n121 vn_p.t613 756.008
R552 vn_p.n119 vn_p.t1402 756.008
R553 vn_p.n119 vn_p.t1157 756.008
R554 vn_p.n117 vn_p.t1049 756.008
R555 vn_p.n117 vn_p.t816 756.008
R556 vn_p.n115 vn_p.t1349 756.008
R557 vn_p.n115 vn_p.t1101 756.008
R558 vn_p.n113 vn_p.t389 756.008
R559 vn_p.n113 vn_p.t159 756.008
R560 vn_p.n111 vn_p.t47 756.008
R561 vn_p.n111 vn_p.t1307 756.008
R562 vn_p.n109 vn_p.t596 756.008
R563 vn_p.n109 vn_p.t352 756.008
R564 vn_p.n107 vn_p.t248 756.008
R565 vn_p.n107 vn_p.t7 756.008
R566 vn_p.n105 vn_p.t1434 756.008
R567 vn_p.n105 vn_p.t1191 756.008
R568 vn_p.n103 vn_p.t1083 756.008
R569 vn_p.n103 vn_p.t853 756.008
R570 vn_p.n101 vn_p.t744 756.008
R571 vn_p.n101 vn_p.t499 756.008
R572 vn_p.n99 vn_p.t1289 756.008
R573 vn_p.n99 vn_p.t1051 756.008
R574 vn_p.n97 vn_p.t944 756.008
R575 vn_p.n97 vn_p.t704 756.008
R576 vn_p.n95 vn_p.t1273 756.008
R577 vn_p.n95 vn_p.t1041 756.008
R578 vn_p.n93 vn_p.t928 756.008
R579 vn_p.n93 vn_p.t697 756.008
R580 vn_p.n91 vn_p.t585 756.008
R581 vn_p.n91 vn_p.t341 756.008
R582 vn_p.n89 vn_p.t1128 756.008
R583 vn_p.n89 vn_p.t892 756.008
R584 vn_p.n87 vn_p.t791 756.008
R585 vn_p.n87 vn_p.t542 756.008
R586 vn_p.n85 vn_p.t478 756.008
R587 vn_p.n85 vn_p.t240 756.008
R588 vn_p.n83 vn_p.t132 756.008
R589 vn_p.n83 vn_p.t1395 756.008
R590 vn_p.n81 vn_p.t673 756.008
R591 vn_p.n81 vn_p.t441 756.008
R592 vn_p.n79 vn_p.t323 756.008
R593 vn_p.n79 vn_p.t93 756.008
R594 vn_p.n77 vn_p.t1475 756.008
R595 vn_p.n77 vn_p.t1237 756.008
R596 vn_p.n75 vn_p.t1167 756.008
R597 vn_p.n75 vn_p.t933 756.008
R598 vn_p.n74 vn_p.t828 756.008
R599 vn_p.n74 vn_p.t586 756.008
R600 vn_p.n970 vn_p.t712 756.008
R601 vn_p.n970 vn_p.t1269 756.008
R602 vn_p.n968 vn_p.t361 756.008
R603 vn_p.n968 vn_p.t923 756.008
R604 vn_p.n966 vn_p.t908 756.008
R605 vn_p.n966 vn_p.t1465 756.008
R606 vn_p.n964 vn_p.t564 756.008
R607 vn_p.n964 vn_p.t1123 756.008
R608 vn_p.n962 vn_p.t251 756.008
R609 vn_p.n962 vn_p.t820 756.008
R610 vn_p.n960 vn_p.t1412 756.008
R611 vn_p.n960 vn_p.t474 756.008
R612 vn_p.n958 vn_p.t1058 756.008
R613 vn_p.n958 vn_p.t127 756.008
R614 vn_p.n956 vn_p.t112 756.008
R615 vn_p.n956 vn_p.t668 756.008
R616 vn_p.n954 vn_p.t1261 756.008
R617 vn_p.n954 vn_p.t319 756.008
R618 vn_p.n952 vn_p.t950 756.008
R619 vn_p.n952 vn_p.t13 756.008
R620 vn_p.n950 vn_p.t606 756.008
R621 vn_p.n950 vn_p.t1163 756.008
R622 vn_p.n948 vn_p.t1148 756.008
R623 vn_p.n948 vn_p.t218 756.008
R624 vn_p.n946 vn_p.t808 756.008
R625 vn_p.n946 vn_p.t1374 756.008
R626 vn_p.n944 vn_p.t466 756.008
R627 vn_p.n944 vn_p.t1024 756.008
R628 vn_p.n942 vn_p.t150 756.008
R629 vn_p.n942 vn_p.t711 756.008
R630 vn_p.n940 vn_p.t1299 756.008
R631 vn_p.n940 vn_p.t360 756.008
R632 vn_p.n938 vn_p.t1389 756.008
R633 vn_p.n938 vn_p.t451 756.008
R634 vn_p.n936 vn_p.t1037 756.008
R635 vn_p.n936 vn_p.t104 756.008
R636 vn_p.n934 vn_p.t693 756.008
R637 vn_p.n934 vn_p.t1248 756.008
R638 vn_p.n932 vn_p.t371 756.008
R639 vn_p.n932 vn_p.t942 756.008
R640 vn_p.n930 vn_p.t30 756.008
R641 vn_p.n930 vn_p.t598 756.008
R642 vn_p.n928 vn_p.t578 756.008
R643 vn_p.n928 vn_p.t1142 756.008
R644 vn_p.n926 vn_p.t234 756.008
R645 vn_p.n926 vn_p.t803 756.008
R646 vn_p.n924 vn_p.t782 756.008
R647 vn_p.n924 vn_p.t1343 756.008
R648 vn_p.n922 vn_p.t1067 756.008
R649 vn_p.n922 vn_p.t143 756.008
R650 vn_p.n920 vn_p.t729 756.008
R651 vn_p.n920 vn_p.t1291 756.008
R652 vn_p.n918 vn_p.t1270 756.008
R653 vn_p.n918 vn_p.t335 756.008
R654 vn_p.n916 vn_p.t926 756.008
R655 vn_p.n916 vn_p.t1489 756.008
R656 vn_p.n914 vn_p.t1468 756.008
R657 vn_p.n914 vn_p.t535 756.008
R658 vn_p.n912 vn_p.t264 756.008
R659 vn_p.n912 vn_p.t837 756.008
R660 vn_p.n910 vn_p.t822 756.008
R661 vn_p.n910 vn_p.t1387 756.008
R662 vn_p.n908 vn_p.t476 756.008
R663 vn_p.n908 vn_p.t1036 756.008
R664 vn_p.n906 vn_p.t130 756.008
R665 vn_p.n906 vn_p.t692 756.008
R666 vn_p.n904 vn_p.t670 756.008
R667 vn_p.n904 vn_p.t1229 756.008
R668 vn_p.n902 vn_p.t968 756.008
R669 vn_p.n902 vn_p.t28 756.008
R670 vn_p.n900 vn_p.t15 756.008
R671 vn_p.n900 vn_p.t577 756.008
R672 vn_p.n898 vn_p.t1164 756.008
R673 vn_p.n898 vn_p.t233 756.008
R674 vn_p.n896 vn_p.t826 756.008
R675 vn_p.n896 vn_p.t1393 756.008
R676 vn_p.n894 vn_p.t1376 756.008
R677 vn_p.n894 vn_p.t436 756.008
R678 vn_p.n892 vn_p.t168 756.008
R679 vn_p.n892 vn_p.t727 756.008
R680 vn_p.n890 vn_p.t1362 756.008
R681 vn_p.n890 vn_p.t423 756.008
R682 vn_p.n888 vn_p.t1013 756.008
R683 vn_p.n888 vn_p.t76 756.008
R684 vn_p.n886 vn_p.t57 756.008
R685 vn_p.n886 vn_p.t619 756.008
R686 vn_p.n884 vn_p.t1200 756.008
R687 vn_p.n884 vn_p.t269 756.008
R688 vn_p.n882 vn_p.t1 756.008
R689 vn_p.n882 vn_p.t570 756.008
R690 vn_p.n880 vn_p.t547 756.008
R691 vn_p.n880 vn_p.t1112 756.008
R692 vn_p.n878 vn_p.t210 756.008
R693 vn_p.n878 vn_p.t773 756.008
R694 vn_p.n876 vn_p.t754 756.008
R695 vn_p.n876 vn_p.t1318 756.008
R696 vn_p.n874 vn_p.t405 756.008
R697 vn_p.n874 vn_p.t972 756.008
R698 vn_p.n872 vn_p.t100 756.008
R699 vn_p.n872 vn_p.t653 756.008
R700 vn_p.n870 vn_p.t1243 756.008
R701 vn_p.n870 vn_p.t304 756.008
R702 vn_p.n868 vn_p.t901 756.008
R703 vn_p.n868 vn_p.t1460 756.008
R704 vn_p.n866 vn_p.t1444 756.008
R705 vn_p.n866 vn_p.t508 756.008
R706 vn_p.n864 vn_p.t1096 756.008
R707 vn_p.n864 vn_p.t175 756.008
R708 vn_p.n862 vn_p.t798 756.008
R709 vn_p.n862 vn_p.t1360 756.008
R710 vn_p.n860 vn_p.t452 756.008
R711 vn_p.n860 vn_p.t1012 756.008
R712 vn_p.n858 vn_p.t105 756.008
R713 vn_p.n858 vn_p.t660 756.008
R714 vn_p.n856 vn_p.t641 756.008
R715 vn_p.n856 vn_p.t1199 756.008
R716 vn_p.n854 vn_p.t295 756.008
R717 vn_p.n854 vn_p.t867 756.008
R718 vn_p.n852 vn_p.t1484 756.008
R719 vn_p.n852 vn_p.t546 756.008
R720 vn_p.n850 vn_p.t1143 756.008
R721 vn_p.n850 vn_p.t209 756.008
R722 vn_p.n848 vn_p.t194 756.008
R723 vn_p.n848 vn_p.t752 756.008
R724 vn_p.n846 vn_p.t1344 756.008
R725 vn_p.n846 vn_p.t403 756.008
R726 vn_p.n844 vn_p.t1001 756.008
R727 vn_p.n844 vn_p.t63 756.008
R728 vn_p.n842 vn_p.t1328 756.008
R729 vn_p.n842 vn_p.t390 756.008
R730 vn_p.n840 vn_p.t987 756.008
R731 vn_p.n840 vn_p.t48 756.008
R732 vn_p.n838 vn_p.t29 756.008
R733 vn_p.n838 vn_p.t597 756.008
R734 vn_p.n836 vn_p.t1176 756.008
R735 vn_p.n836 vn_p.t249 756.008
R736 vn_p.n834 vn_p.t842 756.008
R737 vn_p.n834 vn_p.t1404 756.008
R738 vn_p.n832 vn_p.t518 756.008
R739 vn_p.n832 vn_p.t1084 756.008
R740 vn_p.n830 vn_p.t185 756.008
R741 vn_p.n830 vn_p.t746 756.008
R742 vn_p.n828 vn_p.t728 756.008
R743 vn_p.n828 vn_p.t1290 756.008
R744 vn_p.n826 vn_p.t377 756.008
R745 vn_p.n826 vn_p.t945 756.008
R746 vn_p.n824 vn_p.t924 756.008
R747 vn_p.n824 vn_p.t1487 756.008
R748 vn_p.n823 vn_p.t1215 756.008
R749 vn_p.n823 vn_p.t280 756.008
R750 vn_p.n1119 vn_p.t344 756.008
R751 vn_p.n1119 vn_p.t916 756.008
R752 vn_p.n1117 vn_p.t895 756.008
R753 vn_p.n1117 vn_p.t1459 756.008
R754 vn_p.n1115 vn_p.t545 756.008
R755 vn_p.n1115 vn_p.t1114 756.008
R756 vn_p.n1113 vn_p.t847 756.008
R757 vn_p.n1113 vn_p.t1416 756.008
R758 vn_p.n1111 vn_p.t1398 756.008
R759 vn_p.n1111 vn_p.t469 756.008
R760 vn_p.n1109 vn_p.t1046 756.008
R761 vn_p.n1109 vn_p.t119 756.008
R762 vn_p.n1107 vn_p.t97 756.008
R763 vn_p.n1107 vn_p.t657 756.008
R764 vn_p.n1105 vn_p.t1241 756.008
R765 vn_p.n1105 vn_p.t307 756.008
R766 vn_p.n1103 vn_p.t936 756.008
R767 vn_p.n1103 vn_p.t1499 756.008
R768 vn_p.n1101 vn_p.t591 756.008
R769 vn_p.n1101 vn_p.t1156 756.008
R770 vn_p.n1099 vn_p.t245 756.008
R771 vn_p.n1099 vn_p.t814 756.008
R772 vn_p.n1097 vn_p.t796 756.008
R773 vn_p.n1097 vn_p.t1365 756.008
R774 vn_p.n1095 vn_p.t450 756.008
R775 vn_p.n1095 vn_p.t1014 756.008
R776 vn_p.n1093 vn_p.t139 756.008
R777 vn_p.n1093 vn_p.t701 756.008
R778 vn_p.n1091 vn_p.t1284 756.008
R779 vn_p.n1091 vn_p.t349 756.008
R780 vn_p.n1089 vn_p.t941 756.008
R781 vn_p.n1089 vn_p.t5 756.008
R782 vn_p.n1087 vn_p.t1026 756.008
R783 vn_p.n1087 vn_p.t94 756.008
R784 vn_p.n1085 vn_p.t675 756.008
R785 vn_p.n1085 vn_p.t1238 756.008
R786 vn_p.n1083 vn_p.t362 756.008
R787 vn_p.n1083 vn_p.t932 756.008
R788 vn_p.n1081 vn_p.t18 756.008
R789 vn_p.n1081 vn_p.t588 756.008
R790 vn_p.n1079 vn_p.t565 756.008
R791 vn_p.n1079 vn_p.t1130 756.008
R792 vn_p.n1077 vn_p.t224 756.008
R793 vn_p.n1077 vn_p.t792 756.008
R794 vn_p.n1075 vn_p.t1380 756.008
R795 vn_p.n1075 vn_p.t445 756.008
R796 vn_p.n1073 vn_p.t1059 756.008
R797 vn_p.n1073 vn_p.t134 756.008
R798 vn_p.n1071 vn_p.t717 756.008
R799 vn_p.n1071 vn_p.t1280 756.008
R800 vn_p.n1069 vn_p.t1262 756.008
R801 vn_p.n1069 vn_p.t325 756.008
R802 vn_p.n1067 vn_p.t914 756.008
R803 vn_p.n1067 vn_p.t1476 756.008
R804 vn_p.n1065 vn_p.t571 756.008
R805 vn_p.n1065 vn_p.t1136 756.008
R806 vn_p.n1063 vn_p.t255 756.008
R807 vn_p.n1063 vn_p.t831 756.008
R808 vn_p.n1061 vn_p.t1414 756.008
R809 vn_p.n1061 vn_p.t483 756.008
R810 vn_p.n1059 vn_p.t465 756.008
R811 vn_p.n1059 vn_p.t1029 756.008
R812 vn_p.n1057 vn_p.t116 756.008
R813 vn_p.n1057 vn_p.t678 756.008
R814 vn_p.n1055 vn_p.t654 756.008
R815 vn_p.n1055 vn_p.t1219 756.008
R816 vn_p.n1053 vn_p.t952 756.008
R817 vn_p.n1053 vn_p.t22 756.008
R818 vn_p.n1051 vn_p.t607 756.008
R819 vn_p.n1051 vn_p.t1170 756.008
R820 vn_p.n1049 vn_p.t1150 756.008
R821 vn_p.n1049 vn_p.t226 756.008
R822 vn_p.n1047 vn_p.t811 756.008
R823 vn_p.n1047 vn_p.t1382 756.008
R824 vn_p.n1045 vn_p.t1361 756.008
R825 vn_p.n1045 vn_p.t427 756.008
R826 vn_p.n1043 vn_p.t152 756.008
R827 vn_p.n1043 vn_p.t721 756.008
R828 vn_p.n1041 vn_p.t1342 756.008
R829 vn_p.n1041 vn_p.t409 756.008
R830 vn_p.n1039 vn_p.t1000 756.008
R831 vn_p.n1039 vn_p.t67 756.008
R832 vn_p.n1037 vn_p.t647 756.008
R833 vn_p.n1037 vn_p.t1209 756.008
R834 vn_p.n1035 vn_p.t1190 756.008
R835 vn_p.n1035 vn_p.t262 756.008
R836 vn_p.n1033 vn_p.t1488 756.008
R837 vn_p.n1033 vn_p.t558 756.008
R838 vn_p.n1031 vn_p.t536 756.008
R839 vn_p.n1031 vn_p.t1103 756.008
R840 vn_p.n1029 vn_p.t199 756.008
R841 vn_p.n1029 vn_p.t762 756.008
R842 vn_p.n1027 vn_p.t1351 756.008
R843 vn_p.n1027 vn_p.t417 756.008
R844 vn_p.n1025 vn_p.t391 756.008
R845 vn_p.n1025 vn_p.t962 756.008
R846 vn_p.n1023 vn_p.t691 756.008
R847 vn_p.n1023 vn_p.t1253 756.008
R848 vn_p.n1021 vn_p.t1228 756.008
R849 vn_p.n1021 vn_p.t296 756.008
R850 vn_p.n1019 vn_p.t888 756.008
R851 vn_p.n1019 vn_p.t1452 756.008
R852 vn_p.n1017 vn_p.t1435 756.008
R853 vn_p.n1017 vn_p.t500 756.008
R854 vn_p.n1015 vn_p.t1085 756.008
R855 vn_p.n1015 vn_p.t162 756.008
R856 vn_p.n1013 vn_p.t1392 756.008
R857 vn_p.n1013 vn_p.t460 756.008
R858 vn_p.n1011 vn_p.t435 756.008
R859 vn_p.n1011 vn_p.t1003 756.008
R860 vn_p.n1009 vn_p.t89 756.008
R861 vn_p.n1009 vn_p.t649 756.008
R862 vn_p.n1007 vn_p.t629 756.008
R863 vn_p.n1007 vn_p.t1192 756.008
R864 vn_p.n1005 vn_p.t281 756.008
R865 vn_p.n1005 vn_p.t856 756.008
R866 vn_p.n1003 vn_p.t1466 756.008
R867 vn_p.n1003 vn_p.t539 756.008
R868 vn_p.n1001 vn_p.t1124 756.008
R869 vn_p.n1001 vn_p.t202 756.008
R870 vn_p.n999 vn_p.t786 756.008
R871 vn_p.n999 vn_p.t1355 756.008
R872 vn_p.n997 vn_p.t1327 756.008
R873 vn_p.n997 vn_p.t394 756.008
R874 vn_p.n995 vn_p.t985 756.008
R875 vn_p.n995 vn_p.t52 756.008
R876 vn_p.n993 vn_p.t1317 756.008
R877 vn_p.n993 vn_p.t379 756.008
R878 vn_p.n991 vn_p.t973 756.008
R879 vn_p.n991 vn_p.t40 756.008
R880 vn_p.n989 vn_p.t622 756.008
R881 vn_p.n989 vn_p.t1184 756.008
R882 vn_p.n987 vn_p.t1169 756.008
R883 vn_p.n987 vn_p.t243 756.008
R884 vn_p.n985 vn_p.t830 756.008
R885 vn_p.n985 vn_p.t1399 756.008
R886 vn_p.n983 vn_p.t509 756.008
R887 vn_p.n983 vn_p.t1075 756.008
R888 vn_p.n981 vn_p.t174 756.008
R889 vn_p.n981 vn_p.t738 756.008
R890 vn_p.n979 vn_p.t716 756.008
R891 vn_p.n979 vn_p.t1279 756.008
R892 vn_p.n977 vn_p.t364 756.008
R893 vn_p.n977 vn_p.t937 756.008
R894 vn_p.n975 vn_p.t21 756.008
R895 vn_p.n975 vn_p.t592 756.008
R896 vn_p.n973 vn_p.t1198 756.008
R897 vn_p.n973 vn_p.t271 756.008
R898 vn_p.n972 vn_p.t866 756.008
R899 vn_p.n972 vn_p.t1429 756.008
R900 vn_p.n1268 vn_p.t336 756.008
R901 vn_p.n1268 vn_p.t470 756.008
R902 vn_p.n1266 vn_p.t1491 756.008
R903 vn_p.n1266 vn_p.t123 756.008
R904 vn_p.n1264 vn_p.t537 756.008
R905 vn_p.n1264 vn_p.t661 756.008
R906 vn_p.n1262 vn_p.t201 756.008
R907 vn_p.n1262 vn_p.t312 756.008
R908 vn_p.n1260 vn_p.t1391 756.008
R909 vn_p.n1260 vn_p.t0 756.008
R910 vn_p.n1258 vn_p.t1040 756.008
R911 vn_p.n1258 vn_p.t1158 756.008
R912 vn_p.n1256 vn_p.t694 756.008
R913 vn_p.n1256 vn_p.t817 756.008
R914 vn_p.n1254 vn_p.t1232 756.008
R915 vn_p.n1254 vn_p.t1367 756.008
R916 vn_p.n1252 vn_p.t891 756.008
R917 vn_p.n1252 vn_p.t1020 756.008
R918 vn_p.n1250 vn_p.t582 756.008
R919 vn_p.n1250 vn_p.t702 756.008
R920 vn_p.n1248 vn_p.t238 756.008
R921 vn_p.n1248 vn_p.t353 756.008
R922 vn_p.n1246 vn_p.t785 756.008
R923 vn_p.n1246 vn_p.t900 756.008
R924 vn_p.n1244 vn_p.t440 756.008
R925 vn_p.n1244 vn_p.t555 756.008
R926 vn_p.n1242 vn_p.t92 756.008
R927 vn_p.n1242 vn_p.t216 756.008
R928 vn_p.n1240 vn_p.t1276 756.008
R929 vn_p.n1240 vn_p.t1403 756.008
R930 vn_p.n1238 vn_p.t931 756.008
R931 vn_p.n1238 vn_p.t1052 756.008
R932 vn_p.n1236 vn_p.t1018 756.008
R933 vn_p.n1236 vn_p.t1133 756.008
R934 vn_p.n1234 vn_p.t665 756.008
R935 vn_p.n1234 vn_p.t793 756.008
R936 vn_p.n1232 vn_p.t316 756.008
R937 vn_p.n1232 vn_p.t446 756.008
R938 vn_p.n1230 vn_p.t8 756.008
R939 vn_p.n1230 vn_p.t136 756.008
R940 vn_p.n1228 vn_p.t1160 756.008
R941 vn_p.n1228 vn_p.t1282 756.008
R942 vn_p.n1226 vn_p.t215 756.008
R943 vn_p.n1226 vn_p.t326 756.008
R944 vn_p.n1224 vn_p.t1370 756.008
R945 vn_p.n1224 vn_p.t1477 756.008
R946 vn_p.n1222 vn_p.t410 756.008
R947 vn_p.n1222 vn_p.t525 756.008
R948 vn_p.n1220 vn_p.t705 756.008
R949 vn_p.n1220 vn_p.t832 756.008
R950 vn_p.n1218 vn_p.t355 756.008
R951 vn_p.n1218 vn_p.t485 756.008
R952 vn_p.n1216 vn_p.t904 756.008
R953 vn_p.n1216 vn_p.t1030 756.008
R954 vn_p.n1214 vn_p.t559 756.008
R955 vn_p.n1214 vn_p.t681 756.008
R956 vn_p.n1212 vn_p.t1100 756.008
R957 vn_p.n1212 vn_p.t1221 756.008
R958 vn_p.n1210 vn_p.t1405 756.008
R959 vn_p.n1210 vn_p.t24 756.008
R960 vn_p.n1208 vn_p.t456 756.008
R961 vn_p.n1208 vn_p.t572 756.008
R962 vn_p.n1206 vn_p.t107 756.008
R963 vn_p.n1206 vn_p.t227 756.008
R964 vn_p.n1204 vn_p.t1254 756.008
R965 vn_p.n1204 vn_p.t1385 756.008
R966 vn_p.n1202 vn_p.t297 756.008
R967 vn_p.n1202 vn_p.t429 756.008
R968 vn_p.n1200 vn_p.t600 756.008
R969 vn_p.n1200 vn_p.t723 756.008
R970 vn_p.n1198 vn_p.t1144 756.008
R971 vn_p.n1198 vn_p.t1265 756.008
R972 vn_p.n1196 vn_p.t804 756.008
R973 vn_p.n1196 vn_p.t919 756.008
R974 vn_p.n1194 vn_p.t461 756.008
R975 vn_p.n1194 vn_p.t576 756.008
R976 vn_p.n1192 vn_p.t1004 756.008
R977 vn_p.n1192 vn_p.t1117 756.008
R978 vn_p.n1190 vn_p.t1295 756.008
R979 vn_p.n1190 vn_p.t1420 756.008
R980 vn_p.n1188 vn_p.t991 756.008
R981 vn_p.n1188 vn_p.t1104 756.008
R982 vn_p.n1186 vn_p.t637 756.008
R983 vn_p.n1186 vn_p.t763 756.008
R984 vn_p.n1184 vn_p.t1181 756.008
R985 vn_p.n1184 vn_p.t1308 756.008
R986 vn_p.n1182 vn_p.t845 756.008
R987 vn_p.n1182 vn_p.t963 756.008
R988 vn_p.n1180 vn_p.t1135 756.008
R989 vn_p.n1180 vn_p.t1257 756.008
R990 vn_p.n1178 vn_p.t188 756.008
R991 vn_p.n1178 vn_p.t298 756.008
R992 vn_p.n1176 vn_p.t1338 756.008
R993 vn_p.n1176 vn_p.t1454 756.008
R994 vn_p.n1174 vn_p.t380 756.008
R995 vn_p.n1174 vn_p.t501 756.008
R996 vn_p.n1172 vn_p.t39 756.008
R997 vn_p.n1172 vn_p.t164 756.008
R998 vn_p.n1170 vn_p.t1218 756.008
R999 vn_p.n1170 vn_p.t1352 756.008
R1000 vn_p.n1168 vn_p.t878 756.008
R1001 vn_p.n1168 vn_p.t1005 756.008
R1002 vn_p.n1166 vn_p.t528 756.008
R1003 vn_p.n1166 vn_p.t651 756.008
R1004 vn_p.n1164 vn_p.t1074 756.008
R1005 vn_p.n1164 vn_p.t1194 756.008
R1006 vn_p.n1162 vn_p.t739 756.008
R1007 vn_p.n1162 vn_p.t859 756.008
R1008 vn_p.n1160 vn_p.t426 756.008
R1009 vn_p.n1160 vn_p.t541 756.008
R1010 vn_p.n1158 vn_p.t78 756.008
R1011 vn_p.n1158 vn_p.t203 756.008
R1012 vn_p.n1156 vn_p.t1224 756.008
R1013 vn_p.n1156 vn_p.t1357 756.008
R1014 vn_p.n1154 vn_p.t272 756.008
R1015 vn_p.n1154 vn_p.t397 756.008
R1016 vn_p.n1152 vn_p.t1430 756.008
R1017 vn_p.n1152 vn_p.t54 756.008
R1018 vn_p.n1150 vn_p.t1115 756.008
R1019 vn_p.n1150 vn_p.t1236 756.008
R1020 vn_p.n1148 vn_p.t775 756.008
R1021 vn_p.n1148 vn_p.t893 756.008
R1022 vn_p.n1146 vn_p.t1321 756.008
R1023 vn_p.n1146 vn_p.t1440 756.008
R1024 vn_p.n1144 vn_p.t976 756.008
R1025 vn_p.n1144 vn_p.t1089 756.008
R1026 vn_p.n1142 vn_p.t627 756.008
R1027 vn_p.n1142 vn_p.t750 756.008
R1028 vn_p.n1140 vn_p.t961 756.008
R1029 vn_p.n1140 vn_p.t1076 756.008
R1030 vn_p.n1138 vn_p.t615 756.008
R1031 vn_p.n1138 vn_p.t740 756.008
R1032 vn_p.n1136 vn_p.t1159 756.008
R1033 vn_p.n1136 vn_p.t1281 756.008
R1034 vn_p.n1134 vn_p.t821 756.008
R1035 vn_p.n1134 vn_p.t938 756.008
R1036 vn_p.n1132 vn_p.t475 756.008
R1037 vn_p.n1132 vn_p.t593 756.008
R1038 vn_p.n1130 vn_p.t161 756.008
R1039 vn_p.n1130 vn_p.t273 756.008
R1040 vn_p.n1128 vn_p.t1311 756.008
R1041 vn_p.n1128 vn_p.t1432 756.008
R1042 vn_p.n1126 vn_p.t354 756.008
R1043 vn_p.n1126 vn_p.t484 756.008
R1044 vn_p.n1124 vn_p.t12 756.008
R1045 vn_p.n1124 vn_p.t140 756.008
R1046 vn_p.n1122 vn_p.t557 756.008
R1047 vn_p.n1122 vn_p.t679 756.008
R1048 vn_p.n1121 vn_p.t855 756.008
R1049 vn_p.n1121 vn_p.t978 756.008
R1050 vn_p.n1417 vn_p.t1043 756.008
R1051 vn_p.n1417 vn_p.t1322 756.008
R1052 vn_p.n1415 vn_p.t90 756.008
R1053 vn_p.n1415 vn_p.t365 756.008
R1054 vn_p.n1413 vn_p.t1234 756.008
R1055 vn_p.n1413 vn_p.t23 756.008
R1056 vn_p.n1411 vn_p.t37 756.008
R1057 vn_p.n1411 vn_p.t314 756.008
R1058 vn_p.n1409 vn_p.t583 756.008
R1059 vn_p.n1409 vn_p.t869 756.008
R1060 vn_p.n1407 vn_p.t241 756.008
R1061 vn_p.n1407 vn_p.t513 756.008
R1062 vn_p.n1405 vn_p.t788 756.008
R1063 vn_p.n1405 vn_p.t1062 756.008
R1064 vn_p.n1403 vn_p.t443 756.008
R1065 vn_p.n1403 vn_p.t722 756.008
R1066 vn_p.n1401 vn_p.t128 756.008
R1067 vn_p.n1401 vn_p.t407 756.008
R1068 vn_p.n1399 vn_p.t1277 756.008
R1069 vn_p.n1399 vn_p.t66 756.008
R1070 vn_p.n1397 vn_p.t935 756.008
R1071 vn_p.n1397 vn_p.t1207 756.008
R1072 vn_p.n1395 vn_p.t1473 756.008
R1073 vn_p.n1395 vn_p.t261 756.008
R1074 vn_p.n1393 vn_p.t1132 756.008
R1075 vn_p.n1393 vn_p.t1419 756.008
R1076 vn_p.n1391 vn_p.t825 756.008
R1077 vn_p.n1391 vn_p.t1098 756.008
R1078 vn_p.n1389 vn_p.t482 756.008
R1079 vn_p.n1389 vn_p.t760 756.008
R1080 vn_p.n1387 vn_p.t135 756.008
R1081 vn_p.n1387 vn_p.t413 756.008
R1082 vn_p.n1385 vn_p.t217 756.008
R1083 vn_p.n1385 vn_p.t494 756.008
R1084 vn_p.n1383 vn_p.t1371 756.008
R1085 vn_p.n1383 vn_p.t151 756.008
R1086 vn_p.n1381 vn_p.t1053 756.008
R1087 vn_p.n1381 vn_p.t1336 756.008
R1088 vn_p.n1379 vn_p.t706 756.008
R1089 vn_p.n1379 vn_p.t992 756.008
R1090 vn_p.n1377 vn_p.t1250 756.008
R1091 vn_p.n1377 vn_p.t38 756.008
R1092 vn_p.n1375 vn_p.t905 756.008
R1093 vn_p.n1375 vn_p.t1183 756.008
R1094 vn_p.n1373 vn_p.t560 756.008
R1095 vn_p.n1373 vn_p.t846 756.008
R1096 vn_p.n1371 vn_p.t250 756.008
R1097 vn_p.n1371 vn_p.t526 756.008
R1098 vn_p.n1369 vn_p.t1407 756.008
R1099 vn_p.n1369 vn_p.t192 756.008
R1100 vn_p.n1367 vn_p.t458 756.008
R1101 vn_p.n1367 vn_p.t735 756.008
R1102 vn_p.n1365 vn_p.t108 756.008
R1103 vn_p.n1365 vn_p.t384 756.008
R1104 vn_p.n1363 vn_p.t1255 756.008
R1105 vn_p.n1363 vn_p.t42 756.008
R1106 vn_p.n1361 vn_p.t947 756.008
R1107 vn_p.n1361 vn_p.t1223 756.008
R1108 vn_p.n1359 vn_p.t602 756.008
R1109 vn_p.n1359 vn_p.t882 756.008
R1110 vn_p.n1357 vn_p.t1145 756.008
R1111 vn_p.n1357 vn_p.t1428 756.008
R1112 vn_p.n1355 vn_p.t805 756.008
R1113 vn_p.n1355 vn_p.t1078 756.008
R1114 vn_p.n1353 vn_p.t1353 756.008
R1115 vn_p.n1353 vn_p.t138 756.008
R1116 vn_p.n1351 vn_p.t148 756.008
R1117 vn_p.n1351 vn_p.t431 756.008
R1118 vn_p.n1349 vn_p.t1297 756.008
R1119 vn_p.n1349 vn_p.t80 756.008
R1120 vn_p.n1347 vn_p.t339 756.008
R1121 vn_p.n1347 vn_p.t626 756.008
R1122 vn_p.n1345 vn_p.t1494 756.008
R1123 vn_p.n1345 vn_p.t275 756.008
R1124 vn_p.n1343 vn_p.t540 756.008
R1125 vn_p.n1343 vn_p.t834 756.008
R1126 vn_p.n1341 vn_p.t844 756.008
R1127 vn_p.n1341 vn_p.t1119 756.008
R1128 vn_p.n1339 vn_p.t524 756.008
R1129 vn_p.n1339 vn_p.t818 756.008
R1130 vn_p.n1337 vn_p.t189 756.008
R1131 vn_p.n1337 vn_p.t473 756.008
R1132 vn_p.n1335 vn_p.t1339 756.008
R1133 vn_p.n1335 vn_p.t126 756.008
R1134 vn_p.n1333 vn_p.t382 756.008
R1135 vn_p.n1333 vn_p.t667 756.008
R1136 vn_p.n1331 vn_p.t680 756.008
R1137 vn_p.n1331 vn_p.t964 756.008
R1138 vn_p.n1329 vn_p.t1220 756.008
R1139 vn_p.n1329 vn_p.t9 756.008
R1140 vn_p.n1327 vn_p.t879 756.008
R1141 vn_p.n1327 vn_p.t1161 756.008
R1142 vn_p.n1325 vn_p.t531 756.008
R1143 vn_p.n1325 vn_p.t824 756.008
R1144 vn_p.n1323 vn_p.t1077 756.008
R1145 vn_p.n1323 vn_p.t1372 756.008
R1146 vn_p.n1321 vn_p.t1384 756.008
R1147 vn_p.n1321 vn_p.t167 756.008
R1148 vn_p.n1319 vn_p.t428 756.008
R1149 vn_p.n1319 vn_p.t708 756.008
R1150 vn_p.n1317 vn_p.t79 756.008
R1151 vn_p.n1317 vn_p.t359 756.008
R1152 vn_p.n1315 vn_p.t623 756.008
R1153 vn_p.n1315 vn_p.t906 756.008
R1154 vn_p.n1313 vn_p.t274 756.008
R1155 vn_p.n1313 vn_p.t562 756.008
R1156 vn_p.n1311 vn_p.t575 756.008
R1157 vn_p.n1311 vn_p.t862 756.008
R1158 vn_p.n1309 vn_p.t1116 756.008
R1159 vn_p.n1309 vn_p.t1411 756.008
R1160 vn_p.n1307 vn_p.t777 756.008
R1161 vn_p.n1307 vn_p.t1056 756.008
R1162 vn_p.n1305 vn_p.t1323 756.008
R1163 vn_p.n1305 vn_p.t110 756.008
R1164 vn_p.n1303 vn_p.t977 756.008
R1165 vn_p.n1303 vn_p.t1258 756.008
R1166 vn_p.n1301 vn_p.t663 756.008
R1167 vn_p.n1301 vn_p.t949 756.008
R1168 vn_p.n1299 vn_p.t315 756.008
R1169 vn_p.n1299 vn_p.t604 756.008
R1170 vn_p.n1297 vn_p.t1464 756.008
R1171 vn_p.n1297 vn_p.t252 756.008
R1172 vn_p.n1295 vn_p.t514 756.008
R1173 vn_p.n1295 vn_p.t806 756.008
R1174 vn_p.n1293 vn_p.t178 756.008
R1175 vn_p.n1293 vn_p.t464 756.008
R1176 vn_p.n1291 vn_p.t502 756.008
R1177 vn_p.n1291 vn_p.t795 756.008
R1178 vn_p.n1289 vn_p.t163 756.008
R1179 vn_p.n1289 vn_p.t449 756.008
R1180 vn_p.n1287 vn_p.t1312 756.008
R1181 vn_p.n1287 vn_p.t102 756.008
R1182 vn_p.n1285 vn_p.t356 756.008
R1183 vn_p.n1285 vn_p.t638 756.008
R1184 vn_p.n1283 vn_p.t14 756.008
R1185 vn_p.n1283 vn_p.t290 756.008
R1186 vn_p.n1281 vn_p.t1193 756.008
R1187 vn_p.n1281 vn_p.t1479 756.008
R1188 vn_p.n1279 vn_p.t858 756.008
R1189 vn_p.n1279 vn_p.t1140 756.008
R1190 vn_p.n1277 vn_p.t1406 756.008
R1191 vn_p.n1277 vn_p.t190 756.008
R1192 vn_p.n1275 vn_p.t1054 756.008
R1193 vn_p.n1275 vn_p.t1340 756.008
R1194 vn_p.n1273 vn_p.t713 756.008
R1195 vn_p.n1273 vn_p.t998 756.008
R1196 vn_p.n1271 vn_p.t396 756.008
R1197 vn_p.n1271 vn_p.t683 756.008
R1198 vn_p.n1270 vn_p.t53 756.008
R1199 vn_p.n1270 vn_p.t334 756.008
R1200 vn_p.n670 vn_p.t1423 706.013
R1201 vn_p.n749 vn_p.t294 706.013
R1202 vn_p.n1419 vn_p.t1259 706.013
R1203 vn_p.n0 vn_p.t6 705.989
R1204 vn_p.n743 vn_p.t909 704.872
R1205 vn_p.n742 vn_p.t1453 704.872
R1206 vn_p.n741 vn_p.t1107 704.872
R1207 vn_p.n740 vn_p.t1413 704.872
R1208 vn_p.n739 vn_p.t462 704.872
R1209 vn_p.n738 vn_p.t113 704.872
R1210 vn_p.n737 vn_p.t650 704.872
R1211 vn_p.n736 vn_p.t301 704.872
R1212 vn_p.n735 vn_p.t1493 704.872
R1213 vn_p.n734 vn_p.t1149 704.872
R1214 vn_p.n733 vn_p.t809 704.872
R1215 vn_p.n732 vn_p.t1356 704.872
R1216 vn_p.n731 vn_p.t1008 704.872
R1217 vn_p.n730 vn_p.t698 704.872
R1218 vn_p.n729 vn_p.t343 704.872
R1219 vn_p.n728 vn_p.t1496 704.872
R1220 vn_p.n727 vn_p.t84 704.872
R1221 vn_p.n726 vn_p.t1230 704.872
R1222 vn_p.n725 vn_p.t922 704.872
R1223 vn_p.n724 vn_p.t579 704.872
R1224 vn_p.n723 vn_p.t1121 704.872
R1225 vn_p.n722 vn_p.t783 704.872
R1226 vn_p.n721 vn_p.t438 704.872
R1227 vn_p.n720 vn_p.t125 704.872
R1228 vn_p.n719 vn_p.t1271 704.872
R1229 vn_p.n718 vn_p.t317 704.872
R1230 vn_p.n717 vn_p.t1469 704.872
R1231 vn_p.n716 vn_p.t1126 704.872
R1232 vn_p.n715 vn_p.t823 704.872
R1233 vn_p.n714 vn_p.t477 704.872
R1234 vn_p.n713 vn_p.t1022 704.872
R1235 vn_p.n712 vn_p.t672 704.872
R1236 vn_p.n711 vn_p.t1210 704.872
R1237 vn_p.n710 vn_p.t16 704.872
R1238 vn_p.n709 vn_p.t1166 704.872
R1239 vn_p.n708 vn_p.t220 704.872
R1240 vn_p.n707 vn_p.t1378 704.872
R1241 vn_p.n706 vn_p.t419 704.872
R1242 vn_p.n705 vn_p.t714 704.872
R1243 vn_p.n704 vn_p.t401 704.872
R1244 vn_p.n703 vn_p.t58 704.872
R1245 vn_p.n702 vn_p.t1201 704.872
R1246 vn_p.n701 vn_p.t256 704.872
R1247 vn_p.n700 vn_p.t549 704.872
R1248 vn_p.n699 vn_p.t1092 704.872
R1249 vn_p.n698 vn_p.t755 704.872
R1250 vn_p.n697 vn_p.t406 704.872
R1251 vn_p.n696 vn_p.t954 704.872
R1252 vn_p.n695 vn_p.t1245 704.872
R1253 vn_p.n694 vn_p.t289 704.872
R1254 vn_p.n693 vn_p.t1445 704.872
R1255 vn_p.n692 vn_p.t496 704.872
R1256 vn_p.n691 vn_p.t155 704.872
R1257 vn_p.n690 vn_p.t455 704.872
R1258 vn_p.n689 vn_p.t996 704.872
R1259 vn_p.n688 vn_p.t643 704.872
R1260 vn_p.n687 vn_p.t1186 704.872
R1261 vn_p.n686 vn_p.t849 704.872
R1262 vn_p.n685 vn_p.t532 704.872
R1263 vn_p.n684 vn_p.t196 704.872
R1264 vn_p.n683 vn_p.t1346 704.872
R1265 vn_p.n682 vn_p.t386 704.872
R1266 vn_p.n681 vn_p.t45 704.872
R1267 vn_p.n680 vn_p.t373 704.872
R1268 vn_p.n679 vn_p.t32 704.872
R1269 vn_p.n678 vn_p.t1177 704.872
R1270 vn_p.n677 vn_p.t235 704.872
R1271 vn_p.n676 vn_p.t1394 704.872
R1272 vn_p.n675 vn_p.t1069 704.872
R1273 vn_p.n674 vn_p.t731 704.872
R1274 vn_p.n673 vn_p.t1272 704.872
R1275 vn_p.n672 vn_p.t927 704.872
R1276 vn_p.n671 vn_p.t584 704.872
R1277 vn_p.n670 vn_p.t266 704.872
R1278 vn_p.n0 vn_p.t1204 704.872
R1279 vn_p.n1 vn_p.t664 704.872
R1280 vn_p.n2 vn_p.t1017 704.872
R1281 vn_p.n3 vn_p.t472 704.872
R1282 vn_p.n4 vn_p.t815 704.872
R1283 vn_p.n5 vn_p.t1120 704.872
R1284 vn_p.n6 vn_p.t1461 704.872
R1285 vn_p.n7 vn_p.t310 704.872
R1286 vn_p.n8 vn_p.t1267 704.872
R1287 vn_p.n9 vn_p.t121 704.872
R1288 vn_p.n10 vn_p.t1278 704.872
R1289 vn_p.n11 vn_p.t133 704.872
R1290 vn_p.n12 vn_p.t481 704.872
R1291 vn_p.n13 vn_p.t1425 704.872
R1292 vn_p.n14 vn_p.t270 704.872
R1293 vn_p.n15 vn_p.t587 704.872
R1294 vn_p.n16 vn_p.t934 704.872
R1295 vn_p.n17 vn_p.t381 704.872
R1296 vn_p.n18 vn_p.t734 704.872
R1297 vn_p.n19 vn_p.t1072 704.872
R1298 vn_p.n20 vn_p.t1396 704.872
R1299 vn_p.n21 vn_p.t239 704.872
R1300 vn_p.n22 vn_p.t1182 704.872
R1301 vn_p.n23 vn_p.t35 704.872
R1302 vn_p.n24 vn_p.t375 704.872
R1303 vn_p.n25 vn_p.t695 704.872
R1304 vn_p.n26 vn_p.t1042 704.872
R1305 vn_p.n27 vn_p.t491 704.872
R1306 vn_p.n28 vn_p.t841 704.872
R1307 vn_p.n29 vn_p.t285 704.872
R1308 vn_p.n30 vn_p.t1492 704.872
R1309 vn_p.n31 vn_p.t338 704.872
R1310 vn_p.n32 vn_p.t1294 704.872
R1311 vn_p.n33 vn_p.t146 704.872
R1312 vn_p.n34 vn_p.t457 704.872
R1313 vn_p.n35 vn_p.t160 704.872
R1314 vn_p.n36 vn_p.t1102 704.872
R1315 vn_p.n37 vn_p.t1450 704.872
R1316 vn_p.n38 vn_p.t292 704.872
R1317 vn_p.n39 vn_p.t1249 704.872
R1318 vn_p.n40 vn_p.t959 704.872
R1319 vn_p.n41 vn_p.t412 704.872
R1320 vn_p.n42 vn_p.t759 704.872
R1321 vn_p.n43 vn_p.t1094 704.872
R1322 vn_p.n44 vn_p.t554 704.872
R1323 vn_p.n45 vn_p.t258 704.872
R1324 vn_p.n46 vn_p.t1206 704.872
R1325 vn_p.n47 vn_p.t62 704.872
R1326 vn_p.n48 vn_p.t1019 704.872
R1327 vn_p.n49 vn_p.t1366 704.872
R1328 vn_p.n50 vn_p.t1061 704.872
R1329 vn_p.n51 vn_p.t511 704.872
R1330 vn_p.n52 vn_p.t865 704.872
R1331 vn_p.n53 vn_p.t311 704.872
R1332 vn_p.n54 vn_p.t659 704.872
R1333 vn_p.n55 vn_p.t975 704.872
R1334 vn_p.n56 vn_p.t1320 704.872
R1335 vn_p.n57 vn_p.t173 704.872
R1336 vn_p.n58 vn_p.t87 704.872
R1337 vn_p.n59 vn_p.t434 704.872
R1338 vn_p.n60 vn_p.t742 704.872
R1339 vn_p.n61 vn_p.t1082 704.872
R1340 vn_p.n62 vn_p.t1433 704.872
R1341 vn_p.n63 vn_p.t887 704.872
R1342 vn_p.n64 vn_p.t1227 704.872
R1343 vn_p.n65 vn_p.t46 704.872
R1344 vn_p.n66 vn_p.t387 704.872
R1345 vn_p.n67 vn_p.t1348 704.872
R1346 vn_p.n68 vn_p.t197 704.872
R1347 vn_p.n69 vn_p.t533 704.872
R1348 vn_p.n70 vn_p.t851 704.872
R1349 vn_p.n71 vn_p.t1187 704.872
R1350 vn_p.n72 vn_p.t644 704.872
R1351 vn_p.n73 vn_p.t997 704.872
R1352 vn_p.n749 vn_p.t640 704.872
R1353 vn_p.n750 vn_p.t960 704.872
R1354 vn_p.n751 vn_p.t1303 704.872
R1355 vn_p.n752 vn_p.t153 704.872
R1356 vn_p.n753 vn_p.t1095 704.872
R1357 vn_p.n754 vn_p.t1443 704.872
R1358 vn_p.n755 vn_p.t260 704.872
R1359 vn_p.n756 vn_p.t608 704.872
R1360 vn_p.n757 vn_p.t64 704.872
R1361 vn_p.n758 vn_p.t404 704.872
R1362 vn_p.n759 vn_p.t753 704.872
R1363 vn_p.n760 vn_p.t424 704.872
R1364 vn_p.n761 vn_p.t768 704.872
R1365 vn_p.n762 vn_p.t225 704.872
R1366 vn_p.n763 vn_p.t567 704.872
R1367 vn_p.n764 vn_p.t910 704.872
R1368 vn_p.n765 vn_p.t1216 704.872
R1369 vn_p.n766 vn_p.t71 704.872
R1370 vn_p.n767 vn_p.t1027 704.872
R1371 vn_p.n768 vn_p.t1375 704.872
R1372 vn_p.n769 vn_p.t827 704.872
R1373 vn_p.n770 vn_p.t517 704.872
R1374 vn_p.n771 vn_p.t871 704.872
R1375 vn_p.n772 vn_p.t321 704.872
R1376 vn_p.n773 vn_p.t669 704.872
R1377 vn_p.n774 vn_p.t129 704.872
R1378 vn_p.n775 vn_p.t1329 704.872
R1379 vn_p.n776 vn_p.t789 704.872
R1380 vn_p.n777 vn_p.t1125 704.872
R1381 vn_p.n778 vn_p.t1467 704.872
R1382 vn_p.n779 vn_p.t925 704.872
R1383 vn_p.n780 vn_p.t630 704.872
R1384 vn_p.n781 vn_p.t91 704.872
R1385 vn_p.n782 vn_p.t437 704.872
R1386 vn_p.n783 vn_p.t781 704.872
R1387 vn_p.n784 vn_p.t1081 704.872
R1388 vn_p.n785 vn_p.t799 704.872
R1389 vn_p.n786 vn_p.t246 704.872
R1390 vn_p.n787 vn_p.t594 704.872
R1391 vn_p.n788 vn_p.t44 704.872
R1392 vn_p.n789 vn_p.t385 704.872
R1393 vn_p.n790 vn_p.t98 704.872
R1394 vn_p.n791 vn_p.t1047 704.872
R1395 vn_p.n792 vn_p.t1400 704.872
R1396 vn_p.n793 vn_p.t848 704.872
R1397 vn_p.n794 vn_p.t1185 704.872
R1398 vn_p.n795 vn_p.t2 704.872
R1399 vn_p.n796 vn_p.t345 704.872
R1400 vn_p.n797 vn_p.t699 704.872
R1401 vn_p.n798 vn_p.t154 704.872
R1402 vn_p.n799 vn_p.t495 704.872
R1403 vn_p.n800 vn_p.t812 704.872
R1404 vn_p.n801 vn_p.t1151 704.872
R1405 vn_p.n802 vn_p.t1497 704.872
R1406 vn_p.n803 vn_p.t953 704.872
R1407 vn_p.n804 vn_p.t1300 704.872
R1408 vn_p.n805 vn_p.t117 704.872
R1409 vn_p.n806 vn_p.t467 704.872
R1410 vn_p.n807 vn_p.t370 704.872
R1411 vn_p.n808 vn_p.t725 704.872
R1412 vn_p.n809 vn_p.t1065 704.872
R1413 vn_p.n810 vn_p.t1388 704.872
R1414 vn_p.n811 vn_p.t231 704.872
R1415 vn_p.n812 vn_p.t1174 704.872
R1416 vn_p.n813 vn_p.t27 704.872
R1417 vn_p.n814 vn_p.t368 704.872
R1418 vn_p.n815 vn_p.t686 704.872
R1419 vn_p.n816 vn_p.t1032 704.872
R1420 vn_p.n817 vn_p.t489 704.872
R1421 vn_p.n818 vn_p.t836 704.872
R1422 vn_p.n819 vn_p.t277 704.872
R1423 vn_p.n820 vn_p.t1482 704.872
R1424 vn_p.n821 vn_p.t329 704.872
R1425 vn_p.n822 vn_p.t1287 704.872
R1426 vn_p.n1419 vn_p.t965 704.872
R1427 vn_p.n1420 vn_p.t421 704.872
R1428 vn_p.n1421 vn_p.t764 704.872
R1429 vn_p.n1422 vn_p.t221 704.872
R1430 vn_p.n1423 vn_p.t563 704.872
R1431 vn_p.n1424 vn_p.t874 704.872
R1432 vn_p.n1425 vn_p.t1213 704.872
R1433 vn_p.n1426 vn_p.t68 704.872
R1434 vn_p.n1427 vn_p.t1023 704.872
R1435 vn_p.n1428 vn_p.t1373 704.872
R1436 vn_p.n1429 vn_p.t1035 704.872
R1437 vn_p.n1430 vn_p.t1386 704.872
R1438 vn_p.n1431 vn_p.t229 704.872
R1439 vn_p.n1432 vn_p.t1171 704.872
R1440 vn_p.n1433 vn_p.t25 704.872
R1441 vn_p.n1434 vn_p.t332 704.872
R1442 vn_p.n1435 vn_p.t682 704.872
R1443 vn_p.n1436 vn_p.t141 704.872
R1444 vn_p.n1437 vn_p.t486 704.872
R1445 vn_p.n1438 vn_p.t835 704.872
R1446 vn_p.n1439 vn_p.t1139 704.872
R1447 vn_p.n1440 vn_p.t1478 704.872
R1448 vn_p.n1441 vn_p.t939 704.872
R1449 vn_p.n1442 vn_p.t1283 704.872
R1450 vn_p.n1443 vn_p.t137 704.872
R1451 vn_p.n1444 vn_p.t448 704.872
R1452 vn_p.n1445 vn_p.t794 704.872
R1453 vn_p.n1446 vn_p.t244 704.872
R1454 vn_p.n1447 vn_p.t590 704.872
R1455 vn_p.n1448 vn_p.t41 704.872
R1456 vn_p.n1449 vn_p.t1240 704.872
R1457 vn_p.n1450 vn_p.t96 704.872
R1458 vn_p.n1451 vn_p.t1045 704.872
R1459 vn_p.n1452 vn_p.t1397 704.872
R1460 vn_p.n1453 vn_p.t205 704.872
R1461 vn_p.n1454 vn_p.t1408 704.872
R1462 vn_p.n1455 vn_p.t861 704.872
R1463 vn_p.n1456 vn_p.t1195 704.872
R1464 vn_p.n1457 vn_p.t49 704.872
R1465 vn_p.n1458 vn_p.t1006 704.872
R1466 vn_p.n1459 vn_p.t707 704.872
R1467 vn_p.n1460 vn_p.t165 704.872
R1468 vn_p.n1461 vn_p.t503 704.872
R1469 vn_p.n1462 vn_p.t854 704.872
R1470 vn_p.n1463 vn_p.t299 704.872
R1471 vn_p.n1464 vn_p.t10 704.872
R1472 vn_p.n1465 vn_p.t966 704.872
R1473 vn_p.n1466 vn_p.t1309 704.872
R1474 vn_p.n1467 vn_p.t765 704.872
R1475 vn_p.n1468 vn_p.t1106 704.872
R1476 vn_p.n1469 vn_p.t819 704.872
R1477 vn_p.n1470 vn_p.t263 704.872
R1478 vn_p.n1471 vn_p.t614 704.872
R1479 vn_p.n1472 vn_p.t69 704.872
R1480 vn_p.n1473 vn_p.t416 704.872
R1481 vn_p.n1474 vn_p.t726 704.872
R1482 vn_p.n1475 vn_p.t1066 704.872
R1483 vn_p.n1476 vn_p.t1421 704.872
R1484 vn_p.n1477 vn_p.t1335 704.872
R1485 vn_p.n1478 vn_p.t186 704.872
R1486 vn_p.n1479 vn_p.t493 704.872
R1487 vn_p.n1480 vn_p.t843 704.872
R1488 vn_p.n1481 vn_p.t1178 704.872
R1489 vn_p.n1482 vn_p.t635 704.872
R1490 vn_p.n1483 vn_p.t988 704.872
R1491 vn_p.n1484 vn_p.t1296 704.872
R1492 vn_p.n1485 vn_p.t147 704.872
R1493 vn_p.n1486 vn_p.t1088 704.872
R1494 vn_p.n1487 vn_p.t1438 704.872
R1495 vn_p.n1488 vn_p.t282 704.872
R1496 vn_p.n1489 vn_p.t601 704.872
R1497 vn_p.n1490 vn_p.t946 704.872
R1498 vn_p.n1491 vn_p.t395 704.872
R1499 vn_p.n1492 vn_p.t747 704.872
R1500 vn_p.n744 vn_p.n743 1.225
R1501 vn_p.n671 vn_p.n670 1.141
R1502 vn_p.n672 vn_p.n671 1.141
R1503 vn_p.n673 vn_p.n672 1.141
R1504 vn_p.n674 vn_p.n673 1.141
R1505 vn_p.n675 vn_p.n674 1.141
R1506 vn_p.n676 vn_p.n675 1.141
R1507 vn_p.n677 vn_p.n676 1.141
R1508 vn_p.n678 vn_p.n677 1.141
R1509 vn_p.n679 vn_p.n678 1.141
R1510 vn_p.n680 vn_p.n679 1.141
R1511 vn_p.n681 vn_p.n680 1.141
R1512 vn_p.n682 vn_p.n681 1.141
R1513 vn_p.n683 vn_p.n682 1.141
R1514 vn_p.n684 vn_p.n683 1.141
R1515 vn_p.n685 vn_p.n684 1.141
R1516 vn_p.n686 vn_p.n685 1.141
R1517 vn_p.n687 vn_p.n686 1.141
R1518 vn_p.n688 vn_p.n687 1.141
R1519 vn_p.n689 vn_p.n688 1.141
R1520 vn_p.n690 vn_p.n689 1.141
R1521 vn_p.n691 vn_p.n690 1.141
R1522 vn_p.n692 vn_p.n691 1.141
R1523 vn_p.n693 vn_p.n692 1.141
R1524 vn_p.n694 vn_p.n693 1.141
R1525 vn_p.n695 vn_p.n694 1.141
R1526 vn_p.n696 vn_p.n695 1.141
R1527 vn_p.n697 vn_p.n696 1.141
R1528 vn_p.n698 vn_p.n697 1.141
R1529 vn_p.n699 vn_p.n698 1.141
R1530 vn_p.n700 vn_p.n699 1.141
R1531 vn_p.n701 vn_p.n700 1.141
R1532 vn_p.n702 vn_p.n701 1.141
R1533 vn_p.n703 vn_p.n702 1.141
R1534 vn_p.n704 vn_p.n703 1.141
R1535 vn_p.n705 vn_p.n704 1.141
R1536 vn_p.n706 vn_p.n705 1.141
R1537 vn_p.n707 vn_p.n706 1.141
R1538 vn_p.n708 vn_p.n707 1.141
R1539 vn_p.n709 vn_p.n708 1.141
R1540 vn_p.n710 vn_p.n709 1.141
R1541 vn_p.n711 vn_p.n710 1.141
R1542 vn_p.n712 vn_p.n711 1.141
R1543 vn_p.n713 vn_p.n712 1.141
R1544 vn_p.n714 vn_p.n713 1.141
R1545 vn_p.n715 vn_p.n714 1.141
R1546 vn_p.n716 vn_p.n715 1.141
R1547 vn_p.n717 vn_p.n716 1.141
R1548 vn_p.n718 vn_p.n717 1.141
R1549 vn_p.n719 vn_p.n718 1.141
R1550 vn_p.n720 vn_p.n719 1.141
R1551 vn_p.n721 vn_p.n720 1.141
R1552 vn_p.n722 vn_p.n721 1.141
R1553 vn_p.n723 vn_p.n722 1.141
R1554 vn_p.n724 vn_p.n723 1.141
R1555 vn_p.n725 vn_p.n724 1.141
R1556 vn_p.n726 vn_p.n725 1.141
R1557 vn_p.n727 vn_p.n726 1.141
R1558 vn_p.n728 vn_p.n727 1.141
R1559 vn_p.n729 vn_p.n728 1.141
R1560 vn_p.n730 vn_p.n729 1.141
R1561 vn_p.n731 vn_p.n730 1.141
R1562 vn_p.n732 vn_p.n731 1.141
R1563 vn_p.n733 vn_p.n732 1.141
R1564 vn_p.n734 vn_p.n733 1.141
R1565 vn_p.n735 vn_p.n734 1.141
R1566 vn_p.n736 vn_p.n735 1.141
R1567 vn_p.n737 vn_p.n736 1.141
R1568 vn_p.n738 vn_p.n737 1.141
R1569 vn_p.n739 vn_p.n738 1.141
R1570 vn_p.n740 vn_p.n739 1.141
R1571 vn_p.n741 vn_p.n740 1.141
R1572 vn_p.n742 vn_p.n741 1.141
R1573 vn_p.n743 vn_p.n742 1.141
R1574 vn_p.n750 vn_p.n749 1.141
R1575 vn_p.n751 vn_p.n750 1.141
R1576 vn_p.n752 vn_p.n751 1.141
R1577 vn_p.n753 vn_p.n752 1.141
R1578 vn_p.n754 vn_p.n753 1.141
R1579 vn_p.n755 vn_p.n754 1.141
R1580 vn_p.n756 vn_p.n755 1.141
R1581 vn_p.n757 vn_p.n756 1.141
R1582 vn_p.n758 vn_p.n757 1.141
R1583 vn_p.n759 vn_p.n758 1.141
R1584 vn_p.n760 vn_p.n759 1.141
R1585 vn_p.n761 vn_p.n760 1.141
R1586 vn_p.n762 vn_p.n761 1.141
R1587 vn_p.n763 vn_p.n762 1.141
R1588 vn_p.n764 vn_p.n763 1.141
R1589 vn_p.n765 vn_p.n764 1.141
R1590 vn_p.n766 vn_p.n765 1.141
R1591 vn_p.n767 vn_p.n766 1.141
R1592 vn_p.n768 vn_p.n767 1.141
R1593 vn_p.n769 vn_p.n768 1.141
R1594 vn_p.n770 vn_p.n769 1.141
R1595 vn_p.n771 vn_p.n770 1.141
R1596 vn_p.n772 vn_p.n771 1.141
R1597 vn_p.n773 vn_p.n772 1.141
R1598 vn_p.n774 vn_p.n773 1.141
R1599 vn_p.n775 vn_p.n774 1.141
R1600 vn_p.n776 vn_p.n775 1.141
R1601 vn_p.n777 vn_p.n776 1.141
R1602 vn_p.n778 vn_p.n777 1.141
R1603 vn_p.n779 vn_p.n778 1.141
R1604 vn_p.n780 vn_p.n779 1.141
R1605 vn_p.n781 vn_p.n780 1.141
R1606 vn_p.n782 vn_p.n781 1.141
R1607 vn_p.n783 vn_p.n782 1.141
R1608 vn_p.n784 vn_p.n783 1.141
R1609 vn_p.n785 vn_p.n784 1.141
R1610 vn_p.n786 vn_p.n785 1.141
R1611 vn_p.n787 vn_p.n786 1.141
R1612 vn_p.n788 vn_p.n787 1.141
R1613 vn_p.n789 vn_p.n788 1.141
R1614 vn_p.n790 vn_p.n789 1.141
R1615 vn_p.n791 vn_p.n790 1.141
R1616 vn_p.n792 vn_p.n791 1.141
R1617 vn_p.n793 vn_p.n792 1.141
R1618 vn_p.n794 vn_p.n793 1.141
R1619 vn_p.n795 vn_p.n794 1.141
R1620 vn_p.n796 vn_p.n795 1.141
R1621 vn_p.n797 vn_p.n796 1.141
R1622 vn_p.n798 vn_p.n797 1.141
R1623 vn_p.n799 vn_p.n798 1.141
R1624 vn_p.n800 vn_p.n799 1.141
R1625 vn_p.n801 vn_p.n800 1.141
R1626 vn_p.n802 vn_p.n801 1.141
R1627 vn_p.n803 vn_p.n802 1.141
R1628 vn_p.n804 vn_p.n803 1.141
R1629 vn_p.n805 vn_p.n804 1.141
R1630 vn_p.n806 vn_p.n805 1.141
R1631 vn_p.n807 vn_p.n806 1.141
R1632 vn_p.n808 vn_p.n807 1.141
R1633 vn_p.n809 vn_p.n808 1.141
R1634 vn_p.n810 vn_p.n809 1.141
R1635 vn_p.n811 vn_p.n810 1.141
R1636 vn_p.n812 vn_p.n811 1.141
R1637 vn_p.n813 vn_p.n812 1.141
R1638 vn_p.n814 vn_p.n813 1.141
R1639 vn_p.n815 vn_p.n814 1.141
R1640 vn_p.n816 vn_p.n815 1.141
R1641 vn_p.n817 vn_p.n816 1.141
R1642 vn_p.n818 vn_p.n817 1.141
R1643 vn_p.n819 vn_p.n818 1.141
R1644 vn_p.n820 vn_p.n819 1.141
R1645 vn_p.n821 vn_p.n820 1.141
R1646 vn_p.n822 vn_p.n821 1.141
R1647 vn_p.n1420 vn_p.n1419 1.141
R1648 vn_p.n1421 vn_p.n1420 1.141
R1649 vn_p.n1422 vn_p.n1421 1.141
R1650 vn_p.n1423 vn_p.n1422 1.141
R1651 vn_p.n1424 vn_p.n1423 1.141
R1652 vn_p.n1425 vn_p.n1424 1.141
R1653 vn_p.n1426 vn_p.n1425 1.141
R1654 vn_p.n1427 vn_p.n1426 1.141
R1655 vn_p.n1428 vn_p.n1427 1.141
R1656 vn_p.n1429 vn_p.n1428 1.141
R1657 vn_p.n1430 vn_p.n1429 1.141
R1658 vn_p.n1431 vn_p.n1430 1.141
R1659 vn_p.n1432 vn_p.n1431 1.141
R1660 vn_p.n1433 vn_p.n1432 1.141
R1661 vn_p.n1434 vn_p.n1433 1.141
R1662 vn_p.n1435 vn_p.n1434 1.141
R1663 vn_p.n1436 vn_p.n1435 1.141
R1664 vn_p.n1437 vn_p.n1436 1.141
R1665 vn_p.n1438 vn_p.n1437 1.141
R1666 vn_p.n1439 vn_p.n1438 1.141
R1667 vn_p.n1440 vn_p.n1439 1.141
R1668 vn_p.n1441 vn_p.n1440 1.141
R1669 vn_p.n1442 vn_p.n1441 1.141
R1670 vn_p.n1443 vn_p.n1442 1.141
R1671 vn_p.n1444 vn_p.n1443 1.141
R1672 vn_p.n1445 vn_p.n1444 1.141
R1673 vn_p.n1446 vn_p.n1445 1.141
R1674 vn_p.n1447 vn_p.n1446 1.141
R1675 vn_p.n1448 vn_p.n1447 1.141
R1676 vn_p.n1449 vn_p.n1448 1.141
R1677 vn_p.n1450 vn_p.n1449 1.141
R1678 vn_p.n1451 vn_p.n1450 1.141
R1679 vn_p.n1452 vn_p.n1451 1.141
R1680 vn_p.n1453 vn_p.n1452 1.141
R1681 vn_p.n1454 vn_p.n1453 1.141
R1682 vn_p.n1455 vn_p.n1454 1.141
R1683 vn_p.n1456 vn_p.n1455 1.141
R1684 vn_p.n1457 vn_p.n1456 1.141
R1685 vn_p.n1458 vn_p.n1457 1.141
R1686 vn_p.n1459 vn_p.n1458 1.141
R1687 vn_p.n1460 vn_p.n1459 1.141
R1688 vn_p.n1461 vn_p.n1460 1.141
R1689 vn_p.n1462 vn_p.n1461 1.141
R1690 vn_p.n1463 vn_p.n1462 1.141
R1691 vn_p.n1464 vn_p.n1463 1.141
R1692 vn_p.n1465 vn_p.n1464 1.141
R1693 vn_p.n1466 vn_p.n1465 1.141
R1694 vn_p.n1467 vn_p.n1466 1.141
R1695 vn_p.n1468 vn_p.n1467 1.141
R1696 vn_p.n1469 vn_p.n1468 1.141
R1697 vn_p.n1470 vn_p.n1469 1.141
R1698 vn_p.n1471 vn_p.n1470 1.141
R1699 vn_p.n1472 vn_p.n1471 1.141
R1700 vn_p.n1473 vn_p.n1472 1.141
R1701 vn_p.n1474 vn_p.n1473 1.141
R1702 vn_p.n1475 vn_p.n1474 1.141
R1703 vn_p.n1476 vn_p.n1475 1.141
R1704 vn_p.n1477 vn_p.n1476 1.141
R1705 vn_p.n1478 vn_p.n1477 1.141
R1706 vn_p.n1479 vn_p.n1478 1.141
R1707 vn_p.n1480 vn_p.n1479 1.141
R1708 vn_p.n1481 vn_p.n1480 1.141
R1709 vn_p.n1482 vn_p.n1481 1.141
R1710 vn_p.n1483 vn_p.n1482 1.141
R1711 vn_p.n1484 vn_p.n1483 1.141
R1712 vn_p.n1485 vn_p.n1484 1.141
R1713 vn_p.n1486 vn_p.n1485 1.141
R1714 vn_p.n1487 vn_p.n1486 1.141
R1715 vn_p.n1488 vn_p.n1487 1.141
R1716 vn_p.n1489 vn_p.n1488 1.141
R1717 vn_p.n1490 vn_p.n1489 1.141
R1718 vn_p.n1491 vn_p.n1490 1.141
R1719 vn_p.n1492 vn_p.n1491 1.141
R1720 vn_p.n1 vn_p.n0 1.117
R1721 vn_p.n2 vn_p.n1 1.117
R1722 vn_p.n3 vn_p.n2 1.117
R1723 vn_p.n4 vn_p.n3 1.117
R1724 vn_p.n5 vn_p.n4 1.117
R1725 vn_p.n6 vn_p.n5 1.117
R1726 vn_p.n7 vn_p.n6 1.117
R1727 vn_p.n8 vn_p.n7 1.117
R1728 vn_p.n9 vn_p.n8 1.117
R1729 vn_p.n10 vn_p.n9 1.117
R1730 vn_p.n11 vn_p.n10 1.117
R1731 vn_p.n12 vn_p.n11 1.117
R1732 vn_p.n13 vn_p.n12 1.117
R1733 vn_p.n14 vn_p.n13 1.117
R1734 vn_p.n15 vn_p.n14 1.117
R1735 vn_p.n16 vn_p.n15 1.117
R1736 vn_p.n17 vn_p.n16 1.117
R1737 vn_p.n18 vn_p.n17 1.117
R1738 vn_p.n19 vn_p.n18 1.117
R1739 vn_p.n20 vn_p.n19 1.117
R1740 vn_p.n21 vn_p.n20 1.117
R1741 vn_p.n22 vn_p.n21 1.117
R1742 vn_p.n23 vn_p.n22 1.117
R1743 vn_p.n24 vn_p.n23 1.117
R1744 vn_p.n25 vn_p.n24 1.117
R1745 vn_p.n26 vn_p.n25 1.117
R1746 vn_p.n27 vn_p.n26 1.117
R1747 vn_p.n28 vn_p.n27 1.117
R1748 vn_p.n29 vn_p.n28 1.117
R1749 vn_p.n30 vn_p.n29 1.117
R1750 vn_p.n31 vn_p.n30 1.117
R1751 vn_p.n32 vn_p.n31 1.117
R1752 vn_p.n33 vn_p.n32 1.117
R1753 vn_p.n34 vn_p.n33 1.117
R1754 vn_p.n35 vn_p.n34 1.117
R1755 vn_p.n36 vn_p.n35 1.117
R1756 vn_p.n37 vn_p.n36 1.117
R1757 vn_p.n38 vn_p.n37 1.117
R1758 vn_p.n39 vn_p.n38 1.117
R1759 vn_p.n40 vn_p.n39 1.117
R1760 vn_p.n41 vn_p.n40 1.117
R1761 vn_p.n42 vn_p.n41 1.117
R1762 vn_p.n43 vn_p.n42 1.117
R1763 vn_p.n44 vn_p.n43 1.117
R1764 vn_p.n45 vn_p.n44 1.117
R1765 vn_p.n46 vn_p.n45 1.117
R1766 vn_p.n47 vn_p.n46 1.117
R1767 vn_p.n48 vn_p.n47 1.117
R1768 vn_p.n49 vn_p.n48 1.117
R1769 vn_p.n50 vn_p.n49 1.117
R1770 vn_p.n51 vn_p.n50 1.117
R1771 vn_p.n52 vn_p.n51 1.117
R1772 vn_p.n53 vn_p.n52 1.117
R1773 vn_p.n54 vn_p.n53 1.117
R1774 vn_p.n55 vn_p.n54 1.117
R1775 vn_p.n56 vn_p.n55 1.117
R1776 vn_p.n57 vn_p.n56 1.117
R1777 vn_p.n58 vn_p.n57 1.117
R1778 vn_p.n59 vn_p.n58 1.117
R1779 vn_p.n60 vn_p.n59 1.117
R1780 vn_p.n61 vn_p.n60 1.117
R1781 vn_p.n62 vn_p.n61 1.117
R1782 vn_p.n63 vn_p.n62 1.117
R1783 vn_p.n64 vn_p.n63 1.117
R1784 vn_p.n65 vn_p.n64 1.117
R1785 vn_p.n66 vn_p.n65 1.117
R1786 vn_p.n67 vn_p.n66 1.117
R1787 vn_p.n68 vn_p.n67 1.117
R1788 vn_p.n69 vn_p.n68 1.117
R1789 vn_p.n70 vn_p.n69 1.117
R1790 vn_p.n71 vn_p.n70 1.117
R1791 vn_p.n72 vn_p.n71 1.117
R1792 vn_p.n73 vn_p.n72 1.117
R1793 vn_p.n1497 vn_p.n822 1.084
R1794 vn_p.n1493 vn_p.n1492 0.654
R1795 vn_p.n748 vn_p.n73 0.509
R1796 vn_p.n523 vn_p.n521 0.356
R1797 vn_p.n374 vn_p.n372 0.356
R1798 vn_p.n225 vn_p.n223 0.356
R1799 vn_p.n76 vn_p.n74 0.356
R1800 vn_p.n825 vn_p.n823 0.356
R1801 vn_p.n974 vn_p.n972 0.356
R1802 vn_p.n1123 vn_p.n1121 0.356
R1803 vn_p.n1272 vn_p.n1270 0.356
R1804 vn_p.n745 vn_p.n520 0.319
R1805 vn_p.n747 vn_p.n222 0.319
R1806 vn_p.n1495 vn_p.n1120 0.319
R1807 vn_p.n1493 vn_p.n1418 0.319
R1808 vn_p.n525 vn_p.n523 0.316
R1809 vn_p.n527 vn_p.n525 0.316
R1810 vn_p.n529 vn_p.n527 0.316
R1811 vn_p.n531 vn_p.n529 0.316
R1812 vn_p.n533 vn_p.n531 0.316
R1813 vn_p.n535 vn_p.n533 0.316
R1814 vn_p.n537 vn_p.n535 0.316
R1815 vn_p.n539 vn_p.n537 0.316
R1816 vn_p.n541 vn_p.n539 0.316
R1817 vn_p.n543 vn_p.n541 0.316
R1818 vn_p.n545 vn_p.n543 0.316
R1819 vn_p.n547 vn_p.n545 0.316
R1820 vn_p.n549 vn_p.n547 0.316
R1821 vn_p.n551 vn_p.n549 0.316
R1822 vn_p.n553 vn_p.n551 0.316
R1823 vn_p.n555 vn_p.n553 0.316
R1824 vn_p.n557 vn_p.n555 0.316
R1825 vn_p.n559 vn_p.n557 0.316
R1826 vn_p.n561 vn_p.n559 0.316
R1827 vn_p.n563 vn_p.n561 0.316
R1828 vn_p.n565 vn_p.n563 0.316
R1829 vn_p.n567 vn_p.n565 0.316
R1830 vn_p.n569 vn_p.n567 0.316
R1831 vn_p.n571 vn_p.n569 0.316
R1832 vn_p.n573 vn_p.n571 0.316
R1833 vn_p.n575 vn_p.n573 0.316
R1834 vn_p.n577 vn_p.n575 0.316
R1835 vn_p.n579 vn_p.n577 0.316
R1836 vn_p.n581 vn_p.n579 0.316
R1837 vn_p.n583 vn_p.n581 0.316
R1838 vn_p.n585 vn_p.n583 0.316
R1839 vn_p.n587 vn_p.n585 0.316
R1840 vn_p.n589 vn_p.n587 0.316
R1841 vn_p.n591 vn_p.n589 0.316
R1842 vn_p.n593 vn_p.n591 0.316
R1843 vn_p.n595 vn_p.n593 0.316
R1844 vn_p.n597 vn_p.n595 0.316
R1845 vn_p.n599 vn_p.n597 0.316
R1846 vn_p.n601 vn_p.n599 0.316
R1847 vn_p.n603 vn_p.n601 0.316
R1848 vn_p.n605 vn_p.n603 0.316
R1849 vn_p.n607 vn_p.n605 0.316
R1850 vn_p.n609 vn_p.n607 0.316
R1851 vn_p.n611 vn_p.n609 0.316
R1852 vn_p.n613 vn_p.n611 0.316
R1853 vn_p.n615 vn_p.n613 0.316
R1854 vn_p.n617 vn_p.n615 0.316
R1855 vn_p.n619 vn_p.n617 0.316
R1856 vn_p.n621 vn_p.n619 0.316
R1857 vn_p.n623 vn_p.n621 0.316
R1858 vn_p.n625 vn_p.n623 0.316
R1859 vn_p.n627 vn_p.n625 0.316
R1860 vn_p.n629 vn_p.n627 0.316
R1861 vn_p.n631 vn_p.n629 0.316
R1862 vn_p.n633 vn_p.n631 0.316
R1863 vn_p.n635 vn_p.n633 0.316
R1864 vn_p.n637 vn_p.n635 0.316
R1865 vn_p.n639 vn_p.n637 0.316
R1866 vn_p.n641 vn_p.n639 0.316
R1867 vn_p.n643 vn_p.n641 0.316
R1868 vn_p.n645 vn_p.n643 0.316
R1869 vn_p.n647 vn_p.n645 0.316
R1870 vn_p.n649 vn_p.n647 0.316
R1871 vn_p.n651 vn_p.n649 0.316
R1872 vn_p.n653 vn_p.n651 0.316
R1873 vn_p.n655 vn_p.n653 0.316
R1874 vn_p.n657 vn_p.n655 0.316
R1875 vn_p.n659 vn_p.n657 0.316
R1876 vn_p.n661 vn_p.n659 0.316
R1877 vn_p.n663 vn_p.n661 0.316
R1878 vn_p.n665 vn_p.n663 0.316
R1879 vn_p.n667 vn_p.n665 0.316
R1880 vn_p.n669 vn_p.n667 0.316
R1881 vn_p.n376 vn_p.n374 0.316
R1882 vn_p.n378 vn_p.n376 0.316
R1883 vn_p.n380 vn_p.n378 0.316
R1884 vn_p.n382 vn_p.n380 0.316
R1885 vn_p.n384 vn_p.n382 0.316
R1886 vn_p.n386 vn_p.n384 0.316
R1887 vn_p.n388 vn_p.n386 0.316
R1888 vn_p.n390 vn_p.n388 0.316
R1889 vn_p.n392 vn_p.n390 0.316
R1890 vn_p.n394 vn_p.n392 0.316
R1891 vn_p.n396 vn_p.n394 0.316
R1892 vn_p.n398 vn_p.n396 0.316
R1893 vn_p.n400 vn_p.n398 0.316
R1894 vn_p.n402 vn_p.n400 0.316
R1895 vn_p.n404 vn_p.n402 0.316
R1896 vn_p.n406 vn_p.n404 0.316
R1897 vn_p.n408 vn_p.n406 0.316
R1898 vn_p.n410 vn_p.n408 0.316
R1899 vn_p.n412 vn_p.n410 0.316
R1900 vn_p.n414 vn_p.n412 0.316
R1901 vn_p.n416 vn_p.n414 0.316
R1902 vn_p.n418 vn_p.n416 0.316
R1903 vn_p.n420 vn_p.n418 0.316
R1904 vn_p.n422 vn_p.n420 0.316
R1905 vn_p.n424 vn_p.n422 0.316
R1906 vn_p.n426 vn_p.n424 0.316
R1907 vn_p.n428 vn_p.n426 0.316
R1908 vn_p.n430 vn_p.n428 0.316
R1909 vn_p.n432 vn_p.n430 0.316
R1910 vn_p.n434 vn_p.n432 0.316
R1911 vn_p.n436 vn_p.n434 0.316
R1912 vn_p.n438 vn_p.n436 0.316
R1913 vn_p.n440 vn_p.n438 0.316
R1914 vn_p.n442 vn_p.n440 0.316
R1915 vn_p.n444 vn_p.n442 0.316
R1916 vn_p.n446 vn_p.n444 0.316
R1917 vn_p.n448 vn_p.n446 0.316
R1918 vn_p.n450 vn_p.n448 0.316
R1919 vn_p.n452 vn_p.n450 0.316
R1920 vn_p.n454 vn_p.n452 0.316
R1921 vn_p.n456 vn_p.n454 0.316
R1922 vn_p.n458 vn_p.n456 0.316
R1923 vn_p.n460 vn_p.n458 0.316
R1924 vn_p.n462 vn_p.n460 0.316
R1925 vn_p.n464 vn_p.n462 0.316
R1926 vn_p.n466 vn_p.n464 0.316
R1927 vn_p.n468 vn_p.n466 0.316
R1928 vn_p.n470 vn_p.n468 0.316
R1929 vn_p.n472 vn_p.n470 0.316
R1930 vn_p.n474 vn_p.n472 0.316
R1931 vn_p.n476 vn_p.n474 0.316
R1932 vn_p.n478 vn_p.n476 0.316
R1933 vn_p.n480 vn_p.n478 0.316
R1934 vn_p.n482 vn_p.n480 0.316
R1935 vn_p.n484 vn_p.n482 0.316
R1936 vn_p.n486 vn_p.n484 0.316
R1937 vn_p.n488 vn_p.n486 0.316
R1938 vn_p.n490 vn_p.n488 0.316
R1939 vn_p.n492 vn_p.n490 0.316
R1940 vn_p.n494 vn_p.n492 0.316
R1941 vn_p.n496 vn_p.n494 0.316
R1942 vn_p.n498 vn_p.n496 0.316
R1943 vn_p.n500 vn_p.n498 0.316
R1944 vn_p.n502 vn_p.n500 0.316
R1945 vn_p.n504 vn_p.n502 0.316
R1946 vn_p.n506 vn_p.n504 0.316
R1947 vn_p.n508 vn_p.n506 0.316
R1948 vn_p.n510 vn_p.n508 0.316
R1949 vn_p.n512 vn_p.n510 0.316
R1950 vn_p.n514 vn_p.n512 0.316
R1951 vn_p.n516 vn_p.n514 0.316
R1952 vn_p.n518 vn_p.n516 0.316
R1953 vn_p.n520 vn_p.n518 0.316
R1954 vn_p.n227 vn_p.n225 0.316
R1955 vn_p.n229 vn_p.n227 0.316
R1956 vn_p.n231 vn_p.n229 0.316
R1957 vn_p.n233 vn_p.n231 0.316
R1958 vn_p.n235 vn_p.n233 0.316
R1959 vn_p.n237 vn_p.n235 0.316
R1960 vn_p.n239 vn_p.n237 0.316
R1961 vn_p.n241 vn_p.n239 0.316
R1962 vn_p.n243 vn_p.n241 0.316
R1963 vn_p.n245 vn_p.n243 0.316
R1964 vn_p.n247 vn_p.n245 0.316
R1965 vn_p.n249 vn_p.n247 0.316
R1966 vn_p.n251 vn_p.n249 0.316
R1967 vn_p.n253 vn_p.n251 0.316
R1968 vn_p.n255 vn_p.n253 0.316
R1969 vn_p.n257 vn_p.n255 0.316
R1970 vn_p.n259 vn_p.n257 0.316
R1971 vn_p.n261 vn_p.n259 0.316
R1972 vn_p.n263 vn_p.n261 0.316
R1973 vn_p.n265 vn_p.n263 0.316
R1974 vn_p.n267 vn_p.n265 0.316
R1975 vn_p.n269 vn_p.n267 0.316
R1976 vn_p.n271 vn_p.n269 0.316
R1977 vn_p.n273 vn_p.n271 0.316
R1978 vn_p.n275 vn_p.n273 0.316
R1979 vn_p.n277 vn_p.n275 0.316
R1980 vn_p.n279 vn_p.n277 0.316
R1981 vn_p.n281 vn_p.n279 0.316
R1982 vn_p.n283 vn_p.n281 0.316
R1983 vn_p.n285 vn_p.n283 0.316
R1984 vn_p.n287 vn_p.n285 0.316
R1985 vn_p.n289 vn_p.n287 0.316
R1986 vn_p.n291 vn_p.n289 0.316
R1987 vn_p.n293 vn_p.n291 0.316
R1988 vn_p.n295 vn_p.n293 0.316
R1989 vn_p.n297 vn_p.n295 0.316
R1990 vn_p.n299 vn_p.n297 0.316
R1991 vn_p.n301 vn_p.n299 0.316
R1992 vn_p.n303 vn_p.n301 0.316
R1993 vn_p.n305 vn_p.n303 0.316
R1994 vn_p.n307 vn_p.n305 0.316
R1995 vn_p.n309 vn_p.n307 0.316
R1996 vn_p.n311 vn_p.n309 0.316
R1997 vn_p.n313 vn_p.n311 0.316
R1998 vn_p.n315 vn_p.n313 0.316
R1999 vn_p.n317 vn_p.n315 0.316
R2000 vn_p.n319 vn_p.n317 0.316
R2001 vn_p.n321 vn_p.n319 0.316
R2002 vn_p.n323 vn_p.n321 0.316
R2003 vn_p.n325 vn_p.n323 0.316
R2004 vn_p.n327 vn_p.n325 0.316
R2005 vn_p.n329 vn_p.n327 0.316
R2006 vn_p.n331 vn_p.n329 0.316
R2007 vn_p.n333 vn_p.n331 0.316
R2008 vn_p.n335 vn_p.n333 0.316
R2009 vn_p.n337 vn_p.n335 0.316
R2010 vn_p.n339 vn_p.n337 0.316
R2011 vn_p.n341 vn_p.n339 0.316
R2012 vn_p.n343 vn_p.n341 0.316
R2013 vn_p.n345 vn_p.n343 0.316
R2014 vn_p.n347 vn_p.n345 0.316
R2015 vn_p.n349 vn_p.n347 0.316
R2016 vn_p.n351 vn_p.n349 0.316
R2017 vn_p.n353 vn_p.n351 0.316
R2018 vn_p.n355 vn_p.n353 0.316
R2019 vn_p.n357 vn_p.n355 0.316
R2020 vn_p.n359 vn_p.n357 0.316
R2021 vn_p.n361 vn_p.n359 0.316
R2022 vn_p.n363 vn_p.n361 0.316
R2023 vn_p.n365 vn_p.n363 0.316
R2024 vn_p.n367 vn_p.n365 0.316
R2025 vn_p.n369 vn_p.n367 0.316
R2026 vn_p.n371 vn_p.n369 0.316
R2027 vn_p.n78 vn_p.n76 0.316
R2028 vn_p.n80 vn_p.n78 0.316
R2029 vn_p.n82 vn_p.n80 0.316
R2030 vn_p.n84 vn_p.n82 0.316
R2031 vn_p.n86 vn_p.n84 0.316
R2032 vn_p.n88 vn_p.n86 0.316
R2033 vn_p.n90 vn_p.n88 0.316
R2034 vn_p.n92 vn_p.n90 0.316
R2035 vn_p.n94 vn_p.n92 0.316
R2036 vn_p.n96 vn_p.n94 0.316
R2037 vn_p.n98 vn_p.n96 0.316
R2038 vn_p.n100 vn_p.n98 0.316
R2039 vn_p.n102 vn_p.n100 0.316
R2040 vn_p.n104 vn_p.n102 0.316
R2041 vn_p.n106 vn_p.n104 0.316
R2042 vn_p.n108 vn_p.n106 0.316
R2043 vn_p.n110 vn_p.n108 0.316
R2044 vn_p.n112 vn_p.n110 0.316
R2045 vn_p.n114 vn_p.n112 0.316
R2046 vn_p.n116 vn_p.n114 0.316
R2047 vn_p.n118 vn_p.n116 0.316
R2048 vn_p.n120 vn_p.n118 0.316
R2049 vn_p.n122 vn_p.n120 0.316
R2050 vn_p.n124 vn_p.n122 0.316
R2051 vn_p.n126 vn_p.n124 0.316
R2052 vn_p.n128 vn_p.n126 0.316
R2053 vn_p.n130 vn_p.n128 0.316
R2054 vn_p.n132 vn_p.n130 0.316
R2055 vn_p.n134 vn_p.n132 0.316
R2056 vn_p.n136 vn_p.n134 0.316
R2057 vn_p.n138 vn_p.n136 0.316
R2058 vn_p.n140 vn_p.n138 0.316
R2059 vn_p.n142 vn_p.n140 0.316
R2060 vn_p.n144 vn_p.n142 0.316
R2061 vn_p.n146 vn_p.n144 0.316
R2062 vn_p.n148 vn_p.n146 0.316
R2063 vn_p.n150 vn_p.n148 0.316
R2064 vn_p.n152 vn_p.n150 0.316
R2065 vn_p.n154 vn_p.n152 0.316
R2066 vn_p.n156 vn_p.n154 0.316
R2067 vn_p.n158 vn_p.n156 0.316
R2068 vn_p.n160 vn_p.n158 0.316
R2069 vn_p.n162 vn_p.n160 0.316
R2070 vn_p.n164 vn_p.n162 0.316
R2071 vn_p.n166 vn_p.n164 0.316
R2072 vn_p.n168 vn_p.n166 0.316
R2073 vn_p.n170 vn_p.n168 0.316
R2074 vn_p.n172 vn_p.n170 0.316
R2075 vn_p.n174 vn_p.n172 0.316
R2076 vn_p.n176 vn_p.n174 0.316
R2077 vn_p.n178 vn_p.n176 0.316
R2078 vn_p.n180 vn_p.n178 0.316
R2079 vn_p.n182 vn_p.n180 0.316
R2080 vn_p.n184 vn_p.n182 0.316
R2081 vn_p.n186 vn_p.n184 0.316
R2082 vn_p.n188 vn_p.n186 0.316
R2083 vn_p.n190 vn_p.n188 0.316
R2084 vn_p.n192 vn_p.n190 0.316
R2085 vn_p.n194 vn_p.n192 0.316
R2086 vn_p.n196 vn_p.n194 0.316
R2087 vn_p.n198 vn_p.n196 0.316
R2088 vn_p.n200 vn_p.n198 0.316
R2089 vn_p.n202 vn_p.n200 0.316
R2090 vn_p.n204 vn_p.n202 0.316
R2091 vn_p.n206 vn_p.n204 0.316
R2092 vn_p.n208 vn_p.n206 0.316
R2093 vn_p.n210 vn_p.n208 0.316
R2094 vn_p.n212 vn_p.n210 0.316
R2095 vn_p.n214 vn_p.n212 0.316
R2096 vn_p.n216 vn_p.n214 0.316
R2097 vn_p.n218 vn_p.n216 0.316
R2098 vn_p.n220 vn_p.n218 0.316
R2099 vn_p.n222 vn_p.n220 0.316
R2100 vn_p.n827 vn_p.n825 0.316
R2101 vn_p.n829 vn_p.n827 0.316
R2102 vn_p.n831 vn_p.n829 0.316
R2103 vn_p.n833 vn_p.n831 0.316
R2104 vn_p.n835 vn_p.n833 0.316
R2105 vn_p.n837 vn_p.n835 0.316
R2106 vn_p.n839 vn_p.n837 0.316
R2107 vn_p.n841 vn_p.n839 0.316
R2108 vn_p.n843 vn_p.n841 0.316
R2109 vn_p.n845 vn_p.n843 0.316
R2110 vn_p.n847 vn_p.n845 0.316
R2111 vn_p.n849 vn_p.n847 0.316
R2112 vn_p.n851 vn_p.n849 0.316
R2113 vn_p.n853 vn_p.n851 0.316
R2114 vn_p.n855 vn_p.n853 0.316
R2115 vn_p.n857 vn_p.n855 0.316
R2116 vn_p.n859 vn_p.n857 0.316
R2117 vn_p.n861 vn_p.n859 0.316
R2118 vn_p.n863 vn_p.n861 0.316
R2119 vn_p.n865 vn_p.n863 0.316
R2120 vn_p.n867 vn_p.n865 0.316
R2121 vn_p.n869 vn_p.n867 0.316
R2122 vn_p.n871 vn_p.n869 0.316
R2123 vn_p.n873 vn_p.n871 0.316
R2124 vn_p.n875 vn_p.n873 0.316
R2125 vn_p.n877 vn_p.n875 0.316
R2126 vn_p.n879 vn_p.n877 0.316
R2127 vn_p.n881 vn_p.n879 0.316
R2128 vn_p.n883 vn_p.n881 0.316
R2129 vn_p.n885 vn_p.n883 0.316
R2130 vn_p.n887 vn_p.n885 0.316
R2131 vn_p.n889 vn_p.n887 0.316
R2132 vn_p.n891 vn_p.n889 0.316
R2133 vn_p.n893 vn_p.n891 0.316
R2134 vn_p.n895 vn_p.n893 0.316
R2135 vn_p.n897 vn_p.n895 0.316
R2136 vn_p.n899 vn_p.n897 0.316
R2137 vn_p.n901 vn_p.n899 0.316
R2138 vn_p.n903 vn_p.n901 0.316
R2139 vn_p.n905 vn_p.n903 0.316
R2140 vn_p.n907 vn_p.n905 0.316
R2141 vn_p.n909 vn_p.n907 0.316
R2142 vn_p.n911 vn_p.n909 0.316
R2143 vn_p.n913 vn_p.n911 0.316
R2144 vn_p.n915 vn_p.n913 0.316
R2145 vn_p.n917 vn_p.n915 0.316
R2146 vn_p.n919 vn_p.n917 0.316
R2147 vn_p.n921 vn_p.n919 0.316
R2148 vn_p.n923 vn_p.n921 0.316
R2149 vn_p.n925 vn_p.n923 0.316
R2150 vn_p.n927 vn_p.n925 0.316
R2151 vn_p.n929 vn_p.n927 0.316
R2152 vn_p.n931 vn_p.n929 0.316
R2153 vn_p.n933 vn_p.n931 0.316
R2154 vn_p.n935 vn_p.n933 0.316
R2155 vn_p.n937 vn_p.n935 0.316
R2156 vn_p.n939 vn_p.n937 0.316
R2157 vn_p.n941 vn_p.n939 0.316
R2158 vn_p.n943 vn_p.n941 0.316
R2159 vn_p.n945 vn_p.n943 0.316
R2160 vn_p.n947 vn_p.n945 0.316
R2161 vn_p.n949 vn_p.n947 0.316
R2162 vn_p.n951 vn_p.n949 0.316
R2163 vn_p.n953 vn_p.n951 0.316
R2164 vn_p.n955 vn_p.n953 0.316
R2165 vn_p.n957 vn_p.n955 0.316
R2166 vn_p.n959 vn_p.n957 0.316
R2167 vn_p.n961 vn_p.n959 0.316
R2168 vn_p.n963 vn_p.n961 0.316
R2169 vn_p.n965 vn_p.n963 0.316
R2170 vn_p.n967 vn_p.n965 0.316
R2171 vn_p.n969 vn_p.n967 0.316
R2172 vn_p.n971 vn_p.n969 0.316
R2173 vn_p.n976 vn_p.n974 0.316
R2174 vn_p.n978 vn_p.n976 0.316
R2175 vn_p.n980 vn_p.n978 0.316
R2176 vn_p.n982 vn_p.n980 0.316
R2177 vn_p.n984 vn_p.n982 0.316
R2178 vn_p.n986 vn_p.n984 0.316
R2179 vn_p.n988 vn_p.n986 0.316
R2180 vn_p.n990 vn_p.n988 0.316
R2181 vn_p.n992 vn_p.n990 0.316
R2182 vn_p.n994 vn_p.n992 0.316
R2183 vn_p.n996 vn_p.n994 0.316
R2184 vn_p.n998 vn_p.n996 0.316
R2185 vn_p.n1000 vn_p.n998 0.316
R2186 vn_p.n1002 vn_p.n1000 0.316
R2187 vn_p.n1004 vn_p.n1002 0.316
R2188 vn_p.n1006 vn_p.n1004 0.316
R2189 vn_p.n1008 vn_p.n1006 0.316
R2190 vn_p.n1010 vn_p.n1008 0.316
R2191 vn_p.n1012 vn_p.n1010 0.316
R2192 vn_p.n1014 vn_p.n1012 0.316
R2193 vn_p.n1016 vn_p.n1014 0.316
R2194 vn_p.n1018 vn_p.n1016 0.316
R2195 vn_p.n1020 vn_p.n1018 0.316
R2196 vn_p.n1022 vn_p.n1020 0.316
R2197 vn_p.n1024 vn_p.n1022 0.316
R2198 vn_p.n1026 vn_p.n1024 0.316
R2199 vn_p.n1028 vn_p.n1026 0.316
R2200 vn_p.n1030 vn_p.n1028 0.316
R2201 vn_p.n1032 vn_p.n1030 0.316
R2202 vn_p.n1034 vn_p.n1032 0.316
R2203 vn_p.n1036 vn_p.n1034 0.316
R2204 vn_p.n1038 vn_p.n1036 0.316
R2205 vn_p.n1040 vn_p.n1038 0.316
R2206 vn_p.n1042 vn_p.n1040 0.316
R2207 vn_p.n1044 vn_p.n1042 0.316
R2208 vn_p.n1046 vn_p.n1044 0.316
R2209 vn_p.n1048 vn_p.n1046 0.316
R2210 vn_p.n1050 vn_p.n1048 0.316
R2211 vn_p.n1052 vn_p.n1050 0.316
R2212 vn_p.n1054 vn_p.n1052 0.316
R2213 vn_p.n1056 vn_p.n1054 0.316
R2214 vn_p.n1058 vn_p.n1056 0.316
R2215 vn_p.n1060 vn_p.n1058 0.316
R2216 vn_p.n1062 vn_p.n1060 0.316
R2217 vn_p.n1064 vn_p.n1062 0.316
R2218 vn_p.n1066 vn_p.n1064 0.316
R2219 vn_p.n1068 vn_p.n1066 0.316
R2220 vn_p.n1070 vn_p.n1068 0.316
R2221 vn_p.n1072 vn_p.n1070 0.316
R2222 vn_p.n1074 vn_p.n1072 0.316
R2223 vn_p.n1076 vn_p.n1074 0.316
R2224 vn_p.n1078 vn_p.n1076 0.316
R2225 vn_p.n1080 vn_p.n1078 0.316
R2226 vn_p.n1082 vn_p.n1080 0.316
R2227 vn_p.n1084 vn_p.n1082 0.316
R2228 vn_p.n1086 vn_p.n1084 0.316
R2229 vn_p.n1088 vn_p.n1086 0.316
R2230 vn_p.n1090 vn_p.n1088 0.316
R2231 vn_p.n1092 vn_p.n1090 0.316
R2232 vn_p.n1094 vn_p.n1092 0.316
R2233 vn_p.n1096 vn_p.n1094 0.316
R2234 vn_p.n1098 vn_p.n1096 0.316
R2235 vn_p.n1100 vn_p.n1098 0.316
R2236 vn_p.n1102 vn_p.n1100 0.316
R2237 vn_p.n1104 vn_p.n1102 0.316
R2238 vn_p.n1106 vn_p.n1104 0.316
R2239 vn_p.n1108 vn_p.n1106 0.316
R2240 vn_p.n1110 vn_p.n1108 0.316
R2241 vn_p.n1112 vn_p.n1110 0.316
R2242 vn_p.n1114 vn_p.n1112 0.316
R2243 vn_p.n1116 vn_p.n1114 0.316
R2244 vn_p.n1118 vn_p.n1116 0.316
R2245 vn_p.n1120 vn_p.n1118 0.316
R2246 vn_p.n1125 vn_p.n1123 0.316
R2247 vn_p.n1127 vn_p.n1125 0.316
R2248 vn_p.n1129 vn_p.n1127 0.316
R2249 vn_p.n1131 vn_p.n1129 0.316
R2250 vn_p.n1133 vn_p.n1131 0.316
R2251 vn_p.n1135 vn_p.n1133 0.316
R2252 vn_p.n1137 vn_p.n1135 0.316
R2253 vn_p.n1139 vn_p.n1137 0.316
R2254 vn_p.n1141 vn_p.n1139 0.316
R2255 vn_p.n1143 vn_p.n1141 0.316
R2256 vn_p.n1145 vn_p.n1143 0.316
R2257 vn_p.n1147 vn_p.n1145 0.316
R2258 vn_p.n1149 vn_p.n1147 0.316
R2259 vn_p.n1151 vn_p.n1149 0.316
R2260 vn_p.n1153 vn_p.n1151 0.316
R2261 vn_p.n1155 vn_p.n1153 0.316
R2262 vn_p.n1157 vn_p.n1155 0.316
R2263 vn_p.n1159 vn_p.n1157 0.316
R2264 vn_p.n1161 vn_p.n1159 0.316
R2265 vn_p.n1163 vn_p.n1161 0.316
R2266 vn_p.n1165 vn_p.n1163 0.316
R2267 vn_p.n1167 vn_p.n1165 0.316
R2268 vn_p.n1169 vn_p.n1167 0.316
R2269 vn_p.n1171 vn_p.n1169 0.316
R2270 vn_p.n1173 vn_p.n1171 0.316
R2271 vn_p.n1175 vn_p.n1173 0.316
R2272 vn_p.n1177 vn_p.n1175 0.316
R2273 vn_p.n1179 vn_p.n1177 0.316
R2274 vn_p.n1181 vn_p.n1179 0.316
R2275 vn_p.n1183 vn_p.n1181 0.316
R2276 vn_p.n1185 vn_p.n1183 0.316
R2277 vn_p.n1187 vn_p.n1185 0.316
R2278 vn_p.n1189 vn_p.n1187 0.316
R2279 vn_p.n1191 vn_p.n1189 0.316
R2280 vn_p.n1193 vn_p.n1191 0.316
R2281 vn_p.n1195 vn_p.n1193 0.316
R2282 vn_p.n1197 vn_p.n1195 0.316
R2283 vn_p.n1199 vn_p.n1197 0.316
R2284 vn_p.n1201 vn_p.n1199 0.316
R2285 vn_p.n1203 vn_p.n1201 0.316
R2286 vn_p.n1205 vn_p.n1203 0.316
R2287 vn_p.n1207 vn_p.n1205 0.316
R2288 vn_p.n1209 vn_p.n1207 0.316
R2289 vn_p.n1211 vn_p.n1209 0.316
R2290 vn_p.n1213 vn_p.n1211 0.316
R2291 vn_p.n1215 vn_p.n1213 0.316
R2292 vn_p.n1217 vn_p.n1215 0.316
R2293 vn_p.n1219 vn_p.n1217 0.316
R2294 vn_p.n1221 vn_p.n1219 0.316
R2295 vn_p.n1223 vn_p.n1221 0.316
R2296 vn_p.n1225 vn_p.n1223 0.316
R2297 vn_p.n1227 vn_p.n1225 0.316
R2298 vn_p.n1229 vn_p.n1227 0.316
R2299 vn_p.n1231 vn_p.n1229 0.316
R2300 vn_p.n1233 vn_p.n1231 0.316
R2301 vn_p.n1235 vn_p.n1233 0.316
R2302 vn_p.n1237 vn_p.n1235 0.316
R2303 vn_p.n1239 vn_p.n1237 0.316
R2304 vn_p.n1241 vn_p.n1239 0.316
R2305 vn_p.n1243 vn_p.n1241 0.316
R2306 vn_p.n1245 vn_p.n1243 0.316
R2307 vn_p.n1247 vn_p.n1245 0.316
R2308 vn_p.n1249 vn_p.n1247 0.316
R2309 vn_p.n1251 vn_p.n1249 0.316
R2310 vn_p.n1253 vn_p.n1251 0.316
R2311 vn_p.n1255 vn_p.n1253 0.316
R2312 vn_p.n1257 vn_p.n1255 0.316
R2313 vn_p.n1259 vn_p.n1257 0.316
R2314 vn_p.n1261 vn_p.n1259 0.316
R2315 vn_p.n1263 vn_p.n1261 0.316
R2316 vn_p.n1265 vn_p.n1263 0.316
R2317 vn_p.n1267 vn_p.n1265 0.316
R2318 vn_p.n1269 vn_p.n1267 0.316
R2319 vn_p.n1274 vn_p.n1272 0.316
R2320 vn_p.n1276 vn_p.n1274 0.316
R2321 vn_p.n1278 vn_p.n1276 0.316
R2322 vn_p.n1280 vn_p.n1278 0.316
R2323 vn_p.n1282 vn_p.n1280 0.316
R2324 vn_p.n1284 vn_p.n1282 0.316
R2325 vn_p.n1286 vn_p.n1284 0.316
R2326 vn_p.n1288 vn_p.n1286 0.316
R2327 vn_p.n1290 vn_p.n1288 0.316
R2328 vn_p.n1292 vn_p.n1290 0.316
R2329 vn_p.n1294 vn_p.n1292 0.316
R2330 vn_p.n1296 vn_p.n1294 0.316
R2331 vn_p.n1298 vn_p.n1296 0.316
R2332 vn_p.n1300 vn_p.n1298 0.316
R2333 vn_p.n1302 vn_p.n1300 0.316
R2334 vn_p.n1304 vn_p.n1302 0.316
R2335 vn_p.n1306 vn_p.n1304 0.316
R2336 vn_p.n1308 vn_p.n1306 0.316
R2337 vn_p.n1310 vn_p.n1308 0.316
R2338 vn_p.n1312 vn_p.n1310 0.316
R2339 vn_p.n1314 vn_p.n1312 0.316
R2340 vn_p.n1316 vn_p.n1314 0.316
R2341 vn_p.n1318 vn_p.n1316 0.316
R2342 vn_p.n1320 vn_p.n1318 0.316
R2343 vn_p.n1322 vn_p.n1320 0.316
R2344 vn_p.n1324 vn_p.n1322 0.316
R2345 vn_p.n1326 vn_p.n1324 0.316
R2346 vn_p.n1328 vn_p.n1326 0.316
R2347 vn_p.n1330 vn_p.n1328 0.316
R2348 vn_p.n1332 vn_p.n1330 0.316
R2349 vn_p.n1334 vn_p.n1332 0.316
R2350 vn_p.n1336 vn_p.n1334 0.316
R2351 vn_p.n1338 vn_p.n1336 0.316
R2352 vn_p.n1340 vn_p.n1338 0.316
R2353 vn_p.n1342 vn_p.n1340 0.316
R2354 vn_p.n1344 vn_p.n1342 0.316
R2355 vn_p.n1346 vn_p.n1344 0.316
R2356 vn_p.n1348 vn_p.n1346 0.316
R2357 vn_p.n1350 vn_p.n1348 0.316
R2358 vn_p.n1352 vn_p.n1350 0.316
R2359 vn_p.n1354 vn_p.n1352 0.316
R2360 vn_p.n1356 vn_p.n1354 0.316
R2361 vn_p.n1358 vn_p.n1356 0.316
R2362 vn_p.n1360 vn_p.n1358 0.316
R2363 vn_p.n1362 vn_p.n1360 0.316
R2364 vn_p.n1364 vn_p.n1362 0.316
R2365 vn_p.n1366 vn_p.n1364 0.316
R2366 vn_p.n1368 vn_p.n1366 0.316
R2367 vn_p.n1370 vn_p.n1368 0.316
R2368 vn_p.n1372 vn_p.n1370 0.316
R2369 vn_p.n1374 vn_p.n1372 0.316
R2370 vn_p.n1376 vn_p.n1374 0.316
R2371 vn_p.n1378 vn_p.n1376 0.316
R2372 vn_p.n1380 vn_p.n1378 0.316
R2373 vn_p.n1382 vn_p.n1380 0.316
R2374 vn_p.n1384 vn_p.n1382 0.316
R2375 vn_p.n1386 vn_p.n1384 0.316
R2376 vn_p.n1388 vn_p.n1386 0.316
R2377 vn_p.n1390 vn_p.n1388 0.316
R2378 vn_p.n1392 vn_p.n1390 0.316
R2379 vn_p.n1394 vn_p.n1392 0.316
R2380 vn_p.n1396 vn_p.n1394 0.316
R2381 vn_p.n1398 vn_p.n1396 0.316
R2382 vn_p.n1400 vn_p.n1398 0.316
R2383 vn_p.n1402 vn_p.n1400 0.316
R2384 vn_p.n1404 vn_p.n1402 0.316
R2385 vn_p.n1406 vn_p.n1404 0.316
R2386 vn_p.n1408 vn_p.n1406 0.316
R2387 vn_p.n1410 vn_p.n1408 0.316
R2388 vn_p.n1412 vn_p.n1410 0.316
R2389 vn_p.n1414 vn_p.n1412 0.316
R2390 vn_p.n1416 vn_p.n1414 0.316
R2391 vn_p.n1418 vn_p.n1416 0.316
R2392 vn_p.n745 vn_p.n744 0.149
R2393 vn_p.n746 vn_p.n745 0.149
R2394 vn_p.n747 vn_p.n746 0.149
R2395 vn_p.n1496 vn_p.n1495 0.149
R2396 vn_p.n1494 vn_p.n1493 0.149
R2397 vn_p.n748 vn_p.n747 0.141
R2398 vn_p.n1497 vn_p.n1496 0.141
R2399 vn_p.n744 vn_p.n669 0.134
R2400 vn_p.n746 vn_p.n371 0.134
R2401 vn_p.n1496 vn_p.n971 0.134
R2402 vn_p.n1494 vn_p.n1269 0.134
R2403 vn_p.n1495 vn_p 0.121
R2404 vn_p.n669 vn_p.n668 0.04
R2405 vn_p.n667 vn_p.n666 0.04
R2406 vn_p.n665 vn_p.n664 0.04
R2407 vn_p.n663 vn_p.n662 0.04
R2408 vn_p.n661 vn_p.n660 0.04
R2409 vn_p.n659 vn_p.n658 0.04
R2410 vn_p.n657 vn_p.n656 0.04
R2411 vn_p.n655 vn_p.n654 0.04
R2412 vn_p.n653 vn_p.n652 0.04
R2413 vn_p.n651 vn_p.n650 0.04
R2414 vn_p.n649 vn_p.n648 0.04
R2415 vn_p.n647 vn_p.n646 0.04
R2416 vn_p.n645 vn_p.n644 0.04
R2417 vn_p.n643 vn_p.n642 0.04
R2418 vn_p.n641 vn_p.n640 0.04
R2419 vn_p.n639 vn_p.n638 0.04
R2420 vn_p.n637 vn_p.n636 0.04
R2421 vn_p.n635 vn_p.n634 0.04
R2422 vn_p.n633 vn_p.n632 0.04
R2423 vn_p.n631 vn_p.n630 0.04
R2424 vn_p.n629 vn_p.n628 0.04
R2425 vn_p.n627 vn_p.n626 0.04
R2426 vn_p.n625 vn_p.n624 0.04
R2427 vn_p.n623 vn_p.n622 0.04
R2428 vn_p.n621 vn_p.n620 0.04
R2429 vn_p.n619 vn_p.n618 0.04
R2430 vn_p.n617 vn_p.n616 0.04
R2431 vn_p.n615 vn_p.n614 0.04
R2432 vn_p.n613 vn_p.n612 0.04
R2433 vn_p.n611 vn_p.n610 0.04
R2434 vn_p.n609 vn_p.n608 0.04
R2435 vn_p.n607 vn_p.n606 0.04
R2436 vn_p.n605 vn_p.n604 0.04
R2437 vn_p.n603 vn_p.n602 0.04
R2438 vn_p.n601 vn_p.n600 0.04
R2439 vn_p.n599 vn_p.n598 0.04
R2440 vn_p.n597 vn_p.n596 0.04
R2441 vn_p.n595 vn_p.n594 0.04
R2442 vn_p.n593 vn_p.n592 0.04
R2443 vn_p.n591 vn_p.n590 0.04
R2444 vn_p.n589 vn_p.n588 0.04
R2445 vn_p.n587 vn_p.n586 0.04
R2446 vn_p.n585 vn_p.n584 0.04
R2447 vn_p.n583 vn_p.n582 0.04
R2448 vn_p.n581 vn_p.n580 0.04
R2449 vn_p.n579 vn_p.n578 0.04
R2450 vn_p.n577 vn_p.n576 0.04
R2451 vn_p.n575 vn_p.n574 0.04
R2452 vn_p.n573 vn_p.n572 0.04
R2453 vn_p.n571 vn_p.n570 0.04
R2454 vn_p.n569 vn_p.n568 0.04
R2455 vn_p.n567 vn_p.n566 0.04
R2456 vn_p.n565 vn_p.n564 0.04
R2457 vn_p.n563 vn_p.n562 0.04
R2458 vn_p.n561 vn_p.n560 0.04
R2459 vn_p.n559 vn_p.n558 0.04
R2460 vn_p.n557 vn_p.n556 0.04
R2461 vn_p.n555 vn_p.n554 0.04
R2462 vn_p.n553 vn_p.n552 0.04
R2463 vn_p.n551 vn_p.n550 0.04
R2464 vn_p.n549 vn_p.n548 0.04
R2465 vn_p.n547 vn_p.n546 0.04
R2466 vn_p.n545 vn_p.n544 0.04
R2467 vn_p.n543 vn_p.n542 0.04
R2468 vn_p.n541 vn_p.n540 0.04
R2469 vn_p.n539 vn_p.n538 0.04
R2470 vn_p.n537 vn_p.n536 0.04
R2471 vn_p.n535 vn_p.n534 0.04
R2472 vn_p.n533 vn_p.n532 0.04
R2473 vn_p.n531 vn_p.n530 0.04
R2474 vn_p.n529 vn_p.n528 0.04
R2475 vn_p.n527 vn_p.n526 0.04
R2476 vn_p.n525 vn_p.n524 0.04
R2477 vn_p.n523 vn_p.n522 0.04
R2478 vn_p.n520 vn_p.n519 0.04
R2479 vn_p.n518 vn_p.n517 0.04
R2480 vn_p.n516 vn_p.n515 0.04
R2481 vn_p.n514 vn_p.n513 0.04
R2482 vn_p.n512 vn_p.n511 0.04
R2483 vn_p.n510 vn_p.n509 0.04
R2484 vn_p.n508 vn_p.n507 0.04
R2485 vn_p.n506 vn_p.n505 0.04
R2486 vn_p.n504 vn_p.n503 0.04
R2487 vn_p.n502 vn_p.n501 0.04
R2488 vn_p.n500 vn_p.n499 0.04
R2489 vn_p.n498 vn_p.n497 0.04
R2490 vn_p.n496 vn_p.n495 0.04
R2491 vn_p.n494 vn_p.n493 0.04
R2492 vn_p.n492 vn_p.n491 0.04
R2493 vn_p.n490 vn_p.n489 0.04
R2494 vn_p.n488 vn_p.n487 0.04
R2495 vn_p.n486 vn_p.n485 0.04
R2496 vn_p.n484 vn_p.n483 0.04
R2497 vn_p.n482 vn_p.n481 0.04
R2498 vn_p.n480 vn_p.n479 0.04
R2499 vn_p.n478 vn_p.n477 0.04
R2500 vn_p.n476 vn_p.n475 0.04
R2501 vn_p.n474 vn_p.n473 0.04
R2502 vn_p.n472 vn_p.n471 0.04
R2503 vn_p.n470 vn_p.n469 0.04
R2504 vn_p.n468 vn_p.n467 0.04
R2505 vn_p.n466 vn_p.n465 0.04
R2506 vn_p.n464 vn_p.n463 0.04
R2507 vn_p.n462 vn_p.n461 0.04
R2508 vn_p.n460 vn_p.n459 0.04
R2509 vn_p.n458 vn_p.n457 0.04
R2510 vn_p.n456 vn_p.n455 0.04
R2511 vn_p.n454 vn_p.n453 0.04
R2512 vn_p.n452 vn_p.n451 0.04
R2513 vn_p.n450 vn_p.n449 0.04
R2514 vn_p.n448 vn_p.n447 0.04
R2515 vn_p.n446 vn_p.n445 0.04
R2516 vn_p.n444 vn_p.n443 0.04
R2517 vn_p.n442 vn_p.n441 0.04
R2518 vn_p.n440 vn_p.n439 0.04
R2519 vn_p.n438 vn_p.n437 0.04
R2520 vn_p.n436 vn_p.n435 0.04
R2521 vn_p.n434 vn_p.n433 0.04
R2522 vn_p.n432 vn_p.n431 0.04
R2523 vn_p.n430 vn_p.n429 0.04
R2524 vn_p.n428 vn_p.n427 0.04
R2525 vn_p.n426 vn_p.n425 0.04
R2526 vn_p.n424 vn_p.n423 0.04
R2527 vn_p.n422 vn_p.n421 0.04
R2528 vn_p.n420 vn_p.n419 0.04
R2529 vn_p.n418 vn_p.n417 0.04
R2530 vn_p.n416 vn_p.n415 0.04
R2531 vn_p.n414 vn_p.n413 0.04
R2532 vn_p.n412 vn_p.n411 0.04
R2533 vn_p.n410 vn_p.n409 0.04
R2534 vn_p.n408 vn_p.n407 0.04
R2535 vn_p.n406 vn_p.n405 0.04
R2536 vn_p.n404 vn_p.n403 0.04
R2537 vn_p.n402 vn_p.n401 0.04
R2538 vn_p.n400 vn_p.n399 0.04
R2539 vn_p.n398 vn_p.n397 0.04
R2540 vn_p.n396 vn_p.n395 0.04
R2541 vn_p.n394 vn_p.n393 0.04
R2542 vn_p.n392 vn_p.n391 0.04
R2543 vn_p.n390 vn_p.n389 0.04
R2544 vn_p.n388 vn_p.n387 0.04
R2545 vn_p.n386 vn_p.n385 0.04
R2546 vn_p.n384 vn_p.n383 0.04
R2547 vn_p.n382 vn_p.n381 0.04
R2548 vn_p.n380 vn_p.n379 0.04
R2549 vn_p.n378 vn_p.n377 0.04
R2550 vn_p.n376 vn_p.n375 0.04
R2551 vn_p.n374 vn_p.n373 0.04
R2552 vn_p.n371 vn_p.n370 0.04
R2553 vn_p.n369 vn_p.n368 0.04
R2554 vn_p.n367 vn_p.n366 0.04
R2555 vn_p.n365 vn_p.n364 0.04
R2556 vn_p.n363 vn_p.n362 0.04
R2557 vn_p.n361 vn_p.n360 0.04
R2558 vn_p.n359 vn_p.n358 0.04
R2559 vn_p.n357 vn_p.n356 0.04
R2560 vn_p.n355 vn_p.n354 0.04
R2561 vn_p.n353 vn_p.n352 0.04
R2562 vn_p.n351 vn_p.n350 0.04
R2563 vn_p.n349 vn_p.n348 0.04
R2564 vn_p.n347 vn_p.n346 0.04
R2565 vn_p.n345 vn_p.n344 0.04
R2566 vn_p.n343 vn_p.n342 0.04
R2567 vn_p.n341 vn_p.n340 0.04
R2568 vn_p.n339 vn_p.n338 0.04
R2569 vn_p.n337 vn_p.n336 0.04
R2570 vn_p.n335 vn_p.n334 0.04
R2571 vn_p.n333 vn_p.n332 0.04
R2572 vn_p.n331 vn_p.n330 0.04
R2573 vn_p.n329 vn_p.n328 0.04
R2574 vn_p.n327 vn_p.n326 0.04
R2575 vn_p.n325 vn_p.n324 0.04
R2576 vn_p.n323 vn_p.n322 0.04
R2577 vn_p.n321 vn_p.n320 0.04
R2578 vn_p.n319 vn_p.n318 0.04
R2579 vn_p.n317 vn_p.n316 0.04
R2580 vn_p.n315 vn_p.n314 0.04
R2581 vn_p.n313 vn_p.n312 0.04
R2582 vn_p.n311 vn_p.n310 0.04
R2583 vn_p.n309 vn_p.n308 0.04
R2584 vn_p.n307 vn_p.n306 0.04
R2585 vn_p.n305 vn_p.n304 0.04
R2586 vn_p.n303 vn_p.n302 0.04
R2587 vn_p.n301 vn_p.n300 0.04
R2588 vn_p.n299 vn_p.n298 0.04
R2589 vn_p.n297 vn_p.n296 0.04
R2590 vn_p.n295 vn_p.n294 0.04
R2591 vn_p.n293 vn_p.n292 0.04
R2592 vn_p.n291 vn_p.n290 0.04
R2593 vn_p.n289 vn_p.n288 0.04
R2594 vn_p.n287 vn_p.n286 0.04
R2595 vn_p.n285 vn_p.n284 0.04
R2596 vn_p.n283 vn_p.n282 0.04
R2597 vn_p.n281 vn_p.n280 0.04
R2598 vn_p.n279 vn_p.n278 0.04
R2599 vn_p.n277 vn_p.n276 0.04
R2600 vn_p.n275 vn_p.n274 0.04
R2601 vn_p.n273 vn_p.n272 0.04
R2602 vn_p.n271 vn_p.n270 0.04
R2603 vn_p.n269 vn_p.n268 0.04
R2604 vn_p.n267 vn_p.n266 0.04
R2605 vn_p.n265 vn_p.n264 0.04
R2606 vn_p.n263 vn_p.n262 0.04
R2607 vn_p.n261 vn_p.n260 0.04
R2608 vn_p.n259 vn_p.n258 0.04
R2609 vn_p.n257 vn_p.n256 0.04
R2610 vn_p.n255 vn_p.n254 0.04
R2611 vn_p.n253 vn_p.n252 0.04
R2612 vn_p.n251 vn_p.n250 0.04
R2613 vn_p.n249 vn_p.n248 0.04
R2614 vn_p.n247 vn_p.n246 0.04
R2615 vn_p.n245 vn_p.n244 0.04
R2616 vn_p.n243 vn_p.n242 0.04
R2617 vn_p.n241 vn_p.n240 0.04
R2618 vn_p.n239 vn_p.n238 0.04
R2619 vn_p.n237 vn_p.n236 0.04
R2620 vn_p.n235 vn_p.n234 0.04
R2621 vn_p.n233 vn_p.n232 0.04
R2622 vn_p.n231 vn_p.n230 0.04
R2623 vn_p.n229 vn_p.n228 0.04
R2624 vn_p.n227 vn_p.n226 0.04
R2625 vn_p.n225 vn_p.n224 0.04
R2626 vn_p.n222 vn_p.n221 0.04
R2627 vn_p.n220 vn_p.n219 0.04
R2628 vn_p.n218 vn_p.n217 0.04
R2629 vn_p.n216 vn_p.n215 0.04
R2630 vn_p.n214 vn_p.n213 0.04
R2631 vn_p.n212 vn_p.n211 0.04
R2632 vn_p.n210 vn_p.n209 0.04
R2633 vn_p.n208 vn_p.n207 0.04
R2634 vn_p.n206 vn_p.n205 0.04
R2635 vn_p.n204 vn_p.n203 0.04
R2636 vn_p.n202 vn_p.n201 0.04
R2637 vn_p.n200 vn_p.n199 0.04
R2638 vn_p.n198 vn_p.n197 0.04
R2639 vn_p.n196 vn_p.n195 0.04
R2640 vn_p.n194 vn_p.n193 0.04
R2641 vn_p.n192 vn_p.n191 0.04
R2642 vn_p.n190 vn_p.n189 0.04
R2643 vn_p.n188 vn_p.n187 0.04
R2644 vn_p.n186 vn_p.n185 0.04
R2645 vn_p.n184 vn_p.n183 0.04
R2646 vn_p.n182 vn_p.n181 0.04
R2647 vn_p.n180 vn_p.n179 0.04
R2648 vn_p.n178 vn_p.n177 0.04
R2649 vn_p.n176 vn_p.n175 0.04
R2650 vn_p.n174 vn_p.n173 0.04
R2651 vn_p.n172 vn_p.n171 0.04
R2652 vn_p.n170 vn_p.n169 0.04
R2653 vn_p.n168 vn_p.n167 0.04
R2654 vn_p.n166 vn_p.n165 0.04
R2655 vn_p.n164 vn_p.n163 0.04
R2656 vn_p.n162 vn_p.n161 0.04
R2657 vn_p.n160 vn_p.n159 0.04
R2658 vn_p.n158 vn_p.n157 0.04
R2659 vn_p.n156 vn_p.n155 0.04
R2660 vn_p.n154 vn_p.n153 0.04
R2661 vn_p.n152 vn_p.n151 0.04
R2662 vn_p.n150 vn_p.n149 0.04
R2663 vn_p.n148 vn_p.n147 0.04
R2664 vn_p.n146 vn_p.n145 0.04
R2665 vn_p.n144 vn_p.n143 0.04
R2666 vn_p.n142 vn_p.n141 0.04
R2667 vn_p.n140 vn_p.n139 0.04
R2668 vn_p.n138 vn_p.n137 0.04
R2669 vn_p.n136 vn_p.n135 0.04
R2670 vn_p.n134 vn_p.n133 0.04
R2671 vn_p.n132 vn_p.n131 0.04
R2672 vn_p.n130 vn_p.n129 0.04
R2673 vn_p.n128 vn_p.n127 0.04
R2674 vn_p.n126 vn_p.n125 0.04
R2675 vn_p.n124 vn_p.n123 0.04
R2676 vn_p.n122 vn_p.n121 0.04
R2677 vn_p.n120 vn_p.n119 0.04
R2678 vn_p.n118 vn_p.n117 0.04
R2679 vn_p.n116 vn_p.n115 0.04
R2680 vn_p.n114 vn_p.n113 0.04
R2681 vn_p.n112 vn_p.n111 0.04
R2682 vn_p.n110 vn_p.n109 0.04
R2683 vn_p.n108 vn_p.n107 0.04
R2684 vn_p.n106 vn_p.n105 0.04
R2685 vn_p.n104 vn_p.n103 0.04
R2686 vn_p.n102 vn_p.n101 0.04
R2687 vn_p.n100 vn_p.n99 0.04
R2688 vn_p.n98 vn_p.n97 0.04
R2689 vn_p.n96 vn_p.n95 0.04
R2690 vn_p.n94 vn_p.n93 0.04
R2691 vn_p.n92 vn_p.n91 0.04
R2692 vn_p.n90 vn_p.n89 0.04
R2693 vn_p.n88 vn_p.n87 0.04
R2694 vn_p.n86 vn_p.n85 0.04
R2695 vn_p.n84 vn_p.n83 0.04
R2696 vn_p.n82 vn_p.n81 0.04
R2697 vn_p.n80 vn_p.n79 0.04
R2698 vn_p.n78 vn_p.n77 0.04
R2699 vn_p.n76 vn_p.n75 0.04
R2700 vn_p.n971 vn_p.n970 0.04
R2701 vn_p.n969 vn_p.n968 0.04
R2702 vn_p.n967 vn_p.n966 0.04
R2703 vn_p.n965 vn_p.n964 0.04
R2704 vn_p.n963 vn_p.n962 0.04
R2705 vn_p.n961 vn_p.n960 0.04
R2706 vn_p.n959 vn_p.n958 0.04
R2707 vn_p.n957 vn_p.n956 0.04
R2708 vn_p.n955 vn_p.n954 0.04
R2709 vn_p.n953 vn_p.n952 0.04
R2710 vn_p.n951 vn_p.n950 0.04
R2711 vn_p.n949 vn_p.n948 0.04
R2712 vn_p.n947 vn_p.n946 0.04
R2713 vn_p.n945 vn_p.n944 0.04
R2714 vn_p.n943 vn_p.n942 0.04
R2715 vn_p.n941 vn_p.n940 0.04
R2716 vn_p.n939 vn_p.n938 0.04
R2717 vn_p.n937 vn_p.n936 0.04
R2718 vn_p.n935 vn_p.n934 0.04
R2719 vn_p.n933 vn_p.n932 0.04
R2720 vn_p.n931 vn_p.n930 0.04
R2721 vn_p.n929 vn_p.n928 0.04
R2722 vn_p.n927 vn_p.n926 0.04
R2723 vn_p.n925 vn_p.n924 0.04
R2724 vn_p.n923 vn_p.n922 0.04
R2725 vn_p.n921 vn_p.n920 0.04
R2726 vn_p.n919 vn_p.n918 0.04
R2727 vn_p.n917 vn_p.n916 0.04
R2728 vn_p.n915 vn_p.n914 0.04
R2729 vn_p.n913 vn_p.n912 0.04
R2730 vn_p.n911 vn_p.n910 0.04
R2731 vn_p.n909 vn_p.n908 0.04
R2732 vn_p.n907 vn_p.n906 0.04
R2733 vn_p.n905 vn_p.n904 0.04
R2734 vn_p.n903 vn_p.n902 0.04
R2735 vn_p.n901 vn_p.n900 0.04
R2736 vn_p.n899 vn_p.n898 0.04
R2737 vn_p.n897 vn_p.n896 0.04
R2738 vn_p.n895 vn_p.n894 0.04
R2739 vn_p.n893 vn_p.n892 0.04
R2740 vn_p.n891 vn_p.n890 0.04
R2741 vn_p.n889 vn_p.n888 0.04
R2742 vn_p.n887 vn_p.n886 0.04
R2743 vn_p.n885 vn_p.n884 0.04
R2744 vn_p.n883 vn_p.n882 0.04
R2745 vn_p.n881 vn_p.n880 0.04
R2746 vn_p.n879 vn_p.n878 0.04
R2747 vn_p.n877 vn_p.n876 0.04
R2748 vn_p.n875 vn_p.n874 0.04
R2749 vn_p.n873 vn_p.n872 0.04
R2750 vn_p.n871 vn_p.n870 0.04
R2751 vn_p.n869 vn_p.n868 0.04
R2752 vn_p.n867 vn_p.n866 0.04
R2753 vn_p.n865 vn_p.n864 0.04
R2754 vn_p.n863 vn_p.n862 0.04
R2755 vn_p.n861 vn_p.n860 0.04
R2756 vn_p.n859 vn_p.n858 0.04
R2757 vn_p.n857 vn_p.n856 0.04
R2758 vn_p.n855 vn_p.n854 0.04
R2759 vn_p.n853 vn_p.n852 0.04
R2760 vn_p.n851 vn_p.n850 0.04
R2761 vn_p.n849 vn_p.n848 0.04
R2762 vn_p.n847 vn_p.n846 0.04
R2763 vn_p.n845 vn_p.n844 0.04
R2764 vn_p.n843 vn_p.n842 0.04
R2765 vn_p.n841 vn_p.n840 0.04
R2766 vn_p.n839 vn_p.n838 0.04
R2767 vn_p.n837 vn_p.n836 0.04
R2768 vn_p.n835 vn_p.n834 0.04
R2769 vn_p.n833 vn_p.n832 0.04
R2770 vn_p.n831 vn_p.n830 0.04
R2771 vn_p.n829 vn_p.n828 0.04
R2772 vn_p.n827 vn_p.n826 0.04
R2773 vn_p.n825 vn_p.n824 0.04
R2774 vn_p.n1120 vn_p.n1119 0.04
R2775 vn_p.n1118 vn_p.n1117 0.04
R2776 vn_p.n1116 vn_p.n1115 0.04
R2777 vn_p.n1114 vn_p.n1113 0.04
R2778 vn_p.n1112 vn_p.n1111 0.04
R2779 vn_p.n1110 vn_p.n1109 0.04
R2780 vn_p.n1108 vn_p.n1107 0.04
R2781 vn_p.n1106 vn_p.n1105 0.04
R2782 vn_p.n1104 vn_p.n1103 0.04
R2783 vn_p.n1102 vn_p.n1101 0.04
R2784 vn_p.n1100 vn_p.n1099 0.04
R2785 vn_p.n1098 vn_p.n1097 0.04
R2786 vn_p.n1096 vn_p.n1095 0.04
R2787 vn_p.n1094 vn_p.n1093 0.04
R2788 vn_p.n1092 vn_p.n1091 0.04
R2789 vn_p.n1090 vn_p.n1089 0.04
R2790 vn_p.n1088 vn_p.n1087 0.04
R2791 vn_p.n1086 vn_p.n1085 0.04
R2792 vn_p.n1084 vn_p.n1083 0.04
R2793 vn_p.n1082 vn_p.n1081 0.04
R2794 vn_p.n1080 vn_p.n1079 0.04
R2795 vn_p.n1078 vn_p.n1077 0.04
R2796 vn_p.n1076 vn_p.n1075 0.04
R2797 vn_p.n1074 vn_p.n1073 0.04
R2798 vn_p.n1072 vn_p.n1071 0.04
R2799 vn_p.n1070 vn_p.n1069 0.04
R2800 vn_p.n1068 vn_p.n1067 0.04
R2801 vn_p.n1066 vn_p.n1065 0.04
R2802 vn_p.n1064 vn_p.n1063 0.04
R2803 vn_p.n1062 vn_p.n1061 0.04
R2804 vn_p.n1060 vn_p.n1059 0.04
R2805 vn_p.n1058 vn_p.n1057 0.04
R2806 vn_p.n1056 vn_p.n1055 0.04
R2807 vn_p.n1054 vn_p.n1053 0.04
R2808 vn_p.n1052 vn_p.n1051 0.04
R2809 vn_p.n1050 vn_p.n1049 0.04
R2810 vn_p.n1048 vn_p.n1047 0.04
R2811 vn_p.n1046 vn_p.n1045 0.04
R2812 vn_p.n1044 vn_p.n1043 0.04
R2813 vn_p.n1042 vn_p.n1041 0.04
R2814 vn_p.n1040 vn_p.n1039 0.04
R2815 vn_p.n1038 vn_p.n1037 0.04
R2816 vn_p.n1036 vn_p.n1035 0.04
R2817 vn_p.n1034 vn_p.n1033 0.04
R2818 vn_p.n1032 vn_p.n1031 0.04
R2819 vn_p.n1030 vn_p.n1029 0.04
R2820 vn_p.n1028 vn_p.n1027 0.04
R2821 vn_p.n1026 vn_p.n1025 0.04
R2822 vn_p.n1024 vn_p.n1023 0.04
R2823 vn_p.n1022 vn_p.n1021 0.04
R2824 vn_p.n1020 vn_p.n1019 0.04
R2825 vn_p.n1018 vn_p.n1017 0.04
R2826 vn_p.n1016 vn_p.n1015 0.04
R2827 vn_p.n1014 vn_p.n1013 0.04
R2828 vn_p.n1012 vn_p.n1011 0.04
R2829 vn_p.n1010 vn_p.n1009 0.04
R2830 vn_p.n1008 vn_p.n1007 0.04
R2831 vn_p.n1006 vn_p.n1005 0.04
R2832 vn_p.n1004 vn_p.n1003 0.04
R2833 vn_p.n1002 vn_p.n1001 0.04
R2834 vn_p.n1000 vn_p.n999 0.04
R2835 vn_p.n998 vn_p.n997 0.04
R2836 vn_p.n996 vn_p.n995 0.04
R2837 vn_p.n994 vn_p.n993 0.04
R2838 vn_p.n992 vn_p.n991 0.04
R2839 vn_p.n990 vn_p.n989 0.04
R2840 vn_p.n988 vn_p.n987 0.04
R2841 vn_p.n986 vn_p.n985 0.04
R2842 vn_p.n984 vn_p.n983 0.04
R2843 vn_p.n982 vn_p.n981 0.04
R2844 vn_p.n980 vn_p.n979 0.04
R2845 vn_p.n978 vn_p.n977 0.04
R2846 vn_p.n976 vn_p.n975 0.04
R2847 vn_p.n974 vn_p.n973 0.04
R2848 vn_p.n1269 vn_p.n1268 0.04
R2849 vn_p.n1267 vn_p.n1266 0.04
R2850 vn_p.n1265 vn_p.n1264 0.04
R2851 vn_p.n1263 vn_p.n1262 0.04
R2852 vn_p.n1261 vn_p.n1260 0.04
R2853 vn_p.n1259 vn_p.n1258 0.04
R2854 vn_p.n1257 vn_p.n1256 0.04
R2855 vn_p.n1255 vn_p.n1254 0.04
R2856 vn_p.n1253 vn_p.n1252 0.04
R2857 vn_p.n1251 vn_p.n1250 0.04
R2858 vn_p.n1249 vn_p.n1248 0.04
R2859 vn_p.n1247 vn_p.n1246 0.04
R2860 vn_p.n1245 vn_p.n1244 0.04
R2861 vn_p.n1243 vn_p.n1242 0.04
R2862 vn_p.n1241 vn_p.n1240 0.04
R2863 vn_p.n1239 vn_p.n1238 0.04
R2864 vn_p.n1237 vn_p.n1236 0.04
R2865 vn_p.n1235 vn_p.n1234 0.04
R2866 vn_p.n1233 vn_p.n1232 0.04
R2867 vn_p.n1231 vn_p.n1230 0.04
R2868 vn_p.n1229 vn_p.n1228 0.04
R2869 vn_p.n1227 vn_p.n1226 0.04
R2870 vn_p.n1225 vn_p.n1224 0.04
R2871 vn_p.n1223 vn_p.n1222 0.04
R2872 vn_p.n1221 vn_p.n1220 0.04
R2873 vn_p.n1219 vn_p.n1218 0.04
R2874 vn_p.n1217 vn_p.n1216 0.04
R2875 vn_p.n1215 vn_p.n1214 0.04
R2876 vn_p.n1213 vn_p.n1212 0.04
R2877 vn_p.n1211 vn_p.n1210 0.04
R2878 vn_p.n1209 vn_p.n1208 0.04
R2879 vn_p.n1207 vn_p.n1206 0.04
R2880 vn_p.n1205 vn_p.n1204 0.04
R2881 vn_p.n1203 vn_p.n1202 0.04
R2882 vn_p.n1201 vn_p.n1200 0.04
R2883 vn_p.n1199 vn_p.n1198 0.04
R2884 vn_p.n1197 vn_p.n1196 0.04
R2885 vn_p.n1195 vn_p.n1194 0.04
R2886 vn_p.n1193 vn_p.n1192 0.04
R2887 vn_p.n1191 vn_p.n1190 0.04
R2888 vn_p.n1189 vn_p.n1188 0.04
R2889 vn_p.n1187 vn_p.n1186 0.04
R2890 vn_p.n1185 vn_p.n1184 0.04
R2891 vn_p.n1183 vn_p.n1182 0.04
R2892 vn_p.n1181 vn_p.n1180 0.04
R2893 vn_p.n1179 vn_p.n1178 0.04
R2894 vn_p.n1177 vn_p.n1176 0.04
R2895 vn_p.n1175 vn_p.n1174 0.04
R2896 vn_p.n1173 vn_p.n1172 0.04
R2897 vn_p.n1171 vn_p.n1170 0.04
R2898 vn_p.n1169 vn_p.n1168 0.04
R2899 vn_p.n1167 vn_p.n1166 0.04
R2900 vn_p.n1165 vn_p.n1164 0.04
R2901 vn_p.n1163 vn_p.n1162 0.04
R2902 vn_p.n1161 vn_p.n1160 0.04
R2903 vn_p.n1159 vn_p.n1158 0.04
R2904 vn_p.n1157 vn_p.n1156 0.04
R2905 vn_p.n1155 vn_p.n1154 0.04
R2906 vn_p.n1153 vn_p.n1152 0.04
R2907 vn_p.n1151 vn_p.n1150 0.04
R2908 vn_p.n1149 vn_p.n1148 0.04
R2909 vn_p.n1147 vn_p.n1146 0.04
R2910 vn_p.n1145 vn_p.n1144 0.04
R2911 vn_p.n1143 vn_p.n1142 0.04
R2912 vn_p.n1141 vn_p.n1140 0.04
R2913 vn_p.n1139 vn_p.n1138 0.04
R2914 vn_p.n1137 vn_p.n1136 0.04
R2915 vn_p.n1135 vn_p.n1134 0.04
R2916 vn_p.n1133 vn_p.n1132 0.04
R2917 vn_p.n1131 vn_p.n1130 0.04
R2918 vn_p.n1129 vn_p.n1128 0.04
R2919 vn_p.n1127 vn_p.n1126 0.04
R2920 vn_p.n1125 vn_p.n1124 0.04
R2921 vn_p.n1123 vn_p.n1122 0.04
R2922 vn_p.n1418 vn_p.n1417 0.04
R2923 vn_p.n1416 vn_p.n1415 0.04
R2924 vn_p.n1414 vn_p.n1413 0.04
R2925 vn_p.n1412 vn_p.n1411 0.04
R2926 vn_p.n1410 vn_p.n1409 0.04
R2927 vn_p.n1408 vn_p.n1407 0.04
R2928 vn_p.n1406 vn_p.n1405 0.04
R2929 vn_p.n1404 vn_p.n1403 0.04
R2930 vn_p.n1402 vn_p.n1401 0.04
R2931 vn_p.n1400 vn_p.n1399 0.04
R2932 vn_p.n1398 vn_p.n1397 0.04
R2933 vn_p.n1396 vn_p.n1395 0.04
R2934 vn_p.n1394 vn_p.n1393 0.04
R2935 vn_p.n1392 vn_p.n1391 0.04
R2936 vn_p.n1390 vn_p.n1389 0.04
R2937 vn_p.n1388 vn_p.n1387 0.04
R2938 vn_p.n1386 vn_p.n1385 0.04
R2939 vn_p.n1384 vn_p.n1383 0.04
R2940 vn_p.n1382 vn_p.n1381 0.04
R2941 vn_p.n1380 vn_p.n1379 0.04
R2942 vn_p.n1378 vn_p.n1377 0.04
R2943 vn_p.n1376 vn_p.n1375 0.04
R2944 vn_p.n1374 vn_p.n1373 0.04
R2945 vn_p.n1372 vn_p.n1371 0.04
R2946 vn_p.n1370 vn_p.n1369 0.04
R2947 vn_p.n1368 vn_p.n1367 0.04
R2948 vn_p.n1366 vn_p.n1365 0.04
R2949 vn_p.n1364 vn_p.n1363 0.04
R2950 vn_p.n1362 vn_p.n1361 0.04
R2951 vn_p.n1360 vn_p.n1359 0.04
R2952 vn_p.n1358 vn_p.n1357 0.04
R2953 vn_p.n1356 vn_p.n1355 0.04
R2954 vn_p.n1354 vn_p.n1353 0.04
R2955 vn_p.n1352 vn_p.n1351 0.04
R2956 vn_p.n1350 vn_p.n1349 0.04
R2957 vn_p.n1348 vn_p.n1347 0.04
R2958 vn_p.n1346 vn_p.n1345 0.04
R2959 vn_p.n1344 vn_p.n1343 0.04
R2960 vn_p.n1342 vn_p.n1341 0.04
R2961 vn_p.n1340 vn_p.n1339 0.04
R2962 vn_p.n1338 vn_p.n1337 0.04
R2963 vn_p.n1336 vn_p.n1335 0.04
R2964 vn_p.n1334 vn_p.n1333 0.04
R2965 vn_p.n1332 vn_p.n1331 0.04
R2966 vn_p.n1330 vn_p.n1329 0.04
R2967 vn_p.n1328 vn_p.n1327 0.04
R2968 vn_p.n1326 vn_p.n1325 0.04
R2969 vn_p.n1324 vn_p.n1323 0.04
R2970 vn_p.n1322 vn_p.n1321 0.04
R2971 vn_p.n1320 vn_p.n1319 0.04
R2972 vn_p.n1318 vn_p.n1317 0.04
R2973 vn_p.n1316 vn_p.n1315 0.04
R2974 vn_p.n1314 vn_p.n1313 0.04
R2975 vn_p.n1312 vn_p.n1311 0.04
R2976 vn_p.n1310 vn_p.n1309 0.04
R2977 vn_p.n1308 vn_p.n1307 0.04
R2978 vn_p.n1306 vn_p.n1305 0.04
R2979 vn_p.n1304 vn_p.n1303 0.04
R2980 vn_p.n1302 vn_p.n1301 0.04
R2981 vn_p.n1300 vn_p.n1299 0.04
R2982 vn_p.n1298 vn_p.n1297 0.04
R2983 vn_p.n1296 vn_p.n1295 0.04
R2984 vn_p.n1294 vn_p.n1293 0.04
R2985 vn_p.n1292 vn_p.n1291 0.04
R2986 vn_p.n1290 vn_p.n1289 0.04
R2987 vn_p.n1288 vn_p.n1287 0.04
R2988 vn_p.n1286 vn_p.n1285 0.04
R2989 vn_p.n1284 vn_p.n1283 0.04
R2990 vn_p.n1282 vn_p.n1281 0.04
R2991 vn_p.n1280 vn_p.n1279 0.04
R2992 vn_p.n1278 vn_p.n1277 0.04
R2993 vn_p.n1276 vn_p.n1275 0.04
R2994 vn_p.n1274 vn_p.n1273 0.04
R2995 vn_p.n1272 vn_p.n1271 0.04
R2996 vn_p vn_p.n1497 0.028
R2997 vn_p vn_p.n1494 0.027
R2998 vn_p vn_p.n748 0.005
R2999 vdd2.n440 vdd2.n439 9250.59
R3000 vdd2.n434 vdd2.n429 9250.59
R3001 vdd2.n433 vdd2.n432 2878.29
R3002 vdd2.n438 vdd2.n437 2869.55
R3003 vdd2.n441 vdd2.n434 2247.42
R3004 vdd2.n441 vdd2.n440 2247.42
R3005 vdd2.n433 vdd2.n430 940.477
R3006 vdd2.n438 vdd2.n435 940.476
R3007 vdd2.n434 vdd2.n433 940.476
R3008 vdd2.n440 vdd2.n438 940.476
R3009 vdd2.n502 vdd2.t752 10.284
R3010 vdd2.n23 vdd2.t1165 8.711
R3011 vdd2.n31 vdd2.t76 8.131
R3012 vdd2.n30 vdd2.t320 8.131
R3013 vdd2.n29 vdd2.t1246 8.131
R3014 vdd2.n28 vdd2.t671 8.131
R3015 vdd2.n27 vdd2.t913 8.131
R3016 vdd2.n26 vdd2.t1205 8.131
R3017 vdd2.n25 vdd2.t633 8.131
R3018 vdd2.n24 vdd2.t70 8.131
R3019 vdd2.n23 vdd2.t1446 8.131
R3020 vdd2.n510 vdd2.t1169 8.126
R3021 vdd2.n509 vdd2.t1400 8.126
R3022 vdd2.n508 vdd2.t837 8.126
R3023 vdd2.n507 vdd2.t273 8.126
R3024 vdd2.n506 vdd2.t502 8.126
R3025 vdd2.n505 vdd2.t787 8.126
R3026 vdd2.n504 vdd2.t230 8.126
R3027 vdd2.n503 vdd2.t1163 8.126
R3028 vdd2.n502 vdd2.t1029 8.126
R3029 vdd2.n511 vdd2.t177 8.126
R3030 vdd2.n511 vdd2.t1104 8.126
R3031 vdd2.n512 vdd2.t456 8.126
R3032 vdd2.n512 vdd2.t1376 8.126
R3033 vdd2.n513 vdd2.t583 8.126
R3034 vdd2.n513 vdd2.t8 8.126
R3035 vdd2.n514 vdd2.t1155 8.126
R3036 vdd2.n514 vdd2.t576 8.126
R3037 vdd2.n515 vdd2.t212 8.126
R3038 vdd2.n515 vdd2.t1138 8.126
R3039 vdd2.n516 vdd2.t1425 8.126
R3040 vdd2.n516 vdd2.t855 8.126
R3041 vdd2.n517 vdd2.t1197 8.126
R3042 vdd2.n517 vdd2.t614 8.126
R3043 vdd2.n518 vdd2.t264 8.126
R3044 vdd2.n518 vdd2.t1186 8.126
R3045 vdd2.n519 vdd2.t828 8.126
R3046 vdd2.n519 vdd2.t257 8.126
R3047 vdd2.n520 vdd2.t590 8.126
R3048 vdd2.n520 vdd2.t16 8.126
R3049 vdd2.n522 vdd2.t1134 8.126
R3050 vdd2.n522 vdd2.t553 8.126
R3051 vdd2.n523 vdd2.t1409 8.126
R3052 vdd2.n523 vdd2.t838 8.126
R3053 vdd2.n524 vdd2.t40 8.126
R3054 vdd2.n524 vdd2.t962 8.126
R3055 vdd2.n525 vdd2.t604 8.126
R3056 vdd2.n525 vdd2.t34 8.126
R3057 vdd2.n526 vdd2.t1170 8.126
R3058 vdd2.n526 vdd2.t591 8.126
R3059 vdd2.n527 vdd2.t883 8.126
R3060 vdd2.n527 vdd2.t312 8.126
R3061 vdd2.n528 vdd2.t642 8.126
R3062 vdd2.n528 vdd2.t68 8.126
R3063 vdd2.n529 vdd2.t1216 8.126
R3064 vdd2.n529 vdd2.t631 8.126
R3065 vdd2.n530 vdd2.t288 8.126
R3066 vdd2.n530 vdd2.t1212 8.126
R3067 vdd2.n531 vdd2.t46 8.126
R3068 vdd2.n531 vdd2.t970 8.126
R3069 vdd2.n533 vdd2.t1476 8.126
R3070 vdd2.n533 vdd2.t898 8.126
R3071 vdd2.n534 vdd2.t265 8.126
R3072 vdd2.n534 vdd2.t1187 8.126
R3073 vdd2.n535 vdd2.t385 8.126
R3074 vdd2.n535 vdd2.t1298 8.126
R3075 vdd2.n536 vdd2.t954 8.126
R3076 vdd2.n536 vdd2.t376 8.126
R3077 vdd2.n537 vdd2.t17 8.126
R3078 vdd2.n537 vdd2.t935 8.126
R3079 vdd2.n538 vdd2.t1232 8.126
R3080 vdd2.n538 vdd2.t648 8.126
R3081 vdd2.n539 vdd2.t994 8.126
R3082 vdd2.n539 vdd2.t419 8.126
R3083 vdd2.n540 vdd2.t60 8.126
R3084 vdd2.n540 vdd2.t987 8.126
R3085 vdd2.n541 vdd2.t627 8.126
R3086 vdd2.n541 vdd2.t57 8.126
R3087 vdd2.n542 vdd2.t392 8.126
R3088 vdd2.n542 vdd2.t1306 8.126
R3089 vdd2.n544 vdd2.t1185 8.126
R3090 vdd2.n544 vdd2.t1217 8.126
R3091 vdd2.n545 vdd2.t1462 8.126
R3092 vdd2.n545 vdd2.t1499 8.126
R3093 vdd2.n546 vdd2.t83 8.126
R3094 vdd2.n546 vdd2.t108 8.126
R3095 vdd2.n547 vdd2.t652 8.126
R3096 vdd2.n547 vdd2.t679 8.126
R3097 vdd2.n548 vdd2.t1222 8.126
R3098 vdd2.n548 vdd2.t1248 8.126
R3099 vdd2.n549 vdd2.t931 8.126
R3100 vdd2.n549 vdd2.t966 8.126
R3101 vdd2.n550 vdd2.t689 8.126
R3102 vdd2.n550 vdd2.t721 8.126
R3103 vdd2.n551 vdd2.t1257 8.126
R3104 vdd2.n551 vdd2.t1288 8.126
R3105 vdd2.n552 vdd2.t334 8.126
R3106 vdd2.n552 vdd2.t362 8.126
R3107 vdd2.n553 vdd2.t86 8.126
R3108 vdd2.n553 vdd2.t116 8.126
R3109 vdd2.n555 vdd2.t630 8.126
R3110 vdd2.n555 vdd2.t61 8.126
R3111 vdd2.n556 vdd2.t916 8.126
R3112 vdd2.n556 vdd2.t341 8.126
R3113 vdd2.n557 vdd2.t1030 8.126
R3114 vdd2.n557 vdd2.t459 8.126
R3115 vdd2.n558 vdd2.t101 8.126
R3116 vdd2.n558 vdd2.t1025 8.126
R3117 vdd2.n559 vdd2.t663 8.126
R3118 vdd2.n559 vdd2.t87 8.126
R3119 vdd2.n560 vdd2.t389 8.126
R3120 vdd2.n560 vdd2.t1302 8.126
R3121 vdd2.n561 vdd2.t141 8.126
R3122 vdd2.n561 vdd2.t1066 8.126
R3123 vdd2.n562 vdd2.t709 8.126
R3124 vdd2.n562 vdd2.t131 8.126
R3125 vdd2.n563 vdd2.t1280 8.126
R3126 vdd2.n563 vdd2.t702 8.126
R3127 vdd2.n564 vdd2.t1037 8.126
R3128 vdd2.n564 vdd2.t466 8.126
R3129 vdd2.n566 vdd2.t986 8.126
R3130 vdd2.n566 vdd2.t411 8.126
R3131 vdd2.n567 vdd2.t1258 8.126
R3132 vdd2.n567 vdd2.t682 8.126
R3133 vdd2.n568 vdd2.t1380 8.126
R3134 vdd2.n568 vdd2.t805 8.126
R3135 vdd2.n569 vdd2.t453 8.126
R3136 vdd2.n569 vdd2.t1372 8.126
R3137 vdd2.n570 vdd2.t1010 8.126
R3138 vdd2.n570 vdd2.t441 8.126
R3139 vdd2.n571 vdd2.t729 8.126
R3140 vdd2.n571 vdd2.t151 8.126
R3141 vdd2.n572 vdd2.t489 8.126
R3142 vdd2.n572 vdd2.t1414 8.126
R3143 vdd2.n573 vdd2.t1055 8.126
R3144 vdd2.n573 vdd2.t478 8.126
R3145 vdd2.n574 vdd2.t122 8.126
R3146 vdd2.n574 vdd2.t1045 8.126
R3147 vdd2.n575 vdd2.t1386 8.126
R3148 vdd2.n575 vdd2.t812 8.126
R3149 vdd2.n577 vdd2.t437 8.126
R3150 vdd2.n577 vdd2.t1352 8.126
R3151 vdd2.n578 vdd2.t711 8.126
R3152 vdd2.n578 vdd2.t132 8.126
R3153 vdd2.n579 vdd2.t842 8.126
R3154 vdd2.n579 vdd2.t267 8.126
R3155 vdd2.n580 vdd2.t1402 8.126
R3156 vdd2.n580 vdd2.t831 8.126
R3157 vdd2.n581 vdd2.t467 8.126
R3158 vdd2.n581 vdd2.t1387 8.126
R3159 vdd2.n582 vdd2.t185 8.126
R3160 vdd2.n582 vdd2.t1112 8.126
R3161 vdd2.n583 vdd2.t1444 8.126
R3162 vdd2.n583 vdd2.t871 8.126
R3163 vdd2.n584 vdd2.t510 8.126
R3164 vdd2.n584 vdd2.t1434 8.126
R3165 vdd2.n585 vdd2.t1081 8.126
R3166 vdd2.n585 vdd2.t505 8.126
R3167 vdd2.n586 vdd2.t849 8.126
R3168 vdd2.n586 vdd2.t274 8.126
R3169 vdd2.n588 vdd2.t777 8.126
R3170 vdd2.n588 vdd2.t203 8.126
R3171 vdd2.n589 vdd2.t1056 8.126
R3172 vdd2.n589 vdd2.t479 8.126
R3173 vdd2.n590 vdd2.t1192 8.126
R3174 vdd2.n590 vdd2.t608 8.126
R3175 vdd2.n591 vdd2.t258 8.126
R3176 vdd2.n591 vdd2.t1180 8.126
R3177 vdd2.n592 vdd2.t813 8.126
R3178 vdd2.n592 vdd2.t238 8.126
R3179 vdd2.n593 vdd2.t529 8.126
R3180 vdd2.n593 vdd2.t1453 8.126
R3181 vdd2.n594 vdd2.t302 8.126
R3182 vdd2.n594 vdd2.t1221 8.126
R3183 vdd2.n595 vdd2.t863 8.126
R3184 vdd2.n595 vdd2.t291 8.126
R3185 vdd2.n596 vdd2.t1427 8.126
R3186 vdd2.n596 vdd2.t857 8.126
R3187 vdd2.n597 vdd2.t1198 8.126
R3188 vdd2.n597 vdd2.t615 8.126
R3189 vdd2.n599 vdd2.t1092 8.126
R3190 vdd2.n599 vdd2.t511 8.126
R3191 vdd2.n600 vdd2.t1371 8.126
R3192 vdd2.n600 vdd2.t797 8.126
R3193 vdd2.n601 vdd2.t0 8.126
R3194 vdd2.n601 vdd2.t917 8.126
R3195 vdd2.n602 vdd2.t563 8.126
R3196 vdd2.n602 vdd2.t1486 8.126
R3197 vdd2.n603 vdd2.t1131 8.126
R3198 vdd2.n603 vdd2.t549 8.126
R3199 vdd2.n604 vdd2.t847 8.126
R3200 vdd2.n604 vdd2.t272 8.126
R3201 vdd2.n605 vdd2.t605 8.126
R3202 vdd2.n605 vdd2.t36 8.126
R3203 vdd2.n606 vdd2.t1177 8.126
R3204 vdd2.n606 vdd2.t597 8.126
R3205 vdd2.n607 vdd2.t243 8.126
R3206 vdd2.n607 vdd2.t1168 8.126
R3207 vdd2.n608 vdd2.t6 8.126
R3208 vdd2.n608 vdd2.t925 8.126
R3209 vdd2.n610 vdd2.t1433 8.126
R3210 vdd2.n610 vdd2.t864 8.126
R3211 vdd2.n611 vdd2.t222 8.126
R3212 vdd2.n611 vdd2.t1146 8.126
R3213 vdd2.n612 vdd2.t343 8.126
R3214 vdd2.n612 vdd2.t1261 8.126
R3215 vdd2.n613 vdd2.t908 8.126
R3216 vdd2.n613 vdd2.t336 8.126
R3217 vdd2.n614 vdd2.t1472 8.126
R3218 vdd2.n614 vdd2.t893 8.126
R3219 vdd2.n615 vdd2.t1196 8.126
R3220 vdd2.n615 vdd2.t612 8.126
R3221 vdd2.n616 vdd2.t955 8.126
R3222 vdd2.n616 vdd2.t377 8.126
R3223 vdd2.n617 vdd2.t25 8.126
R3224 vdd2.n617 vdd2.t943 8.126
R3225 vdd2.n618 vdd2.t588 8.126
R3226 vdd2.n618 vdd2.t14 8.126
R3227 vdd2.n619 vdd2.t350 8.126
R3228 vdd2.n619 vdd2.t1267 8.126
R3229 vdd2.n621 vdd2.t292 8.126
R3230 vdd2.n621 vdd2.t321 8.126
R3231 vdd2.n622 vdd2.t564 8.126
R3232 vdd2.n622 vdd2.t599 8.126
R3233 vdd2.n623 vdd2.t685 8.126
R3234 vdd2.n623 vdd2.t714 8.126
R3235 vdd2.n624 vdd2.t1254 8.126
R3236 vdd2.n624 vdd2.t1281 8.126
R3237 vdd2.n625 vdd2.t325 8.126
R3238 vdd2.n625 vdd2.t351 8.126
R3239 vdd2.n626 vdd2.t42 8.126
R3240 vdd2.n626 vdd2.t66 8.126
R3241 vdd2.n627 vdd2.t1293 8.126
R3242 vdd2.n627 vdd2.t1322 8.126
R3243 vdd2.n628 vdd2.t365 8.126
R3244 vdd2.n628 vdd2.t402 8.126
R3245 vdd2.n629 vdd2.t933 8.126
R3246 vdd2.n629 vdd2.t969 8.126
R3247 vdd2.n630 vdd2.t690 8.126
R3248 vdd2.n630 vdd2.t723 8.126
R3249 vdd2.n632 vdd2.t1238 8.126
R3250 vdd2.n632 vdd2.t656 8.126
R3251 vdd2.n633 vdd2.t26 8.126
R3252 vdd2.n633 vdd2.t944 8.126
R3253 vdd2.n634 vdd2.t134 8.126
R3254 vdd2.n634 vdd2.t1059 8.126
R3255 vdd2.n635 vdd2.t703 8.126
R3256 vdd2.n635 vdd2.t125 8.126
R3257 vdd2.n636 vdd2.t1268 8.126
R3258 vdd2.n636 vdd2.t691 8.126
R3259 vdd2.n637 vdd2.t993 8.126
R3260 vdd2.n637 vdd2.t417 8.126
R3261 vdd2.n638 vdd2.t748 8.126
R3262 vdd2.n638 vdd2.t173 8.126
R3263 vdd2.n639 vdd2.t1312 8.126
R3264 vdd2.n639 vdd2.t738 8.126
R3265 vdd2.n640 vdd2.t391 8.126
R3266 vdd2.n640 vdd2.t1304 8.126
R3267 vdd2.n641 vdd2.t143 8.126
R3268 vdd2.n641 vdd2.t1067 8.126
R3269 vdd2.n643 vdd2.t80 8.126
R3270 vdd2.n643 vdd2.t1006 8.126
R3271 vdd2.n644 vdd2.t367 8.126
R3272 vdd2.n644 vdd2.t1283 8.126
R3273 vdd2.n645 vdd2.t485 8.126
R3274 vdd2.n645 vdd2.t1407 8.126
R3275 vdd2.n646 vdd2.t1049 8.126
R3276 vdd2.n646 vdd2.t475 8.126
R3277 vdd2.n647 vdd2.t111 8.126
R3278 vdd2.n647 vdd2.t1033 8.126
R3279 vdd2.n648 vdd2.t1330 8.126
R3280 vdd2.n648 vdd2.t757 8.126
R3281 vdd2.n649 vdd2.t1100 8.126
R3282 vdd2.n649 vdd2.t518 8.126
R3283 vdd2.n650 vdd2.t165 8.126
R3284 vdd2.n650 vdd2.t1085 8.126
R3285 vdd2.n651 vdd2.t732 8.126
R3286 vdd2.n651 vdd2.t154 8.126
R3287 vdd2.n652 vdd2.t491 8.126
R3288 vdd2.n652 vdd2.t1416 8.126
R3289 vdd2.n654 vdd2.t401 8.126
R3290 vdd2.n654 vdd2.t1313 8.126
R3291 vdd2.n655 vdd2.t674 8.126
R3292 vdd2.n655 vdd2.t96 8.126
R3293 vdd2.n656 vdd2.t798 8.126
R3294 vdd2.n656 vdd2.t223 8.126
R3295 vdd2.n657 vdd2.t1360 8.126
R3296 vdd2.n657 vdd2.t788 8.126
R3297 vdd2.n658 vdd2.t434 8.126
R3298 vdd2.n658 vdd2.t1349 8.126
R3299 vdd2.n659 vdd2.t140 8.126
R3300 vdd2.n659 vdd2.t1065 8.126
R3301 vdd2.n660 vdd2.t1404 8.126
R3302 vdd2.n660 vdd2.t833 8.126
R3303 vdd2.n661 vdd2.t471 8.126
R3304 vdd2.n661 vdd2.t1393 8.126
R3305 vdd2.n662 vdd2.t1036 8.126
R3306 vdd2.n662 vdd2.t465 8.126
R3307 vdd2.n663 vdd2.t801 8.126
R3308 vdd2.n663 vdd2.t231 8.126
R3309 vdd2.n665 vdd2.t739 8.126
R3310 vdd2.n665 vdd2.t164 8.126
R3311 vdd2.n666 vdd2.t1017 8.126
R3312 vdd2.n666 vdd2.t447 8.126
R3313 vdd2.n667 vdd2.t1150 8.126
R3314 vdd2.n667 vdd2.t568 8.126
R3315 vdd2.n668 vdd2.t215 8.126
R3316 vdd2.n668 vdd2.t1139 8.126
R3317 vdd2.n669 vdd2.t774 8.126
R3318 vdd2.n669 vdd2.t200 8.126
R3319 vdd2.n670 vdd2.t488 8.126
R3320 vdd2.n670 vdd2.t1412 8.126
R3321 vdd2.n671 vdd2.t260 8.126
R3322 vdd2.n671 vdd2.t1181 8.126
R3323 vdd2.n672 vdd2.t822 8.126
R3324 vdd2.n672 vdd2.t248 8.126
R3325 vdd2.n673 vdd2.t1385 8.126
R3326 vdd2.n673 vdd2.t811 8.126
R3327 vdd2.n674 vdd2.t1156 8.126
R3328 vdd2.n674 vdd2.t578 8.126
R3329 vdd2.n676 vdd2.t1086 8.126
R3330 vdd2.n676 vdd2.t78 8.126
R3331 vdd2.n677 vdd2.t1364 8.126
R3332 vdd2.n677 vdd2.t366 8.126
R3333 vdd2.n678 vdd2.t1494 8.126
R3334 vdd2.n678 vdd2.t481 8.126
R3335 vdd2.n679 vdd2.t558 8.126
R3336 vdd2.n679 vdd2.t1048 8.126
R3337 vdd2.n680 vdd2.t1129 8.126
R3338 vdd2.n680 vdd2.t110 8.126
R3339 vdd2.n681 vdd2.t841 8.126
R3340 vdd2.n681 vdd2.t1326 8.126
R3341 vdd2.n682 vdd2.t603 8.126
R3342 vdd2.n682 vdd2.t1097 8.126
R3343 vdd2.n683 vdd2.t1172 8.126
R3344 vdd2.n683 vdd2.t162 8.126
R3345 vdd2.n684 vdd2.t236 8.126
R3346 vdd2.n684 vdd2.t728 8.126
R3347 vdd2.n685 vdd2.t3 8.126
R3348 vdd2.n685 vdd2.t490 8.126
R3349 vdd2.n687 vdd2.t1005 8.126
R3350 vdd2.n687 vdd2.t433 8.126
R3351 vdd2.n688 vdd2.t1282 8.126
R3352 vdd2.n688 vdd2.t706 8.126
R3353 vdd2.n689 vdd2.t1405 8.126
R3354 vdd2.n689 vdd2.t834 8.126
R3355 vdd2.n690 vdd2.t473 8.126
R3356 vdd2.n690 vdd2.t1395 8.126
R3357 vdd2.n691 vdd2.t1032 8.126
R3358 vdd2.n691 vdd2.t462 8.126
R3359 vdd2.n692 vdd2.t754 8.126
R3360 vdd2.n692 vdd2.t179 8.126
R3361 vdd2.n693 vdd2.t517 8.126
R3362 vdd2.n693 vdd2.t1439 8.126
R3363 vdd2.n694 vdd2.t1084 8.126
R3364 vdd2.n694 vdd2.t506 8.126
R3365 vdd2.n695 vdd2.t152 8.126
R3366 vdd2.n695 vdd2.t1074 8.126
R3367 vdd2.n696 vdd2.t1415 8.126
R3368 vdd2.n696 vdd2.t844 8.126
R3369 vdd2.n698 vdd2.t1348 8.126
R3370 vdd2.n698 vdd2.t773 8.126
R3371 vdd2.n699 vdd2.t128 8.126
R3372 vdd2.n699 vdd2.t1053 8.126
R3373 vdd2.n700 vdd2.t261 8.126
R3374 vdd2.n700 vdd2.t1183 8.126
R3375 vdd2.n701 vdd2.t824 8.126
R3376 vdd2.n701 vdd2.t251 8.126
R3377 vdd2.n702 vdd2.t1382 8.126
R3378 vdd2.n702 vdd2.t806 8.126
R3379 vdd2.n703 vdd2.t1106 8.126
R3380 vdd2.n703 vdd2.t524 8.126
R3381 vdd2.n704 vdd2.t867 8.126
R3382 vdd2.n704 vdd2.t297 8.126
R3383 vdd2.n705 vdd2.t1429 8.126
R3384 vdd2.n705 vdd2.t860 8.126
R3385 vdd2.n706 vdd2.t497 8.126
R3386 vdd2.n706 vdd2.t1422 8.126
R3387 vdd2.n707 vdd2.t269 8.126
R3388 vdd2.n707 vdd2.t1194 8.126
R3389 vdd2.n709 vdd2.t163 8.126
R3390 vdd2.n709 vdd2.t1083 8.126
R3391 vdd2.n710 vdd2.t446 8.126
R3392 vdd2.n710 vdd2.t1363 8.126
R3393 vdd2.n711 vdd2.t567 8.126
R3394 vdd2.n711 vdd2.t1491 8.126
R3395 vdd2.n712 vdd2.t1137 8.126
R3396 vdd2.n712 vdd2.t557 8.126
R3397 vdd2.n713 vdd2.t199 8.126
R3398 vdd2.n713 vdd2.t1128 8.126
R3399 vdd2.n714 vdd2.t1411 8.126
R3400 vdd2.n714 vdd2.t840 8.126
R3401 vdd2.n715 vdd2.t1179 8.126
R3402 vdd2.n715 vdd2.t600 8.126
R3403 vdd2.n716 vdd2.t247 8.126
R3404 vdd2.n716 vdd2.t1171 8.126
R3405 vdd2.n717 vdd2.t810 8.126
R3406 vdd2.n717 vdd2.t235 8.126
R3407 vdd2.n718 vdd2.t577 8.126
R3408 vdd2.n718 vdd2.t1 8.126
R3409 vdd2.n720 vdd2.t507 8.126
R3410 vdd2.n720 vdd2.t1430 8.126
R3411 vdd2.n721 vdd2.t793 8.126
R3412 vdd2.n721 vdd2.t217 8.126
R3413 vdd2.n722 vdd2.t911 8.126
R3414 vdd2.n722 vdd2.t339 8.126
R3415 vdd2.n723 vdd2.t1481 8.126
R3416 vdd2.n723 vdd2.t901 8.126
R3417 vdd2.n724 vdd2.t546 8.126
R3418 vdd2.n724 vdd2.t1469 8.126
R3419 vdd2.n725 vdd2.t266 8.126
R3420 vdd2.n725 vdd2.t1188 8.126
R3421 vdd2.n726 vdd2.t29 8.126
R3422 vdd2.n726 vdd2.t947 8.126
R3423 vdd2.n727 vdd2.t592 8.126
R3424 vdd2.n727 vdd2.t18 8.126
R3425 vdd2.n728 vdd2.t1162 8.126
R3426 vdd2.n728 vdd2.t584 8.126
R3427 vdd2.n729 vdd2.t920 8.126
R3428 vdd2.n729 vdd2.t346 8.126
R3429 vdd2.n731 vdd2.t1461 8.126
R3430 vdd2.n731 vdd2.t885 8.126
R3431 vdd2.n732 vdd2.t249 8.126
R3432 vdd2.n732 vdd2.t1173 8.126
R3433 vdd2.n733 vdd2.t369 8.126
R3434 vdd2.n733 vdd2.t1284 8.126
R3435 vdd2.n734 vdd2.t934 8.126
R3436 vdd2.n734 vdd2.t357 8.126
R3437 vdd2.n735 vdd2.t2 8.126
R3438 vdd2.n735 vdd2.t921 8.126
R3439 vdd2.n736 vdd2.t1220 8.126
R3440 vdd2.n736 vdd2.t634 8.126
R3441 vdd2.n737 vdd2.t983 8.126
R3442 vdd2.n737 vdd2.t406 8.126
R3443 vdd2.n738 vdd2.t48 8.126
R3444 vdd2.n738 vdd2.t972 8.126
R3445 vdd2.n739 vdd2.t613 8.126
R3446 vdd2.n739 vdd2.t41 8.126
R3447 vdd2.n740 vdd2.t378 8.126
R3448 vdd2.n740 vdd2.t1292 8.126
R3449 vdd2.n742 vdd2.t316 8.126
R3450 vdd2.n742 vdd2.t1236 8.126
R3451 vdd2.n743 vdd2.t594 8.126
R3452 vdd2.n743 vdd2.t22 8.126
R3453 vdd2.n744 vdd2.t707 8.126
R3454 vdd2.n744 vdd2.t129 8.126
R3455 vdd2.n745 vdd2.t1275 8.126
R3456 vdd2.n745 vdd2.t696 8.126
R3457 vdd2.n746 vdd2.t348 8.126
R3458 vdd2.n746 vdd2.t1265 8.126
R3459 vdd2.n747 vdd2.t62 8.126
R3460 vdd2.n747 vdd2.t988 8.126
R3461 vdd2.n748 vdd2.t1318 8.126
R3462 vdd2.n748 vdd2.t743 8.126
R3463 vdd2.n749 vdd2.t394 8.126
R3464 vdd2.n749 vdd2.t1308 8.126
R3465 vdd2.n750 vdd2.t961 8.126
R3466 vdd2.n750 vdd2.t386 8.126
R3467 vdd2.n751 vdd2.t716 8.126
R3468 vdd2.n751 vdd2.t136 8.126
R3469 vdd2.n753 vdd2.t653 8.126
R3470 vdd2.n753 vdd2.t680 8.126
R3471 vdd2.n754 vdd2.t939 8.126
R3472 vdd2.n754 vdd2.t974 8.126
R3473 vdd2.n755 vdd2.t1054 8.126
R3474 vdd2.n755 vdd2.t1089 8.126
R3475 vdd2.n756 vdd2.t119 8.126
R3476 vdd2.n756 vdd2.t156 8.126
R3477 vdd2.n757 vdd2.t687 8.126
R3478 vdd2.n757 vdd2.t717 8.126
R3479 vdd2.n758 vdd2.t412 8.126
R3480 vdd2.n758 vdd2.t438 8.126
R3481 vdd2.n759 vdd2.t167 8.126
R3482 vdd2.n759 vdd2.t197 8.126
R3483 vdd2.n760 vdd2.t733 8.126
R3484 vdd2.n760 vdd2.t762 8.126
R3485 vdd2.n761 vdd2.t1299 8.126
R3486 vdd2.n761 vdd2.t1329 8.126
R3487 vdd2.n762 vdd2.t1061 8.126
R3488 vdd2.n762 vdd2.t1099 8.126
R3489 vdd2.n764 vdd2.t973 8.126
R3490 vdd2.n764 vdd2.t393 8.126
R3491 vdd2.n765 vdd2.t1249 8.126
R3492 vdd2.n765 vdd2.t667 8.126
R3493 vdd2.n766 vdd2.t1365 8.126
R3494 vdd2.n766 vdd2.t794 8.126
R3495 vdd2.n767 vdd2.t440 8.126
R3496 vdd2.n767 vdd2.t1356 8.126
R3497 vdd2.n768 vdd2.t1004 8.126
R3498 vdd2.n768 vdd2.t432 8.126
R3499 vdd2.n769 vdd2.t712 8.126
R3500 vdd2.n769 vdd2.t133 8.126
R3501 vdd2.n770 vdd2.t474 8.126
R3502 vdd2.n770 vdd2.t1396 8.126
R3503 vdd2.n771 vdd2.t1040 8.126
R3504 vdd2.n771 vdd2.t468 8.126
R3505 vdd2.n772 vdd2.t109 8.126
R3506 vdd2.n772 vdd2.t1031 8.126
R3507 vdd2.n773 vdd2.t1374 8.126
R3508 vdd2.n773 vdd2.t799 8.126
R3509 vdd2.n775 vdd2.t1307 8.126
R3510 vdd2.n775 vdd2.t734 8.126
R3511 vdd2.n776 vdd2.t92 8.126
R3512 vdd2.n776 vdd2.t1014 8.126
R3513 vdd2.n777 vdd2.t219 8.126
R3514 vdd2.n777 vdd2.t1144 8.126
R3515 vdd2.n778 vdd2.t782 8.126
R3516 vdd2.n778 vdd2.t208 8.126
R3517 vdd2.n779 vdd2.t1345 8.126
R3518 vdd2.n779 vdd2.t770 8.126
R3519 vdd2.n780 vdd2.t1057 8.126
R3520 vdd2.n780 vdd2.t480 8.126
R3521 vdd2.n781 vdd2.t825 8.126
R3522 vdd2.n781 vdd2.t252 8.126
R3523 vdd2.n782 vdd2.t1388 8.126
R3524 vdd2.n782 vdd2.t814 8.126
R3525 vdd2.n783 vdd2.t460 8.126
R3526 vdd2.n783 vdd2.t1381 8.126
R3527 vdd2.n784 vdd2.t228 8.126
R3528 vdd2.n784 vdd2.t1153 8.126
R3529 vdd2.n786 vdd2.t764 8.126
R3530 vdd2.n786 vdd2.t190 8.126
R3531 vdd2.n787 vdd2.t1041 8.126
R3532 vdd2.n787 vdd2.t469 8.126
R3533 vdd2.n788 vdd2.t1174 8.126
R3534 vdd2.n788 vdd2.t595 8.126
R3535 vdd2.n789 vdd2.t237 8.126
R3536 vdd2.n789 vdd2.t1164 8.126
R3537 vdd2.n790 vdd2.t800 8.126
R3538 vdd2.n790 vdd2.t229 8.126
R3539 vdd2.n791 vdd2.t513 8.126
R3540 vdd2.n791 vdd2.t1437 8.126
R3541 vdd2.n792 vdd2.t285 8.126
R3542 vdd2.n792 vdd2.t1208 8.126
R3543 vdd2.n793 vdd2.t851 8.126
R3544 vdd2.n793 vdd2.t277 8.126
R3545 vdd2.n794 vdd2.t1413 8.126
R3546 vdd2.n794 vdd2.t843 8.126
R3547 vdd2.n795 vdd2.t1182 8.126
R3548 vdd2.n795 vdd2.t602 8.126
R3549 vdd2.n797 vdd2.t1115 8.126
R3550 vdd2.n797 vdd2.t533 8.126
R3551 vdd2.n798 vdd2.t1391 8.126
R3552 vdd2.n798 vdd2.t818 8.126
R3553 vdd2.n799 vdd2.t23 8.126
R3554 vdd2.n799 vdd2.t940 8.126
R3555 vdd2.n800 vdd2.t585 8.126
R3556 vdd2.n800 vdd2.t10 8.126
R3557 vdd2.n801 vdd2.t1154 8.126
R3558 vdd2.n801 vdd2.t573 8.126
R3559 vdd2.n802 vdd2.t865 8.126
R3560 vdd2.n802 vdd2.t293 8.126
R3561 vdd2.n803 vdd2.t624 8.126
R3562 vdd2.n803 vdd2.t51 8.126
R3563 vdd2.n804 vdd2.t1199 8.126
R3564 vdd2.n804 vdd2.t618 8.126
R3565 vdd2.n805 vdd2.t268 8.126
R3566 vdd2.n805 vdd2.t1193 8.126
R3567 vdd2.n806 vdd2.t30 8.126
R3568 vdd2.n806 vdd2.t951 8.126
R3569 vdd2.n808 vdd2.t1457 8.126
R3570 vdd2.n808 vdd2.t1489 8.126
R3571 vdd2.n809 vdd2.t244 8.126
R3572 vdd2.n809 vdd2.t278 8.126
R3573 vdd2.n810 vdd2.t363 8.126
R3574 vdd2.n810 vdd2.t399 8.126
R3575 vdd2.n811 vdd2.t928 8.126
R3576 vdd2.n811 vdd2.t964 8.126
R3577 vdd2.n812 vdd2.t1497 8.126
R3578 vdd2.n812 vdd2.t31 8.126
R3579 vdd2.n813 vdd2.t1213 8.126
R3580 vdd2.n813 vdd2.t1241 8.126
R3581 vdd2.n814 vdd2.t978 8.126
R3582 vdd2.n814 vdd2.t1001 8.126
R3583 vdd2.n815 vdd2.t43 8.126
R3584 vdd2.n815 vdd2.t72 8.126
R3585 vdd2.n816 vdd2.t610 8.126
R3586 vdd2.n816 vdd2.t636 8.126
R3587 vdd2.n817 vdd2.t373 8.126
R3588 vdd2.n817 vdd2.t408 8.126
R3589 vdd2.n819 vdd2.t276 8.126
R3590 vdd2.n819 vdd2.t1200 8.126
R3591 vdd2.n820 vdd2.t552 8.126
R3592 vdd2.n820 vdd2.t1475 8.126
R3593 vdd2.n821 vdd2.t668 8.126
R3594 vdd2.n821 vdd2.t94 8.126
R3595 vdd2.n822 vdd2.t1244 8.126
R3596 vdd2.n822 vdd2.t662 8.126
R3597 vdd2.n823 vdd2.t314 8.126
R3598 vdd2.n823 vdd2.t1235 8.126
R3599 vdd2.n824 vdd2.t27 8.126
R3600 vdd2.n824 vdd2.t945 8.126
R3601 vdd2.n825 vdd2.t1276 8.126
R3602 vdd2.n825 vdd2.t697 8.126
R3603 vdd2.n826 vdd2.t352 8.126
R3604 vdd2.n826 vdd2.t1269 8.126
R3605 vdd2.n827 vdd2.t918 8.126
R3606 vdd2.n827 vdd2.t344 8.126
R3607 vdd2.n828 vdd2.t676 8.126
R3608 vdd2.n828 vdd2.t98 8.126
R3609 vdd2.n830 vdd2.t617 8.126
R3610 vdd2.n830 vdd2.t645 8.126
R3611 vdd2.n831 vdd2.t897 8.126
R3612 vdd2.n831 vdd2.t927 8.126
R3613 vdd2.n832 vdd2.t1016 8.126
R3614 vdd2.n832 vdd2.t1043 8.126
R3615 vdd2.n833 vdd2.t85 8.126
R3616 vdd2.n833 vdd2.t112 8.126
R3617 vdd2.n834 vdd2.t651 8.126
R3618 vdd2.n834 vdd2.t677 8.126
R3619 vdd2.n835 vdd2.t368 8.126
R3620 vdd2.n835 vdd2.t405 8.126
R3621 vdd2.n836 vdd2.t120 8.126
R3622 vdd2.n836 vdd2.t158 8.126
R3623 vdd2.n837 vdd2.t692 8.126
R3624 vdd2.n837 vdd2.t725 8.126
R3625 vdd2.n838 vdd2.t1262 8.126
R3626 vdd2.n838 vdd2.t1291 8.126
R3627 vdd2.n839 vdd2.t1022 8.126
R3628 vdd2.n839 vdd2.t1052 8.126
R3629 vdd2.n841 vdd2.t71 8.126
R3630 vdd2.n841 vdd2.t996 8.126
R3631 vdd2.n842 vdd2.t354 8.126
R3632 vdd2.n842 vdd2.t1272 8.126
R3633 vdd2.n843 vdd2.t470 8.126
R3634 vdd2.n843 vdd2.t1392 8.126
R3635 vdd2.n844 vdd2.t1034 8.126
R3636 vdd2.n844 vdd2.t463 8.126
R3637 vdd2.n845 vdd2.t99 8.126
R3638 vdd2.n845 vdd2.t1023 8.126
R3639 vdd2.n846 vdd2.t1315 8.126
R3640 vdd2.n846 vdd2.t740 8.126
R3641 vdd2.n847 vdd2.t1077 8.126
R3642 vdd2.n847 vdd2.t500 8.126
R3643 vdd2.n848 vdd2.t145 8.126
R3644 vdd2.n848 vdd2.t1069 8.126
R3645 vdd2.n849 vdd2.t715 8.126
R3646 vdd2.n849 vdd2.t135 8.126
R3647 vdd2.n850 vdd2.t477 8.126
R3648 vdd2.n850 vdd2.t1398 8.126
R3649 vdd2.n491 vdd2.t421 8.126
R3650 vdd2.n491 vdd2.t1334 8.126
R3651 vdd2.n492 vdd2.t694 8.126
R3652 vdd2.n492 vdd2.t114 8.126
R3653 vdd2.n493 vdd2.t821 8.126
R3654 vdd2.n493 vdd2.t245 8.126
R3655 vdd2.n494 vdd2.t1383 8.126
R3656 vdd2.n494 vdd2.t807 8.126
R3657 vdd2.n495 vdd2.t452 8.126
R3658 vdd2.n495 vdd2.t1369 8.126
R3659 vdd2.n496 vdd2.t166 8.126
R3660 vdd2.n496 vdd2.t1087 8.126
R3661 vdd2.n497 vdd2.t1424 8.126
R3662 vdd2.n497 vdd2.t854 8.126
R3663 vdd2.n498 vdd2.t492 8.126
R3664 vdd2.n498 vdd2.t1417 8.126
R3665 vdd2.n499 vdd2.t1060 8.126
R3666 vdd2.n499 vdd2.t484 8.126
R3667 vdd2.n500 vdd2.t827 8.126
R3668 vdd2.n500 vdd2.t255 8.126
R3669 vdd2.n32 vdd2.t816 8.126
R3670 vdd2.n32 vdd2.t240 8.126
R3671 vdd2.n33 vdd2.t1103 8.126
R3672 vdd2.n33 vdd2.t521 8.126
R3673 vdd2.n34 vdd2.t1228 8.126
R3674 vdd2.n34 vdd2.t644 8.126
R3675 vdd2.n35 vdd2.t301 8.126
R3676 vdd2.n35 vdd2.t1219 8.126
R3677 vdd2.n36 vdd2.t859 8.126
R3678 vdd2.n36 vdd2.t284 8.126
R3679 vdd2.n37 vdd2.t566 8.126
R3680 vdd2.n37 vdd2.t1493 8.126
R3681 vdd2.n38 vdd2.t332 8.126
R3682 vdd2.n38 vdd2.t1252 8.126
R3683 vdd2.n39 vdd2.t894 8.126
R3684 vdd2.n39 vdd2.t327 8.126
R3685 vdd2.n40 vdd2.t1463 8.126
R3686 vdd2.n40 vdd2.t888 8.126
R3687 vdd2.n41 vdd2.t1233 8.126
R3688 vdd2.n41 vdd2.t649 8.126
R3689 vdd2.n43 vdd2.t501 8.126
R3690 vdd2.n43 vdd2.t534 8.126
R3691 vdd2.n44 vdd2.t786 8.126
R3692 vdd2.n44 vdd2.t820 8.126
R3693 vdd2.n45 vdd2.t907 8.126
R3694 vdd2.n45 vdd2.t942 8.126
R3695 vdd2.n46 vdd2.t1478 8.126
R3696 vdd2.n46 vdd2.t12 8.126
R3697 vdd2.n47 vdd2.t539 8.126
R3698 vdd2.n47 vdd2.t575 8.126
R3699 vdd2.n48 vdd2.t262 8.126
R3700 vdd2.n48 vdd2.t295 8.126
R3701 vdd2.n49 vdd2.t24 8.126
R3702 vdd2.n49 vdd2.t53 8.126
R3703 vdd2.n50 vdd2.t587 8.126
R3704 vdd2.n50 vdd2.t619 8.126
R3705 vdd2.n51 vdd2.t1159 8.126
R3706 vdd2.n51 vdd2.t1191 8.126
R3707 vdd2.n52 vdd2.t915 8.126
R3708 vdd2.n52 vdd2.t949 8.126
R3709 vdd2.n54 vdd2.t159 8.126
R3710 vdd2.n54 vdd2.t1078 8.126
R3711 vdd2.n55 vdd2.t445 8.126
R3712 vdd2.n55 vdd2.t1359 8.126
R3713 vdd2.n56 vdd2.t562 8.126
R3714 vdd2.n56 vdd2.t1487 8.126
R3715 vdd2.n57 vdd2.t1135 8.126
R3716 vdd2.n57 vdd2.t554 8.126
R3717 vdd2.n58 vdd2.t196 8.126
R3718 vdd2.n58 vdd2.t1122 8.126
R3719 vdd2.n59 vdd2.t1406 8.126
R3720 vdd2.n59 vdd2.t835 8.126
R3721 vdd2.n60 vdd2.t1176 8.126
R3722 vdd2.n60 vdd2.t596 8.126
R3723 vdd2.n61 vdd2.t239 8.126
R3724 vdd2.n61 vdd2.t1166 8.126
R3725 vdd2.n62 vdd2.t803 8.126
R3726 vdd2.n62 vdd2.t233 8.126
R3727 vdd2.n63 vdd2.t572 8.126
R3728 vdd2.n63 vdd2.t1496 8.126
R3729 vdd2.n65 vdd2.t1309 8.126
R3730 vdd2.n65 vdd2.t735 8.126
R3731 vdd2.n66 vdd2.t93 8.126
R3732 vdd2.n66 vdd2.t1015 8.126
R3733 vdd2.n67 vdd2.t220 8.126
R3734 vdd2.n67 vdd2.t1145 8.126
R3735 vdd2.n68 vdd2.t783 8.126
R3736 vdd2.n68 vdd2.t209 8.126
R3737 vdd2.n69 vdd2.t1346 8.126
R3738 vdd2.n69 vdd2.t771 8.126
R3739 vdd2.n70 vdd2.t1058 8.126
R3740 vdd2.n70 vdd2.t482 8.126
R3741 vdd2.n71 vdd2.t826 8.126
R3742 vdd2.n71 vdd2.t253 8.126
R3743 vdd2.n72 vdd2.t1390 8.126
R3744 vdd2.n72 vdd2.t815 8.126
R3745 vdd2.n73 vdd2.t461 8.126
R3746 vdd2.n73 vdd2.t1379 8.126
R3747 vdd2.n74 vdd2.t227 8.126
R3748 vdd2.n74 vdd2.t1152 8.126
R3749 vdd2.n76 vdd2.t359 8.126
R3750 vdd2.n76 vdd2.t1278 8.126
R3751 vdd2.n77 vdd2.t641 8.126
R3752 vdd2.n77 vdd2.t67 8.126
R3753 vdd2.n78 vdd2.t761 8.126
R3754 vdd2.n78 vdd2.t188 8.126
R3755 vdd2.n79 vdd2.t1325 8.126
R3756 vdd2.n79 vdd2.t753 8.126
R3757 vdd2.n80 vdd2.t404 8.126
R3758 vdd2.n80 vdd2.t1314 8.126
R3759 vdd2.n81 vdd2.t104 8.126
R3760 vdd2.n81 vdd2.t1027 8.126
R3761 vdd2.n82 vdd2.t1367 8.126
R3762 vdd2.n82 vdd2.t796 8.126
R3763 vdd2.n83 vdd2.t442 8.126
R3764 vdd2.n83 vdd2.t1357 8.126
R3765 vdd2.n84 vdd2.t1007 8.126
R3766 vdd2.n84 vdd2.t436 8.126
R3767 vdd2.n85 vdd2.t768 8.126
R3768 vdd2.n85 vdd2.t195 8.126
R3769 vdd2.n87 vdd2.t20 8.126
R3770 vdd2.n87 vdd2.t936 8.126
R3771 vdd2.n88 vdd2.t306 8.126
R3772 vdd2.n88 vdd2.t1226 8.126
R3773 vdd2.n89 vdd2.t424 8.126
R3774 vdd2.n89 vdd2.t1338 8.126
R3775 vdd2.n90 vdd2.t990 8.126
R3776 vdd2.n90 vdd2.t415 8.126
R3777 vdd2.n91 vdd2.t56 8.126
R3778 vdd2.n91 vdd2.t981 8.126
R3779 vdd2.n92 vdd2.t1259 8.126
R3780 vdd2.n92 vdd2.t684 8.126
R3781 vdd2.n93 vdd2.t1021 8.126
R3782 vdd2.n93 vdd2.t451 8.126
R3783 vdd2.n94 vdd2.t90 8.126
R3784 vdd2.n94 vdd2.t1012 8.126
R3785 vdd2.n95 vdd2.t659 8.126
R3786 vdd2.n95 vdd2.t82 8.126
R3787 vdd2.n96 vdd2.t430 8.126
R3788 vdd2.n96 vdd2.t1343 8.126
R3789 vdd2.n98 vdd2.t1209 8.126
R3790 vdd2.n98 vdd2.t625 8.126
R3791 vdd2.n99 vdd2.t1485 8.126
R3792 vdd2.n99 vdd2.t906 8.126
R3793 vdd2.n100 vdd2.t100 8.126
R3794 vdd2.n100 vdd2.t1024 8.126
R3795 vdd2.n101 vdd2.t669 8.126
R3796 vdd2.n101 vdd2.t95 8.126
R3797 vdd2.n102 vdd2.t1239 8.126
R3798 vdd2.n102 vdd2.t657 8.126
R3799 vdd2.n103 vdd2.t957 8.126
R3800 vdd2.n103 vdd2.t379 8.126
R3801 vdd2.n104 vdd2.t708 8.126
R3802 vdd2.n104 vdd2.t130 8.126
R3803 vdd2.n105 vdd2.t1277 8.126
R3804 vdd2.n105 vdd2.t698 8.126
R3805 vdd2.n106 vdd2.t353 8.126
R3806 vdd2.n106 vdd2.t1271 8.126
R3807 vdd2.n107 vdd2.t105 8.126
R3808 vdd2.n107 vdd2.t1028 8.126
R3809 vdd2.n109 vdd2.t861 8.126
R3810 vdd2.n109 vdd2.t286 8.126
R3811 vdd2.n110 vdd2.t1143 8.126
R3812 vdd2.n110 vdd2.t561 8.126
R3813 vdd2.n111 vdd2.t1256 8.126
R3814 vdd2.n111 vdd2.t678 8.126
R3815 vdd2.n112 vdd2.t330 8.126
R3816 vdd2.n112 vdd2.t1250 8.126
R3817 vdd2.n113 vdd2.t891 8.126
R3818 vdd2.n113 vdd2.t323 8.126
R3819 vdd2.n114 vdd2.t607 8.126
R3820 vdd2.n114 vdd2.t38 8.126
R3821 vdd2.n115 vdd2.t371 8.126
R3822 vdd2.n115 vdd2.t1287 8.126
R3823 vdd2.n116 vdd2.t938 8.126
R3824 vdd2.n116 vdd2.t358 8.126
R3825 vdd2.n117 vdd2.t9 8.126
R3826 vdd2.n117 vdd2.t926 8.126
R3827 vdd2.n118 vdd2.t1264 8.126
R3828 vdd2.n118 vdd2.t686 8.126
R3829 vdd2.n120 vdd2.t1397 8.126
R3830 vdd2.n120 vdd2.t1431 8.126
R3831 vdd2.n121 vdd2.t187 8.126
R3832 vdd2.n121 vdd2.t218 8.126
R3833 vdd2.n122 vdd2.t315 8.126
R3834 vdd2.n122 vdd2.t340 8.126
R3835 vdd2.n123 vdd2.t877 8.126
R3836 vdd2.n123 vdd2.t902 8.126
R3837 vdd2.n124 vdd2.t1435 8.126
R3838 vdd2.n124 vdd2.t1470 8.126
R3839 vdd2.n125 vdd2.t1158 8.126
R3840 vdd2.n125 vdd2.t1189 8.126
R3841 vdd2.n126 vdd2.t914 8.126
R3842 vdd2.n126 vdd2.t948 8.126
R3843 vdd2.n127 vdd2.t1482 8.126
R3844 vdd2.n127 vdd2.t19 8.126
R3845 vdd2.n128 vdd2.t551 8.126
R3846 vdd2.n128 vdd2.t582 8.126
R3847 vdd2.n129 vdd2.t322 8.126
R3848 vdd2.n129 vdd2.t347 8.126
R3849 vdd2.n131 vdd2.t1050 8.126
R3850 vdd2.n131 vdd2.t476 8.126
R3851 vdd2.n132 vdd2.t1336 8.126
R3852 vdd2.n132 vdd2.t759 8.126
R3853 vdd2.n133 vdd2.t1459 8.126
R3854 vdd2.n133 vdd2.t884 8.126
R3855 vdd2.n134 vdd2.t526 8.126
R3856 vdd2.n134 vdd2.t1451 8.126
R3857 vdd2.n135 vdd2.t1095 8.126
R3858 vdd2.n135 vdd2.t512 8.126
R3859 vdd2.n136 vdd2.t802 8.126
R3860 vdd2.n136 vdd2.t232 8.126
R3861 vdd2.n137 vdd2.t571 8.126
R3862 vdd2.n137 vdd2.t1495 8.126
R3863 vdd2.n138 vdd2.t1142 8.126
R3864 vdd2.n138 vdd2.t559 8.126
R3865 vdd2.n139 vdd2.t206 8.126
R3866 vdd2.n139 vdd2.t1133 8.126
R3867 vdd2.n140 vdd2.t1467 8.126
R3868 vdd2.n140 vdd2.t890 8.126
R3869 vdd2.n142 vdd2.t704 8.126
R3870 vdd2.n142 vdd2.t126 8.126
R3871 vdd2.n143 vdd2.t997 8.126
R3872 vdd2.n143 vdd2.t423 8.126
R3873 vdd2.n144 vdd2.t1120 8.126
R3874 vdd2.n144 vdd2.t538 8.126
R3875 vdd2.n145 vdd2.t182 8.126
R3876 vdd2.n145 vdd2.t1109 8.126
R3877 vdd2.n146 vdd2.t746 8.126
R3878 vdd2.n146 vdd2.t171 8.126
R3879 vdd2.n147 vdd2.t458 8.126
R3880 vdd2.n147 vdd2.t1378 8.126
R3881 vdd2.n148 vdd2.t226 8.126
R3882 vdd2.n148 vdd2.t1149 8.126
R3883 vdd2.n149 vdd2.t790 8.126
R3884 vdd2.n149 vdd2.t214 8.126
R3885 vdd2.n150 vdd2.t1354 8.126
R3886 vdd2.n150 vdd2.t780 8.126
R3887 vdd2.n151 vdd2.t1126 8.126
R3888 vdd2.n151 vdd2.t544 8.126
R3889 vdd2.n153 vdd2.t1035 8.126
R3890 vdd2.n153 vdd2.t464 8.126
R3891 vdd2.n154 vdd2.t1321 8.126
R3892 vdd2.n154 vdd2.t749 8.126
R3893 vdd2.n155 vdd2.t1447 8.126
R3894 vdd2.n155 vdd2.t872 8.126
R3895 vdd2.n156 vdd2.t514 8.126
R3896 vdd2.n156 vdd2.t1436 8.126
R3897 vdd2.n157 vdd2.t1075 8.126
R3898 vdd2.n157 vdd2.t498 8.126
R3899 vdd2.n158 vdd2.t795 8.126
R3900 vdd2.n158 vdd2.t221 8.126
R3901 vdd2.n159 vdd2.t555 8.126
R3902 vdd2.n159 vdd2.t1479 8.126
R3903 vdd2.n160 vdd2.t1130 8.126
R3904 vdd2.n160 vdd2.t548 8.126
R3905 vdd2.n161 vdd2.t193 8.126
R3906 vdd2.n161 vdd2.t1121 8.126
R3907 vdd2.n162 vdd2.t1454 8.126
R3908 vdd2.n162 vdd2.t879 8.126
R3909 vdd2.n164 vdd2.t693 8.126
R3910 vdd2.n164 vdd2.t113 8.126
R3911 vdd2.n165 vdd2.t985 8.126
R3912 vdd2.n165 vdd2.t410 8.126
R3913 vdd2.n166 vdd2.t1105 8.126
R3914 vdd2.n166 vdd2.t523 8.126
R3915 vdd2.n167 vdd2.t172 8.126
R3916 vdd2.n167 vdd2.t1096 8.126
R3917 vdd2.n168 vdd2.t731 8.126
R3918 vdd2.n168 vdd2.t155 8.126
R3919 vdd2.n169 vdd2.t448 8.126
R3920 vdd2.n169 vdd2.t1366 8.126
R3921 vdd2.n170 vdd2.t210 8.126
R3922 vdd2.n170 vdd2.t1136 8.126
R3923 vdd2.n171 vdd2.t775 8.126
R3924 vdd2.n171 vdd2.t201 8.126
R3925 vdd2.n172 vdd2.t1341 8.126
R3926 vdd2.n172 vdd2.t766 8.126
R3927 vdd2.n173 vdd2.t1113 8.126
R3928 vdd2.n173 vdd2.t530 8.126
R3929 vdd2.n175 vdd2.t1247 8.126
R3930 vdd2.n175 vdd2.t1270 8.126
R3931 vdd2.n176 vdd2.t35 8.126
R3932 vdd2.n176 vdd2.t59 8.126
R3933 vdd2.n177 vdd2.t144 8.126
R3934 vdd2.n177 vdd2.t178 8.126
R3935 vdd2.n178 vdd2.t713 8.126
R3936 vdd2.n178 vdd2.t747 8.126
R3937 vdd2.n179 vdd2.t1274 8.126
R3938 vdd2.n179 vdd2.t1305 8.126
R3939 vdd2.n180 vdd2.t1000 8.126
R3940 vdd2.n180 vdd2.t1018 8.126
R3941 vdd2.n181 vdd2.t755 8.126
R3942 vdd2.n181 vdd2.t784 8.126
R3943 vdd2.n182 vdd2.t1320 8.126
R3944 vdd2.n182 vdd2.t1350 8.126
R3945 vdd2.n183 vdd2.t400 8.126
R3946 vdd2.n183 vdd2.t428 8.126
R3947 vdd2.n184 vdd2.t153 8.126
R3948 vdd2.n184 vdd2.t186 8.126
R3949 vdd2.n186 vdd2.t895 8.126
R3950 vdd2.n186 vdd2.t328 8.126
R3951 vdd2.n187 vdd2.t1184 8.126
R3952 vdd2.n187 vdd2.t606 8.126
R3953 vdd2.n188 vdd2.t1297 8.126
R3954 vdd2.n188 vdd2.t724 8.126
R3955 vdd2.n189 vdd2.t375 8.126
R3956 vdd2.n189 vdd2.t1290 8.126
R3957 vdd2.n190 vdd2.t932 8.126
R3958 vdd2.n190 vdd2.t356 8.126
R3959 vdd2.n191 vdd2.t646 8.126
R3960 vdd2.n191 vdd2.t74 8.126
R3961 vdd2.n192 vdd2.t416 8.126
R3962 vdd2.n192 vdd2.t1327 8.126
R3963 vdd2.n193 vdd2.t984 8.126
R3964 vdd2.n193 vdd2.t409 8.126
R3965 vdd2.n194 vdd2.t50 8.126
R3966 vdd2.n194 vdd2.t976 8.126
R3967 vdd2.n195 vdd2.t1303 8.126
R3968 vdd2.n195 vdd2.t730 8.126
R3969 vdd2.n197 vdd2.t550 8.126
R3970 vdd2.n197 vdd2.t1474 8.126
R3971 vdd2.n198 vdd2.t836 8.126
R3972 vdd2.n198 vdd2.t263 8.126
R3973 vdd2.n199 vdd2.t960 8.126
R3974 vdd2.n199 vdd2.t384 8.126
R3975 vdd2.n200 vdd2.t33 8.126
R3976 vdd2.n200 vdd2.t953 8.126
R3977 vdd2.n201 vdd2.t589 8.126
R3978 vdd2.n201 vdd2.t15 8.126
R3979 vdd2.n202 vdd2.t308 8.126
R3980 vdd2.n202 vdd2.t1229 8.126
R3981 vdd2.n203 vdd2.t65 8.126
R3982 vdd2.n203 vdd2.t992 8.126
R3983 vdd2.n204 vdd2.t629 8.126
R3984 vdd2.n204 vdd2.t58 8.126
R3985 vdd2.n205 vdd2.t1206 8.126
R3986 vdd2.n205 vdd2.t623 8.126
R3987 vdd2.n206 vdd2.t967 8.126
R3988 vdd2.n206 vdd2.t390 8.126
R3989 vdd2.n208 vdd2.t241 8.126
R3990 vdd2.n208 vdd2.t1167 8.126
R3991 vdd2.n209 vdd2.t522 8.126
R3992 vdd2.n209 vdd2.t1445 8.126
R3993 vdd2.n210 vdd2.t643 8.126
R3994 vdd2.n210 vdd2.t69 8.126
R3995 vdd2.n211 vdd2.t1218 8.126
R3996 vdd2.n211 vdd2.t632 8.126
R3997 vdd2.n212 vdd2.t283 8.126
R3998 vdd2.n212 vdd2.t1204 8.126
R3999 vdd2.n213 vdd2.t1492 8.126
R4000 vdd2.n213 vdd2.t912 8.126
R4001 vdd2.n214 vdd2.t1251 8.126
R4002 vdd2.n214 vdd2.t670 8.126
R4003 vdd2.n215 vdd2.t326 8.126
R4004 vdd2.n215 vdd2.t1245 8.126
R4005 vdd2.n216 vdd2.t887 8.126
R4006 vdd2.n216 vdd2.t319 8.126
R4007 vdd2.n217 vdd2.t650 8.126
R4008 vdd2.n217 vdd2.t77 8.126
R4009 vdd2.n219 vdd2.t1389 8.126
R4010 vdd2.n219 vdd2.t817 8.126
R4011 vdd2.n220 vdd2.t176 8.126
R4012 vdd2.n220 vdd2.t1102 8.126
R4013 vdd2.n221 vdd2.t307 8.126
R4014 vdd2.n221 vdd2.t1227 8.126
R4015 vdd2.n222 vdd2.t870 8.126
R4016 vdd2.n222 vdd2.t300 8.126
R4017 vdd2.n223 vdd2.t1428 8.126
R4018 vdd2.n223 vdd2.t858 8.126
R4019 vdd2.n224 vdd2.t1147 8.126
R4020 vdd2.n224 vdd2.t565 8.126
R4021 vdd2.n225 vdd2.t903 8.126
R4022 vdd2.n225 vdd2.t331 8.126
R4023 vdd2.n226 vdd2.t1473 8.126
R4024 vdd2.n226 vdd2.t896 8.126
R4025 vdd2.n227 vdd2.t542 8.126
R4026 vdd2.n227 vdd2.t1465 8.126
R4027 vdd2.n228 vdd2.t313 8.126
R4028 vdd2.n228 vdd2.t1234 8.126
R4029 vdd2.n230 vdd2.t443 8.126
R4030 vdd2.n230 vdd2.t1358 8.126
R4031 vdd2.n231 vdd2.t722 8.126
R4032 vdd2.n231 vdd2.t142 8.126
R4033 vdd2.n232 vdd2.t850 8.126
R4034 vdd2.n232 vdd2.t275 8.126
R4035 vdd2.n233 vdd2.t1410 8.126
R4036 vdd2.n233 vdd2.t839 8.126
R4037 vdd2.n234 vdd2.t472 8.126
R4038 vdd2.n234 vdd2.t1394 8.126
R4039 vdd2.n235 vdd2.t192 8.126
R4040 vdd2.n235 vdd2.t1118 8.126
R4041 vdd2.n236 vdd2.t1452 8.126
R4042 vdd2.n236 vdd2.t878 8.126
R4043 vdd2.n237 vdd2.t520 8.126
R4044 vdd2.n237 vdd2.t1443 8.126
R4045 vdd2.n238 vdd2.t1091 8.126
R4046 vdd2.n238 vdd2.t509 8.126
R4047 vdd2.n239 vdd2.t856 8.126
R4048 vdd2.n239 vdd2.t282 8.126
R4049 vdd2.n241 vdd2.t88 8.126
R4050 vdd2.n241 vdd2.t1013 8.126
R4051 vdd2.n242 vdd2.t383 8.126
R4052 vdd2.n242 vdd2.t1296 8.126
R4053 vdd2.n243 vdd2.t496 8.126
R4054 vdd2.n243 vdd2.t1421 8.126
R4055 vdd2.n244 vdd2.t1064 8.126
R4056 vdd2.n244 vdd2.t487 8.126
R4057 vdd2.n245 vdd2.t124 8.126
R4058 vdd2.n245 vdd2.t1047 8.126
R4059 vdd2.n246 vdd2.t1340 8.126
R4060 vdd2.n246 vdd2.t765 8.126
R4061 vdd2.n247 vdd2.t1110 8.126
R4062 vdd2.n247 vdd2.t528 8.126
R4063 vdd2.n248 vdd2.t174 8.126
R4064 vdd2.n248 vdd2.t1101 8.126
R4065 vdd2.n249 vdd2.t741 8.126
R4066 vdd2.n249 vdd2.t168 8.126
R4067 vdd2.n250 vdd2.t503 8.126
R4068 vdd2.n250 vdd2.t1426 8.126
R4069 vdd2.n252 vdd2.t637 8.126
R4070 vdd2.n252 vdd2.t664 8.126
R4071 vdd2.n253 vdd2.t924 8.126
R4072 vdd2.n253 vdd2.t958 8.126
R4073 vdd2.n254 vdd2.t1039 8.126
R4074 vdd2.n254 vdd2.t1073 8.126
R4075 vdd2.n255 vdd2.t107 8.126
R4076 vdd2.n255 vdd2.t139 8.126
R4077 vdd2.n256 vdd2.t672 8.126
R4078 vdd2.n256 vdd2.t701 8.126
R4079 vdd2.n257 vdd2.t398 8.126
R4080 vdd2.n257 vdd2.t427 8.126
R4081 vdd2.n258 vdd2.t150 8.126
R4082 vdd2.n258 vdd2.t184 8.126
R4083 vdd2.n259 vdd2.t720 8.126
R4084 vdd2.n259 vdd2.t751 8.126
R4085 vdd2.n260 vdd2.t1285 8.126
R4086 vdd2.n260 vdd2.t1316 8.126
R4087 vdd2.n261 vdd2.t1044 8.126
R4088 vdd2.n261 vdd2.t1079 8.126
R4089 vdd2.n263 vdd2.t937 8.126
R4090 vdd2.n263 vdd2.t360 8.126
R4091 vdd2.n264 vdd2.t1225 8.126
R4092 vdd2.n264 vdd2.t640 8.126
R4093 vdd2.n265 vdd2.t1337 8.126
R4094 vdd2.n265 vdd2.t760 8.126
R4095 vdd2.n266 vdd2.t414 8.126
R4096 vdd2.n266 vdd2.t1324 8.126
R4097 vdd2.n267 vdd2.t982 8.126
R4098 vdd2.n267 vdd2.t403 8.126
R4099 vdd2.n268 vdd2.t683 8.126
R4100 vdd2.n268 vdd2.t103 8.126
R4101 vdd2.n269 vdd2.t450 8.126
R4102 vdd2.n269 vdd2.t1368 8.126
R4103 vdd2.n270 vdd2.t1011 8.126
R4104 vdd2.n270 vdd2.t444 8.126
R4105 vdd2.n271 vdd2.t84 8.126
R4106 vdd2.n271 vdd2.t1009 8.126
R4107 vdd2.n272 vdd2.t1344 8.126
R4108 vdd2.n272 vdd2.t769 8.126
R4109 vdd2.n274 vdd2.t593 8.126
R4110 vdd2.n274 vdd2.t21 8.126
R4111 vdd2.n275 vdd2.t876 8.126
R4112 vdd2.n275 vdd2.t305 8.126
R4113 vdd2.n276 vdd2.t999 8.126
R4114 vdd2.n276 vdd2.t425 8.126
R4115 vdd2.n277 vdd2.t64 8.126
R4116 vdd2.n277 vdd2.t991 8.126
R4117 vdd2.n278 vdd2.t628 8.126
R4118 vdd2.n278 vdd2.t55 8.126
R4119 vdd2.n279 vdd2.t342 8.126
R4120 vdd2.n279 vdd2.t1260 8.126
R4121 vdd2.n280 vdd2.t97 8.126
R4122 vdd2.n280 vdd2.t1020 8.126
R4123 vdd2.n281 vdd2.t666 8.126
R4124 vdd2.n281 vdd2.t89 8.126
R4125 vdd2.n282 vdd2.t1242 8.126
R4126 vdd2.n282 vdd2.t660 8.126
R4127 vdd2.n283 vdd2.t1003 8.126
R4128 vdd2.n283 vdd2.t431 8.126
R4129 vdd2.n285 vdd2.t1140 8.126
R4130 vdd2.n285 vdd2.t560 8.126
R4131 vdd2.n286 vdd2.t1420 8.126
R4132 vdd2.n286 vdd2.t848 8.126
R4133 vdd2.n287 vdd2.t47 8.126
R4134 vdd2.n287 vdd2.t971 8.126
R4135 vdd2.n288 vdd2.t611 8.126
R4136 vdd2.n288 vdd2.t39 8.126
R4137 vdd2.n289 vdd2.t1178 8.126
R4138 vdd2.n289 vdd2.t598 8.126
R4139 vdd2.n290 vdd2.t886 8.126
R4140 vdd2.n290 vdd2.t317 8.126
R4141 vdd2.n291 vdd2.t647 8.126
R4142 vdd2.n291 vdd2.t75 8.126
R4143 vdd2.n292 vdd2.t1223 8.126
R4144 vdd2.n292 vdd2.t639 8.126
R4145 vdd2.n293 vdd2.t296 8.126
R4146 vdd2.n293 vdd2.t1215 8.126
R4147 vdd2.n294 vdd2.t54 8.126
R4148 vdd2.n294 vdd2.t980 8.126
R4149 vdd2.n296 vdd2.t791 8.126
R4150 vdd2.n296 vdd2.t216 8.126
R4151 vdd2.n297 vdd2.t1071 8.126
R4152 vdd2.n297 vdd2.t494 8.126
R4153 vdd2.n298 vdd2.t1203 8.126
R4154 vdd2.n298 vdd2.t621 8.126
R4155 vdd2.n299 vdd2.t271 8.126
R4156 vdd2.n299 vdd2.t1195 8.126
R4157 vdd2.n300 vdd2.t830 8.126
R4158 vdd2.n300 vdd2.t256 8.126
R4159 vdd2.n301 vdd2.t541 8.126
R4160 vdd2.n301 vdd2.t1464 8.126
R4161 vdd2.n302 vdd2.t311 8.126
R4162 vdd2.n302 vdd2.t1231 8.126
R4163 vdd2.n303 vdd2.t875 8.126
R4164 vdd2.n303 vdd2.t303 8.126
R4165 vdd2.n304 vdd2.t1438 8.126
R4166 vdd2.n304 vdd2.t866 8.126
R4167 vdd2.n305 vdd2.t1210 8.126
R4168 vdd2.n305 vdd2.t626 8.126
R4169 vdd2.n307 vdd2.t1332 8.126
R4170 vdd2.n307 vdd2.t1362 8.126
R4171 vdd2.n308 vdd2.t115 8.126
R4172 vdd2.n308 vdd2.t147 8.126
R4173 vdd2.n309 vdd2.t246 8.126
R4174 vdd2.n309 vdd2.t281 8.126
R4175 vdd2.n310 vdd2.t808 8.126
R4176 vdd2.n310 vdd2.t846 8.126
R4177 vdd2.n311 vdd2.t1370 8.126
R4178 vdd2.n311 vdd2.t1399 8.126
R4179 vdd2.n312 vdd2.t1088 8.126
R4180 vdd2.n312 vdd2.t1124 8.126
R4181 vdd2.n313 vdd2.t853 8.126
R4182 vdd2.n313 vdd2.t882 8.126
R4183 vdd2.n314 vdd2.t1418 8.126
R4184 vdd2.n314 vdd2.t1449 8.126
R4185 vdd2.n315 vdd2.t483 8.126
R4186 vdd2.n315 vdd2.t515 8.126
R4187 vdd2.n316 vdd2.t254 8.126
R4188 vdd2.n316 vdd2.t287 8.126
R4189 vdd2.n318 vdd2.t127 8.126
R4190 vdd2.n318 vdd2.t1051 8.126
R4191 vdd2.n319 vdd2.t422 8.126
R4192 vdd2.n319 vdd2.t1335 8.126
R4193 vdd2.n320 vdd2.t537 8.126
R4194 vdd2.n320 vdd2.t1460 8.126
R4195 vdd2.n321 vdd2.t1108 8.126
R4196 vdd2.n321 vdd2.t527 8.126
R4197 vdd2.n322 vdd2.t170 8.126
R4198 vdd2.n322 vdd2.t1094 8.126
R4199 vdd2.n323 vdd2.t1377 8.126
R4200 vdd2.n323 vdd2.t804 8.126
R4201 vdd2.n324 vdd2.t1151 8.126
R4202 vdd2.n324 vdd2.t570 8.126
R4203 vdd2.n325 vdd2.t213 8.126
R4204 vdd2.n325 vdd2.t1141 8.126
R4205 vdd2.n326 vdd2.t781 8.126
R4206 vdd2.n326 vdd2.t207 8.126
R4207 vdd2.n327 vdd2.t545 8.126
R4208 vdd2.n327 vdd2.t1468 8.126
R4209 vdd2.n329 vdd2.t675 8.126
R4210 vdd2.n329 vdd2.t705 8.126
R4211 vdd2.n330 vdd2.t968 8.126
R4212 vdd2.n330 vdd2.t998 8.126
R4213 vdd2.n331 vdd2.t1082 8.126
R4214 vdd2.n331 vdd2.t1119 8.126
R4215 vdd2.n332 vdd2.t148 8.126
R4216 vdd2.n332 vdd2.t181 8.126
R4217 vdd2.n333 vdd2.t710 8.126
R4218 vdd2.n333 vdd2.t745 8.126
R4219 vdd2.n334 vdd2.t435 8.126
R4220 vdd2.n334 vdd2.t457 8.126
R4221 vdd2.n335 vdd2.t194 8.126
R4222 vdd2.n335 vdd2.t225 8.126
R4223 vdd2.n336 vdd2.t758 8.126
R4224 vdd2.n336 vdd2.t789 8.126
R4225 vdd2.n337 vdd2.t1323 8.126
R4226 vdd2.n337 vdd2.t1355 8.126
R4227 vdd2.n338 vdd2.t1093 8.126
R4228 vdd2.n338 vdd2.t1127 8.126
R4229 vdd2.n340 vdd2.t338 8.126
R4230 vdd2.n340 vdd2.t1255 8.126
R4231 vdd2.n341 vdd2.t620 8.126
R4232 vdd2.n341 vdd2.t45 8.126
R4233 vdd2.n342 vdd2.t737 8.126
R4234 vdd2.n342 vdd2.t161 8.126
R4235 vdd2.n343 vdd2.t1300 8.126
R4236 vdd2.n343 vdd2.t726 8.126
R4237 vdd2.n344 vdd2.t374 8.126
R4238 vdd2.n344 vdd2.t1289 8.126
R4239 vdd2.n345 vdd2.t81 8.126
R4240 vdd2.n345 vdd2.t1008 8.126
R4241 vdd2.n346 vdd2.t1342 8.126
R4242 vdd2.n346 vdd2.t767 8.126
R4243 vdd2.n347 vdd2.t420 8.126
R4244 vdd2.n347 vdd2.t1333 8.126
R4245 vdd2.n348 vdd2.t989 8.126
R4246 vdd2.n348 vdd2.t413 8.126
R4247 vdd2.n349 vdd2.t744 8.126
R4248 vdd2.n349 vdd2.t169 8.126
R4249 vdd2.n351 vdd2.t1490 8.126
R4250 vdd2.n351 vdd2.t909 8.126
R4251 vdd2.n352 vdd2.t279 8.126
R4252 vdd2.n352 vdd2.t1201 8.126
R4253 vdd2.n353 vdd2.t396 8.126
R4254 vdd2.n353 vdd2.t1311 8.126
R4255 vdd2.n354 vdd2.t963 8.126
R4256 vdd2.n354 vdd2.t387 8.126
R4257 vdd2.n355 vdd2.t32 8.126
R4258 vdd2.n355 vdd2.t952 8.126
R4259 vdd2.n356 vdd2.t1240 8.126
R4260 vdd2.n356 vdd2.t658 8.126
R4261 vdd2.n357 vdd2.t1002 8.126
R4262 vdd2.n357 vdd2.t429 8.126
R4263 vdd2.n358 vdd2.t73 8.126
R4264 vdd2.n358 vdd2.t995 8.126
R4265 vdd2.n359 vdd2.t635 8.126
R4266 vdd2.n359 vdd2.t63 8.126
R4267 vdd2.n360 vdd2.t407 8.126
R4268 vdd2.n360 vdd2.t1319 8.126
R4269 vdd2.n362 vdd2.t535 8.126
R4270 vdd2.n362 vdd2.t1458 8.126
R4271 vdd2.n363 vdd2.t819 8.126
R4272 vdd2.n363 vdd2.t242 8.126
R4273 vdd2.n364 vdd2.t941 8.126
R4274 vdd2.n364 vdd2.t364 8.126
R4275 vdd2.n365 vdd2.t11 8.126
R4276 vdd2.n365 vdd2.t929 8.126
R4277 vdd2.n366 vdd2.t574 8.126
R4278 vdd2.n366 vdd2.t1498 8.126
R4279 vdd2.n367 vdd2.t294 8.126
R4280 vdd2.n367 vdd2.t1214 8.126
R4281 vdd2.n368 vdd2.t52 8.126
R4282 vdd2.n368 vdd2.t979 8.126
R4283 vdd2.n369 vdd2.t616 8.126
R4284 vdd2.n369 vdd2.t44 8.126
R4285 vdd2.n370 vdd2.t1190 8.126
R4286 vdd2.n370 vdd2.t609 8.126
R4287 vdd2.n371 vdd2.t950 8.126
R4288 vdd2.n371 vdd2.t372 8.126
R4289 vdd2.n373 vdd2.t832 8.126
R4290 vdd2.n373 vdd2.t259 8.126
R4291 vdd2.n374 vdd2.t1117 8.126
R4292 vdd2.n374 vdd2.t536 8.126
R4293 vdd2.n375 vdd2.t1237 8.126
R4294 vdd2.n375 vdd2.t654 8.126
R4295 vdd2.n376 vdd2.t309 8.126
R4296 vdd2.n376 vdd2.t1230 8.126
R4297 vdd2.n377 vdd2.t869 8.126
R4298 vdd2.n377 vdd2.t299 8.126
R4299 vdd2.n378 vdd2.t581 8.126
R4300 vdd2.n378 vdd2.t7 8.126
R4301 vdd2.n379 vdd2.t345 8.126
R4302 vdd2.n379 vdd2.t1263 8.126
R4303 vdd2.n380 vdd2.t910 8.126
R4304 vdd2.n380 vdd2.t337 8.126
R4305 vdd2.n381 vdd2.t1480 8.126
R4306 vdd2.n381 vdd2.t900 8.126
R4307 vdd2.n382 vdd2.t1243 8.126
R4308 vdd2.n382 vdd2.t661 8.126
R4309 vdd2.n384 vdd2.t1373 8.126
R4310 vdd2.n384 vdd2.t1403 8.126
R4311 vdd2.n385 vdd2.t160 8.126
R4312 vdd2.n385 vdd2.t191 8.126
R4313 vdd2.n386 vdd2.t290 8.126
R4314 vdd2.n386 vdd2.t318 8.126
R4315 vdd2.n387 vdd2.t852 8.126
R4316 vdd2.n387 vdd2.t880 8.126
R4317 vdd2.n388 vdd2.t1408 8.126
R4318 vdd2.n388 vdd2.t1442 8.126
R4319 vdd2.n389 vdd2.t1132 8.126
R4320 vdd2.n389 vdd2.t1161 8.126
R4321 vdd2.n390 vdd2.t889 8.126
R4322 vdd2.n390 vdd2.t919 8.126
R4323 vdd2.n391 vdd2.t1456 8.126
R4324 vdd2.n391 vdd2.t1488 8.126
R4325 vdd2.n392 vdd2.t525 8.126
R4326 vdd2.n392 vdd2.t556 8.126
R4327 vdd2.n393 vdd2.t298 8.126
R4328 vdd2.n393 vdd2.t324 8.126
R4329 vdd2.n12 vdd2.t1026 8.126
R4330 vdd2.n12 vdd2.t454 8.126
R4331 vdd2.n13 vdd2.t1310 8.126
R4332 vdd2.n13 vdd2.t736 8.126
R4333 vdd2.n14 vdd2.t1432 8.126
R4334 vdd2.n14 vdd2.t862 8.126
R4335 vdd2.n15 vdd2.t499 8.126
R4336 vdd2.n15 vdd2.t1423 8.126
R4337 vdd2.n16 vdd2.t1062 8.126
R4338 vdd2.n16 vdd2.t486 8.126
R4339 vdd2.n17 vdd2.t779 8.126
R4340 vdd2.n17 vdd2.t205 8.126
R4341 vdd2.n18 vdd2.t543 8.126
R4342 vdd2.n18 vdd2.t1466 8.126
R4343 vdd2.n19 vdd2.t1116 8.126
R4344 vdd2.n19 vdd2.t532 8.126
R4345 vdd2.n20 vdd2.t180 8.126
R4346 vdd2.n20 vdd2.t1107 8.126
R4347 vdd2.n21 vdd2.t1441 8.126
R4348 vdd2.n21 vdd2.t868 8.126
R4349 vdd2.n396 vdd2.t681 8.126
R4350 vdd2.n396 vdd2.t102 8.126
R4351 vdd2.n397 vdd2.t975 8.126
R4352 vdd2.n397 vdd2.t395 8.126
R4353 vdd2.n398 vdd2.t1090 8.126
R4354 vdd2.n398 vdd2.t508 8.126
R4355 vdd2.n399 vdd2.t157 8.126
R4356 vdd2.n399 vdd2.t1076 8.126
R4357 vdd2.n400 vdd2.t718 8.126
R4358 vdd2.n400 vdd2.t137 8.126
R4359 vdd2.n401 vdd2.t439 8.126
R4360 vdd2.n401 vdd2.t1353 8.126
R4361 vdd2.n402 vdd2.t198 8.126
R4362 vdd2.n402 vdd2.t1125 8.126
R4363 vdd2.n403 vdd2.t763 8.126
R4364 vdd2.n403 vdd2.t189 8.126
R4365 vdd2.n404 vdd2.t1328 8.126
R4366 vdd2.n404 vdd2.t756 8.126
R4367 vdd2.n405 vdd2.t1098 8.126
R4368 vdd2.n405 vdd2.t519 8.126
R4369 vdd2.n407 vdd2.t380 8.126
R4370 vdd2.n407 vdd2.t1294 8.126
R4371 vdd2.n408 vdd2.t655 8.126
R4372 vdd2.n408 vdd2.t79 8.126
R4373 vdd2.n409 vdd2.t778 8.126
R4374 vdd2.n409 vdd2.t204 8.126
R4375 vdd2.n410 vdd2.t1347 8.126
R4376 vdd2.n410 vdd2.t772 8.126
R4377 vdd2.n411 vdd2.t418 8.126
R4378 vdd2.n411 vdd2.t1331 8.126
R4379 vdd2.n412 vdd2.t118 8.126
R4380 vdd2.n412 vdd2.t1042 8.126
R4381 vdd2.n413 vdd2.t1384 8.126
R4382 vdd2.n413 vdd2.t809 8.126
R4383 vdd2.n414 vdd2.t455 8.126
R4384 vdd2.n414 vdd2.t1375 8.126
R4385 vdd2.n415 vdd2.t1019 8.126
R4386 vdd2.n415 vdd2.t449 8.126
R4387 vdd2.n416 vdd2.t785 8.126
R4388 vdd2.n416 vdd2.t211 8.126
R4389 vdd2.n418 vdd2.t665 8.126
R4390 vdd2.n418 vdd2.t91 8.126
R4391 vdd2.n419 vdd2.t959 8.126
R4392 vdd2.n419 vdd2.t382 8.126
R4393 vdd2.n420 vdd2.t1072 8.126
R4394 vdd2.n420 vdd2.t495 8.126
R4395 vdd2.n421 vdd2.t138 8.126
R4396 vdd2.n421 vdd2.t1063 8.126
R4397 vdd2.n422 vdd2.t700 8.126
R4398 vdd2.n422 vdd2.t123 8.126
R4399 vdd2.n423 vdd2.t426 8.126
R4400 vdd2.n423 vdd2.t1339 8.126
R4401 vdd2.n424 vdd2.t183 8.126
R4402 vdd2.n424 vdd2.t1111 8.126
R4403 vdd2.n425 vdd2.t750 8.126
R4404 vdd2.n425 vdd2.t175 8.126
R4405 vdd2.n426 vdd2.t1317 8.126
R4406 vdd2.n426 vdd2.t742 8.126
R4407 vdd2.n427 vdd2.t1080 8.126
R4408 vdd2.n427 vdd2.t504 8.126
R4409 vdd2.n444 vdd2.t1224 8.126
R4410 vdd2.n444 vdd2.t638 8.126
R4411 vdd2.n445 vdd2.t5 8.126
R4412 vdd2.n445 vdd2.t923 8.126
R4413 vdd2.n446 vdd2.t117 8.126
R4414 vdd2.n446 vdd2.t1038 8.126
R4415 vdd2.n447 vdd2.t688 8.126
R4416 vdd2.n447 vdd2.t106 8.126
R4417 vdd2.n448 vdd2.t1253 8.126
R4418 vdd2.n448 vdd2.t673 8.126
R4419 vdd2.n449 vdd2.t977 8.126
R4420 vdd2.n449 vdd2.t397 8.126
R4421 vdd2.n450 vdd2.t727 8.126
R4422 vdd2.n450 vdd2.t149 8.126
R4423 vdd2.n451 vdd2.t1295 8.126
R4424 vdd2.n451 vdd2.t719 8.126
R4425 vdd2.n452 vdd2.t370 8.126
R4426 vdd2.n452 vdd2.t1286 8.126
R4427 vdd2.n453 vdd2.t121 8.126
R4428 vdd2.n453 vdd2.t1046 8.126
R4429 vdd2.n456 vdd2.t873 8.126
R4430 vdd2.n456 vdd2.t304 8.126
R4431 vdd2.n457 vdd2.t1160 8.126
R4432 vdd2.n457 vdd2.t580 8.126
R4433 vdd2.n458 vdd2.t1273 8.126
R4434 vdd2.n458 vdd2.t695 8.126
R4435 vdd2.n459 vdd2.t349 8.126
R4436 vdd2.n459 vdd2.t1266 8.126
R4437 vdd2.n460 vdd2.t905 8.126
R4438 vdd2.n460 vdd2.t335 8.126
R4439 vdd2.n461 vdd2.t622 8.126
R4440 vdd2.n461 vdd2.t49 8.126
R4441 vdd2.n462 vdd2.t388 8.126
R4442 vdd2.n462 vdd2.t1301 8.126
R4443 vdd2.n463 vdd2.t956 8.126
R4444 vdd2.n463 vdd2.t381 8.126
R4445 vdd2.n464 vdd2.t28 8.126
R4446 vdd2.n464 vdd2.t946 8.126
R4447 vdd2.n465 vdd2.t1279 8.126
R4448 vdd2.n465 vdd2.t699 8.126
R4449 vdd2.n467 vdd2.t1419 8.126
R4450 vdd2.n467 vdd2.t1450 8.126
R4451 vdd2.n468 vdd2.t202 8.126
R4452 vdd2.n468 vdd2.t234 8.126
R4453 vdd2.n469 vdd2.t329 8.126
R4454 vdd2.n469 vdd2.t355 8.126
R4455 vdd2.n470 vdd2.t892 8.126
R4456 vdd2.n470 vdd2.t922 8.126
R4457 vdd2.n471 vdd2.t1455 8.126
R4458 vdd2.n471 vdd2.t1484 8.126
R4459 vdd2.n472 vdd2.t1175 8.126
R4460 vdd2.n472 vdd2.t1207 8.126
R4461 vdd2.n473 vdd2.t930 8.126
R4462 vdd2.n473 vdd2.t965 8.126
R4463 vdd2.n474 vdd2.t4 8.126
R4464 vdd2.n474 vdd2.t37 8.126
R4465 vdd2.n475 vdd2.t569 8.126
R4466 vdd2.n475 vdd2.t601 8.126
R4467 vdd2.n476 vdd2.t333 8.126
R4468 vdd2.n476 vdd2.t361 8.126
R4469 vdd2.n478 vdd2.t1068 8.126
R4470 vdd2.n478 vdd2.t493 8.126
R4471 vdd2.n479 vdd2.t1351 8.126
R4472 vdd2.n479 vdd2.t776 8.126
R4473 vdd2.n480 vdd2.t1477 8.126
R4474 vdd2.n480 vdd2.t899 8.126
R4475 vdd2.n481 vdd2.t547 8.126
R4476 vdd2.n481 vdd2.t1471 8.126
R4477 vdd2.n482 vdd2.t1114 8.126
R4478 vdd2.n482 vdd2.t531 8.126
R4479 vdd2.n483 vdd2.t823 8.126
R4480 vdd2.n483 vdd2.t250 8.126
R4481 vdd2.n484 vdd2.t586 8.126
R4482 vdd2.n484 vdd2.t13 8.126
R4483 vdd2.n485 vdd2.t1157 8.126
R4484 vdd2.n485 vdd2.t579 8.126
R4485 vdd2.n486 vdd2.t224 8.126
R4486 vdd2.n486 vdd2.t1148 8.126
R4487 vdd2.n487 vdd2.t1483 8.126
R4488 vdd2.n487 vdd2.t904 8.126
R4489 vdd2.n0 vdd2.t1361 8.126
R4490 vdd2.n0 vdd2.t792 8.126
R4491 vdd2.n1 vdd2.t146 8.126
R4492 vdd2.n1 vdd2.t1070 8.126
R4493 vdd2.n2 vdd2.t280 8.126
R4494 vdd2.n2 vdd2.t1202 8.126
R4495 vdd2.n3 vdd2.t845 8.126
R4496 vdd2.n3 vdd2.t270 8.126
R4497 vdd2.n4 vdd2.t1401 8.126
R4498 vdd2.n4 vdd2.t829 8.126
R4499 vdd2.n5 vdd2.t1123 8.126
R4500 vdd2.n5 vdd2.t540 8.126
R4501 vdd2.n6 vdd2.t881 8.126
R4502 vdd2.n6 vdd2.t310 8.126
R4503 vdd2.n7 vdd2.t1448 8.126
R4504 vdd2.n7 vdd2.t874 8.126
R4505 vdd2.n8 vdd2.t516 8.126
R4506 vdd2.n8 vdd2.t1440 8.126
R4507 vdd2.n9 vdd2.t289 8.126
R4508 vdd2.n9 vdd2.t1211 8.126
R4509 vdd2.n437 vdd2.n436 7.5
R4510 vdd2.n432 vdd2.n431 3.75
R4511 vdd2.n506 vdd2.n505 2.427
R4512 vdd2.n510 vdd2.n509 2.158
R4513 vdd2.n509 vdd2.n508 2.158
R4514 vdd2.n508 vdd2.n507 2.158
R4515 vdd2.n507 vdd2.n506 2.158
R4516 vdd2.n505 vdd2.n504 2.158
R4517 vdd2.n504 vdd2.n503 2.158
R4518 vdd2.n503 vdd2.n502 2.158
R4519 vdd2.n521 vdd2.n510 1.212
R4520 vdd2.n516 vdd2.n515 0.866
R4521 vdd2.n527 vdd2.n526 0.849
R4522 vdd2.n538 vdd2.n537 0.849
R4523 vdd2.n549 vdd2.n548 0.849
R4524 vdd2.n560 vdd2.n559 0.849
R4525 vdd2.n571 vdd2.n570 0.849
R4526 vdd2.n582 vdd2.n581 0.849
R4527 vdd2.n593 vdd2.n592 0.849
R4528 vdd2.n604 vdd2.n603 0.849
R4529 vdd2.n615 vdd2.n614 0.849
R4530 vdd2.n626 vdd2.n625 0.849
R4531 vdd2.n637 vdd2.n636 0.849
R4532 vdd2.n648 vdd2.n647 0.849
R4533 vdd2.n659 vdd2.n658 0.849
R4534 vdd2.n670 vdd2.n669 0.849
R4535 vdd2.n681 vdd2.n680 0.849
R4536 vdd2.n692 vdd2.n691 0.849
R4537 vdd2.n703 vdd2.n702 0.849
R4538 vdd2.n714 vdd2.n713 0.849
R4539 vdd2.n725 vdd2.n724 0.849
R4540 vdd2.n736 vdd2.n735 0.849
R4541 vdd2.n747 vdd2.n746 0.849
R4542 vdd2.n758 vdd2.n757 0.849
R4543 vdd2.n769 vdd2.n768 0.849
R4544 vdd2.n780 vdd2.n779 0.849
R4545 vdd2.n791 vdd2.n790 0.849
R4546 vdd2.n802 vdd2.n801 0.849
R4547 vdd2.n813 vdd2.n812 0.849
R4548 vdd2.n824 vdd2.n823 0.849
R4549 vdd2.n835 vdd2.n834 0.849
R4550 vdd2.n846 vdd2.n845 0.849
R4551 vdd2.n496 vdd2.n495 0.849
R4552 vdd2.n37 vdd2.n36 0.849
R4553 vdd2.n48 vdd2.n47 0.849
R4554 vdd2.n59 vdd2.n58 0.849
R4555 vdd2.n70 vdd2.n69 0.849
R4556 vdd2.n81 vdd2.n80 0.849
R4557 vdd2.n92 vdd2.n91 0.849
R4558 vdd2.n103 vdd2.n102 0.849
R4559 vdd2.n114 vdd2.n113 0.849
R4560 vdd2.n125 vdd2.n124 0.849
R4561 vdd2.n136 vdd2.n135 0.849
R4562 vdd2.n147 vdd2.n146 0.849
R4563 vdd2.n158 vdd2.n157 0.849
R4564 vdd2.n169 vdd2.n168 0.849
R4565 vdd2.n180 vdd2.n179 0.849
R4566 vdd2.n191 vdd2.n190 0.849
R4567 vdd2.n202 vdd2.n201 0.849
R4568 vdd2.n213 vdd2.n212 0.849
R4569 vdd2.n224 vdd2.n223 0.849
R4570 vdd2.n235 vdd2.n234 0.849
R4571 vdd2.n246 vdd2.n245 0.849
R4572 vdd2.n257 vdd2.n256 0.849
R4573 vdd2.n268 vdd2.n267 0.849
R4574 vdd2.n279 vdd2.n278 0.849
R4575 vdd2.n290 vdd2.n289 0.849
R4576 vdd2.n301 vdd2.n300 0.849
R4577 vdd2.n312 vdd2.n311 0.849
R4578 vdd2.n323 vdd2.n322 0.849
R4579 vdd2.n334 vdd2.n333 0.849
R4580 vdd2.n345 vdd2.n344 0.849
R4581 vdd2.n356 vdd2.n355 0.849
R4582 vdd2.n367 vdd2.n366 0.849
R4583 vdd2.n378 vdd2.n377 0.849
R4584 vdd2.n389 vdd2.n388 0.849
R4585 vdd2.n17 vdd2.n16 0.849
R4586 vdd2.n401 vdd2.n400 0.849
R4587 vdd2.n412 vdd2.n411 0.849
R4588 vdd2.n423 vdd2.n422 0.849
R4589 vdd2.n449 vdd2.n448 0.849
R4590 vdd2.n461 vdd2.n460 0.849
R4591 vdd2.n472 vdd2.n471 0.849
R4592 vdd2.n483 vdd2.n482 0.849
R4593 vdd2.n5 vdd2.n4 0.849
R4594 vdd2.n520 vdd2.n519 0.77
R4595 vdd2.n519 vdd2.n518 0.77
R4596 vdd2.n518 vdd2.n517 0.77
R4597 vdd2.n517 vdd2.n516 0.77
R4598 vdd2.n515 vdd2.n514 0.77
R4599 vdd2.n514 vdd2.n513 0.77
R4600 vdd2.n513 vdd2.n512 0.77
R4601 vdd2.n512 vdd2.n511 0.77
R4602 vdd2.n531 vdd2.n530 0.753
R4603 vdd2.n530 vdd2.n529 0.753
R4604 vdd2.n529 vdd2.n528 0.753
R4605 vdd2.n528 vdd2.n527 0.753
R4606 vdd2.n526 vdd2.n525 0.753
R4607 vdd2.n525 vdd2.n524 0.753
R4608 vdd2.n524 vdd2.n523 0.753
R4609 vdd2.n523 vdd2.n522 0.753
R4610 vdd2.n542 vdd2.n541 0.753
R4611 vdd2.n541 vdd2.n540 0.753
R4612 vdd2.n540 vdd2.n539 0.753
R4613 vdd2.n539 vdd2.n538 0.753
R4614 vdd2.n537 vdd2.n536 0.753
R4615 vdd2.n536 vdd2.n535 0.753
R4616 vdd2.n535 vdd2.n534 0.753
R4617 vdd2.n534 vdd2.n533 0.753
R4618 vdd2.n553 vdd2.n552 0.753
R4619 vdd2.n552 vdd2.n551 0.753
R4620 vdd2.n551 vdd2.n550 0.753
R4621 vdd2.n550 vdd2.n549 0.753
R4622 vdd2.n548 vdd2.n547 0.753
R4623 vdd2.n547 vdd2.n546 0.753
R4624 vdd2.n546 vdd2.n545 0.753
R4625 vdd2.n545 vdd2.n544 0.753
R4626 vdd2.n564 vdd2.n563 0.753
R4627 vdd2.n563 vdd2.n562 0.753
R4628 vdd2.n562 vdd2.n561 0.753
R4629 vdd2.n561 vdd2.n560 0.753
R4630 vdd2.n559 vdd2.n558 0.753
R4631 vdd2.n558 vdd2.n557 0.753
R4632 vdd2.n557 vdd2.n556 0.753
R4633 vdd2.n556 vdd2.n555 0.753
R4634 vdd2.n575 vdd2.n574 0.753
R4635 vdd2.n574 vdd2.n573 0.753
R4636 vdd2.n573 vdd2.n572 0.753
R4637 vdd2.n572 vdd2.n571 0.753
R4638 vdd2.n570 vdd2.n569 0.753
R4639 vdd2.n569 vdd2.n568 0.753
R4640 vdd2.n568 vdd2.n567 0.753
R4641 vdd2.n567 vdd2.n566 0.753
R4642 vdd2.n586 vdd2.n585 0.753
R4643 vdd2.n585 vdd2.n584 0.753
R4644 vdd2.n584 vdd2.n583 0.753
R4645 vdd2.n583 vdd2.n582 0.753
R4646 vdd2.n581 vdd2.n580 0.753
R4647 vdd2.n580 vdd2.n579 0.753
R4648 vdd2.n579 vdd2.n578 0.753
R4649 vdd2.n578 vdd2.n577 0.753
R4650 vdd2.n597 vdd2.n596 0.753
R4651 vdd2.n596 vdd2.n595 0.753
R4652 vdd2.n595 vdd2.n594 0.753
R4653 vdd2.n594 vdd2.n593 0.753
R4654 vdd2.n592 vdd2.n591 0.753
R4655 vdd2.n591 vdd2.n590 0.753
R4656 vdd2.n590 vdd2.n589 0.753
R4657 vdd2.n589 vdd2.n588 0.753
R4658 vdd2.n608 vdd2.n607 0.753
R4659 vdd2.n607 vdd2.n606 0.753
R4660 vdd2.n606 vdd2.n605 0.753
R4661 vdd2.n605 vdd2.n604 0.753
R4662 vdd2.n603 vdd2.n602 0.753
R4663 vdd2.n602 vdd2.n601 0.753
R4664 vdd2.n601 vdd2.n600 0.753
R4665 vdd2.n600 vdd2.n599 0.753
R4666 vdd2.n619 vdd2.n618 0.753
R4667 vdd2.n618 vdd2.n617 0.753
R4668 vdd2.n617 vdd2.n616 0.753
R4669 vdd2.n616 vdd2.n615 0.753
R4670 vdd2.n614 vdd2.n613 0.753
R4671 vdd2.n613 vdd2.n612 0.753
R4672 vdd2.n612 vdd2.n611 0.753
R4673 vdd2.n611 vdd2.n610 0.753
R4674 vdd2.n630 vdd2.n629 0.753
R4675 vdd2.n629 vdd2.n628 0.753
R4676 vdd2.n628 vdd2.n627 0.753
R4677 vdd2.n627 vdd2.n626 0.753
R4678 vdd2.n625 vdd2.n624 0.753
R4679 vdd2.n624 vdd2.n623 0.753
R4680 vdd2.n623 vdd2.n622 0.753
R4681 vdd2.n622 vdd2.n621 0.753
R4682 vdd2.n641 vdd2.n640 0.753
R4683 vdd2.n640 vdd2.n639 0.753
R4684 vdd2.n639 vdd2.n638 0.753
R4685 vdd2.n638 vdd2.n637 0.753
R4686 vdd2.n636 vdd2.n635 0.753
R4687 vdd2.n635 vdd2.n634 0.753
R4688 vdd2.n634 vdd2.n633 0.753
R4689 vdd2.n633 vdd2.n632 0.753
R4690 vdd2.n652 vdd2.n651 0.753
R4691 vdd2.n651 vdd2.n650 0.753
R4692 vdd2.n650 vdd2.n649 0.753
R4693 vdd2.n649 vdd2.n648 0.753
R4694 vdd2.n647 vdd2.n646 0.753
R4695 vdd2.n646 vdd2.n645 0.753
R4696 vdd2.n645 vdd2.n644 0.753
R4697 vdd2.n644 vdd2.n643 0.753
R4698 vdd2.n663 vdd2.n662 0.753
R4699 vdd2.n662 vdd2.n661 0.753
R4700 vdd2.n661 vdd2.n660 0.753
R4701 vdd2.n660 vdd2.n659 0.753
R4702 vdd2.n658 vdd2.n657 0.753
R4703 vdd2.n657 vdd2.n656 0.753
R4704 vdd2.n656 vdd2.n655 0.753
R4705 vdd2.n655 vdd2.n654 0.753
R4706 vdd2.n674 vdd2.n673 0.753
R4707 vdd2.n673 vdd2.n672 0.753
R4708 vdd2.n672 vdd2.n671 0.753
R4709 vdd2.n671 vdd2.n670 0.753
R4710 vdd2.n669 vdd2.n668 0.753
R4711 vdd2.n668 vdd2.n667 0.753
R4712 vdd2.n667 vdd2.n666 0.753
R4713 vdd2.n666 vdd2.n665 0.753
R4714 vdd2.n685 vdd2.n684 0.753
R4715 vdd2.n684 vdd2.n683 0.753
R4716 vdd2.n683 vdd2.n682 0.753
R4717 vdd2.n682 vdd2.n681 0.753
R4718 vdd2.n680 vdd2.n679 0.753
R4719 vdd2.n679 vdd2.n678 0.753
R4720 vdd2.n678 vdd2.n677 0.753
R4721 vdd2.n677 vdd2.n676 0.753
R4722 vdd2.n696 vdd2.n695 0.753
R4723 vdd2.n695 vdd2.n694 0.753
R4724 vdd2.n694 vdd2.n693 0.753
R4725 vdd2.n693 vdd2.n692 0.753
R4726 vdd2.n691 vdd2.n690 0.753
R4727 vdd2.n690 vdd2.n689 0.753
R4728 vdd2.n689 vdd2.n688 0.753
R4729 vdd2.n688 vdd2.n687 0.753
R4730 vdd2.n707 vdd2.n706 0.753
R4731 vdd2.n706 vdd2.n705 0.753
R4732 vdd2.n705 vdd2.n704 0.753
R4733 vdd2.n704 vdd2.n703 0.753
R4734 vdd2.n702 vdd2.n701 0.753
R4735 vdd2.n701 vdd2.n700 0.753
R4736 vdd2.n700 vdd2.n699 0.753
R4737 vdd2.n699 vdd2.n698 0.753
R4738 vdd2.n718 vdd2.n717 0.753
R4739 vdd2.n717 vdd2.n716 0.753
R4740 vdd2.n716 vdd2.n715 0.753
R4741 vdd2.n715 vdd2.n714 0.753
R4742 vdd2.n713 vdd2.n712 0.753
R4743 vdd2.n712 vdd2.n711 0.753
R4744 vdd2.n711 vdd2.n710 0.753
R4745 vdd2.n710 vdd2.n709 0.753
R4746 vdd2.n729 vdd2.n728 0.753
R4747 vdd2.n728 vdd2.n727 0.753
R4748 vdd2.n727 vdd2.n726 0.753
R4749 vdd2.n726 vdd2.n725 0.753
R4750 vdd2.n724 vdd2.n723 0.753
R4751 vdd2.n723 vdd2.n722 0.753
R4752 vdd2.n722 vdd2.n721 0.753
R4753 vdd2.n721 vdd2.n720 0.753
R4754 vdd2.n740 vdd2.n739 0.753
R4755 vdd2.n739 vdd2.n738 0.753
R4756 vdd2.n738 vdd2.n737 0.753
R4757 vdd2.n737 vdd2.n736 0.753
R4758 vdd2.n735 vdd2.n734 0.753
R4759 vdd2.n734 vdd2.n733 0.753
R4760 vdd2.n733 vdd2.n732 0.753
R4761 vdd2.n732 vdd2.n731 0.753
R4762 vdd2.n751 vdd2.n750 0.753
R4763 vdd2.n750 vdd2.n749 0.753
R4764 vdd2.n749 vdd2.n748 0.753
R4765 vdd2.n748 vdd2.n747 0.753
R4766 vdd2.n746 vdd2.n745 0.753
R4767 vdd2.n745 vdd2.n744 0.753
R4768 vdd2.n744 vdd2.n743 0.753
R4769 vdd2.n743 vdd2.n742 0.753
R4770 vdd2.n762 vdd2.n761 0.753
R4771 vdd2.n761 vdd2.n760 0.753
R4772 vdd2.n760 vdd2.n759 0.753
R4773 vdd2.n759 vdd2.n758 0.753
R4774 vdd2.n757 vdd2.n756 0.753
R4775 vdd2.n756 vdd2.n755 0.753
R4776 vdd2.n755 vdd2.n754 0.753
R4777 vdd2.n754 vdd2.n753 0.753
R4778 vdd2.n773 vdd2.n772 0.753
R4779 vdd2.n772 vdd2.n771 0.753
R4780 vdd2.n771 vdd2.n770 0.753
R4781 vdd2.n770 vdd2.n769 0.753
R4782 vdd2.n768 vdd2.n767 0.753
R4783 vdd2.n767 vdd2.n766 0.753
R4784 vdd2.n766 vdd2.n765 0.753
R4785 vdd2.n765 vdd2.n764 0.753
R4786 vdd2.n784 vdd2.n783 0.753
R4787 vdd2.n783 vdd2.n782 0.753
R4788 vdd2.n782 vdd2.n781 0.753
R4789 vdd2.n781 vdd2.n780 0.753
R4790 vdd2.n779 vdd2.n778 0.753
R4791 vdd2.n778 vdd2.n777 0.753
R4792 vdd2.n777 vdd2.n776 0.753
R4793 vdd2.n776 vdd2.n775 0.753
R4794 vdd2.n795 vdd2.n794 0.753
R4795 vdd2.n794 vdd2.n793 0.753
R4796 vdd2.n793 vdd2.n792 0.753
R4797 vdd2.n792 vdd2.n791 0.753
R4798 vdd2.n790 vdd2.n789 0.753
R4799 vdd2.n789 vdd2.n788 0.753
R4800 vdd2.n788 vdd2.n787 0.753
R4801 vdd2.n787 vdd2.n786 0.753
R4802 vdd2.n806 vdd2.n805 0.753
R4803 vdd2.n805 vdd2.n804 0.753
R4804 vdd2.n804 vdd2.n803 0.753
R4805 vdd2.n803 vdd2.n802 0.753
R4806 vdd2.n801 vdd2.n800 0.753
R4807 vdd2.n800 vdd2.n799 0.753
R4808 vdd2.n799 vdd2.n798 0.753
R4809 vdd2.n798 vdd2.n797 0.753
R4810 vdd2.n817 vdd2.n816 0.753
R4811 vdd2.n816 vdd2.n815 0.753
R4812 vdd2.n815 vdd2.n814 0.753
R4813 vdd2.n814 vdd2.n813 0.753
R4814 vdd2.n812 vdd2.n811 0.753
R4815 vdd2.n811 vdd2.n810 0.753
R4816 vdd2.n810 vdd2.n809 0.753
R4817 vdd2.n809 vdd2.n808 0.753
R4818 vdd2.n828 vdd2.n827 0.753
R4819 vdd2.n827 vdd2.n826 0.753
R4820 vdd2.n826 vdd2.n825 0.753
R4821 vdd2.n825 vdd2.n824 0.753
R4822 vdd2.n823 vdd2.n822 0.753
R4823 vdd2.n822 vdd2.n821 0.753
R4824 vdd2.n821 vdd2.n820 0.753
R4825 vdd2.n820 vdd2.n819 0.753
R4826 vdd2.n839 vdd2.n838 0.753
R4827 vdd2.n838 vdd2.n837 0.753
R4828 vdd2.n837 vdd2.n836 0.753
R4829 vdd2.n836 vdd2.n835 0.753
R4830 vdd2.n834 vdd2.n833 0.753
R4831 vdd2.n833 vdd2.n832 0.753
R4832 vdd2.n832 vdd2.n831 0.753
R4833 vdd2.n831 vdd2.n830 0.753
R4834 vdd2.n850 vdd2.n849 0.753
R4835 vdd2.n849 vdd2.n848 0.753
R4836 vdd2.n848 vdd2.n847 0.753
R4837 vdd2.n847 vdd2.n846 0.753
R4838 vdd2.n845 vdd2.n844 0.753
R4839 vdd2.n844 vdd2.n843 0.753
R4840 vdd2.n843 vdd2.n842 0.753
R4841 vdd2.n842 vdd2.n841 0.753
R4842 vdd2.n500 vdd2.n499 0.753
R4843 vdd2.n499 vdd2.n498 0.753
R4844 vdd2.n498 vdd2.n497 0.753
R4845 vdd2.n497 vdd2.n496 0.753
R4846 vdd2.n495 vdd2.n494 0.753
R4847 vdd2.n494 vdd2.n493 0.753
R4848 vdd2.n493 vdd2.n492 0.753
R4849 vdd2.n492 vdd2.n491 0.753
R4850 vdd2.n41 vdd2.n40 0.753
R4851 vdd2.n40 vdd2.n39 0.753
R4852 vdd2.n39 vdd2.n38 0.753
R4853 vdd2.n38 vdd2.n37 0.753
R4854 vdd2.n36 vdd2.n35 0.753
R4855 vdd2.n35 vdd2.n34 0.753
R4856 vdd2.n34 vdd2.n33 0.753
R4857 vdd2.n33 vdd2.n32 0.753
R4858 vdd2.n52 vdd2.n51 0.753
R4859 vdd2.n51 vdd2.n50 0.753
R4860 vdd2.n50 vdd2.n49 0.753
R4861 vdd2.n49 vdd2.n48 0.753
R4862 vdd2.n47 vdd2.n46 0.753
R4863 vdd2.n46 vdd2.n45 0.753
R4864 vdd2.n45 vdd2.n44 0.753
R4865 vdd2.n44 vdd2.n43 0.753
R4866 vdd2.n63 vdd2.n62 0.753
R4867 vdd2.n62 vdd2.n61 0.753
R4868 vdd2.n61 vdd2.n60 0.753
R4869 vdd2.n60 vdd2.n59 0.753
R4870 vdd2.n58 vdd2.n57 0.753
R4871 vdd2.n57 vdd2.n56 0.753
R4872 vdd2.n56 vdd2.n55 0.753
R4873 vdd2.n55 vdd2.n54 0.753
R4874 vdd2.n74 vdd2.n73 0.753
R4875 vdd2.n73 vdd2.n72 0.753
R4876 vdd2.n72 vdd2.n71 0.753
R4877 vdd2.n71 vdd2.n70 0.753
R4878 vdd2.n69 vdd2.n68 0.753
R4879 vdd2.n68 vdd2.n67 0.753
R4880 vdd2.n67 vdd2.n66 0.753
R4881 vdd2.n66 vdd2.n65 0.753
R4882 vdd2.n85 vdd2.n84 0.753
R4883 vdd2.n84 vdd2.n83 0.753
R4884 vdd2.n83 vdd2.n82 0.753
R4885 vdd2.n82 vdd2.n81 0.753
R4886 vdd2.n80 vdd2.n79 0.753
R4887 vdd2.n79 vdd2.n78 0.753
R4888 vdd2.n78 vdd2.n77 0.753
R4889 vdd2.n77 vdd2.n76 0.753
R4890 vdd2.n96 vdd2.n95 0.753
R4891 vdd2.n95 vdd2.n94 0.753
R4892 vdd2.n94 vdd2.n93 0.753
R4893 vdd2.n93 vdd2.n92 0.753
R4894 vdd2.n91 vdd2.n90 0.753
R4895 vdd2.n90 vdd2.n89 0.753
R4896 vdd2.n89 vdd2.n88 0.753
R4897 vdd2.n88 vdd2.n87 0.753
R4898 vdd2.n107 vdd2.n106 0.753
R4899 vdd2.n106 vdd2.n105 0.753
R4900 vdd2.n105 vdd2.n104 0.753
R4901 vdd2.n104 vdd2.n103 0.753
R4902 vdd2.n102 vdd2.n101 0.753
R4903 vdd2.n101 vdd2.n100 0.753
R4904 vdd2.n100 vdd2.n99 0.753
R4905 vdd2.n99 vdd2.n98 0.753
R4906 vdd2.n118 vdd2.n117 0.753
R4907 vdd2.n117 vdd2.n116 0.753
R4908 vdd2.n116 vdd2.n115 0.753
R4909 vdd2.n115 vdd2.n114 0.753
R4910 vdd2.n113 vdd2.n112 0.753
R4911 vdd2.n112 vdd2.n111 0.753
R4912 vdd2.n111 vdd2.n110 0.753
R4913 vdd2.n110 vdd2.n109 0.753
R4914 vdd2.n129 vdd2.n128 0.753
R4915 vdd2.n128 vdd2.n127 0.753
R4916 vdd2.n127 vdd2.n126 0.753
R4917 vdd2.n126 vdd2.n125 0.753
R4918 vdd2.n124 vdd2.n123 0.753
R4919 vdd2.n123 vdd2.n122 0.753
R4920 vdd2.n122 vdd2.n121 0.753
R4921 vdd2.n121 vdd2.n120 0.753
R4922 vdd2.n140 vdd2.n139 0.753
R4923 vdd2.n139 vdd2.n138 0.753
R4924 vdd2.n138 vdd2.n137 0.753
R4925 vdd2.n137 vdd2.n136 0.753
R4926 vdd2.n135 vdd2.n134 0.753
R4927 vdd2.n134 vdd2.n133 0.753
R4928 vdd2.n133 vdd2.n132 0.753
R4929 vdd2.n132 vdd2.n131 0.753
R4930 vdd2.n151 vdd2.n150 0.753
R4931 vdd2.n150 vdd2.n149 0.753
R4932 vdd2.n149 vdd2.n148 0.753
R4933 vdd2.n148 vdd2.n147 0.753
R4934 vdd2.n146 vdd2.n145 0.753
R4935 vdd2.n145 vdd2.n144 0.753
R4936 vdd2.n144 vdd2.n143 0.753
R4937 vdd2.n143 vdd2.n142 0.753
R4938 vdd2.n162 vdd2.n161 0.753
R4939 vdd2.n161 vdd2.n160 0.753
R4940 vdd2.n160 vdd2.n159 0.753
R4941 vdd2.n159 vdd2.n158 0.753
R4942 vdd2.n157 vdd2.n156 0.753
R4943 vdd2.n156 vdd2.n155 0.753
R4944 vdd2.n155 vdd2.n154 0.753
R4945 vdd2.n154 vdd2.n153 0.753
R4946 vdd2.n173 vdd2.n172 0.753
R4947 vdd2.n172 vdd2.n171 0.753
R4948 vdd2.n171 vdd2.n170 0.753
R4949 vdd2.n170 vdd2.n169 0.753
R4950 vdd2.n168 vdd2.n167 0.753
R4951 vdd2.n167 vdd2.n166 0.753
R4952 vdd2.n166 vdd2.n165 0.753
R4953 vdd2.n165 vdd2.n164 0.753
R4954 vdd2.n184 vdd2.n183 0.753
R4955 vdd2.n183 vdd2.n182 0.753
R4956 vdd2.n182 vdd2.n181 0.753
R4957 vdd2.n181 vdd2.n180 0.753
R4958 vdd2.n179 vdd2.n178 0.753
R4959 vdd2.n178 vdd2.n177 0.753
R4960 vdd2.n177 vdd2.n176 0.753
R4961 vdd2.n176 vdd2.n175 0.753
R4962 vdd2.n195 vdd2.n194 0.753
R4963 vdd2.n194 vdd2.n193 0.753
R4964 vdd2.n193 vdd2.n192 0.753
R4965 vdd2.n192 vdd2.n191 0.753
R4966 vdd2.n190 vdd2.n189 0.753
R4967 vdd2.n189 vdd2.n188 0.753
R4968 vdd2.n188 vdd2.n187 0.753
R4969 vdd2.n187 vdd2.n186 0.753
R4970 vdd2.n206 vdd2.n205 0.753
R4971 vdd2.n205 vdd2.n204 0.753
R4972 vdd2.n204 vdd2.n203 0.753
R4973 vdd2.n203 vdd2.n202 0.753
R4974 vdd2.n201 vdd2.n200 0.753
R4975 vdd2.n200 vdd2.n199 0.753
R4976 vdd2.n199 vdd2.n198 0.753
R4977 vdd2.n198 vdd2.n197 0.753
R4978 vdd2.n217 vdd2.n216 0.753
R4979 vdd2.n216 vdd2.n215 0.753
R4980 vdd2.n215 vdd2.n214 0.753
R4981 vdd2.n214 vdd2.n213 0.753
R4982 vdd2.n212 vdd2.n211 0.753
R4983 vdd2.n211 vdd2.n210 0.753
R4984 vdd2.n210 vdd2.n209 0.753
R4985 vdd2.n209 vdd2.n208 0.753
R4986 vdd2.n228 vdd2.n227 0.753
R4987 vdd2.n227 vdd2.n226 0.753
R4988 vdd2.n226 vdd2.n225 0.753
R4989 vdd2.n225 vdd2.n224 0.753
R4990 vdd2.n223 vdd2.n222 0.753
R4991 vdd2.n222 vdd2.n221 0.753
R4992 vdd2.n221 vdd2.n220 0.753
R4993 vdd2.n220 vdd2.n219 0.753
R4994 vdd2.n239 vdd2.n238 0.753
R4995 vdd2.n238 vdd2.n237 0.753
R4996 vdd2.n237 vdd2.n236 0.753
R4997 vdd2.n236 vdd2.n235 0.753
R4998 vdd2.n234 vdd2.n233 0.753
R4999 vdd2.n233 vdd2.n232 0.753
R5000 vdd2.n232 vdd2.n231 0.753
R5001 vdd2.n231 vdd2.n230 0.753
R5002 vdd2.n250 vdd2.n249 0.753
R5003 vdd2.n249 vdd2.n248 0.753
R5004 vdd2.n248 vdd2.n247 0.753
R5005 vdd2.n247 vdd2.n246 0.753
R5006 vdd2.n245 vdd2.n244 0.753
R5007 vdd2.n244 vdd2.n243 0.753
R5008 vdd2.n243 vdd2.n242 0.753
R5009 vdd2.n242 vdd2.n241 0.753
R5010 vdd2.n261 vdd2.n260 0.753
R5011 vdd2.n260 vdd2.n259 0.753
R5012 vdd2.n259 vdd2.n258 0.753
R5013 vdd2.n258 vdd2.n257 0.753
R5014 vdd2.n256 vdd2.n255 0.753
R5015 vdd2.n255 vdd2.n254 0.753
R5016 vdd2.n254 vdd2.n253 0.753
R5017 vdd2.n253 vdd2.n252 0.753
R5018 vdd2.n272 vdd2.n271 0.753
R5019 vdd2.n271 vdd2.n270 0.753
R5020 vdd2.n270 vdd2.n269 0.753
R5021 vdd2.n269 vdd2.n268 0.753
R5022 vdd2.n267 vdd2.n266 0.753
R5023 vdd2.n266 vdd2.n265 0.753
R5024 vdd2.n265 vdd2.n264 0.753
R5025 vdd2.n264 vdd2.n263 0.753
R5026 vdd2.n283 vdd2.n282 0.753
R5027 vdd2.n282 vdd2.n281 0.753
R5028 vdd2.n281 vdd2.n280 0.753
R5029 vdd2.n280 vdd2.n279 0.753
R5030 vdd2.n278 vdd2.n277 0.753
R5031 vdd2.n277 vdd2.n276 0.753
R5032 vdd2.n276 vdd2.n275 0.753
R5033 vdd2.n275 vdd2.n274 0.753
R5034 vdd2.n294 vdd2.n293 0.753
R5035 vdd2.n293 vdd2.n292 0.753
R5036 vdd2.n292 vdd2.n291 0.753
R5037 vdd2.n291 vdd2.n290 0.753
R5038 vdd2.n289 vdd2.n288 0.753
R5039 vdd2.n288 vdd2.n287 0.753
R5040 vdd2.n287 vdd2.n286 0.753
R5041 vdd2.n286 vdd2.n285 0.753
R5042 vdd2.n305 vdd2.n304 0.753
R5043 vdd2.n304 vdd2.n303 0.753
R5044 vdd2.n303 vdd2.n302 0.753
R5045 vdd2.n302 vdd2.n301 0.753
R5046 vdd2.n300 vdd2.n299 0.753
R5047 vdd2.n299 vdd2.n298 0.753
R5048 vdd2.n298 vdd2.n297 0.753
R5049 vdd2.n297 vdd2.n296 0.753
R5050 vdd2.n316 vdd2.n315 0.753
R5051 vdd2.n315 vdd2.n314 0.753
R5052 vdd2.n314 vdd2.n313 0.753
R5053 vdd2.n313 vdd2.n312 0.753
R5054 vdd2.n311 vdd2.n310 0.753
R5055 vdd2.n310 vdd2.n309 0.753
R5056 vdd2.n309 vdd2.n308 0.753
R5057 vdd2.n308 vdd2.n307 0.753
R5058 vdd2.n327 vdd2.n326 0.753
R5059 vdd2.n326 vdd2.n325 0.753
R5060 vdd2.n325 vdd2.n324 0.753
R5061 vdd2.n324 vdd2.n323 0.753
R5062 vdd2.n322 vdd2.n321 0.753
R5063 vdd2.n321 vdd2.n320 0.753
R5064 vdd2.n320 vdd2.n319 0.753
R5065 vdd2.n319 vdd2.n318 0.753
R5066 vdd2.n338 vdd2.n337 0.753
R5067 vdd2.n337 vdd2.n336 0.753
R5068 vdd2.n336 vdd2.n335 0.753
R5069 vdd2.n335 vdd2.n334 0.753
R5070 vdd2.n333 vdd2.n332 0.753
R5071 vdd2.n332 vdd2.n331 0.753
R5072 vdd2.n331 vdd2.n330 0.753
R5073 vdd2.n330 vdd2.n329 0.753
R5074 vdd2.n349 vdd2.n348 0.753
R5075 vdd2.n348 vdd2.n347 0.753
R5076 vdd2.n347 vdd2.n346 0.753
R5077 vdd2.n346 vdd2.n345 0.753
R5078 vdd2.n344 vdd2.n343 0.753
R5079 vdd2.n343 vdd2.n342 0.753
R5080 vdd2.n342 vdd2.n341 0.753
R5081 vdd2.n341 vdd2.n340 0.753
R5082 vdd2.n360 vdd2.n359 0.753
R5083 vdd2.n359 vdd2.n358 0.753
R5084 vdd2.n358 vdd2.n357 0.753
R5085 vdd2.n357 vdd2.n356 0.753
R5086 vdd2.n355 vdd2.n354 0.753
R5087 vdd2.n354 vdd2.n353 0.753
R5088 vdd2.n353 vdd2.n352 0.753
R5089 vdd2.n352 vdd2.n351 0.753
R5090 vdd2.n371 vdd2.n370 0.753
R5091 vdd2.n370 vdd2.n369 0.753
R5092 vdd2.n369 vdd2.n368 0.753
R5093 vdd2.n368 vdd2.n367 0.753
R5094 vdd2.n366 vdd2.n365 0.753
R5095 vdd2.n365 vdd2.n364 0.753
R5096 vdd2.n364 vdd2.n363 0.753
R5097 vdd2.n363 vdd2.n362 0.753
R5098 vdd2.n382 vdd2.n381 0.753
R5099 vdd2.n381 vdd2.n380 0.753
R5100 vdd2.n380 vdd2.n379 0.753
R5101 vdd2.n379 vdd2.n378 0.753
R5102 vdd2.n377 vdd2.n376 0.753
R5103 vdd2.n376 vdd2.n375 0.753
R5104 vdd2.n375 vdd2.n374 0.753
R5105 vdd2.n374 vdd2.n373 0.753
R5106 vdd2.n393 vdd2.n392 0.753
R5107 vdd2.n392 vdd2.n391 0.753
R5108 vdd2.n391 vdd2.n390 0.753
R5109 vdd2.n390 vdd2.n389 0.753
R5110 vdd2.n388 vdd2.n387 0.753
R5111 vdd2.n387 vdd2.n386 0.753
R5112 vdd2.n386 vdd2.n385 0.753
R5113 vdd2.n385 vdd2.n384 0.753
R5114 vdd2.n21 vdd2.n20 0.753
R5115 vdd2.n20 vdd2.n19 0.753
R5116 vdd2.n19 vdd2.n18 0.753
R5117 vdd2.n18 vdd2.n17 0.753
R5118 vdd2.n16 vdd2.n15 0.753
R5119 vdd2.n15 vdd2.n14 0.753
R5120 vdd2.n14 vdd2.n13 0.753
R5121 vdd2.n13 vdd2.n12 0.753
R5122 vdd2.n405 vdd2.n404 0.753
R5123 vdd2.n404 vdd2.n403 0.753
R5124 vdd2.n403 vdd2.n402 0.753
R5125 vdd2.n402 vdd2.n401 0.753
R5126 vdd2.n400 vdd2.n399 0.753
R5127 vdd2.n399 vdd2.n398 0.753
R5128 vdd2.n398 vdd2.n397 0.753
R5129 vdd2.n397 vdd2.n396 0.753
R5130 vdd2.n416 vdd2.n415 0.753
R5131 vdd2.n415 vdd2.n414 0.753
R5132 vdd2.n414 vdd2.n413 0.753
R5133 vdd2.n413 vdd2.n412 0.753
R5134 vdd2.n411 vdd2.n410 0.753
R5135 vdd2.n410 vdd2.n409 0.753
R5136 vdd2.n409 vdd2.n408 0.753
R5137 vdd2.n408 vdd2.n407 0.753
R5138 vdd2.n427 vdd2.n426 0.753
R5139 vdd2.n426 vdd2.n425 0.753
R5140 vdd2.n425 vdd2.n424 0.753
R5141 vdd2.n424 vdd2.n423 0.753
R5142 vdd2.n422 vdd2.n421 0.753
R5143 vdd2.n421 vdd2.n420 0.753
R5144 vdd2.n420 vdd2.n419 0.753
R5145 vdd2.n419 vdd2.n418 0.753
R5146 vdd2.n453 vdd2.n452 0.753
R5147 vdd2.n452 vdd2.n451 0.753
R5148 vdd2.n451 vdd2.n450 0.753
R5149 vdd2.n450 vdd2.n449 0.753
R5150 vdd2.n448 vdd2.n447 0.753
R5151 vdd2.n447 vdd2.n446 0.753
R5152 vdd2.n446 vdd2.n445 0.753
R5153 vdd2.n445 vdd2.n444 0.753
R5154 vdd2.n465 vdd2.n464 0.753
R5155 vdd2.n464 vdd2.n463 0.753
R5156 vdd2.n463 vdd2.n462 0.753
R5157 vdd2.n462 vdd2.n461 0.753
R5158 vdd2.n460 vdd2.n459 0.753
R5159 vdd2.n459 vdd2.n458 0.753
R5160 vdd2.n458 vdd2.n457 0.753
R5161 vdd2.n457 vdd2.n456 0.753
R5162 vdd2.n476 vdd2.n475 0.753
R5163 vdd2.n475 vdd2.n474 0.753
R5164 vdd2.n474 vdd2.n473 0.753
R5165 vdd2.n473 vdd2.n472 0.753
R5166 vdd2.n471 vdd2.n470 0.753
R5167 vdd2.n470 vdd2.n469 0.753
R5168 vdd2.n469 vdd2.n468 0.753
R5169 vdd2.n468 vdd2.n467 0.753
R5170 vdd2.n487 vdd2.n486 0.753
R5171 vdd2.n486 vdd2.n485 0.753
R5172 vdd2.n485 vdd2.n484 0.753
R5173 vdd2.n484 vdd2.n483 0.753
R5174 vdd2.n482 vdd2.n481 0.753
R5175 vdd2.n481 vdd2.n480 0.753
R5176 vdd2.n480 vdd2.n479 0.753
R5177 vdd2.n479 vdd2.n478 0.753
R5178 vdd2.n9 vdd2.n8 0.753
R5179 vdd2.n8 vdd2.n7 0.753
R5180 vdd2.n7 vdd2.n6 0.753
R5181 vdd2.n6 vdd2.n5 0.753
R5182 vdd2.n4 vdd2.n3 0.753
R5183 vdd2.n3 vdd2.n2 0.753
R5184 vdd2.n2 vdd2.n1 0.753
R5185 vdd2.n1 vdd2.n0 0.753
R5186 vdd2.n27 vdd2.n26 0.726
R5187 vdd2.n24 vdd2.n23 0.58
R5188 vdd2.n25 vdd2.n24 0.58
R5189 vdd2.n26 vdd2.n25 0.58
R5190 vdd2.n28 vdd2.n27 0.58
R5191 vdd2.n29 vdd2.n28 0.58
R5192 vdd2.n30 vdd2.n29 0.58
R5193 vdd2.n31 vdd2.n30 0.58
R5194 vdd2.n42 vdd2.n31 0.515
R5195 vdd2.n521 vdd2.n520 0.427
R5196 vdd2.n532 vdd2.n531 0.427
R5197 vdd2.n543 vdd2.n542 0.427
R5198 vdd2.n554 vdd2.n553 0.427
R5199 vdd2.n565 vdd2.n564 0.427
R5200 vdd2.n576 vdd2.n575 0.427
R5201 vdd2.n587 vdd2.n586 0.427
R5202 vdd2.n598 vdd2.n597 0.427
R5203 vdd2.n609 vdd2.n608 0.427
R5204 vdd2.n620 vdd2.n619 0.427
R5205 vdd2.n631 vdd2.n630 0.427
R5206 vdd2.n642 vdd2.n641 0.427
R5207 vdd2.n653 vdd2.n652 0.427
R5208 vdd2.n664 vdd2.n663 0.427
R5209 vdd2.n675 vdd2.n674 0.427
R5210 vdd2.n686 vdd2.n685 0.427
R5211 vdd2.n697 vdd2.n696 0.427
R5212 vdd2.n708 vdd2.n707 0.427
R5213 vdd2.n719 vdd2.n718 0.427
R5214 vdd2.n730 vdd2.n729 0.427
R5215 vdd2.n741 vdd2.n740 0.427
R5216 vdd2.n752 vdd2.n751 0.427
R5217 vdd2.n763 vdd2.n762 0.427
R5218 vdd2.n774 vdd2.n773 0.427
R5219 vdd2.n785 vdd2.n784 0.427
R5220 vdd2.n796 vdd2.n795 0.427
R5221 vdd2.n807 vdd2.n806 0.427
R5222 vdd2.n818 vdd2.n817 0.427
R5223 vdd2.n829 vdd2.n828 0.427
R5224 vdd2.n840 vdd2.n839 0.427
R5225 vdd2.n851 vdd2.n850 0.427
R5226 vdd2.n53 vdd2.n52 0.427
R5227 vdd2.n64 vdd2.n63 0.427
R5228 vdd2.n75 vdd2.n74 0.427
R5229 vdd2.n86 vdd2.n85 0.427
R5230 vdd2.n97 vdd2.n96 0.427
R5231 vdd2.n108 vdd2.n107 0.427
R5232 vdd2.n119 vdd2.n118 0.427
R5233 vdd2.n130 vdd2.n129 0.427
R5234 vdd2.n141 vdd2.n140 0.427
R5235 vdd2.n152 vdd2.n151 0.427
R5236 vdd2.n163 vdd2.n162 0.427
R5237 vdd2.n174 vdd2.n173 0.427
R5238 vdd2.n185 vdd2.n184 0.427
R5239 vdd2.n196 vdd2.n195 0.427
R5240 vdd2.n207 vdd2.n206 0.427
R5241 vdd2.n218 vdd2.n217 0.427
R5242 vdd2.n229 vdd2.n228 0.427
R5243 vdd2.n240 vdd2.n239 0.427
R5244 vdd2.n251 vdd2.n250 0.427
R5245 vdd2.n262 vdd2.n261 0.427
R5246 vdd2.n273 vdd2.n272 0.427
R5247 vdd2.n284 vdd2.n283 0.427
R5248 vdd2.n295 vdd2.n294 0.427
R5249 vdd2.n306 vdd2.n305 0.427
R5250 vdd2.n317 vdd2.n316 0.427
R5251 vdd2.n328 vdd2.n327 0.427
R5252 vdd2.n339 vdd2.n338 0.427
R5253 vdd2.n350 vdd2.n349 0.427
R5254 vdd2.n361 vdd2.n360 0.427
R5255 vdd2.n372 vdd2.n371 0.427
R5256 vdd2.n383 vdd2.n382 0.427
R5257 vdd2.n394 vdd2.n393 0.427
R5258 vdd2.n406 vdd2.n405 0.427
R5259 vdd2.n417 vdd2.n416 0.427
R5260 vdd2.n428 vdd2.n427 0.427
R5261 vdd2.n466 vdd2.n465 0.427
R5262 vdd2.n477 vdd2.n476 0.427
R5263 vdd2.n488 vdd2.n487 0.427
R5264 vdd2.n42 vdd2.n41 0.427
R5265 vdd2.n501 vdd2.n500 0.427
R5266 vdd2.n454 vdd2.n453 0.427
R5267 vdd2.n22 vdd2.n21 0.426
R5268 vdd2.n10 vdd2.n9 0.426
R5269 vdd2 vdd2.n11 0.224
R5270 vdd2.n22 vdd2.n11 0.16
R5271 vdd2.n395 vdd2.n11 0.094
R5272 vdd2.n490 vdd2.n489 0.094
R5273 vdd2.n443 vdd2.n442 0.093
R5274 vdd2.n53 vdd2.n42 0.004
R5275 vdd2.n532 vdd2.n521 0.004
R5276 vdd2.n543 vdd2.n532 0.004
R5277 vdd2.n554 vdd2.n543 0.004
R5278 vdd2.n565 vdd2.n554 0.004
R5279 vdd2.n576 vdd2.n565 0.004
R5280 vdd2.n587 vdd2.n576 0.004
R5281 vdd2.n598 vdd2.n587 0.004
R5282 vdd2.n609 vdd2.n598 0.004
R5283 vdd2.n620 vdd2.n609 0.004
R5284 vdd2.n631 vdd2.n620 0.004
R5285 vdd2.n642 vdd2.n631 0.004
R5286 vdd2.n653 vdd2.n642 0.004
R5287 vdd2.n664 vdd2.n653 0.004
R5288 vdd2.n675 vdd2.n664 0.004
R5289 vdd2.n686 vdd2.n675 0.004
R5290 vdd2.n697 vdd2.n686 0.004
R5291 vdd2.n708 vdd2.n697 0.004
R5292 vdd2.n719 vdd2.n708 0.004
R5293 vdd2.n730 vdd2.n719 0.004
R5294 vdd2.n741 vdd2.n730 0.004
R5295 vdd2.n752 vdd2.n741 0.004
R5296 vdd2.n763 vdd2.n752 0.004
R5297 vdd2.n774 vdd2.n763 0.004
R5298 vdd2.n785 vdd2.n774 0.004
R5299 vdd2.n796 vdd2.n785 0.004
R5300 vdd2.n807 vdd2.n796 0.004
R5301 vdd2.n818 vdd2.n807 0.004
R5302 vdd2.n829 vdd2.n818 0.004
R5303 vdd2.n840 vdd2.n829 0.004
R5304 vdd2.n851 vdd2.n840 0.004
R5305 vdd2.n64 vdd2.n53 0.004
R5306 vdd2.n75 vdd2.n64 0.004
R5307 vdd2.n86 vdd2.n75 0.004
R5308 vdd2.n97 vdd2.n86 0.004
R5309 vdd2.n108 vdd2.n97 0.004
R5310 vdd2.n119 vdd2.n108 0.004
R5311 vdd2.n130 vdd2.n119 0.004
R5312 vdd2.n141 vdd2.n130 0.004
R5313 vdd2.n152 vdd2.n141 0.004
R5314 vdd2.n163 vdd2.n152 0.004
R5315 vdd2.n174 vdd2.n163 0.004
R5316 vdd2.n185 vdd2.n174 0.004
R5317 vdd2.n196 vdd2.n185 0.004
R5318 vdd2.n207 vdd2.n196 0.004
R5319 vdd2.n218 vdd2.n207 0.004
R5320 vdd2.n229 vdd2.n218 0.004
R5321 vdd2.n240 vdd2.n229 0.004
R5322 vdd2.n251 vdd2.n240 0.004
R5323 vdd2.n262 vdd2.n251 0.004
R5324 vdd2.n273 vdd2.n262 0.004
R5325 vdd2.n284 vdd2.n273 0.004
R5326 vdd2.n295 vdd2.n284 0.004
R5327 vdd2.n306 vdd2.n295 0.004
R5328 vdd2.n317 vdd2.n306 0.004
R5329 vdd2.n328 vdd2.n317 0.004
R5330 vdd2.n339 vdd2.n328 0.004
R5331 vdd2.n350 vdd2.n339 0.004
R5332 vdd2.n361 vdd2.n350 0.004
R5333 vdd2.n372 vdd2.n361 0.004
R5334 vdd2.n383 vdd2.n372 0.004
R5335 vdd2.n394 vdd2.n383 0.004
R5336 vdd2.n417 vdd2.n406 0.004
R5337 vdd2.n428 vdd2.n417 0.004
R5338 vdd2.n477 vdd2.n466 0.004
R5339 vdd2.n488 vdd2.n477 0.004
R5340 vdd2.n406 vdd2 0.003
R5341 vdd2.n466 vdd2.n455 0.003
R5342 vdd2.n852 vdd2.n851 0.003
R5343 vdd2 vdd2.n395 0.002
R5344 vdd2.n455 vdd2.n443 0.002
R5345 vdd2.n853 vdd2.n490 0.002
R5346 vdd2.n853 vdd2.n852 0.002
R5347 vdd2.n852 vdd2.n501 0.001
R5348 vdd2.n455 vdd2.n454 0.001
R5349 vdd2 vdd2.n22 0.001
R5350 vdd2.n853 vdd2.n10 0.001
R5351 vdd2.n442 vdd2.n441 0.001
R5352 vdd2.n395 vdd2.n394 0.001
R5353 vdd2.n443 vdd2.n428 0.001
R5354 vdd2.n490 vdd2.n488 0.001
R5355 vdd2.n854 vdd2.n853 0.001
R5356 out_n.n619 out_n.t1014 8.126
R5357 out_n.n619 out_n.t439 8.126
R5358 out_n.n618 out_n.t1291 8.126
R5359 out_n.n618 out_n.t718 8.126
R5360 out_n.n617 out_n.t1425 8.126
R5361 out_n.n617 out_n.t845 8.126
R5362 out_n.n616 out_n.t492 8.126
R5363 out_n.n616 out_n.t1417 8.126
R5364 out_n.n615 out_n.t1049 8.126
R5365 out_n.n615 out_n.t474 8.126
R5366 out_n.n614 out_n.t764 8.126
R5367 out_n.n614 out_n.t1687 8.126
R5368 out_n.n613 out_n.t535 8.126
R5369 out_n.n613 out_n.t1459 8.126
R5370 out_n.n612 out_n.t1099 8.126
R5371 out_n.n612 out_n.t526 8.126
R5372 out_n.n611 out_n.t1662 8.126
R5373 out_n.n611 out_n.t1090 8.126
R5374 out_n.n610 out_n.t1431 8.126
R5375 out_n.n610 out_n.t852 8.126
R5376 out_n.n600 out_n.t278 8.126
R5377 out_n.n600 out_n.t308 8.126
R5378 out_n.n601 out_n.t519 8.126
R5379 out_n.n601 out_n.t550 8.126
R5380 out_n.n602 out_n.t1448 8.126
R5381 out_n.n602 out_n.t1478 8.126
R5382 out_n.n603 out_n.t876 8.126
R5383 out_n.n603 out_n.t904 8.126
R5384 out_n.n604 out_n.t1117 8.126
R5385 out_n.n604 out_n.t1145 8.126
R5386 out_n.n605 out_n.t1400 8.126
R5387 out_n.n605 out_n.t1432 8.126
R5388 out_n.n606 out_n.t838 8.126
R5389 out_n.n606 out_n.t866 8.126
R5390 out_n.n607 out_n.t270 8.126
R5391 out_n.n607 out_n.t302 8.126
R5392 out_n.n608 out_n.t1638 8.126
R5393 out_n.n608 out_n.t1671 8.126
R5394 out_n.n609 out_n.t1366 8.126
R5395 out_n.n609 out_n.t1396 8.126
R5396 out_n.n590 out_n.t1232 8.126
R5397 out_n.n590 out_n.t654 8.126
R5398 out_n.n591 out_n.t1474 8.126
R5399 out_n.n591 out_n.t889 8.126
R5400 out_n.n592 out_n.t893 8.126
R5401 out_n.n592 out_n.t322 8.126
R5402 out_n.n593 out_n.t330 8.126
R5403 out_n.n593 out_n.t1256 8.126
R5404 out_n.n594 out_n.t574 8.126
R5405 out_n.n594 out_n.t1494 8.126
R5406 out_n.n595 out_n.t853 8.126
R5407 out_n.n595 out_n.t279 8.126
R5408 out_n.n596 out_n.t296 8.126
R5409 out_n.n596 out_n.t1216 8.126
R5410 out_n.n597 out_n.t1224 8.126
R5411 out_n.n597 out_n.t647 8.126
R5412 out_n.n598 out_n.t1100 8.126
R5413 out_n.n598 out_n.t527 8.126
R5414 out_n.n599 out_n.t815 8.126
R5415 out_n.n599 out_n.t1738 8.126
R5416 out_n.n580 out_n.t1568 8.126
R5417 out_n.n580 out_n.t348 8.126
R5418 out_n.n581 out_n.t319 8.126
R5419 out_n.n581 out_n.t596 8.126
R5420 out_n.n582 out_n.t1249 8.126
R5421 out_n.n582 out_n.t1519 8.126
R5422 out_n.n583 out_n.t681 8.126
R5423 out_n.n583 out_n.t951 8.126
R5424 out_n.n584 out_n.t910 8.126
R5425 out_n.n584 out_n.t1193 8.126
R5426 out_n.n585 out_n.t1197 8.126
R5427 out_n.n585 out_n.t1484 8.126
R5428 out_n.n586 out_n.t638 8.126
R5429 out_n.n586 out_n.t914 8.126
R5430 out_n.n587 out_n.t1560 8.126
R5431 out_n.n587 out_n.t345 8.126
R5432 out_n.n588 out_n.t1449 8.126
R5433 out_n.n588 out_n.t1724 8.126
R5434 out_n.n589 out_n.t1160 8.126
R5435 out_n.n589 out_n.t1447 8.126
R5436 out_n.n570 out_n.t378 8.126
R5437 out_n.n570 out_n.t1299 8.126
R5438 out_n.n571 out_n.t624 8.126
R5439 out_n.n571 out_n.t1542 8.126
R5440 out_n.n572 out_n.t1550 8.126
R5441 out_n.n572 out_n.t971 8.126
R5442 out_n.n573 out_n.t983 8.126
R5443 out_n.n573 out_n.t403 8.126
R5444 out_n.n574 out_n.t1228 8.126
R5445 out_n.n574 out_n.t651 8.126
R5446 out_n.n575 out_n.t1510 8.126
R5447 out_n.n575 out_n.t925 8.126
R5448 out_n.n576 out_n.t941 8.126
R5449 out_n.n576 out_n.t363 8.126
R5450 out_n.n577 out_n.t370 8.126
R5451 out_n.n577 out_n.t1292 8.126
R5452 out_n.n578 out_n.t1761 8.126
R5453 out_n.n578 out_n.t1178 8.126
R5454 out_n.n579 out_n.t1479 8.126
R5455 out_n.n579 out_n.t892 8.126
R5456 out_n.n560 out_n.t728 8.126
R5457 out_n.n560 out_n.t1648 8.126
R5458 out_n.n561 out_n.t964 8.126
R5459 out_n.n561 out_n.t384 8.126
R5460 out_n.n562 out_n.t393 8.126
R5461 out_n.n562 out_n.t1317 8.126
R5462 out_n.n563 out_n.t1328 8.126
R5463 out_n.n563 out_n.t751 8.126
R5464 out_n.n564 out_n.t1564 8.126
R5465 out_n.n564 out_n.t991 8.126
R5466 out_n.n565 out_n.t349 8.126
R5467 out_n.n565 out_n.t1272 8.126
R5468 out_n.n566 out_n.t1287 8.126
R5469 out_n.n566 out_n.t715 8.126
R5470 out_n.n567 out_n.t721 8.126
R5471 out_n.n567 out_n.t1642 8.126
R5472 out_n.n568 out_n.t603 8.126
R5473 out_n.n568 out_n.t1520 8.126
R5474 out_n.n569 out_n.t323 8.126
R5475 out_n.n569 out_n.t1248 8.126
R5476 out_n.n550 out_n.t1074 8.126
R5477 out_n.n550 out_n.t1111 8.126
R5478 out_n.n551 out_n.t1307 8.126
R5479 out_n.n551 out_n.t1343 8.126
R5480 out_n.n552 out_n.t740 8.126
R5481 out_n.n552 out_n.t772 8.126
R5482 out_n.n553 out_n.t1676 8.126
R5483 out_n.n553 out_n.t1706 8.126
R5484 out_n.n554 out_n.t413 8.126
R5485 out_n.n554 out_n.t447 8.126
R5486 out_n.n555 out_n.t703 8.126
R5487 out_n.n555 out_n.t729 8.126
R5488 out_n.n556 out_n.t1634 8.126
R5489 out_n.n556 out_n.t1664 8.126
R5490 out_n.n557 out_n.t1067 8.126
R5491 out_n.n557 out_n.t1104 8.126
R5492 out_n.n558 out_n.t944 8.126
R5493 out_n.n558 out_n.t973 8.126
R5494 out_n.n559 out_n.t673 8.126
R5495 out_n.n559 out_n.t699 8.126
R5496 out_n.n540 out_n.t536 8.126
R5497 out_n.n540 out_n.t1460 8.126
R5498 out_n.n541 out_n.t767 8.126
R5499 out_n.n541 out_n.t1689 8.126
R5500 out_n.n542 out_n.t1696 8.126
R5501 out_n.n542 out_n.t1125 8.126
R5502 out_n.n543 out_n.t1133 8.126
R5503 out_n.n543 out_n.t564 8.126
R5504 out_n.n544 out_n.t1374 8.126
R5505 out_n.n544 out_n.t791 8.126
R5506 out_n.n545 out_n.t1649 8.126
R5507 out_n.n545 out_n.t1075 8.126
R5508 out_n.n546 out_n.t1093 8.126
R5509 out_n.n546 out_n.t520 8.126
R5510 out_n.n547 out_n.t529 8.126
R5511 out_n.n547 out_n.t1454 8.126
R5512 out_n.n548 out_n.t394 8.126
R5513 out_n.n548 out_n.t1318 8.126
R5514 out_n.n549 out_n.t1614 8.126
R5515 out_n.n549 out_n.t1039 8.126
R5516 out_n.n530 out_n.t877 8.126
R5517 out_n.n530 out_n.t268 8.126
R5518 out_n.n531 out_n.t1119 8.126
R5519 out_n.n531 out_n.t505 8.126
R5520 out_n.n532 out_n.t553 8.126
R5521 out_n.n532 out_n.t1439 8.126
R5522 out_n.n533 out_n.t1483 8.126
R5523 out_n.n533 out_n.t867 8.126
R5524 out_n.n534 out_n.t1715 8.126
R5525 out_n.n534 out_n.t1109 8.126
R5526 out_n.n535 out_n.t500 8.126
R5527 out_n.n535 out_n.t1393 8.126
R5528 out_n.n536 out_n.t1442 8.126
R5529 out_n.n536 out_n.t825 8.126
R5530 out_n.n537 out_n.t870 8.126
R5531 out_n.n537 out_n.t262 8.126
R5532 out_n.n538 out_n.t741 8.126
R5533 out_n.n538 out_n.t1633 8.126
R5534 out_n.n539 out_n.t465 8.126
R5535 out_n.n539 out_n.t1354 8.126
R5536 out_n.n520 out_n.t1187 8.126
R5537 out_n.n520 out_n.t612 8.126
R5538 out_n.n521 out_n.t1430 8.126
R5539 out_n.n521 out_n.t850 8.126
R5540 out_n.n522 out_n.t859 8.126
R5541 out_n.n522 out_n.t287 8.126
R5542 out_n.n523 out_n.t298 8.126
R5543 out_n.n523 out_n.t1217 8.126
R5544 out_n.n524 out_n.t534 8.126
R5545 out_n.n524 out_n.t1458 8.126
R5546 out_n.n525 out_n.t811 8.126
R5547 out_n.n525 out_n.t1734 8.126
R5548 out_n.n526 out_n.t1748 8.126
R5549 out_n.n526 out_n.t1170 8.126
R5550 out_n.n527 out_n.t1179 8.126
R5551 out_n.n527 out_n.t605 8.126
R5552 out_n.n528 out_n.t1059 8.126
R5553 out_n.n528 out_n.t484 8.126
R5554 out_n.n529 out_n.t773 8.126
R5555 out_n.n529 out_n.t1695 8.126
R5556 out_n.n510 out_n.t1529 8.126
R5557 out_n.n510 out_n.t952 8.126
R5558 out_n.n511 out_n.t276 8.126
R5559 out_n.n511 out_n.t1195 8.126
R5560 out_n.n512 out_n.t1205 8.126
R5561 out_n.n512 out_n.t627 8.126
R5562 out_n.n513 out_n.t639 8.126
R5563 out_n.n513 out_n.t1555 8.126
R5564 out_n.n514 out_n.t874 8.126
R5565 out_n.n514 out_n.t304 8.126
R5566 out_n.n515 out_n.t1155 8.126
R5567 out_n.n515 out_n.t587 8.126
R5568 out_n.n516 out_n.t598 8.126
R5569 out_n.n516 out_n.t1516 8.126
R5570 out_n.n517 out_n.t1523 8.126
R5571 out_n.n517 out_n.t947 8.126
R5572 out_n.n518 out_n.t1408 8.126
R5573 out_n.n518 out_n.t826 8.126
R5574 out_n.n519 out_n.t1126 8.126
R5575 out_n.n519 out_n.t554 8.126
R5576 out_n.n500 out_n.t985 8.126
R5577 out_n.n500 out_n.t405 8.126
R5578 out_n.n501 out_n.t1231 8.126
R5579 out_n.n501 out_n.t653 8.126
R5580 out_n.n502 out_n.t664 8.126
R5581 out_n.n502 out_n.t1574 8.126
R5582 out_n.n503 out_n.t1584 8.126
R5583 out_n.n503 out_n.t1010 8.126
R5584 out_n.n504 out_n.t328 8.126
R5585 out_n.n504 out_n.t1255 8.126
R5586 out_n.n505 out_n.t613 8.126
R5587 out_n.n505 out_n.t1530 8.126
R5588 out_n.n506 out_n.t1543 8.126
R5589 out_n.n506 out_n.t965 8.126
R5590 out_n.n507 out_n.t976 8.126
R5591 out_n.n507 out_n.t396 8.126
R5592 out_n.n508 out_n.t861 8.126
R5593 out_n.n508 out_n.t288 8.126
R5594 out_n.n509 out_n.t583 8.126
R5595 out_n.n509 out_n.t1500 8.126
R5596 out_n.n490 out_n.t1329 8.126
R5597 out_n.n490 out_n.t753 8.126
R5598 out_n.n491 out_n.t1566 8.126
R5599 out_n.n491 out_n.t994 8.126
R5600 out_n.n492 out_n.t1000 8.126
R5601 out_n.n492 out_n.t427 8.126
R5602 out_n.n493 out_n.t435 8.126
R5603 out_n.n493 out_n.t1362 8.126
R5604 out_n.n494 out_n.t679 8.126
R5605 out_n.n494 out_n.t1592 8.126
R5606 out_n.n495 out_n.t953 8.126
R5607 out_n.n495 out_n.t373 8.126
R5608 out_n.n496 out_n.t387 8.126
R5609 out_n.n496 out_n.t1311 8.126
R5610 out_n.n497 out_n.t1321 8.126
R5611 out_n.n497 out_n.t747 8.126
R5612 out_n.n498 out_n.t1206 8.126
R5613 out_n.n498 out_n.t629 8.126
R5614 out_n.n499 out_n.t918 8.126
R5615 out_n.n499 out_n.t342 8.126
R5616 out_n.n480 out_n.t1678 8.126
R5617 out_n.n480 out_n.t1063 8.126
R5618 out_n.n481 out_n.t416 8.126
R5619 out_n.n481 out_n.t1298 8.126
R5620 out_n.n482 out_n.t1347 8.126
R5621 out_n.n482 out_n.t733 8.126
R5622 out_n.n483 out_n.t780 8.126
R5623 out_n.n483 out_n.t1666 8.126
R5624 out_n.n484 out_n.t1019 8.126
R5625 out_n.n484 out_n.t402 8.126
R5626 out_n.n485 out_n.t1295 8.126
R5627 out_n.n485 out_n.t696 8.126
R5628 out_n.n486 out_n.t737 8.126
R5629 out_n.n486 out_n.t1622 8.126
R5630 out_n.n487 out_n.t1669 8.126
R5631 out_n.n487 out_n.t1060 8.126
R5632 out_n.n488 out_n.t1545 8.126
R5633 out_n.n488 out_n.t936 8.126
R5634 out_n.n489 out_n.t1268 8.126
R5635 out_n.n489 out_n.t663 8.126
R5636 out_n.n470 out_n.t493 8.126
R5637 out_n.n470 out_n.t1418 8.126
R5638 out_n.n471 out_n.t727 8.126
R5639 out_n.n471 out_n.t1647 8.126
R5640 out_n.n472 out_n.t1655 8.126
R5641 out_n.n472 out_n.t1084 8.126
R5642 out_n.n473 out_n.t1095 8.126
R5643 out_n.n473 out_n.t522 8.126
R5644 out_n.n474 out_n.t1327 8.126
R5645 out_n.n474 out_n.t750 8.126
R5646 out_n.n475 out_n.t1611 8.126
R5647 out_n.n475 out_n.t1036 8.126
R5648 out_n.n476 out_n.t1050 8.126
R5649 out_n.n476 out_n.t477 8.126
R5650 out_n.n477 out_n.t485 8.126
R5651 out_n.n477 out_n.t1412 8.126
R5652 out_n.n478 out_n.t358 8.126
R5653 out_n.n478 out_n.t1279 8.126
R5654 out_n.n479 out_n.t1575 8.126
R5655 out_n.n479 out_n.t1001 8.126
R5656 out_n.n460 out_n.t840 8.126
R5657 out_n.n460 out_n.t265 8.126
R5658 out_n.n461 out_n.t1073 8.126
R5659 out_n.n461 out_n.t498 8.126
R5660 out_n.n462 out_n.t510 8.126
R5661 out_n.n462 out_n.t1434 8.126
R5662 out_n.n463 out_n.t1443 8.126
R5663 out_n.n463 out_n.t865 8.126
R5664 out_n.n464 out_n.t1674 8.126
R5665 out_n.n464 out_n.t1103 8.126
R5666 out_n.n465 out_n.t462 8.126
R5667 out_n.n465 out_n.t1391 8.126
R5668 out_n.n466 out_n.t1401 8.126
R5669 out_n.n466 out_n.t820 8.126
R5670 out_n.n467 out_n.t830 8.126
R5671 out_n.n467 out_n.t1756 8.126
R5672 out_n.n468 out_n.t709 8.126
R5673 out_n.n468 out_n.t1626 8.126
R5674 out_n.n469 out_n.t426 8.126
R5675 out_n.n469 out_n.t1348 8.126
R5676 out_n.n450 out_n.t752 8.126
R5677 out_n.n450 out_n.t1677 8.126
R5678 out_n.n451 out_n.t990 8.126
R5679 out_n.n451 out_n.t414 8.126
R5680 out_n.n452 out_n.t424 8.126
R5681 out_n.n452 out_n.t1346 8.126
R5682 out_n.n453 out_n.t1359 8.126
R5683 out_n.n453 out_n.t779 8.126
R5684 out_n.n454 out_n.t1588 8.126
R5685 out_n.n454 out_n.t1016 8.126
R5686 out_n.n455 out_n.t372 8.126
R5687 out_n.n455 out_n.t1294 8.126
R5688 out_n.n456 out_n.t1310 8.126
R5689 out_n.n456 out_n.t735 8.126
R5690 out_n.n457 out_n.t743 8.126
R5691 out_n.n457 out_n.t1667 8.126
R5692 out_n.n458 out_n.t628 8.126
R5693 out_n.n458 out_n.t1544 8.126
R5694 out_n.n459 out_n.t340 8.126
R5695 out_n.n459 out_n.t1267 8.126
R5696 out_n.n440 out_n.t1106 8.126
R5697 out_n.n440 out_n.t531 8.126
R5698 out_n.n441 out_n.t1336 8.126
R5699 out_n.n441 out_n.t759 8.126
R5700 out_n.n442 out_n.t768 8.126
R5701 out_n.n442 out_n.t1691 8.126
R5702 out_n.n443 out_n.t1701 8.126
R5703 out_n.n443 out_n.t1129 8.126
R5704 out_n.n444 out_n.t441 8.126
R5705 out_n.n444 out_n.t1368 8.126
R5706 out_n.n445 out_n.t724 8.126
R5707 out_n.n445 out_n.t1644 8.126
R5708 out_n.n446 out_n.t1657 8.126
R5709 out_n.n446 out_n.t1086 8.126
R5710 out_n.n447 out_n.t1096 8.126
R5711 out_n.n447 out_n.t523 8.126
R5712 out_n.n448 out_n.t968 8.126
R5713 out_n.n448 out_n.t390 8.126
R5714 out_n.n449 out_n.t695 8.126
R5715 out_n.n449 out_n.t1610 8.126
R5716 out_n.n430 out_n.t1456 8.126
R5717 out_n.n430 out_n.t839 8.126
R5718 out_n.n431 out_n.t1684 8.126
R5719 out_n.n431 out_n.t1072 8.126
R5720 out_n.n432 out_n.t1122 8.126
R5721 out_n.n432 out_n.t509 8.126
R5722 out_n.n433 out_n.t559 8.126
R5723 out_n.n433 out_n.t1441 8.126
R5724 out_n.n434 out_n.t786 8.126
R5725 out_n.n434 out_n.t1673 8.126
R5726 out_n.n435 out_n.t1068 8.126
R5727 out_n.n435 out_n.t461 8.126
R5728 out_n.n436 out_n.t513 8.126
R5729 out_n.n436 out_n.t1399 8.126
R5730 out_n.n437 out_n.t1445 8.126
R5731 out_n.n437 out_n.t829 8.126
R5732 out_n.n438 out_n.t1315 8.126
R5733 out_n.n438 out_n.t708 8.126
R5734 out_n.n439 out_n.t1035 8.126
R5735 out_n.n439 out_n.t425 8.126
R5736 out_n.n420 out_n.t263 8.126
R5737 out_n.n420 out_n.t1182 8.126
R5738 out_n.n421 out_n.t497 8.126
R5739 out_n.n421 out_n.t1424 8.126
R5740 out_n.n422 out_n.t1433 8.126
R5741 out_n.n422 out_n.t854 8.126
R5742 out_n.n423 out_n.t862 8.126
R5743 out_n.n423 out_n.t291 8.126
R5744 out_n.n424 out_n.t1102 8.126
R5745 out_n.n424 out_n.t528 8.126
R5746 out_n.n425 out_n.t1390 8.126
R5747 out_n.n425 out_n.t808 8.126
R5748 out_n.n426 out_n.t819 8.126
R5749 out_n.n426 out_n.t1743 8.126
R5750 out_n.n427 out_n.t1753 8.126
R5751 out_n.n427 out_n.t1173 8.126
R5752 out_n.n428 out_n.t1625 8.126
R5753 out_n.n428 out_n.t1055 8.126
R5754 out_n.n429 out_n.t1345 8.126
R5755 out_n.n429 out_n.t769 8.126
R5756 out_n.n410 out_n.t608 8.126
R5757 out_n.n410 out_n.t640 8.126
R5758 out_n.n411 out_n.t846 8.126
R5759 out_n.n411 out_n.t875 8.126
R5760 out_n.n412 out_n.t280 8.126
R5761 out_n.n412 out_n.t310 8.126
R5762 out_n.n413 out_n.t1209 8.126
R5763 out_n.n413 out_n.t1245 8.126
R5764 out_n.n414 out_n.t1450 8.126
R5765 out_n.n414 out_n.t1482 8.126
R5766 out_n.n415 out_n.t1731 8.126
R5767 out_n.n415 out_n.t264 8.126
R5768 out_n.n416 out_n.t1163 8.126
R5769 out_n.n416 out_n.t1196 8.126
R5770 out_n.n417 out_n.t601 8.126
R5771 out_n.n417 out_n.t631 8.126
R5772 out_n.n418 out_n.t479 8.126
R5773 out_n.n418 out_n.t511 8.126
R5774 out_n.n419 out_n.t1692 8.126
R5775 out_n.n419 out_n.t1723 8.126
R5776 out_n.n400 out_n.t1554 8.126
R5777 out_n.n400 out_n.t978 8.126
R5778 out_n.n401 out_n.t303 8.126
R5779 out_n.n401 out_n.t1223 8.126
R5780 out_n.n402 out_n.t1234 8.126
R5781 out_n.n402 out_n.t656 8.126
R5782 out_n.n403 out_n.t668 8.126
R5783 out_n.n403 out_n.t1580 8.126
R5784 out_n.n404 out_n.t896 8.126
R5785 out_n.n404 out_n.t324 8.126
R5786 out_n.n405 out_n.t1183 8.126
R5787 out_n.n405 out_n.t610 8.126
R5788 out_n.n406 out_n.t619 8.126
R5789 out_n.n406 out_n.t1537 8.126
R5790 out_n.n407 out_n.t1546 8.126
R5791 out_n.n407 out_n.t969 8.126
R5792 out_n.n408 out_n.t1435 8.126
R5793 out_n.n408 out_n.t856 8.126
R5794 out_n.n409 out_n.t1147 8.126
R5795 out_n.n409 out_n.t578 8.126
R5796 out_n.n390 out_n.t398 8.126
R5797 out_n.n390 out_n.t1323 8.126
R5798 out_n.n391 out_n.t648 8.126
R5799 out_n.n391 out_n.t1561 8.126
R5800 out_n.n392 out_n.t1570 8.126
R5801 out_n.n392 out_n.t995 8.126
R5802 out_n.n393 out_n.t1005 8.126
R5803 out_n.n393 out_n.t429 8.126
R5804 out_n.n394 out_n.t1250 8.126
R5805 out_n.n394 out_n.t674 8.126
R5806 out_n.n395 out_n.t1527 8.126
R5807 out_n.n395 out_n.t949 8.126
R5808 out_n.n396 out_n.t958 8.126
R5809 out_n.n396 out_n.t381 8.126
R5810 out_n.n397 out_n.t391 8.126
R5811 out_n.n397 out_n.t1316 8.126
R5812 out_n.n398 out_n.t284 8.126
R5813 out_n.n398 out_n.t1201 8.126
R5814 out_n.n399 out_n.t1498 8.126
R5815 out_n.n399 out_n.t915 8.126
R5816 out_n.n380 out_n.t1361 8.126
R5817 out_n.n380 out_n.t1636 8.126
R5818 out_n.n381 out_n.t1591 8.126
R5819 out_n.n381 out_n.t371 8.126
R5820 out_n.n382 out_n.t1024 8.126
R5821 out_n.n382 out_n.t1302 8.126
R5822 out_n.n383 out_n.t459 8.126
R5823 out_n.n383 out_n.t736 8.126
R5824 out_n.n384 out_n.t700 8.126
R5825 out_n.n384 out_n.t974 8.126
R5826 out_n.n385 out_n.t979 8.126
R5827 out_n.n385 out_n.t1266 8.126
R5828 out_n.n386 out_n.t418 8.126
R5829 out_n.n386 out_n.t702 8.126
R5830 out_n.n387 out_n.t1351 8.126
R5831 out_n.n387 out_n.t1627 8.126
R5832 out_n.n388 out_n.t1236 8.126
R5833 out_n.n388 out_n.t1511 8.126
R5834 out_n.n389 out_n.t942 8.126
R5835 out_n.n389 out_n.t1235 8.126
R5836 out_n.n370 out_n.t1061 8.126
R5837 out_n.n370 out_n.t490 8.126
R5838 out_n.n371 out_n.t1293 8.126
R5839 out_n.n371 out_n.t722 8.126
R5840 out_n.n372 out_n.t730 8.126
R5841 out_n.n372 out_n.t1650 8.126
R5842 out_n.n373 out_n.t1658 8.126
R5843 out_n.n373 out_n.t1087 8.126
R5844 out_n.n374 out_n.t395 8.126
R5845 out_n.n374 out_n.t1319 8.126
R5846 out_n.n375 out_n.t694 8.126
R5847 out_n.n375 out_n.t1607 8.126
R5848 out_n.n376 out_n.t1618 8.126
R5849 out_n.n376 out_n.t1044 8.126
R5850 out_n.n377 out_n.t1056 8.126
R5851 out_n.n377 out_n.t481 8.126
R5852 out_n.n378 out_n.t929 8.126
R5853 out_n.n378 out_n.t354 8.126
R5854 out_n.n379 out_n.t655 8.126
R5855 out_n.n379 out_n.t1569 8.126
R5856 out_n.n360 out_n.t1415 8.126
R5857 out_n.n360 out_n.t1444 8.126
R5858 out_n.n361 out_n.t1643 8.126
R5859 out_n.n361 out_n.t1675 8.126
R5860 out_n.n362 out_n.t1076 8.126
R5861 out_n.n362 out_n.t1113 8.126
R5862 out_n.n363 out_n.t514 8.126
R5863 out_n.n363 out_n.t547 8.126
R5864 out_n.n364 out_n.t742 8.126
R5865 out_n.n364 out_n.t775 8.126
R5866 out_n.n365 out_n.t1032 8.126
R5867 out_n.n365 out_n.t1062 8.126
R5868 out_n.n366 out_n.t470 8.126
R5869 out_n.n366 out_n.t499 8.126
R5870 out_n.n367 out_n.t1406 8.126
R5871 out_n.n367 out_n.t1436 8.126
R5872 out_n.n368 out_n.t1276 8.126
R5873 out_n.n368 out_n.t1303 8.126
R5874 out_n.n369 out_n.t996 8.126
R5875 out_n.n369 out_n.t1026 8.126
R5876 out_n.n350 out_n.t864 8.126
R5877 out_n.n350 out_n.t292 8.126
R5878 out_n.n351 out_n.t1105 8.126
R5879 out_n.n351 out_n.t530 8.126
R5880 out_n.n352 out_n.t539 8.126
R5881 out_n.n352 out_n.t1461 8.126
R5882 out_n.n353 out_n.t1470 8.126
R5883 out_n.n353 out_n.t886 8.126
R5884 out_n.n354 out_n.t1699 8.126
R5885 out_n.n354 out_n.t1127 8.126
R5886 out_n.n355 out_n.t491 8.126
R5887 out_n.n355 out_n.t1416 8.126
R5888 out_n.n356 out_n.t1426 8.126
R5889 out_n.n356 out_n.t847 8.126
R5890 out_n.n357 out_n.t857 8.126
R5891 out_n.n357 out_n.t285 8.126
R5892 out_n.n358 out_n.t731 8.126
R5893 out_n.n358 out_n.t1653 8.126
R5894 out_n.n359 out_n.t452 8.126
R5895 out_n.n359 out_n.t1377 8.126
R5896 out_n.n340 out_n.t1213 8.126
R5897 out_n.n340 out_n.t635 8.126
R5898 out_n.n341 out_n.t1455 8.126
R5899 out_n.n341 out_n.t872 8.126
R5900 out_n.n342 out_n.t880 8.126
R5901 out_n.n342 out_n.t305 8.126
R5902 out_n.n343 out_n.t313 8.126
R5903 out_n.n343 out_n.t1240 8.126
R5904 out_n.n344 out_n.t555 8.126
R5905 out_n.n344 out_n.t1475 8.126
R5906 out_n.n345 out_n.t835 8.126
R5907 out_n.n345 out_n.t1759 8.126
R5908 out_n.n346 out_n.t272 8.126
R5909 out_n.n346 out_n.t1190 8.126
R5910 out_n.n347 out_n.t1202 8.126
R5911 out_n.n347 out_n.t625 8.126
R5912 out_n.n348 out_n.t1080 8.126
R5913 out_n.n348 out_n.t506 8.126
R5914 out_n.n349 out_n.t795 8.126
R5915 out_n.n349 out_n.t1719 8.126
R5916 out_n.n330 out_n.t670 8.126
R5917 out_n.n330 out_n.t938 8.126
R5918 out_n.n331 out_n.t898 8.126
R5919 out_n.n331 out_n.t1180 8.126
R5920 out_n.n332 out_n.t334 8.126
R5921 out_n.n332 out_n.t614 8.126
R5922 out_n.n333 out_n.t1263 8.126
R5923 out_n.n333 out_n.t1538 8.126
R5924 out_n.n334 out_n.t1503 8.126
R5925 out_n.n334 out_n.t289 8.126
R5926 out_n.n335 out_n.t293 8.126
R5927 out_n.n335 out_n.t576 8.126
R5928 out_n.n336 out_n.t1226 8.126
R5929 out_n.n336 out_n.t1506 8.126
R5930 out_n.n337 out_n.t661 8.126
R5931 out_n.n337 out_n.t930 8.126
R5932 out_n.n338 out_n.t540 8.126
R5933 out_n.n338 out_n.t814 8.126
R5934 out_n.n339 out_n.t1751 8.126
R5935 out_n.n339 out_n.t538 8.126
R5936 out_n.n320 out_n.t360 8.126
R5937 out_n.n320 out_n.t1284 8.126
R5938 out_n.n321 out_n.t606 8.126
R5939 out_n.n321 out_n.t1524 8.126
R5940 out_n.n322 out_n.t1531 8.126
R5941 out_n.n322 out_n.t954 8.126
R5942 out_n.n323 out_n.t959 8.126
R5943 out_n.n323 out_n.t382 8.126
R5944 out_n.n324 out_n.t1207 8.126
R5945 out_n.n324 out_n.t630 8.126
R5946 out_n.n325 out_n.t1497 8.126
R5947 out_n.n325 out_n.t913 8.126
R5948 out_n.n326 out_n.t924 8.126
R5949 out_n.n326 out_n.t347 8.126
R5950 out_n.n327 out_n.t356 8.126
R5951 out_n.n327 out_n.t1278 8.126
R5952 out_n.n328 out_n.t1737 8.126
R5953 out_n.n328 out_n.t1159 8.126
R5954 out_n.n329 out_n.t1462 8.126
R5955 out_n.n329 out_n.t879 8.126
R5956 out_n.n310 out_n.t1314 8.126
R5957 out_n.n310 out_n.t739 8.126
R5958 out_n.n311 out_n.t1553 8.126
R5959 out_n.n311 out_n.t977 8.126
R5960 out_n.n312 out_n.t987 8.126
R5961 out_n.n312 out_n.t407 8.126
R5962 out_n.n313 out_n.t420 8.126
R5963 out_n.n313 out_n.t1339 8.126
R5964 out_n.n314 out_n.t667 8.126
R5965 out_n.n314 out_n.t1577 8.126
R5966 out_n.n315 out_n.t939 8.126
R5967 out_n.n315 out_n.t361 8.126
R5968 out_n.n316 out_n.t374 8.126
R5969 out_n.n316 out_n.t1296 8.126
R5970 out_n.n317 out_n.t1305 8.126
R5971 out_n.n317 out_n.t732 8.126
R5972 out_n.n318 out_n.t1189 8.126
R5973 out_n.n318 out_n.t616 8.126
R5974 out_n.n319 out_n.t907 8.126
R5975 out_n.n319 out_n.t333 8.126
R5976 out_n.n300 out_n.t1660 8.126
R5977 out_n.n300 out_n.t1089 8.126
R5978 out_n.n301 out_n.t397 8.126
R5979 out_n.n301 out_n.t1322 8.126
R5980 out_n.n302 out_n.t1331 8.126
R5981 out_n.n302 out_n.t754 8.126
R5982 out_n.n303 out_n.t762 8.126
R5983 out_n.n303 out_n.t1686 8.126
R5984 out_n.n304 out_n.t1002 8.126
R5985 out_n.n304 out_n.t428 8.126
R5986 out_n.n305 out_n.t1285 8.126
R5987 out_n.n305 out_n.t714 8.126
R5988 out_n.n306 out_n.t725 8.126
R5989 out_n.n306 out_n.t1645 8.126
R5990 out_n.n307 out_n.t1654 8.126
R5991 out_n.n307 out_n.t1083 8.126
R5992 out_n.n308 out_n.t1534 8.126
R5993 out_n.n308 out_n.t956 8.126
R5994 out_n.n309 out_n.t1258 8.126
R5995 out_n.n309 out_n.t683 8.126
R5996 out_n.n290 out_n.t517 8.126
R5997 out_n.n290 out_n.t551 8.126
R5998 out_n.n291 out_n.t746 8.126
R5999 out_n.n291 out_n.t778 8.126
R6000 out_n.n292 out_n.t1679 8.126
R6001 out_n.n292 out_n.t1710 8.126
R6002 out_n.n293 out_n.t1116 8.126
R6003 out_n.n293 out_n.t1143 8.126
R6004 out_n.n294 out_n.t1349 8.126
R6005 out_n.n294 out_n.t1385 8.126
R6006 out_n.n295 out_n.t1631 8.126
R6007 out_n.n295 out_n.t1663 8.126
R6008 out_n.n296 out_n.t1069 8.126
R6009 out_n.n296 out_n.t1107 8.126
R6010 out_n.n297 out_n.t507 8.126
R6011 out_n.n297 out_n.t542 8.126
R6012 out_n.n298 out_n.t376 8.126
R6013 out_n.n298 out_n.t408 8.126
R6014 out_n.n299 out_n.t1596 8.126
R6015 out_n.n299 out_n.t1623 8.126
R6016 out_n.n280 out_n.t1473 8.126
R6017 out_n.n280 out_n.t1745 8.126
R6018 out_n.n281 out_n.t1702 8.126
R6019 out_n.n281 out_n.t486 8.126
R6020 out_n.n282 out_n.t1136 8.126
R6021 out_n.n282 out_n.t1419 8.126
R6022 out_n.n283 out_n.t572 8.126
R6023 out_n.n283 out_n.t848 8.126
R6024 out_n.n284 out_n.t802 8.126
R6025 out_n.n284 out_n.t1085 8.126
R6026 out_n.n285 out_n.t1091 8.126
R6027 out_n.n285 out_n.t1376 8.126
R6028 out_n.n286 out_n.t532 8.126
R6029 out_n.n286 out_n.t809 8.126
R6030 out_n.n287 out_n.t1464 8.126
R6031 out_n.n287 out_n.t1739 8.126
R6032 out_n.n288 out_n.t1332 8.126
R6033 out_n.n288 out_n.t1613 8.126
R6034 out_n.n289 out_n.t1054 8.126
R6035 out_n.n289 out_n.t1330 8.126
R6036 out_n.n270 out_n.t1166 8.126
R6037 out_n.n270 out_n.t595 8.126
R6038 out_n.n271 out_n.t1410 8.126
R6039 out_n.n271 out_n.t831 8.126
R6040 out_n.n272 out_n.t841 8.126
R6041 out_n.n272 out_n.t266 8.126
R6042 out_n.n273 out_n.t275 8.126
R6043 out_n.n273 out_n.t1192 8.126
R6044 out_n.n274 out_n.t512 8.126
R6045 out_n.n274 out_n.t1437 8.126
R6046 out_n.n275 out_n.t793 8.126
R6047 out_n.n275 out_n.t1717 8.126
R6048 out_n.n276 out_n.t1733 8.126
R6049 out_n.n276 out_n.t1154 8.126
R6050 out_n.n277 out_n.t1161 8.126
R6051 out_n.n277 out_n.t591 8.126
R6052 out_n.n278 out_n.t1038 8.126
R6053 out_n.n278 out_n.t464 8.126
R6054 out_n.n279 out_n.t755 8.126
R6055 out_n.n279 out_n.t1681 8.126
R6056 out_n.n260 out_n.t623 8.126
R6057 out_n.n260 out_n.t1541 8.126
R6058 out_n.n261 out_n.t863 8.126
R6059 out_n.n261 out_n.t290 8.126
R6060 out_n.n262 out_n.t299 8.126
R6061 out_n.n262 out_n.t1218 8.126
R6062 out_n.n263 out_n.t1227 8.126
R6063 out_n.n263 out_n.t650 8.126
R6064 out_n.n264 out_n.t1469 8.126
R6065 out_n.n264 out_n.t884 8.126
R6066 out_n.n265 out_n.t1746 8.126
R6067 out_n.n265 out_n.t1167 8.126
R6068 out_n.n266 out_n.t1184 8.126
R6069 out_n.n266 out_n.t611 8.126
R6070 out_n.n267 out_n.t617 8.126
R6071 out_n.n267 out_n.t1535 8.126
R6072 out_n.n268 out_n.t496 8.126
R6073 out_n.n268 out_n.t1422 8.126
R6074 out_n.n269 out_n.t1712 8.126
R6075 out_n.n269 out_n.t1135 8.126
R6076 out_n.n250 out_n.t961 8.126
R6077 out_n.n250 out_n.t383 8.126
R6078 out_n.n251 out_n.t1208 8.126
R6079 out_n.n251 out_n.t632 8.126
R6080 out_n.n252 out_n.t643 8.126
R6081 out_n.n252 out_n.t1557 8.126
R6082 out_n.n253 out_n.t1563 8.126
R6083 out_n.n253 out_n.t989 8.126
R6084 out_n.n254 out_n.t311 8.126
R6085 out_n.n254 out_n.t1239 8.126
R6086 out_n.n255 out_n.t597 8.126
R6087 out_n.n255 out_n.t1515 8.126
R6088 out_n.n256 out_n.t1528 8.126
R6089 out_n.n256 out_n.t950 8.126
R6090 out_n.n257 out_n.t957 8.126
R6091 out_n.n257 out_n.t379 8.126
R6092 out_n.n258 out_n.t842 8.126
R6093 out_n.n258 out_n.t267 8.126
R6094 out_n.n259 out_n.t566 8.126
R6095 out_n.n259 out_n.t1486 8.126
R6096 out_n.n240 out_n.t1308 8.126
R6097 out_n.n240 out_n.t1342 8.126
R6098 out_n.n241 out_n.t1548 8.126
R6099 out_n.n241 out_n.t1579 8.126
R6100 out_n.n242 out_n.t981 8.126
R6101 out_n.n242 out_n.t1012 8.126
R6102 out_n.n243 out_n.t411 8.126
R6103 out_n.n243 out_n.t445 8.126
R6104 out_n.n244 out_n.t659 8.126
R6105 out_n.n244 out_n.t688 8.126
R6106 out_n.n245 out_n.t935 8.126
R6107 out_n.n245 out_n.t962 8.126
R6108 out_n.n246 out_n.t368 8.126
R6109 out_n.n246 out_n.t400 8.126
R6110 out_n.n247 out_n.t1300 8.126
R6111 out_n.n247 out_n.t1334 8.126
R6112 out_n.n248 out_n.t1185 8.126
R6113 out_n.n248 out_n.t1221 8.126
R6114 out_n.n249 out_n.t900 8.126
R6115 out_n.n249 out_n.t927 8.126
R6116 out_n.n230 out_n.t766 8.126
R6117 out_n.n230 out_n.t1047 8.126
R6118 out_n.n231 out_n.t1004 8.126
R6119 out_n.n231 out_n.t1281 8.126
R6120 out_n.n232 out_n.t437 8.126
R6121 out_n.n232 out_n.t717 8.126
R6122 out_n.n233 out_n.t1373 8.126
R6123 out_n.n233 out_n.t1646 8.126
R6124 out_n.n234 out_n.t1601 8.126
R6125 out_n.n234 out_n.t380 8.126
R6126 out_n.n235 out_n.t385 8.126
R6127 out_n.n235 out_n.t680 8.126
R6128 out_n.n236 out_n.t1325 8.126
R6129 out_n.n236 out_n.t1609 8.126
R6130 out_n.n237 out_n.t757 8.126
R6131 out_n.n237 out_n.t1040 8.126
R6132 out_n.n238 out_n.t644 8.126
R6133 out_n.n238 out_n.t917 8.126
R6134 out_n.n239 out_n.t353 8.126
R6135 out_n.n239 out_n.t642 8.126
R6136 out_n.n220 out_n.t473 8.126
R6137 out_n.n220 out_n.t1360 8.126
R6138 out_n.n221 out_n.t711 8.126
R6139 out_n.n221 out_n.t1590 8.126
R6140 out_n.n222 out_n.t1637 8.126
R6141 out_n.n222 out_n.t1025 8.126
R6142 out_n.n223 out_n.t1071 8.126
R6143 out_n.n223 out_n.t460 8.126
R6144 out_n.n224 out_n.t1304 8.126
R6145 out_n.n224 out_n.t701 8.126
R6146 out_n.n225 out_n.t1593 8.126
R6147 out_n.n225 out_n.t980 8.126
R6148 out_n.n226 out_n.t1034 8.126
R6149 out_n.n226 out_n.t419 8.126
R6150 out_n.n227 out_n.t466 8.126
R6151 out_n.n227 out_n.t1352 8.126
R6152 out_n.n228 out_n.t341 8.126
R6153 out_n.n228 out_n.t1237 8.126
R6154 out_n.n229 out_n.t1556 8.126
R6155 out_n.n229 out_n.t943 8.126
R6156 out_n.n210 out_n.t781 8.126
R6157 out_n.n210 out_n.t1703 8.126
R6158 out_n.n211 out_n.t1018 8.126
R6159 out_n.n211 out_n.t442 8.126
R6160 out_n.n212 out_n.t451 8.126
R6161 out_n.n212 out_n.t1378 8.126
R6162 out_n.n213 out_n.t1387 8.126
R6163 out_n.n213 out_n.t805 8.126
R6164 out_n.n214 out_n.t1615 8.126
R6165 out_n.n214 out_n.t1041 8.126
R6166 out_n.n215 out_n.t399 8.126
R6167 out_n.n215 out_n.t1324 8.126
R6168 out_n.n216 out_n.t1338 8.126
R6169 out_n.n216 out_n.t761 8.126
R6170 out_n.n217 out_n.t770 8.126
R6171 out_n.n217 out_n.t1694 8.126
R6172 out_n.n218 out_n.t657 8.126
R6173 out_n.n218 out_n.t1572 8.126
R6174 out_n.n219 out_n.t364 8.126
R6175 out_n.n219 out_n.t1288 8.126
R6176 out_n.n200 out_n.t1130 8.126
R6177 out_n.n200 out_n.t560 8.126
R6178 out_n.n201 out_n.t1369 8.126
R6179 out_n.n201 out_n.t787 8.126
R6180 out_n.n202 out_n.t794 8.126
R6181 out_n.n202 out_n.t1718 8.126
R6182 out_n.n203 out_n.t1728 8.126
R6183 out_n.n203 out_n.t1151 8.126
R6184 out_n.n204 out_n.t467 8.126
R6185 out_n.n204 out_n.t1394 8.126
R6186 out_n.n205 out_n.t748 8.126
R6187 out_n.n205 out_n.t1670 8.126
R6188 out_n.n206 out_n.t1685 8.126
R6189 out_n.n206 out_n.t1114 8.126
R6190 out_n.n207 out_n.t1124 8.126
R6191 out_n.n207 out_n.t552 8.126
R6192 out_n.n208 out_n.t998 8.126
R6193 out_n.n208 out_n.t422 8.126
R6194 out_n.n209 out_n.t716 8.126
R6195 out_n.n209 out_n.t1635 8.126
R6196 out_n.n190 out_n.t586 8.126
R6197 out_n.n190 out_n.t1505 8.126
R6198 out_n.n191 out_n.t818 8.126
R6199 out_n.n191 out_n.t1742 8.126
R6200 out_n.n192 out_n.t1750 8.126
R6201 out_n.n192 out_n.t1172 8.126
R6202 out_n.n193 out_n.t1181 8.126
R6203 out_n.n193 out_n.t607 8.126
R6204 out_n.n194 out_n.t1423 8.126
R6205 out_n.n194 out_n.t843 8.126
R6206 out_n.n195 out_n.t1704 8.126
R6207 out_n.n195 out_n.t1131 8.126
R6208 out_n.n196 out_n.t1142 8.126
R6209 out_n.n196 out_n.t571 8.126
R6210 out_n.n197 out_n.t580 8.126
R6211 out_n.n197 out_n.t1499 8.126
R6212 out_n.n198 out_n.t453 8.126
R6213 out_n.n198 out_n.t1379 8.126
R6214 out_n.n199 out_n.t1665 8.126
R6215 out_n.n199 out_n.t1094 8.126
R6216 out_n.n180 out_n.t923 8.126
R6217 out_n.n180 out_n.t1212 8.126
R6218 out_n.n181 out_n.t1162 8.126
R6219 out_n.n181 out_n.t1452 8.126
R6220 out_n.n182 out_n.t599 8.126
R6221 out_n.n182 out_n.t878 8.126
R6222 out_n.n183 out_n.t1525 8.126
R6223 out_n.n183 out_n.t314 8.126
R6224 out_n.n184 out_n.t269 8.126
R6225 out_n.n184 out_n.t556 8.126
R6226 out_n.n185 out_n.t561 8.126
R6227 out_n.n185 out_n.t836 8.126
R6228 out_n.n186 out_n.t1492 8.126
R6229 out_n.n186 out_n.t273 8.126
R6230 out_n.n187 out_n.t916 8.126
R6231 out_n.n187 out_n.t1203 8.126
R6232 out_n.n188 out_n.t798 8.126
R6233 out_n.n188 out_n.t1081 8.126
R6234 out_n.n189 out_n.t521 8.126
R6235 out_n.n189 out_n.t797 8.126
R6236 out_n.n170 out_n.t634 8.126
R6237 out_n.n170 out_n.t669 8.126
R6238 out_n.n171 out_n.t871 8.126
R6239 out_n.n171 out_n.t897 8.126
R6240 out_n.n172 out_n.t306 8.126
R6241 out_n.n172 out_n.t335 8.126
R6242 out_n.n173 out_n.t1241 8.126
R6243 out_n.n173 out_n.t1264 8.126
R6244 out_n.n174 out_n.t1476 8.126
R6245 out_n.n174 out_n.t1502 8.126
R6246 out_n.n175 out_n.t1760 8.126
R6247 out_n.n175 out_n.t294 8.126
R6248 out_n.n176 out_n.t1191 8.126
R6249 out_n.n176 out_n.t1225 8.126
R6250 out_n.n177 out_n.t626 8.126
R6251 out_n.n177 out_n.t658 8.126
R6252 out_n.n178 out_n.t504 8.126
R6253 out_n.n178 out_n.t541 8.126
R6254 out_n.n179 out_n.t1720 8.126
R6255 out_n.n179 out_n.t1752 8.126
R6256 out_n.n160 out_n.t1581 8.126
R6257 out_n.n160 out_n.t1006 8.126
R6258 out_n.n161 out_n.t325 8.126
R6259 out_n.n161 out_n.t1251 8.126
R6260 out_n.n162 out_n.t1257 8.126
R6261 out_n.n162 out_n.t682 8.126
R6262 out_n.n163 out_n.t691 8.126
R6263 out_n.n163 out_n.t1604 8.126
R6264 out_n.n164 out_n.t920 8.126
R6265 out_n.n164 out_n.t343 8.126
R6266 out_n.n165 out_n.t1214 8.126
R6267 out_n.n165 out_n.t636 8.126
R6268 out_n.n166 out_n.t649 8.126
R6269 out_n.n166 out_n.t1562 8.126
R6270 out_n.n167 out_n.t1573 8.126
R6271 out_n.n167 out_n.t999 8.126
R6272 out_n.n168 out_n.t1463 8.126
R6273 out_n.n168 out_n.t882 8.126
R6274 out_n.n169 out_n.t1171 8.126
R6275 out_n.n169 out_n.t600 8.126
R6276 out_n.n150 out_n.t431 8.126
R6277 out_n.n150 out_n.t1355 8.126
R6278 out_n.n151 out_n.t675 8.126
R6279 out_n.n151 out_n.t1585 8.126
R6280 out_n.n152 out_n.t1595 8.126
R6281 out_n.n152 out_n.t1020 8.126
R6282 out_n.n153 out_n.t1029 8.126
R6283 out_n.n153 out_n.t456 8.126
R6284 out_n.n154 out_n.t1270 8.126
R6285 out_n.n154 out_n.t697 8.126
R6286 out_n.n155 out_n.t1551 8.126
R6287 out_n.n155 out_n.t972 8.126
R6288 out_n.n156 out_n.t988 8.126
R6289 out_n.n156 out_n.t410 8.126
R6290 out_n.n157 out_n.t423 8.126
R6291 out_n.n157 out_n.t1344 8.126
R6292 out_n.n158 out_n.t307 8.126
R6293 out_n.n158 out_n.t1230 8.126
R6294 out_n.n159 out_n.t1517 8.126
R6295 out_n.n159 out_n.t937 8.126
R6296 out_n.n140 out_n.t1389 8.126
R6297 out_n.n140 out_n.t807 8.126
R6298 out_n.n141 out_n.t1617 8.126
R6299 out_n.n141 out_n.t1043 8.126
R6300 out_n.n142 out_n.t1051 8.126
R6301 out_n.n142 out_n.t475 8.126
R6302 out_n.n143 out_n.t487 8.126
R6303 out_n.n143 out_n.t1413 8.126
R6304 out_n.n144 out_n.t719 8.126
R6305 out_n.n144 out_n.t1639 8.126
R6306 out_n.n145 out_n.t1007 8.126
R6307 out_n.n145 out_n.t432 8.126
R6308 out_n.n146 out_n.t443 8.126
R6309 out_n.n146 out_n.t1370 8.126
R6310 out_n.n147 out_n.t1381 8.126
R6311 out_n.n147 out_n.t799 8.126
R6312 out_n.n148 out_n.t1260 8.126
R6313 out_n.n148 out_n.t684 8.126
R6314 out_n.n149 out_n.t967 8.126
R6315 out_n.n149 out_n.t389 8.126
R6316 out_n.n130 out_n.t1730 8.126
R6317 out_n.n130 out_n.t516 8.126
R6318 out_n.n131 out_n.t469 8.126
R6319 out_n.n131 out_n.t745 8.126
R6320 out_n.n132 out_n.t1403 8.126
R6321 out_n.n132 out_n.t1680 8.126
R6322 out_n.n133 out_n.t832 8.126
R6323 out_n.n133 out_n.t1115 8.126
R6324 out_n.n134 out_n.t1066 8.126
R6325 out_n.n134 out_n.t1350 8.126
R6326 out_n.n135 out_n.t1356 8.126
R6327 out_n.n135 out_n.t1632 8.126
R6328 out_n.n136 out_n.t789 8.126
R6329 out_n.n136 out_n.t1070 8.126
R6330 out_n.n137 out_n.t1722 8.126
R6331 out_n.n137 out_n.t508 8.126
R6332 out_n.n138 out_n.t1597 8.126
R6333 out_n.n138 out_n.t377 8.126
R6334 out_n.n139 out_n.t1313 8.126
R6335 out_n.n139 out_n.t1594 8.126
R6336 out_n.n120 out_n.t549 8.126
R6337 out_n.n120 out_n.t1472 8.126
R6338 out_n.n121 out_n.t777 8.126
R6339 out_n.n121 out_n.t1700 8.126
R6340 out_n.n122 out_n.t1711 8.126
R6341 out_n.n122 out_n.t1137 8.126
R6342 out_n.n123 out_n.t1144 8.126
R6343 out_n.n123 out_n.t573 8.126
R6344 out_n.n124 out_n.t1386 8.126
R6345 out_n.n124 out_n.t803 8.126
R6346 out_n.n125 out_n.t1661 8.126
R6347 out_n.n125 out_n.t1092 8.126
R6348 out_n.n126 out_n.t1108 8.126
R6349 out_n.n126 out_n.t533 8.126
R6350 out_n.n127 out_n.t543 8.126
R6351 out_n.n127 out_n.t1465 8.126
R6352 out_n.n128 out_n.t409 8.126
R6353 out_n.n128 out_n.t1333 8.126
R6354 out_n.n129 out_n.t1624 8.126
R6355 out_n.n129 out_n.t1053 8.126
R6356 out_n.n110 out_n.t888 8.126
R6357 out_n.n110 out_n.t316 8.126
R6358 out_n.n111 out_n.t1128 8.126
R6359 out_n.n111 out_n.t558 8.126
R6360 out_n.n112 out_n.t565 8.126
R6361 out_n.n112 out_n.t1485 8.126
R6362 out_n.n113 out_n.t1493 8.126
R6363 out_n.n113 out_n.t909 8.126
R6364 out_n.n114 out_n.t1726 8.126
R6365 out_n.n114 out_n.t1148 8.126
R6366 out_n.n115 out_n.t518 8.126
R6367 out_n.n115 out_n.t1440 8.126
R6368 out_n.n116 out_n.t1457 8.126
R6369 out_n.n116 out_n.t873 8.126
R6370 out_n.n117 out_n.t883 8.126
R6371 out_n.n117 out_n.t309 8.126
R6372 out_n.n118 out_n.t756 8.126
R6373 out_n.n118 out_n.t1682 8.126
R6374 out_n.n119 out_n.t478 8.126
R6375 out_n.n119 out_n.t1402 8.126
R6376 out_n.n100 out_n.t1242 8.126
R6377 out_n.n100 out_n.t1265 8.126
R6378 out_n.n101 out_n.t1477 8.126
R6379 out_n.n101 out_n.t1504 8.126
R6380 out_n.n102 out_n.t901 8.126
R6381 out_n.n102 out_n.t928 8.126
R6382 out_n.n103 out_n.t337 8.126
R6383 out_n.n103 out_n.t359 8.126
R6384 out_n.n104 out_n.t579 8.126
R6385 out_n.n104 out_n.t604 8.126
R6386 out_n.n105 out_n.t860 8.126
R6387 out_n.n105 out_n.t890 8.126
R6388 out_n.n106 out_n.t301 8.126
R6389 out_n.n106 out_n.t326 8.126
R6390 out_n.n107 out_n.t1233 8.126
R6391 out_n.n107 out_n.t1261 8.126
R6392 out_n.n108 out_n.t1110 8.126
R6393 out_n.n108 out_n.t1138 8.126
R6394 out_n.n109 out_n.t822 8.126
R6395 out_n.n109 out_n.t855 8.126
R6396 out_n.n90 out_n.t693 8.126
R6397 out_n.n90 out_n.t1606 8.126
R6398 out_n.n91 out_n.t922 8.126
R6399 out_n.n91 out_n.t346 8.126
R6400 out_n.n92 out_n.t351 8.126
R6401 out_n.n92 out_n.t1273 8.126
R6402 out_n.n93 out_n.t1282 8.126
R6403 out_n.n93 out_n.t712 8.126
R6404 out_n.n94 out_n.t1522 8.126
R6405 out_n.n94 out_n.t945 8.126
R6406 out_n.n95 out_n.t317 8.126
R6407 out_n.n95 out_n.t1244 8.126
R6408 out_n.n96 out_n.t1253 8.126
R6409 out_n.n96 out_n.t676 8.126
R6410 out_n.n97 out_n.t687 8.126
R6411 out_n.n97 out_n.t1599 8.126
R6412 out_n.n98 out_n.t567 8.126
R6413 out_n.n98 out_n.t1487 8.126
R6414 out_n.n99 out_n.t283 8.126
R6415 out_n.n99 out_n.t1199 8.126
R6416 out_n.n80 out_n.t1031 8.126
R6417 out_n.n80 out_n.t1306 8.126
R6418 out_n.n81 out_n.t1271 8.126
R6419 out_n.n81 out_n.t1547 8.126
R6420 out_n.n82 out_n.t706 8.126
R6421 out_n.n82 out_n.t982 8.126
R6422 out_n.n83 out_n.t1630 8.126
R6423 out_n.n83 out_n.t412 8.126
R6424 out_n.n84 out_n.t365 8.126
R6425 out_n.n84 out_n.t660 8.126
R6426 out_n.n85 out_n.t665 8.126
R6427 out_n.n85 out_n.t934 8.126
R6428 out_n.n86 out_n.t1586 8.126
R6429 out_n.n86 out_n.t369 8.126
R6430 out_n.n87 out_n.t1022 8.126
R6431 out_n.n87 out_n.t1301 8.126
R6432 out_n.n88 out_n.t902 8.126
R6433 out_n.n88 out_n.t1186 8.126
R6434 out_n.n89 out_n.t622 8.126
R6435 out_n.n89 out_n.t899 8.126
R6436 out_n.n70 out_n.t1341 8.126
R6437 out_n.n70 out_n.t765 8.126
R6438 out_n.n71 out_n.t1578 8.126
R6439 out_n.n71 out_n.t1003 8.126
R6440 out_n.n72 out_n.t1013 8.126
R6441 out_n.n72 out_n.t436 8.126
R6442 out_n.n73 out_n.t446 8.126
R6443 out_n.n73 out_n.t1372 8.126
R6444 out_n.n74 out_n.t689 8.126
R6445 out_n.n74 out_n.t1602 8.126
R6446 out_n.n75 out_n.t963 8.126
R6447 out_n.n75 out_n.t386 8.126
R6448 out_n.n76 out_n.t401 8.126
R6449 out_n.n76 out_n.t1326 8.126
R6450 out_n.n77 out_n.t1335 8.126
R6451 out_n.n77 out_n.t758 8.126
R6452 out_n.n78 out_n.t1220 8.126
R6453 out_n.n78 out_n.t645 8.126
R6454 out_n.n79 out_n.t926 8.126
R6455 out_n.n79 out_n.t350 8.126
R6456 out_n.n60 out_n.t1688 8.126
R6457 out_n.n60 out_n.t1118 8.126
R6458 out_n.n61 out_n.t430 8.126
R6459 out_n.n61 out_n.t1353 8.126
R6460 out_n.n62 out_n.t1363 8.126
R6461 out_n.n62 out_n.t782 8.126
R6462 out_n.n63 out_n.t790 8.126
R6463 out_n.n63 out_n.t1714 8.126
R6464 out_n.n64 out_n.t1027 8.126
R6465 out_n.n64 out_n.t454 8.126
R6466 out_n.n65 out_n.t1309 8.126
R6467 out_n.n65 out_n.t734 8.126
R6468 out_n.n66 out_n.t749 8.126
R6469 out_n.n66 out_n.t1672 8.126
R6470 out_n.n67 out_n.t1683 8.126
R6471 out_n.n67 out_n.t1112 8.126
R6472 out_n.n68 out_n.t1558 8.126
R6473 out_n.n68 out_n.t984 8.126
R6474 out_n.n69 out_n.t1275 8.126
R6475 out_n.n69 out_n.t705 8.126
R6476 out_n.n50 out_n.t544 8.126
R6477 out_n.n50 out_n.t575 8.126
R6478 out_n.n51 out_n.t771 8.126
R6479 out_n.n51 out_n.t804 8.126
R6480 out_n.n52 out_n.t1705 8.126
R6481 out_n.n52 out_n.t1735 8.126
R6482 out_n.n53 out_n.t1140 8.126
R6483 out_n.n53 out_n.t1165 8.126
R6484 out_n.n54 out_n.t1380 8.126
R6485 out_n.n54 out_n.t1409 8.126
R6486 out_n.n55 out_n.t1656 8.126
R6487 out_n.n55 out_n.t1690 8.126
R6488 out_n.n56 out_n.t1101 8.126
R6489 out_n.n56 out_n.t1132 8.126
R6490 out_n.n57 out_n.t537 8.126
R6491 out_n.n57 out_n.t569 8.126
R6492 out_n.n58 out_n.t404 8.126
R6493 out_n.n58 out_n.t438 8.126
R6494 out_n.n59 out_n.t1620 8.126
R6495 out_n.n59 out_n.t1651 8.126
R6496 out_n.n40 out_n.t1496 8.126
R6497 out_n.n40 out_n.t912 8.126
R6498 out_n.n41 out_n.t1727 8.126
R6499 out_n.n41 out_n.t1149 8.126
R6500 out_n.n42 out_n.t1158 8.126
R6501 out_n.n42 out_n.t588 8.126
R6502 out_n.n43 out_n.t593 8.126
R6503 out_n.n43 out_n.t1513 8.126
R6504 out_n.n44 out_n.t827 8.126
R6505 out_n.n44 out_n.t1754 8.126
R6506 out_n.n45 out_n.t1120 8.126
R6507 out_n.n45 out_n.t545 8.126
R6508 out_n.n46 out_n.t562 8.126
R6509 out_n.n46 out_n.t1480 8.126
R6510 out_n.n47 out_n.t1489 8.126
R6511 out_n.n47 out_n.t905 8.126
R6512 out_n.n48 out_n.t1364 8.126
R6513 out_n.n48 out_n.t784 8.126
R6514 out_n.n49 out_n.t1079 8.126
R6515 out_n.n49 out_n.t503 8.126
R6516 out_n.n30 out_n.t339 8.126
R6517 out_n.n30 out_n.t1229 8.126
R6518 out_n.n31 out_n.t581 8.126
R6519 out_n.n31 out_n.t1468 8.126
R6520 out_n.n32 out_n.t1507 8.126
R6521 out_n.n32 out_n.t891 8.126
R6522 out_n.n33 out_n.t932 8.126
R6523 out_n.n33 out_n.t327 8.126
R6524 out_n.n34 out_n.t1174 8.126
R6525 out_n.n34 out_n.t570 8.126
R6526 out_n.n35 out_n.t1466 8.126
R6527 out_n.n35 out_n.t851 8.126
R6528 out_n.n36 out_n.t894 8.126
R6529 out_n.n36 out_n.t295 8.126
R6530 out_n.n37 out_n.t331 8.126
R6531 out_n.n37 out_n.t1222 8.126
R6532 out_n.n38 out_n.t1707 8.126
R6533 out_n.n38 out_n.t1098 8.126
R6534 out_n.n39 out_n.t1429 8.126
R6535 out_n.n39 out_n.t812 8.126
R6536 out_n.n20 out_n.t652 8.126
R6537 out_n.n20 out_n.t1565 8.126
R6538 out_n.n21 out_n.t885 8.126
R6539 out_n.n21 out_n.t312 8.126
R6540 out_n.n22 out_n.t320 8.126
R6541 out_n.n22 out_n.t1246 8.126
R6542 out_n.n23 out_n.t1254 8.126
R6543 out_n.n23 out_n.t678 8.126
R6544 out_n.n24 out_n.t1491 8.126
R6545 out_n.n24 out_n.t908 8.126
R6546 out_n.n25 out_n.t277 8.126
R6547 out_n.n25 out_n.t1194 8.126
R6548 out_n.n26 out_n.t1215 8.126
R6549 out_n.n26 out_n.t637 8.126
R6550 out_n.n27 out_n.t646 8.126
R6551 out_n.n27 out_n.t1559 8.126
R6552 out_n.n28 out_n.t525 8.126
R6553 out_n.n28 out_n.t1446 8.126
R6554 out_n.n29 out_n.t1736 8.126
R6555 out_n.n29 out_n.t1157 8.126
R6556 out_n.n10 out_n.t992 8.126
R6557 out_n.n10 out_n.t415 8.126
R6558 out_n.n11 out_n.t1238 8.126
R6559 out_n.n11 out_n.t662 8.126
R6560 out_n.n12 out_n.t671 8.126
R6561 out_n.n12 out_n.t1582 8.126
R6562 out_n.n13 out_n.t1589 8.126
R6563 out_n.n13 out_n.t1017 8.126
R6564 out_n.n14 out_n.t336 8.126
R6565 out_n.n14 out_n.t1262 8.126
R6566 out_n.n15 out_n.t618 8.126
R6567 out_n.n15 out_n.t1536 8.126
R6568 out_n.n16 out_n.t1552 8.126
R6569 out_n.n16 out_n.t975 8.126
R6570 out_n.n17 out_n.t986 8.126
R6571 out_n.n17 out_n.t406 8.126
R6572 out_n.n18 out_n.t868 8.126
R6573 out_n.n18 out_n.t297 8.126
R6574 out_n.n19 out_n.t590 8.126
R6575 out_n.n19 out_n.t1509 8.126
R6576 out_n.n805 out_n.t792 8.126
R6577 out_n.n805 out_n.t1716 8.126
R6578 out_n.n806 out_n.t1028 8.126
R6579 out_n.n806 out_n.t455 8.126
R6580 out_n.n807 out_n.t463 8.126
R6581 out_n.n807 out_n.t1392 8.126
R6582 out_n.n808 out_n.t1398 8.126
R6583 out_n.n808 out_n.t817 8.126
R6584 out_n.n809 out_n.t1628 8.126
R6585 out_n.n809 out_n.t1057 8.126
R6586 out_n.n810 out_n.t417 8.126
R6587 out_n.n810 out_n.t1337 8.126
R6588 out_n.n811 out_n.t1358 8.126
R6589 out_n.n811 out_n.t776 8.126
R6590 out_n.n812 out_n.t785 8.126
R6591 out_n.n812 out_n.t1709 8.126
R6592 out_n.n813 out_n.t672 8.126
R6593 out_n.n813 out_n.t1583 8.126
R6594 out_n.n814 out_n.t375 8.126
R6595 out_n.n814 out_n.t1297 8.126
R6596 out_n.n815 out_n.t1141 8.126
R6597 out_n.n815 out_n.t1388 8.126
R6598 out_n.n816 out_n.t1383 8.126
R6599 out_n.n816 out_n.t1616 8.126
R6600 out_n.n817 out_n.t810 8.126
R6601 out_n.n817 out_n.t1052 8.126
R6602 out_n.n818 out_n.t1741 8.126
R6603 out_n.n818 out_n.t488 8.126
R6604 out_n.n819 out_n.t483 8.126
R6605 out_n.n819 out_n.t720 8.126
R6606 out_n.n820 out_n.t760 8.126
R6607 out_n.n820 out_n.t1008 8.126
R6608 out_n.n821 out_n.t1698 8.126
R6609 out_n.n821 out_n.t444 8.126
R6610 out_n.n822 out_n.t1134 8.126
R6611 out_n.n822 out_n.t1382 8.126
R6612 out_n.n823 out_n.t1011 8.126
R6613 out_n.n823 out_n.t1259 8.126
R6614 out_n.n824 out_n.t726 8.126
R6615 out_n.n824 out_n.t966 8.126
R6616 out_n.n827 out_n.t806 8.126
R6617 out_n.n827 out_n.t1729 8.126
R6618 out_n.n828 out_n.t1042 8.126
R6619 out_n.n828 out_n.t468 8.126
R6620 out_n.n829 out_n.t476 8.126
R6621 out_n.n829 out_n.t1404 8.126
R6622 out_n.n830 out_n.t1411 8.126
R6623 out_n.n830 out_n.t833 8.126
R6624 out_n.n831 out_n.t1640 8.126
R6625 out_n.n831 out_n.t1064 8.126
R6626 out_n.n832 out_n.t433 8.126
R6627 out_n.n832 out_n.t1357 8.126
R6628 out_n.n833 out_n.t1371 8.126
R6629 out_n.n833 out_n.t788 8.126
R6630 out_n.n834 out_n.t800 8.126
R6631 out_n.n834 out_n.t1721 8.126
R6632 out_n.n835 out_n.t685 8.126
R6633 out_n.n835 out_n.t1598 8.126
R6634 out_n.n836 out_n.t388 8.126
R6635 out_n.n836 out_n.t1312 8.126
R6636 out_n.n839 out_n.t1152 8.126
R6637 out_n.n839 out_n.t584 8.126
R6638 out_n.n840 out_n.t1395 8.126
R6639 out_n.n840 out_n.t813 8.126
R6640 out_n.n841 out_n.t821 8.126
R6641 out_n.n841 out_n.t1744 8.126
R6642 out_n.n842 out_n.t1757 8.126
R6643 out_n.n842 out_n.t1176 8.126
R6644 out_n.n843 out_n.t494 8.126
R6645 out_n.n843 out_n.t1420 8.126
R6646 out_n.n844 out_n.t774 8.126
R6647 out_n.n844 out_n.t1697 8.126
R6648 out_n.n845 out_n.t1713 8.126
R6649 out_n.n845 out_n.t1139 8.126
R6650 out_n.n846 out_n.t1146 8.126
R6651 out_n.n846 out_n.t577 8.126
R6652 out_n.n847 out_n.t1021 8.126
R6653 out_n.n847 out_n.t449 8.126
R6654 out_n.n848 out_n.t738 8.126
R6655 out_n.n848 out_n.t1659 8.126
R6656 out_n.n851 out_n.t609 8.126
R6657 out_n.n851 out_n.t1526 8.126
R6658 out_n.n852 out_n.t844 8.126
R6659 out_n.n852 out_n.t271 8.126
R6660 out_n.n853 out_n.t281 8.126
R6661 out_n.n853 out_n.t1200 8.126
R6662 out_n.n854 out_n.t1210 8.126
R6663 out_n.n854 out_n.t633 8.126
R6664 out_n.n855 out_n.t1451 8.126
R6665 out_n.n855 out_n.t869 8.126
R6666 out_n.n856 out_n.t1732 8.126
R6667 out_n.n856 out_n.t1153 8.126
R6668 out_n.n857 out_n.t1164 8.126
R6669 out_n.n857 out_n.t592 8.126
R6670 out_n.n858 out_n.t602 8.126
R6671 out_n.n858 out_n.t1518 8.126
R6672 out_n.n859 out_n.t480 8.126
R6673 out_n.n859 out_n.t1405 8.126
R6674 out_n.n860 out_n.t1693 8.126
R6675 out_n.n860 out_n.t1123 8.126
R6676 out_n.n863 out_n.t948 8.126
R6677 out_n.n863 out_n.t367 8.126
R6678 out_n.n864 out_n.t1188 8.126
R6679 out_n.n864 out_n.t615 8.126
R6680 out_n.n865 out_n.t620 8.126
R6681 out_n.n865 out_n.t1539 8.126
R6682 out_n.n866 out_n.t1549 8.126
R6683 out_n.n866 out_n.t970 8.126
R6684 out_n.n867 out_n.t300 8.126
R6685 out_n.n867 out_n.t1219 8.126
R6686 out_n.n868 out_n.t585 8.126
R6687 out_n.n868 out_n.t1501 8.126
R6688 out_n.n869 out_n.t1512 8.126
R6689 out_n.n869 out_n.t931 8.126
R6690 out_n.n870 out_n.t940 8.126
R6691 out_n.n870 out_n.t362 8.126
R6692 out_n.n871 out_n.t823 8.126
R6693 out_n.n871 out_n.t1747 8.126
R6694 out_n.n872 out_n.t548 8.126
R6695 out_n.n872 out_n.t1471 8.126
R6696 out_n.n875 out_n.t1290 8.126
R6697 out_n.n875 out_n.t692 8.126
R6698 out_n.n876 out_n.t1533 8.126
R6699 out_n.n876 out_n.t921 8.126
R6700 out_n.n877 out_n.t960 8.126
R6701 out_n.n877 out_n.t352 8.126
R6702 out_n.n878 out_n.t392 8.126
R6703 out_n.n878 out_n.t1283 8.126
R6704 out_n.n879 out_n.t641 8.126
R6705 out_n.n879 out_n.t1521 8.126
R6706 out_n.n880 out_n.t919 8.126
R6707 out_n.n880 out_n.t318 8.126
R6708 out_n.n881 out_n.t357 8.126
R6709 out_n.n881 out_n.t1252 8.126
R6710 out_n.n882 out_n.t1286 8.126
R6711 out_n.n882 out_n.t686 8.126
R6712 out_n.n883 out_n.t1168 8.126
R6713 out_n.n883 out_n.t568 8.126
R6714 out_n.n884 out_n.t887 8.126
R6715 out_n.n884 out_n.t282 8.126
R6716 out_n.n887 out_n.t1605 8.126
R6717 out_n.n887 out_n.t1030 8.126
R6718 out_n.n888 out_n.t344 8.126
R6719 out_n.n888 out_n.t1269 8.126
R6720 out_n.n889 out_n.t1274 8.126
R6721 out_n.n889 out_n.t704 8.126
R6722 out_n.n890 out_n.t713 8.126
R6723 out_n.n890 out_n.t1629 8.126
R6724 out_n.n891 out_n.t946 8.126
R6725 out_n.n891 out_n.t366 8.126
R6726 out_n.n892 out_n.t1243 8.126
R6727 out_n.n892 out_n.t666 8.126
R6728 out_n.n893 out_n.t677 8.126
R6729 out_n.n893 out_n.t1587 8.126
R6730 out_n.n894 out_n.t1600 8.126
R6731 out_n.n894 out_n.t1023 8.126
R6732 out_n.n895 out_n.t1488 8.126
R6733 out_n.n895 out_n.t903 8.126
R6734 out_n.n896 out_n.t1198 8.126
R6735 out_n.n896 out_n.t621 8.126
R6736 out_n.n899 out_n.t457 8.126
R6737 out_n.n899 out_n.t489 8.126
R6738 out_n.n900 out_n.t698 8.126
R6739 out_n.n900 out_n.t723 8.126
R6740 out_n.n901 out_n.t1619 8.126
R6741 out_n.n901 out_n.t1652 8.126
R6742 out_n.n902 out_n.t1058 8.126
R6743 out_n.n902 out_n.t1088 8.126
R6744 out_n.n903 out_n.t1289 8.126
R6745 out_n.n903 out_n.t1320 8.126
R6746 out_n.n904 out_n.t1576 8.126
R6747 out_n.n904 out_n.t1608 8.126
R6748 out_n.n905 out_n.t1015 8.126
R6749 out_n.n905 out_n.t1045 8.126
R6750 out_n.n906 out_n.t450 8.126
R6751 out_n.n906 out_n.t482 8.126
R6752 out_n.n907 out_n.t329 8.126
R6753 out_n.n907 out_n.t355 8.126
R6754 out_n.n908 out_n.t1540 8.126
R6755 out_n.n908 out_n.t1571 8.126
R6756 out_n.n911 out_n.t1414 8.126
R6757 out_n.n911 out_n.t834 8.126
R6758 out_n.n912 out_n.t1641 8.126
R6759 out_n.n912 out_n.t1065 8.126
R6760 out_n.n913 out_n.t1077 8.126
R6761 out_n.n913 out_n.t501 8.126
R6762 out_n.n914 out_n.t515 8.126
R6763 out_n.n914 out_n.t1438 8.126
R6764 out_n.n915 out_n.t744 8.126
R6765 out_n.n915 out_n.t1668 8.126
R6766 out_n.n916 out_n.t1033 8.126
R6767 out_n.n916 out_n.t458 8.126
R6768 out_n.n917 out_n.t471 8.126
R6769 out_n.n917 out_n.t1397 8.126
R6770 out_n.n918 out_n.t1407 8.126
R6771 out_n.n918 out_n.t824 8.126
R6772 out_n.n919 out_n.t1277 8.126
R6773 out_n.n919 out_n.t707 8.126
R6774 out_n.n920 out_n.t997 8.126
R6775 out_n.n920 out_n.t421 8.126
R6776 out_n.n923 out_n.t1758 8.126
R6777 out_n.n923 out_n.t1177 8.126
R6778 out_n.n924 out_n.t495 8.126
R6779 out_n.n924 out_n.t1421 8.126
R6780 out_n.n925 out_n.t1428 8.126
R6781 out_n.n925 out_n.t849 8.126
R6782 out_n.n926 out_n.t858 8.126
R6783 out_n.n926 out_n.t286 8.126
R6784 out_n.n927 out_n.t1097 8.126
R6785 out_n.n927 out_n.t524 8.126
R6786 out_n.n928 out_n.t1384 8.126
R6787 out_n.n928 out_n.t801 8.126
R6788 out_n.n929 out_n.t816 8.126
R6789 out_n.n929 out_n.t1740 8.126
R6790 out_n.n930 out_n.t1749 8.126
R6791 out_n.n930 out_n.t1169 8.126
R6792 out_n.n931 out_n.t1621 8.126
R6793 out_n.n931 out_n.t1048 8.126
R6794 out_n.n932 out_n.t1340 8.126
R6795 out_n.n932 out_n.t763 8.126
R6796 out_n.n935 out_n.t1211 8.126
R6797 out_n.n935 out_n.t1495 8.126
R6798 out_n.n936 out_n.t1453 8.126
R6799 out_n.n936 out_n.t1725 8.126
R6800 out_n.n937 out_n.t881 8.126
R6801 out_n.n937 out_n.t1156 8.126
R6802 out_n.n938 out_n.t315 8.126
R6803 out_n.n938 out_n.t594 8.126
R6804 out_n.n939 out_n.t557 8.126
R6805 out_n.n939 out_n.t828 8.126
R6806 out_n.n940 out_n.t837 8.126
R6807 out_n.n940 out_n.t1121 8.126
R6808 out_n.n941 out_n.t274 8.126
R6809 out_n.n941 out_n.t563 8.126
R6810 out_n.n942 out_n.t1204 8.126
R6811 out_n.n942 out_n.t1490 8.126
R6812 out_n.n943 out_n.t1082 8.126
R6813 out_n.n943 out_n.t1365 8.126
R6814 out_n.n944 out_n.t796 8.126
R6815 out_n.n944 out_n.t1078 8.126
R6816 out_n.n947 out_n.t911 8.126
R6817 out_n.n947 out_n.t338 8.126
R6818 out_n.n948 out_n.t1150 8.126
R6819 out_n.n948 out_n.t582 8.126
R6820 out_n.n949 out_n.t589 8.126
R6821 out_n.n949 out_n.t1508 8.126
R6822 out_n.n950 out_n.t1514 8.126
R6823 out_n.n950 out_n.t933 8.126
R6824 out_n.n951 out_n.t1755 8.126
R6825 out_n.n951 out_n.t1175 8.126
R6826 out_n.n952 out_n.t546 8.126
R6827 out_n.n952 out_n.t1467 8.126
R6828 out_n.n953 out_n.t1481 8.126
R6829 out_n.n953 out_n.t895 8.126
R6830 out_n.n954 out_n.t906 8.126
R6831 out_n.n954 out_n.t332 8.126
R6832 out_n.n955 out_n.t783 8.126
R6833 out_n.n955 out_n.t1708 8.126
R6834 out_n.n956 out_n.t502 8.126
R6835 out_n.n956 out_n.t1427 8.126
R6836 out_n.n0 out_n.t448 8.126
R6837 out_n.n0 out_n.t1375 8.126
R6838 out_n.n1 out_n.t690 8.126
R6839 out_n.n1 out_n.t1603 8.126
R6840 out_n.n2 out_n.t1612 8.126
R6841 out_n.n2 out_n.t1037 8.126
R6842 out_n.n3 out_n.t1046 8.126
R6843 out_n.n3 out_n.t472 8.126
R6844 out_n.n4 out_n.t1280 8.126
R6845 out_n.n4 out_n.t710 8.126
R6846 out_n.n5 out_n.t1567 8.126
R6847 out_n.n5 out_n.t993 8.126
R6848 out_n.n6 out_n.t1009 8.126
R6849 out_n.n6 out_n.t434 8.126
R6850 out_n.n7 out_n.t440 8.126
R6851 out_n.n7 out_n.t1367 8.126
R6852 out_n.n8 out_n.t321 8.126
R6853 out_n.n8 out_n.t1247 8.126
R6854 out_n.n9 out_n.t1532 8.126
R6855 out_n.n9 out_n.t955 8.126
R6856 out_n.n957 out_n.t195 4.95
R6857 out_n.n957 out_n.t57 4.95
R6858 out_n.n958 out_n.t203 4.95
R6859 out_n.n958 out_n.t256 4.95
R6860 out_n.n945 out_n.t229 4.95
R6861 out_n.n945 out_n.t207 4.95
R6862 out_n.n946 out_n.t74 4.95
R6863 out_n.n946 out_n.t118 4.95
R6864 out_n.n933 out_n.t83 4.95
R6865 out_n.n933 out_n.t92 4.95
R6866 out_n.n934 out_n.t23 4.95
R6867 out_n.n934 out_n.t163 4.95
R6868 out_n.n921 out_n.t143 4.95
R6869 out_n.n921 out_n.t249 4.95
R6870 out_n.n922 out_n.t172 4.95
R6871 out_n.n922 out_n.t211 4.95
R6872 out_n.n909 out_n.t30 4.95
R6873 out_n.n909 out_n.t61 4.95
R6874 out_n.n910 out_n.t183 4.95
R6875 out_n.n910 out_n.t97 4.95
R6876 out_n.n897 out_n.t244 4.95
R6877 out_n.n897 out_n.t124 4.95
R6878 out_n.n898 out_n.t1792 4.95
R6879 out_n.n898 out_n.t107 4.95
R6880 out_n.n885 out_n.t218 4.95
R6881 out_n.n885 out_n.t4 4.95
R6882 out_n.n886 out_n.t155 4.95
R6883 out_n.n886 out_n.t70 4.95
R6884 out_n.n873 out_n.t190 4.95
R6885 out_n.n873 out_n.t257 4.95
R6886 out_n.n874 out_n.t214 4.95
R6887 out_n.n874 out_n.t1777 4.95
R6888 out_n.n861 out_n.t147 4.95
R6889 out_n.n861 out_n.t77 4.95
R6890 out_n.n862 out_n.t131 4.95
R6891 out_n.n862 out_n.t261 4.95
R6892 out_n.n849 out_n.t137 4.95
R6893 out_n.n849 out_n.t114 4.95
R6894 out_n.n850 out_n.t232 4.95
R6895 out_n.n850 out_n.t29 4.95
R6896 out_n.n837 out_n.t151 4.95
R6897 out_n.n837 out_n.t88 4.95
R6898 out_n.n838 out_n.t46 4.95
R6899 out_n.n838 out_n.t9 4.95
R6900 out_n.n825 out_n.t174 4.95
R6901 out_n.n825 out_n.t1798 4.95
R6902 out_n.n826 out_n.t90 4.95
R6903 out_n.n826 out_n.t39 4.95
R6904 out_n.n803 out_n.t164 4.95
R6905 out_n.n803 out_n.t1764 4.95
R6906 out_n.n804 out_n.t48 4.95
R6907 out_n.n804 out_n.t12 4.95
R6908 out_n.n800 out_n.t215 4.95
R6909 out_n.n800 out_n.t1778 4.95
R6910 out_n.n801 out_n.t123 4.95
R6911 out_n.n801 out_n.t65 4.95
R6912 out_n.n797 out_n.t133 4.95
R6913 out_n.n797 out_n.t50 4.95
R6914 out_n.n798 out_n.t3 4.95
R6915 out_n.n798 out_n.t243 4.95
R6916 out_n.n794 out_n.t58 4.95
R6917 out_n.n794 out_n.t162 4.95
R6918 out_n.n795 out_n.t255 4.95
R6919 out_n.n795 out_n.t222 4.95
R6920 out_n.n791 out_n.t206 4.95
R6921 out_n.n791 out_n.t196 4.95
R6922 out_n.n792 out_n.t117 4.95
R6923 out_n.n792 out_n.t202 4.95
R6924 out_n.n788 out_n.t95 4.95
R6925 out_n.n788 out_n.t1783 4.95
R6926 out_n.n789 out_n.t112 4.95
R6927 out_n.n789 out_n.t144 4.95
R6928 out_n.n785 out_n.t1768 4.95
R6929 out_n.n785 out_n.t178 4.95
R6930 out_n.n786 out_n.t86 4.95
R6931 out_n.n786 out_n.t136 4.95
R6932 out_n.n782 out_n.t240 4.95
R6933 out_n.n782 out_n.t168 4.95
R6934 out_n.n783 out_n.t1797 4.95
R6935 out_n.n783 out_n.t150 4.95
R6936 out_n.n779 out_n.t223 4.95
R6937 out_n.n779 out_n.t234 4.95
R6938 out_n.n780 out_n.t106 4.95
R6939 out_n.n780 out_n.t14 4.95
R6940 out_n.n776 out_n.t5 4.95
R6941 out_n.n776 out_n.t245 4.95
R6942 out_n.n777 out_n.t69 4.95
R6943 out_n.n777 out_n.t1791 4.95
R6944 out_n.n773 out_n.t76 4.95
R6945 out_n.n773 out_n.t72 4.95
R6946 out_n.n774 out_n.t220 4.95
R6947 out_n.n774 out_n.t236 4.95
R6948 out_n.n770 out_n.t208 4.95
R6949 out_n.n770 out_n.t18 4.95
R6950 out_n.n771 out_n.t192 4.95
R6951 out_n.n771 out_n.t54 4.95
R6952 out_n.n767 out_n.t1787 4.95
R6953 out_n.n767 out_n.t43 4.95
R6954 out_n.n768 out_n.t111 4.95
R6955 out_n.n768 out_n.t79 4.95
R6956 out_n.n764 out_n.t87 4.95
R6957 out_n.n764 out_n.t181 4.95
R6958 out_n.n765 out_n.t8 4.95
R6959 out_n.n765 out_n.t1785 4.95
R6960 out_n.n761 out_n.t1799 4.95
R6961 out_n.n761 out_n.t152 4.95
R6962 out_n.n762 out_n.t38 4.95
R6963 out_n.n762 out_n.t45 4.95
R6964 out_n.n758 out_n.t35 4.95
R6965 out_n.n758 out_n.t238 4.95
R6966 out_n.n759 out_n.t63 4.95
R6967 out_n.n759 out_n.t128 4.95
R6968 out_n.n755 out_n.t259 4.95
R6969 out_n.n755 out_n.t227 4.95
R6970 out_n.n756 out_n.t1795 4.95
R6971 out_n.n756 out_n.t121 4.95
R6972 out_n.n752 out_n.t25 4.95
R6973 out_n.n752 out_n.t1774 4.95
R6974 out_n.n753 out_n.t1772 4.95
R6975 out_n.n753 out_n.t1 4.95
R6976 out_n.n749 out_n.t193 4.95
R6977 out_n.n749 out_n.t230 4.95
R6978 out_n.n750 out_n.t200 4.95
R6979 out_n.n750 out_n.t75 4.95
R6980 out_n.n746 out_n.t113 4.95
R6981 out_n.n746 out_n.t80 4.95
R6982 out_n.n747 out_n.t27 4.95
R6983 out_n.n747 out_n.t52 4.95
R6984 out_n.n743 out_n.t176 4.95
R6985 out_n.n743 out_n.t1786 4.95
R6986 out_n.n744 out_n.t93 4.95
R6987 out_n.n744 out_n.t148 4.95
R6988 out_n.n740 out_n.t166 4.95
R6989 out_n.n740 out_n.t1766 4.95
R6990 out_n.n741 out_n.t250 4.95
R6991 out_n.n741 out_n.t84 4.95
R6992 out_n.n737 out_n.t64 4.95
R6993 out_n.n737 out_n.t16 4.95
R6994 out_n.n738 out_n.t180 4.95
R6995 out_n.n738 out_n.t127 4.95
R6996 out_n.n734 out_n.t169 4.95
R6997 out_n.n734 out_n.t122 4.95
R6998 out_n.n735 out_n.t251 4.95
R6999 out_n.n735 out_n.t104 4.95
R7000 out_n.n731 out_n.t235 4.95
R7001 out_n.n731 out_n.t241 4.95
R7002 out_n.n732 out_n.t13 4.95
R7003 out_n.n732 out_n.t1796 4.95
R7004 out_n.n728 out_n.t201 4.95
R7005 out_n.n728 out_n.t253 4.95
R7006 out_n.n729 out_n.t226 4.95
R7007 out_n.n729 out_n.t34 4.95
R7008 out_n.n725 out_n.t28 4.95
R7009 out_n.n725 out_n.t116 4.95
R7010 out_n.n726 out_n.t1773 4.95
R7011 out_n.n726 out_n.t258 4.95
R7012 out_n.n722 out_n.t135 4.95
R7013 out_n.n722 out_n.t149 4.95
R7014 out_n.n723 out_n.t228 4.95
R7015 out_n.n723 out_n.t134 4.95
R7016 out_n.n719 out_n.t42 4.95
R7017 out_n.n719 out_n.t85 4.95
R7018 out_n.n720 out_n.t78 4.95
R7019 out_n.n720 out_n.t6 4.95
R7020 out_n.n716 out_n.t182 4.95
R7021 out_n.n716 out_n.t94 4.95
R7022 out_n.n717 out_n.t1784 4.95
R7023 out_n.n717 out_n.t110 4.95
R7024 out_n.n713 out_n.t1790 4.95
R7025 out_n.n713 out_n.t105 4.95
R7026 out_n.n714 out_n.t1765 4.95
R7027 out_n.n714 out_n.t175 4.95
R7028 out_n.n710 out_n.t233 4.95
R7029 out_n.n710 out_n.t68 4.95
R7030 out_n.n711 out_n.t188 4.95
R7031 out_n.n711 out_n.t165 4.95
R7032 out_n.n707 out_n.t53 4.95
R7033 out_n.n707 out_n.t219 4.95
R7034 out_n.n708 out_n.t1779 4.95
R7035 out_n.n708 out_n.t156 4.95
R7036 out_n.n704 out_n.t1775 4.95
R7037 out_n.n704 out_n.t191 4.95
R7038 out_n.n705 out_n.t0 4.95
R7039 out_n.n705 out_n.t216 4.95
R7040 out_n.n701 out_n.t231 4.95
R7041 out_n.n701 out_n.t26 4.95
R7042 out_n.n702 out_n.t73 4.95
R7043 out_n.n702 out_n.t1771 4.95
R7044 out_n.n698 out_n.t44 4.95
R7045 out_n.n698 out_n.t7 4.95
R7046 out_n.n699 out_n.t197 4.95
R7047 out_n.n699 out_n.t59 4.95
R7048 out_n.n695 out_n.t125 4.95
R7049 out_n.n695 out_n.t37 4.95
R7050 out_n.n696 out_n.t171 4.95
R7051 out_n.n696 out_n.t40 4.95
R7052 out_n.n692 out_n.t120 4.95
R7053 out_n.n692 out_n.t62 4.95
R7054 out_n.n693 out_n.t101 4.95
R7055 out_n.n693 out_n.t98 4.95
R7056 out_n.n689 out_n.t15 4.95
R7057 out_n.n689 out_n.t1794 4.95
R7058 out_n.n690 out_n.t126 4.95
R7059 out_n.n690 out_n.t1769 4.95
R7060 out_n.n686 out_n.t1781 4.95
R7061 out_n.n686 out_n.t158 4.95
R7062 out_n.n687 out_n.t32 4.95
R7063 out_n.n687 out_n.t186 4.95
R7064 out_n.n683 out_n.t51 4.95
R7065 out_n.n683 out_n.t199 4.95
R7066 out_n.n684 out_n.t246 4.95
R7067 out_n.n684 out_n.t225 4.95
R7068 out_n.n680 out_n.t146 4.95
R7069 out_n.n680 out_n.t24 4.95
R7070 out_n.n681 out_n.t130 4.95
R7071 out_n.n681 out_n.t1770 4.95
R7072 out_n.n677 out_n.t82 4.95
R7073 out_n.n677 out_n.t91 4.95
R7074 out_n.n678 out_n.t21 4.95
R7075 out_n.n678 out_n.t160 4.95
R7076 out_n.n674 out_n.t36 4.95
R7077 out_n.n674 out_n.t248 4.95
R7078 out_n.n675 out_n.t205 4.95
R7079 out_n.n675 out_n.t210 4.95
R7080 out_n.n671 out_n.t103 4.95
R7081 out_n.n671 out_n.t179 4.95
R7082 out_n.n672 out_n.t139 4.95
R7083 out_n.n672 out_n.t1782 4.95
R7084 out_n.n668 out_n.t67 4.95
R7085 out_n.n668 out_n.t1789 4.95
R7086 out_n.n669 out_n.t154 4.95
R7087 out_n.n669 out_n.t1763 4.95
R7088 out_n.n665 out_n.t247 4.95
R7089 out_n.n665 out_n.t81 4.95
R7090 out_n.n666 out_n.t209 4.95
R7091 out_n.n666 out_n.t20 4.95
R7092 out_n.n662 out_n.t60 4.95
R7093 out_n.n662 out_n.t142 4.95
R7094 out_n.n663 out_n.t96 4.95
R7095 out_n.n663 out_n.t170 4.95
R7096 out_n.n659 out_n.t1788 4.95
R7097 out_n.n659 out_n.t109 4.95
R7098 out_n.n660 out_n.t1762 4.95
R7099 out_n.n660 out_n.t100 4.95
R7100 out_n.n656 out_n.t157 4.95
R7101 out_n.n656 out_n.t66 4.95
R7102 out_n.n657 out_n.t185 4.95
R7103 out_n.n657 out_n.t153 4.95
R7104 out_n.n653 out_n.t217 4.95
R7105 out_n.n653 out_n.t1780 4.95
R7106 out_n.n654 out_n.t224 4.95
R7107 out_n.n654 out_n.t31 4.95
R7108 out_n.n650 out_n.t119 4.95
R7109 out_n.n650 out_n.t189 4.95
R7110 out_n.n651 out_n.t260 4.95
R7111 out_n.n651 out_n.t213 4.95
R7112 out_n.n647 out_n.t89 4.95
R7113 out_n.n647 out_n.t145 4.95
R7114 out_n.n648 out_n.t159 4.95
R7115 out_n.n648 out_n.t129 4.95
R7116 out_n.n644 out_n.t212 4.95
R7117 out_n.n644 out_n.t11 4.95
R7118 out_n.n645 out_n.t194 4.95
R7119 out_n.n645 out_n.t19 4.95
R7120 out_n.n641 out_n.t99 4.95
R7121 out_n.n641 out_n.t173 4.95
R7122 out_n.n642 out_n.t115 4.95
R7123 out_n.n642 out_n.t204 4.95
R7124 out_n.n638 out_n.t108 4.95
R7125 out_n.n638 out_n.t102 4.95
R7126 out_n.n639 out_n.t177 4.95
R7127 out_n.n639 out_n.t138 4.95
R7128 out_n.n635 out_n.t71 4.95
R7129 out_n.n635 out_n.t1793 4.95
R7130 out_n.n636 out_n.t167 4.95
R7131 out_n.n636 out_n.t1767 4.95
R7132 out_n.n632 out_n.t254 4.95
R7133 out_n.n632 out_n.t237 4.95
R7134 out_n.n633 out_n.t1776 4.95
R7135 out_n.n633 out_n.t239 4.95
R7136 out_n.n629 out_n.t49 4.95
R7137 out_n.n629 out_n.t55 4.95
R7138 out_n.n630 out_n.t242 4.95
R7139 out_n.n630 out_n.t252 4.95
R7140 out_n.n626 out_n.t161 4.95
R7141 out_n.n626 out_n.t132 4.95
R7142 out_n.n627 out_n.t221 4.95
R7143 out_n.n627 out_n.t2 4.95
R7144 out_n.n623 out_n.t10 4.95
R7145 out_n.n623 out_n.t22 4.95
R7146 out_n.n624 out_n.t17 4.95
R7147 out_n.n624 out_n.t56 4.95
R7148 out_n.n620 out_n.t140 4.95
R7149 out_n.n620 out_n.t47 4.95
R7150 out_n.n621 out_n.t41 4.95
R7151 out_n.n621 out_n.t198 4.95
R7152 out_n.n971 out_n.t33 4.95
R7153 out_n.n971 out_n.t187 4.95
R7154 out_n.n972 out_n.t184 4.95
R7155 out_n.n972 out_n.t141 4.95
R7156 out_n.n615 out_n.n614 0.866
R7157 out_n.n605 out_n.n604 0.849
R7158 out_n.n595 out_n.n594 0.849
R7159 out_n.n585 out_n.n584 0.849
R7160 out_n.n575 out_n.n574 0.849
R7161 out_n.n565 out_n.n564 0.849
R7162 out_n.n555 out_n.n554 0.849
R7163 out_n.n545 out_n.n544 0.849
R7164 out_n.n535 out_n.n534 0.849
R7165 out_n.n525 out_n.n524 0.849
R7166 out_n.n515 out_n.n514 0.849
R7167 out_n.n505 out_n.n504 0.849
R7168 out_n.n495 out_n.n494 0.849
R7169 out_n.n485 out_n.n484 0.849
R7170 out_n.n475 out_n.n474 0.849
R7171 out_n.n465 out_n.n464 0.849
R7172 out_n.n455 out_n.n454 0.849
R7173 out_n.n445 out_n.n444 0.849
R7174 out_n.n435 out_n.n434 0.849
R7175 out_n.n425 out_n.n424 0.849
R7176 out_n.n415 out_n.n414 0.849
R7177 out_n.n405 out_n.n404 0.849
R7178 out_n.n395 out_n.n394 0.849
R7179 out_n.n385 out_n.n384 0.849
R7180 out_n.n375 out_n.n374 0.849
R7181 out_n.n365 out_n.n364 0.849
R7182 out_n.n355 out_n.n354 0.849
R7183 out_n.n345 out_n.n344 0.849
R7184 out_n.n335 out_n.n334 0.849
R7185 out_n.n325 out_n.n324 0.849
R7186 out_n.n315 out_n.n314 0.849
R7187 out_n.n305 out_n.n304 0.849
R7188 out_n.n295 out_n.n294 0.849
R7189 out_n.n285 out_n.n284 0.849
R7190 out_n.n275 out_n.n274 0.849
R7191 out_n.n265 out_n.n264 0.849
R7192 out_n.n255 out_n.n254 0.849
R7193 out_n.n245 out_n.n244 0.849
R7194 out_n.n235 out_n.n234 0.849
R7195 out_n.n225 out_n.n224 0.849
R7196 out_n.n215 out_n.n214 0.849
R7197 out_n.n205 out_n.n204 0.849
R7198 out_n.n195 out_n.n194 0.849
R7199 out_n.n185 out_n.n184 0.849
R7200 out_n.n175 out_n.n174 0.849
R7201 out_n.n165 out_n.n164 0.849
R7202 out_n.n155 out_n.n154 0.849
R7203 out_n.n145 out_n.n144 0.849
R7204 out_n.n135 out_n.n134 0.849
R7205 out_n.n125 out_n.n124 0.849
R7206 out_n.n115 out_n.n114 0.849
R7207 out_n.n105 out_n.n104 0.849
R7208 out_n.n95 out_n.n94 0.849
R7209 out_n.n85 out_n.n84 0.849
R7210 out_n.n75 out_n.n74 0.849
R7211 out_n.n65 out_n.n64 0.849
R7212 out_n.n55 out_n.n54 0.849
R7213 out_n.n45 out_n.n44 0.849
R7214 out_n.n35 out_n.n34 0.849
R7215 out_n.n25 out_n.n24 0.849
R7216 out_n.n15 out_n.n14 0.849
R7217 out_n.n810 out_n.n809 0.849
R7218 out_n.n820 out_n.n819 0.849
R7219 out_n.n832 out_n.n831 0.849
R7220 out_n.n844 out_n.n843 0.849
R7221 out_n.n856 out_n.n855 0.849
R7222 out_n.n868 out_n.n867 0.849
R7223 out_n.n880 out_n.n879 0.849
R7224 out_n.n892 out_n.n891 0.849
R7225 out_n.n904 out_n.n903 0.849
R7226 out_n.n916 out_n.n915 0.849
R7227 out_n.n928 out_n.n927 0.849
R7228 out_n.n940 out_n.n939 0.849
R7229 out_n.n952 out_n.n951 0.849
R7230 out_n.n5 out_n.n4 0.849
R7231 out_n.n611 out_n.n610 0.77
R7232 out_n.n612 out_n.n611 0.77
R7233 out_n.n613 out_n.n612 0.77
R7234 out_n.n614 out_n.n613 0.77
R7235 out_n.n616 out_n.n615 0.77
R7236 out_n.n617 out_n.n616 0.77
R7237 out_n.n618 out_n.n617 0.77
R7238 out_n.n619 out_n.n618 0.77
R7239 out_n.n958 out_n.n957 0.76
R7240 out_n.n946 out_n.n945 0.76
R7241 out_n.n934 out_n.n933 0.76
R7242 out_n.n922 out_n.n921 0.76
R7243 out_n.n910 out_n.n909 0.76
R7244 out_n.n898 out_n.n897 0.76
R7245 out_n.n886 out_n.n885 0.76
R7246 out_n.n874 out_n.n873 0.76
R7247 out_n.n862 out_n.n861 0.76
R7248 out_n.n850 out_n.n849 0.76
R7249 out_n.n838 out_n.n837 0.76
R7250 out_n.n826 out_n.n825 0.76
R7251 out_n.n804 out_n.n803 0.76
R7252 out_n.n801 out_n.n800 0.76
R7253 out_n.n798 out_n.n797 0.76
R7254 out_n.n795 out_n.n794 0.76
R7255 out_n.n792 out_n.n791 0.76
R7256 out_n.n789 out_n.n788 0.76
R7257 out_n.n786 out_n.n785 0.76
R7258 out_n.n783 out_n.n782 0.76
R7259 out_n.n780 out_n.n779 0.76
R7260 out_n.n777 out_n.n776 0.76
R7261 out_n.n774 out_n.n773 0.76
R7262 out_n.n771 out_n.n770 0.76
R7263 out_n.n768 out_n.n767 0.76
R7264 out_n.n765 out_n.n764 0.76
R7265 out_n.n762 out_n.n761 0.76
R7266 out_n.n759 out_n.n758 0.76
R7267 out_n.n756 out_n.n755 0.76
R7268 out_n.n753 out_n.n752 0.76
R7269 out_n.n750 out_n.n749 0.76
R7270 out_n.n747 out_n.n746 0.76
R7271 out_n.n744 out_n.n743 0.76
R7272 out_n.n741 out_n.n740 0.76
R7273 out_n.n738 out_n.n737 0.76
R7274 out_n.n735 out_n.n734 0.76
R7275 out_n.n732 out_n.n731 0.76
R7276 out_n.n729 out_n.n728 0.76
R7277 out_n.n726 out_n.n725 0.76
R7278 out_n.n723 out_n.n722 0.76
R7279 out_n.n720 out_n.n719 0.76
R7280 out_n.n717 out_n.n716 0.76
R7281 out_n.n714 out_n.n713 0.76
R7282 out_n.n711 out_n.n710 0.76
R7283 out_n.n708 out_n.n707 0.76
R7284 out_n.n705 out_n.n704 0.76
R7285 out_n.n702 out_n.n701 0.76
R7286 out_n.n699 out_n.n698 0.76
R7287 out_n.n696 out_n.n695 0.76
R7288 out_n.n693 out_n.n692 0.76
R7289 out_n.n690 out_n.n689 0.76
R7290 out_n.n687 out_n.n686 0.76
R7291 out_n.n684 out_n.n683 0.76
R7292 out_n.n681 out_n.n680 0.76
R7293 out_n.n678 out_n.n677 0.76
R7294 out_n.n675 out_n.n674 0.76
R7295 out_n.n672 out_n.n671 0.76
R7296 out_n.n669 out_n.n668 0.76
R7297 out_n.n666 out_n.n665 0.76
R7298 out_n.n663 out_n.n662 0.76
R7299 out_n.n660 out_n.n659 0.76
R7300 out_n.n657 out_n.n656 0.76
R7301 out_n.n654 out_n.n653 0.76
R7302 out_n.n651 out_n.n650 0.76
R7303 out_n.n648 out_n.n647 0.76
R7304 out_n.n645 out_n.n644 0.76
R7305 out_n.n642 out_n.n641 0.76
R7306 out_n.n639 out_n.n638 0.76
R7307 out_n.n636 out_n.n635 0.76
R7308 out_n.n633 out_n.n632 0.76
R7309 out_n.n630 out_n.n629 0.76
R7310 out_n.n627 out_n.n626 0.76
R7311 out_n.n624 out_n.n623 0.76
R7312 out_n.n621 out_n.n620 0.76
R7313 out_n.n972 out_n.n971 0.76
R7314 out_n.n601 out_n.n600 0.753
R7315 out_n.n602 out_n.n601 0.753
R7316 out_n.n603 out_n.n602 0.753
R7317 out_n.n604 out_n.n603 0.753
R7318 out_n.n606 out_n.n605 0.753
R7319 out_n.n607 out_n.n606 0.753
R7320 out_n.n608 out_n.n607 0.753
R7321 out_n.n609 out_n.n608 0.753
R7322 out_n.n591 out_n.n590 0.753
R7323 out_n.n592 out_n.n591 0.753
R7324 out_n.n593 out_n.n592 0.753
R7325 out_n.n594 out_n.n593 0.753
R7326 out_n.n596 out_n.n595 0.753
R7327 out_n.n597 out_n.n596 0.753
R7328 out_n.n598 out_n.n597 0.753
R7329 out_n.n599 out_n.n598 0.753
R7330 out_n.n581 out_n.n580 0.753
R7331 out_n.n582 out_n.n581 0.753
R7332 out_n.n583 out_n.n582 0.753
R7333 out_n.n584 out_n.n583 0.753
R7334 out_n.n586 out_n.n585 0.753
R7335 out_n.n587 out_n.n586 0.753
R7336 out_n.n588 out_n.n587 0.753
R7337 out_n.n589 out_n.n588 0.753
R7338 out_n.n571 out_n.n570 0.753
R7339 out_n.n572 out_n.n571 0.753
R7340 out_n.n573 out_n.n572 0.753
R7341 out_n.n574 out_n.n573 0.753
R7342 out_n.n576 out_n.n575 0.753
R7343 out_n.n577 out_n.n576 0.753
R7344 out_n.n578 out_n.n577 0.753
R7345 out_n.n579 out_n.n578 0.753
R7346 out_n.n561 out_n.n560 0.753
R7347 out_n.n562 out_n.n561 0.753
R7348 out_n.n563 out_n.n562 0.753
R7349 out_n.n564 out_n.n563 0.753
R7350 out_n.n566 out_n.n565 0.753
R7351 out_n.n567 out_n.n566 0.753
R7352 out_n.n568 out_n.n567 0.753
R7353 out_n.n569 out_n.n568 0.753
R7354 out_n.n551 out_n.n550 0.753
R7355 out_n.n552 out_n.n551 0.753
R7356 out_n.n553 out_n.n552 0.753
R7357 out_n.n554 out_n.n553 0.753
R7358 out_n.n556 out_n.n555 0.753
R7359 out_n.n557 out_n.n556 0.753
R7360 out_n.n558 out_n.n557 0.753
R7361 out_n.n559 out_n.n558 0.753
R7362 out_n.n541 out_n.n540 0.753
R7363 out_n.n542 out_n.n541 0.753
R7364 out_n.n543 out_n.n542 0.753
R7365 out_n.n544 out_n.n543 0.753
R7366 out_n.n546 out_n.n545 0.753
R7367 out_n.n547 out_n.n546 0.753
R7368 out_n.n548 out_n.n547 0.753
R7369 out_n.n549 out_n.n548 0.753
R7370 out_n.n531 out_n.n530 0.753
R7371 out_n.n532 out_n.n531 0.753
R7372 out_n.n533 out_n.n532 0.753
R7373 out_n.n534 out_n.n533 0.753
R7374 out_n.n536 out_n.n535 0.753
R7375 out_n.n537 out_n.n536 0.753
R7376 out_n.n538 out_n.n537 0.753
R7377 out_n.n539 out_n.n538 0.753
R7378 out_n.n521 out_n.n520 0.753
R7379 out_n.n522 out_n.n521 0.753
R7380 out_n.n523 out_n.n522 0.753
R7381 out_n.n524 out_n.n523 0.753
R7382 out_n.n526 out_n.n525 0.753
R7383 out_n.n527 out_n.n526 0.753
R7384 out_n.n528 out_n.n527 0.753
R7385 out_n.n529 out_n.n528 0.753
R7386 out_n.n511 out_n.n510 0.753
R7387 out_n.n512 out_n.n511 0.753
R7388 out_n.n513 out_n.n512 0.753
R7389 out_n.n514 out_n.n513 0.753
R7390 out_n.n516 out_n.n515 0.753
R7391 out_n.n517 out_n.n516 0.753
R7392 out_n.n518 out_n.n517 0.753
R7393 out_n.n519 out_n.n518 0.753
R7394 out_n.n501 out_n.n500 0.753
R7395 out_n.n502 out_n.n501 0.753
R7396 out_n.n503 out_n.n502 0.753
R7397 out_n.n504 out_n.n503 0.753
R7398 out_n.n506 out_n.n505 0.753
R7399 out_n.n507 out_n.n506 0.753
R7400 out_n.n508 out_n.n507 0.753
R7401 out_n.n509 out_n.n508 0.753
R7402 out_n.n491 out_n.n490 0.753
R7403 out_n.n492 out_n.n491 0.753
R7404 out_n.n493 out_n.n492 0.753
R7405 out_n.n494 out_n.n493 0.753
R7406 out_n.n496 out_n.n495 0.753
R7407 out_n.n497 out_n.n496 0.753
R7408 out_n.n498 out_n.n497 0.753
R7409 out_n.n499 out_n.n498 0.753
R7410 out_n.n481 out_n.n480 0.753
R7411 out_n.n482 out_n.n481 0.753
R7412 out_n.n483 out_n.n482 0.753
R7413 out_n.n484 out_n.n483 0.753
R7414 out_n.n486 out_n.n485 0.753
R7415 out_n.n487 out_n.n486 0.753
R7416 out_n.n488 out_n.n487 0.753
R7417 out_n.n489 out_n.n488 0.753
R7418 out_n.n471 out_n.n470 0.753
R7419 out_n.n472 out_n.n471 0.753
R7420 out_n.n473 out_n.n472 0.753
R7421 out_n.n474 out_n.n473 0.753
R7422 out_n.n476 out_n.n475 0.753
R7423 out_n.n477 out_n.n476 0.753
R7424 out_n.n478 out_n.n477 0.753
R7425 out_n.n479 out_n.n478 0.753
R7426 out_n.n461 out_n.n460 0.753
R7427 out_n.n462 out_n.n461 0.753
R7428 out_n.n463 out_n.n462 0.753
R7429 out_n.n464 out_n.n463 0.753
R7430 out_n.n466 out_n.n465 0.753
R7431 out_n.n467 out_n.n466 0.753
R7432 out_n.n468 out_n.n467 0.753
R7433 out_n.n469 out_n.n468 0.753
R7434 out_n.n451 out_n.n450 0.753
R7435 out_n.n452 out_n.n451 0.753
R7436 out_n.n453 out_n.n452 0.753
R7437 out_n.n454 out_n.n453 0.753
R7438 out_n.n456 out_n.n455 0.753
R7439 out_n.n457 out_n.n456 0.753
R7440 out_n.n458 out_n.n457 0.753
R7441 out_n.n459 out_n.n458 0.753
R7442 out_n.n441 out_n.n440 0.753
R7443 out_n.n442 out_n.n441 0.753
R7444 out_n.n443 out_n.n442 0.753
R7445 out_n.n444 out_n.n443 0.753
R7446 out_n.n446 out_n.n445 0.753
R7447 out_n.n447 out_n.n446 0.753
R7448 out_n.n448 out_n.n447 0.753
R7449 out_n.n449 out_n.n448 0.753
R7450 out_n.n431 out_n.n430 0.753
R7451 out_n.n432 out_n.n431 0.753
R7452 out_n.n433 out_n.n432 0.753
R7453 out_n.n434 out_n.n433 0.753
R7454 out_n.n436 out_n.n435 0.753
R7455 out_n.n437 out_n.n436 0.753
R7456 out_n.n438 out_n.n437 0.753
R7457 out_n.n439 out_n.n438 0.753
R7458 out_n.n421 out_n.n420 0.753
R7459 out_n.n422 out_n.n421 0.753
R7460 out_n.n423 out_n.n422 0.753
R7461 out_n.n424 out_n.n423 0.753
R7462 out_n.n426 out_n.n425 0.753
R7463 out_n.n427 out_n.n426 0.753
R7464 out_n.n428 out_n.n427 0.753
R7465 out_n.n429 out_n.n428 0.753
R7466 out_n.n411 out_n.n410 0.753
R7467 out_n.n412 out_n.n411 0.753
R7468 out_n.n413 out_n.n412 0.753
R7469 out_n.n414 out_n.n413 0.753
R7470 out_n.n416 out_n.n415 0.753
R7471 out_n.n417 out_n.n416 0.753
R7472 out_n.n418 out_n.n417 0.753
R7473 out_n.n419 out_n.n418 0.753
R7474 out_n.n401 out_n.n400 0.753
R7475 out_n.n402 out_n.n401 0.753
R7476 out_n.n403 out_n.n402 0.753
R7477 out_n.n404 out_n.n403 0.753
R7478 out_n.n406 out_n.n405 0.753
R7479 out_n.n407 out_n.n406 0.753
R7480 out_n.n408 out_n.n407 0.753
R7481 out_n.n409 out_n.n408 0.753
R7482 out_n.n391 out_n.n390 0.753
R7483 out_n.n392 out_n.n391 0.753
R7484 out_n.n393 out_n.n392 0.753
R7485 out_n.n394 out_n.n393 0.753
R7486 out_n.n396 out_n.n395 0.753
R7487 out_n.n397 out_n.n396 0.753
R7488 out_n.n398 out_n.n397 0.753
R7489 out_n.n399 out_n.n398 0.753
R7490 out_n.n381 out_n.n380 0.753
R7491 out_n.n382 out_n.n381 0.753
R7492 out_n.n383 out_n.n382 0.753
R7493 out_n.n384 out_n.n383 0.753
R7494 out_n.n386 out_n.n385 0.753
R7495 out_n.n387 out_n.n386 0.753
R7496 out_n.n388 out_n.n387 0.753
R7497 out_n.n389 out_n.n388 0.753
R7498 out_n.n371 out_n.n370 0.753
R7499 out_n.n372 out_n.n371 0.753
R7500 out_n.n373 out_n.n372 0.753
R7501 out_n.n374 out_n.n373 0.753
R7502 out_n.n376 out_n.n375 0.753
R7503 out_n.n377 out_n.n376 0.753
R7504 out_n.n378 out_n.n377 0.753
R7505 out_n.n379 out_n.n378 0.753
R7506 out_n.n361 out_n.n360 0.753
R7507 out_n.n362 out_n.n361 0.753
R7508 out_n.n363 out_n.n362 0.753
R7509 out_n.n364 out_n.n363 0.753
R7510 out_n.n366 out_n.n365 0.753
R7511 out_n.n367 out_n.n366 0.753
R7512 out_n.n368 out_n.n367 0.753
R7513 out_n.n369 out_n.n368 0.753
R7514 out_n.n351 out_n.n350 0.753
R7515 out_n.n352 out_n.n351 0.753
R7516 out_n.n353 out_n.n352 0.753
R7517 out_n.n354 out_n.n353 0.753
R7518 out_n.n356 out_n.n355 0.753
R7519 out_n.n357 out_n.n356 0.753
R7520 out_n.n358 out_n.n357 0.753
R7521 out_n.n359 out_n.n358 0.753
R7522 out_n.n341 out_n.n340 0.753
R7523 out_n.n342 out_n.n341 0.753
R7524 out_n.n343 out_n.n342 0.753
R7525 out_n.n344 out_n.n343 0.753
R7526 out_n.n346 out_n.n345 0.753
R7527 out_n.n347 out_n.n346 0.753
R7528 out_n.n348 out_n.n347 0.753
R7529 out_n.n349 out_n.n348 0.753
R7530 out_n.n331 out_n.n330 0.753
R7531 out_n.n332 out_n.n331 0.753
R7532 out_n.n333 out_n.n332 0.753
R7533 out_n.n334 out_n.n333 0.753
R7534 out_n.n336 out_n.n335 0.753
R7535 out_n.n337 out_n.n336 0.753
R7536 out_n.n338 out_n.n337 0.753
R7537 out_n.n339 out_n.n338 0.753
R7538 out_n.n321 out_n.n320 0.753
R7539 out_n.n322 out_n.n321 0.753
R7540 out_n.n323 out_n.n322 0.753
R7541 out_n.n324 out_n.n323 0.753
R7542 out_n.n326 out_n.n325 0.753
R7543 out_n.n327 out_n.n326 0.753
R7544 out_n.n328 out_n.n327 0.753
R7545 out_n.n329 out_n.n328 0.753
R7546 out_n.n311 out_n.n310 0.753
R7547 out_n.n312 out_n.n311 0.753
R7548 out_n.n313 out_n.n312 0.753
R7549 out_n.n314 out_n.n313 0.753
R7550 out_n.n316 out_n.n315 0.753
R7551 out_n.n317 out_n.n316 0.753
R7552 out_n.n318 out_n.n317 0.753
R7553 out_n.n319 out_n.n318 0.753
R7554 out_n.n301 out_n.n300 0.753
R7555 out_n.n302 out_n.n301 0.753
R7556 out_n.n303 out_n.n302 0.753
R7557 out_n.n304 out_n.n303 0.753
R7558 out_n.n306 out_n.n305 0.753
R7559 out_n.n307 out_n.n306 0.753
R7560 out_n.n308 out_n.n307 0.753
R7561 out_n.n309 out_n.n308 0.753
R7562 out_n.n291 out_n.n290 0.753
R7563 out_n.n292 out_n.n291 0.753
R7564 out_n.n293 out_n.n292 0.753
R7565 out_n.n294 out_n.n293 0.753
R7566 out_n.n296 out_n.n295 0.753
R7567 out_n.n297 out_n.n296 0.753
R7568 out_n.n298 out_n.n297 0.753
R7569 out_n.n299 out_n.n298 0.753
R7570 out_n.n281 out_n.n280 0.753
R7571 out_n.n282 out_n.n281 0.753
R7572 out_n.n283 out_n.n282 0.753
R7573 out_n.n284 out_n.n283 0.753
R7574 out_n.n286 out_n.n285 0.753
R7575 out_n.n287 out_n.n286 0.753
R7576 out_n.n288 out_n.n287 0.753
R7577 out_n.n289 out_n.n288 0.753
R7578 out_n.n271 out_n.n270 0.753
R7579 out_n.n272 out_n.n271 0.753
R7580 out_n.n273 out_n.n272 0.753
R7581 out_n.n274 out_n.n273 0.753
R7582 out_n.n276 out_n.n275 0.753
R7583 out_n.n277 out_n.n276 0.753
R7584 out_n.n278 out_n.n277 0.753
R7585 out_n.n279 out_n.n278 0.753
R7586 out_n.n261 out_n.n260 0.753
R7587 out_n.n262 out_n.n261 0.753
R7588 out_n.n263 out_n.n262 0.753
R7589 out_n.n264 out_n.n263 0.753
R7590 out_n.n266 out_n.n265 0.753
R7591 out_n.n267 out_n.n266 0.753
R7592 out_n.n268 out_n.n267 0.753
R7593 out_n.n269 out_n.n268 0.753
R7594 out_n.n251 out_n.n250 0.753
R7595 out_n.n252 out_n.n251 0.753
R7596 out_n.n253 out_n.n252 0.753
R7597 out_n.n254 out_n.n253 0.753
R7598 out_n.n256 out_n.n255 0.753
R7599 out_n.n257 out_n.n256 0.753
R7600 out_n.n258 out_n.n257 0.753
R7601 out_n.n259 out_n.n258 0.753
R7602 out_n.n241 out_n.n240 0.753
R7603 out_n.n242 out_n.n241 0.753
R7604 out_n.n243 out_n.n242 0.753
R7605 out_n.n244 out_n.n243 0.753
R7606 out_n.n246 out_n.n245 0.753
R7607 out_n.n247 out_n.n246 0.753
R7608 out_n.n248 out_n.n247 0.753
R7609 out_n.n249 out_n.n248 0.753
R7610 out_n.n231 out_n.n230 0.753
R7611 out_n.n232 out_n.n231 0.753
R7612 out_n.n233 out_n.n232 0.753
R7613 out_n.n234 out_n.n233 0.753
R7614 out_n.n236 out_n.n235 0.753
R7615 out_n.n237 out_n.n236 0.753
R7616 out_n.n238 out_n.n237 0.753
R7617 out_n.n239 out_n.n238 0.753
R7618 out_n.n221 out_n.n220 0.753
R7619 out_n.n222 out_n.n221 0.753
R7620 out_n.n223 out_n.n222 0.753
R7621 out_n.n224 out_n.n223 0.753
R7622 out_n.n226 out_n.n225 0.753
R7623 out_n.n227 out_n.n226 0.753
R7624 out_n.n228 out_n.n227 0.753
R7625 out_n.n229 out_n.n228 0.753
R7626 out_n.n211 out_n.n210 0.753
R7627 out_n.n212 out_n.n211 0.753
R7628 out_n.n213 out_n.n212 0.753
R7629 out_n.n214 out_n.n213 0.753
R7630 out_n.n216 out_n.n215 0.753
R7631 out_n.n217 out_n.n216 0.753
R7632 out_n.n218 out_n.n217 0.753
R7633 out_n.n219 out_n.n218 0.753
R7634 out_n.n201 out_n.n200 0.753
R7635 out_n.n202 out_n.n201 0.753
R7636 out_n.n203 out_n.n202 0.753
R7637 out_n.n204 out_n.n203 0.753
R7638 out_n.n206 out_n.n205 0.753
R7639 out_n.n207 out_n.n206 0.753
R7640 out_n.n208 out_n.n207 0.753
R7641 out_n.n209 out_n.n208 0.753
R7642 out_n.n191 out_n.n190 0.753
R7643 out_n.n192 out_n.n191 0.753
R7644 out_n.n193 out_n.n192 0.753
R7645 out_n.n194 out_n.n193 0.753
R7646 out_n.n196 out_n.n195 0.753
R7647 out_n.n197 out_n.n196 0.753
R7648 out_n.n198 out_n.n197 0.753
R7649 out_n.n199 out_n.n198 0.753
R7650 out_n.n181 out_n.n180 0.753
R7651 out_n.n182 out_n.n181 0.753
R7652 out_n.n183 out_n.n182 0.753
R7653 out_n.n184 out_n.n183 0.753
R7654 out_n.n186 out_n.n185 0.753
R7655 out_n.n187 out_n.n186 0.753
R7656 out_n.n188 out_n.n187 0.753
R7657 out_n.n189 out_n.n188 0.753
R7658 out_n.n171 out_n.n170 0.753
R7659 out_n.n172 out_n.n171 0.753
R7660 out_n.n173 out_n.n172 0.753
R7661 out_n.n174 out_n.n173 0.753
R7662 out_n.n176 out_n.n175 0.753
R7663 out_n.n177 out_n.n176 0.753
R7664 out_n.n178 out_n.n177 0.753
R7665 out_n.n179 out_n.n178 0.753
R7666 out_n.n161 out_n.n160 0.753
R7667 out_n.n162 out_n.n161 0.753
R7668 out_n.n163 out_n.n162 0.753
R7669 out_n.n164 out_n.n163 0.753
R7670 out_n.n166 out_n.n165 0.753
R7671 out_n.n167 out_n.n166 0.753
R7672 out_n.n168 out_n.n167 0.753
R7673 out_n.n169 out_n.n168 0.753
R7674 out_n.n151 out_n.n150 0.753
R7675 out_n.n152 out_n.n151 0.753
R7676 out_n.n153 out_n.n152 0.753
R7677 out_n.n154 out_n.n153 0.753
R7678 out_n.n156 out_n.n155 0.753
R7679 out_n.n157 out_n.n156 0.753
R7680 out_n.n158 out_n.n157 0.753
R7681 out_n.n159 out_n.n158 0.753
R7682 out_n.n141 out_n.n140 0.753
R7683 out_n.n142 out_n.n141 0.753
R7684 out_n.n143 out_n.n142 0.753
R7685 out_n.n144 out_n.n143 0.753
R7686 out_n.n146 out_n.n145 0.753
R7687 out_n.n147 out_n.n146 0.753
R7688 out_n.n148 out_n.n147 0.753
R7689 out_n.n149 out_n.n148 0.753
R7690 out_n.n131 out_n.n130 0.753
R7691 out_n.n132 out_n.n131 0.753
R7692 out_n.n133 out_n.n132 0.753
R7693 out_n.n134 out_n.n133 0.753
R7694 out_n.n136 out_n.n135 0.753
R7695 out_n.n137 out_n.n136 0.753
R7696 out_n.n138 out_n.n137 0.753
R7697 out_n.n139 out_n.n138 0.753
R7698 out_n.n121 out_n.n120 0.753
R7699 out_n.n122 out_n.n121 0.753
R7700 out_n.n123 out_n.n122 0.753
R7701 out_n.n124 out_n.n123 0.753
R7702 out_n.n126 out_n.n125 0.753
R7703 out_n.n127 out_n.n126 0.753
R7704 out_n.n128 out_n.n127 0.753
R7705 out_n.n129 out_n.n128 0.753
R7706 out_n.n111 out_n.n110 0.753
R7707 out_n.n112 out_n.n111 0.753
R7708 out_n.n113 out_n.n112 0.753
R7709 out_n.n114 out_n.n113 0.753
R7710 out_n.n116 out_n.n115 0.753
R7711 out_n.n117 out_n.n116 0.753
R7712 out_n.n118 out_n.n117 0.753
R7713 out_n.n119 out_n.n118 0.753
R7714 out_n.n101 out_n.n100 0.753
R7715 out_n.n102 out_n.n101 0.753
R7716 out_n.n103 out_n.n102 0.753
R7717 out_n.n104 out_n.n103 0.753
R7718 out_n.n106 out_n.n105 0.753
R7719 out_n.n107 out_n.n106 0.753
R7720 out_n.n108 out_n.n107 0.753
R7721 out_n.n109 out_n.n108 0.753
R7722 out_n.n91 out_n.n90 0.753
R7723 out_n.n92 out_n.n91 0.753
R7724 out_n.n93 out_n.n92 0.753
R7725 out_n.n94 out_n.n93 0.753
R7726 out_n.n96 out_n.n95 0.753
R7727 out_n.n97 out_n.n96 0.753
R7728 out_n.n98 out_n.n97 0.753
R7729 out_n.n99 out_n.n98 0.753
R7730 out_n.n81 out_n.n80 0.753
R7731 out_n.n82 out_n.n81 0.753
R7732 out_n.n83 out_n.n82 0.753
R7733 out_n.n84 out_n.n83 0.753
R7734 out_n.n86 out_n.n85 0.753
R7735 out_n.n87 out_n.n86 0.753
R7736 out_n.n88 out_n.n87 0.753
R7737 out_n.n89 out_n.n88 0.753
R7738 out_n.n71 out_n.n70 0.753
R7739 out_n.n72 out_n.n71 0.753
R7740 out_n.n73 out_n.n72 0.753
R7741 out_n.n74 out_n.n73 0.753
R7742 out_n.n76 out_n.n75 0.753
R7743 out_n.n77 out_n.n76 0.753
R7744 out_n.n78 out_n.n77 0.753
R7745 out_n.n79 out_n.n78 0.753
R7746 out_n.n61 out_n.n60 0.753
R7747 out_n.n62 out_n.n61 0.753
R7748 out_n.n63 out_n.n62 0.753
R7749 out_n.n64 out_n.n63 0.753
R7750 out_n.n66 out_n.n65 0.753
R7751 out_n.n67 out_n.n66 0.753
R7752 out_n.n68 out_n.n67 0.753
R7753 out_n.n69 out_n.n68 0.753
R7754 out_n.n51 out_n.n50 0.753
R7755 out_n.n52 out_n.n51 0.753
R7756 out_n.n53 out_n.n52 0.753
R7757 out_n.n54 out_n.n53 0.753
R7758 out_n.n56 out_n.n55 0.753
R7759 out_n.n57 out_n.n56 0.753
R7760 out_n.n58 out_n.n57 0.753
R7761 out_n.n59 out_n.n58 0.753
R7762 out_n.n41 out_n.n40 0.753
R7763 out_n.n42 out_n.n41 0.753
R7764 out_n.n43 out_n.n42 0.753
R7765 out_n.n44 out_n.n43 0.753
R7766 out_n.n46 out_n.n45 0.753
R7767 out_n.n47 out_n.n46 0.753
R7768 out_n.n48 out_n.n47 0.753
R7769 out_n.n49 out_n.n48 0.753
R7770 out_n.n31 out_n.n30 0.753
R7771 out_n.n32 out_n.n31 0.753
R7772 out_n.n33 out_n.n32 0.753
R7773 out_n.n34 out_n.n33 0.753
R7774 out_n.n36 out_n.n35 0.753
R7775 out_n.n37 out_n.n36 0.753
R7776 out_n.n38 out_n.n37 0.753
R7777 out_n.n39 out_n.n38 0.753
R7778 out_n.n21 out_n.n20 0.753
R7779 out_n.n22 out_n.n21 0.753
R7780 out_n.n23 out_n.n22 0.753
R7781 out_n.n24 out_n.n23 0.753
R7782 out_n.n26 out_n.n25 0.753
R7783 out_n.n27 out_n.n26 0.753
R7784 out_n.n28 out_n.n27 0.753
R7785 out_n.n29 out_n.n28 0.753
R7786 out_n.n11 out_n.n10 0.753
R7787 out_n.n12 out_n.n11 0.753
R7788 out_n.n13 out_n.n12 0.753
R7789 out_n.n14 out_n.n13 0.753
R7790 out_n.n16 out_n.n15 0.753
R7791 out_n.n17 out_n.n16 0.753
R7792 out_n.n18 out_n.n17 0.753
R7793 out_n.n19 out_n.n18 0.753
R7794 out_n.n806 out_n.n805 0.753
R7795 out_n.n807 out_n.n806 0.753
R7796 out_n.n808 out_n.n807 0.753
R7797 out_n.n809 out_n.n808 0.753
R7798 out_n.n811 out_n.n810 0.753
R7799 out_n.n812 out_n.n811 0.753
R7800 out_n.n813 out_n.n812 0.753
R7801 out_n.n814 out_n.n813 0.753
R7802 out_n.n816 out_n.n815 0.753
R7803 out_n.n817 out_n.n816 0.753
R7804 out_n.n818 out_n.n817 0.753
R7805 out_n.n819 out_n.n818 0.753
R7806 out_n.n821 out_n.n820 0.753
R7807 out_n.n822 out_n.n821 0.753
R7808 out_n.n823 out_n.n822 0.753
R7809 out_n.n824 out_n.n823 0.753
R7810 out_n.n828 out_n.n827 0.753
R7811 out_n.n829 out_n.n828 0.753
R7812 out_n.n830 out_n.n829 0.753
R7813 out_n.n831 out_n.n830 0.753
R7814 out_n.n833 out_n.n832 0.753
R7815 out_n.n834 out_n.n833 0.753
R7816 out_n.n835 out_n.n834 0.753
R7817 out_n.n836 out_n.n835 0.753
R7818 out_n.n840 out_n.n839 0.753
R7819 out_n.n841 out_n.n840 0.753
R7820 out_n.n842 out_n.n841 0.753
R7821 out_n.n843 out_n.n842 0.753
R7822 out_n.n845 out_n.n844 0.753
R7823 out_n.n846 out_n.n845 0.753
R7824 out_n.n847 out_n.n846 0.753
R7825 out_n.n848 out_n.n847 0.753
R7826 out_n.n852 out_n.n851 0.753
R7827 out_n.n853 out_n.n852 0.753
R7828 out_n.n854 out_n.n853 0.753
R7829 out_n.n855 out_n.n854 0.753
R7830 out_n.n857 out_n.n856 0.753
R7831 out_n.n858 out_n.n857 0.753
R7832 out_n.n859 out_n.n858 0.753
R7833 out_n.n860 out_n.n859 0.753
R7834 out_n.n864 out_n.n863 0.753
R7835 out_n.n865 out_n.n864 0.753
R7836 out_n.n866 out_n.n865 0.753
R7837 out_n.n867 out_n.n866 0.753
R7838 out_n.n869 out_n.n868 0.753
R7839 out_n.n870 out_n.n869 0.753
R7840 out_n.n871 out_n.n870 0.753
R7841 out_n.n872 out_n.n871 0.753
R7842 out_n.n876 out_n.n875 0.753
R7843 out_n.n877 out_n.n876 0.753
R7844 out_n.n878 out_n.n877 0.753
R7845 out_n.n879 out_n.n878 0.753
R7846 out_n.n881 out_n.n880 0.753
R7847 out_n.n882 out_n.n881 0.753
R7848 out_n.n883 out_n.n882 0.753
R7849 out_n.n884 out_n.n883 0.753
R7850 out_n.n888 out_n.n887 0.753
R7851 out_n.n889 out_n.n888 0.753
R7852 out_n.n890 out_n.n889 0.753
R7853 out_n.n891 out_n.n890 0.753
R7854 out_n.n893 out_n.n892 0.753
R7855 out_n.n894 out_n.n893 0.753
R7856 out_n.n895 out_n.n894 0.753
R7857 out_n.n896 out_n.n895 0.753
R7858 out_n.n900 out_n.n899 0.753
R7859 out_n.n901 out_n.n900 0.753
R7860 out_n.n902 out_n.n901 0.753
R7861 out_n.n903 out_n.n902 0.753
R7862 out_n.n905 out_n.n904 0.753
R7863 out_n.n906 out_n.n905 0.753
R7864 out_n.n907 out_n.n906 0.753
R7865 out_n.n908 out_n.n907 0.753
R7866 out_n.n912 out_n.n911 0.753
R7867 out_n.n913 out_n.n912 0.753
R7868 out_n.n914 out_n.n913 0.753
R7869 out_n.n915 out_n.n914 0.753
R7870 out_n.n917 out_n.n916 0.753
R7871 out_n.n918 out_n.n917 0.753
R7872 out_n.n919 out_n.n918 0.753
R7873 out_n.n920 out_n.n919 0.753
R7874 out_n.n924 out_n.n923 0.753
R7875 out_n.n925 out_n.n924 0.753
R7876 out_n.n926 out_n.n925 0.753
R7877 out_n.n927 out_n.n926 0.753
R7878 out_n.n929 out_n.n928 0.753
R7879 out_n.n930 out_n.n929 0.753
R7880 out_n.n931 out_n.n930 0.753
R7881 out_n.n932 out_n.n931 0.753
R7882 out_n.n936 out_n.n935 0.753
R7883 out_n.n937 out_n.n936 0.753
R7884 out_n.n938 out_n.n937 0.753
R7885 out_n.n939 out_n.n938 0.753
R7886 out_n.n941 out_n.n940 0.753
R7887 out_n.n942 out_n.n941 0.753
R7888 out_n.n943 out_n.n942 0.753
R7889 out_n.n944 out_n.n943 0.753
R7890 out_n.n948 out_n.n947 0.753
R7891 out_n.n949 out_n.n948 0.753
R7892 out_n.n950 out_n.n949 0.753
R7893 out_n.n951 out_n.n950 0.753
R7894 out_n.n953 out_n.n952 0.753
R7895 out_n.n954 out_n.n953 0.753
R7896 out_n.n955 out_n.n954 0.753
R7897 out_n.n956 out_n.n955 0.753
R7898 out_n.n1 out_n.n0 0.753
R7899 out_n.n2 out_n.n1 0.753
R7900 out_n.n3 out_n.n2 0.753
R7901 out_n.n4 out_n.n3 0.753
R7902 out_n.n6 out_n.n5 0.753
R7903 out_n.n7 out_n.n6 0.753
R7904 out_n.n8 out_n.n7 0.753
R7905 out_n.n9 out_n.n8 0.753
R7906 out_n.n959 out_n.n958 0.554
R7907 out_n.n960 out_n.n946 0.554
R7908 out_n.n961 out_n.n934 0.554
R7909 out_n.n962 out_n.n922 0.554
R7910 out_n.n963 out_n.n910 0.554
R7911 out_n.n964 out_n.n898 0.554
R7912 out_n.n965 out_n.n886 0.554
R7913 out_n.n966 out_n.n874 0.554
R7914 out_n.n967 out_n.n862 0.554
R7915 out_n.n968 out_n.n850 0.554
R7916 out_n.n969 out_n.n838 0.554
R7917 out_n.n970 out_n.n826 0.554
R7918 out_n out_n.n804 0.554
R7919 out_n.n802 out_n.n801 0.554
R7920 out_n.n799 out_n.n798 0.554
R7921 out_n.n796 out_n.n795 0.554
R7922 out_n.n793 out_n.n792 0.554
R7923 out_n.n790 out_n.n789 0.554
R7924 out_n.n787 out_n.n786 0.554
R7925 out_n.n784 out_n.n783 0.554
R7926 out_n.n781 out_n.n780 0.554
R7927 out_n.n778 out_n.n777 0.554
R7928 out_n.n775 out_n.n774 0.554
R7929 out_n.n772 out_n.n771 0.554
R7930 out_n.n769 out_n.n768 0.554
R7931 out_n.n766 out_n.n765 0.554
R7932 out_n.n763 out_n.n762 0.554
R7933 out_n.n760 out_n.n759 0.554
R7934 out_n.n757 out_n.n756 0.554
R7935 out_n.n754 out_n.n753 0.554
R7936 out_n.n751 out_n.n750 0.554
R7937 out_n.n748 out_n.n747 0.554
R7938 out_n.n745 out_n.n744 0.554
R7939 out_n.n742 out_n.n741 0.554
R7940 out_n.n739 out_n.n738 0.554
R7941 out_n.n736 out_n.n735 0.554
R7942 out_n.n733 out_n.n732 0.554
R7943 out_n.n730 out_n.n729 0.554
R7944 out_n.n727 out_n.n726 0.554
R7945 out_n.n724 out_n.n723 0.554
R7946 out_n.n721 out_n.n720 0.554
R7947 out_n.n718 out_n.n717 0.554
R7948 out_n.n715 out_n.n714 0.554
R7949 out_n.n712 out_n.n711 0.554
R7950 out_n.n709 out_n.n708 0.554
R7951 out_n.n706 out_n.n705 0.554
R7952 out_n.n703 out_n.n702 0.554
R7953 out_n.n700 out_n.n699 0.554
R7954 out_n.n697 out_n.n696 0.554
R7955 out_n.n694 out_n.n693 0.554
R7956 out_n.n691 out_n.n690 0.554
R7957 out_n.n688 out_n.n687 0.554
R7958 out_n.n685 out_n.n684 0.554
R7959 out_n.n682 out_n.n681 0.554
R7960 out_n.n679 out_n.n678 0.554
R7961 out_n.n676 out_n.n675 0.554
R7962 out_n.n673 out_n.n672 0.554
R7963 out_n.n670 out_n.n669 0.554
R7964 out_n.n667 out_n.n666 0.554
R7965 out_n.n664 out_n.n663 0.554
R7966 out_n.n661 out_n.n660 0.554
R7967 out_n.n658 out_n.n657 0.554
R7968 out_n.n655 out_n.n654 0.554
R7969 out_n.n652 out_n.n651 0.554
R7970 out_n.n649 out_n.n648 0.554
R7971 out_n.n646 out_n.n645 0.554
R7972 out_n.n643 out_n.n642 0.554
R7973 out_n.n640 out_n.n639 0.554
R7974 out_n.n637 out_n.n636 0.554
R7975 out_n.n634 out_n.n633 0.554
R7976 out_n.n631 out_n.n630 0.554
R7977 out_n.n628 out_n.n627 0.554
R7978 out_n.n625 out_n.n624 0.554
R7979 out_n.n622 out_n.n621 0.554
R7980 out_n.n973 out_n.n972 0.554
R7981 out_n.n622 out_n.n619 0.541
R7982 out_n.n625 out_n.n609 0.523
R7983 out_n.n628 out_n.n599 0.523
R7984 out_n.n631 out_n.n589 0.523
R7985 out_n.n634 out_n.n579 0.523
R7986 out_n.n637 out_n.n569 0.523
R7987 out_n.n640 out_n.n559 0.523
R7988 out_n.n643 out_n.n549 0.523
R7989 out_n.n646 out_n.n539 0.523
R7990 out_n.n649 out_n.n529 0.523
R7991 out_n.n652 out_n.n519 0.523
R7992 out_n.n655 out_n.n509 0.523
R7993 out_n.n658 out_n.n499 0.523
R7994 out_n.n661 out_n.n489 0.523
R7995 out_n.n664 out_n.n479 0.523
R7996 out_n.n667 out_n.n469 0.523
R7997 out_n.n670 out_n.n459 0.523
R7998 out_n.n673 out_n.n449 0.523
R7999 out_n.n676 out_n.n439 0.523
R8000 out_n.n679 out_n.n429 0.523
R8001 out_n.n682 out_n.n419 0.523
R8002 out_n.n685 out_n.n409 0.523
R8003 out_n.n688 out_n.n399 0.523
R8004 out_n.n691 out_n.n389 0.523
R8005 out_n.n694 out_n.n379 0.523
R8006 out_n.n697 out_n.n369 0.523
R8007 out_n.n700 out_n.n359 0.523
R8008 out_n.n703 out_n.n349 0.523
R8009 out_n.n706 out_n.n339 0.523
R8010 out_n.n709 out_n.n329 0.523
R8011 out_n.n712 out_n.n319 0.523
R8012 out_n.n715 out_n.n309 0.523
R8013 out_n.n718 out_n.n299 0.523
R8014 out_n.n721 out_n.n289 0.523
R8015 out_n.n724 out_n.n279 0.523
R8016 out_n.n727 out_n.n269 0.523
R8017 out_n.n730 out_n.n259 0.523
R8018 out_n.n733 out_n.n249 0.523
R8019 out_n.n736 out_n.n239 0.523
R8020 out_n.n739 out_n.n229 0.523
R8021 out_n.n742 out_n.n219 0.523
R8022 out_n.n745 out_n.n209 0.523
R8023 out_n.n748 out_n.n199 0.523
R8024 out_n.n751 out_n.n189 0.523
R8025 out_n.n754 out_n.n179 0.523
R8026 out_n.n757 out_n.n169 0.523
R8027 out_n.n760 out_n.n159 0.523
R8028 out_n.n763 out_n.n149 0.523
R8029 out_n.n766 out_n.n139 0.523
R8030 out_n.n769 out_n.n129 0.523
R8031 out_n.n772 out_n.n119 0.523
R8032 out_n.n775 out_n.n109 0.523
R8033 out_n.n778 out_n.n99 0.523
R8034 out_n.n781 out_n.n89 0.523
R8035 out_n.n784 out_n.n79 0.523
R8036 out_n.n787 out_n.n69 0.523
R8037 out_n.n790 out_n.n59 0.523
R8038 out_n.n793 out_n.n49 0.523
R8039 out_n.n796 out_n.n39 0.523
R8040 out_n.n799 out_n.n29 0.523
R8041 out_n.n802 out_n.n19 0.523
R8042 out_n out_n.n814 0.523
R8043 out_n.n970 out_n.n824 0.523
R8044 out_n.n969 out_n.n836 0.523
R8045 out_n.n968 out_n.n848 0.523
R8046 out_n.n967 out_n.n860 0.523
R8047 out_n.n966 out_n.n872 0.523
R8048 out_n.n965 out_n.n884 0.523
R8049 out_n.n964 out_n.n896 0.523
R8050 out_n.n963 out_n.n908 0.523
R8051 out_n.n962 out_n.n920 0.523
R8052 out_n.n961 out_n.n932 0.523
R8053 out_n.n960 out_n.n944 0.523
R8054 out_n.n959 out_n.n956 0.523
R8055 out_n.n973 out_n.n9 0.523
R8056 out_n.n960 out_n.n959 0.002
R8057 out_n.n961 out_n.n960 0.002
R8058 out_n.n962 out_n.n961 0.002
R8059 out_n.n963 out_n.n962 0.002
R8060 out_n.n964 out_n.n963 0.002
R8061 out_n.n965 out_n.n964 0.002
R8062 out_n.n966 out_n.n965 0.002
R8063 out_n.n967 out_n.n966 0.002
R8064 out_n.n968 out_n.n967 0.002
R8065 out_n.n969 out_n.n968 0.002
R8066 out_n.n970 out_n.n969 0.002
R8067 out_n out_n.n970 0.002
R8068 out_n.n973 out_n 0.002
R8069 out_n.n973 out_n.n802 0.002
R8070 out_n.n802 out_n.n799 0.002
R8071 out_n.n799 out_n.n796 0.002
R8072 out_n.n796 out_n.n793 0.002
R8073 out_n.n793 out_n.n790 0.002
R8074 out_n.n790 out_n.n787 0.002
R8075 out_n.n787 out_n.n784 0.002
R8076 out_n.n784 out_n.n781 0.002
R8077 out_n.n781 out_n.n778 0.002
R8078 out_n.n778 out_n.n775 0.002
R8079 out_n.n775 out_n.n772 0.002
R8080 out_n.n772 out_n.n769 0.002
R8081 out_n.n769 out_n.n766 0.002
R8082 out_n.n766 out_n.n763 0.002
R8083 out_n.n763 out_n.n760 0.002
R8084 out_n.n760 out_n.n757 0.002
R8085 out_n.n757 out_n.n754 0.002
R8086 out_n.n754 out_n.n751 0.002
R8087 out_n.n751 out_n.n748 0.002
R8088 out_n.n748 out_n.n745 0.002
R8089 out_n.n745 out_n.n742 0.002
R8090 out_n.n742 out_n.n739 0.002
R8091 out_n.n739 out_n.n736 0.002
R8092 out_n.n736 out_n.n733 0.002
R8093 out_n.n733 out_n.n730 0.002
R8094 out_n.n730 out_n.n727 0.002
R8095 out_n.n727 out_n.n724 0.002
R8096 out_n.n724 out_n.n721 0.002
R8097 out_n.n721 out_n.n718 0.002
R8098 out_n.n718 out_n.n715 0.002
R8099 out_n.n715 out_n.n712 0.002
R8100 out_n.n712 out_n.n709 0.002
R8101 out_n.n709 out_n.n706 0.002
R8102 out_n.n706 out_n.n703 0.002
R8103 out_n.n703 out_n.n700 0.002
R8104 out_n.n700 out_n.n697 0.002
R8105 out_n.n697 out_n.n694 0.002
R8106 out_n.n694 out_n.n691 0.002
R8107 out_n.n691 out_n.n688 0.002
R8108 out_n.n688 out_n.n685 0.002
R8109 out_n.n685 out_n.n682 0.002
R8110 out_n.n682 out_n.n679 0.002
R8111 out_n.n679 out_n.n676 0.002
R8112 out_n.n676 out_n.n673 0.002
R8113 out_n.n673 out_n.n670 0.002
R8114 out_n.n670 out_n.n667 0.002
R8115 out_n.n667 out_n.n664 0.002
R8116 out_n.n664 out_n.n661 0.002
R8117 out_n.n661 out_n.n658 0.002
R8118 out_n.n658 out_n.n655 0.002
R8119 out_n.n655 out_n.n652 0.002
R8120 out_n.n652 out_n.n649 0.002
R8121 out_n.n649 out_n.n646 0.002
R8122 out_n.n646 out_n.n643 0.002
R8123 out_n.n643 out_n.n640 0.002
R8124 out_n.n640 out_n.n637 0.002
R8125 out_n.n637 out_n.n634 0.002
R8126 out_n.n634 out_n.n631 0.002
R8127 out_n.n631 out_n.n628 0.002
R8128 out_n.n628 out_n.n625 0.002
R8129 out_n.n625 out_n.n622 0.002
R8130 vp_p.n668 vp_p.t1390 756.008
R8131 vp_p.n668 vp_p.t466 756.008
R8132 vp_p.n666 vp_p.t124 756.008
R8133 vp_p.n666 vp_p.t707 756.008
R8134 vp_p.n664 vp_p.t1219 756.008
R8135 vp_p.n664 vp_p.t290 756.008
R8136 vp_p.n662 vp_p.t650 756.008
R8137 vp_p.n662 vp_p.t1209 756.008
R8138 vp_p.n660 vp_p.t879 756.008
R8139 vp_p.n660 vp_p.t1443 756.008
R8140 vp_p.n658 vp_p.t475 756.008
R8141 vp_p.n658 vp_p.t1039 756.008
R8142 vp_p.n656 vp_p.t713 756.008
R8143 vp_p.n656 vp_p.t1273 756.008
R8144 vp_p.n654 vp_p.t299 756.008
R8145 vp_p.n654 vp_p.t866 756.008
R8146 vp_p.n652 vp_p.t362 756.008
R8147 vp_p.n652 vp_p.t930 756.008
R8148 vp_p.n650 vp_p.t1451 756.008
R8149 vp_p.n650 vp_p.t531 756.008
R8150 vp_p.n648 vp_p.t1052 756.008
R8151 vp_p.n648 vp_p.t112 756.008
R8152 vp_p.n646 vp_p.t1277 756.008
R8153 vp_p.n646 vp_p.t356 756.008
R8154 vp_p.n644 vp_p.t876 756.008
R8155 vp_p.n644 vp_p.t1435 756.008
R8156 vp_p.n642 vp_p.t933 756.008
R8157 vp_p.n642 vp_p.t1499 756.008
R8158 vp_p.n640 vp_p.t536 756.008
R8159 vp_p.n640 vp_p.t1105 756.008
R8160 vp_p.n638 vp_p.t120 756.008
R8161 vp_p.n638 vp_p.t699 756.008
R8162 vp_p.n636 vp_p.t142 756.008
R8163 vp_p.n636 vp_p.t718 756.008
R8164 vp_p.n634 vp_p.t1228 756.008
R8165 vp_p.n634 vp_p.t303 756.008
R8166 vp_p.n632 vp_p.t1300 756.008
R8167 vp_p.n632 vp_p.t372 756.008
R8168 vp_p.n630 vp_p.t898 756.008
R8169 vp_p.n630 vp_p.t1458 756.008
R8170 vp_p.n628 vp_p.t1132 756.008
R8171 vp_p.n628 vp_p.t192 756.008
R8172 vp_p.n626 vp_p.t726 756.008
R8173 vp_p.n626 vp_p.t1281 756.008
R8174 vp_p.n624 vp_p.t308 756.008
R8175 vp_p.n624 vp_p.t882 756.008
R8176 vp_p.n622 vp_p.t387 756.008
R8177 vp_p.n622 vp_p.t943 756.008
R8178 vp_p.n620 vp_p.t1466 756.008
R8179 vp_p.n620 vp_p.t542 756.008
R8180 vp_p.n618 vp_p.t205 756.008
R8181 vp_p.n618 vp_p.t778 756.008
R8182 vp_p.n616 vp_p.t1291 756.008
R8183 vp_p.n616 vp_p.t366 756.008
R8184 vp_p.n614 vp_p.t888 756.008
R8185 vp_p.n614 vp_p.t1453 756.008
R8186 vp_p.n612 vp_p.t956 756.008
R8187 vp_p.n612 vp_p.t14 756.008
R8188 vp_p.n610 vp_p.t551 756.008
R8189 vp_p.n610 vp_p.t1113 756.008
R8190 vp_p.n608 vp_p.t790 756.008
R8191 vp_p.n608 vp_p.t1343 756.008
R8192 vp_p.n606 vp_p.t378 756.008
R8193 vp_p.n606 vp_p.t936 756.008
R8194 vp_p.n604 vp_p.t614 756.008
R8195 vp_p.n604 vp_p.t1173 756.008
R8196 vp_p.n602 vp_p.t25 756.008
R8197 vp_p.n602 vp_p.t600 756.008
R8198 vp_p.n600 vp_p.t1123 756.008
R8199 vp_p.n600 vp_p.t183 756.008
R8200 vp_p.n598 vp_p.t1356 756.008
R8201 vp_p.n598 vp_p.t428 756.008
R8202 vp_p.n596 vp_p.t947 756.008
R8203 vp_p.n596 vp_p.t4 756.008
R8204 vp_p.n594 vp_p.t1188 756.008
R8205 vp_p.n594 vp_p.t249 756.008
R8206 vp_p.n592 vp_p.t615 756.008
R8207 vp_p.n592 vp_p.t1176 756.008
R8208 vp_p.n590 vp_p.t238 756.008
R8209 vp_p.n590 vp_p.t809 756.008
R8210 vp_p.n588 vp_p.t1330 756.008
R8211 vp_p.n588 vp_p.t401 756.008
R8212 vp_p.n586 vp_p.t918 756.008
R8213 vp_p.n586 vp_p.t1476 756.008
R8214 vp_p.n584 vp_p.t1153 756.008
R8215 vp_p.n584 vp_p.t217 756.008
R8216 vp_p.n582 vp_p.t581 756.008
R8217 vp_p.n582 vp_p.t1141 756.008
R8218 vp_p.n580 vp_p.t819 756.008
R8219 vp_p.n580 vp_p.t1377 756.008
R8220 vp_p.n578 vp_p.t411 756.008
R8221 vp_p.n578 vp_p.t967 756.008
R8222 vp_p.n576 vp_p.t1483 756.008
R8223 vp_p.n576 vp_p.t562 756.008
R8224 vp_p.n574 vp_p.t231 756.008
R8225 vp_p.n574 vp_p.t802 756.008
R8226 vp_p.n572 vp_p.t1154 756.008
R8227 vp_p.n572 vp_p.t218 756.008
R8228 vp_p.n570 vp_p.t1389 756.008
R8229 vp_p.n570 vp_p.t464 756.008
R8230 vp_p.n568 vp_p.t981 756.008
R8231 vp_p.n568 vp_p.t38 756.008
R8232 vp_p.n566 vp_p.t1217 756.008
R8233 vp_p.n566 vp_p.t285 756.008
R8234 vp_p.n564 vp_p.t814 756.008
R8235 vp_p.n564 vp_p.t1368 756.008
R8236 vp_p.n562 vp_p.t232 756.008
R8237 vp_p.n562 vp_p.t803 756.008
R8238 vp_p.n560 vp_p.t474 756.008
R8239 vp_p.n560 vp_p.t1036 756.008
R8240 vp_p.n558 vp_p.t49 756.008
R8241 vp_p.n558 vp_p.t628 756.008
R8242 vp_p.n556 vp_p.t297 756.008
R8243 vp_p.n556 vp_p.t862 756.008
R8244 vp_p.n554 vp_p.t1382 756.008
R8245 vp_p.n554 vp_p.t454 756.008
R8246 vp_p.n552 vp_p.t1450 756.008
R8247 vp_p.n552 vp_p.t529 756.008
R8248 vp_p.n550 vp_p.t1049 756.008
R8249 vp_p.n550 vp_p.t107 756.008
R8250 vp_p.n548 vp_p.t643 756.008
R8251 vp_p.n548 vp_p.t1200 756.008
R8252 vp_p.n546 vp_p.t874 756.008
R8253 vp_p.n546 vp_p.t1429 756.008
R8254 vp_p.n544 vp_p.t468 756.008
R8255 vp_p.n544 vp_p.t1028 756.008
R8256 vp_p.n542 vp_p.t1419 756.008
R8257 vp_p.n542 vp_p.t499 756.008
R8258 vp_p.n540 vp_p.t1015 756.008
R8259 vp_p.n540 vp_p.t76 756.008
R8260 vp_p.n538 vp_p.t609 756.008
R8261 vp_p.n538 vp_p.t1168 756.008
R8262 vp_p.n536 vp_p.t846 756.008
R8263 vp_p.n536 vp_p.t1403 756.008
R8264 vp_p.n534 vp_p.t438 756.008
R8265 vp_p.n534 vp_p.t997 756.008
R8266 vp_p.n532 vp_p.t508 756.008
R8267 vp_p.n532 vp_p.t1072 756.008
R8268 vp_p.n530 vp_p.t88 756.008
R8269 vp_p.n530 vp_p.t662 756.008
R8270 vp_p.n528 vp_p.t329 756.008
R8271 vp_p.n528 vp_p.t896 756.008
R8272 vp_p.n526 vp_p.t1413 756.008
R8273 vp_p.n526 vp_p.t489 756.008
R8274 vp_p.n524 vp_p.t1007 756.008
R8275 vp_p.n524 vp_p.t68 756.008
R8276 vp_p.n522 vp_p.t1081 756.008
R8277 vp_p.n522 vp_p.t140 756.008
R8278 vp_p.n521 vp_p.t676 756.008
R8279 vp_p.n521 vp_p.t1229 756.008
R8280 vp_p.n519 vp_p.t673 756.008
R8281 vp_p.n519 vp_p.t794 756.008
R8282 vp_p.n517 vp_p.t252 756.008
R8283 vp_p.n517 vp_p.t386 756.008
R8284 vp_p.n515 vp_p.t501 756.008
R8285 vp_p.n515 vp_p.t620 756.008
R8286 vp_p.n513 vp_p.t77 756.008
R8287 vp_p.n513 vp_p.t206 756.008
R8288 vp_p.n511 vp_p.t149 756.008
R8289 vp_p.n511 vp_p.t270 756.008
R8290 vp_p.n509 vp_p.t1241 756.008
R8291 vp_p.n509 vp_p.t1362 756.008
R8292 vp_p.n507 vp_p.t835 756.008
R8293 vp_p.n507 vp_p.t957 756.008
R8294 vp_p.n505 vp_p.t1074 756.008
R8295 vp_p.n505 vp_p.t1192 756.008
R8296 vp_p.n503 vp_p.t663 756.008
R8297 vp_p.n503 vp_p.t789 756.008
R8298 vp_p.n501 vp_p.t734 756.008
R8299 vp_p.n501 vp_p.t851 756.008
R8300 vp_p.n499 vp_p.t322 756.008
R8301 vp_p.n499 vp_p.t445 756.008
R8302 vp_p.n497 vp_p.t558 756.008
R8303 vp_p.n497 vp_p.t684 756.008
R8304 vp_p.n495 vp_p.t143 756.008
R8305 vp_p.n495 vp_p.t267 756.008
R8306 vp_p.n493 vp_p.t1231 756.008
R8307 vp_p.n493 vp_p.t1355 756.008
R8308 vp_p.n491 vp_p.t1301 756.008
R8309 vp_p.n491 vp_p.t1421 756.008
R8310 vp_p.n489 vp_p.t899 756.008
R8311 vp_p.n489 vp_p.t1018 756.008
R8312 vp_p.n487 vp_p.t914 756.008
R8313 vp_p.n487 vp_p.t1041 756.008
R8314 vp_p.n485 vp_p.t514 756.008
R8315 vp_p.n485 vp_p.t632 756.008
R8316 vp_p.n483 vp_p.t96 756.008
R8317 vp_p.n483 vp_p.t212 756.008
R8318 vp_p.n481 vp_p.t162 756.008
R8319 vp_p.n481 vp_p.t291 756.008
R8320 vp_p.n479 vp_p.t1255 756.008
R8321 vp_p.n479 vp_p.t1374 756.008
R8322 vp_p.n477 vp_p.t1481 756.008
R8323 vp_p.n477 vp_p.t116 756.008
R8324 vp_p.n475 vp_p.t1087 756.008
R8325 vp_p.n475 vp_p.t1205 756.008
R8326 vp_p.n473 vp_p.t1315 756.008
R8327 vp_p.n473 vp_p.t1437 756.008
R8328 vp_p.n471 vp_p.t746 756.008
R8329 vp_p.n471 vp_p.t868 756.008
R8330 vp_p.n469 vp_p.t336 756.008
R8331 vp_p.n469 vp_p.t461 756.008
R8332 vp_p.n467 vp_p.t567 756.008
R8333 vp_p.n467 vp_p.t703 756.008
R8334 vp_p.n465 vp_p.t156 756.008
R8335 vp_p.n465 vp_p.t282 756.008
R8336 vp_p.n463 vp_p.t397 756.008
R8337 vp_p.n463 vp_p.t522 756.008
R8338 vp_p.n461 vp_p.t1316 756.008
R8339 vp_p.n461 vp_p.t1438 756.008
R8340 vp_p.n459 vp_p.t44 756.008
R8341 vp_p.n459 vp_p.t174 756.008
R8342 vp_p.n457 vp_p.t1139 756.008
R8343 vp_p.n457 vp_p.t1265 756.008
R8344 vp_p.n455 vp_p.t740 756.008
R8345 vp_p.n455 vp_p.t860 756.008
R8346 vp_p.n453 vp_p.t964 756.008
R8347 vp_p.n453 vp_p.t1095 756.008
R8348 vp_p.n451 vp_p.t398 756.008
R8349 vp_p.n451 vp_p.t523 756.008
R8350 vp_p.n449 vp_p.t635 756.008
R8351 vp_p.n449 vp_p.t762 756.008
R8352 vp_p.n447 vp_p.t215 756.008
R8353 vp_p.n447 vp_p.t347 756.008
R8354 vp_p.n445 vp_p.t1307 756.008
R8355 vp_p.n445 vp_p.t1426 756.008
R8356 vp_p.n443 vp_p.t36 756.008
R8357 vp_p.n443 vp_p.t167 756.008
R8358 vp_p.n441 vp_p.t966 756.008
R8359 vp_p.n441 vp_p.t1098 756.008
R8360 vp_p.n439 vp_p.t603 756.008
R8361 vp_p.n439 vp_p.t728 756.008
R8362 vp_p.n437 vp_p.t184 756.008
R8363 vp_p.n437 vp_p.t317 756.008
R8364 vp_p.n435 vp_p.t432 756.008
R8365 vp_p.n435 vp_p.t554 756.008
R8366 vp_p.n433 vp_p.t5 756.008
R8367 vp_p.n433 vp_p.t135 756.008
R8368 vp_p.n431 vp_p.t938 756.008
R8369 vp_p.n431 vp_p.t1068 756.008
R8370 vp_p.n429 vp_p.t1177 756.008
R8371 vp_p.n429 vp_p.t1298 756.008
R8372 vp_p.n427 vp_p.t770 756.008
R8373 vp_p.n427 vp_p.t893 756.008
R8374 vp_p.n425 vp_p.t1003 756.008
R8375 vp_p.n425 vp_p.t1127 756.008
R8376 vp_p.n423 vp_p.t592 756.008
R8377 vp_p.n423 vp_p.t724 756.008
R8378 vp_p.n421 vp_p.t670 756.008
R8379 vp_p.n421 vp_p.t791 756.008
R8380 vp_p.n419 vp_p.t251 756.008
R8381 vp_p.n419 vp_p.t383 756.008
R8382 vp_p.n417 vp_p.t1337 756.008
R8383 vp_p.n417 vp_p.t1464 756.008
R8384 vp_p.n415 vp_p.t74 756.008
R8385 vp_p.n415 vp_p.t199 756.008
R8386 vp_p.n413 vp_p.t1167 756.008
R8387 vp_p.n413 vp_p.t1287 756.008
R8388 vp_p.n411 vp_p.t1239 756.008
R8389 vp_p.n411 vp_p.t1358 756.008
R8390 vp_p.n409 vp_p.t832 756.008
R8391 vp_p.n409 vp_p.t952 756.008
R8392 vp_p.n407 vp_p.t424 756.008
R8393 vp_p.n407 vp_p.t550 756.008
R8394 vp_p.n405 vp_p.t660 756.008
R8395 vp_p.n405 vp_p.t783 756.008
R8396 vp_p.n403 vp_p.t244 756.008
R8397 vp_p.n403 vp_p.t376 756.008
R8398 vp_p.n401 vp_p.t316 756.008
R8399 vp_p.n401 vp_p.t443 756.008
R8400 vp_p.n399 vp_p.t1401 756.008
R8401 vp_p.n399 vp_p.t20 756.008
R8402 vp_p.n397 vp_p.t138 756.008
R8403 vp_p.n397 vp_p.t263 756.008
R8404 vp_p.n395 vp_p.t1227 756.008
R8405 vp_p.n395 vp_p.t1350 756.008
R8406 vp_p.n393 vp_p.t827 756.008
R8407 vp_p.n393 vp_p.t946 756.008
R8408 vp_p.n391 vp_p.t287 756.008
R8409 vp_p.n391 vp_p.t416 756.008
R8410 vp_p.n389 vp_p.t1370 756.008
R8411 vp_p.n389 vp_p.t1490 756.008
R8412 vp_p.n387 vp_p.t111 756.008
R8413 vp_p.n387 vp_p.t235 756.008
R8414 vp_p.n385 vp_p.t1202 756.008
R8415 vp_p.n385 vp_p.t1325 756.008
R8416 vp_p.n383 vp_p.t799 756.008
R8417 vp_p.n383 vp_p.t917 756.008
R8418 vp_p.n381 vp_p.t864 756.008
R8419 vp_p.n381 vp_p.t984 756.008
R8420 vp_p.n379 vp_p.t455 756.008
R8421 vp_p.n379 vp_p.t578 756.008
R8422 vp_p.n377 vp_p.t696 756.008
R8423 vp_p.n377 vp_p.t816 756.008
R8424 vp_p.n375 vp_p.t279 756.008
R8425 vp_p.n375 vp_p.t407 756.008
R8426 vp_p.n373 vp_p.t518 756.008
R8427 vp_p.n373 vp_p.t646 756.008
R8428 vp_p.n372 vp_p.t1431 756.008
R8429 vp_p.n372 vp_p.t53 756.008
R8430 vp_p.n370 vp_p.t587 756.008
R8431 vp_p.n370 vp_p.t797 756.008
R8432 vp_p.n368 vp_p.t821 756.008
R8433 vp_p.n368 vp_p.t1023 756.008
R8434 vp_p.n366 vp_p.t418 756.008
R8435 vp_p.n366 vp_p.t624 756.008
R8436 vp_p.n364 vp_p.t1333 756.008
R8437 vp_p.n364 vp_p.t31 756.008
R8438 vp_p.n362 vp_p.t61 756.008
R8439 vp_p.n362 vp_p.t273 756.008
R8440 vp_p.n360 vp_p.t1161 756.008
R8441 vp_p.n360 vp_p.t1364 756.008
R8442 vp_p.n358 vp_p.t1391 756.008
R8443 vp_p.n358 vp_p.t97 756.008
R8444 vp_p.n356 vp_p.t987 756.008
R8445 vp_p.n356 vp_p.t1196 756.008
R8446 vp_p.n354 vp_p.t1056 756.008
R8447 vp_p.n354 vp_p.t1253 756.008
R8448 vp_p.n352 vp_p.t652 756.008
R8449 vp_p.n352 vp_p.t853 756.008
R8450 vp_p.n350 vp_p.t237 756.008
R8451 vp_p.n350 vp_p.t449 756.008
R8452 vp_p.n348 vp_p.t477 756.008
R8453 vp_p.n348 vp_p.t685 756.008
R8454 vp_p.n346 vp_p.t56 756.008
R8455 vp_p.n346 vp_p.t272 756.008
R8456 vp_p.n344 vp_p.t125 756.008
R8457 vp_p.n344 vp_p.t337 756.008
R8458 vp_p.n342 vp_p.t1220 756.008
R8459 vp_p.n342 vp_p.t1422 756.008
R8460 vp_p.n340 vp_p.t818 756.008
R8461 vp_p.n340 vp_p.t1022 756.008
R8462 vp_p.n338 vp_p.t837 756.008
R8463 vp_p.n338 vp_p.t1045 756.008
R8464 vp_p.n336 vp_p.t429 756.008
R8465 vp_p.n336 vp_p.t641 756.008
R8466 vp_p.n334 vp_p.t502 756.008
R8467 vp_p.n334 vp_p.t709 756.008
R8468 vp_p.n332 vp_p.t79 756.008
R8469 vp_p.n332 vp_p.t294 756.008
R8470 vp_p.n330 vp_p.t324 756.008
R8471 vp_p.n330 vp_p.t535 756.008
R8472 vp_p.n328 vp_p.t1408 756.008
R8473 vp_p.n328 vp_p.t118 756.008
R8474 vp_p.n326 vp_p.t1000 756.008
R8475 vp_p.n326 vp_p.t1211 756.008
R8476 vp_p.n324 vp_p.t1076 756.008
R8477 vp_p.n324 vp_p.t1276 756.008
R8478 vp_p.n322 vp_p.t667 756.008
R8479 vp_p.n322 vp_p.t873 756.008
R8480 vp_p.n320 vp_p.t901 756.008
R8481 vp_p.n320 vp_p.t1108 756.008
R8482 vp_p.n318 vp_p.t494 756.008
R8483 vp_p.n318 vp_p.t708 756.008
R8484 vp_p.n316 vp_p.t71 756.008
R8485 vp_p.n316 vp_p.t292 756.008
R8486 vp_p.n314 vp_p.t145 756.008
R8487 vp_p.n314 vp_p.t360 756.008
R8488 vp_p.n312 vp_p.t1235 756.008
R8489 vp_p.n312 vp_p.t1444 756.008
R8490 vp_p.n310 vp_p.t1468 756.008
R8491 vp_p.n310 vp_p.t179 756.008
R8492 vp_p.n308 vp_p.t1065 756.008
R8493 vp_p.n308 vp_p.t1274 756.008
R8494 vp_p.n306 vp_p.t1293 756.008
R8495 vp_p.n306 vp_p.t0 756.008
R8496 vp_p.n304 vp_p.t727 756.008
R8497 vp_p.n304 vp_p.t931 756.008
R8498 vp_p.n302 vp_p.t313 756.008
R8499 vp_p.n302 vp_p.t532 756.008
R8500 vp_p.n300 vp_p.t553 756.008
R8501 vp_p.n300 vp_p.t767 756.008
R8502 vp_p.n298 vp_p.t133 756.008
R8503 vp_p.n298 vp_p.t357 756.008
R8504 vp_p.n296 vp_p.t381 756.008
R8505 vp_p.n296 vp_p.t588 756.008
R8506 vp_p.n294 vp_p.t1294 756.008
R8507 vp_p.n294 vp_p.t1 756.008
R8508 vp_p.n292 vp_p.t926 756.008
R8509 vp_p.n292 vp_p.t1136 756.008
R8510 vp_p.n290 vp_p.t525 756.008
R8511 vp_p.n290 vp_p.t737 756.008
R8512 vp_p.n288 vp_p.t108 756.008
R8513 vp_p.n288 vp_p.t326 756.008
R8514 vp_p.n286 vp_p.t348 756.008
R8515 vp_p.n286 vp_p.t560 756.008
R8516 vp_p.n284 vp_p.t1267 756.008
R8517 vp_p.n284 vp_p.t1474 756.008
R8518 vp_p.n282 vp_p.t1493 756.008
R8519 vp_p.n282 vp_p.t211 756.008
R8520 vp_p.n280 vp_p.t1099 756.008
R8521 vp_p.n280 vp_p.t1304 756.008
R8522 vp_p.n278 vp_p.t693 756.008
R8523 vp_p.n278 vp_p.t903 756.008
R8524 vp_p.n276 vp_p.t922 756.008
R8525 vp_p.n276 vp_p.t1133 756.008
R8526 vp_p.n274 vp_p.t350 756.008
R8527 vp_p.n274 vp_p.t561 756.008
R8528 vp_p.n272 vp_p.t583 756.008
R8529 vp_p.n272 vp_p.t796 756.008
R8530 vp_p.n270 vp_p.t169 756.008
R8531 vp_p.n270 vp_p.t390 756.008
R8532 vp_p.n268 vp_p.t413 756.008
R8533 vp_p.n268 vp_p.t622 756.008
R8534 vp_p.n266 vp_p.t1486 756.008
R8535 vp_p.n266 vp_p.t208 756.008
R8536 vp_p.n264 vp_p.t923 756.008
R8537 vp_p.n264 vp_p.t1134 756.008
R8538 vp_p.n262 vp_p.t1157 756.008
R8539 vp_p.n262 vp_p.t1363 756.008
R8540 vp_p.n260 vp_p.t755 756.008
R8541 vp_p.n260 vp_p.t959 756.008
R8542 vp_p.n258 vp_p.t982 756.008
R8543 vp_p.n258 vp_p.t1194 756.008
R8544 vp_p.n256 vp_p.t576 756.008
R8545 vp_p.n256 vp_p.t793 756.008
R8546 vp_p.n254 vp_p.t651 756.008
R8547 vp_p.n254 vp_p.t852 756.008
R8548 vp_p.n252 vp_p.t234 756.008
R8549 vp_p.n252 vp_p.t447 756.008
R8550 vp_p.n250 vp_p.t1323 756.008
R8551 vp_p.n250 vp_p.t28 756.008
R8552 vp_p.n248 vp_p.t51 756.008
R8553 vp_p.n248 vp_p.t269 756.008
R8554 vp_p.n246 vp_p.t1149 756.008
R8555 vp_p.n246 vp_p.t1361 756.008
R8556 vp_p.n244 vp_p.t618 756.008
R8557 vp_p.n244 vp_p.t823 756.008
R8558 vp_p.n242 vp_p.t203 756.008
R8559 vp_p.n242 vp_p.t421 756.008
R8560 vp_p.n240 vp_p.t1289 756.008
R8561 vp_p.n240 vp_p.t1497 756.008
R8562 vp_p.n238 vp_p.t22 756.008
R8563 vp_p.n238 vp_p.t241 756.008
R8564 vp_p.n236 vp_p.t1122 756.008
R8565 vp_p.n236 vp_p.t1334 756.008
R8566 vp_p.n234 vp_p.t1193 756.008
R8567 vp_p.n234 vp_p.t1392 756.008
R8568 vp_p.n232 vp_p.t786 756.008
R8569 vp_p.n232 vp_p.t990 756.008
R8570 vp_p.n230 vp_p.t1017 756.008
R8571 vp_p.n230 vp_p.t1221 756.008
R8572 vp_p.n228 vp_p.t610 756.008
R8573 vp_p.n228 vp_p.t822 756.008
R8574 vp_p.n226 vp_p.t195 756.008
R8575 vp_p.n226 vp_p.t419 756.008
R8576 vp_p.n224 vp_p.t265 756.008
R8577 vp_p.n224 vp_p.t480 756.008
R8578 vp_p.n223 vp_p.t1352 756.008
R8579 vp_p.n223 vp_p.t62 756.008
R8580 vp_p.n221 vp_p.t993 756.008
R8581 vp_p.n221 vp_p.t54 756.008
R8582 vp_p.n219 vp_p.t590 756.008
R8583 vp_p.n219 vp_p.t1150 756.008
R8584 vp_p.n217 vp_p.t824 756.008
R8585 vp_p.n217 vp_p.t1386 756.008
R8586 vp_p.n215 vp_p.t422 756.008
R8587 vp_p.n215 vp_p.t978 756.008
R8588 vp_p.n213 vp_p.t483 756.008
R8589 vp_p.n213 vp_p.t1053 756.008
R8590 vp_p.n211 vp_p.t65 756.008
R8591 vp_p.n211 vp_p.t647 756.008
R8592 vp_p.n209 vp_p.t1164 756.008
R8593 vp_p.n209 vp_p.t230 756.008
R8594 vp_p.n207 vp_p.t1393 756.008
R8595 vp_p.n207 vp_p.t471 756.008
R8596 vp_p.n205 vp_p.t991 756.008
R8597 vp_p.n205 vp_p.t47 756.008
R8598 vp_p.n203 vp_p.t1057 756.008
R8599 vp_p.n203 vp_p.t122 756.008
R8600 vp_p.n201 vp_p.t654 756.008
R8601 vp_p.n201 vp_p.t1215 756.008
R8602 vp_p.n199 vp_p.t881 756.008
R8603 vp_p.n199 vp_p.t1446 756.008
R8604 vp_p.n197 vp_p.t481 756.008
R8605 vp_p.n197 vp_p.t1046 756.008
R8606 vp_p.n195 vp_p.t63 756.008
R8607 vp_p.n195 vp_p.t642 756.008
R8608 vp_p.n193 vp_p.t126 756.008
R8609 vp_p.n193 vp_p.t710 756.008
R8610 vp_p.n191 vp_p.t1222 756.008
R8611 vp_p.n191 vp_p.t295 756.008
R8612 vp_p.n189 vp_p.t1242 756.008
R8613 vp_p.n189 vp_p.t309 756.008
R8614 vp_p.n187 vp_p.t842 756.008
R8615 vp_p.n187 vp_p.t1397 756.008
R8616 vp_p.n185 vp_p.t437 756.008
R8617 vp_p.n185 vp_p.t995 756.008
R8618 vp_p.n183 vp_p.t504 756.008
R8619 vp_p.n183 vp_p.t1063 756.008
R8620 vp_p.n181 vp_p.t84 756.008
R8621 vp_p.n181 vp_p.t657 756.008
R8622 vp_p.n179 vp_p.t327 756.008
R8623 vp_p.n179 vp_p.t890 756.008
R8624 vp_p.n177 vp_p.t1412 756.008
R8625 vp_p.n177 vp_p.t487 756.008
R8626 vp_p.n175 vp_p.t150 756.008
R8627 vp_p.n175 vp_p.t720 756.008
R8628 vp_p.n173 vp_p.t1079 756.008
R8629 vp_p.n173 vp_p.t134 756.008
R8630 vp_p.n171 vp_p.t674 756.008
R8631 vp_p.n171 vp_p.t1225 756.008
R8632 vp_p.n169 vp_p.t906 756.008
R8633 vp_p.n169 vp_p.t1461 756.008
R8634 vp_p.n167 vp_p.t503 756.008
R8635 vp_p.n167 vp_p.t1061 756.008
R8636 vp_p.n165 vp_p.t735 756.008
R8637 vp_p.n165 vp_p.t1284 756.008
R8638 vp_p.n163 vp_p.t151 756.008
R8639 vp_p.n163 vp_p.t721 756.008
R8640 vp_p.n161 vp_p.t391 756.008
R8641 vp_p.n161 vp_p.t949 756.008
R8642 vp_p.n159 vp_p.t1473 756.008
R8643 vp_p.n159 vp_p.t547 756.008
R8644 vp_p.n157 vp_p.t1077 756.008
R8645 vp_p.n157 vp_p.t131 756.008
R8646 vp_p.n155 vp_p.t1302 756.008
R8647 vp_p.n155 vp_p.t373 756.008
R8648 vp_p.n153 vp_p.t736 756.008
R8649 vp_p.n153 vp_p.t1285 756.008
R8650 vp_p.n151 vp_p.t960 756.008
R8651 vp_p.n151 vp_p.t18 756.008
R8652 vp_p.n149 vp_p.t559 756.008
R8653 vp_p.n149 vp_p.t1118 756.008
R8654 vp_p.n147 vp_p.t146 756.008
R8655 vp_p.n147 vp_p.t719 756.008
R8656 vp_p.n145 vp_p.t388 756.008
R8657 vp_p.n145 vp_p.t944 756.008
R8658 vp_p.n143 vp_p.t1303 756.008
R8659 vp_p.n143 vp_p.t374 756.008
R8660 vp_p.n141 vp_p.t932 756.008
R8661 vp_p.n141 vp_p.t1487 756.008
R8662 vp_p.n139 vp_p.t534 756.008
R8663 vp_p.n139 vp_p.t1092 756.008
R8664 vp_p.n137 vp_p.t768 756.008
R8665 vp_p.n137 vp_p.t1322 756.008
R8666 vp_p.n135 vp_p.t358 756.008
R8667 vp_p.n135 vp_p.t916 756.008
R8668 vp_p.n133 vp_p.t1275 756.008
R8669 vp_p.n133 vp_p.t344 756.008
R8670 vp_p.n131 vp_p.t2 756.008
R8671 vp_p.n131 vp_p.t577 756.008
R8672 vp_p.n129 vp_p.t1106 756.008
R8673 vp_p.n129 vp_p.t163 756.008
R8674 vp_p.n127 vp_p.t1335 756.008
R8675 vp_p.n127 vp_p.t406 756.008
R8676 vp_p.n125 vp_p.t928 756.008
R8677 vp_p.n125 vp_p.t1482 756.008
R8678 vp_p.n123 vp_p.t992 756.008
R8679 vp_p.n123 vp_p.t50 756.008
R8680 vp_p.n121 vp_p.t589 756.008
R8681 vp_p.n121 vp_p.t1148 756.008
R8682 vp_p.n119 vp_p.t178 756.008
R8683 vp_p.n119 vp_p.t750 756.008
R8684 vp_p.n117 vp_p.t420 756.008
R8685 vp_p.n117 vp_p.t975 756.008
R8686 vp_p.n115 vp_p.t1494 756.008
R8687 vp_p.n115 vp_p.t569 756.008
R8688 vp_p.n113 vp_p.t64 756.008
R8689 vp_p.n113 vp_p.t645 756.008
R8690 vp_p.n111 vp_p.t1163 756.008
R8691 vp_p.n111 vp_p.t228 756.008
R8692 vp_p.n109 vp_p.t765 756.008
R8693 vp_p.n109 vp_p.t1320 756.008
R8694 vp_p.n107 vp_p.t989 756.008
R8695 vp_p.n107 vp_p.t45 756.008
R8696 vp_p.n105 vp_p.t586 756.008
R8697 vp_p.n105 vp_p.t1145 756.008
R8698 vp_p.n103 vp_p.t653 756.008
R8699 vp_p.n103 vp_p.t1213 756.008
R8700 vp_p.n101 vp_p.t239 756.008
R8701 vp_p.n101 vp_p.t810 756.008
R8702 vp_p.n99 vp_p.t479 756.008
R8703 vp_p.n99 vp_p.t1043 756.008
R8704 vp_p.n97 vp_p.t60 756.008
R8705 vp_p.n97 vp_p.t638 756.008
R8706 vp_p.n95 vp_p.t1160 756.008
R8707 vp_p.n95 vp_p.t224 756.008
R8708 vp_p.n93 vp_p.t623 756.008
R8709 vp_p.n93 vp_p.t1184 756.008
R8710 vp_p.n91 vp_p.t209 756.008
R8711 vp_p.n91 vp_p.t781 756.008
R8712 vp_p.n89 vp_p.t448 756.008
R8713 vp_p.n89 vp_p.t1010 756.008
R8714 vp_p.n87 vp_p.t30 756.008
R8715 vp_p.n87 vp_p.t606 756.008
R8716 vp_p.n85 vp_p.t1131 756.008
R8717 vp_p.n85 vp_p.t190 756.008
R8718 vp_p.n83 vp_p.t1195 756.008
R8719 vp_p.n83 vp_p.t258 756.008
R8720 vp_p.n81 vp_p.t795 756.008
R8721 vp_p.n81 vp_p.t1347 756.008
R8722 vp_p.n79 vp_p.t1021 756.008
R8723 vp_p.n79 vp_p.t83 756.008
R8724 vp_p.n77 vp_p.t621 756.008
R8725 vp_p.n77 vp_p.t1181 756.008
R8726 vp_p.n75 vp_p.t850 756.008
R8727 vp_p.n75 vp_p.t1411 756.008
R8728 vp_p.n74 vp_p.t271 756.008
R8729 vp_p.n74 vp_p.t841 756.008
R8730 vp_p.n970 vp_p.t268 756.008
R8731 vp_p.n970 vp_p.t839 756.008
R8732 vp_p.n968 vp_p.t510 756.008
R8733 vp_p.n968 vp_p.t1078 756.008
R8734 vp_p.n966 vp_p.t94 756.008
R8735 vp_p.n966 vp_p.t671 756.008
R8736 vp_p.n964 vp_p.t1019 756.008
R8737 vp_p.n964 vp_p.t80 756.008
R8738 vp_p.n962 vp_p.t1249 756.008
R8739 vp_p.n962 vp_p.t325 756.008
R8740 vp_p.n960 vp_p.t849 756.008
R8741 vp_p.n960 vp_p.t1409 756.008
R8742 vp_p.n958 vp_p.t1083 756.008
R8743 vp_p.n958 vp_p.t147 756.008
R8744 vp_p.n956 vp_p.t681 756.008
R8745 vp_p.n956 vp_p.t1237 756.008
R8746 vp_p.n954 vp_p.t739 756.008
R8747 vp_p.n954 vp_p.t1305 756.008
R8748 vp_p.n952 vp_p.t333 756.008
R8749 vp_p.n952 vp_p.t904 756.008
R8750 vp_p.n950 vp_p.t1418 756.008
R8751 vp_p.n950 vp_p.t496 756.008
R8752 vp_p.n948 vp_p.t152 756.008
R8753 vp_p.n948 vp_p.t730 756.008
R8754 vp_p.n946 vp_p.t1246 756.008
R8755 vp_p.n946 vp_p.t319 756.008
R8756 vp_p.n944 vp_p.t1306 756.008
R8757 vp_p.n944 vp_p.t389 756.008
R8758 vp_p.n942 vp_p.t908 756.008
R8759 vp_p.n942 vp_p.t1470 756.008
R8760 vp_p.n940 vp_p.t507 756.008
R8761 vp_p.n940 vp_p.t1070 756.008
R8762 vp_p.n938 vp_p.t526 756.008
R8763 vp_p.n938 vp_p.t1089 756.008
R8764 vp_p.n936 vp_p.t104 756.008
R8765 vp_p.n936 vp_p.t687 756.008
R8766 vp_p.n934 vp_p.t175 756.008
R8767 vp_p.n934 vp_p.t748 756.008
R8768 vp_p.n932 vp_p.t1268 756.008
R8769 vp_p.n932 vp_p.t340 756.008
R8770 vp_p.n930 vp_p.t1495 756.008
R8771 vp_p.n930 vp_p.t570 756.008
R8772 vp_p.n928 vp_p.t1100 756.008
R8773 vp_p.n928 vp_p.t159 756.008
R8774 vp_p.n926 vp_p.t694 756.008
R8775 vp_p.n926 vp_p.t1252 756.008
R8776 vp_p.n924 vp_p.t763 756.008
R8777 vp_p.n924 vp_p.t1318 756.008
R8778 vp_p.n922 vp_p.t351 756.008
R8779 vp_p.n922 vp_p.t911 756.008
R8780 vp_p.n920 vp_p.t584 756.008
R8781 vp_p.n920 vp_p.t1143 756.008
R8782 vp_p.n918 vp_p.t170 756.008
R8783 vp_p.n918 vp_p.t743 756.008
R8784 vp_p.n916 vp_p.t1260 756.008
R8785 vp_p.n916 vp_p.t335 756.008
R8786 vp_p.n914 vp_p.t1331 756.008
R8787 vp_p.n914 vp_p.t402 756.008
R8788 vp_p.n912 vp_p.t924 756.008
R8789 vp_p.n912 vp_p.t1479 756.008
R8790 vp_p.n910 vp_p.t1158 756.008
R8791 vp_p.n910 vp_p.t221 756.008
R8792 vp_p.n908 vp_p.t756 756.008
R8793 vp_p.n908 vp_p.t1311 756.008
R8794 vp_p.n906 vp_p.t983 756.008
R8795 vp_p.n906 vp_p.t39 756.008
R8796 vp_p.n904 vp_p.t414 756.008
R8797 vp_p.n904 vp_p.t969 756.008
R8798 vp_p.n902 vp_p.t1488 756.008
R8799 vp_p.n902 vp_p.t564 756.008
R8800 vp_p.n900 vp_p.t233 756.008
R8801 vp_p.n900 vp_p.t804 756.008
R8802 vp_p.n898 vp_p.t1324 756.008
R8803 vp_p.n898 vp_p.t393 756.008
R8804 vp_p.n896 vp_p.t52 756.008
R8805 vp_p.n896 vp_p.t629 756.008
R8806 vp_p.n894 vp_p.t985 756.008
R8807 vp_p.n894 vp_p.t41 756.008
R8808 vp_p.n892 vp_p.t619 756.008
R8809 vp_p.n892 vp_p.t1180 756.008
R8810 vp_p.n890 vp_p.t204 756.008
R8811 vp_p.n890 vp_p.t776 756.008
R8812 vp_p.n888 vp_p.t1290 756.008
R8813 vp_p.n888 vp_p.t364 756.008
R8814 vp_p.n886 vp_p.t23 756.008
R8815 vp_p.n886 vp_p.t596 756.008
R8816 vp_p.n884 vp_p.t955 756.008
R8817 vp_p.n884 vp_p.t11 756.008
R8818 vp_p.n882 vp_p.t1191 756.008
R8819 vp_p.n882 vp_p.t253 756.008
R8820 vp_p.n880 vp_p.t788 756.008
R8821 vp_p.n880 vp_p.t1341 756.008
R8822 vp_p.n878 vp_p.t377 756.008
R8823 vp_p.n878 vp_p.t934 756.008
R8824 vp_p.n876 vp_p.t612 756.008
R8825 vp_p.n876 vp_p.t1170 756.008
R8826 vp_p.n874 vp_p.t24 756.008
R8827 vp_p.n874 vp_p.t597 756.008
R8828 vp_p.n872 vp_p.t266 756.008
R8829 vp_p.n872 vp_p.t836 756.008
R8830 vp_p.n870 vp_p.t1354 756.008
R8831 vp_p.n870 vp_p.t426 756.008
R8832 vp_p.n868 vp_p.t91 756.008
R8833 vp_p.n868 vp_p.t665 756.008
R8834 vp_p.n866 vp_p.t1185 756.008
R8835 vp_p.n866 vp_p.t246 756.008
R8836 vp_p.n864 vp_p.t613 756.008
R8837 vp_p.n864 vp_p.t1171 756.008
R8838 vp_p.n862 vp_p.t848 756.008
R8839 vp_p.n862 vp_p.t1406 756.008
R8840 vp_p.n860 vp_p.t440 756.008
R8841 vp_p.n860 vp_p.t998 756.008
R8842 vp_p.n858 vp_p.t678 756.008
R8843 vp_p.n858 vp_p.t1232 756.008
R8844 vp_p.n856 vp_p.t260 756.008
R8845 vp_p.n856 vp_p.t829 756.008
R8846 vp_p.n854 vp_p.t332 756.008
R8847 vp_p.n854 vp_p.t902 756.008
R8848 vp_p.n852 vp_p.t1415 756.008
R8849 vp_p.n852 vp_p.t492 756.008
R8850 vp_p.n850 vp_p.t1011 756.008
R8851 vp_p.n850 vp_p.t69 756.008
R8852 vp_p.n848 vp_p.t1244 756.008
R8853 vp_p.n848 vp_p.t310 756.008
R8854 vp_p.n846 vp_p.t844 756.008
R8855 vp_p.n846 vp_p.t1398 756.008
R8856 vp_p.n844 vp_p.t300 756.008
R8857 vp_p.n844 vp_p.t869 756.008
R8858 vp_p.n842 vp_p.t1387 756.008
R8859 vp_p.n842 vp_p.t458 756.008
R8860 vp_p.n840 vp_p.t979 756.008
R8861 vp_p.n840 vp_p.t35 756.008
R8862 vp_p.n838 vp_p.t1216 756.008
R8863 vp_p.n838 vp_p.t283 756.008
R8864 vp_p.n836 vp_p.t813 756.008
R8865 vp_p.n836 vp_p.t1366 756.008
R8866 vp_p.n834 vp_p.t877 756.008
R8867 vp_p.n834 vp_p.t1439 756.008
R8868 vp_p.n832 vp_p.t472 756.008
R8869 vp_p.n832 vp_p.t1033 756.008
R8870 vp_p.n830 vp_p.t711 756.008
R8871 vp_p.n830 vp_p.t1266 756.008
R8872 vp_p.n828 vp_p.t296 756.008
R8873 vp_p.n828 vp_p.t858 756.008
R8874 vp_p.n826 vp_p.t1381 756.008
R8875 vp_p.n826 vp_p.t452 756.008
R8876 vp_p.n824 vp_p.t1448 756.008
R8877 vp_p.n824 vp_p.t524 756.008
R8878 vp_p.n823 vp_p.t1048 756.008
R8879 vp_p.n823 vp_p.t105 756.008
R8880 vp_p.n1119 vp_p.t1042 756.008
R8881 vp_p.n1119 vp_p.t177 756.008
R8882 vp_p.n1117 vp_p.t636 756.008
R8883 vp_p.n1117 vp_p.t1270 756.008
R8884 vp_p.n1115 vp_p.t871 756.008
R8885 vp_p.n1115 vp_p.t1496 756.008
R8886 vp_p.n1113 vp_p.t462 756.008
R8887 vp_p.n1113 vp_p.t1101 756.008
R8888 vp_p.n1111 vp_p.t533 756.008
R8889 vp_p.n1111 vp_p.t1162 756.008
R8890 vp_p.n1109 vp_p.t117 756.008
R8891 vp_p.n1109 vp_p.t764 756.008
R8892 vp_p.n1107 vp_p.t1208 756.008
R8893 vp_p.n1107 vp_p.t352 756.008
R8894 vp_p.n1105 vp_p.t1440 756.008
R8895 vp_p.n1105 vp_p.t585 756.008
R8896 vp_p.n1103 vp_p.t1034 756.008
R8897 vp_p.n1103 vp_p.t171 756.008
R8898 vp_p.n1101 vp_p.t1107 756.008
R8899 vp_p.n1101 vp_p.t240 756.008
R8900 vp_p.n1099 vp_p.t704 756.008
R8901 vp_p.n1099 vp_p.t1332 756.008
R8902 vp_p.n1097 vp_p.t927 756.008
R8903 vp_p.n1097 vp_p.t59 756.008
R8904 vp_p.n1095 vp_p.t527 756.008
R8905 vp_p.n1095 vp_p.t1159 756.008
R8906 vp_p.n1093 vp_p.t109 756.008
R8907 vp_p.n1093 vp_p.t757 756.008
R8908 vp_p.n1091 vp_p.t176 756.008
R8909 vp_p.n1091 vp_p.t820 756.008
R8910 vp_p.n1089 vp_p.t1269 756.008
R8911 vp_p.n1089 vp_p.t415 756.008
R8912 vp_p.n1087 vp_p.t1282 756.008
R8913 vp_p.n1087 vp_p.t434 756.008
R8914 vp_p.n1085 vp_p.t885 756.008
R8915 vp_p.n1085 vp_p.t7 756.008
R8916 vp_p.n1083 vp_p.t482 756.008
R8917 vp_p.n1083 vp_p.t1112 756.008
R8918 vp_p.n1081 vp_p.t544 756.008
R8919 vp_p.n1081 vp_p.t1178 756.008
R8920 vp_p.n1079 vp_p.t129 756.008
R8921 vp_p.n1079 vp_p.t774 756.008
R8922 vp_p.n1077 vp_p.t369 756.008
R8923 vp_p.n1077 vp_p.t1004 756.008
R8924 vp_p.n1075 vp_p.t1456 756.008
R8925 vp_p.n1075 vp_p.t595 756.008
R8926 vp_p.n1073 vp_p.t187 756.008
R8927 vp_p.n1073 vp_p.t833 756.008
R8928 vp_p.n1071 vp_p.t1115 756.008
R8929 vp_p.n1071 vp_p.t254 756.008
R8930 vp_p.n1069 vp_p.t715 756.008
R8931 vp_p.n1069 vp_p.t1340 756.008
R8932 vp_p.n1067 vp_p.t940 756.008
R8933 vp_p.n1067 vp_p.t78 756.008
R8934 vp_p.n1065 vp_p.t540 756.008
R8935 vp_p.n1065 vp_p.t1169 756.008
R8936 vp_p.n1063 vp_p.t771 756.008
R8937 vp_p.n1063 vp_p.t1404 756.008
R8938 vp_p.n1061 vp_p.t188 756.008
R8939 vp_p.n1061 vp_p.t834 756.008
R8940 vp_p.n1059 vp_p.t433 756.008
R8941 vp_p.n1059 vp_p.t1075 756.008
R8942 vp_p.n1057 vp_p.t9 756.008
R8943 vp_p.n1057 vp_p.t664 756.008
R8944 vp_p.n1055 vp_p.t1111 756.008
R8945 vp_p.n1055 vp_p.t245 756.008
R8946 vp_p.n1053 vp_p.t1338 756.008
R8947 vp_p.n1053 vp_p.t490 756.008
R8948 vp_p.n1051 vp_p.t773 756.008
R8949 vp_p.n1051 vp_p.t1405 756.008
R8950 vp_p.n1049 vp_p.t1005 756.008
R8951 vp_p.n1049 vp_p.t144 756.008
R8952 vp_p.n1047 vp_p.t594 756.008
R8953 vp_p.n1047 vp_p.t1230 756.008
R8954 vp_p.n1045 vp_p.t181 756.008
R8955 vp_p.n1045 vp_p.t828 756.008
R8956 vp_p.n1043 vp_p.t425 756.008
R8957 vp_p.n1043 vp_p.t1062 756.008
R8958 vp_p.n1041 vp_p.t1339 756.008
R8959 vp_p.n1041 vp_p.t491 756.008
R8960 vp_p.n1039 vp_p.t973 756.008
R8961 vp_p.n1039 vp_p.t115 756.008
R8962 vp_p.n1037 vp_p.t565 756.008
R8963 vp_p.n1037 vp_p.t1204 756.008
R8964 vp_p.n1035 vp_p.t806 756.008
R8965 vp_p.n1035 vp_p.t1436 756.008
R8966 vp_p.n1033 vp_p.t395 756.008
R8967 vp_p.n1033 vp_p.t1032 756.008
R8968 vp_p.n1031 vp_p.t1313 756.008
R8969 vp_p.n1031 vp_p.t459 756.008
R8970 vp_p.n1029 vp_p.t42 756.008
R8971 vp_p.n1029 vp_p.t702 756.008
R8972 vp_p.n1027 vp_p.t1137 756.008
R8973 vp_p.n1027 vp_p.t281 756.008
R8974 vp_p.n1025 vp_p.t1372 756.008
R8975 vp_p.n1025 vp_p.t521 756.008
R8976 vp_p.n1023 vp_p.t962 756.008
R8977 vp_p.n1023 vp_p.t101 756.008
R8978 vp_p.n1021 vp_p.t1040 756.008
R8979 vp_p.n1021 vp_p.t173 756.008
R8980 vp_p.n1019 vp_p.t631 756.008
R8981 vp_p.n1019 vp_p.t1264 756.008
R8982 vp_p.n1017 vp_p.t213 756.008
R8983 vp_p.n1017 vp_p.t859 756.008
R8984 vp_p.n1015 vp_p.t456 756.008
R8985 vp_p.n1015 vp_p.t1094 756.008
R8986 vp_p.n1013 vp_p.t34 756.008
R8987 vp_p.n1013 vp_p.t690 756.008
R8988 vp_p.n1011 vp_p.t114 756.008
R8989 vp_p.n1011 vp_p.t761 756.008
R8990 vp_p.n1009 vp_p.t1206 756.008
R8991 vp_p.n1009 vp_p.t346 756.008
R8992 vp_p.n1007 vp_p.t800 756.008
R8993 vp_p.n1007 vp_p.t1425 756.008
R8994 vp_p.n1005 vp_p.t1031 756.008
R8995 vp_p.n1005 vp_p.t166 756.008
R8996 vp_p.n1003 vp_p.t626 756.008
R8997 vp_p.n1003 vp_p.t1259 756.008
R8998 vp_p.n1001 vp_p.t700 756.008
R8999 vp_p.n1001 vp_p.t1329 756.008
R9000 vp_p.n999 vp_p.t280 756.008
R9001 vp_p.n999 vp_p.t919 756.008
R9002 vp_p.n997 vp_p.t520 756.008
R9003 vp_p.n997 vp_p.t1155 756.008
R9004 vp_p.n995 vp_p.t103 756.008
R9005 vp_p.n995 vp_p.t753 756.008
R9006 vp_p.n993 vp_p.t1198 756.008
R9007 vp_p.n993 vp_p.t342 756.008
R9008 vp_p.n991 vp_p.t668 756.008
R9009 vp_p.n991 vp_p.t1297 756.008
R9010 vp_p.n989 vp_p.t247 756.008
R9011 vp_p.n989 vp_p.t892 756.008
R9012 vp_p.n987 vp_p.t495 756.008
R9013 vp_p.n987 vp_p.t1126 756.008
R9014 vp_p.n985 vp_p.t72 756.008
R9015 vp_p.n985 vp_p.t723 756.008
R9016 vp_p.n983 vp_p.t1166 756.008
R9017 vp_p.n983 vp_p.t307 756.008
R9018 vp_p.n981 vp_p.t1236 756.008
R9019 vp_p.n981 vp_p.t382 756.008
R9020 vp_p.n979 vp_p.t830 756.008
R9021 vp_p.n979 vp_p.t1463 756.008
R9022 vp_p.n977 vp_p.t1066 756.008
R9023 vp_p.n977 vp_p.t198 756.008
R9024 vp_p.n975 vp_p.t658 756.008
R9025 vp_p.n975 vp_p.t1286 756.008
R9026 vp_p.n973 vp_p.t891 756.008
R9027 vp_p.n973 vp_p.t19 756.008
R9028 vp_p.n972 vp_p.t314 756.008
R9029 vp_p.n972 vp_p.t951 756.008
R9030 vp_p.n1268 vp_p.t1471 756.008
R9031 vp_p.n1268 vp_p.t545 756.008
R9032 vp_p.n1266 vp_p.t207 756.008
R9033 vp_p.n1266 vp_p.t780 756.008
R9034 vp_p.n1264 vp_p.t1296 756.008
R9035 vp_p.n1264 vp_p.t370 756.008
R9036 vp_p.n1262 vp_p.t731 756.008
R9037 vp_p.n1262 vp_p.t1283 756.008
R9038 vp_p.n1260 vp_p.t958 756.008
R9039 vp_p.n1260 vp_p.t15 756.008
R9040 vp_p.n1258 vp_p.t556 756.008
R9041 vp_p.n1258 vp_p.t1116 756.008
R9042 vp_p.n1256 vp_p.t792 756.008
R9043 vp_p.n1256 vp_p.t1345 756.008
R9044 vp_p.n1254 vp_p.t385 756.008
R9045 vp_p.n1254 vp_p.t941 756.008
R9046 vp_p.n1252 vp_p.t446 756.008
R9047 vp_p.n1252 vp_p.t1008 756.008
R9048 vp_p.n1250 vp_p.t29 756.008
R9049 vp_p.n1250 vp_p.t605 756.008
R9050 vp_p.n1248 vp_p.t1130 756.008
R9051 vp_p.n1248 vp_p.t189 756.008
R9052 vp_p.n1246 vp_p.t1360 756.008
R9053 vp_p.n1246 vp_p.t435 756.008
R9054 vp_p.n1244 vp_p.t954 756.008
R9055 vp_p.n1244 vp_p.t10 756.008
R9056 vp_p.n1242 vp_p.t1020 756.008
R9057 vp_p.n1242 vp_p.t82 756.008
R9058 vp_p.n1240 vp_p.t617 756.008
R9059 vp_p.n1240 vp_p.t1179 756.008
R9060 vp_p.n1238 vp_p.t202 756.008
R9061 vp_p.n1238 vp_p.t775 756.008
R9062 vp_p.n1236 vp_p.t222 756.008
R9063 vp_p.n1236 vp_p.t798 756.008
R9064 vp_p.n1234 vp_p.t1309 756.008
R9065 vp_p.n1234 vp_p.t392 756.008
R9066 vp_p.n1232 vp_p.t1378 756.008
R9067 vp_p.n1232 vp_p.t451 756.008
R9068 vp_p.n1230 vp_p.t970 756.008
R9069 vp_p.n1230 vp_p.t33 756.008
R9070 vp_p.n1228 vp_p.t1210 756.008
R9071 vp_p.n1228 vp_p.t276 756.008
R9072 vp_p.n1226 vp_p.t805 756.008
R9073 vp_p.n1226 vp_p.t1365 756.008
R9074 vp_p.n1224 vp_p.t394 756.008
R9075 vp_p.n1224 vp_p.t961 756.008
R9076 vp_p.n1222 vp_p.t467 756.008
R9077 vp_p.n1222 vp_p.t1026 756.008
R9078 vp_p.n1220 vp_p.t40 756.008
R9079 vp_p.n1220 vp_p.t625 756.008
R9080 vp_p.n1218 vp_p.t288 756.008
R9081 vp_p.n1218 vp_p.t855 756.008
R9082 vp_p.n1216 vp_p.t1371 756.008
R9083 vp_p.n1216 vp_p.t450 756.008
R9084 vp_p.n1214 vp_p.t963 756.008
R9085 vp_p.n1214 vp_p.t32 756.008
R9086 vp_p.n1212 vp_p.t1037 756.008
R9087 vp_p.n1212 vp_p.t100 756.008
R9088 vp_p.n1210 vp_p.t630 756.008
R9089 vp_p.n1210 vp_p.t1197 756.008
R9090 vp_p.n1208 vp_p.t867 756.008
R9091 vp_p.n1208 vp_p.t1424 756.008
R9092 vp_p.n1206 vp_p.t457 756.008
R9093 vp_p.n1206 vp_p.t1024 756.008
R9094 vp_p.n1204 vp_p.t697 756.008
R9095 vp_p.n1204 vp_p.t1254 756.008
R9096 vp_p.n1202 vp_p.t113 756.008
R9097 vp_p.n1202 vp_p.t688 756.008
R9098 vp_p.n1200 vp_p.t1203 756.008
R9099 vp_p.n1200 vp_p.t274 756.008
R9100 vp_p.n1198 vp_p.t1432 756.008
R9101 vp_p.n1198 vp_p.t512 756.008
R9102 vp_p.n1196 vp_p.t1030 756.008
R9103 vp_p.n1196 vp_p.t98 756.008
R9104 vp_p.n1194 vp_p.t1262 756.008
R9105 vp_p.n1194 vp_p.t338 756.008
R9106 vp_p.n1192 vp_p.t701 756.008
R9107 vp_p.n1192 vp_p.t1256 756.008
R9108 vp_p.n1190 vp_p.t323 756.008
R9109 vp_p.n1190 vp_p.t886 756.008
R9110 vp_p.n1188 vp_p.t1407 756.008
R9111 vp_p.n1188 vp_p.t486 756.008
R9112 vp_p.n1186 vp_p.t999 756.008
R9113 vp_p.n1186 vp_p.t66 756.008
R9114 vp_p.n1184 vp_p.t1233 756.008
R9115 vp_p.n1184 vp_p.t305 756.008
R9116 vp_p.n1182 vp_p.t666 756.008
R9117 vp_p.n1182 vp_p.t1224 756.008
R9118 vp_p.n1180 vp_p.t900 756.008
R9119 vp_p.n1180 vp_p.t1459 756.008
R9120 vp_p.n1178 vp_p.t493 756.008
R9121 vp_p.n1178 vp_p.t1060 756.008
R9122 vp_p.n1176 vp_p.t70 756.008
R9123 vp_p.n1176 vp_p.t655 756.008
R9124 vp_p.n1174 vp_p.t311 756.008
R9125 vp_p.n1174 vp_p.t883 756.008
R9126 vp_p.n1172 vp_p.t1234 756.008
R9127 vp_p.n1172 vp_p.t306 756.008
R9128 vp_p.n1170 vp_p.t1467 756.008
R9129 vp_p.n1170 vp_p.t543 756.008
R9130 vp_p.n1168 vp_p.t1064 756.008
R9131 vp_p.n1168 vp_p.t128 756.008
R9132 vp_p.n1166 vp_p.t1292 756.008
R9133 vp_p.n1166 vp_p.t367 756.008
R9134 vp_p.n1164 vp_p.t889 756.008
R9135 vp_p.n1164 vp_p.t1454 756.008
R9136 vp_p.n1162 vp_p.t312 756.008
R9137 vp_p.n1162 vp_p.t884 756.008
R9138 vp_p.n1160 vp_p.t552 756.008
R9139 vp_p.n1160 vp_p.t1114 756.008
R9140 vp_p.n1158 vp_p.t132 756.008
R9141 vp_p.n1158 vp_p.t714 756.008
R9142 vp_p.n1156 vp_p.t379 756.008
R9143 vp_p.n1156 vp_p.t937 756.008
R9144 vp_p.n1154 vp_p.t1462 756.008
R9145 vp_p.n1154 vp_p.t538 756.008
R9146 vp_p.n1152 vp_p.t27 756.008
R9147 vp_p.n1152 vp_p.t601 756.008
R9148 vp_p.n1150 vp_p.t1125 756.008
R9149 vp_p.n1150 vp_p.t185 756.008
R9150 vp_p.n1148 vp_p.t722 756.008
R9151 vp_p.n1148 vp_p.t1278 756.008
R9152 vp_p.n1146 vp_p.t950 756.008
R9153 vp_p.n1146 vp_p.t6 756.008
R9154 vp_p.n1144 vp_p.t546 756.008
R9155 vp_p.n1144 vp_p.t1110 756.008
R9156 vp_p.n1142 vp_p.t1492 756.008
R9157 vp_p.n1142 vp_p.t568 756.008
R9158 vp_p.n1140 vp_p.t1097 756.008
R9159 vp_p.n1140 vp_p.t158 756.008
R9160 vp_p.n1138 vp_p.t692 756.008
R9161 vp_p.n1138 vp_p.t1251 756.008
R9162 vp_p.n1136 vp_p.t921 756.008
R9163 vp_p.n1136 vp_p.t1478 756.008
R9164 vp_p.n1134 vp_p.t517 756.008
R9165 vp_p.n1134 vp_p.t1085 756.008
R9166 vp_p.n1132 vp_p.t582 756.008
R9167 vp_p.n1132 vp_p.t1142 756.008
R9168 vp_p.n1130 vp_p.t168 756.008
R9169 vp_p.n1130 vp_p.t742 756.008
R9170 vp_p.n1128 vp_p.t412 756.008
R9171 vp_p.n1128 vp_p.t968 756.008
R9172 vp_p.n1126 vp_p.t1485 756.008
R9173 vp_p.n1126 vp_p.t563 756.008
R9174 vp_p.n1124 vp_p.t1091 756.008
R9175 vp_p.n1124 vp_p.t154 756.008
R9176 vp_p.n1122 vp_p.t1156 756.008
R9177 vp_p.n1122 vp_p.t220 756.008
R9178 vp_p.n1121 vp_p.t754 756.008
R9179 vp_p.n1121 vp_p.t1310 756.008
R9180 vp_p.n1417 vp_p.t749 756.008
R9181 vp_p.n1417 vp_p.t872 756.008
R9182 vp_p.n1415 vp_p.t341 756.008
R9183 vp_p.n1415 vp_p.t465 756.008
R9184 vp_p.n1413 vp_p.t571 756.008
R9185 vp_p.n1413 vp_p.t706 756.008
R9186 vp_p.n1411 vp_p.t160 756.008
R9187 vp_p.n1411 vp_p.t289 756.008
R9188 vp_p.n1409 vp_p.t226 756.008
R9189 vp_p.n1409 vp_p.t359 756.008
R9190 vp_p.n1407 vp_p.t1319 756.008
R9191 vp_p.n1407 vp_p.t1442 756.008
R9192 vp_p.n1405 vp_p.t912 756.008
R9193 vp_p.n1405 vp_p.t1038 756.008
R9194 vp_p.n1403 vp_p.t1144 756.008
R9195 vp_p.n1403 vp_p.t1272 756.008
R9196 vp_p.n1401 vp_p.t744 756.008
R9197 vp_p.n1401 vp_p.t865 756.008
R9198 vp_p.n1399 vp_p.t811 756.008
R9199 vp_p.n1399 vp_p.t929 756.008
R9200 vp_p.n1397 vp_p.t403 756.008
R9201 vp_p.n1397 vp_p.t530 756.008
R9202 vp_p.n1395 vp_p.t637 756.008
R9203 vp_p.n1395 vp_p.t766 756.008
R9204 vp_p.n1393 vp_p.t223 756.008
R9205 vp_p.n1393 vp_p.t354 756.008
R9206 vp_p.n1391 vp_p.t1312 756.008
R9207 vp_p.n1391 vp_p.t1433 756.008
R9208 vp_p.n1389 vp_p.t1379 756.008
R9209 vp_p.n1389 vp_p.t1498 756.008
R9210 vp_p.n1387 vp_p.t971 756.008
R9211 vp_p.n1387 vp_p.t1103 756.008
R9212 vp_p.n1385 vp_p.t994 756.008
R9213 vp_p.n1385 vp_p.t1117 756.008
R9214 vp_p.n1383 vp_p.t591 756.008
R9215 vp_p.n1383 vp_p.t717 756.008
R9216 vp_p.n1381 vp_p.t180 756.008
R9217 vp_p.n1381 vp_p.t302 756.008
R9218 vp_p.n1379 vp_p.t243 756.008
R9219 vp_p.n1379 vp_p.t371 756.008
R9220 vp_p.n1377 vp_p.t1336 756.008
R9221 vp_p.n1377 vp_p.t1457 756.008
R9222 vp_p.n1375 vp_p.t67 756.008
R9223 vp_p.n1375 vp_p.t191 756.008
R9224 vp_p.n1373 vp_p.t1165 756.008
R9225 vp_p.n1373 vp_p.t1280 756.008
R9226 vp_p.n1371 vp_p.t1395 756.008
R9227 vp_p.n1371 vp_p.t12 756.008
R9228 vp_p.n1369 vp_p.t826 756.008
R9229 vp_p.n1369 vp_p.t942 756.008
R9230 vp_p.n1367 vp_p.t423 756.008
R9231 vp_p.n1367 vp_p.t541 756.008
R9232 vp_p.n1365 vp_p.t656 756.008
R9233 vp_p.n1365 vp_p.t777 756.008
R9234 vp_p.n1363 vp_p.t242 756.008
R9235 vp_p.n1363 vp_p.t365 756.008
R9236 vp_p.n1361 vp_p.t484 756.008
R9237 vp_p.n1361 vp_p.t598 756.008
R9238 vp_p.n1359 vp_p.t1396 756.008
R9239 vp_p.n1359 vp_p.t13 756.008
R9240 vp_p.n1357 vp_p.t130 756.008
R9241 vp_p.n1357 vp_p.t255 756.008
R9242 vp_p.n1355 vp_p.t1223 756.008
R9243 vp_p.n1355 vp_p.t1342 756.008
R9244 vp_p.n1353 vp_p.t825 756.008
R9245 vp_p.n1353 vp_p.t935 756.008
R9246 vp_p.n1351 vp_p.t1058 756.008
R9247 vp_p.n1351 vp_p.t1172 756.008
R9248 vp_p.n1349 vp_p.t485 756.008
R9249 vp_p.n1349 vp_p.t599 756.008
R9250 vp_p.n1347 vp_p.t716 756.008
R9251 vp_p.n1347 vp_p.t838 756.008
R9252 vp_p.n1345 vp_p.t304 756.008
R9253 vp_p.n1345 vp_p.t427 756.008
R9254 vp_p.n1343 vp_p.t1394 756.008
R9255 vp_p.n1343 vp_p.t3 756.008
R9256 vp_p.n1341 vp_p.t127 756.008
R9257 vp_p.n1341 vp_p.t248 756.008
R9258 vp_p.n1339 vp_p.t1059 756.008
R9259 vp_p.n1339 vp_p.t1174 756.008
R9260 vp_p.n1337 vp_p.t689 756.008
R9261 vp_p.n1337 vp_p.t808 756.008
R9262 vp_p.n1335 vp_p.t275 756.008
R9263 vp_p.n1335 vp_p.t400 756.008
R9264 vp_p.n1333 vp_p.t515 756.008
R9265 vp_p.n1333 vp_p.t634 756.008
R9266 vp_p.n1331 vp_p.t99 756.008
R9267 vp_p.n1331 vp_p.t216 756.008
R9268 vp_p.n1329 vp_p.t1025 756.008
R9269 vp_p.n1329 vp_p.t1140 756.008
R9270 vp_p.n1327 vp_p.t1257 756.008
R9271 vp_p.n1327 vp_p.t1376 756.008
R9272 vp_p.n1325 vp_p.t854 756.008
R9273 vp_p.n1325 vp_p.t965 756.008
R9274 vp_p.n1323 vp_p.t1088 756.008
R9275 vp_p.n1323 vp_p.t1207 756.008
R9276 vp_p.n1321 vp_p.t686 756.008
R9277 vp_p.n1321 vp_p.t801 756.008
R9278 vp_p.n1319 vp_p.t747 756.008
R9279 vp_p.n1319 vp_p.t870 756.008
R9280 vp_p.n1317 vp_p.t339 756.008
R9281 vp_p.n1317 vp_p.t463 756.008
R9282 vp_p.n1315 vp_p.t1423 756.008
R9283 vp_p.n1315 vp_p.t37 756.008
R9284 vp_p.n1313 vp_p.t157 756.008
R9285 vp_p.n1313 vp_p.t284 756.008
R9286 vp_p.n1311 vp_p.t1250 756.008
R9287 vp_p.n1311 vp_p.t1367 756.008
R9288 vp_p.n1309 vp_p.t1317 756.008
R9289 vp_p.n1309 vp_p.t1441 756.008
R9290 vp_p.n1307 vp_p.t910 756.008
R9291 vp_p.n1307 vp_p.t1035 756.008
R9292 vp_p.n1305 vp_p.t511 756.008
R9293 vp_p.n1305 vp_p.t627 756.008
R9294 vp_p.n1303 vp_p.t741 756.008
R9295 vp_p.n1303 vp_p.t861 756.008
R9296 vp_p.n1301 vp_p.t334 756.008
R9297 vp_p.n1301 vp_p.t453 756.008
R9298 vp_p.n1299 vp_p.t399 756.008
R9299 vp_p.n1299 vp_p.t528 756.008
R9300 vp_p.n1297 vp_p.t1477 756.008
R9301 vp_p.n1297 vp_p.t106 756.008
R9302 vp_p.n1295 vp_p.t219 756.008
R9303 vp_p.n1295 vp_p.t349 756.008
R9304 vp_p.n1293 vp_p.t1308 756.008
R9305 vp_p.n1293 vp_p.t1428 756.008
R9306 vp_p.n1291 vp_p.t909 756.008
R9307 vp_p.n1291 vp_p.t1027 756.008
R9308 vp_p.n1289 vp_p.t368 756.008
R9309 vp_p.n1289 vp_p.t498 756.008
R9310 vp_p.n1287 vp_p.t1455 756.008
R9311 vp_p.n1287 vp_p.t75 756.008
R9312 vp_p.n1285 vp_p.t186 756.008
R9313 vp_p.n1285 vp_p.t320 756.008
R9314 vp_p.n1283 vp_p.t1279 756.008
R9315 vp_p.n1283 vp_p.t1402 756.008
R9316 vp_p.n1281 vp_p.t880 756.008
R9317 vp_p.n1281 vp_p.t996 756.008
R9318 vp_p.n1279 vp_p.t939 756.008
R9319 vp_p.n1279 vp_p.t1071 756.008
R9320 vp_p.n1277 vp_p.t539 756.008
R9321 vp_p.n1277 vp_p.t661 756.008
R9322 vp_p.n1275 vp_p.t772 756.008
R9323 vp_p.n1275 vp_p.t895 756.008
R9324 vp_p.n1273 vp_p.t363 756.008
R9325 vp_p.n1273 vp_p.t488 756.008
R9326 vp_p.n1271 vp_p.t593 756.008
R9327 vp_p.n1271 vp_p.t725 756.008
R9328 vp_p.n1270 vp_p.t8 756.008
R9329 vp_p.n1270 vp_p.t139 756.008
R9330 vp_p.n670 vp_p.t875 706.013
R9331 vp_p.n0 vp_p.t639 706.013
R9332 vp_p.n1419 vp_p.t1430 706.013
R9333 vp_p.n749 vp_p.t1245 705.989
R9334 vp_p.n743 vp_p.t95 704.872
R9335 vp_p.n742 vp_p.t1190 704.872
R9336 vp_p.n741 vp_p.t1420 704.872
R9337 vp_p.n740 vp_p.t1016 704.872
R9338 vp_p.n739 vp_p.t1084 704.872
R9339 vp_p.n738 vp_p.t683 704.872
R9340 vp_p.n737 vp_p.t264 704.872
R9341 vp_p.n736 vp_p.t509 704.872
R9342 vp_p.n735 vp_p.t89 704.872
R9343 vp_p.n734 vp_p.t153 704.872
R9344 vp_p.n733 vp_p.t1248 704.872
R9345 vp_p.n732 vp_p.t1475 704.872
R9346 vp_p.n731 vp_p.t1082 704.872
R9347 vp_p.n730 vp_p.t677 704.872
R9348 vp_p.n729 vp_p.t738 704.872
R9349 vp_p.n728 vp_p.t330 704.872
R9350 vp_p.n727 vp_p.t355 704.872
R9351 vp_p.n726 vp_p.t1434 704.872
R9352 vp_p.n725 vp_p.t1029 704.872
R9353 vp_p.n724 vp_p.t1104 704.872
R9354 vp_p.n723 vp_p.t698 704.872
R9355 vp_p.n722 vp_p.t925 704.872
R9356 vp_p.n721 vp_p.t519 704.872
R9357 vp_p.n720 vp_p.t759 704.872
R9358 vp_p.n719 vp_p.t172 704.872
R9359 vp_p.n718 vp_p.t1261 704.872
R9360 vp_p.n717 vp_p.t1491 704.872
R9361 vp_p.n716 vp_p.t1093 704.872
R9362 vp_p.n715 vp_p.t1327 704.872
R9363 vp_p.n714 vp_p.t760 704.872
R9364 vp_p.n713 vp_p.t988 704.872
R9365 vp_p.n712 vp_p.t580 704.872
R9366 vp_p.n711 vp_p.t164 704.872
R9367 vp_p.n710 vp_p.t409 704.872
R9368 vp_p.n709 vp_p.t1328 704.872
R9369 vp_p.n708 vp_p.t57 704.872
R9370 vp_p.n707 vp_p.t1152 704.872
R9371 vp_p.n706 vp_p.t751 704.872
R9372 vp_p.n705 vp_p.t980 704.872
R9373 vp_p.n704 vp_p.t410 704.872
R9374 vp_p.n703 vp_p.t26 704.872
R9375 vp_p.n702 vp_p.t1124 704.872
R9376 vp_p.n701 vp_p.t1357 704.872
R9377 vp_p.n700 vp_p.t948 704.872
R9378 vp_p.n699 vp_p.t380 704.872
R9379 vp_p.n698 vp_p.t616 704.872
R9380 vp_p.n697 vp_p.t196 704.872
R9381 vp_p.n696 vp_p.t442 704.872
R9382 vp_p.n695 vp_p.t17 704.872
R9383 vp_p.n694 vp_p.t93 704.872
R9384 vp_p.n693 vp_p.t1189 704.872
R9385 vp_p.n692 vp_p.t782 704.872
R9386 vp_p.n691 vp_p.t1014 704.872
R9387 vp_p.n690 vp_p.t608 704.872
R9388 vp_p.n689 vp_p.t682 704.872
R9389 vp_p.n688 vp_p.t262 704.872
R9390 vp_p.n687 vp_p.t1348 704.872
R9391 vp_p.n686 vp_p.t87 704.872
R9392 vp_p.n685 vp_p.t1182 704.872
R9393 vp_p.n684 vp_p.t1247 704.872
R9394 vp_p.n683 vp_p.t845 704.872
R9395 vp_p.n682 vp_p.t1080 704.872
R9396 vp_p.n681 vp_p.t675 704.872
R9397 vp_p.n680 vp_p.t256 704.872
R9398 vp_p.n679 vp_p.t1218 704.872
R9399 vp_p.n678 vp_p.t815 704.872
R9400 vp_p.n677 vp_p.t1051 704.872
R9401 vp_p.n676 vp_p.t644 704.872
R9402 vp_p.n675 vp_p.t227 704.872
R9403 vp_p.n674 vp_p.t298 704.872
R9404 vp_p.n673 vp_p.t1383 704.872
R9405 vp_p.n672 vp_p.t119 704.872
R9406 vp_p.n671 vp_p.t1212 704.872
R9407 vp_p.n670 vp_p.t1445 704.872
R9408 vp_p.n0 vp_p.t1044 704.872
R9409 vp_p.n1 vp_p.t972 704.872
R9410 vp_p.n2 vp_p.t1380 704.872
R9411 vp_p.n3 vp_p.t293 704.872
R9412 vp_p.n4 vp_p.t46 704.872
R9413 vp_p.n5 vp_p.t469 704.872
R9414 vp_p.n6 vp_p.t404 704.872
R9415 vp_p.n7 vp_p.t812 704.872
R9416 vp_p.n8 vp_p.t572 704.872
R9417 vp_p.n9 vp_p.t976 704.872
R9418 vp_p.n10 vp_p.t1384 704.872
R9419 vp_p.n11 vp_p.t436 704.872
R9420 vp_p.n12 vp_p.t840 704.872
R9421 vp_p.n13 vp_p.t604 704.872
R9422 vp_p.n14 vp_p.t1009 704.872
R9423 vp_p.n15 vp_p.t1414 704.872
R9424 vp_p.n16 vp_p.t1346 704.872
R9425 vp_p.n17 vp_p.t257 704.872
R9426 vp_p.n18 vp_p.t16 704.872
R9427 vp_p.n19 vp_p.t439 704.872
R9428 vp_p.n20 vp_p.t194 704.872
R9429 vp_p.n21 vp_p.t779 704.872
R9430 vp_p.n22 vp_p.t1183 704.872
R9431 vp_p.n23 vp_p.t945 704.872
R9432 vp_p.n24 vp_p.t1349 704.872
R9433 vp_p.n25 vp_p.t1120 704.872
R9434 vp_p.n26 vp_p.t193 704.872
R9435 vp_p.n27 vp_p.t1460 704.872
R9436 vp_p.n28 vp_p.t375 704.872
R9437 vp_p.n29 vp_p.t784 704.872
R9438 vp_p.n30 vp_p.t548 704.872
R9439 vp_p.n31 vp_p.t1119 704.872
R9440 vp_p.n32 vp_p.t887 704.872
R9441 vp_p.n33 vp_p.t1288 704.872
R9442 vp_p.n34 vp_p.t197 704.872
R9443 vp_p.n35 vp_p.t575 704.872
R9444 vp_p.n36 vp_p.t1147 704.872
R9445 vp_p.n37 vp_p.t915 704.872
R9446 vp_p.n38 vp_p.t1321 704.872
R9447 vp_p.n39 vp_p.t1090 704.872
R9448 vp_p.n40 vp_p.t1484 704.872
R9449 vp_p.n41 vp_p.t574 704.872
R9450 vp_p.n42 vp_p.t343 704.872
R9451 vp_p.n43 vp_p.t752 704.872
R9452 vp_p.n44 vp_p.t516 704.872
R9453 vp_p.n45 vp_p.t920 704.872
R9454 vp_p.n46 vp_p.t856 704.872
R9455 vp_p.n47 vp_p.t1258 704.872
R9456 vp_p.n48 vp_p.t165 704.872
R9457 vp_p.n49 vp_p.t1427 704.872
R9458 vp_p.n50 vp_p.t345 704.872
R9459 vp_p.n51 vp_p.t277 704.872
R9460 vp_p.n52 vp_p.t691 704.872
R9461 vp_p.n53 vp_p.t1096 704.872
R9462 vp_p.n54 vp_p.t857 704.872
R9463 vp_p.n55 vp_p.t1263 704.872
R9464 vp_p.n56 vp_p.t1199 704.872
R9465 vp_p.n57 vp_p.t102 704.872
R9466 vp_p.n58 vp_p.t85 704.872
R9467 vp_p.n59 vp_p.t505 704.872
R9468 vp_p.n60 vp_p.t907 704.872
R9469 vp_p.n61 vp_p.t843 704.872
R9470 vp_p.n62 vp_p.t1243 704.872
R9471 vp_p.n63 vp_p.t1012 704.872
R9472 vp_p.n64 vp_p.t1416 704.872
R9473 vp_p.n65 vp_p.t331 704.872
R9474 vp_p.n66 vp_p.t259 704.872
R9475 vp_p.n67 vp_p.t679 704.872
R9476 vp_p.n68 vp_p.t441 704.872
R9477 vp_p.n69 vp_p.t847 704.872
R9478 vp_p.n70 vp_p.t611 704.872
R9479 vp_p.n71 vp_p.t1186 704.872
R9480 vp_p.n72 vp_p.t90 704.872
R9481 vp_p.n73 vp_p.t1353 704.872
R9482 vp_p.n749 vp_p.t328 704.872
R9483 vp_p.n750 vp_p.t86 704.872
R9484 vp_p.n751 vp_p.t506 704.872
R9485 vp_p.n752 vp_p.t261 704.872
R9486 vp_p.n753 vp_p.t680 704.872
R9487 vp_p.n754 vp_p.t607 704.872
R9488 vp_p.n755 vp_p.t1013 704.872
R9489 vp_p.n756 vp_p.t1417 704.872
R9490 vp_p.n757 vp_p.t1187 704.872
R9491 vp_p.n758 vp_p.t92 704.872
R9492 vp_p.n759 vp_p.t640 704.872
R9493 vp_p.n760 vp_p.t1047 704.872
R9494 vp_p.n761 vp_p.t1447 704.872
R9495 vp_p.n762 vp_p.t1214 704.872
R9496 vp_p.n763 vp_p.t121 704.872
R9497 vp_p.n764 vp_p.t48 704.872
R9498 vp_p.n765 vp_p.t470 704.872
R9499 vp_p.n766 vp_p.t229 704.872
R9500 vp_p.n767 vp_p.t648 704.872
R9501 vp_p.n768 vp_p.t1054 704.872
R9502 vp_p.n769 vp_p.t977 704.872
R9503 vp_p.n770 vp_p.t1385 704.872
R9504 vp_p.n771 vp_p.t1151 704.872
R9505 vp_p.n772 vp_p.t55 704.872
R9506 vp_p.n773 vp_p.t476 704.872
R9507 vp_p.n774 vp_p.t408 704.872
R9508 vp_p.n775 vp_p.t817 704.872
R9509 vp_p.n776 vp_p.t579 704.872
R9510 vp_p.n777 vp_p.t986 704.872
R9511 vp_p.n778 vp_p.t758 704.872
R9512 vp_p.n779 vp_p.t1326 704.872
R9513 vp_p.n780 vp_p.t236 704.872
R9514 vp_p.n781 vp_p.t1489 704.872
R9515 vp_p.n782 vp_p.t417 704.872
R9516 vp_p.n783 vp_p.t787 704.872
R9517 vp_p.n784 vp_p.t1351 704.872
R9518 vp_p.n785 vp_p.t1121 704.872
R9519 vp_p.n786 vp_p.t21 704.872
R9520 vp_p.n787 vp_p.t444 704.872
R9521 vp_p.n788 vp_p.t201 704.872
R9522 vp_p.n789 vp_p.t785 704.872
R9523 vp_p.n790 vp_p.t549 704.872
R9524 vp_p.n791 vp_p.t953 704.872
R9525 vp_p.n792 vp_p.t1359 704.872
R9526 vp_p.n793 vp_p.t1129 704.872
R9527 vp_p.n794 vp_p.t200 704.872
R9528 vp_p.n795 vp_p.t1465 704.872
R9529 vp_p.n796 vp_p.t384 704.872
R9530 vp_p.n797 vp_p.t136 704.872
R9531 vp_p.n798 vp_p.t555 704.872
R9532 vp_p.n799 vp_p.t1128 704.872
R9533 vp_p.n800 vp_p.t894 704.872
R9534 vp_p.n801 vp_p.t1295 704.872
R9535 vp_p.n802 vp_p.t1069 704.872
R9536 vp_p.n803 vp_p.t1469 704.872
R9537 vp_p.n804 vp_p.t1399 704.872
R9538 vp_p.n805 vp_p.t318 704.872
R9539 vp_p.n806 vp_p.t729 704.872
R9540 vp_p.n807 vp_p.t712 704.872
R9541 vp_p.n808 vp_p.t1109 704.872
R9542 vp_p.n809 vp_p.t1050 704.872
R9543 vp_p.n810 vp_p.t1449 704.872
R9544 vp_p.n811 vp_p.t361 704.872
R9545 vp_p.n812 vp_p.t123 704.872
R9546 vp_p.n813 vp_p.t537 704.872
R9547 vp_p.n814 vp_p.t473 704.872
R9548 vp_p.n815 vp_p.t878 704.872
R9549 vp_p.n816 vp_p.t649 704.872
R9550 vp_p.n817 vp_p.t1055 704.872
R9551 vp_p.n818 vp_p.t1452 704.872
R9552 vp_p.n819 vp_p.t1388 704.872
R9553 vp_p.n820 vp_p.t301 704.872
R9554 vp_p.n821 vp_p.t58 704.872
R9555 vp_p.n822 vp_p.t478 704.872
R9556 vp_p.n1419 vp_p.t353 704.872
R9557 vp_p.n1420 vp_p.t278 704.872
R9558 vp_p.n1421 vp_p.t695 704.872
R9559 vp_p.n1422 vp_p.t1102 704.872
R9560 vp_p.n1423 vp_p.t863 704.872
R9561 vp_p.n1424 vp_p.t1271 704.872
R9562 vp_p.n1425 vp_p.t1201 704.872
R9563 vp_p.n1426 vp_p.t110 704.872
R9564 vp_p.n1427 vp_p.t1369 704.872
R9565 vp_p.n1428 vp_p.t286 704.872
R9566 vp_p.n1429 vp_p.t705 704.872
R9567 vp_p.n1430 vp_p.t1226 704.872
R9568 vp_p.n1431 vp_p.t137 704.872
R9569 vp_p.n1432 vp_p.t1400 704.872
R9570 vp_p.n1433 vp_p.t315 704.872
R9571 vp_p.n1434 vp_p.t732 704.872
R9572 vp_p.n1435 vp_p.t659 704.872
R9573 vp_p.n1436 vp_p.t1067 704.872
R9574 vp_p.n1437 vp_p.t831 704.872
R9575 vp_p.n1438 vp_p.t1238 704.872
R9576 vp_p.n1439 vp_p.t1002 704.872
R9577 vp_p.n1440 vp_p.t73 704.872
R9578 vp_p.n1441 vp_p.t497 704.872
R9579 vp_p.n1442 vp_p.t250 704.872
R9580 vp_p.n1443 vp_p.t669 704.872
R9581 vp_p.n1444 vp_p.t431 704.872
R9582 vp_p.n1445 vp_p.t1001 704.872
R9583 vp_p.n1446 vp_p.t769 704.872
R9584 vp_p.n1447 vp_p.t1175 704.872
R9585 vp_p.n1448 vp_p.t81 704.872
R9586 vp_p.n1449 vp_p.t1344 704.872
R9587 vp_p.n1450 vp_p.t430 704.872
R9588 vp_p.n1451 vp_p.t182 704.872
R9589 vp_p.n1452 vp_p.t602 704.872
R9590 vp_p.n1453 vp_p.t1006 704.872
R9591 vp_p.n1454 vp_p.t1375 704.872
R9592 vp_p.n1455 vp_p.t460 704.872
R9593 vp_p.n1456 vp_p.t214 704.872
R9594 vp_p.n1457 vp_p.t633 704.872
R9595 vp_p.n1458 vp_p.t396 704.872
R9596 vp_p.n1459 vp_p.t807 704.872
R9597 vp_p.n1460 vp_p.t1373 704.872
R9598 vp_p.n1461 vp_p.t1138 704.872
R9599 vp_p.n1462 vp_p.t43 704.872
R9600 vp_p.n1463 vp_p.t1314 704.872
R9601 vp_p.n1464 vp_p.t225 704.872
R9602 vp_p.n1465 vp_p.t155 704.872
R9603 vp_p.n1466 vp_p.t566 704.872
R9604 vp_p.n1467 vp_p.t974 704.872
R9605 vp_p.n1468 vp_p.t745 704.872
R9606 vp_p.n1469 vp_p.t1146 704.872
R9607 vp_p.n1470 vp_p.t1086 704.872
R9608 vp_p.n1471 vp_p.t1480 704.872
R9609 vp_p.n1472 vp_p.t405 704.872
R9610 vp_p.n1473 vp_p.t161 704.872
R9611 vp_p.n1474 vp_p.t573 704.872
R9612 vp_p.n1475 vp_p.t513 704.872
R9613 vp_p.n1476 vp_p.t913 704.872
R9614 vp_p.n1477 vp_p.t897 704.872
R9615 vp_p.n1478 vp_p.t1299 704.872
R9616 vp_p.n1479 vp_p.t210 704.872
R9617 vp_p.n1480 vp_p.t141 704.872
R9618 vp_p.n1481 vp_p.t557 704.872
R9619 vp_p.n1482 vp_p.t321 704.872
R9620 vp_p.n1483 vp_p.t733 704.872
R9621 vp_p.n1484 vp_p.t1135 704.872
R9622 vp_p.n1485 vp_p.t1073 704.872
R9623 vp_p.n1486 vp_p.t1472 704.872
R9624 vp_p.n1487 vp_p.t1240 704.872
R9625 vp_p.n1488 vp_p.t148 704.872
R9626 vp_p.n1489 vp_p.t1410 704.872
R9627 vp_p.n1490 vp_p.t500 704.872
R9628 vp_p.n1491 vp_p.t905 704.872
R9629 vp_p.n1492 vp_p.t672 704.872
R9630 vp_p.n1493 vp_p.n1492 1.225
R9631 vp_p.n671 vp_p.n670 1.141
R9632 vp_p.n672 vp_p.n671 1.141
R9633 vp_p.n673 vp_p.n672 1.141
R9634 vp_p.n674 vp_p.n673 1.141
R9635 vp_p.n675 vp_p.n674 1.141
R9636 vp_p.n676 vp_p.n675 1.141
R9637 vp_p.n677 vp_p.n676 1.141
R9638 vp_p.n678 vp_p.n677 1.141
R9639 vp_p.n679 vp_p.n678 1.141
R9640 vp_p.n680 vp_p.n679 1.141
R9641 vp_p.n681 vp_p.n680 1.141
R9642 vp_p.n682 vp_p.n681 1.141
R9643 vp_p.n683 vp_p.n682 1.141
R9644 vp_p.n684 vp_p.n683 1.141
R9645 vp_p.n685 vp_p.n684 1.141
R9646 vp_p.n686 vp_p.n685 1.141
R9647 vp_p.n687 vp_p.n686 1.141
R9648 vp_p.n688 vp_p.n687 1.141
R9649 vp_p.n689 vp_p.n688 1.141
R9650 vp_p.n690 vp_p.n689 1.141
R9651 vp_p.n691 vp_p.n690 1.141
R9652 vp_p.n692 vp_p.n691 1.141
R9653 vp_p.n693 vp_p.n692 1.141
R9654 vp_p.n694 vp_p.n693 1.141
R9655 vp_p.n695 vp_p.n694 1.141
R9656 vp_p.n696 vp_p.n695 1.141
R9657 vp_p.n697 vp_p.n696 1.141
R9658 vp_p.n698 vp_p.n697 1.141
R9659 vp_p.n699 vp_p.n698 1.141
R9660 vp_p.n700 vp_p.n699 1.141
R9661 vp_p.n701 vp_p.n700 1.141
R9662 vp_p.n702 vp_p.n701 1.141
R9663 vp_p.n703 vp_p.n702 1.141
R9664 vp_p.n704 vp_p.n703 1.141
R9665 vp_p.n705 vp_p.n704 1.141
R9666 vp_p.n706 vp_p.n705 1.141
R9667 vp_p.n707 vp_p.n706 1.141
R9668 vp_p.n708 vp_p.n707 1.141
R9669 vp_p.n709 vp_p.n708 1.141
R9670 vp_p.n710 vp_p.n709 1.141
R9671 vp_p.n711 vp_p.n710 1.141
R9672 vp_p.n712 vp_p.n711 1.141
R9673 vp_p.n713 vp_p.n712 1.141
R9674 vp_p.n714 vp_p.n713 1.141
R9675 vp_p.n715 vp_p.n714 1.141
R9676 vp_p.n716 vp_p.n715 1.141
R9677 vp_p.n717 vp_p.n716 1.141
R9678 vp_p.n718 vp_p.n717 1.141
R9679 vp_p.n719 vp_p.n718 1.141
R9680 vp_p.n720 vp_p.n719 1.141
R9681 vp_p.n721 vp_p.n720 1.141
R9682 vp_p.n722 vp_p.n721 1.141
R9683 vp_p.n723 vp_p.n722 1.141
R9684 vp_p.n724 vp_p.n723 1.141
R9685 vp_p.n725 vp_p.n724 1.141
R9686 vp_p.n726 vp_p.n725 1.141
R9687 vp_p.n727 vp_p.n726 1.141
R9688 vp_p.n728 vp_p.n727 1.141
R9689 vp_p.n729 vp_p.n728 1.141
R9690 vp_p.n730 vp_p.n729 1.141
R9691 vp_p.n731 vp_p.n730 1.141
R9692 vp_p.n732 vp_p.n731 1.141
R9693 vp_p.n733 vp_p.n732 1.141
R9694 vp_p.n734 vp_p.n733 1.141
R9695 vp_p.n735 vp_p.n734 1.141
R9696 vp_p.n736 vp_p.n735 1.141
R9697 vp_p.n737 vp_p.n736 1.141
R9698 vp_p.n738 vp_p.n737 1.141
R9699 vp_p.n739 vp_p.n738 1.141
R9700 vp_p.n740 vp_p.n739 1.141
R9701 vp_p.n741 vp_p.n740 1.141
R9702 vp_p.n742 vp_p.n741 1.141
R9703 vp_p.n743 vp_p.n742 1.141
R9704 vp_p.n1 vp_p.n0 1.141
R9705 vp_p.n2 vp_p.n1 1.141
R9706 vp_p.n3 vp_p.n2 1.141
R9707 vp_p.n4 vp_p.n3 1.141
R9708 vp_p.n5 vp_p.n4 1.141
R9709 vp_p.n6 vp_p.n5 1.141
R9710 vp_p.n7 vp_p.n6 1.141
R9711 vp_p.n8 vp_p.n7 1.141
R9712 vp_p.n9 vp_p.n8 1.141
R9713 vp_p.n10 vp_p.n9 1.141
R9714 vp_p.n11 vp_p.n10 1.141
R9715 vp_p.n12 vp_p.n11 1.141
R9716 vp_p.n13 vp_p.n12 1.141
R9717 vp_p.n14 vp_p.n13 1.141
R9718 vp_p.n15 vp_p.n14 1.141
R9719 vp_p.n16 vp_p.n15 1.141
R9720 vp_p.n17 vp_p.n16 1.141
R9721 vp_p.n18 vp_p.n17 1.141
R9722 vp_p.n19 vp_p.n18 1.141
R9723 vp_p.n20 vp_p.n19 1.141
R9724 vp_p.n21 vp_p.n20 1.141
R9725 vp_p.n22 vp_p.n21 1.141
R9726 vp_p.n23 vp_p.n22 1.141
R9727 vp_p.n24 vp_p.n23 1.141
R9728 vp_p.n25 vp_p.n24 1.141
R9729 vp_p.n26 vp_p.n25 1.141
R9730 vp_p.n27 vp_p.n26 1.141
R9731 vp_p.n28 vp_p.n27 1.141
R9732 vp_p.n29 vp_p.n28 1.141
R9733 vp_p.n30 vp_p.n29 1.141
R9734 vp_p.n31 vp_p.n30 1.141
R9735 vp_p.n32 vp_p.n31 1.141
R9736 vp_p.n33 vp_p.n32 1.141
R9737 vp_p.n34 vp_p.n33 1.141
R9738 vp_p.n35 vp_p.n34 1.141
R9739 vp_p.n36 vp_p.n35 1.141
R9740 vp_p.n37 vp_p.n36 1.141
R9741 vp_p.n38 vp_p.n37 1.141
R9742 vp_p.n39 vp_p.n38 1.141
R9743 vp_p.n40 vp_p.n39 1.141
R9744 vp_p.n41 vp_p.n40 1.141
R9745 vp_p.n42 vp_p.n41 1.141
R9746 vp_p.n43 vp_p.n42 1.141
R9747 vp_p.n44 vp_p.n43 1.141
R9748 vp_p.n45 vp_p.n44 1.141
R9749 vp_p.n46 vp_p.n45 1.141
R9750 vp_p.n47 vp_p.n46 1.141
R9751 vp_p.n48 vp_p.n47 1.141
R9752 vp_p.n49 vp_p.n48 1.141
R9753 vp_p.n50 vp_p.n49 1.141
R9754 vp_p.n51 vp_p.n50 1.141
R9755 vp_p.n52 vp_p.n51 1.141
R9756 vp_p.n53 vp_p.n52 1.141
R9757 vp_p.n54 vp_p.n53 1.141
R9758 vp_p.n55 vp_p.n54 1.141
R9759 vp_p.n56 vp_p.n55 1.141
R9760 vp_p.n57 vp_p.n56 1.141
R9761 vp_p.n58 vp_p.n57 1.141
R9762 vp_p.n59 vp_p.n58 1.141
R9763 vp_p.n60 vp_p.n59 1.141
R9764 vp_p.n61 vp_p.n60 1.141
R9765 vp_p.n62 vp_p.n61 1.141
R9766 vp_p.n63 vp_p.n62 1.141
R9767 vp_p.n64 vp_p.n63 1.141
R9768 vp_p.n65 vp_p.n64 1.141
R9769 vp_p.n66 vp_p.n65 1.141
R9770 vp_p.n67 vp_p.n66 1.141
R9771 vp_p.n68 vp_p.n67 1.141
R9772 vp_p.n69 vp_p.n68 1.141
R9773 vp_p.n70 vp_p.n69 1.141
R9774 vp_p.n71 vp_p.n70 1.141
R9775 vp_p.n72 vp_p.n71 1.141
R9776 vp_p.n73 vp_p.n72 1.141
R9777 vp_p.n1420 vp_p.n1419 1.141
R9778 vp_p.n1421 vp_p.n1420 1.141
R9779 vp_p.n1422 vp_p.n1421 1.141
R9780 vp_p.n1423 vp_p.n1422 1.141
R9781 vp_p.n1424 vp_p.n1423 1.141
R9782 vp_p.n1425 vp_p.n1424 1.141
R9783 vp_p.n1426 vp_p.n1425 1.141
R9784 vp_p.n1427 vp_p.n1426 1.141
R9785 vp_p.n1428 vp_p.n1427 1.141
R9786 vp_p.n1429 vp_p.n1428 1.141
R9787 vp_p.n1430 vp_p.n1429 1.141
R9788 vp_p.n1431 vp_p.n1430 1.141
R9789 vp_p.n1432 vp_p.n1431 1.141
R9790 vp_p.n1433 vp_p.n1432 1.141
R9791 vp_p.n1434 vp_p.n1433 1.141
R9792 vp_p.n1435 vp_p.n1434 1.141
R9793 vp_p.n1436 vp_p.n1435 1.141
R9794 vp_p.n1437 vp_p.n1436 1.141
R9795 vp_p.n1438 vp_p.n1437 1.141
R9796 vp_p.n1439 vp_p.n1438 1.141
R9797 vp_p.n1440 vp_p.n1439 1.141
R9798 vp_p.n1441 vp_p.n1440 1.141
R9799 vp_p.n1442 vp_p.n1441 1.141
R9800 vp_p.n1443 vp_p.n1442 1.141
R9801 vp_p.n1444 vp_p.n1443 1.141
R9802 vp_p.n1445 vp_p.n1444 1.141
R9803 vp_p.n1446 vp_p.n1445 1.141
R9804 vp_p.n1447 vp_p.n1446 1.141
R9805 vp_p.n1448 vp_p.n1447 1.141
R9806 vp_p.n1449 vp_p.n1448 1.141
R9807 vp_p.n1450 vp_p.n1449 1.141
R9808 vp_p.n1451 vp_p.n1450 1.141
R9809 vp_p.n1452 vp_p.n1451 1.141
R9810 vp_p.n1453 vp_p.n1452 1.141
R9811 vp_p.n1454 vp_p.n1453 1.141
R9812 vp_p.n1455 vp_p.n1454 1.141
R9813 vp_p.n1456 vp_p.n1455 1.141
R9814 vp_p.n1457 vp_p.n1456 1.141
R9815 vp_p.n1458 vp_p.n1457 1.141
R9816 vp_p.n1459 vp_p.n1458 1.141
R9817 vp_p.n1460 vp_p.n1459 1.141
R9818 vp_p.n1461 vp_p.n1460 1.141
R9819 vp_p.n1462 vp_p.n1461 1.141
R9820 vp_p.n1463 vp_p.n1462 1.141
R9821 vp_p.n1464 vp_p.n1463 1.141
R9822 vp_p.n1465 vp_p.n1464 1.141
R9823 vp_p.n1466 vp_p.n1465 1.141
R9824 vp_p.n1467 vp_p.n1466 1.141
R9825 vp_p.n1468 vp_p.n1467 1.141
R9826 vp_p.n1469 vp_p.n1468 1.141
R9827 vp_p.n1470 vp_p.n1469 1.141
R9828 vp_p.n1471 vp_p.n1470 1.141
R9829 vp_p.n1472 vp_p.n1471 1.141
R9830 vp_p.n1473 vp_p.n1472 1.141
R9831 vp_p.n1474 vp_p.n1473 1.141
R9832 vp_p.n1475 vp_p.n1474 1.141
R9833 vp_p.n1476 vp_p.n1475 1.141
R9834 vp_p.n1477 vp_p.n1476 1.141
R9835 vp_p.n1478 vp_p.n1477 1.141
R9836 vp_p.n1479 vp_p.n1478 1.141
R9837 vp_p.n1480 vp_p.n1479 1.141
R9838 vp_p.n1481 vp_p.n1480 1.141
R9839 vp_p.n1482 vp_p.n1481 1.141
R9840 vp_p.n1483 vp_p.n1482 1.141
R9841 vp_p.n1484 vp_p.n1483 1.141
R9842 vp_p.n1485 vp_p.n1484 1.141
R9843 vp_p.n1486 vp_p.n1485 1.141
R9844 vp_p.n1487 vp_p.n1486 1.141
R9845 vp_p.n1488 vp_p.n1487 1.141
R9846 vp_p.n1489 vp_p.n1488 1.141
R9847 vp_p.n1490 vp_p.n1489 1.141
R9848 vp_p.n1491 vp_p.n1490 1.141
R9849 vp_p.n1492 vp_p.n1491 1.141
R9850 vp_p.n750 vp_p.n749 1.117
R9851 vp_p.n751 vp_p.n750 1.117
R9852 vp_p.n752 vp_p.n751 1.117
R9853 vp_p.n753 vp_p.n752 1.117
R9854 vp_p.n754 vp_p.n753 1.117
R9855 vp_p.n755 vp_p.n754 1.117
R9856 vp_p.n756 vp_p.n755 1.117
R9857 vp_p.n757 vp_p.n756 1.117
R9858 vp_p.n758 vp_p.n757 1.117
R9859 vp_p.n759 vp_p.n758 1.117
R9860 vp_p.n760 vp_p.n759 1.117
R9861 vp_p.n761 vp_p.n760 1.117
R9862 vp_p.n762 vp_p.n761 1.117
R9863 vp_p.n763 vp_p.n762 1.117
R9864 vp_p.n764 vp_p.n763 1.117
R9865 vp_p.n765 vp_p.n764 1.117
R9866 vp_p.n766 vp_p.n765 1.117
R9867 vp_p.n767 vp_p.n766 1.117
R9868 vp_p.n768 vp_p.n767 1.117
R9869 vp_p.n769 vp_p.n768 1.117
R9870 vp_p.n770 vp_p.n769 1.117
R9871 vp_p.n771 vp_p.n770 1.117
R9872 vp_p.n772 vp_p.n771 1.117
R9873 vp_p.n773 vp_p.n772 1.117
R9874 vp_p.n774 vp_p.n773 1.117
R9875 vp_p.n775 vp_p.n774 1.117
R9876 vp_p.n776 vp_p.n775 1.117
R9877 vp_p.n777 vp_p.n776 1.117
R9878 vp_p.n778 vp_p.n777 1.117
R9879 vp_p.n779 vp_p.n778 1.117
R9880 vp_p.n780 vp_p.n779 1.117
R9881 vp_p.n781 vp_p.n780 1.117
R9882 vp_p.n782 vp_p.n781 1.117
R9883 vp_p.n783 vp_p.n782 1.117
R9884 vp_p.n784 vp_p.n783 1.117
R9885 vp_p.n785 vp_p.n784 1.117
R9886 vp_p.n786 vp_p.n785 1.117
R9887 vp_p.n787 vp_p.n786 1.117
R9888 vp_p.n788 vp_p.n787 1.117
R9889 vp_p.n789 vp_p.n788 1.117
R9890 vp_p.n790 vp_p.n789 1.117
R9891 vp_p.n791 vp_p.n790 1.117
R9892 vp_p.n792 vp_p.n791 1.117
R9893 vp_p.n793 vp_p.n792 1.117
R9894 vp_p.n794 vp_p.n793 1.117
R9895 vp_p.n795 vp_p.n794 1.117
R9896 vp_p.n796 vp_p.n795 1.117
R9897 vp_p.n797 vp_p.n796 1.117
R9898 vp_p.n798 vp_p.n797 1.117
R9899 vp_p.n799 vp_p.n798 1.117
R9900 vp_p.n800 vp_p.n799 1.117
R9901 vp_p.n801 vp_p.n800 1.117
R9902 vp_p.n802 vp_p.n801 1.117
R9903 vp_p.n803 vp_p.n802 1.117
R9904 vp_p.n804 vp_p.n803 1.117
R9905 vp_p.n805 vp_p.n804 1.117
R9906 vp_p.n806 vp_p.n805 1.117
R9907 vp_p.n807 vp_p.n806 1.117
R9908 vp_p.n808 vp_p.n807 1.117
R9909 vp_p.n809 vp_p.n808 1.117
R9910 vp_p.n810 vp_p.n809 1.117
R9911 vp_p.n811 vp_p.n810 1.117
R9912 vp_p.n812 vp_p.n811 1.117
R9913 vp_p.n813 vp_p.n812 1.117
R9914 vp_p.n814 vp_p.n813 1.117
R9915 vp_p.n815 vp_p.n814 1.117
R9916 vp_p.n816 vp_p.n815 1.117
R9917 vp_p.n817 vp_p.n816 1.117
R9918 vp_p.n818 vp_p.n817 1.117
R9919 vp_p.n819 vp_p.n818 1.117
R9920 vp_p.n820 vp_p.n819 1.117
R9921 vp_p.n821 vp_p.n820 1.117
R9922 vp_p.n822 vp_p.n821 1.117
R9923 vp_p.n748 vp_p.n73 1.084
R9924 vp_p.n744 vp_p.n743 0.654
R9925 vp_p.n1497 vp_p.n822 0.509
R9926 vp_p.n523 vp_p.n521 0.356
R9927 vp_p.n374 vp_p.n372 0.356
R9928 vp_p.n225 vp_p.n223 0.356
R9929 vp_p.n76 vp_p.n74 0.356
R9930 vp_p.n825 vp_p.n823 0.356
R9931 vp_p.n974 vp_p.n972 0.356
R9932 vp_p.n1123 vp_p.n1121 0.356
R9933 vp_p.n1272 vp_p.n1270 0.356
R9934 vp_p.n744 vp_p.n669 0.319
R9935 vp_p.n746 vp_p.n371 0.319
R9936 vp_p.n1496 vp_p.n971 0.319
R9937 vp_p.n1494 vp_p.n1269 0.319
R9938 vp_p.n525 vp_p.n523 0.316
R9939 vp_p.n527 vp_p.n525 0.316
R9940 vp_p.n529 vp_p.n527 0.316
R9941 vp_p.n531 vp_p.n529 0.316
R9942 vp_p.n533 vp_p.n531 0.316
R9943 vp_p.n535 vp_p.n533 0.316
R9944 vp_p.n537 vp_p.n535 0.316
R9945 vp_p.n539 vp_p.n537 0.316
R9946 vp_p.n541 vp_p.n539 0.316
R9947 vp_p.n543 vp_p.n541 0.316
R9948 vp_p.n545 vp_p.n543 0.316
R9949 vp_p.n547 vp_p.n545 0.316
R9950 vp_p.n549 vp_p.n547 0.316
R9951 vp_p.n551 vp_p.n549 0.316
R9952 vp_p.n553 vp_p.n551 0.316
R9953 vp_p.n555 vp_p.n553 0.316
R9954 vp_p.n557 vp_p.n555 0.316
R9955 vp_p.n559 vp_p.n557 0.316
R9956 vp_p.n561 vp_p.n559 0.316
R9957 vp_p.n563 vp_p.n561 0.316
R9958 vp_p.n565 vp_p.n563 0.316
R9959 vp_p.n567 vp_p.n565 0.316
R9960 vp_p.n569 vp_p.n567 0.316
R9961 vp_p.n571 vp_p.n569 0.316
R9962 vp_p.n573 vp_p.n571 0.316
R9963 vp_p.n575 vp_p.n573 0.316
R9964 vp_p.n577 vp_p.n575 0.316
R9965 vp_p.n579 vp_p.n577 0.316
R9966 vp_p.n581 vp_p.n579 0.316
R9967 vp_p.n583 vp_p.n581 0.316
R9968 vp_p.n585 vp_p.n583 0.316
R9969 vp_p.n587 vp_p.n585 0.316
R9970 vp_p.n589 vp_p.n587 0.316
R9971 vp_p.n591 vp_p.n589 0.316
R9972 vp_p.n593 vp_p.n591 0.316
R9973 vp_p.n595 vp_p.n593 0.316
R9974 vp_p.n597 vp_p.n595 0.316
R9975 vp_p.n599 vp_p.n597 0.316
R9976 vp_p.n601 vp_p.n599 0.316
R9977 vp_p.n603 vp_p.n601 0.316
R9978 vp_p.n605 vp_p.n603 0.316
R9979 vp_p.n607 vp_p.n605 0.316
R9980 vp_p.n609 vp_p.n607 0.316
R9981 vp_p.n611 vp_p.n609 0.316
R9982 vp_p.n613 vp_p.n611 0.316
R9983 vp_p.n615 vp_p.n613 0.316
R9984 vp_p.n617 vp_p.n615 0.316
R9985 vp_p.n619 vp_p.n617 0.316
R9986 vp_p.n621 vp_p.n619 0.316
R9987 vp_p.n623 vp_p.n621 0.316
R9988 vp_p.n625 vp_p.n623 0.316
R9989 vp_p.n627 vp_p.n625 0.316
R9990 vp_p.n629 vp_p.n627 0.316
R9991 vp_p.n631 vp_p.n629 0.316
R9992 vp_p.n633 vp_p.n631 0.316
R9993 vp_p.n635 vp_p.n633 0.316
R9994 vp_p.n637 vp_p.n635 0.316
R9995 vp_p.n639 vp_p.n637 0.316
R9996 vp_p.n641 vp_p.n639 0.316
R9997 vp_p.n643 vp_p.n641 0.316
R9998 vp_p.n645 vp_p.n643 0.316
R9999 vp_p.n647 vp_p.n645 0.316
R10000 vp_p.n649 vp_p.n647 0.316
R10001 vp_p.n651 vp_p.n649 0.316
R10002 vp_p.n653 vp_p.n651 0.316
R10003 vp_p.n655 vp_p.n653 0.316
R10004 vp_p.n657 vp_p.n655 0.316
R10005 vp_p.n659 vp_p.n657 0.316
R10006 vp_p.n661 vp_p.n659 0.316
R10007 vp_p.n663 vp_p.n661 0.316
R10008 vp_p.n665 vp_p.n663 0.316
R10009 vp_p.n667 vp_p.n665 0.316
R10010 vp_p.n669 vp_p.n667 0.316
R10011 vp_p.n376 vp_p.n374 0.316
R10012 vp_p.n378 vp_p.n376 0.316
R10013 vp_p.n380 vp_p.n378 0.316
R10014 vp_p.n382 vp_p.n380 0.316
R10015 vp_p.n384 vp_p.n382 0.316
R10016 vp_p.n386 vp_p.n384 0.316
R10017 vp_p.n388 vp_p.n386 0.316
R10018 vp_p.n390 vp_p.n388 0.316
R10019 vp_p.n392 vp_p.n390 0.316
R10020 vp_p.n394 vp_p.n392 0.316
R10021 vp_p.n396 vp_p.n394 0.316
R10022 vp_p.n398 vp_p.n396 0.316
R10023 vp_p.n400 vp_p.n398 0.316
R10024 vp_p.n402 vp_p.n400 0.316
R10025 vp_p.n404 vp_p.n402 0.316
R10026 vp_p.n406 vp_p.n404 0.316
R10027 vp_p.n408 vp_p.n406 0.316
R10028 vp_p.n410 vp_p.n408 0.316
R10029 vp_p.n412 vp_p.n410 0.316
R10030 vp_p.n414 vp_p.n412 0.316
R10031 vp_p.n416 vp_p.n414 0.316
R10032 vp_p.n418 vp_p.n416 0.316
R10033 vp_p.n420 vp_p.n418 0.316
R10034 vp_p.n422 vp_p.n420 0.316
R10035 vp_p.n424 vp_p.n422 0.316
R10036 vp_p.n426 vp_p.n424 0.316
R10037 vp_p.n428 vp_p.n426 0.316
R10038 vp_p.n430 vp_p.n428 0.316
R10039 vp_p.n432 vp_p.n430 0.316
R10040 vp_p.n434 vp_p.n432 0.316
R10041 vp_p.n436 vp_p.n434 0.316
R10042 vp_p.n438 vp_p.n436 0.316
R10043 vp_p.n440 vp_p.n438 0.316
R10044 vp_p.n442 vp_p.n440 0.316
R10045 vp_p.n444 vp_p.n442 0.316
R10046 vp_p.n446 vp_p.n444 0.316
R10047 vp_p.n448 vp_p.n446 0.316
R10048 vp_p.n450 vp_p.n448 0.316
R10049 vp_p.n452 vp_p.n450 0.316
R10050 vp_p.n454 vp_p.n452 0.316
R10051 vp_p.n456 vp_p.n454 0.316
R10052 vp_p.n458 vp_p.n456 0.316
R10053 vp_p.n460 vp_p.n458 0.316
R10054 vp_p.n462 vp_p.n460 0.316
R10055 vp_p.n464 vp_p.n462 0.316
R10056 vp_p.n466 vp_p.n464 0.316
R10057 vp_p.n468 vp_p.n466 0.316
R10058 vp_p.n470 vp_p.n468 0.316
R10059 vp_p.n472 vp_p.n470 0.316
R10060 vp_p.n474 vp_p.n472 0.316
R10061 vp_p.n476 vp_p.n474 0.316
R10062 vp_p.n478 vp_p.n476 0.316
R10063 vp_p.n480 vp_p.n478 0.316
R10064 vp_p.n482 vp_p.n480 0.316
R10065 vp_p.n484 vp_p.n482 0.316
R10066 vp_p.n486 vp_p.n484 0.316
R10067 vp_p.n488 vp_p.n486 0.316
R10068 vp_p.n490 vp_p.n488 0.316
R10069 vp_p.n492 vp_p.n490 0.316
R10070 vp_p.n494 vp_p.n492 0.316
R10071 vp_p.n496 vp_p.n494 0.316
R10072 vp_p.n498 vp_p.n496 0.316
R10073 vp_p.n500 vp_p.n498 0.316
R10074 vp_p.n502 vp_p.n500 0.316
R10075 vp_p.n504 vp_p.n502 0.316
R10076 vp_p.n506 vp_p.n504 0.316
R10077 vp_p.n508 vp_p.n506 0.316
R10078 vp_p.n510 vp_p.n508 0.316
R10079 vp_p.n512 vp_p.n510 0.316
R10080 vp_p.n514 vp_p.n512 0.316
R10081 vp_p.n516 vp_p.n514 0.316
R10082 vp_p.n518 vp_p.n516 0.316
R10083 vp_p.n520 vp_p.n518 0.316
R10084 vp_p.n227 vp_p.n225 0.316
R10085 vp_p.n229 vp_p.n227 0.316
R10086 vp_p.n231 vp_p.n229 0.316
R10087 vp_p.n233 vp_p.n231 0.316
R10088 vp_p.n235 vp_p.n233 0.316
R10089 vp_p.n237 vp_p.n235 0.316
R10090 vp_p.n239 vp_p.n237 0.316
R10091 vp_p.n241 vp_p.n239 0.316
R10092 vp_p.n243 vp_p.n241 0.316
R10093 vp_p.n245 vp_p.n243 0.316
R10094 vp_p.n247 vp_p.n245 0.316
R10095 vp_p.n249 vp_p.n247 0.316
R10096 vp_p.n251 vp_p.n249 0.316
R10097 vp_p.n253 vp_p.n251 0.316
R10098 vp_p.n255 vp_p.n253 0.316
R10099 vp_p.n257 vp_p.n255 0.316
R10100 vp_p.n259 vp_p.n257 0.316
R10101 vp_p.n261 vp_p.n259 0.316
R10102 vp_p.n263 vp_p.n261 0.316
R10103 vp_p.n265 vp_p.n263 0.316
R10104 vp_p.n267 vp_p.n265 0.316
R10105 vp_p.n269 vp_p.n267 0.316
R10106 vp_p.n271 vp_p.n269 0.316
R10107 vp_p.n273 vp_p.n271 0.316
R10108 vp_p.n275 vp_p.n273 0.316
R10109 vp_p.n277 vp_p.n275 0.316
R10110 vp_p.n279 vp_p.n277 0.316
R10111 vp_p.n281 vp_p.n279 0.316
R10112 vp_p.n283 vp_p.n281 0.316
R10113 vp_p.n285 vp_p.n283 0.316
R10114 vp_p.n287 vp_p.n285 0.316
R10115 vp_p.n289 vp_p.n287 0.316
R10116 vp_p.n291 vp_p.n289 0.316
R10117 vp_p.n293 vp_p.n291 0.316
R10118 vp_p.n295 vp_p.n293 0.316
R10119 vp_p.n297 vp_p.n295 0.316
R10120 vp_p.n299 vp_p.n297 0.316
R10121 vp_p.n301 vp_p.n299 0.316
R10122 vp_p.n303 vp_p.n301 0.316
R10123 vp_p.n305 vp_p.n303 0.316
R10124 vp_p.n307 vp_p.n305 0.316
R10125 vp_p.n309 vp_p.n307 0.316
R10126 vp_p.n311 vp_p.n309 0.316
R10127 vp_p.n313 vp_p.n311 0.316
R10128 vp_p.n315 vp_p.n313 0.316
R10129 vp_p.n317 vp_p.n315 0.316
R10130 vp_p.n319 vp_p.n317 0.316
R10131 vp_p.n321 vp_p.n319 0.316
R10132 vp_p.n323 vp_p.n321 0.316
R10133 vp_p.n325 vp_p.n323 0.316
R10134 vp_p.n327 vp_p.n325 0.316
R10135 vp_p.n329 vp_p.n327 0.316
R10136 vp_p.n331 vp_p.n329 0.316
R10137 vp_p.n333 vp_p.n331 0.316
R10138 vp_p.n335 vp_p.n333 0.316
R10139 vp_p.n337 vp_p.n335 0.316
R10140 vp_p.n339 vp_p.n337 0.316
R10141 vp_p.n341 vp_p.n339 0.316
R10142 vp_p.n343 vp_p.n341 0.316
R10143 vp_p.n345 vp_p.n343 0.316
R10144 vp_p.n347 vp_p.n345 0.316
R10145 vp_p.n349 vp_p.n347 0.316
R10146 vp_p.n351 vp_p.n349 0.316
R10147 vp_p.n353 vp_p.n351 0.316
R10148 vp_p.n355 vp_p.n353 0.316
R10149 vp_p.n357 vp_p.n355 0.316
R10150 vp_p.n359 vp_p.n357 0.316
R10151 vp_p.n361 vp_p.n359 0.316
R10152 vp_p.n363 vp_p.n361 0.316
R10153 vp_p.n365 vp_p.n363 0.316
R10154 vp_p.n367 vp_p.n365 0.316
R10155 vp_p.n369 vp_p.n367 0.316
R10156 vp_p.n371 vp_p.n369 0.316
R10157 vp_p.n78 vp_p.n76 0.316
R10158 vp_p.n80 vp_p.n78 0.316
R10159 vp_p.n82 vp_p.n80 0.316
R10160 vp_p.n84 vp_p.n82 0.316
R10161 vp_p.n86 vp_p.n84 0.316
R10162 vp_p.n88 vp_p.n86 0.316
R10163 vp_p.n90 vp_p.n88 0.316
R10164 vp_p.n92 vp_p.n90 0.316
R10165 vp_p.n94 vp_p.n92 0.316
R10166 vp_p.n96 vp_p.n94 0.316
R10167 vp_p.n98 vp_p.n96 0.316
R10168 vp_p.n100 vp_p.n98 0.316
R10169 vp_p.n102 vp_p.n100 0.316
R10170 vp_p.n104 vp_p.n102 0.316
R10171 vp_p.n106 vp_p.n104 0.316
R10172 vp_p.n108 vp_p.n106 0.316
R10173 vp_p.n110 vp_p.n108 0.316
R10174 vp_p.n112 vp_p.n110 0.316
R10175 vp_p.n114 vp_p.n112 0.316
R10176 vp_p.n116 vp_p.n114 0.316
R10177 vp_p.n118 vp_p.n116 0.316
R10178 vp_p.n120 vp_p.n118 0.316
R10179 vp_p.n122 vp_p.n120 0.316
R10180 vp_p.n124 vp_p.n122 0.316
R10181 vp_p.n126 vp_p.n124 0.316
R10182 vp_p.n128 vp_p.n126 0.316
R10183 vp_p.n130 vp_p.n128 0.316
R10184 vp_p.n132 vp_p.n130 0.316
R10185 vp_p.n134 vp_p.n132 0.316
R10186 vp_p.n136 vp_p.n134 0.316
R10187 vp_p.n138 vp_p.n136 0.316
R10188 vp_p.n140 vp_p.n138 0.316
R10189 vp_p.n142 vp_p.n140 0.316
R10190 vp_p.n144 vp_p.n142 0.316
R10191 vp_p.n146 vp_p.n144 0.316
R10192 vp_p.n148 vp_p.n146 0.316
R10193 vp_p.n150 vp_p.n148 0.316
R10194 vp_p.n152 vp_p.n150 0.316
R10195 vp_p.n154 vp_p.n152 0.316
R10196 vp_p.n156 vp_p.n154 0.316
R10197 vp_p.n158 vp_p.n156 0.316
R10198 vp_p.n160 vp_p.n158 0.316
R10199 vp_p.n162 vp_p.n160 0.316
R10200 vp_p.n164 vp_p.n162 0.316
R10201 vp_p.n166 vp_p.n164 0.316
R10202 vp_p.n168 vp_p.n166 0.316
R10203 vp_p.n170 vp_p.n168 0.316
R10204 vp_p.n172 vp_p.n170 0.316
R10205 vp_p.n174 vp_p.n172 0.316
R10206 vp_p.n176 vp_p.n174 0.316
R10207 vp_p.n178 vp_p.n176 0.316
R10208 vp_p.n180 vp_p.n178 0.316
R10209 vp_p.n182 vp_p.n180 0.316
R10210 vp_p.n184 vp_p.n182 0.316
R10211 vp_p.n186 vp_p.n184 0.316
R10212 vp_p.n188 vp_p.n186 0.316
R10213 vp_p.n190 vp_p.n188 0.316
R10214 vp_p.n192 vp_p.n190 0.316
R10215 vp_p.n194 vp_p.n192 0.316
R10216 vp_p.n196 vp_p.n194 0.316
R10217 vp_p.n198 vp_p.n196 0.316
R10218 vp_p.n200 vp_p.n198 0.316
R10219 vp_p.n202 vp_p.n200 0.316
R10220 vp_p.n204 vp_p.n202 0.316
R10221 vp_p.n206 vp_p.n204 0.316
R10222 vp_p.n208 vp_p.n206 0.316
R10223 vp_p.n210 vp_p.n208 0.316
R10224 vp_p.n212 vp_p.n210 0.316
R10225 vp_p.n214 vp_p.n212 0.316
R10226 vp_p.n216 vp_p.n214 0.316
R10227 vp_p.n218 vp_p.n216 0.316
R10228 vp_p.n220 vp_p.n218 0.316
R10229 vp_p.n222 vp_p.n220 0.316
R10230 vp_p.n827 vp_p.n825 0.316
R10231 vp_p.n829 vp_p.n827 0.316
R10232 vp_p.n831 vp_p.n829 0.316
R10233 vp_p.n833 vp_p.n831 0.316
R10234 vp_p.n835 vp_p.n833 0.316
R10235 vp_p.n837 vp_p.n835 0.316
R10236 vp_p.n839 vp_p.n837 0.316
R10237 vp_p.n841 vp_p.n839 0.316
R10238 vp_p.n843 vp_p.n841 0.316
R10239 vp_p.n845 vp_p.n843 0.316
R10240 vp_p.n847 vp_p.n845 0.316
R10241 vp_p.n849 vp_p.n847 0.316
R10242 vp_p.n851 vp_p.n849 0.316
R10243 vp_p.n853 vp_p.n851 0.316
R10244 vp_p.n855 vp_p.n853 0.316
R10245 vp_p.n857 vp_p.n855 0.316
R10246 vp_p.n859 vp_p.n857 0.316
R10247 vp_p.n861 vp_p.n859 0.316
R10248 vp_p.n863 vp_p.n861 0.316
R10249 vp_p.n865 vp_p.n863 0.316
R10250 vp_p.n867 vp_p.n865 0.316
R10251 vp_p.n869 vp_p.n867 0.316
R10252 vp_p.n871 vp_p.n869 0.316
R10253 vp_p.n873 vp_p.n871 0.316
R10254 vp_p.n875 vp_p.n873 0.316
R10255 vp_p.n877 vp_p.n875 0.316
R10256 vp_p.n879 vp_p.n877 0.316
R10257 vp_p.n881 vp_p.n879 0.316
R10258 vp_p.n883 vp_p.n881 0.316
R10259 vp_p.n885 vp_p.n883 0.316
R10260 vp_p.n887 vp_p.n885 0.316
R10261 vp_p.n889 vp_p.n887 0.316
R10262 vp_p.n891 vp_p.n889 0.316
R10263 vp_p.n893 vp_p.n891 0.316
R10264 vp_p.n895 vp_p.n893 0.316
R10265 vp_p.n897 vp_p.n895 0.316
R10266 vp_p.n899 vp_p.n897 0.316
R10267 vp_p.n901 vp_p.n899 0.316
R10268 vp_p.n903 vp_p.n901 0.316
R10269 vp_p.n905 vp_p.n903 0.316
R10270 vp_p.n907 vp_p.n905 0.316
R10271 vp_p.n909 vp_p.n907 0.316
R10272 vp_p.n911 vp_p.n909 0.316
R10273 vp_p.n913 vp_p.n911 0.316
R10274 vp_p.n915 vp_p.n913 0.316
R10275 vp_p.n917 vp_p.n915 0.316
R10276 vp_p.n919 vp_p.n917 0.316
R10277 vp_p.n921 vp_p.n919 0.316
R10278 vp_p.n923 vp_p.n921 0.316
R10279 vp_p.n925 vp_p.n923 0.316
R10280 vp_p.n927 vp_p.n925 0.316
R10281 vp_p.n929 vp_p.n927 0.316
R10282 vp_p.n931 vp_p.n929 0.316
R10283 vp_p.n933 vp_p.n931 0.316
R10284 vp_p.n935 vp_p.n933 0.316
R10285 vp_p.n937 vp_p.n935 0.316
R10286 vp_p.n939 vp_p.n937 0.316
R10287 vp_p.n941 vp_p.n939 0.316
R10288 vp_p.n943 vp_p.n941 0.316
R10289 vp_p.n945 vp_p.n943 0.316
R10290 vp_p.n947 vp_p.n945 0.316
R10291 vp_p.n949 vp_p.n947 0.316
R10292 vp_p.n951 vp_p.n949 0.316
R10293 vp_p.n953 vp_p.n951 0.316
R10294 vp_p.n955 vp_p.n953 0.316
R10295 vp_p.n957 vp_p.n955 0.316
R10296 vp_p.n959 vp_p.n957 0.316
R10297 vp_p.n961 vp_p.n959 0.316
R10298 vp_p.n963 vp_p.n961 0.316
R10299 vp_p.n965 vp_p.n963 0.316
R10300 vp_p.n967 vp_p.n965 0.316
R10301 vp_p.n969 vp_p.n967 0.316
R10302 vp_p.n971 vp_p.n969 0.316
R10303 vp_p.n976 vp_p.n974 0.316
R10304 vp_p.n978 vp_p.n976 0.316
R10305 vp_p.n980 vp_p.n978 0.316
R10306 vp_p.n982 vp_p.n980 0.316
R10307 vp_p.n984 vp_p.n982 0.316
R10308 vp_p.n986 vp_p.n984 0.316
R10309 vp_p.n988 vp_p.n986 0.316
R10310 vp_p.n990 vp_p.n988 0.316
R10311 vp_p.n992 vp_p.n990 0.316
R10312 vp_p.n994 vp_p.n992 0.316
R10313 vp_p.n996 vp_p.n994 0.316
R10314 vp_p.n998 vp_p.n996 0.316
R10315 vp_p.n1000 vp_p.n998 0.316
R10316 vp_p.n1002 vp_p.n1000 0.316
R10317 vp_p.n1004 vp_p.n1002 0.316
R10318 vp_p.n1006 vp_p.n1004 0.316
R10319 vp_p.n1008 vp_p.n1006 0.316
R10320 vp_p.n1010 vp_p.n1008 0.316
R10321 vp_p.n1012 vp_p.n1010 0.316
R10322 vp_p.n1014 vp_p.n1012 0.316
R10323 vp_p.n1016 vp_p.n1014 0.316
R10324 vp_p.n1018 vp_p.n1016 0.316
R10325 vp_p.n1020 vp_p.n1018 0.316
R10326 vp_p.n1022 vp_p.n1020 0.316
R10327 vp_p.n1024 vp_p.n1022 0.316
R10328 vp_p.n1026 vp_p.n1024 0.316
R10329 vp_p.n1028 vp_p.n1026 0.316
R10330 vp_p.n1030 vp_p.n1028 0.316
R10331 vp_p.n1032 vp_p.n1030 0.316
R10332 vp_p.n1034 vp_p.n1032 0.316
R10333 vp_p.n1036 vp_p.n1034 0.316
R10334 vp_p.n1038 vp_p.n1036 0.316
R10335 vp_p.n1040 vp_p.n1038 0.316
R10336 vp_p.n1042 vp_p.n1040 0.316
R10337 vp_p.n1044 vp_p.n1042 0.316
R10338 vp_p.n1046 vp_p.n1044 0.316
R10339 vp_p.n1048 vp_p.n1046 0.316
R10340 vp_p.n1050 vp_p.n1048 0.316
R10341 vp_p.n1052 vp_p.n1050 0.316
R10342 vp_p.n1054 vp_p.n1052 0.316
R10343 vp_p.n1056 vp_p.n1054 0.316
R10344 vp_p.n1058 vp_p.n1056 0.316
R10345 vp_p.n1060 vp_p.n1058 0.316
R10346 vp_p.n1062 vp_p.n1060 0.316
R10347 vp_p.n1064 vp_p.n1062 0.316
R10348 vp_p.n1066 vp_p.n1064 0.316
R10349 vp_p.n1068 vp_p.n1066 0.316
R10350 vp_p.n1070 vp_p.n1068 0.316
R10351 vp_p.n1072 vp_p.n1070 0.316
R10352 vp_p.n1074 vp_p.n1072 0.316
R10353 vp_p.n1076 vp_p.n1074 0.316
R10354 vp_p.n1078 vp_p.n1076 0.316
R10355 vp_p.n1080 vp_p.n1078 0.316
R10356 vp_p.n1082 vp_p.n1080 0.316
R10357 vp_p.n1084 vp_p.n1082 0.316
R10358 vp_p.n1086 vp_p.n1084 0.316
R10359 vp_p.n1088 vp_p.n1086 0.316
R10360 vp_p.n1090 vp_p.n1088 0.316
R10361 vp_p.n1092 vp_p.n1090 0.316
R10362 vp_p.n1094 vp_p.n1092 0.316
R10363 vp_p.n1096 vp_p.n1094 0.316
R10364 vp_p.n1098 vp_p.n1096 0.316
R10365 vp_p.n1100 vp_p.n1098 0.316
R10366 vp_p.n1102 vp_p.n1100 0.316
R10367 vp_p.n1104 vp_p.n1102 0.316
R10368 vp_p.n1106 vp_p.n1104 0.316
R10369 vp_p.n1108 vp_p.n1106 0.316
R10370 vp_p.n1110 vp_p.n1108 0.316
R10371 vp_p.n1112 vp_p.n1110 0.316
R10372 vp_p.n1114 vp_p.n1112 0.316
R10373 vp_p.n1116 vp_p.n1114 0.316
R10374 vp_p.n1118 vp_p.n1116 0.316
R10375 vp_p.n1120 vp_p.n1118 0.316
R10376 vp_p.n1125 vp_p.n1123 0.316
R10377 vp_p.n1127 vp_p.n1125 0.316
R10378 vp_p.n1129 vp_p.n1127 0.316
R10379 vp_p.n1131 vp_p.n1129 0.316
R10380 vp_p.n1133 vp_p.n1131 0.316
R10381 vp_p.n1135 vp_p.n1133 0.316
R10382 vp_p.n1137 vp_p.n1135 0.316
R10383 vp_p.n1139 vp_p.n1137 0.316
R10384 vp_p.n1141 vp_p.n1139 0.316
R10385 vp_p.n1143 vp_p.n1141 0.316
R10386 vp_p.n1145 vp_p.n1143 0.316
R10387 vp_p.n1147 vp_p.n1145 0.316
R10388 vp_p.n1149 vp_p.n1147 0.316
R10389 vp_p.n1151 vp_p.n1149 0.316
R10390 vp_p.n1153 vp_p.n1151 0.316
R10391 vp_p.n1155 vp_p.n1153 0.316
R10392 vp_p.n1157 vp_p.n1155 0.316
R10393 vp_p.n1159 vp_p.n1157 0.316
R10394 vp_p.n1161 vp_p.n1159 0.316
R10395 vp_p.n1163 vp_p.n1161 0.316
R10396 vp_p.n1165 vp_p.n1163 0.316
R10397 vp_p.n1167 vp_p.n1165 0.316
R10398 vp_p.n1169 vp_p.n1167 0.316
R10399 vp_p.n1171 vp_p.n1169 0.316
R10400 vp_p.n1173 vp_p.n1171 0.316
R10401 vp_p.n1175 vp_p.n1173 0.316
R10402 vp_p.n1177 vp_p.n1175 0.316
R10403 vp_p.n1179 vp_p.n1177 0.316
R10404 vp_p.n1181 vp_p.n1179 0.316
R10405 vp_p.n1183 vp_p.n1181 0.316
R10406 vp_p.n1185 vp_p.n1183 0.316
R10407 vp_p.n1187 vp_p.n1185 0.316
R10408 vp_p.n1189 vp_p.n1187 0.316
R10409 vp_p.n1191 vp_p.n1189 0.316
R10410 vp_p.n1193 vp_p.n1191 0.316
R10411 vp_p.n1195 vp_p.n1193 0.316
R10412 vp_p.n1197 vp_p.n1195 0.316
R10413 vp_p.n1199 vp_p.n1197 0.316
R10414 vp_p.n1201 vp_p.n1199 0.316
R10415 vp_p.n1203 vp_p.n1201 0.316
R10416 vp_p.n1205 vp_p.n1203 0.316
R10417 vp_p.n1207 vp_p.n1205 0.316
R10418 vp_p.n1209 vp_p.n1207 0.316
R10419 vp_p.n1211 vp_p.n1209 0.316
R10420 vp_p.n1213 vp_p.n1211 0.316
R10421 vp_p.n1215 vp_p.n1213 0.316
R10422 vp_p.n1217 vp_p.n1215 0.316
R10423 vp_p.n1219 vp_p.n1217 0.316
R10424 vp_p.n1221 vp_p.n1219 0.316
R10425 vp_p.n1223 vp_p.n1221 0.316
R10426 vp_p.n1225 vp_p.n1223 0.316
R10427 vp_p.n1227 vp_p.n1225 0.316
R10428 vp_p.n1229 vp_p.n1227 0.316
R10429 vp_p.n1231 vp_p.n1229 0.316
R10430 vp_p.n1233 vp_p.n1231 0.316
R10431 vp_p.n1235 vp_p.n1233 0.316
R10432 vp_p.n1237 vp_p.n1235 0.316
R10433 vp_p.n1239 vp_p.n1237 0.316
R10434 vp_p.n1241 vp_p.n1239 0.316
R10435 vp_p.n1243 vp_p.n1241 0.316
R10436 vp_p.n1245 vp_p.n1243 0.316
R10437 vp_p.n1247 vp_p.n1245 0.316
R10438 vp_p.n1249 vp_p.n1247 0.316
R10439 vp_p.n1251 vp_p.n1249 0.316
R10440 vp_p.n1253 vp_p.n1251 0.316
R10441 vp_p.n1255 vp_p.n1253 0.316
R10442 vp_p.n1257 vp_p.n1255 0.316
R10443 vp_p.n1259 vp_p.n1257 0.316
R10444 vp_p.n1261 vp_p.n1259 0.316
R10445 vp_p.n1263 vp_p.n1261 0.316
R10446 vp_p.n1265 vp_p.n1263 0.316
R10447 vp_p.n1267 vp_p.n1265 0.316
R10448 vp_p.n1269 vp_p.n1267 0.316
R10449 vp_p.n1274 vp_p.n1272 0.316
R10450 vp_p.n1276 vp_p.n1274 0.316
R10451 vp_p.n1278 vp_p.n1276 0.316
R10452 vp_p.n1280 vp_p.n1278 0.316
R10453 vp_p.n1282 vp_p.n1280 0.316
R10454 vp_p.n1284 vp_p.n1282 0.316
R10455 vp_p.n1286 vp_p.n1284 0.316
R10456 vp_p.n1288 vp_p.n1286 0.316
R10457 vp_p.n1290 vp_p.n1288 0.316
R10458 vp_p.n1292 vp_p.n1290 0.316
R10459 vp_p.n1294 vp_p.n1292 0.316
R10460 vp_p.n1296 vp_p.n1294 0.316
R10461 vp_p.n1298 vp_p.n1296 0.316
R10462 vp_p.n1300 vp_p.n1298 0.316
R10463 vp_p.n1302 vp_p.n1300 0.316
R10464 vp_p.n1304 vp_p.n1302 0.316
R10465 vp_p.n1306 vp_p.n1304 0.316
R10466 vp_p.n1308 vp_p.n1306 0.316
R10467 vp_p.n1310 vp_p.n1308 0.316
R10468 vp_p.n1312 vp_p.n1310 0.316
R10469 vp_p.n1314 vp_p.n1312 0.316
R10470 vp_p.n1316 vp_p.n1314 0.316
R10471 vp_p.n1318 vp_p.n1316 0.316
R10472 vp_p.n1320 vp_p.n1318 0.316
R10473 vp_p.n1322 vp_p.n1320 0.316
R10474 vp_p.n1324 vp_p.n1322 0.316
R10475 vp_p.n1326 vp_p.n1324 0.316
R10476 vp_p.n1328 vp_p.n1326 0.316
R10477 vp_p.n1330 vp_p.n1328 0.316
R10478 vp_p.n1332 vp_p.n1330 0.316
R10479 vp_p.n1334 vp_p.n1332 0.316
R10480 vp_p.n1336 vp_p.n1334 0.316
R10481 vp_p.n1338 vp_p.n1336 0.316
R10482 vp_p.n1340 vp_p.n1338 0.316
R10483 vp_p.n1342 vp_p.n1340 0.316
R10484 vp_p.n1344 vp_p.n1342 0.316
R10485 vp_p.n1346 vp_p.n1344 0.316
R10486 vp_p.n1348 vp_p.n1346 0.316
R10487 vp_p.n1350 vp_p.n1348 0.316
R10488 vp_p.n1352 vp_p.n1350 0.316
R10489 vp_p.n1354 vp_p.n1352 0.316
R10490 vp_p.n1356 vp_p.n1354 0.316
R10491 vp_p.n1358 vp_p.n1356 0.316
R10492 vp_p.n1360 vp_p.n1358 0.316
R10493 vp_p.n1362 vp_p.n1360 0.316
R10494 vp_p.n1364 vp_p.n1362 0.316
R10495 vp_p.n1366 vp_p.n1364 0.316
R10496 vp_p.n1368 vp_p.n1366 0.316
R10497 vp_p.n1370 vp_p.n1368 0.316
R10498 vp_p.n1372 vp_p.n1370 0.316
R10499 vp_p.n1374 vp_p.n1372 0.316
R10500 vp_p.n1376 vp_p.n1374 0.316
R10501 vp_p.n1378 vp_p.n1376 0.316
R10502 vp_p.n1380 vp_p.n1378 0.316
R10503 vp_p.n1382 vp_p.n1380 0.316
R10504 vp_p.n1384 vp_p.n1382 0.316
R10505 vp_p.n1386 vp_p.n1384 0.316
R10506 vp_p.n1388 vp_p.n1386 0.316
R10507 vp_p.n1390 vp_p.n1388 0.316
R10508 vp_p.n1392 vp_p.n1390 0.316
R10509 vp_p.n1394 vp_p.n1392 0.316
R10510 vp_p.n1396 vp_p.n1394 0.316
R10511 vp_p.n1398 vp_p.n1396 0.316
R10512 vp_p.n1400 vp_p.n1398 0.316
R10513 vp_p.n1402 vp_p.n1400 0.316
R10514 vp_p.n1404 vp_p.n1402 0.316
R10515 vp_p.n1406 vp_p.n1404 0.316
R10516 vp_p.n1408 vp_p.n1406 0.316
R10517 vp_p.n1410 vp_p.n1408 0.316
R10518 vp_p.n1412 vp_p.n1410 0.316
R10519 vp_p.n1414 vp_p.n1412 0.316
R10520 vp_p.n1416 vp_p.n1414 0.316
R10521 vp_p.n1418 vp_p.n1416 0.316
R10522 vp_p.n745 vp_p.n744 0.149
R10523 vp_p.n747 vp_p.n746 0.149
R10524 vp_p.n1496 vp_p.n1495 0.149
R10525 vp_p.n1495 vp_p.n1494 0.149
R10526 vp_p.n1494 vp_p.n1493 0.149
R10527 vp_p.n748 vp_p.n747 0.141
R10528 vp_p.n1497 vp_p.n1496 0.141
R10529 vp_p.n746 vp_p 0.137
R10530 vp_p.n745 vp_p.n520 0.134
R10531 vp_p.n747 vp_p.n222 0.134
R10532 vp_p.n1495 vp_p.n1120 0.134
R10533 vp_p.n1493 vp_p.n1418 0.134
R10534 vp_p.n669 vp_p.n668 0.04
R10535 vp_p.n667 vp_p.n666 0.04
R10536 vp_p.n665 vp_p.n664 0.04
R10537 vp_p.n663 vp_p.n662 0.04
R10538 vp_p.n661 vp_p.n660 0.04
R10539 vp_p.n659 vp_p.n658 0.04
R10540 vp_p.n657 vp_p.n656 0.04
R10541 vp_p.n655 vp_p.n654 0.04
R10542 vp_p.n653 vp_p.n652 0.04
R10543 vp_p.n651 vp_p.n650 0.04
R10544 vp_p.n649 vp_p.n648 0.04
R10545 vp_p.n647 vp_p.n646 0.04
R10546 vp_p.n645 vp_p.n644 0.04
R10547 vp_p.n643 vp_p.n642 0.04
R10548 vp_p.n641 vp_p.n640 0.04
R10549 vp_p.n639 vp_p.n638 0.04
R10550 vp_p.n637 vp_p.n636 0.04
R10551 vp_p.n635 vp_p.n634 0.04
R10552 vp_p.n633 vp_p.n632 0.04
R10553 vp_p.n631 vp_p.n630 0.04
R10554 vp_p.n629 vp_p.n628 0.04
R10555 vp_p.n627 vp_p.n626 0.04
R10556 vp_p.n625 vp_p.n624 0.04
R10557 vp_p.n623 vp_p.n622 0.04
R10558 vp_p.n621 vp_p.n620 0.04
R10559 vp_p.n619 vp_p.n618 0.04
R10560 vp_p.n617 vp_p.n616 0.04
R10561 vp_p.n615 vp_p.n614 0.04
R10562 vp_p.n613 vp_p.n612 0.04
R10563 vp_p.n611 vp_p.n610 0.04
R10564 vp_p.n609 vp_p.n608 0.04
R10565 vp_p.n607 vp_p.n606 0.04
R10566 vp_p.n605 vp_p.n604 0.04
R10567 vp_p.n603 vp_p.n602 0.04
R10568 vp_p.n601 vp_p.n600 0.04
R10569 vp_p.n599 vp_p.n598 0.04
R10570 vp_p.n597 vp_p.n596 0.04
R10571 vp_p.n595 vp_p.n594 0.04
R10572 vp_p.n593 vp_p.n592 0.04
R10573 vp_p.n591 vp_p.n590 0.04
R10574 vp_p.n589 vp_p.n588 0.04
R10575 vp_p.n587 vp_p.n586 0.04
R10576 vp_p.n585 vp_p.n584 0.04
R10577 vp_p.n583 vp_p.n582 0.04
R10578 vp_p.n581 vp_p.n580 0.04
R10579 vp_p.n579 vp_p.n578 0.04
R10580 vp_p.n577 vp_p.n576 0.04
R10581 vp_p.n575 vp_p.n574 0.04
R10582 vp_p.n573 vp_p.n572 0.04
R10583 vp_p.n571 vp_p.n570 0.04
R10584 vp_p.n569 vp_p.n568 0.04
R10585 vp_p.n567 vp_p.n566 0.04
R10586 vp_p.n565 vp_p.n564 0.04
R10587 vp_p.n563 vp_p.n562 0.04
R10588 vp_p.n561 vp_p.n560 0.04
R10589 vp_p.n559 vp_p.n558 0.04
R10590 vp_p.n557 vp_p.n556 0.04
R10591 vp_p.n555 vp_p.n554 0.04
R10592 vp_p.n553 vp_p.n552 0.04
R10593 vp_p.n551 vp_p.n550 0.04
R10594 vp_p.n549 vp_p.n548 0.04
R10595 vp_p.n547 vp_p.n546 0.04
R10596 vp_p.n545 vp_p.n544 0.04
R10597 vp_p.n543 vp_p.n542 0.04
R10598 vp_p.n541 vp_p.n540 0.04
R10599 vp_p.n539 vp_p.n538 0.04
R10600 vp_p.n537 vp_p.n536 0.04
R10601 vp_p.n535 vp_p.n534 0.04
R10602 vp_p.n533 vp_p.n532 0.04
R10603 vp_p.n531 vp_p.n530 0.04
R10604 vp_p.n529 vp_p.n528 0.04
R10605 vp_p.n527 vp_p.n526 0.04
R10606 vp_p.n525 vp_p.n524 0.04
R10607 vp_p.n523 vp_p.n522 0.04
R10608 vp_p.n520 vp_p.n519 0.04
R10609 vp_p.n518 vp_p.n517 0.04
R10610 vp_p.n516 vp_p.n515 0.04
R10611 vp_p.n514 vp_p.n513 0.04
R10612 vp_p.n512 vp_p.n511 0.04
R10613 vp_p.n510 vp_p.n509 0.04
R10614 vp_p.n508 vp_p.n507 0.04
R10615 vp_p.n506 vp_p.n505 0.04
R10616 vp_p.n504 vp_p.n503 0.04
R10617 vp_p.n502 vp_p.n501 0.04
R10618 vp_p.n500 vp_p.n499 0.04
R10619 vp_p.n498 vp_p.n497 0.04
R10620 vp_p.n496 vp_p.n495 0.04
R10621 vp_p.n494 vp_p.n493 0.04
R10622 vp_p.n492 vp_p.n491 0.04
R10623 vp_p.n490 vp_p.n489 0.04
R10624 vp_p.n488 vp_p.n487 0.04
R10625 vp_p.n486 vp_p.n485 0.04
R10626 vp_p.n484 vp_p.n483 0.04
R10627 vp_p.n482 vp_p.n481 0.04
R10628 vp_p.n480 vp_p.n479 0.04
R10629 vp_p.n478 vp_p.n477 0.04
R10630 vp_p.n476 vp_p.n475 0.04
R10631 vp_p.n474 vp_p.n473 0.04
R10632 vp_p.n472 vp_p.n471 0.04
R10633 vp_p.n470 vp_p.n469 0.04
R10634 vp_p.n468 vp_p.n467 0.04
R10635 vp_p.n466 vp_p.n465 0.04
R10636 vp_p.n464 vp_p.n463 0.04
R10637 vp_p.n462 vp_p.n461 0.04
R10638 vp_p.n460 vp_p.n459 0.04
R10639 vp_p.n458 vp_p.n457 0.04
R10640 vp_p.n456 vp_p.n455 0.04
R10641 vp_p.n454 vp_p.n453 0.04
R10642 vp_p.n452 vp_p.n451 0.04
R10643 vp_p.n450 vp_p.n449 0.04
R10644 vp_p.n448 vp_p.n447 0.04
R10645 vp_p.n446 vp_p.n445 0.04
R10646 vp_p.n444 vp_p.n443 0.04
R10647 vp_p.n442 vp_p.n441 0.04
R10648 vp_p.n440 vp_p.n439 0.04
R10649 vp_p.n438 vp_p.n437 0.04
R10650 vp_p.n436 vp_p.n435 0.04
R10651 vp_p.n434 vp_p.n433 0.04
R10652 vp_p.n432 vp_p.n431 0.04
R10653 vp_p.n430 vp_p.n429 0.04
R10654 vp_p.n428 vp_p.n427 0.04
R10655 vp_p.n426 vp_p.n425 0.04
R10656 vp_p.n424 vp_p.n423 0.04
R10657 vp_p.n422 vp_p.n421 0.04
R10658 vp_p.n420 vp_p.n419 0.04
R10659 vp_p.n418 vp_p.n417 0.04
R10660 vp_p.n416 vp_p.n415 0.04
R10661 vp_p.n414 vp_p.n413 0.04
R10662 vp_p.n412 vp_p.n411 0.04
R10663 vp_p.n410 vp_p.n409 0.04
R10664 vp_p.n408 vp_p.n407 0.04
R10665 vp_p.n406 vp_p.n405 0.04
R10666 vp_p.n404 vp_p.n403 0.04
R10667 vp_p.n402 vp_p.n401 0.04
R10668 vp_p.n400 vp_p.n399 0.04
R10669 vp_p.n398 vp_p.n397 0.04
R10670 vp_p.n396 vp_p.n395 0.04
R10671 vp_p.n394 vp_p.n393 0.04
R10672 vp_p.n392 vp_p.n391 0.04
R10673 vp_p.n390 vp_p.n389 0.04
R10674 vp_p.n388 vp_p.n387 0.04
R10675 vp_p.n386 vp_p.n385 0.04
R10676 vp_p.n384 vp_p.n383 0.04
R10677 vp_p.n382 vp_p.n381 0.04
R10678 vp_p.n380 vp_p.n379 0.04
R10679 vp_p.n378 vp_p.n377 0.04
R10680 vp_p.n376 vp_p.n375 0.04
R10681 vp_p.n374 vp_p.n373 0.04
R10682 vp_p.n371 vp_p.n370 0.04
R10683 vp_p.n369 vp_p.n368 0.04
R10684 vp_p.n367 vp_p.n366 0.04
R10685 vp_p.n365 vp_p.n364 0.04
R10686 vp_p.n363 vp_p.n362 0.04
R10687 vp_p.n361 vp_p.n360 0.04
R10688 vp_p.n359 vp_p.n358 0.04
R10689 vp_p.n357 vp_p.n356 0.04
R10690 vp_p.n355 vp_p.n354 0.04
R10691 vp_p.n353 vp_p.n352 0.04
R10692 vp_p.n351 vp_p.n350 0.04
R10693 vp_p.n349 vp_p.n348 0.04
R10694 vp_p.n347 vp_p.n346 0.04
R10695 vp_p.n345 vp_p.n344 0.04
R10696 vp_p.n343 vp_p.n342 0.04
R10697 vp_p.n341 vp_p.n340 0.04
R10698 vp_p.n339 vp_p.n338 0.04
R10699 vp_p.n337 vp_p.n336 0.04
R10700 vp_p.n335 vp_p.n334 0.04
R10701 vp_p.n333 vp_p.n332 0.04
R10702 vp_p.n331 vp_p.n330 0.04
R10703 vp_p.n329 vp_p.n328 0.04
R10704 vp_p.n327 vp_p.n326 0.04
R10705 vp_p.n325 vp_p.n324 0.04
R10706 vp_p.n323 vp_p.n322 0.04
R10707 vp_p.n321 vp_p.n320 0.04
R10708 vp_p.n319 vp_p.n318 0.04
R10709 vp_p.n317 vp_p.n316 0.04
R10710 vp_p.n315 vp_p.n314 0.04
R10711 vp_p.n313 vp_p.n312 0.04
R10712 vp_p.n311 vp_p.n310 0.04
R10713 vp_p.n309 vp_p.n308 0.04
R10714 vp_p.n307 vp_p.n306 0.04
R10715 vp_p.n305 vp_p.n304 0.04
R10716 vp_p.n303 vp_p.n302 0.04
R10717 vp_p.n301 vp_p.n300 0.04
R10718 vp_p.n299 vp_p.n298 0.04
R10719 vp_p.n297 vp_p.n296 0.04
R10720 vp_p.n295 vp_p.n294 0.04
R10721 vp_p.n293 vp_p.n292 0.04
R10722 vp_p.n291 vp_p.n290 0.04
R10723 vp_p.n289 vp_p.n288 0.04
R10724 vp_p.n287 vp_p.n286 0.04
R10725 vp_p.n285 vp_p.n284 0.04
R10726 vp_p.n283 vp_p.n282 0.04
R10727 vp_p.n281 vp_p.n280 0.04
R10728 vp_p.n279 vp_p.n278 0.04
R10729 vp_p.n277 vp_p.n276 0.04
R10730 vp_p.n275 vp_p.n274 0.04
R10731 vp_p.n273 vp_p.n272 0.04
R10732 vp_p.n271 vp_p.n270 0.04
R10733 vp_p.n269 vp_p.n268 0.04
R10734 vp_p.n267 vp_p.n266 0.04
R10735 vp_p.n265 vp_p.n264 0.04
R10736 vp_p.n263 vp_p.n262 0.04
R10737 vp_p.n261 vp_p.n260 0.04
R10738 vp_p.n259 vp_p.n258 0.04
R10739 vp_p.n257 vp_p.n256 0.04
R10740 vp_p.n255 vp_p.n254 0.04
R10741 vp_p.n253 vp_p.n252 0.04
R10742 vp_p.n251 vp_p.n250 0.04
R10743 vp_p.n249 vp_p.n248 0.04
R10744 vp_p.n247 vp_p.n246 0.04
R10745 vp_p.n245 vp_p.n244 0.04
R10746 vp_p.n243 vp_p.n242 0.04
R10747 vp_p.n241 vp_p.n240 0.04
R10748 vp_p.n239 vp_p.n238 0.04
R10749 vp_p.n237 vp_p.n236 0.04
R10750 vp_p.n235 vp_p.n234 0.04
R10751 vp_p.n233 vp_p.n232 0.04
R10752 vp_p.n231 vp_p.n230 0.04
R10753 vp_p.n229 vp_p.n228 0.04
R10754 vp_p.n227 vp_p.n226 0.04
R10755 vp_p.n225 vp_p.n224 0.04
R10756 vp_p.n222 vp_p.n221 0.04
R10757 vp_p.n220 vp_p.n219 0.04
R10758 vp_p.n218 vp_p.n217 0.04
R10759 vp_p.n216 vp_p.n215 0.04
R10760 vp_p.n214 vp_p.n213 0.04
R10761 vp_p.n212 vp_p.n211 0.04
R10762 vp_p.n210 vp_p.n209 0.04
R10763 vp_p.n208 vp_p.n207 0.04
R10764 vp_p.n206 vp_p.n205 0.04
R10765 vp_p.n204 vp_p.n203 0.04
R10766 vp_p.n202 vp_p.n201 0.04
R10767 vp_p.n200 vp_p.n199 0.04
R10768 vp_p.n198 vp_p.n197 0.04
R10769 vp_p.n196 vp_p.n195 0.04
R10770 vp_p.n194 vp_p.n193 0.04
R10771 vp_p.n192 vp_p.n191 0.04
R10772 vp_p.n190 vp_p.n189 0.04
R10773 vp_p.n188 vp_p.n187 0.04
R10774 vp_p.n186 vp_p.n185 0.04
R10775 vp_p.n184 vp_p.n183 0.04
R10776 vp_p.n182 vp_p.n181 0.04
R10777 vp_p.n180 vp_p.n179 0.04
R10778 vp_p.n178 vp_p.n177 0.04
R10779 vp_p.n176 vp_p.n175 0.04
R10780 vp_p.n174 vp_p.n173 0.04
R10781 vp_p.n172 vp_p.n171 0.04
R10782 vp_p.n170 vp_p.n169 0.04
R10783 vp_p.n168 vp_p.n167 0.04
R10784 vp_p.n166 vp_p.n165 0.04
R10785 vp_p.n164 vp_p.n163 0.04
R10786 vp_p.n162 vp_p.n161 0.04
R10787 vp_p.n160 vp_p.n159 0.04
R10788 vp_p.n158 vp_p.n157 0.04
R10789 vp_p.n156 vp_p.n155 0.04
R10790 vp_p.n154 vp_p.n153 0.04
R10791 vp_p.n152 vp_p.n151 0.04
R10792 vp_p.n150 vp_p.n149 0.04
R10793 vp_p.n148 vp_p.n147 0.04
R10794 vp_p.n146 vp_p.n145 0.04
R10795 vp_p.n144 vp_p.n143 0.04
R10796 vp_p.n142 vp_p.n141 0.04
R10797 vp_p.n140 vp_p.n139 0.04
R10798 vp_p.n138 vp_p.n137 0.04
R10799 vp_p.n136 vp_p.n135 0.04
R10800 vp_p.n134 vp_p.n133 0.04
R10801 vp_p.n132 vp_p.n131 0.04
R10802 vp_p.n130 vp_p.n129 0.04
R10803 vp_p.n128 vp_p.n127 0.04
R10804 vp_p.n126 vp_p.n125 0.04
R10805 vp_p.n124 vp_p.n123 0.04
R10806 vp_p.n122 vp_p.n121 0.04
R10807 vp_p.n120 vp_p.n119 0.04
R10808 vp_p.n118 vp_p.n117 0.04
R10809 vp_p.n116 vp_p.n115 0.04
R10810 vp_p.n114 vp_p.n113 0.04
R10811 vp_p.n112 vp_p.n111 0.04
R10812 vp_p.n110 vp_p.n109 0.04
R10813 vp_p.n108 vp_p.n107 0.04
R10814 vp_p.n106 vp_p.n105 0.04
R10815 vp_p.n104 vp_p.n103 0.04
R10816 vp_p.n102 vp_p.n101 0.04
R10817 vp_p.n100 vp_p.n99 0.04
R10818 vp_p.n98 vp_p.n97 0.04
R10819 vp_p.n96 vp_p.n95 0.04
R10820 vp_p.n94 vp_p.n93 0.04
R10821 vp_p.n92 vp_p.n91 0.04
R10822 vp_p.n90 vp_p.n89 0.04
R10823 vp_p.n88 vp_p.n87 0.04
R10824 vp_p.n86 vp_p.n85 0.04
R10825 vp_p.n84 vp_p.n83 0.04
R10826 vp_p.n82 vp_p.n81 0.04
R10827 vp_p.n80 vp_p.n79 0.04
R10828 vp_p.n78 vp_p.n77 0.04
R10829 vp_p.n76 vp_p.n75 0.04
R10830 vp_p.n971 vp_p.n970 0.04
R10831 vp_p.n969 vp_p.n968 0.04
R10832 vp_p.n967 vp_p.n966 0.04
R10833 vp_p.n965 vp_p.n964 0.04
R10834 vp_p.n963 vp_p.n962 0.04
R10835 vp_p.n961 vp_p.n960 0.04
R10836 vp_p.n959 vp_p.n958 0.04
R10837 vp_p.n957 vp_p.n956 0.04
R10838 vp_p.n955 vp_p.n954 0.04
R10839 vp_p.n953 vp_p.n952 0.04
R10840 vp_p.n951 vp_p.n950 0.04
R10841 vp_p.n949 vp_p.n948 0.04
R10842 vp_p.n947 vp_p.n946 0.04
R10843 vp_p.n945 vp_p.n944 0.04
R10844 vp_p.n943 vp_p.n942 0.04
R10845 vp_p.n941 vp_p.n940 0.04
R10846 vp_p.n939 vp_p.n938 0.04
R10847 vp_p.n937 vp_p.n936 0.04
R10848 vp_p.n935 vp_p.n934 0.04
R10849 vp_p.n933 vp_p.n932 0.04
R10850 vp_p.n931 vp_p.n930 0.04
R10851 vp_p.n929 vp_p.n928 0.04
R10852 vp_p.n927 vp_p.n926 0.04
R10853 vp_p.n925 vp_p.n924 0.04
R10854 vp_p.n923 vp_p.n922 0.04
R10855 vp_p.n921 vp_p.n920 0.04
R10856 vp_p.n919 vp_p.n918 0.04
R10857 vp_p.n917 vp_p.n916 0.04
R10858 vp_p.n915 vp_p.n914 0.04
R10859 vp_p.n913 vp_p.n912 0.04
R10860 vp_p.n911 vp_p.n910 0.04
R10861 vp_p.n909 vp_p.n908 0.04
R10862 vp_p.n907 vp_p.n906 0.04
R10863 vp_p.n905 vp_p.n904 0.04
R10864 vp_p.n903 vp_p.n902 0.04
R10865 vp_p.n901 vp_p.n900 0.04
R10866 vp_p.n899 vp_p.n898 0.04
R10867 vp_p.n897 vp_p.n896 0.04
R10868 vp_p.n895 vp_p.n894 0.04
R10869 vp_p.n893 vp_p.n892 0.04
R10870 vp_p.n891 vp_p.n890 0.04
R10871 vp_p.n889 vp_p.n888 0.04
R10872 vp_p.n887 vp_p.n886 0.04
R10873 vp_p.n885 vp_p.n884 0.04
R10874 vp_p.n883 vp_p.n882 0.04
R10875 vp_p.n881 vp_p.n880 0.04
R10876 vp_p.n879 vp_p.n878 0.04
R10877 vp_p.n877 vp_p.n876 0.04
R10878 vp_p.n875 vp_p.n874 0.04
R10879 vp_p.n873 vp_p.n872 0.04
R10880 vp_p.n871 vp_p.n870 0.04
R10881 vp_p.n869 vp_p.n868 0.04
R10882 vp_p.n867 vp_p.n866 0.04
R10883 vp_p.n865 vp_p.n864 0.04
R10884 vp_p.n863 vp_p.n862 0.04
R10885 vp_p.n861 vp_p.n860 0.04
R10886 vp_p.n859 vp_p.n858 0.04
R10887 vp_p.n857 vp_p.n856 0.04
R10888 vp_p.n855 vp_p.n854 0.04
R10889 vp_p.n853 vp_p.n852 0.04
R10890 vp_p.n851 vp_p.n850 0.04
R10891 vp_p.n849 vp_p.n848 0.04
R10892 vp_p.n847 vp_p.n846 0.04
R10893 vp_p.n845 vp_p.n844 0.04
R10894 vp_p.n843 vp_p.n842 0.04
R10895 vp_p.n841 vp_p.n840 0.04
R10896 vp_p.n839 vp_p.n838 0.04
R10897 vp_p.n837 vp_p.n836 0.04
R10898 vp_p.n835 vp_p.n834 0.04
R10899 vp_p.n833 vp_p.n832 0.04
R10900 vp_p.n831 vp_p.n830 0.04
R10901 vp_p.n829 vp_p.n828 0.04
R10902 vp_p.n827 vp_p.n826 0.04
R10903 vp_p.n825 vp_p.n824 0.04
R10904 vp_p.n1120 vp_p.n1119 0.04
R10905 vp_p.n1118 vp_p.n1117 0.04
R10906 vp_p.n1116 vp_p.n1115 0.04
R10907 vp_p.n1114 vp_p.n1113 0.04
R10908 vp_p.n1112 vp_p.n1111 0.04
R10909 vp_p.n1110 vp_p.n1109 0.04
R10910 vp_p.n1108 vp_p.n1107 0.04
R10911 vp_p.n1106 vp_p.n1105 0.04
R10912 vp_p.n1104 vp_p.n1103 0.04
R10913 vp_p.n1102 vp_p.n1101 0.04
R10914 vp_p.n1100 vp_p.n1099 0.04
R10915 vp_p.n1098 vp_p.n1097 0.04
R10916 vp_p.n1096 vp_p.n1095 0.04
R10917 vp_p.n1094 vp_p.n1093 0.04
R10918 vp_p.n1092 vp_p.n1091 0.04
R10919 vp_p.n1090 vp_p.n1089 0.04
R10920 vp_p.n1088 vp_p.n1087 0.04
R10921 vp_p.n1086 vp_p.n1085 0.04
R10922 vp_p.n1084 vp_p.n1083 0.04
R10923 vp_p.n1082 vp_p.n1081 0.04
R10924 vp_p.n1080 vp_p.n1079 0.04
R10925 vp_p.n1078 vp_p.n1077 0.04
R10926 vp_p.n1076 vp_p.n1075 0.04
R10927 vp_p.n1074 vp_p.n1073 0.04
R10928 vp_p.n1072 vp_p.n1071 0.04
R10929 vp_p.n1070 vp_p.n1069 0.04
R10930 vp_p.n1068 vp_p.n1067 0.04
R10931 vp_p.n1066 vp_p.n1065 0.04
R10932 vp_p.n1064 vp_p.n1063 0.04
R10933 vp_p.n1062 vp_p.n1061 0.04
R10934 vp_p.n1060 vp_p.n1059 0.04
R10935 vp_p.n1058 vp_p.n1057 0.04
R10936 vp_p.n1056 vp_p.n1055 0.04
R10937 vp_p.n1054 vp_p.n1053 0.04
R10938 vp_p.n1052 vp_p.n1051 0.04
R10939 vp_p.n1050 vp_p.n1049 0.04
R10940 vp_p.n1048 vp_p.n1047 0.04
R10941 vp_p.n1046 vp_p.n1045 0.04
R10942 vp_p.n1044 vp_p.n1043 0.04
R10943 vp_p.n1042 vp_p.n1041 0.04
R10944 vp_p.n1040 vp_p.n1039 0.04
R10945 vp_p.n1038 vp_p.n1037 0.04
R10946 vp_p.n1036 vp_p.n1035 0.04
R10947 vp_p.n1034 vp_p.n1033 0.04
R10948 vp_p.n1032 vp_p.n1031 0.04
R10949 vp_p.n1030 vp_p.n1029 0.04
R10950 vp_p.n1028 vp_p.n1027 0.04
R10951 vp_p.n1026 vp_p.n1025 0.04
R10952 vp_p.n1024 vp_p.n1023 0.04
R10953 vp_p.n1022 vp_p.n1021 0.04
R10954 vp_p.n1020 vp_p.n1019 0.04
R10955 vp_p.n1018 vp_p.n1017 0.04
R10956 vp_p.n1016 vp_p.n1015 0.04
R10957 vp_p.n1014 vp_p.n1013 0.04
R10958 vp_p.n1012 vp_p.n1011 0.04
R10959 vp_p.n1010 vp_p.n1009 0.04
R10960 vp_p.n1008 vp_p.n1007 0.04
R10961 vp_p.n1006 vp_p.n1005 0.04
R10962 vp_p.n1004 vp_p.n1003 0.04
R10963 vp_p.n1002 vp_p.n1001 0.04
R10964 vp_p.n1000 vp_p.n999 0.04
R10965 vp_p.n998 vp_p.n997 0.04
R10966 vp_p.n996 vp_p.n995 0.04
R10967 vp_p.n994 vp_p.n993 0.04
R10968 vp_p.n992 vp_p.n991 0.04
R10969 vp_p.n990 vp_p.n989 0.04
R10970 vp_p.n988 vp_p.n987 0.04
R10971 vp_p.n986 vp_p.n985 0.04
R10972 vp_p.n984 vp_p.n983 0.04
R10973 vp_p.n982 vp_p.n981 0.04
R10974 vp_p.n980 vp_p.n979 0.04
R10975 vp_p.n978 vp_p.n977 0.04
R10976 vp_p.n976 vp_p.n975 0.04
R10977 vp_p.n974 vp_p.n973 0.04
R10978 vp_p.n1269 vp_p.n1268 0.04
R10979 vp_p.n1267 vp_p.n1266 0.04
R10980 vp_p.n1265 vp_p.n1264 0.04
R10981 vp_p.n1263 vp_p.n1262 0.04
R10982 vp_p.n1261 vp_p.n1260 0.04
R10983 vp_p.n1259 vp_p.n1258 0.04
R10984 vp_p.n1257 vp_p.n1256 0.04
R10985 vp_p.n1255 vp_p.n1254 0.04
R10986 vp_p.n1253 vp_p.n1252 0.04
R10987 vp_p.n1251 vp_p.n1250 0.04
R10988 vp_p.n1249 vp_p.n1248 0.04
R10989 vp_p.n1247 vp_p.n1246 0.04
R10990 vp_p.n1245 vp_p.n1244 0.04
R10991 vp_p.n1243 vp_p.n1242 0.04
R10992 vp_p.n1241 vp_p.n1240 0.04
R10993 vp_p.n1239 vp_p.n1238 0.04
R10994 vp_p.n1237 vp_p.n1236 0.04
R10995 vp_p.n1235 vp_p.n1234 0.04
R10996 vp_p.n1233 vp_p.n1232 0.04
R10997 vp_p.n1231 vp_p.n1230 0.04
R10998 vp_p.n1229 vp_p.n1228 0.04
R10999 vp_p.n1227 vp_p.n1226 0.04
R11000 vp_p.n1225 vp_p.n1224 0.04
R11001 vp_p.n1223 vp_p.n1222 0.04
R11002 vp_p.n1221 vp_p.n1220 0.04
R11003 vp_p.n1219 vp_p.n1218 0.04
R11004 vp_p.n1217 vp_p.n1216 0.04
R11005 vp_p.n1215 vp_p.n1214 0.04
R11006 vp_p.n1213 vp_p.n1212 0.04
R11007 vp_p.n1211 vp_p.n1210 0.04
R11008 vp_p.n1209 vp_p.n1208 0.04
R11009 vp_p.n1207 vp_p.n1206 0.04
R11010 vp_p.n1205 vp_p.n1204 0.04
R11011 vp_p.n1203 vp_p.n1202 0.04
R11012 vp_p.n1201 vp_p.n1200 0.04
R11013 vp_p.n1199 vp_p.n1198 0.04
R11014 vp_p.n1197 vp_p.n1196 0.04
R11015 vp_p.n1195 vp_p.n1194 0.04
R11016 vp_p.n1193 vp_p.n1192 0.04
R11017 vp_p.n1191 vp_p.n1190 0.04
R11018 vp_p.n1189 vp_p.n1188 0.04
R11019 vp_p.n1187 vp_p.n1186 0.04
R11020 vp_p.n1185 vp_p.n1184 0.04
R11021 vp_p.n1183 vp_p.n1182 0.04
R11022 vp_p.n1181 vp_p.n1180 0.04
R11023 vp_p.n1179 vp_p.n1178 0.04
R11024 vp_p.n1177 vp_p.n1176 0.04
R11025 vp_p.n1175 vp_p.n1174 0.04
R11026 vp_p.n1173 vp_p.n1172 0.04
R11027 vp_p.n1171 vp_p.n1170 0.04
R11028 vp_p.n1169 vp_p.n1168 0.04
R11029 vp_p.n1167 vp_p.n1166 0.04
R11030 vp_p.n1165 vp_p.n1164 0.04
R11031 vp_p.n1163 vp_p.n1162 0.04
R11032 vp_p.n1161 vp_p.n1160 0.04
R11033 vp_p.n1159 vp_p.n1158 0.04
R11034 vp_p.n1157 vp_p.n1156 0.04
R11035 vp_p.n1155 vp_p.n1154 0.04
R11036 vp_p.n1153 vp_p.n1152 0.04
R11037 vp_p.n1151 vp_p.n1150 0.04
R11038 vp_p.n1149 vp_p.n1148 0.04
R11039 vp_p.n1147 vp_p.n1146 0.04
R11040 vp_p.n1145 vp_p.n1144 0.04
R11041 vp_p.n1143 vp_p.n1142 0.04
R11042 vp_p.n1141 vp_p.n1140 0.04
R11043 vp_p.n1139 vp_p.n1138 0.04
R11044 vp_p.n1137 vp_p.n1136 0.04
R11045 vp_p.n1135 vp_p.n1134 0.04
R11046 vp_p.n1133 vp_p.n1132 0.04
R11047 vp_p.n1131 vp_p.n1130 0.04
R11048 vp_p.n1129 vp_p.n1128 0.04
R11049 vp_p.n1127 vp_p.n1126 0.04
R11050 vp_p.n1125 vp_p.n1124 0.04
R11051 vp_p.n1123 vp_p.n1122 0.04
R11052 vp_p.n1418 vp_p.n1417 0.04
R11053 vp_p.n1416 vp_p.n1415 0.04
R11054 vp_p.n1414 vp_p.n1413 0.04
R11055 vp_p.n1412 vp_p.n1411 0.04
R11056 vp_p.n1410 vp_p.n1409 0.04
R11057 vp_p.n1408 vp_p.n1407 0.04
R11058 vp_p.n1406 vp_p.n1405 0.04
R11059 vp_p.n1404 vp_p.n1403 0.04
R11060 vp_p.n1402 vp_p.n1401 0.04
R11061 vp_p.n1400 vp_p.n1399 0.04
R11062 vp_p.n1398 vp_p.n1397 0.04
R11063 vp_p.n1396 vp_p.n1395 0.04
R11064 vp_p.n1394 vp_p.n1393 0.04
R11065 vp_p.n1392 vp_p.n1391 0.04
R11066 vp_p.n1390 vp_p.n1389 0.04
R11067 vp_p.n1388 vp_p.n1387 0.04
R11068 vp_p.n1386 vp_p.n1385 0.04
R11069 vp_p.n1384 vp_p.n1383 0.04
R11070 vp_p.n1382 vp_p.n1381 0.04
R11071 vp_p.n1380 vp_p.n1379 0.04
R11072 vp_p.n1378 vp_p.n1377 0.04
R11073 vp_p.n1376 vp_p.n1375 0.04
R11074 vp_p.n1374 vp_p.n1373 0.04
R11075 vp_p.n1372 vp_p.n1371 0.04
R11076 vp_p.n1370 vp_p.n1369 0.04
R11077 vp_p.n1368 vp_p.n1367 0.04
R11078 vp_p.n1366 vp_p.n1365 0.04
R11079 vp_p.n1364 vp_p.n1363 0.04
R11080 vp_p.n1362 vp_p.n1361 0.04
R11081 vp_p.n1360 vp_p.n1359 0.04
R11082 vp_p.n1358 vp_p.n1357 0.04
R11083 vp_p.n1356 vp_p.n1355 0.04
R11084 vp_p.n1354 vp_p.n1353 0.04
R11085 vp_p.n1352 vp_p.n1351 0.04
R11086 vp_p.n1350 vp_p.n1349 0.04
R11087 vp_p.n1348 vp_p.n1347 0.04
R11088 vp_p.n1346 vp_p.n1345 0.04
R11089 vp_p.n1344 vp_p.n1343 0.04
R11090 vp_p.n1342 vp_p.n1341 0.04
R11091 vp_p.n1340 vp_p.n1339 0.04
R11092 vp_p.n1338 vp_p.n1337 0.04
R11093 vp_p.n1336 vp_p.n1335 0.04
R11094 vp_p.n1334 vp_p.n1333 0.04
R11095 vp_p.n1332 vp_p.n1331 0.04
R11096 vp_p.n1330 vp_p.n1329 0.04
R11097 vp_p.n1328 vp_p.n1327 0.04
R11098 vp_p.n1326 vp_p.n1325 0.04
R11099 vp_p.n1324 vp_p.n1323 0.04
R11100 vp_p.n1322 vp_p.n1321 0.04
R11101 vp_p.n1320 vp_p.n1319 0.04
R11102 vp_p.n1318 vp_p.n1317 0.04
R11103 vp_p.n1316 vp_p.n1315 0.04
R11104 vp_p.n1314 vp_p.n1313 0.04
R11105 vp_p.n1312 vp_p.n1311 0.04
R11106 vp_p.n1310 vp_p.n1309 0.04
R11107 vp_p.n1308 vp_p.n1307 0.04
R11108 vp_p.n1306 vp_p.n1305 0.04
R11109 vp_p.n1304 vp_p.n1303 0.04
R11110 vp_p.n1302 vp_p.n1301 0.04
R11111 vp_p.n1300 vp_p.n1299 0.04
R11112 vp_p.n1298 vp_p.n1297 0.04
R11113 vp_p.n1296 vp_p.n1295 0.04
R11114 vp_p.n1294 vp_p.n1293 0.04
R11115 vp_p.n1292 vp_p.n1291 0.04
R11116 vp_p.n1290 vp_p.n1289 0.04
R11117 vp_p.n1288 vp_p.n1287 0.04
R11118 vp_p.n1286 vp_p.n1285 0.04
R11119 vp_p.n1284 vp_p.n1283 0.04
R11120 vp_p.n1282 vp_p.n1281 0.04
R11121 vp_p.n1280 vp_p.n1279 0.04
R11122 vp_p.n1278 vp_p.n1277 0.04
R11123 vp_p.n1276 vp_p.n1275 0.04
R11124 vp_p.n1274 vp_p.n1273 0.04
R11125 vp_p.n1272 vp_p.n1271 0.04
R11126 vp_p vp_p.n748 0.028
R11127 vp_p vp_p.n745 0.011
R11128 vp_p vp_p.n1497 0.005
R11129 out_p.n828 out_p.t358 8.126
R11130 out_p.n828 out_p.t1164 8.126
R11131 out_p.n829 out_p.t610 8.126
R11132 out_p.n829 out_p.t1284 8.126
R11133 out_p.n830 out_p.t1643 8.126
R11134 out_p.n830 out_p.t763 8.126
R11135 out_p.n831 out_p.t679 8.126
R11136 out_p.n831 out_p.t441 8.126
R11137 out_p.n832 out_p.t1349 8.126
R11138 out_p.n832 out_p.t1546 8.126
R11139 out_p.n833 out_p.t1753 8.126
R11140 out_p.n833 out_p.t476 8.126
R11141 out_p.n834 out_p.t761 8.126
R11142 out_p.n834 out_p.t497 8.126
R11143 out_p.n835 out_p.t525 8.126
R11144 out_p.n835 out_p.t1242 8.126
R11145 out_p.n836 out_p.t1163 8.126
R11146 out_p.n836 out_p.t1365 8.126
R11147 out_p.n837 out_p.t1719 8.126
R11148 out_p.n837 out_p.t332 8.126
R11149 out_p.n839 out_p.t829 8.126
R11150 out_p.n839 out_p.t1091 8.126
R11151 out_p.n840 out_p.t1083 8.126
R11152 out_p.n840 out_p.t845 8.126
R11153 out_p.n841 out_p.t582 8.126
R11154 out_p.n841 out_p.t1438 8.126
R11155 out_p.n842 out_p.t1703 8.126
R11156 out_p.n842 out_p.t774 8.126
R11157 out_p.n843 out_p.t630 8.126
R11158 out_p.n843 out_p.t1146 8.126
R11159 out_p.n844 out_p.t1183 8.126
R11160 out_p.n844 out_p.t1550 8.126
R11161 out_p.n845 out_p.t1744 8.126
R11162 out_p.n845 out_p.t292 8.126
R11163 out_p.n846 out_p.t443 8.126
R11164 out_p.n846 out_p.t755 8.126
R11165 out_p.n847 out_p.t804 8.126
R11166 out_p.n847 out_p.t372 8.126
R11167 out_p.n848 out_p.t1149 8.126
R11168 out_p.n848 out_p.t1513 8.126
R11169 out_p.n850 out_p.t324 8.126
R11170 out_p.n850 out_p.t737 8.126
R11171 out_p.n851 out_p.t1079 8.126
R11172 out_p.n851 out_p.t339 8.126
R11173 out_p.n852 out_p.t1308 8.126
R11174 out_p.n852 out_p.t1503 8.126
R11175 out_p.n853 out_p.t395 8.126
R11176 out_p.n853 out_p.t418 8.126
R11177 out_p.n854 out_p.t465 8.126
R11178 out_p.n854 out_p.t1213 8.126
R11179 out_p.n855 out_p.t1413 8.126
R11180 out_p.n855 out_p.t1622 8.126
R11181 out_p.n856 out_p.t577 8.126
R11182 out_p.n856 out_p.t586 8.126
R11183 out_p.n857 out_p.t1036 8.126
R11184 out_p.n857 out_p.t895 8.126
R11185 out_p.n858 out_p.t752 8.126
R11186 out_p.n858 out_p.t500 8.126
R11187 out_p.n859 out_p.t1382 8.126
R11188 out_p.n859 out_p.t1587 8.126
R11189 out_p.n861 out_p.t1699 8.126
R11190 out_p.n861 out_p.t930 8.126
R11191 out_p.n862 out_p.t667 8.126
R11192 out_p.n862 out_p.t1029 8.126
R11193 out_p.n863 out_p.t897 8.126
R11194 out_p.n863 out_p.t1109 8.126
R11195 out_p.n864 out_p.t1528 8.126
R11196 out_p.n864 out_p.t1736 8.126
R11197 out_p.n865 out_p.t864 8.126
R11198 out_p.n865 out_p.t711 8.126
R11199 out_p.n866 out_p.t474 8.126
R11200 out_p.n866 out_p.t1214 8.126
R11201 out_p.n867 out_p.t1573 8.126
R11202 out_p.n867 out_p.t266 8.126
R11203 out_p.n868 out_p.t974 8.126
R11204 out_p.n868 out_p.t990 8.126
R11205 out_p.n869 out_p.t929 8.126
R11206 out_p.n869 out_p.t934 8.126
R11207 out_p.n870 out_p.t400 8.126
R11208 out_p.n870 out_p.t1181 8.126
R11209 out_p.n872 out_p.t385 8.126
R11210 out_p.n872 out_p.t1492 8.126
R11211 out_p.n873 out_p.t708 8.126
R11212 out_p.n873 out_p.t1626 8.126
R11213 out_p.n874 out_p.t1131 8.126
R11214 out_p.n874 out_p.t597 8.126
R11215 out_p.n875 out_p.t263 8.126
R11216 out_p.n875 out_p.t1328 8.126
R11217 out_p.n876 out_p.t781 8.126
R11218 out_p.n876 out_p.t870 8.126
R11219 out_p.n877 out_p.t1247 8.126
R11220 out_p.n877 out_p.t707 8.126
R11221 out_p.n878 out_p.t1023 8.126
R11222 out_p.n878 out_p.t1373 8.126
R11223 out_p.n879 out_p.t1028 8.126
R11224 out_p.n879 out_p.t1577 8.126
R11225 out_p.n880 out_p.t452 8.126
R11226 out_p.n880 out_p.t1698 8.126
R11227 out_p.n881 out_p.t1211 8.126
R11228 out_p.n881 out_p.t648 8.126
R11229 out_p.n883 out_p.t1523 8.126
R11230 out_p.n883 out_p.t1731 8.126
R11231 out_p.n884 out_p.t1655 8.126
R11232 out_p.n884 out_p.t803 8.126
R11233 out_p.n885 out_p.t1060 8.126
R11234 out_p.n885 out_p.t294 8.126
R11235 out_p.n886 out_p.t1358 8.126
R11236 out_p.n886 out_p.t1561 8.126
R11237 out_p.n887 out_p.t310 8.126
R11238 out_p.n887 out_p.t325 8.126
R11239 out_p.n888 out_p.t777 8.126
R11240 out_p.n888 out_p.t533 8.126
R11241 out_p.n889 out_p.t1399 8.126
R11242 out_p.n889 out_p.t1604 8.126
R11243 out_p.n890 out_p.t1610 8.126
R11244 out_p.n890 out_p.t637 8.126
R11245 out_p.n891 out_p.t1730 8.126
R11246 out_p.n891 out_p.t373 8.126
R11247 out_p.n892 out_p.t696 8.126
R11248 out_p.n892 out_p.t466 8.126
R11249 out_p.n894 out_p.t1598 8.126
R11250 out_p.n894 out_p.t1323 8.126
R11251 out_p.n895 out_p.t1714 8.126
R11252 out_p.n895 out_p.t1452 8.126
R11253 out_p.n896 out_p.t674 8.126
R11254 out_p.n896 out_p.t953 8.126
R11255 out_p.n897 out_p.t1428 8.126
R11256 out_p.n897 out_p.t1155 8.126
R11257 out_p.n898 out_p.t1009 8.126
R11258 out_p.n898 out_p.t1717 8.126
R11259 out_p.n899 out_p.t905 8.126
R11260 out_p.n899 out_p.t335 8.126
R11261 out_p.n900 out_p.t1463 8.126
R11262 out_p.n900 out_p.t1202 8.126
R11263 out_p.n901 out_p.t1677 8.126
R11264 out_p.n901 out_p.t1401 8.126
R11265 out_p.n902 out_p.t1022 8.126
R11266 out_p.n902 out_p.t1522 8.126
R11267 out_p.n903 out_p.t836 8.126
R11268 out_p.n903 out_p.t854 8.126
R11269 out_p.n905 out_p.t1192 8.126
R11270 out_p.n905 out_p.t1393 8.126
R11271 out_p.n906 out_p.t1315 8.126
R11272 out_p.n906 out_p.t1509 8.126
R11273 out_p.n907 out_p.t830 8.126
R11274 out_p.n907 out_p.t818 8.126
R11275 out_p.n908 out_p.t480 8.126
R11276 out_p.n908 out_p.t1228 8.126
R11277 out_p.n909 out_p.t1581 8.126
R11278 out_p.n909 out_p.t989 8.126
R11279 out_p.n910 out_p.t1015 8.126
R11280 out_p.n910 out_p.t1038 8.126
R11281 out_p.n911 out_p.t569 8.126
R11282 out_p.n911 out_p.t1260 8.126
R11283 out_p.n912 out_p.t1269 8.126
R11284 out_p.n912 out_p.t1472 8.126
R11285 out_p.n913 out_p.t1392 8.126
R11286 out_p.n913 out_p.t1597 8.126
R11287 out_p.n914 out_p.t451 8.126
R11288 out_p.n914 out_p.t479 8.126
R11289 out_p.n916 out_p.t640 8.126
R11290 out_p.n916 out_p.t433 8.126
R11291 out_p.n917 out_p.t931 8.126
R11292 out_p.n917 out_p.t1116 8.126
R11293 out_p.n918 out_p.t1468 8.126
R11294 out_p.n918 out_p.t1673 8.126
R11295 out_p.n919 out_p.t928 8.126
R11296 out_p.n919 out_p.t727 8.126
R11297 out_p.n920 out_p.t1177 8.126
R11298 out_p.n920 out_p.t1378 8.126
R11299 out_p.n921 out_p.t1584 8.126
R11300 out_p.n921 out_p.t1011 8.126
R11301 out_p.n922 out_p.t436 8.126
R11302 out_p.n922 out_p.t821 8.126
R11303 out_p.n923 out_p.t815 8.126
R11304 out_p.n923 out_p.t574 8.126
R11305 out_p.n924 out_p.t421 8.126
R11306 out_p.n924 out_p.t1191 8.126
R11307 out_p.n925 out_p.t1543 8.126
R11308 out_p.n925 out_p.t1748 8.126
R11309 out_p.n927 out_p.t492 8.126
R11310 out_p.n927 out_p.t1225 8.126
R11311 out_p.n928 out_p.t1139 8.126
R11312 out_p.n928 out_p.t1343 8.126
R11313 out_p.n929 out_p.t1702 8.126
R11314 out_p.n929 out_p.t283 8.126
R11315 out_p.n930 out_p.t796 8.126
R11316 out_p.n930 out_p.t560 8.126
R11317 out_p.n931 out_p.t1407 8.126
R11318 out_p.n931 out_p.t1615 8.126
R11319 out_p.n932 out_p.t681 8.126
R11320 out_p.n932 out_p.t975 8.126
R11321 out_p.n933 out_p.t892 8.126
R11322 out_p.n933 out_p.t1097 8.126
R11323 out_p.n934 out_p.t1104 8.126
R11324 out_p.n934 out_p.t1305 8.126
R11325 out_p.n935 out_p.t1224 8.126
R11326 out_p.n935 out_p.t1426 8.126
R11327 out_p.n936 out_p.t971 8.126
R11328 out_p.n936 out_p.t997 8.126
R11329 out_p.n938 out_p.t904 8.126
R11330 out_p.n938 out_p.t731 8.126
R11331 out_p.n939 out_p.t1074 8.126
R11332 out_p.n939 out_p.t315 8.126
R11333 out_p.n940 out_p.t1297 8.126
R11334 out_p.n940 out_p.t1497 8.126
R11335 out_p.n941 out_p.t352 8.126
R11336 out_p.n941 out_p.t388 8.126
R11337 out_p.n942 out_p.t446 8.126
R11338 out_p.n942 out_p.t1207 8.126
R11339 out_p.n943 out_p.t1410 8.126
R11340 out_p.n943 out_p.t1618 8.126
R11341 out_p.n944 out_p.t570 8.126
R11342 out_p.n944 out_p.t595 8.126
R11343 out_p.n945 out_p.t572 8.126
R11344 out_p.n945 out_p.t887 8.126
R11345 out_p.n946 out_p.t716 8.126
R11346 out_p.n946 out_p.t482 8.126
R11347 out_p.n947 out_p.t1376 8.126
R11348 out_p.n947 out_p.t1579 8.126
R11349 out_p.n949 out_p.t1567 8.126
R11350 out_p.n949 out_p.t890 8.126
R11351 out_p.n950 out_p.t1685 8.126
R11352 out_p.n950 out_p.t1000 8.126
R11353 out_p.n951 out_p.t624 8.126
R11354 out_p.n951 out_p.t1102 8.126
R11355 out_p.n952 out_p.t1396 8.126
R11356 out_p.n952 out_p.t1725 8.126
R11357 out_p.n953 out_p.t477 8.126
R11358 out_p.n953 out_p.t683 8.126
R11359 out_p.n954 out_p.t862 8.126
R11360 out_p.n954 out_p.t1210 8.126
R11361 out_p.n955 out_p.t1434 8.126
R11362 out_p.n955 out_p.t273 8.126
R11363 out_p.n956 out_p.t1648 8.126
R11364 out_p.n956 out_p.t603 8.126
R11365 out_p.n957 out_p.t269 8.126
R11366 out_p.n957 out_p.t908 8.126
R11367 out_p.n958 out_p.t791 8.126
R11368 out_p.n958 out_p.t1175 8.126
R11369 out_p.n960 out_p.t1166 8.126
R11370 out_p.n960 out_p.t1368 8.126
R11371 out_p.n961 out_p.t1286 8.126
R11372 out_p.n961 out_p.t1484 8.126
R11373 out_p.n962 out_p.t730 8.126
R11374 out_p.n962 out_p.t650 8.126
R11375 out_p.n963 out_p.t440 8.126
R11376 out_p.n963 out_p.t1196 8.126
R11377 out_p.n964 out_p.t1547 8.126
R11378 out_p.n964 out_p.t1750 8.126
R11379 out_p.n965 out_p.t485 8.126
R11380 out_p.n965 out_p.t487 8.126
R11381 out_p.n966 out_p.t518 8.126
R11382 out_p.n966 out_p.t1233 8.126
R11383 out_p.n967 out_p.t1244 8.126
R11384 out_p.n967 out_p.t1445 8.126
R11385 out_p.n968 out_p.t1367 8.126
R11386 out_p.n968 out_p.t1566 8.126
R11387 out_p.n969 out_p.t344 8.126
R11388 out_p.n969 out_p.t397 8.126
R11389 out_p.n10 out_p.t431 8.126
R11390 out_p.n10 out_p.t1194 8.126
R11391 out_p.n11 out_p.t1117 8.126
R11392 out_p.n11 out_p.t1316 8.126
R11393 out_p.n12 out_p.t1675 8.126
R11394 out_p.n12 out_p.t839 8.126
R11395 out_p.n13 out_p.t725 8.126
R11396 out_p.n13 out_p.t489 8.126
R11397 out_p.n14 out_p.t1380 8.126
R11398 out_p.n14 out_p.t1583 8.126
R11399 out_p.n15 out_p.t1005 8.126
R11400 out_p.n15 out_p.t963 8.126
R11401 out_p.n16 out_p.t832 8.126
R11402 out_p.n16 out_p.t568 8.126
R11403 out_p.n17 out_p.t573 8.126
R11404 out_p.n17 out_p.t1271 8.126
R11405 out_p.n18 out_p.t1193 8.126
R11406 out_p.n18 out_p.t1394 8.126
R11407 out_p.n19 out_p.t1749 8.126
R11408 out_p.n19 out_p.t460 8.126
R11409 out_p.n24 out_p.t754 8.126
R11410 out_p.n24 out_p.t651 8.126
R11411 out_p.n25 out_p.t1043 8.126
R11412 out_p.n25 out_p.t915 8.126
R11413 out_p.n26 out_p.t1265 8.126
R11414 out_p.n26 out_p.t1469 8.126
R11415 out_p.n27 out_p.t910 8.126
R11416 out_p.n27 out_p.t924 8.126
R11417 out_p.n28 out_p.t401 8.126
R11418 out_p.n28 out_p.t1179 8.126
R11419 out_p.n29 out_p.t1381 8.126
R11420 out_p.n29 out_p.t1585 8.126
R11421 out_p.n30 out_p.t404 8.126
R11422 out_p.n30 out_p.t486 8.126
R11423 out_p.n31 out_p.t503 8.126
R11424 out_p.n31 out_p.t842 8.126
R11425 out_p.n32 out_p.t668 8.126
R11426 out_p.n32 out_p.t419 8.126
R11427 out_p.n33 out_p.t1347 8.126
R11428 out_p.n33 out_p.t1545 8.126
R11429 out_p.n36 out_p.t461 8.126
R11430 out_p.n36 out_p.t800 8.126
R11431 out_p.n37 out_p.t649 8.126
R11432 out_p.n37 out_p.t982 8.126
R11433 out_p.n38 out_p.t1335 8.126
R11434 out_p.n38 out_p.t556 8.126
R11435 out_p.n39 out_p.t553 8.126
R11436 out_p.n39 out_p.t1692 8.126
R11437 out_p.n40 out_p.t534 8.126
R11438 out_p.n40 out_p.t634 8.126
R11439 out_p.n41 out_p.t1449 8.126
R11440 out_p.n41 out_p.t1180 8.126
R11441 out_p.n42 out_p.t313 8.126
R11442 out_p.n42 out_p.t1742 8.126
R11443 out_p.n43 out_p.t1066 8.126
R11444 out_p.n43 out_p.t426 8.126
R11445 out_p.n44 out_p.t822 8.126
R11446 out_p.n44 out_p.t758 8.126
R11447 out_p.n45 out_p.t1412 8.126
R11448 out_p.n45 out_p.t1144 8.126
R11449 out_p.n48 out_p.t1733 8.126
R11450 out_p.n48 out_p.t383 8.126
R11451 out_p.n49 out_p.t770 8.126
R11452 out_p.n49 out_p.t704 8.126
R11453 out_p.n50 out_p.t319 8.126
R11454 out_p.n50 out_p.t1132 8.126
R11455 out_p.n51 out_p.t1563 8.126
R11456 out_p.n51 out_p.t259 8.126
R11457 out_p.n52 out_p.t363 8.126
R11458 out_p.n52 out_p.t765 8.126
R11459 out_p.n53 out_p.t543 8.126
R11460 out_p.n53 out_p.t1248 8.126
R11461 out_p.n54 out_p.t1605 8.126
R11462 out_p.n54 out_p.t1010 8.126
R11463 out_p.n55 out_p.t660 8.126
R11464 out_p.n55 out_p.t1084 8.126
R11465 out_p.n56 out_p.t396 8.126
R11466 out_p.n56 out_p.t408 8.126
R11467 out_p.n57 out_p.t454 8.126
R11468 out_p.n57 out_p.t1212 8.126
R11469 out_p.n60 out_p.t544 8.126
R11470 out_p.n60 out_p.t1527 8.126
R11471 out_p.n61 out_p.t848 8.126
R11472 out_p.n61 out_p.t1657 8.126
R11473 out_p.n62 out_p.t1169 8.126
R11474 out_p.n62 out_p.t1063 8.126
R11475 out_p.n63 out_p.t1025 8.126
R11476 out_p.n63 out_p.t1362 8.126
R11477 out_p.n64 out_p.t852 8.126
R11478 out_p.n64 out_p.t333 8.126
R11479 out_p.n65 out_p.t1274 8.126
R11480 out_p.n65 out_p.t776 8.126
R11481 out_p.n66 out_p.t688 8.126
R11482 out_p.n66 out_p.t1400 8.126
R11483 out_p.n67 out_p.t627 8.126
R11484 out_p.n67 out_p.t1612 8.126
R11485 out_p.n68 out_p.t547 8.126
R11486 out_p.n68 out_p.t1732 8.126
R11487 out_p.n69 out_p.t1246 8.126
R11488 out_p.n69 out_p.t695 8.126
R11489 out_p.n72 out_p.t1559 8.126
R11490 out_p.n72 out_p.t260 8.126
R11491 out_p.n73 out_p.t1684 8.126
R11492 out_p.n73 out_p.t860 8.126
R11493 out_p.n74 out_p.t945 8.126
R11494 out_p.n74 out_p.t368 8.126
R11495 out_p.n75 out_p.t1388 8.126
R11496 out_p.n75 out_p.t1596 8.126
R11497 out_p.n76 out_p.t424 8.126
R11498 out_p.n76 out_p.t470 8.126
R11499 out_p.n77 out_p.t837 8.126
R11500 out_p.n77 out_p.t591 8.126
R11501 out_p.n78 out_p.t1431 8.126
R11502 out_p.n78 out_p.t1635 8.126
R11503 out_p.n79 out_p.t1642 8.126
R11504 out_p.n79 out_p.t729 8.126
R11505 out_p.n80 out_p.t271 8.126
R11506 out_p.n80 out_p.t545 8.126
R11507 out_p.n81 out_p.t766 8.126
R11508 out_p.n81 out_p.t523 8.126
R11509 out_p.n84 out_p.t1153 8.126
R11510 out_p.n84 out_p.t1356 8.126
R11511 out_p.n85 out_p.t1277 8.126
R11512 out_p.n85 out_p.t1480 8.126
R11513 out_p.n86 out_p.t709 8.126
R11514 out_p.n86 out_p.t644 8.126
R11515 out_p.n87 out_p.t410 8.126
R11516 out_p.n87 out_p.t1188 8.126
R11517 out_p.n88 out_p.t1540 8.126
R11518 out_p.n88 out_p.t1746 8.126
R11519 out_p.n89 out_p.t442 8.126
R11520 out_p.n89 out_p.t520 8.126
R11521 out_p.n90 out_p.t498 8.126
R11522 out_p.n90 out_p.t1231 8.126
R11523 out_p.n91 out_p.t1236 8.126
R11524 out_p.n91 out_p.t1437 8.126
R11525 out_p.n92 out_p.t1355 8.126
R11526 out_p.n92 out_p.t1558 8.126
R11527 out_p.n93 out_p.t297 8.126
R11528 out_p.n93 out_p.t314 8.126
R11529 out_p.n96 out_p.t1227 8.126
R11530 out_p.n96 out_p.t1592 8.126
R11531 out_p.n97 out_p.t1344 8.126
R11532 out_p.n97 out_p.t1710 8.126
R11533 out_p.n98 out_p.t280 8.126
R11534 out_p.n98 out_p.t664 8.126
R11535 out_p.n99 out_p.t549 8.126
R11536 out_p.n99 out_p.t1423 8.126
R11537 out_p.n100 out_p.t1617 8.126
R11538 out_p.n100 out_p.t972 8.126
R11539 out_p.n101 out_p.t993 8.126
R11540 out_p.n101 out_p.t922 8.126
R11541 out_p.n102 out_p.t1100 8.126
R11542 out_p.n102 out_p.t1460 8.126
R11543 out_p.n103 out_p.t1307 8.126
R11544 out_p.n103 out_p.t1671 8.126
R11545 out_p.n104 out_p.t1427 8.126
R11546 out_p.n104 out_p.t973 8.126
R11547 out_p.n105 out_p.t1003 8.126
R11548 out_p.n105 out_p.t826 8.126
R11549 out_p.n108 out_p.t742 8.126
R11550 out_p.n108 out_p.t491 8.126
R11551 out_p.n109 out_p.t328 8.126
R11552 out_p.n109 out_p.t1140 8.126
R11553 out_p.n110 out_p.t1500 8.126
R11554 out_p.n110 out_p.t1705 8.126
R11555 out_p.n111 out_p.t398 8.126
R11556 out_p.n111 out_p.t811 8.126
R11557 out_p.n112 out_p.t1209 8.126
R11558 out_p.n112 out_p.t1409 8.126
R11559 out_p.n113 out_p.t1619 8.126
R11560 out_p.n113 out_p.t655 8.126
R11561 out_p.n114 out_p.t585 8.126
R11562 out_p.n114 out_p.t877 8.126
R11563 out_p.n115 out_p.t912 8.126
R11564 out_p.n115 out_p.t1108 8.126
R11565 out_p.n116 out_p.t481 8.126
R11566 out_p.n116 out_p.t1226 8.126
R11567 out_p.n117 out_p.t1580 8.126
R11568 out_p.n117 out_p.t968 8.126
R11569 out_p.n120 out_p.t539 8.126
R11570 out_p.n120 out_p.t918 8.126
R11571 out_p.n121 out_p.t1171 8.126
R11572 out_p.n121 out_p.t1075 8.126
R11573 out_p.n122 out_p.t1735 8.126
R11574 out_p.n122 out_p.t1302 8.126
R11575 out_p.n123 out_p.t867 8.126
R11576 out_p.n123 out_p.t362 8.126
R11577 out_p.n124 out_p.t1443 8.126
R11578 out_p.n124 out_p.t456 8.126
R11579 out_p.n125 out_p.t740 8.126
R11580 out_p.n125 out_p.t1411 8.126
R11581 out_p.n126 out_p.t288 8.126
R11582 out_p.n126 out_p.t578 8.126
R11583 out_p.n127 out_p.t1130 8.126
R11584 out_p.n127 out_p.t587 8.126
R11585 out_p.n128 out_p.t1257 8.126
R11586 out_p.n128 out_p.t715 8.126
R11587 out_p.n129 out_p.t671 8.126
R11588 out_p.n129 out_p.t1377 8.126
R11589 out_p.n132 out_p.t417 8.126
R11590 out_p.n132 out_p.t785 8.126
R11591 out_p.n133 out_p.t622 8.126
R11592 out_p.n133 out_p.t392 8.126
R11593 out_p.n134 out_p.t1330 8.126
R11594 out_p.n134 out_p.t1530 8.126
R11595 out_p.n135 out_p.t528 8.126
R11596 out_p.n135 out_p.t530 8.126
R11597 out_p.n136 out_p.t526 8.126
R11598 out_p.n136 out_p.t1240 8.126
R11599 out_p.n137 out_p.t1446 8.126
R11600 out_p.n137 out_p.t1649 8.126
R11601 out_p.n138 out_p.t670 8.126
R11602 out_p.n138 out_p.t1052 8.126
R11603 out_p.n139 out_p.t1059 8.126
R11604 out_p.n139 out_p.t308 8.126
R11605 out_p.n140 out_p.t801 8.126
R11606 out_p.n140 out_p.t551 8.126
R11607 out_p.n141 out_p.t1405 8.126
R11608 out_p.n141 out_p.t1613 8.126
R11609 out_p.n144 out_p.t1724 8.126
R11610 out_p.n144 out_p.t365 8.126
R11611 out_p.n145 out_p.t750 8.126
R11612 out_p.n145 out_p.t686 8.126
R11613 out_p.n146 out_p.t285 8.126
R11614 out_p.n146 out_p.t1127 8.126
R11615 out_p.n147 out_p.t1554 8.126
R11616 out_p.n147 out_p.t265 8.126
R11617 out_p.n148 out_p.t366 8.126
R11618 out_p.n148 out_p.t771 8.126
R11619 out_p.n149 out_p.t535 8.126
R11620 out_p.n149 out_p.t1245 8.126
R11621 out_p.n150 out_p.t1602 8.126
R11622 out_p.n150 out_p.t262 8.126
R11623 out_p.n151 out_p.t998 8.126
R11624 out_p.n151 out_p.t954 8.126
R11625 out_p.n152 out_p.t353 8.126
R11626 out_p.n152 out_p.t356 8.126
R11627 out_p.n153 out_p.t457 8.126
R11628 out_p.n153 out_p.t1205 8.126
R11629 out_p.n156 out_p.t995 8.126
R11630 out_p.n156 out_p.t554 8.126
R11631 out_p.n157 out_p.t301 8.126
R11632 out_p.n157 out_p.t689 8.126
R11633 out_p.n158 out_p.t439 8.126
R11634 out_p.n158 out_p.t1360 8.126
R11635 out_p.n159 out_p.t1632 8.126
R11636 out_p.n159 out_p.t1007 8.126
R11637 out_p.n160 out_p.t1035 8.126
R11638 out_p.n160 out_p.t565 8.126
R11639 out_p.n161 out_p.t1112 8.126
R11640 out_p.n161 out_p.t1474 8.126
R11641 out_p.n162 out_p.t1666 8.126
R11642 out_p.n162 out_p.t959 8.126
R11643 out_p.n163 out_p.t863 8.126
R11644 out_p.n163 out_p.t267 8.126
R11645 out_p.n164 out_p.t960 8.126
R11646 out_p.n164 out_p.t857 8.126
R11647 out_p.n165 out_p.t581 8.126
R11648 out_p.n165 out_p.t1440 8.126
R11649 out_p.n168 out_p.t1387 8.126
R11650 out_p.n168 out_p.t1593 8.126
R11651 out_p.n169 out_p.t1506 8.126
R11652 out_p.n169 out_p.t1711 8.126
R11653 out_p.n170 out_p.t798 8.126
R11654 out_p.n170 out_p.t678 8.126
R11655 out_p.n171 out_p.t1222 8.126
R11656 out_p.n171 out_p.t1424 8.126
R11657 out_p.n172 out_p.t977 8.126
R11658 out_p.n172 out_p.t978 8.126
R11659 out_p.n173 out_p.t1032 8.126
R11660 out_p.n173 out_p.t907 8.126
R11661 out_p.n174 out_p.t1259 8.126
R11662 out_p.n174 out_p.t1461 8.126
R11663 out_p.n175 out_p.t1467 8.126
R11664 out_p.n175 out_p.t1672 8.126
R11665 out_p.n176 out_p.t1591 8.126
R11666 out_p.n176 out_p.t966 8.126
R11667 out_p.n177 out_p.t462 8.126
R11668 out_p.n177 out_p.t841 8.126
R11669 out_p.n180 out_p.t1629 8.126
R11670 out_p.n180 out_p.t713 8.126
R11671 out_p.n181 out_p.t1740 8.126
R11672 out_p.n181 out_p.t405 8.126
R11673 out_p.n182 out_p.t741 8.126
R11674 out_p.n182 out_p.t501 8.126
R11675 out_p.n183 out_p.t1457 8.126
R11676 out_p.n183 out_p.t1660 8.126
R11677 out_p.n184 out_p.t584 8.126
R11678 out_p.n184 out_p.t1065 8.126
R11679 out_p.n185 out_p.t305 8.126
R11680 out_p.n185 out_p.t1134 8.126
R11681 out_p.n186 out_p.t1488 8.126
R11682 out_p.n186 out_p.t1691 8.126
R11683 out_p.n187 out_p.t1701 8.126
R11684 out_p.n187 out_p.t937 8.126
R11685 out_p.n188 out_p.t702 8.126
R11686 out_p.n188 out_p.t1031 8.126
R11687 out_p.n189 out_p.t911 8.126
R11688 out_p.n189 out_p.t1111 8.126
R11689 out_p.n192 out_p.t1218 8.126
R11690 out_p.n192 out_p.t1419 8.126
R11691 out_p.n193 out_p.t1337 8.126
R11692 out_p.n193 out_p.t1534 8.126
R11693 out_p.n194 out_p.t900 8.126
R11694 out_p.n194 out_p.t940 8.126
R11695 out_p.n195 out_p.t531 8.126
R11696 out_p.n195 out_p.t1253 8.126
R11697 out_p.n196 out_p.t1608 8.126
R11698 out_p.n196 out_p.t951 8.126
R11699 out_p.n197 out_p.t609 8.126
R11700 out_p.n197 out_p.t1067 8.126
R11701 out_p.n198 out_p.t1094 8.126
R11702 out_p.n198 out_p.t1290 8.126
R11703 out_p.n199 out_p.t1296 8.126
R11704 out_p.n199 out_p.t1495 8.126
R11705 out_p.n200 out_p.t1417 8.126
R11706 out_p.n200 out_p.t1627 8.126
R11707 out_p.n201 out_p.t611 8.126
R11708 out_p.n201 out_p.t605 8.126
R11709 out_p.n204 out_p.t1454 8.126
R11710 out_p.n204 out_p.t473 8.126
R11711 out_p.n205 out_p.t1569 8.126
R11712 out_p.n205 out_p.t1135 8.126
R11713 out_p.n206 out_p.t435 8.126
R11714 out_p.n206 out_p.t1694 8.126
R11715 out_p.n207 out_p.t1281 8.126
R11716 out_p.n207 out_p.t787 8.126
R11717 out_p.n208 out_p.t719 8.126
R11718 out_p.n208 out_p.t1403 8.126
R11719 out_p.n209 out_p.t943 8.126
R11720 out_p.n209 out_p.t647 8.126
R11721 out_p.n210 out_p.t1319 8.126
R11722 out_p.n210 out_p.t881 8.126
R11723 out_p.n211 out_p.t1526 8.126
R11724 out_p.n211 out_p.t1101 8.126
R11725 out_p.n212 out_p.t1656 8.126
R11726 out_p.n212 out_p.t1217 8.126
R11727 out_p.n213 out_p.t1062 8.126
R11728 out_p.n213 out_p.t983 8.126
R11729 out_p.n216 out_p.t871 8.126
R11730 out_p.n216 out_p.t1250 8.126
R11731 out_p.n217 out_p.t438 8.126
R11732 out_p.n217 out_p.t1370 8.126
R11733 out_p.n218 out_p.t1562 8.126
R11734 out_p.n218 out_p.t375 8.126
R11735 out_p.n219 out_p.t1047 8.126
R11736 out_p.n219 out_p.t601 8.126
R11737 out_p.n220 out_p.t1268 8.126
R11738 out_p.n220 out_p.t1639 8.126
R11739 out_p.n221 out_p.t1678 8.126
R11740 out_p.n221 out_p.t639 8.126
R11741 out_p.n222 out_p.t1093 8.126
R11742 out_p.n222 out_p.t1120 8.126
R11743 out_p.n223 out_p.t382 8.126
R11744 out_p.n223 out_p.t1327 8.126
R11745 out_p.n224 out_p.t608 8.126
R11746 out_p.n224 out_p.t1453 8.126
R11747 out_p.n225 out_p.t1646 8.126
R11748 out_p.n225 out_p.t604 8.126
R11749 out_p.n228 out_p.t511 8.126
R11750 out_p.n228 out_p.t513 8.126
R11751 out_p.n229 out_p.t828 8.126
R11752 out_p.n229 out_p.t673 8.126
R11753 out_p.n230 out_p.t1158 8.126
R11754 out_p.n230 out_p.t1361 8.126
R11755 out_p.n231 out_p.t992 8.126
R11756 out_p.n231 out_p.t1013 8.126
R11757 out_p.n232 out_p.t831 8.126
R11758 out_p.n232 out_p.t575 8.126
R11759 out_p.n233 out_p.t1272 8.126
R11760 out_p.n233 out_p.t1475 8.126
R11761 out_p.n234 out_p.t677 8.126
R11762 out_p.n234 out_p.t955 8.126
R11763 out_p.n235 out_p.t615 8.126
R11764 out_p.n235 out_p.t948 8.126
R11765 out_p.n236 out_p.t504 8.126
R11766 out_p.n236 out_p.t856 8.126
R11767 out_p.n237 out_p.t1237 8.126
R11768 out_p.n237 out_p.t1441 8.126
R11769 out_p.n240 out_p.t1042 8.126
R11770 out_p.n240 out_p.t925 8.126
R11771 out_p.n241 out_p.t735 8.126
R11772 out_p.n241 out_p.t499 8.126
R11773 out_p.n242 out_p.t1390 8.126
R11774 out_p.n242 out_p.t1595 8.126
R11775 out_p.n243 out_p.t1018 8.126
R11776 out_p.n243 out_p.t1078 8.126
R11777 out_p.n244 out_p.t1105 8.126
R11778 out_p.n244 out_p.t1304 8.126
R11779 out_p.n245 out_p.t1502 8.126
R11780 out_p.n245 out_p.t1707 8.126
R11781 out_p.n246 out_p.t724 8.126
R11782 out_p.n246 out_p.t646 8.126
R11783 out_p.n247 out_p.t652 8.126
R11784 out_p.n247 out_p.t432 8.126
R11785 out_p.n248 out_p.t927 8.126
R11786 out_p.n248 out_p.t1118 8.126
R11787 out_p.n249 out_p.t1470 8.126
R11788 out_p.n249 out_p.t1676 8.126
R11789 out_p.n252 out_p.t999 8.126
R11790 out_p.n252 out_p.t976 8.126
R11791 out_p.n253 out_p.t291 8.126
R11792 out_p.n253 out_p.t274 8.126
R11793 out_p.n254 out_p.t423 8.126
R11794 out_p.n254 out_p.t1187 8.126
R11795 out_p.n255 out_p.t1621 8.126
R11796 out_p.n255 out_p.t656 8.126
R11797 out_p.n256 out_p.t614 8.126
R11798 out_p.n256 out_p.t902 8.126
R11799 out_p.n257 out_p.t1107 8.126
R11800 out_p.n257 out_p.t1306 8.126
R11801 out_p.n258 out_p.t1662 8.126
R11802 out_p.n258 out_p.t789 8.126
R11803 out_p.n259 out_p.t819 8.126
R11804 out_p.n259 out_p.t778 8.126
R11805 out_p.n260 out_p.t970 8.126
R11806 out_p.n260 out_p.t1041 8.126
R11807 out_p.n261 out_p.t567 8.126
R11808 out_p.n261 out_p.t1264 8.126
R11809 out_p.n264 out_p.t1420 8.126
R11810 out_p.n264 out_p.t1588 8.126
R11811 out_p.n265 out_p.t1535 8.126
R11812 out_p.n265 out_p.t1708 8.126
R11813 out_p.n266 out_p.t936 8.126
R11814 out_p.n266 out_p.t642 8.126
R11815 out_p.n267 out_p.t1255 8.126
R11816 out_p.n267 out_p.t1414 8.126
R11817 out_p.n268 out_p.t950 8.126
R11818 out_p.n268 out_p.t593 8.126
R11819 out_p.n269 out_p.t1069 8.126
R11820 out_p.n269 out_p.t896 8.126
R11821 out_p.n270 out_p.t1291 8.126
R11822 out_p.n270 out_p.t1458 8.126
R11823 out_p.n271 out_p.t1496 8.126
R11824 out_p.n271 out_p.t1668 8.126
R11825 out_p.n272 out_p.t1628 8.126
R11826 out_p.n272 out_p.t1002 8.126
R11827 out_p.n273 out_p.t1033 8.126
R11828 out_p.n273 out_p.t817 8.126
R11829 out_p.n276 out_p.t797 8.126
R11830 out_p.n276 out_p.t1219 8.126
R11831 out_p.n277 out_p.t378 8.126
R11832 out_p.n277 out_p.t1338 8.126
R11833 out_p.n278 out_p.t1532 8.126
R11834 out_p.n278 out_p.t909 8.126
R11835 out_p.n279 out_p.t538 8.126
R11836 out_p.n279 out_p.t541 8.126
R11837 out_p.n280 out_p.t1243 8.126
R11838 out_p.n280 out_p.t1609 8.126
R11839 out_p.n281 out_p.t1650 8.126
R11840 out_p.n281 out_p.t1087 8.126
R11841 out_p.n282 out_p.t1054 8.126
R11842 out_p.n282 out_p.t1090 8.126
R11843 out_p.n283 out_p.t307 8.126
R11844 out_p.n283 out_p.t1300 8.126
R11845 out_p.n284 out_p.t550 8.126
R11846 out_p.n284 out_p.t1418 8.126
R11847 out_p.n285 out_p.t1614 8.126
R11848 out_p.n285 out_p.t1026 8.126
R11849 out_p.n288 out_p.t606 8.126
R11850 out_p.n288 out_p.t377 8.126
R11851 out_p.n289 out_p.t1200 8.126
R11852 out_p.n289 out_p.t621 8.126
R11853 out_p.n290 out_p.t1020 8.126
R11854 out_p.n290 out_p.t1332 8.126
R11855 out_p.n291 out_p.t279 8.126
R11856 out_p.n291 out_p.t536 8.126
R11857 out_p.n292 out_p.t1473 8.126
R11858 out_p.n292 out_p.t514 8.126
R11859 out_p.n293 out_p.t849 8.126
R11860 out_p.n293 out_p.t1447 8.126
R11861 out_p.n294 out_p.t349 8.126
R11862 out_p.n294 out_p.t303 8.126
R11863 out_p.n295 out_p.t1168 8.126
R11864 out_p.n295 out_p.t1061 8.126
R11865 out_p.n296 out_p.t1287 8.126
R11866 out_p.n296 out_p.t812 8.126
R11867 out_p.n297 out_p.t773 8.126
R11868 out_p.n297 out_p.t1406 8.126
R11869 out_p.n300 out_p.t571 8.126
R11870 out_p.n300 out_p.t882 8.126
R11871 out_p.n301 out_p.t701 8.126
R11872 out_p.n301 out_p.t449 8.126
R11873 out_p.n302 out_p.t1364 8.126
R11874 out_p.n302 out_p.t1564 8.126
R11875 out_p.n303 out_p.t1021 8.126
R11876 out_p.n303 out_p.t1049 8.126
R11877 out_p.n304 out_p.t583 8.126
R11878 out_p.n304 out_p.t1270 8.126
R11879 out_p.n305 out_p.t1476 8.126
R11880 out_p.n305 out_p.t1679 8.126
R11881 out_p.n306 out_p.t958 8.126
R11882 out_p.n306 out_p.t1085 8.126
R11883 out_p.n307 out_p.t947 8.126
R11884 out_p.n307 out_p.t381 8.126
R11885 out_p.n308 out_p.t855 8.126
R11886 out_p.n308 out_p.t607 8.126
R11887 out_p.n309 out_p.t1442 8.126
R11888 out_p.n309 out_p.t1647 8.126
R11889 out_p.n312 out_p.t1756 8.126
R11890 out_p.n312 out_p.t510 8.126
R11891 out_p.n313 out_p.t859 8.126
R11892 out_p.n313 out_p.t834 8.126
R11893 out_p.n314 out_p.t348 8.126
R11894 out_p.n314 out_p.t1162 8.126
R11895 out_p.n315 out_p.t1589 8.126
R11896 out_p.n315 out_p.t979 8.126
R11897 out_p.n316 out_p.t453 8.126
R11898 out_p.n316 out_p.t827 8.126
R11899 out_p.n317 out_p.t592 8.126
R11900 out_p.n317 out_p.t1273 8.126
R11901 out_p.n318 out_p.t1634 8.126
R11902 out_p.n318 out_p.t687 8.126
R11903 out_p.n319 out_p.t699 8.126
R11904 out_p.n319 out_p.t631 8.126
R11905 out_p.n320 out_p.t502 8.126
R11906 out_p.n320 out_p.t521 8.126
R11907 out_p.n321 out_p.t505 8.126
R11908 out_p.n321 out_p.t1238 8.126
R11909 out_p.n324 out_p.t994 8.126
R11910 out_p.n324 out_p.t1046 8.126
R11911 out_p.n325 out_p.t275 8.126
R11912 out_p.n325 out_p.t762 8.126
R11913 out_p.n326 out_p.t1189 8.126
R11914 out_p.n326 out_p.t1391 8.126
R11915 out_p.n327 out_p.t703 8.126
R11916 out_p.n327 out_p.t967 8.126
R11917 out_p.n328 out_p.t901 8.126
R11918 out_p.n328 out_p.t1106 8.126
R11919 out_p.n329 out_p.t1309 8.126
R11920 out_p.n329 out_p.t1504 8.126
R11921 out_p.n330 out_p.t823 8.126
R11922 out_p.n330 out_p.t734 8.126
R11923 out_p.n331 out_p.t788 8.126
R11924 out_p.n331 out_p.t665 8.126
R11925 out_p.n332 out_p.t1044 8.126
R11926 out_p.n332 out_p.t926 8.126
R11927 out_p.n333 out_p.t1266 8.126
R11928 out_p.n333 out_p.t1471 8.126
R11929 out_p.n336 out_p.t1422 8.126
R11930 out_p.n336 out_p.t996 8.126
R11931 out_p.n337 out_p.t1536 8.126
R11932 out_p.n337 out_p.t302 8.126
R11933 out_p.n338 out_p.t935 8.126
R11934 out_p.n338 out_p.t422 8.126
R11935 out_p.n339 out_p.t1256 8.126
R11936 out_p.n339 out_p.t1625 8.126
R11937 out_p.n340 out_p.t661 8.126
R11938 out_p.n340 out_p.t612 8.126
R11939 out_p.n341 out_p.t1070 8.126
R11940 out_p.n341 out_p.t1110 8.126
R11941 out_p.n342 out_p.t1292 8.126
R11942 out_p.n342 out_p.t1663 8.126
R11943 out_p.n343 out_p.t1499 8.126
R11944 out_p.n343 out_p.t853 8.126
R11945 out_p.n344 out_p.t1630 8.126
R11946 out_p.n344 out_p.t988 8.126
R11947 out_p.n345 out_p.t1034 8.126
R11948 out_p.n345 out_p.t566 8.126
R11949 out_p.n348 out_p.t1659 8.126
R11950 out_p.n348 out_p.t1221 8.126
R11951 out_p.n349 out_p.t270 8.126
R11952 out_p.n349 out_p.t1340 8.126
R11953 out_p.n350 out_p.t795 8.126
R11954 out_p.n350 out_p.t920 8.126
R11955 out_p.n351 out_p.t1483 8.126
R11956 out_p.n351 out_p.t540 8.126
R11957 out_p.n352 out_p.t643 8.126
R11958 out_p.n352 out_p.t1611 8.126
R11959 out_p.n353 out_p.t380 8.126
R11960 out_p.n353 out_p.t1030 8.126
R11961 out_p.n354 out_p.t1517 8.126
R11962 out_p.n354 out_p.t946 8.126
R11963 out_p.n355 out_p.t1734 8.126
R11964 out_p.n355 out_p.t1301 8.126
R11965 out_p.n356 out_p.t779 8.126
R11966 out_p.n356 out_p.t1421 8.126
R11967 out_p.n357 out_p.t318 8.126
R11968 out_p.n357 out_p.t965 8.126
R11969 out_p.n360 out_p.t1252 8.126
R11970 out_p.n360 out_p.t1456 8.126
R11971 out_p.n361 out_p.t1371 8.126
R11972 out_p.n361 out_p.t1570 8.126
R11973 out_p.n362 out_p.t374 8.126
R11974 out_p.n362 out_p.t444 8.126
R11975 out_p.n363 out_p.t600 8.126
R11976 out_p.n363 out_p.t1283 8.126
R11977 out_p.n364 out_p.t1641 8.126
R11978 out_p.n364 out_p.t720 8.126
R11979 out_p.n365 out_p.t654 8.126
R11980 out_p.n365 out_p.t942 8.126
R11981 out_p.n366 out_p.t1121 8.126
R11982 out_p.n366 out_p.t1320 8.126
R11983 out_p.n367 out_p.t1329 8.126
R11984 out_p.n367 out_p.t1529 8.126
R11985 out_p.n368 out_p.t1455 8.126
R11986 out_p.n368 out_p.t1658 8.126
R11987 out_p.n369 out_p.t594 8.126
R11988 out_p.n369 out_p.t1064 8.126
R11989 out_p.n372 out_p.t775 8.126
R11990 out_p.n372 out_p.t542 8.126
R11991 out_p.n373 out_p.t393 8.126
R11992 out_p.n373 out_p.t1170 8.126
R11993 out_p.n374 out_p.t1519 8.126
R11994 out_p.n374 out_p.t1727 8.126
R11995 out_p.n375 out_p.t546 8.126
R11996 out_p.n375 out_p.t861 8.126
R11997 out_p.n376 out_p.t1235 8.126
R11998 out_p.n376 out_p.t1436 8.126
R11999 out_p.n377 out_p.t1645 8.126
R12000 out_p.n377 out_p.t739 8.126
R12001 out_p.n378 out_p.t1051 8.126
R12002 out_p.n378 out_p.t277 8.126
R12003 out_p.n379 out_p.t957 8.126
R12004 out_p.n379 out_p.t1126 8.126
R12005 out_p.n380 out_p.t532 8.126
R12006 out_p.n380 out_p.t1251 8.126
R12007 out_p.n381 out_p.t1606 8.126
R12008 out_p.n381 out_p.t991 8.126
R12009 out_p.n384 out_p.t602 8.126
R12010 out_p.n384 out_p.t1280 8.126
R12011 out_p.n385 out_p.t1198 8.126
R12012 out_p.n385 out_p.t1397 8.126
R12013 out_p.n386 out_p.t261 8.126
R12014 out_p.n386 out_p.t527 8.126
R12015 out_p.n387 out_p.t917 8.126
R12016 out_p.n387 out_p.t1115 8.126
R12017 out_p.n388 out_p.t1465 8.126
R12018 out_p.n388 out_p.t1670 8.126
R12019 out_p.n389 out_p.t873 8.126
R12020 out_p.n389 out_p.t814 8.126
R12021 out_p.n390 out_p.t338 8.126
R12022 out_p.n390 out_p.t1150 8.126
R12023 out_p.n391 out_p.t1156 8.126
R12024 out_p.n391 out_p.t1359 8.126
R12025 out_p.n392 out_p.t1278 8.126
R12026 out_p.n392 out_p.t1481 8.126
R12027 out_p.n393 out_p.t743 8.126
R12028 out_p.n393 out_p.t659 8.126
R12029 out_p.n396 out_p.t1001 8.126
R12030 out_p.n396 out_p.t835 8.126
R12031 out_p.n397 out_p.t334 8.126
R12032 out_p.n397 out_p.t450 8.126
R12033 out_p.n398 out_p.t1190 8.126
R12034 out_p.n398 out_p.t1557 8.126
R12035 out_p.n399 out_p.t676 8.126
R12036 out_p.n399 out_p.t1040 8.126
R12037 out_p.n400 out_p.t885 8.126
R12038 out_p.n400 out_p.t1263 8.126
R12039 out_p.n401 out_p.t1310 8.126
R12040 out_p.n401 out_p.t1674 8.126
R12041 out_p.n402 out_p.t790 8.126
R12042 out_p.n402 out_p.t1089 8.126
R12043 out_p.n403 out_p.t784 8.126
R12044 out_p.n403 out_p.t361 8.126
R12045 out_p.n404 out_p.t1045 8.126
R12046 out_p.n404 out_p.t590 8.126
R12047 out_p.n405 out_p.t1267 8.126
R12048 out_p.n405 out_p.t1638 8.126
R12049 out_p.n408 out_p.t1077 8.126
R12050 out_p.n408 out_p.t327 8.126
R12051 out_p.n409 out_p.t806 8.126
R12052 out_p.n409 out_p.t548 8.126
R12053 out_p.n410 out_p.t1425 8.126
R12054 out_p.n410 out_p.t1631 8.126
R12055 out_p.n411 out_p.t693 8.126
R12056 out_p.n411 out_p.t618 8.126
R12057 out_p.n412 out_p.t1129 8.126
R12058 out_p.n412 out_p.t1334 8.126
R12059 out_p.n413 out_p.t1533 8.126
R12060 out_p.n413 out_p.t1738 8.126
R12061 out_p.n414 out_p.t888 8.126
R12062 out_p.n414 out_p.t706 8.126
R12063 out_p.n415 out_p.t726 8.126
R12064 out_p.n415 out_p.t490 8.126
R12065 out_p.n416 out_p.t340 8.126
R12066 out_p.n416 out_p.t1141 8.126
R12067 out_p.n417 out_p.t1501 8.126
R12068 out_p.n417 out_p.t1706 8.126
R12069 out_p.n420 out_p.t692 8.126
R12070 out_p.n420 out_p.t1012 8.126
R12071 out_p.n421 out_p.t394 8.126
R12072 out_p.n421 out_p.t428 8.126
R12073 out_p.n422 out_p.t483 8.126
R12074 out_p.n422 out_p.t1223 8.126
R12075 out_p.n423 out_p.t1654 8.126
R12076 out_p.n423 out_p.t769 8.126
R12077 out_p.n424 out_p.t1058 8.126
R12078 out_p.n424 out_p.t295 8.126
R12079 out_p.n425 out_p.t1133 8.126
R12080 out_p.n425 out_p.t1336 8.126
R12081 out_p.n426 out_p.t1688 8.126
R12082 out_p.n426 out_p.t880 8.126
R12083 out_p.n427 out_p.t933 8.126
R12084 out_p.n427 out_p.t939 8.126
R12085 out_p.n428 out_p.t1006 8.126
R12086 out_p.n428 out_p.t1076 8.126
R12087 out_p.n429 out_p.t1103 8.126
R12088 out_p.n429 out_p.t1303 8.126
R12089 out_p.n432 out_p.t697 8.126
R12090 out_p.n432 out_p.t1620 8.126
R12091 out_p.n433 out_p.t596 8.126
R12092 out_p.n433 out_p.t1739 8.126
R12093 out_p.n434 out_p.t1254 8.126
R12094 out_p.n434 out_p.t717 8.126
R12095 out_p.n435 out_p.t893 8.126
R12096 out_p.n435 out_p.t1451 8.126
R12097 out_p.n436 out_p.t370 8.126
R12098 out_p.n436 out_p.t298 8.126
R12099 out_p.n437 out_p.t1369 8.126
R12100 out_p.n437 out_p.t306 8.126
R12101 out_p.n438 out_p.t331 8.126
R12102 out_p.n438 out_p.t1486 8.126
R12103 out_p.n439 out_p.t427 8.126
R12104 out_p.n439 out_p.t1693 8.126
R12105 out_p.n440 out_p.t619 8.126
R12106 out_p.n440 out_p.t680 8.126
R12107 out_p.n441 out_p.t1333 8.126
R12108 out_p.n441 out_p.t875 8.126
R12109 out_p.n444 out_p.t1652 8.126
R12110 out_p.n444 out_p.t793 8.126
R12111 out_p.n445 out_p.t257 8.126
R12112 out_p.n445 out_p.t562 8.126
R12113 out_p.n446 out_p.t802 8.126
R12114 out_p.n446 out_p.t552 8.126
R12115 out_p.n447 out_p.t1479 8.126
R12116 out_p.n447 out_p.t1683 8.126
R12117 out_p.n448 out_p.t632 8.126
R12118 out_p.n448 out_p.t1027 8.126
R12119 out_p.n449 out_p.t369 8.126
R12120 out_p.n449 out_p.t1167 8.126
R12121 out_p.n450 out_p.t1515 8.126
R12122 out_p.n450 out_p.t1721 8.126
R12123 out_p.n451 out_p.t1726 8.126
R12124 out_p.n451 out_p.t364 8.126
R12125 out_p.n452 out_p.t759 8.126
R12126 out_p.n452 out_p.t682 8.126
R12127 out_p.n453 out_p.t296 8.126
R12128 out_p.n453 out_p.t1128 8.126
R12129 out_p.n456 out_p.t589 8.126
R12130 out_p.n456 out_p.t1448 8.126
R12131 out_p.n457 out_p.t1199 8.126
R12132 out_p.n457 out_p.t1568 8.126
R12133 out_p.n458 out_p.t272 8.126
R12134 out_p.n458 out_p.t346 8.126
R12135 out_p.n459 out_p.t916 8.126
R12136 out_p.n459 out_p.t1276 8.126
R12137 out_p.n460 out_p.t1466 8.126
R12138 out_p.n460 out_p.t733 8.126
R12139 out_p.n461 out_p.t840 8.126
R12140 out_p.n461 out_p.t944 8.126
R12141 out_p.n462 out_p.t351 8.126
R12142 out_p.n462 out_p.t1318 8.126
R12143 out_p.n463 out_p.t1157 8.126
R12144 out_p.n463 out_p.t1518 8.126
R12145 out_p.n464 out_p.t1279 8.126
R12146 out_p.n464 out_p.t1651 8.126
R12147 out_p.n465 out_p.t710 8.126
R12148 out_p.n465 out_p.t1055 8.126
R12149 out_p.n468 out_p.t1314 8.126
R12150 out_p.n468 out_p.t1508 8.126
R12151 out_p.n469 out_p.t1429 8.126
R12152 out_p.n469 out_p.t1633 8.126
R12153 out_p.n470 out_p.t1019 8.126
R12154 out_p.n470 out_p.t1048 8.126
R12155 out_p.n471 out_p.t1138 8.126
R12156 out_p.n471 out_p.t1342 8.126
R12157 out_p.n472 out_p.t1700 8.126
R12158 out_p.n472 out_p.t938 8.126
R12159 out_p.n473 out_p.t300 8.126
R12160 out_p.n473 out_p.t736 8.126
R12161 out_p.n474 out_p.t1182 8.126
R12162 out_p.n474 out_p.t1383 8.126
R12163 out_p.n475 out_p.t1389 8.126
R12164 out_p.n475 out_p.t1594 8.126
R12165 out_p.n476 out_p.t1507 8.126
R12166 out_p.n476 out_p.t1712 8.126
R12167 out_p.n477 out_p.t808 8.126
R12168 out_p.n477 out_p.t675 8.126
R12169 out_p.n480 out_p.t921 8.126
R12170 out_p.n480 out_p.t1114 8.126
R12171 out_p.n481 out_p.t488 8.126
R12172 out_p.n481 out_p.t1229 8.126
R12173 out_p.n482 out_p.t1590 8.126
R12174 out_p.n482 out_p.t1014 8.126
R12175 out_p.n483 out_p.t1073 8.126
R12176 out_p.n483 out_p.t329 8.126
R12177 out_p.n484 out_p.t1299 8.126
R12178 out_p.n484 out_p.t1494 8.126
R12179 out_p.n485 out_p.t1704 8.126
R12180 out_p.n485 out_p.t281 8.126
R12181 out_p.n486 out_p.t629 8.126
R12182 out_p.n486 out_p.t412 8.126
R12183 out_p.n487 out_p.t411 8.126
R12184 out_p.n487 out_p.t1186 8.126
R12185 out_p.n488 out_p.t1113 8.126
R12186 out_p.n488 out_p.t1313 8.126
R12187 out_p.n489 out_p.t1669 8.126
R12188 out_p.n489 out_p.t820 8.126
R12189 out_p.n492 out_p.t1137 8.126
R12190 out_p.n492 out_p.t1037 8.126
R12191 out_p.n493 out_p.t1258 8.126
R12192 out_p.n493 out_p.t751 8.126
R12193 out_p.n494 out_p.t691 8.126
R12194 out_p.n494 out_p.t1384 8.126
R12195 out_p.n495 out_p.t379 8.126
R12196 out_p.n495 out_p.t987 8.126
R12197 out_p.n496 out_p.t1525 8.126
R12198 out_p.n496 out_p.t1099 8.126
R12199 out_p.n497 out_p.t406 8.126
R12200 out_p.n497 out_p.t1498 8.126
R12201 out_p.n498 out_p.t464 8.126
R12202 out_p.n498 out_p.t728 8.126
R12203 out_p.n499 out_p.t1220 8.126
R12204 out_p.n499 out_p.t658 8.126
R12205 out_p.n500 out_p.t1339 8.126
R12206 out_p.n500 out_p.t906 8.126
R12207 out_p.n501 out_p.t941 8.126
R12208 out_p.n501 out_p.t1462 8.126
R12209 out_p.n504 out_p.t1068 8.126
R12210 out_p.n504 out_p.t330 8.126
R12211 out_p.n505 out_p.t807 8.126
R12212 out_p.n505 out_p.t559 8.126
R12213 out_p.n506 out_p.t1416 8.126
R12214 out_p.n506 out_p.t1624 8.126
R12215 out_p.n507 out_p.t672 8.126
R12216 out_p.n507 out_p.t636 8.126
R12217 out_p.n508 out_p.t1125 8.126
R12218 out_p.n508 out_p.t1326 8.126
R12219 out_p.n509 out_p.t1531 8.126
R12220 out_p.n509 out_p.t1737 8.126
R12221 out_p.n510 out_p.t874 8.126
R12222 out_p.n510 out_p.t722 8.126
R12223 out_p.n511 out_p.t721 8.126
R12224 out_p.n511 out_p.t472 8.126
R12225 out_p.n512 out_p.t317 8.126
R12226 out_p.n512 out_p.t1136 8.126
R12227 out_p.n513 out_p.t1490 8.126
R12228 out_p.n513 out_p.t1696 8.126
R12229 out_p.n516 out_p.t684 8.126
R12230 out_p.n516 out_p.t969 8.126
R12231 out_p.n517 out_p.t278 8.126
R12232 out_p.n517 out_p.t469 8.126
R12233 out_p.n518 out_p.t1482 8.126
R12234 out_p.n518 out_p.t1216 8.126
R12235 out_p.n519 out_p.t345 8.126
R12236 out_p.n519 out_p.t783 8.126
R12237 out_p.n520 out_p.t1195 8.126
R12238 out_p.n520 out_p.t286 8.126
R12239 out_p.n521 out_p.t1599 8.126
R12240 out_p.n521 out_p.t1331 8.126
R12241 out_p.n522 out_p.t529 8.126
R12242 out_p.n522 out_p.t913 8.126
R12243 out_p.n523 out_p.t866 8.126
R12244 out_p.n523 out_p.t884 8.126
R12245 out_p.n524 out_p.t448 8.126
R12246 out_p.n524 out_p.t1071 8.126
R12247 out_p.n525 out_p.t1565 8.126
R12248 out_p.n525 out_p.t1294 8.126
R12249 out_p.n528 out_p.t850 8.126
R12250 out_p.n528 out_p.t838 8.126
R12251 out_p.n529 out_p.t952 8.126
R12252 out_p.n529 out_p.t1050 8.126
R12253 out_p.n530 out_p.t599 8.126
R12254 out_p.n530 out_p.t1285 8.126
R12255 out_p.n531 out_p.t1709 8.126
R12256 out_p.n531 out_p.t290 8.126
R12257 out_p.n532 out_p.t653 8.126
R12258 out_p.n532 out_p.t430 8.126
R12259 out_p.n533 out_p.t1197 8.126
R12260 out_p.n533 out_p.t1395 8.126
R12261 out_p.n534 out_p.t1752 8.126
R12262 out_p.n534 out_p.t468 8.126
R12263 out_p.n535 out_p.t519 8.126
R12264 out_p.n535 out_p.t563 8.126
R12265 out_p.n536 out_p.t824 8.126
R12266 out_p.n536 out_p.t685 8.126
R12267 out_p.n537 out_p.t1160 8.126
R12268 out_p.n537 out_p.t1366 8.126
R12269 out_p.n540 out_p.t1477 8.126
R12270 out_p.n540 out_p.t1681 8.126
R12271 out_p.n541 out_p.t1600 8.126
R12272 out_p.n541 out_p.t1017 8.126
R12273 out_p.n542 out_p.t496 8.126
R12274 out_p.n542 out_p.t846 8.126
R12275 out_p.n543 out_p.t1312 8.126
R12276 out_p.n543 out_p.t1505 8.126
R12277 out_p.n544 out_p.t810 8.126
R12278 out_p.n544 out_p.t764 8.126
R12279 out_p.n545 out_p.t690 8.126
R12280 out_p.n545 out_p.t429 8.126
R12281 out_p.n546 out_p.t1352 8.126
R12282 out_p.n546 out_p.t1549 8.126
R12283 out_p.n547 out_p.t1553 8.126
R12284 out_p.n547 out_p.t258 8.126
R12285 out_p.n548 out_p.t1680 8.126
R12286 out_p.n548 out_p.t883 8.126
R12287 out_p.n549 out_p.t1082 8.126
R12288 out_p.n549 out_p.t347 8.126
R12289 out_p.n552 out_p.t1491 8.126
R12290 out_p.n552 out_p.t1697 8.126
R12291 out_p.n553 out_p.t1623 8.126
R12292 out_p.n553 out_p.t666 8.126
R12293 out_p.n554 out_p.t579 8.126
R12294 out_p.n554 out_p.t886 8.126
R12295 out_p.n555 out_p.t1325 8.126
R12296 out_p.n555 out_p.t1524 8.126
R12297 out_p.n556 out_p.t903 8.126
R12298 out_p.n556 out_p.t868 8.126
R12299 out_p.n557 out_p.t694 8.126
R12300 out_p.n557 out_p.t475 8.126
R12301 out_p.n558 out_p.t1372 8.126
R12302 out_p.n558 out_p.t1572 8.126
R12303 out_p.n559 out_p.t1576 8.126
R12304 out_p.n559 out_p.t980 8.126
R12305 out_p.n560 out_p.t1695 8.126
R12306 out_p.n560 out_p.t919 8.126
R12307 out_p.n561 out_p.t616 8.126
R12308 out_p.n561 out_p.t413 8.126
R12309 out_p.n564 out_p.t1096 8.126
R12310 out_p.n564 out_p.t1295 8.126
R12311 out_p.n565 out_p.t1215 8.126
R12312 out_p.n565 out_p.t1415 8.126
R12313 out_p.n566 out_p.t986 8.126
R12314 out_p.n566 out_p.t613 8.126
R12315 out_p.n567 out_p.t287 8.126
R12316 out_p.n567 out_p.t1124 8.126
R12317 out_p.n568 out_p.t1485 8.126
R12318 out_p.n568 out_p.t1686 8.126
R12319 out_p.n569 out_p.t879 8.126
R12320 out_p.n569 out_p.t878 8.126
R12321 out_p.n570 out_p.t391 8.126
R12322 out_p.n570 out_p.t1172 8.126
R12323 out_p.n571 out_p.t1173 8.126
R12324 out_p.n571 out_p.t1374 8.126
R12325 out_p.n572 out_p.t1293 8.126
R12326 out_p.n572 out_p.t1489 8.126
R12327 out_p.n573 out_p.t780 8.126
R12328 out_p.n573 out_p.t714 8.126
R12329 out_p.n576 out_p.t1161 8.126
R12330 out_p.n576 out_p.t865 8.126
R12331 out_p.n577 out_p.t1282 8.126
R12332 out_p.n577 out_p.t463 8.126
R12333 out_p.n578 out_p.t753 8.126
R12334 out_p.n578 out_p.t1574 8.126
R12335 out_p.n579 out_p.t420 8.126
R12336 out_p.n579 out_p.t1053 8.126
R12337 out_p.n580 out_p.t1544 8.126
R12338 out_p.n580 out_p.t1288 8.126
R12339 out_p.n581 out_p.t459 8.126
R12340 out_p.n581 out_p.t1687 8.126
R12341 out_p.n582 out_p.t508 8.126
R12342 out_p.n582 out_p.t635 8.126
R12343 out_p.n583 out_p.t1239 8.126
R12344 out_p.n583 out_p.t403 8.126
R12345 out_p.n584 out_p.t1363 8.126
R12346 out_p.n584 out_p.t1095 8.126
R12347 out_p.n585 out_p.t320 8.126
R12348 out_p.n585 out_p.t1661 8.126
R12349 out_p.n588 out_p.t1086 8.126
R12350 out_p.n588 out_p.t359 8.126
R12351 out_p.n589 out_p.t847 8.126
R12352 out_p.n589 out_p.t588 8.126
R12353 out_p.n590 out_p.t1435 8.126
R12354 out_p.n590 out_p.t1640 8.126
R12355 out_p.n591 out_p.t768 8.126
R12356 out_p.n591 out_p.t669 8.126
R12357 out_p.n592 out_p.t1145 8.126
R12358 out_p.n592 out_p.t1348 8.126
R12359 out_p.n593 out_p.t1548 8.126
R12360 out_p.n593 out_p.t1751 8.126
R12361 out_p.n594 out_p.t321 8.126
R12362 out_p.n594 out_p.t746 8.126
R12363 out_p.n595 out_p.t756 8.126
R12364 out_p.n595 out_p.t516 8.126
R12365 out_p.n596 out_p.t360 8.126
R12366 out_p.n596 out_p.t1159 8.126
R12367 out_p.n597 out_p.t1512 8.126
R12368 out_p.n597 out_p.t1718 8.126
R12369 out_p.n600 out_p.t723 8.126
R12370 out_p.n600 out_p.t625 8.126
R12371 out_p.n601 out_p.t494 8.126
R12372 out_p.n601 out_p.t537 8.126
R12373 out_p.n602 out_p.t506 8.126
R12374 out_p.n602 out_p.t1234 8.126
R12375 out_p.n603 out_p.t1667 8.126
R12376 out_p.n603 out_p.t843 8.126
R12377 out_p.n604 out_p.t1081 8.126
R12378 out_p.n604 out_p.t326 8.126
R12379 out_p.n605 out_p.t1148 8.126
R12380 out_p.n605 out_p.t1351 8.126
R12381 out_p.n606 out_p.t1713 8.126
R12382 out_p.n606 out_p.t312 8.126
R12383 out_p.n607 out_p.t299 8.126
R12384 out_p.n607 out_p.t304 8.126
R12385 out_p.n608 out_p.t626 8.126
R12386 out_p.n608 out_p.t1088 8.126
R12387 out_p.n609 out_p.t1119 8.126
R12388 out_p.n609 out_p.t1317 8.126
R12389 out_p.n612 out_p.t744 8.126
R12390 out_p.n612 out_p.t657 8.126
R12391 out_p.n613 out_p.t1039 8.126
R12392 out_p.n613 out_p.t932 8.126
R12393 out_p.n614 out_p.t1262 8.126
R12394 out_p.n614 out_p.t1464 8.126
R12395 out_p.n615 out_p.t899 8.126
R12396 out_p.n615 out_p.t914 8.126
R12397 out_p.n616 out_p.t402 8.126
R12398 out_p.n616 out_p.t1176 8.126
R12399 out_p.n617 out_p.t1379 8.126
R12400 out_p.n617 out_p.t1582 8.126
R12401 out_p.n618 out_p.t416 8.126
R12402 out_p.n618 out_p.t478 8.126
R12403 out_p.n619 out_p.t495 8.126
R12404 out_p.n619 out_p.t816 8.126
R12405 out_p.n620 out_p.t641 8.126
R12406 out_p.n620 out_p.t409 8.126
R12407 out_p.n621 out_p.t1346 8.126
R12408 out_p.n621 out_p.t1542 8.126
R12409 out_p.n624 out_p.t1665 8.126
R12410 out_p.n624 out_p.t833 8.126
R12411 out_p.n625 out_p.t1008 8.126
R12412 out_p.n625 out_p.t1024 8.126
R12413 out_p.n626 out_p.t805 8.126
R12414 out_p.n626 out_p.t557 8.126
R12415 out_p.n627 out_p.t1487 8.126
R12416 out_p.n627 out_p.t1690 8.126
R12417 out_p.n628 out_p.t718 8.126
R12418 out_p.n628 out_p.t617 8.126
R12419 out_p.n629 out_p.t389 8.126
R12420 out_p.n629 out_p.t1178 8.126
R12421 out_p.n630 out_p.t1537 8.126
R12422 out_p.n630 out_p.t1741 8.126
R12423 out_p.n631 out_p.t1743 8.126
R12424 out_p.n631 out_p.t415 8.126
R12425 out_p.n632 out_p.t799 8.126
R12426 out_p.n632 out_p.t748 8.126
R12427 out_p.n633 out_p.t956 8.126
R12428 out_p.n633 out_p.t1143 8.126
R12429 out_p.n636 out_p.t1729 8.126
R12430 out_p.n636 out_p.t1459 8.126
R12431 out_p.n637 out_p.t760 8.126
R12432 out_p.n637 out_p.t1586 8.126
R12433 out_p.n638 out_p.t309 8.126
R12434 out_p.n638 out_p.t445 8.126
R12435 out_p.n639 out_p.t1560 8.126
R12436 out_p.n639 out_p.t1289 8.126
R12437 out_p.n640 out_p.t376 8.126
R12438 out_p.n640 out_p.t813 8.126
R12439 out_p.n641 out_p.t522 8.126
R12440 out_p.n641 out_p.t633 8.126
R12441 out_p.n642 out_p.t1603 8.126
R12442 out_p.n642 out_p.t1341 8.126
R12443 out_p.n643 out_p.t962 8.126
R12444 out_p.n643 out_p.t1538 8.126
R12445 out_p.n644 out_p.t386 8.126
R12446 out_p.n644 out_p.t1664 8.126
R12447 out_p.n645 out_p.t455 8.126
R12448 out_p.n645 out_p.t1080 8.126
R12449 out_p.n648 out_p.t1322 8.126
R12450 out_p.n648 out_p.t1521 8.126
R12451 out_p.n649 out_p.t1450 8.126
R12452 out_p.n649 out_p.t1653 8.126
R12453 out_p.n650 out_p.t289 8.126
R12454 out_p.n650 out_p.t1057 8.126
R12455 out_p.n651 out_p.t1154 8.126
R12456 out_p.n651 out_p.t1357 8.126
R12457 out_p.n652 out_p.t1716 8.126
R12458 out_p.n652 out_p.t323 8.126
R12459 out_p.n653 out_p.t387 8.126
R12460 out_p.n653 out_p.t792 8.126
R12461 out_p.n654 out_p.t1201 8.126
R12462 out_p.n654 out_p.t1398 8.126
R12463 out_p.n655 out_p.t1402 8.126
R12464 out_p.n655 out_p.t1607 8.126
R12465 out_p.n656 out_p.t1520 8.126
R12466 out_p.n656 out_p.t1728 8.126
R12467 out_p.n657 out_p.t858 8.126
R12468 out_p.n657 out_p.t712 8.126
R12469 out_p.n660 out_p.t1556 8.126
R12470 out_p.n660 out_p.t1122 8.126
R12471 out_p.n661 out_p.t1682 8.126
R12472 out_p.n661 out_p.t1249 8.126
R12473 out_p.n662 out_p.t638 8.126
R12474 out_p.n662 out_p.t1004 8.126
R12475 out_p.n663 out_p.t1386 8.126
R12476 out_p.n663 out_p.t336 8.126
R12477 out_p.n664 out_p.t425 8.126
R12478 out_p.n664 out_p.t1511 8.126
R12479 out_p.n665 out_p.t825 8.126
R12480 out_p.n665 out_p.t322 8.126
R12481 out_p.n666 out_p.t1430 8.126
R12482 out_p.n666 out_p.t437 8.126
R12483 out_p.n667 out_p.t1637 8.126
R12484 out_p.n667 out_p.t1203 8.126
R12485 out_p.n668 out_p.t264 8.126
R12486 out_p.n668 out_p.t1321 8.126
R12487 out_p.n669 out_p.t782 8.126
R12488 out_p.n669 out_p.t869 8.126
R12489 out_p.n672 out_p.t1152 8.126
R12490 out_p.n672 out_p.t1354 8.126
R12491 out_p.n673 out_p.t1275 8.126
R12492 out_p.n673 out_p.t1478 8.126
R12493 out_p.n674 out_p.t698 8.126
R12494 out_p.n674 out_p.t620 8.126
R12495 out_p.n675 out_p.t399 8.126
R12496 out_p.n675 out_p.t1185 8.126
R12497 out_p.n676 out_p.t1539 8.126
R12498 out_p.n676 out_p.t1745 8.126
R12499 out_p.n677 out_p.t434 8.126
R12500 out_p.n677 out_p.t512 8.126
R12501 out_p.n678 out_p.t509 8.126
R12502 out_p.n678 out_p.t1230 8.126
R12503 out_p.n679 out_p.t1232 8.126
R12504 out_p.n679 out_p.t1433 8.126
R12505 out_p.n680 out_p.t1353 8.126
R12506 out_p.n680 out_p.t1555 8.126
R12507 out_p.n681 out_p.t311 8.126
R12508 out_p.n681 out_p.t342 8.126
R12509 out_p.n684 out_p.t1092 8.126
R12510 out_p.n684 out_p.t350 8.126
R12511 out_p.n685 out_p.t851 8.126
R12512 out_p.n685 out_p.t580 8.126
R12513 out_p.n686 out_p.t1432 8.126
R12514 out_p.n686 out_p.t1636 8.126
R12515 out_p.n687 out_p.t738 8.126
R12516 out_p.n687 out_p.t628 8.126
R12517 out_p.n688 out_p.t1142 8.126
R12518 out_p.n688 out_p.t1345 8.126
R12519 out_p.n689 out_p.t1541 8.126
R12520 out_p.n689 out_p.t1747 8.126
R12521 out_p.n690 out_p.t284 8.126
R12522 out_p.n690 out_p.t747 8.126
R12523 out_p.n691 out_p.t745 8.126
R12524 out_p.n691 out_p.t507 8.126
R12525 out_p.n692 out_p.t337 8.126
R12526 out_p.n692 out_p.t1151 8.126
R12527 out_p.n693 out_p.t1510 8.126
R12528 out_p.n693 out_p.t1715 8.126
R12529 out_p.n696 out_p.t732 8.126
R12530 out_p.n696 out_p.t1184 8.126
R12531 out_p.n697 out_p.t316 8.126
R12532 out_p.n697 out_p.t1311 8.126
R12533 out_p.n698 out_p.t1493 8.126
R12534 out_p.n698 out_p.t809 8.126
R12535 out_p.n699 out_p.t367 8.126
R12536 out_p.n699 out_p.t484 8.126
R12537 out_p.n700 out_p.t1206 8.126
R12538 out_p.n700 out_p.t1575 8.126
R12539 out_p.n701 out_p.t1616 8.126
R12540 out_p.n701 out_p.t984 8.126
R12541 out_p.n702 out_p.t555 8.126
R12542 out_p.n702 out_p.t558 8.126
R12543 out_p.n703 out_p.t891 8.126
R12544 out_p.n703 out_p.t1261 8.126
R12545 out_p.n704 out_p.t471 8.126
R12546 out_p.n704 out_p.t1385 8.126
R12547 out_p.n705 out_p.t1578 8.126
R12548 out_p.n705 out_p.t414 8.126
R12549 out_p.n708 out_p.t923 8.126
R12550 out_p.n708 out_p.t894 8.126
R12551 out_p.n709 out_p.t981 8.126
R12552 out_p.n709 out_p.t1072 8.126
R12553 out_p.n710 out_p.t1098 8.126
R12554 out_p.n710 out_p.t1298 8.126
R12555 out_p.n711 out_p.t1723 8.126
R12556 out_p.n711 out_p.t341 8.126
R12557 out_p.n712 out_p.t700 8.126
R12558 out_p.n712 out_p.t447 8.126
R12559 out_p.n713 out_p.t1208 8.126
R12560 out_p.n713 out_p.t1408 8.126
R12561 out_p.n714 out_p.t268 8.126
R12562 out_p.n714 out_p.t561 8.126
R12563 out_p.n715 out_p.t576 8.126
R12564 out_p.n715 out_p.t564 8.126
R12565 out_p.n716 out_p.t898 8.126
R12566 out_p.n716 out_p.t705 8.126
R12567 out_p.n717 out_p.t1174 8.126
R12568 out_p.n717 out_p.t1375 8.126
R12569 out_p.n720 out_p.t384 8.126
R12570 out_p.n720 out_p.t1689 8.126
R12571 out_p.n721 out_p.t623 8.126
R12572 out_p.n721 out_p.t645 8.126
R12573 out_p.n722 out_p.t1324 8.126
R12574 out_p.n722 out_p.t876 8.126
R12575 out_p.n723 out_p.t493 8.126
R12576 out_p.n723 out_p.t1516 8.126
R12577 out_p.n724 out_p.t517 8.126
R12578 out_p.n724 out_p.t844 8.126
R12579 out_p.n725 out_p.t1444 8.126
R12580 out_p.n725 out_p.t467 8.126
R12581 out_p.n726 out_p.t961 8.126
R12582 out_p.n726 out_p.t1571 8.126
R12583 out_p.n727 out_p.t1056 8.126
R12584 out_p.n727 out_p.t964 8.126
R12585 out_p.n728 out_p.t786 8.126
R12586 out_p.n728 out_p.t889 8.126
R12587 out_p.n729 out_p.t1404 8.126
R12588 out_p.n729 out_p.t390 8.126
R12589 out_p.n732 out_p.t1722 8.126
R12590 out_p.n732 out_p.t354 8.126
R12591 out_p.n733 out_p.t749 8.126
R12592 out_p.n733 out_p.t662 8.126
R12593 out_p.n734 out_p.t276 8.126
R12594 out_p.n734 out_p.t1123 8.126
R12595 out_p.n735 out_p.t1552 8.126
R12596 out_p.n735 out_p.t1755 8.126
R12597 out_p.n736 out_p.t355 8.126
R12598 out_p.n736 out_p.t757 8.126
R12599 out_p.n737 out_p.t515 8.126
R12600 out_p.n737 out_p.t1241 8.126
R12601 out_p.n738 out_p.t1601 8.126
R12602 out_p.n738 out_p.t985 8.126
R12603 out_p.n739 out_p.t1016 8.126
R12604 out_p.n739 out_p.t282 8.126
R12605 out_p.n740 out_p.t343 8.126
R12606 out_p.n740 out_p.t407 8.126
R12607 out_p.n741 out_p.t458 8.126
R12608 out_p.n741 out_p.t1204 8.126
R12609 out_p.n0 out_p.t949 8.126
R12610 out_p.n0 out_p.t357 8.126
R12611 out_p.n1 out_p.t872 8.126
R12612 out_p.n1 out_p.t598 8.126
R12613 out_p.n2 out_p.t1439 8.126
R12614 out_p.n2 out_p.t1644 8.126
R12615 out_p.n3 out_p.t794 8.126
R12616 out_p.n3 out_p.t663 8.126
R12617 out_p.n4 out_p.t1147 8.126
R12618 out_p.n4 out_p.t1350 8.126
R12619 out_p.n5 out_p.t1551 8.126
R12620 out_p.n5 out_p.t1754 8.126
R12621 out_p.n6 out_p.t293 8.126
R12622 out_p.n6 out_p.t772 8.126
R12623 out_p.n7 out_p.t767 8.126
R12624 out_p.n7 out_p.t524 8.126
R12625 out_p.n8 out_p.t371 8.126
R12626 out_p.n8 out_p.t1165 8.126
R12627 out_p.n9 out_p.t1514 8.126
R12628 out_p.n9 out_p.t1720 8.126
R12629 out_p.n731 out_p.t185 4.95
R12630 out_p.n731 out_p.t145 4.95
R12631 out_p.n730 out_p.t162 4.95
R12632 out_p.n730 out_p.t49 4.95
R12633 out_p.n718 out_p.t106 4.95
R12634 out_p.n718 out_p.t167 4.95
R12635 out_p.n719 out_p.t93 4.95
R12636 out_p.n719 out_p.t192 4.95
R12637 out_p.n706 out_p.t54 4.95
R12638 out_p.n706 out_p.t114 4.95
R12639 out_p.n707 out_p.t151 4.95
R12640 out_p.n707 out_p.t100 4.95
R12641 out_p.n694 out_p.t239 4.95
R12642 out_p.n694 out_p.t1765 4.95
R12643 out_p.n695 out_p.t29 4.95
R12644 out_p.n695 out_p.t230 4.95
R12645 out_p.n682 out_p.t252 4.95
R12646 out_p.n682 out_p.t210 4.95
R12647 out_p.n683 out_p.t110 4.95
R12648 out_p.n683 out_p.t82 4.95
R12649 out_p.n670 out_p.t1772 4.95
R12650 out_p.n670 out_p.t17 4.95
R12651 out_p.n671 out_p.t197 4.95
R12652 out_p.n671 out_p.t1798 4.95
R12653 out_p.n658 out_p.t195 4.95
R12654 out_p.n658 out_p.t1775 4.95
R12655 out_p.n659 out_p.t3 4.95
R12656 out_p.n659 out_p.t202 4.95
R12657 out_p.n646 out_p.t1782 4.95
R12658 out_p.n646 out_p.t128 4.95
R12659 out_p.n647 out_p.t1762 4.95
R12660 out_p.n647 out_p.t9 4.95
R12661 out_p.n634 out_p.t160 4.95
R12662 out_p.n634 out_p.t137 4.95
R12663 out_p.n635 out_p.t183 4.95
R12664 out_p.n635 out_p.t1780 4.95
R12665 out_p.n622 out_p.t171 4.95
R12666 out_p.n622 out_p.t60 4.95
R12667 out_p.n623 out_p.t125 4.95
R12668 out_p.n623 out_p.t157 4.95
R12669 out_p.n610 out_p.t119 4.95
R12670 out_p.n610 out_p.t245 4.95
R12671 out_p.n611 out_p.t45 4.95
R12672 out_p.n611 out_p.t36 4.95
R12673 out_p.n598 out_p.t40 4.95
R12674 out_p.n598 out_p.t124 4.95
R12675 out_p.n599 out_p.t164 4.95
R12676 out_p.n599 out_p.t51 4.95
R12677 out_p.n586 out_p.t251 4.95
R12678 out_p.n586 out_p.t209 4.95
R12679 out_p.n587 out_p.t109 4.95
R12680 out_p.n587 out_p.t81 4.95
R12681 out_p.n574 out_p.t1770 4.95
R12682 out_p.n574 out_p.t67 4.95
R12683 out_p.n575 out_p.t235 4.95
R12684 out_p.n575 out_p.t248 4.95
R12685 out_p.n562 out_p.t219 4.95
R12686 out_p.n562 out_p.t1787 4.95
R12687 out_p.n563 out_p.t206 4.95
R12688 out_p.n563 out_p.t1767 4.95
R12689 out_p.n550 out_p.t133 4.95
R12690 out_p.n550 out_p.t166 4.95
R12691 out_p.n551 out_p.t14 4.95
R12692 out_p.n551 out_p.t191 4.95
R12693 out_p.n538 out_p.t136 4.95
R12694 out_p.n538 out_p.t170 4.95
R12695 out_p.n539 out_p.t18 4.95
R12696 out_p.n539 out_p.t196 4.95
R12697 out_p.n526 out_p.t57 4.95
R12698 out_p.n526 out_p.t117 4.95
R12699 out_p.n527 out_p.t154 4.95
R12700 out_p.n527 out_p.t104 4.95
R12701 out_p.n514 out_p.t242 4.95
R12702 out_p.n514 out_p.t89 4.95
R12703 out_p.n515 out_p.t33 4.95
R12704 out_p.n515 out_p.t56 4.95
R12705 out_p.n502 out_p.t19 4.95
R12706 out_p.n502 out_p.t215 4.95
R12707 out_p.n503 out_p.t116 4.95
R12708 out_p.n503 out_p.t241 4.95
R12709 out_p.n490 out_p.t1774 4.95
R12710 out_p.n490 out_p.t25 4.95
R12711 out_p.n491 out_p.t201 4.95
R12712 out_p.n491 out_p.t122 4.95
R12713 out_p.n478 out_p.t66 4.95
R12714 out_p.n478 out_p.t218 4.95
R12715 out_p.n479 out_p.t247 4.95
R12716 out_p.n479 out_p.t205 4.95
R12717 out_p.n466 out_p.t1786 4.95
R12718 out_p.n466 out_p.t131 4.95
R12719 out_p.n467 out_p.t1766 4.95
R12720 out_p.n467 out_p.t12 4.95
R12721 out_p.n454 out_p.t226 4.95
R12722 out_p.n454 out_p.t0 4.95
R12723 out_p.n455 out_p.t212 4.95
R12724 out_p.n455 out_p.t1785 4.95
R12725 out_p.n442 out_p.t176 4.95
R12726 out_p.n442 out_p.t39 4.95
R12727 out_p.n443 out_p.t130 4.95
R12728 out_p.n443 out_p.t163 4.95
R12729 out_p.n430 out_p.t123 4.95
R12730 out_p.n430 out_p.t180 4.95
R12731 out_p.n431 out_p.t50 4.95
R12732 out_p.n431 out_p.t135 4.95
R12733 out_p.n418 out_p.t1778 4.95
R12734 out_p.n418 out_p.t88 4.95
R12735 out_p.n419 out_p.t169 4.95
R12736 out_p.n419 out_p.t55 4.95
R12737 out_p.n406 out_p.t256 4.95
R12738 out_p.n406 out_p.t214 4.95
R12739 out_p.n407 out_p.t115 4.95
R12740 out_p.n407 out_p.t240 4.95
R12741 out_p.n394 out_p.t94 4.95
R12742 out_p.n394 out_p.t73 4.95
R12743 out_p.n395 out_p.t61 4.95
R12744 out_p.n395 out_p.t255 4.95
R12745 out_p.n382 out_p.t227 4.95
R12746 out_p.n382 out_p.t1791 4.95
R12747 out_p.n383 out_p.t213 4.95
R12748 out_p.n383 out_p.t1773 4.95
R12749 out_p.n370 out_p.t78 4.95
R12750 out_p.n370 out_p.t232 4.95
R12751 out_p.n371 out_p.t22 4.95
R12752 out_p.n371 out_p.t64 4.95
R12753 out_p.n358 out_p.t1794 4.95
R12754 out_p.n358 out_p.t142 4.95
R12755 out_p.n359 out_p.t1776 4.95
R12756 out_p.n359 out_p.t1783 4.95
R12757 out_p.n346 out_p.t175 4.95
R12758 out_p.n346 out_p.t1758 4.95
R12759 out_p.n347 out_p.t129 4.95
R12760 out_p.n347 out_p.t222 4.95
R12761 out_p.n334 out_p.t4 4.95
R12762 out_p.n334 out_p.t147 4.95
R12763 out_p.n335 out_p.t1788 4.95
R12764 out_p.n335 out_p.t173 4.95
R12765 out_p.n322 out_p.t95 4.95
R12766 out_p.n322 out_p.t23 4.95
R12767 out_p.n323 out_p.t62 4.95
R12768 out_p.n323 out_p.t120 4.95
R12769 out_p.n310 out_p.t153 4.95
R12770 out_p.n310 out_p.t102 4.95
R12771 out_p.n311 out_p.t178 4.95
R12772 out_p.n311 out_p.t42 4.95
R12773 out_p.n298 out_p.t30 4.95
R12774 out_p.n298 out_p.t71 4.95
R12775 out_p.n299 out_p.t85 4.95
R12776 out_p.n299 out_p.t253 4.95
R12777 out_p.n286 out_p.t225 4.95
R12778 out_p.n286 out_p.t38 4.95
R12779 out_p.n287 out_p.t211 4.95
R12780 out_p.n287 out_p.t91 4.95
R12781 out_p.n274 out_p.t76 4.95
R12782 out_p.n274 out_p.t1759 4.95
R12783 out_p.n275 out_p.t20 4.95
R12784 out_p.n275 out_p.t223 4.95
R12785 out_p.n262 out_p.t5 4.95
R12786 out_p.n262 out_p.t189 4.95
R12787 out_p.n263 out_p.t1789 4.95
R12788 out_p.n263 out_p.t141 4.95
R12789 out_p.n250 out_p.t148 4.95
R12790 out_p.n250 out_p.t96 4.95
R12791 out_p.n251 out_p.t174 4.95
R12792 out_p.n251 out_p.t63 4.95
R12793 out_p.n238 out_p.t24 4.95
R12794 out_p.n238 out_p.t65 4.95
R12795 out_p.n239 out_p.t121 4.95
R12796 out_p.n239 out_p.t246 4.95
R12797 out_p.n226 out_p.t103 4.95
R12798 out_p.n226 out_p.t31 4.95
R12799 out_p.n227 out_p.t43 4.95
R12800 out_p.n227 out_p.t86 4.95
R12801 out_p.n214 out_p.t72 4.95
R12802 out_p.n214 out_p.t1795 4.95
R12803 out_p.n215 out_p.t254 4.95
R12804 out_p.n215 out_p.t217 4.95
R12805 out_p.n202 out_p.t143 4.95
R12806 out_p.n202 out_p.t200 4.95
R12807 out_p.n203 out_p.t1784 4.95
R12808 out_p.n203 out_p.t70 4.95
R12809 out_p.n190 out_p.t1760 4.95
R12810 out_p.n190 out_p.t6 4.95
R12811 out_p.n191 out_p.t224 4.95
R12812 out_p.n191 out_p.t1790 4.95
R12813 out_p.n178 out_p.t179 4.95
R12814 out_p.n178 out_p.t1777 4.95
R12815 out_p.n179 out_p.t134 4.95
R12816 out_p.n179 out_p.t168 4.95
R12817 out_p.n166 out_p.t11 4.95
R12818 out_p.n166 out_p.t187 4.95
R12819 out_p.n167 out_p.t1793 4.95
R12820 out_p.n167 out_p.t139 4.95
R12821 out_p.n154 out_p.t146 4.95
R12822 out_p.n154 out_p.t32 4.95
R12823 out_p.n155 out_p.t172 4.95
R12824 out_p.n155 out_p.t87 4.95
R12825 out_p.n142 out_p.t161 4.95
R12826 out_p.n142 out_p.t48 4.95
R12827 out_p.n143 out_p.t184 4.95
R12828 out_p.n143 out_p.t144 4.95
R12829 out_p.n130 out_p.t105 4.95
R12830 out_p.n130 out_p.t77 4.95
R12831 out_p.n131 out_p.t92 4.95
R12832 out_p.n131 out_p.t21 4.95
R12833 out_p.n118 out_p.t231 4.95
R12834 out_p.n118 out_p.t112 4.95
R12835 out_p.n119 out_p.t216 4.95
R12836 out_p.n119 out_p.t98 4.95
R12837 out_p.n106 out_p.t237 4.95
R12838 out_p.n106 out_p.t198 4.95
R12839 out_p.n107 out_p.t27 4.95
R12840 out_p.n107 out_p.t68 4.95
R12841 out_p.n94 out_p.t1799 4.95
R12842 out_p.n94 out_p.t188 4.95
R12843 out_p.n95 out_p.t220 4.95
R12844 out_p.n95 out_p.t140 4.95
R12845 out_p.n82 out_p.t1771 4.95
R12846 out_p.n82 out_p.t16 4.95
R12847 out_p.n83 out_p.t236 4.95
R12848 out_p.n83 out_p.t1797 4.95
R12849 out_p.n70 out_p.t194 4.95
R12850 out_p.n70 out_p.t152 4.95
R12851 out_p.n71 out_p.t2 4.95
R12852 out_p.n71 out_p.t177 4.95
R12853 out_p.n58 out_p.t101 4.95
R12854 out_p.n58 out_p.t126 4.95
R12855 out_p.n59 out_p.t41 4.95
R12856 out_p.n59 out_p.t7 4.95
R12857 out_p.n46 out_p.t158 4.95
R12858 out_p.n46 out_p.t46 4.95
R12859 out_p.n47 out_p.t181 4.95
R12860 out_p.n47 out_p.t1779 4.95
R12861 out_p.n34 out_p.t37 4.95
R12862 out_p.n34 out_p.t59 4.95
R12863 out_p.n35 out_p.t90 4.95
R12864 out_p.n35 out_p.t156 4.95
R12865 out_p.n22 out_p.t118 4.95
R12866 out_p.n22 out_p.t243 4.95
R12867 out_p.n23 out_p.t44 4.95
R12868 out_p.n23 out_p.t34 4.95
R12869 out_p.n20 out_p.t203 4.95
R12870 out_p.n20 out_p.t1763 4.95
R12871 out_p.n21 out_p.t74 4.95
R12872 out_p.n21 out_p.t228 4.95
R12873 out_p.n802 out_p.t1768 4.95
R12874 out_p.n802 out_p.t15 4.95
R12875 out_p.n803 out_p.t233 4.95
R12876 out_p.n803 out_p.t1796 4.95
R12877 out_p.n804 out_p.t193 4.95
R12878 out_p.n804 out_p.t53 4.95
R12879 out_p.n805 out_p.t1 4.95
R12880 out_p.n805 out_p.t150 4.95
R12881 out_p.n806 out_p.t113 4.95
R12882 out_p.n806 out_p.t238 4.95
R12883 out_p.n807 out_p.t99 4.95
R12884 out_p.n807 out_p.t28 4.95
R12885 out_p.n808 out_p.t199 4.95
R12886 out_p.n808 out_p.t1757 4.95
R12887 out_p.n809 out_p.t69 4.95
R12888 out_p.n809 out_p.t221 4.95
R12889 out_p.n810 out_p.t244 4.95
R12890 out_p.n810 out_p.t204 4.95
R12891 out_p.n811 out_p.t35 4.95
R12892 out_p.n811 out_p.t75 4.95
R12893 out_p.n812 out_p.t1764 4.95
R12894 out_p.n812 out_p.t10 4.95
R12895 out_p.n813 out_p.t229 4.95
R12896 out_p.n813 out_p.t1792 4.95
R12897 out_p.n814 out_p.t186 4.95
R12898 out_p.n814 out_p.t1781 4.95
R12899 out_p.n815 out_p.t138 4.95
R12900 out_p.n815 out_p.t1761 4.95
R12901 out_p.n816 out_p.t127 4.95
R12902 out_p.n816 out_p.t159 4.95
R12903 out_p.n817 out_p.t8 4.95
R12904 out_p.n817 out_p.t182 4.95
R12905 out_p.n818 out_p.t47 4.95
R12906 out_p.n818 out_p.t132 4.95
R12907 out_p.n819 out_p.t84 4.95
R12908 out_p.n819 out_p.t13 4.95
R12909 out_p.n820 out_p.t165 4.95
R12910 out_p.n820 out_p.t52 4.95
R12911 out_p.n821 out_p.t190 4.95
R12912 out_p.n821 out_p.t149 4.95
R12913 out_p.n822 out_p.t111 4.95
R12914 out_p.n822 out_p.t83 4.95
R12915 out_p.n823 out_p.t97 4.95
R12916 out_p.n823 out_p.t26 4.95
R12917 out_p.n824 out_p.t58 4.95
R12918 out_p.n824 out_p.t250 4.95
R12919 out_p.n825 out_p.t155 4.95
R12920 out_p.n825 out_p.t108 4.95
R12921 out_p.n826 out_p.t208 4.95
R12922 out_p.n826 out_p.t1769 4.95
R12923 out_p.n827 out_p.t80 4.95
R12924 out_p.n827 out_p.t234 4.95
R12925 out_p.n971 out_p.t249 4.95
R12926 out_p.n971 out_p.t207 4.95
R12927 out_p.n972 out_p.t107 4.95
R12928 out_p.n972 out_p.t79 4.95
R12929 out_p.n737 out_p.n736 0.866
R12930 out_p.n833 out_p.n832 0.85
R12931 out_p.n844 out_p.n843 0.85
R12932 out_p.n855 out_p.n854 0.85
R12933 out_p.n866 out_p.n865 0.85
R12934 out_p.n877 out_p.n876 0.85
R12935 out_p.n888 out_p.n887 0.85
R12936 out_p.n899 out_p.n898 0.85
R12937 out_p.n910 out_p.n909 0.85
R12938 out_p.n921 out_p.n920 0.85
R12939 out_p.n932 out_p.n931 0.85
R12940 out_p.n943 out_p.n942 0.85
R12941 out_p.n954 out_p.n953 0.85
R12942 out_p.n965 out_p.n964 0.85
R12943 out_p.n15 out_p.n14 0.85
R12944 out_p.n29 out_p.n28 0.85
R12945 out_p.n41 out_p.n40 0.85
R12946 out_p.n53 out_p.n52 0.85
R12947 out_p.n65 out_p.n64 0.85
R12948 out_p.n77 out_p.n76 0.85
R12949 out_p.n89 out_p.n88 0.85
R12950 out_p.n101 out_p.n100 0.85
R12951 out_p.n113 out_p.n112 0.85
R12952 out_p.n125 out_p.n124 0.85
R12953 out_p.n137 out_p.n136 0.85
R12954 out_p.n149 out_p.n148 0.85
R12955 out_p.n161 out_p.n160 0.85
R12956 out_p.n173 out_p.n172 0.85
R12957 out_p.n185 out_p.n184 0.85
R12958 out_p.n197 out_p.n196 0.85
R12959 out_p.n209 out_p.n208 0.85
R12960 out_p.n221 out_p.n220 0.85
R12961 out_p.n233 out_p.n232 0.85
R12962 out_p.n245 out_p.n244 0.85
R12963 out_p.n257 out_p.n256 0.85
R12964 out_p.n269 out_p.n268 0.85
R12965 out_p.n281 out_p.n280 0.85
R12966 out_p.n293 out_p.n292 0.85
R12967 out_p.n305 out_p.n304 0.85
R12968 out_p.n317 out_p.n316 0.85
R12969 out_p.n329 out_p.n328 0.85
R12970 out_p.n341 out_p.n340 0.85
R12971 out_p.n353 out_p.n352 0.85
R12972 out_p.n365 out_p.n364 0.85
R12973 out_p.n377 out_p.n376 0.85
R12974 out_p.n389 out_p.n388 0.85
R12975 out_p.n401 out_p.n400 0.85
R12976 out_p.n413 out_p.n412 0.85
R12977 out_p.n425 out_p.n424 0.85
R12978 out_p.n437 out_p.n436 0.85
R12979 out_p.n449 out_p.n448 0.85
R12980 out_p.n461 out_p.n460 0.85
R12981 out_p.n473 out_p.n472 0.85
R12982 out_p.n485 out_p.n484 0.85
R12983 out_p.n497 out_p.n496 0.85
R12984 out_p.n509 out_p.n508 0.85
R12985 out_p.n521 out_p.n520 0.85
R12986 out_p.n533 out_p.n532 0.85
R12987 out_p.n545 out_p.n544 0.85
R12988 out_p.n557 out_p.n556 0.85
R12989 out_p.n569 out_p.n568 0.85
R12990 out_p.n581 out_p.n580 0.85
R12991 out_p.n593 out_p.n592 0.85
R12992 out_p.n605 out_p.n604 0.85
R12993 out_p.n617 out_p.n616 0.85
R12994 out_p.n629 out_p.n628 0.85
R12995 out_p.n641 out_p.n640 0.85
R12996 out_p.n653 out_p.n652 0.85
R12997 out_p.n665 out_p.n664 0.85
R12998 out_p.n677 out_p.n676 0.85
R12999 out_p.n689 out_p.n688 0.85
R13000 out_p.n701 out_p.n700 0.85
R13001 out_p.n713 out_p.n712 0.85
R13002 out_p.n725 out_p.n724 0.85
R13003 out_p.n5 out_p.n4 0.85
R13004 out_p.n741 out_p.n740 0.77
R13005 out_p.n740 out_p.n739 0.77
R13006 out_p.n739 out_p.n738 0.77
R13007 out_p.n738 out_p.n737 0.77
R13008 out_p.n736 out_p.n735 0.77
R13009 out_p.n735 out_p.n734 0.77
R13010 out_p.n734 out_p.n733 0.77
R13011 out_p.n733 out_p.n732 0.77
R13012 out_p.n731 out_p.n730 0.76
R13013 out_p.n719 out_p.n718 0.76
R13014 out_p.n707 out_p.n706 0.76
R13015 out_p.n695 out_p.n694 0.76
R13016 out_p.n683 out_p.n682 0.76
R13017 out_p.n671 out_p.n670 0.76
R13018 out_p.n659 out_p.n658 0.76
R13019 out_p.n647 out_p.n646 0.76
R13020 out_p.n635 out_p.n634 0.76
R13021 out_p.n623 out_p.n622 0.76
R13022 out_p.n611 out_p.n610 0.76
R13023 out_p.n599 out_p.n598 0.76
R13024 out_p.n587 out_p.n586 0.76
R13025 out_p.n575 out_p.n574 0.76
R13026 out_p.n563 out_p.n562 0.76
R13027 out_p.n551 out_p.n550 0.76
R13028 out_p.n539 out_p.n538 0.76
R13029 out_p.n527 out_p.n526 0.76
R13030 out_p.n515 out_p.n514 0.76
R13031 out_p.n503 out_p.n502 0.76
R13032 out_p.n491 out_p.n490 0.76
R13033 out_p.n479 out_p.n478 0.76
R13034 out_p.n467 out_p.n466 0.76
R13035 out_p.n455 out_p.n454 0.76
R13036 out_p.n443 out_p.n442 0.76
R13037 out_p.n431 out_p.n430 0.76
R13038 out_p.n419 out_p.n418 0.76
R13039 out_p.n407 out_p.n406 0.76
R13040 out_p.n395 out_p.n394 0.76
R13041 out_p.n383 out_p.n382 0.76
R13042 out_p.n371 out_p.n370 0.76
R13043 out_p.n359 out_p.n358 0.76
R13044 out_p.n347 out_p.n346 0.76
R13045 out_p.n335 out_p.n334 0.76
R13046 out_p.n323 out_p.n322 0.76
R13047 out_p.n311 out_p.n310 0.76
R13048 out_p.n299 out_p.n298 0.76
R13049 out_p.n287 out_p.n286 0.76
R13050 out_p.n275 out_p.n274 0.76
R13051 out_p.n263 out_p.n262 0.76
R13052 out_p.n251 out_p.n250 0.76
R13053 out_p.n239 out_p.n238 0.76
R13054 out_p.n227 out_p.n226 0.76
R13055 out_p.n215 out_p.n214 0.76
R13056 out_p.n203 out_p.n202 0.76
R13057 out_p.n191 out_p.n190 0.76
R13058 out_p.n179 out_p.n178 0.76
R13059 out_p.n167 out_p.n166 0.76
R13060 out_p.n155 out_p.n154 0.76
R13061 out_p.n143 out_p.n142 0.76
R13062 out_p.n131 out_p.n130 0.76
R13063 out_p.n119 out_p.n118 0.76
R13064 out_p.n107 out_p.n106 0.76
R13065 out_p.n95 out_p.n94 0.76
R13066 out_p.n83 out_p.n82 0.76
R13067 out_p.n71 out_p.n70 0.76
R13068 out_p.n59 out_p.n58 0.76
R13069 out_p.n47 out_p.n46 0.76
R13070 out_p.n35 out_p.n34 0.76
R13071 out_p.n23 out_p.n22 0.76
R13072 out_p.n21 out_p.n20 0.76
R13073 out_p.n803 out_p.n802 0.76
R13074 out_p.n805 out_p.n804 0.76
R13075 out_p.n807 out_p.n806 0.76
R13076 out_p.n809 out_p.n808 0.76
R13077 out_p.n811 out_p.n810 0.76
R13078 out_p.n813 out_p.n812 0.76
R13079 out_p.n815 out_p.n814 0.76
R13080 out_p.n817 out_p.n816 0.76
R13081 out_p.n819 out_p.n818 0.76
R13082 out_p.n821 out_p.n820 0.76
R13083 out_p.n823 out_p.n822 0.76
R13084 out_p.n825 out_p.n824 0.76
R13085 out_p.n827 out_p.n826 0.76
R13086 out_p.n972 out_p.n971 0.76
R13087 out_p.n837 out_p.n836 0.754
R13088 out_p.n836 out_p.n835 0.754
R13089 out_p.n835 out_p.n834 0.754
R13090 out_p.n834 out_p.n833 0.754
R13091 out_p.n832 out_p.n831 0.754
R13092 out_p.n831 out_p.n830 0.754
R13093 out_p.n830 out_p.n829 0.754
R13094 out_p.n829 out_p.n828 0.754
R13095 out_p.n848 out_p.n847 0.754
R13096 out_p.n847 out_p.n846 0.754
R13097 out_p.n846 out_p.n845 0.754
R13098 out_p.n845 out_p.n844 0.754
R13099 out_p.n843 out_p.n842 0.754
R13100 out_p.n842 out_p.n841 0.754
R13101 out_p.n841 out_p.n840 0.754
R13102 out_p.n840 out_p.n839 0.754
R13103 out_p.n859 out_p.n858 0.754
R13104 out_p.n858 out_p.n857 0.754
R13105 out_p.n857 out_p.n856 0.754
R13106 out_p.n856 out_p.n855 0.754
R13107 out_p.n854 out_p.n853 0.754
R13108 out_p.n853 out_p.n852 0.754
R13109 out_p.n852 out_p.n851 0.754
R13110 out_p.n851 out_p.n850 0.754
R13111 out_p.n870 out_p.n869 0.754
R13112 out_p.n869 out_p.n868 0.754
R13113 out_p.n868 out_p.n867 0.754
R13114 out_p.n867 out_p.n866 0.754
R13115 out_p.n865 out_p.n864 0.754
R13116 out_p.n864 out_p.n863 0.754
R13117 out_p.n863 out_p.n862 0.754
R13118 out_p.n862 out_p.n861 0.754
R13119 out_p.n881 out_p.n880 0.754
R13120 out_p.n880 out_p.n879 0.754
R13121 out_p.n879 out_p.n878 0.754
R13122 out_p.n878 out_p.n877 0.754
R13123 out_p.n876 out_p.n875 0.754
R13124 out_p.n875 out_p.n874 0.754
R13125 out_p.n874 out_p.n873 0.754
R13126 out_p.n873 out_p.n872 0.754
R13127 out_p.n892 out_p.n891 0.754
R13128 out_p.n891 out_p.n890 0.754
R13129 out_p.n890 out_p.n889 0.754
R13130 out_p.n889 out_p.n888 0.754
R13131 out_p.n887 out_p.n886 0.754
R13132 out_p.n886 out_p.n885 0.754
R13133 out_p.n885 out_p.n884 0.754
R13134 out_p.n884 out_p.n883 0.754
R13135 out_p.n903 out_p.n902 0.754
R13136 out_p.n902 out_p.n901 0.754
R13137 out_p.n901 out_p.n900 0.754
R13138 out_p.n900 out_p.n899 0.754
R13139 out_p.n898 out_p.n897 0.754
R13140 out_p.n897 out_p.n896 0.754
R13141 out_p.n896 out_p.n895 0.754
R13142 out_p.n895 out_p.n894 0.754
R13143 out_p.n914 out_p.n913 0.754
R13144 out_p.n913 out_p.n912 0.754
R13145 out_p.n912 out_p.n911 0.754
R13146 out_p.n911 out_p.n910 0.754
R13147 out_p.n909 out_p.n908 0.754
R13148 out_p.n908 out_p.n907 0.754
R13149 out_p.n907 out_p.n906 0.754
R13150 out_p.n906 out_p.n905 0.754
R13151 out_p.n925 out_p.n924 0.754
R13152 out_p.n924 out_p.n923 0.754
R13153 out_p.n923 out_p.n922 0.754
R13154 out_p.n922 out_p.n921 0.754
R13155 out_p.n920 out_p.n919 0.754
R13156 out_p.n919 out_p.n918 0.754
R13157 out_p.n918 out_p.n917 0.754
R13158 out_p.n917 out_p.n916 0.754
R13159 out_p.n936 out_p.n935 0.754
R13160 out_p.n935 out_p.n934 0.754
R13161 out_p.n934 out_p.n933 0.754
R13162 out_p.n933 out_p.n932 0.754
R13163 out_p.n931 out_p.n930 0.754
R13164 out_p.n930 out_p.n929 0.754
R13165 out_p.n929 out_p.n928 0.754
R13166 out_p.n928 out_p.n927 0.754
R13167 out_p.n947 out_p.n946 0.754
R13168 out_p.n946 out_p.n945 0.754
R13169 out_p.n945 out_p.n944 0.754
R13170 out_p.n944 out_p.n943 0.754
R13171 out_p.n942 out_p.n941 0.754
R13172 out_p.n941 out_p.n940 0.754
R13173 out_p.n940 out_p.n939 0.754
R13174 out_p.n939 out_p.n938 0.754
R13175 out_p.n958 out_p.n957 0.754
R13176 out_p.n957 out_p.n956 0.754
R13177 out_p.n956 out_p.n955 0.754
R13178 out_p.n955 out_p.n954 0.754
R13179 out_p.n953 out_p.n952 0.754
R13180 out_p.n952 out_p.n951 0.754
R13181 out_p.n951 out_p.n950 0.754
R13182 out_p.n950 out_p.n949 0.754
R13183 out_p.n969 out_p.n968 0.754
R13184 out_p.n968 out_p.n967 0.754
R13185 out_p.n967 out_p.n966 0.754
R13186 out_p.n966 out_p.n965 0.754
R13187 out_p.n964 out_p.n963 0.754
R13188 out_p.n963 out_p.n962 0.754
R13189 out_p.n962 out_p.n961 0.754
R13190 out_p.n961 out_p.n960 0.754
R13191 out_p.n19 out_p.n18 0.754
R13192 out_p.n18 out_p.n17 0.754
R13193 out_p.n17 out_p.n16 0.754
R13194 out_p.n16 out_p.n15 0.754
R13195 out_p.n14 out_p.n13 0.754
R13196 out_p.n13 out_p.n12 0.754
R13197 out_p.n12 out_p.n11 0.754
R13198 out_p.n11 out_p.n10 0.754
R13199 out_p.n33 out_p.n32 0.754
R13200 out_p.n32 out_p.n31 0.754
R13201 out_p.n31 out_p.n30 0.754
R13202 out_p.n30 out_p.n29 0.754
R13203 out_p.n28 out_p.n27 0.754
R13204 out_p.n27 out_p.n26 0.754
R13205 out_p.n26 out_p.n25 0.754
R13206 out_p.n25 out_p.n24 0.754
R13207 out_p.n45 out_p.n44 0.754
R13208 out_p.n44 out_p.n43 0.754
R13209 out_p.n43 out_p.n42 0.754
R13210 out_p.n42 out_p.n41 0.754
R13211 out_p.n40 out_p.n39 0.754
R13212 out_p.n39 out_p.n38 0.754
R13213 out_p.n38 out_p.n37 0.754
R13214 out_p.n37 out_p.n36 0.754
R13215 out_p.n57 out_p.n56 0.754
R13216 out_p.n56 out_p.n55 0.754
R13217 out_p.n55 out_p.n54 0.754
R13218 out_p.n54 out_p.n53 0.754
R13219 out_p.n52 out_p.n51 0.754
R13220 out_p.n51 out_p.n50 0.754
R13221 out_p.n50 out_p.n49 0.754
R13222 out_p.n49 out_p.n48 0.754
R13223 out_p.n69 out_p.n68 0.754
R13224 out_p.n68 out_p.n67 0.754
R13225 out_p.n67 out_p.n66 0.754
R13226 out_p.n66 out_p.n65 0.754
R13227 out_p.n64 out_p.n63 0.754
R13228 out_p.n63 out_p.n62 0.754
R13229 out_p.n62 out_p.n61 0.754
R13230 out_p.n61 out_p.n60 0.754
R13231 out_p.n81 out_p.n80 0.754
R13232 out_p.n80 out_p.n79 0.754
R13233 out_p.n79 out_p.n78 0.754
R13234 out_p.n78 out_p.n77 0.754
R13235 out_p.n76 out_p.n75 0.754
R13236 out_p.n75 out_p.n74 0.754
R13237 out_p.n74 out_p.n73 0.754
R13238 out_p.n73 out_p.n72 0.754
R13239 out_p.n93 out_p.n92 0.754
R13240 out_p.n92 out_p.n91 0.754
R13241 out_p.n91 out_p.n90 0.754
R13242 out_p.n90 out_p.n89 0.754
R13243 out_p.n88 out_p.n87 0.754
R13244 out_p.n87 out_p.n86 0.754
R13245 out_p.n86 out_p.n85 0.754
R13246 out_p.n85 out_p.n84 0.754
R13247 out_p.n105 out_p.n104 0.754
R13248 out_p.n104 out_p.n103 0.754
R13249 out_p.n103 out_p.n102 0.754
R13250 out_p.n102 out_p.n101 0.754
R13251 out_p.n100 out_p.n99 0.754
R13252 out_p.n99 out_p.n98 0.754
R13253 out_p.n98 out_p.n97 0.754
R13254 out_p.n97 out_p.n96 0.754
R13255 out_p.n117 out_p.n116 0.754
R13256 out_p.n116 out_p.n115 0.754
R13257 out_p.n115 out_p.n114 0.754
R13258 out_p.n114 out_p.n113 0.754
R13259 out_p.n112 out_p.n111 0.754
R13260 out_p.n111 out_p.n110 0.754
R13261 out_p.n110 out_p.n109 0.754
R13262 out_p.n109 out_p.n108 0.754
R13263 out_p.n129 out_p.n128 0.754
R13264 out_p.n128 out_p.n127 0.754
R13265 out_p.n127 out_p.n126 0.754
R13266 out_p.n126 out_p.n125 0.754
R13267 out_p.n124 out_p.n123 0.754
R13268 out_p.n123 out_p.n122 0.754
R13269 out_p.n122 out_p.n121 0.754
R13270 out_p.n121 out_p.n120 0.754
R13271 out_p.n141 out_p.n140 0.754
R13272 out_p.n140 out_p.n139 0.754
R13273 out_p.n139 out_p.n138 0.754
R13274 out_p.n138 out_p.n137 0.754
R13275 out_p.n136 out_p.n135 0.754
R13276 out_p.n135 out_p.n134 0.754
R13277 out_p.n134 out_p.n133 0.754
R13278 out_p.n133 out_p.n132 0.754
R13279 out_p.n153 out_p.n152 0.754
R13280 out_p.n152 out_p.n151 0.754
R13281 out_p.n151 out_p.n150 0.754
R13282 out_p.n150 out_p.n149 0.754
R13283 out_p.n148 out_p.n147 0.754
R13284 out_p.n147 out_p.n146 0.754
R13285 out_p.n146 out_p.n145 0.754
R13286 out_p.n145 out_p.n144 0.754
R13287 out_p.n165 out_p.n164 0.754
R13288 out_p.n164 out_p.n163 0.754
R13289 out_p.n163 out_p.n162 0.754
R13290 out_p.n162 out_p.n161 0.754
R13291 out_p.n160 out_p.n159 0.754
R13292 out_p.n159 out_p.n158 0.754
R13293 out_p.n158 out_p.n157 0.754
R13294 out_p.n157 out_p.n156 0.754
R13295 out_p.n177 out_p.n176 0.754
R13296 out_p.n176 out_p.n175 0.754
R13297 out_p.n175 out_p.n174 0.754
R13298 out_p.n174 out_p.n173 0.754
R13299 out_p.n172 out_p.n171 0.754
R13300 out_p.n171 out_p.n170 0.754
R13301 out_p.n170 out_p.n169 0.754
R13302 out_p.n169 out_p.n168 0.754
R13303 out_p.n189 out_p.n188 0.754
R13304 out_p.n188 out_p.n187 0.754
R13305 out_p.n187 out_p.n186 0.754
R13306 out_p.n186 out_p.n185 0.754
R13307 out_p.n184 out_p.n183 0.754
R13308 out_p.n183 out_p.n182 0.754
R13309 out_p.n182 out_p.n181 0.754
R13310 out_p.n181 out_p.n180 0.754
R13311 out_p.n201 out_p.n200 0.754
R13312 out_p.n200 out_p.n199 0.754
R13313 out_p.n199 out_p.n198 0.754
R13314 out_p.n198 out_p.n197 0.754
R13315 out_p.n196 out_p.n195 0.754
R13316 out_p.n195 out_p.n194 0.754
R13317 out_p.n194 out_p.n193 0.754
R13318 out_p.n193 out_p.n192 0.754
R13319 out_p.n213 out_p.n212 0.754
R13320 out_p.n212 out_p.n211 0.754
R13321 out_p.n211 out_p.n210 0.754
R13322 out_p.n210 out_p.n209 0.754
R13323 out_p.n208 out_p.n207 0.754
R13324 out_p.n207 out_p.n206 0.754
R13325 out_p.n206 out_p.n205 0.754
R13326 out_p.n205 out_p.n204 0.754
R13327 out_p.n225 out_p.n224 0.754
R13328 out_p.n224 out_p.n223 0.754
R13329 out_p.n223 out_p.n222 0.754
R13330 out_p.n222 out_p.n221 0.754
R13331 out_p.n220 out_p.n219 0.754
R13332 out_p.n219 out_p.n218 0.754
R13333 out_p.n218 out_p.n217 0.754
R13334 out_p.n217 out_p.n216 0.754
R13335 out_p.n237 out_p.n236 0.754
R13336 out_p.n236 out_p.n235 0.754
R13337 out_p.n235 out_p.n234 0.754
R13338 out_p.n234 out_p.n233 0.754
R13339 out_p.n232 out_p.n231 0.754
R13340 out_p.n231 out_p.n230 0.754
R13341 out_p.n230 out_p.n229 0.754
R13342 out_p.n229 out_p.n228 0.754
R13343 out_p.n249 out_p.n248 0.754
R13344 out_p.n248 out_p.n247 0.754
R13345 out_p.n247 out_p.n246 0.754
R13346 out_p.n246 out_p.n245 0.754
R13347 out_p.n244 out_p.n243 0.754
R13348 out_p.n243 out_p.n242 0.754
R13349 out_p.n242 out_p.n241 0.754
R13350 out_p.n241 out_p.n240 0.754
R13351 out_p.n261 out_p.n260 0.754
R13352 out_p.n260 out_p.n259 0.754
R13353 out_p.n259 out_p.n258 0.754
R13354 out_p.n258 out_p.n257 0.754
R13355 out_p.n256 out_p.n255 0.754
R13356 out_p.n255 out_p.n254 0.754
R13357 out_p.n254 out_p.n253 0.754
R13358 out_p.n253 out_p.n252 0.754
R13359 out_p.n273 out_p.n272 0.754
R13360 out_p.n272 out_p.n271 0.754
R13361 out_p.n271 out_p.n270 0.754
R13362 out_p.n270 out_p.n269 0.754
R13363 out_p.n268 out_p.n267 0.754
R13364 out_p.n267 out_p.n266 0.754
R13365 out_p.n266 out_p.n265 0.754
R13366 out_p.n265 out_p.n264 0.754
R13367 out_p.n285 out_p.n284 0.754
R13368 out_p.n284 out_p.n283 0.754
R13369 out_p.n283 out_p.n282 0.754
R13370 out_p.n282 out_p.n281 0.754
R13371 out_p.n280 out_p.n279 0.754
R13372 out_p.n279 out_p.n278 0.754
R13373 out_p.n278 out_p.n277 0.754
R13374 out_p.n277 out_p.n276 0.754
R13375 out_p.n297 out_p.n296 0.754
R13376 out_p.n296 out_p.n295 0.754
R13377 out_p.n295 out_p.n294 0.754
R13378 out_p.n294 out_p.n293 0.754
R13379 out_p.n292 out_p.n291 0.754
R13380 out_p.n291 out_p.n290 0.754
R13381 out_p.n290 out_p.n289 0.754
R13382 out_p.n289 out_p.n288 0.754
R13383 out_p.n309 out_p.n308 0.754
R13384 out_p.n308 out_p.n307 0.754
R13385 out_p.n307 out_p.n306 0.754
R13386 out_p.n306 out_p.n305 0.754
R13387 out_p.n304 out_p.n303 0.754
R13388 out_p.n303 out_p.n302 0.754
R13389 out_p.n302 out_p.n301 0.754
R13390 out_p.n301 out_p.n300 0.754
R13391 out_p.n321 out_p.n320 0.754
R13392 out_p.n320 out_p.n319 0.754
R13393 out_p.n319 out_p.n318 0.754
R13394 out_p.n318 out_p.n317 0.754
R13395 out_p.n316 out_p.n315 0.754
R13396 out_p.n315 out_p.n314 0.754
R13397 out_p.n314 out_p.n313 0.754
R13398 out_p.n313 out_p.n312 0.754
R13399 out_p.n333 out_p.n332 0.754
R13400 out_p.n332 out_p.n331 0.754
R13401 out_p.n331 out_p.n330 0.754
R13402 out_p.n330 out_p.n329 0.754
R13403 out_p.n328 out_p.n327 0.754
R13404 out_p.n327 out_p.n326 0.754
R13405 out_p.n326 out_p.n325 0.754
R13406 out_p.n325 out_p.n324 0.754
R13407 out_p.n345 out_p.n344 0.754
R13408 out_p.n344 out_p.n343 0.754
R13409 out_p.n343 out_p.n342 0.754
R13410 out_p.n342 out_p.n341 0.754
R13411 out_p.n340 out_p.n339 0.754
R13412 out_p.n339 out_p.n338 0.754
R13413 out_p.n338 out_p.n337 0.754
R13414 out_p.n337 out_p.n336 0.754
R13415 out_p.n357 out_p.n356 0.754
R13416 out_p.n356 out_p.n355 0.754
R13417 out_p.n355 out_p.n354 0.754
R13418 out_p.n354 out_p.n353 0.754
R13419 out_p.n352 out_p.n351 0.754
R13420 out_p.n351 out_p.n350 0.754
R13421 out_p.n350 out_p.n349 0.754
R13422 out_p.n349 out_p.n348 0.754
R13423 out_p.n369 out_p.n368 0.754
R13424 out_p.n368 out_p.n367 0.754
R13425 out_p.n367 out_p.n366 0.754
R13426 out_p.n366 out_p.n365 0.754
R13427 out_p.n364 out_p.n363 0.754
R13428 out_p.n363 out_p.n362 0.754
R13429 out_p.n362 out_p.n361 0.754
R13430 out_p.n361 out_p.n360 0.754
R13431 out_p.n381 out_p.n380 0.754
R13432 out_p.n380 out_p.n379 0.754
R13433 out_p.n379 out_p.n378 0.754
R13434 out_p.n378 out_p.n377 0.754
R13435 out_p.n376 out_p.n375 0.754
R13436 out_p.n375 out_p.n374 0.754
R13437 out_p.n374 out_p.n373 0.754
R13438 out_p.n373 out_p.n372 0.754
R13439 out_p.n393 out_p.n392 0.754
R13440 out_p.n392 out_p.n391 0.754
R13441 out_p.n391 out_p.n390 0.754
R13442 out_p.n390 out_p.n389 0.754
R13443 out_p.n388 out_p.n387 0.754
R13444 out_p.n387 out_p.n386 0.754
R13445 out_p.n386 out_p.n385 0.754
R13446 out_p.n385 out_p.n384 0.754
R13447 out_p.n405 out_p.n404 0.754
R13448 out_p.n404 out_p.n403 0.754
R13449 out_p.n403 out_p.n402 0.754
R13450 out_p.n402 out_p.n401 0.754
R13451 out_p.n400 out_p.n399 0.754
R13452 out_p.n399 out_p.n398 0.754
R13453 out_p.n398 out_p.n397 0.754
R13454 out_p.n397 out_p.n396 0.754
R13455 out_p.n417 out_p.n416 0.754
R13456 out_p.n416 out_p.n415 0.754
R13457 out_p.n415 out_p.n414 0.754
R13458 out_p.n414 out_p.n413 0.754
R13459 out_p.n412 out_p.n411 0.754
R13460 out_p.n411 out_p.n410 0.754
R13461 out_p.n410 out_p.n409 0.754
R13462 out_p.n409 out_p.n408 0.754
R13463 out_p.n429 out_p.n428 0.754
R13464 out_p.n428 out_p.n427 0.754
R13465 out_p.n427 out_p.n426 0.754
R13466 out_p.n426 out_p.n425 0.754
R13467 out_p.n424 out_p.n423 0.754
R13468 out_p.n423 out_p.n422 0.754
R13469 out_p.n422 out_p.n421 0.754
R13470 out_p.n421 out_p.n420 0.754
R13471 out_p.n441 out_p.n440 0.754
R13472 out_p.n440 out_p.n439 0.754
R13473 out_p.n439 out_p.n438 0.754
R13474 out_p.n438 out_p.n437 0.754
R13475 out_p.n436 out_p.n435 0.754
R13476 out_p.n435 out_p.n434 0.754
R13477 out_p.n434 out_p.n433 0.754
R13478 out_p.n433 out_p.n432 0.754
R13479 out_p.n453 out_p.n452 0.754
R13480 out_p.n452 out_p.n451 0.754
R13481 out_p.n451 out_p.n450 0.754
R13482 out_p.n450 out_p.n449 0.754
R13483 out_p.n448 out_p.n447 0.754
R13484 out_p.n447 out_p.n446 0.754
R13485 out_p.n446 out_p.n445 0.754
R13486 out_p.n445 out_p.n444 0.754
R13487 out_p.n465 out_p.n464 0.754
R13488 out_p.n464 out_p.n463 0.754
R13489 out_p.n463 out_p.n462 0.754
R13490 out_p.n462 out_p.n461 0.754
R13491 out_p.n460 out_p.n459 0.754
R13492 out_p.n459 out_p.n458 0.754
R13493 out_p.n458 out_p.n457 0.754
R13494 out_p.n457 out_p.n456 0.754
R13495 out_p.n477 out_p.n476 0.754
R13496 out_p.n476 out_p.n475 0.754
R13497 out_p.n475 out_p.n474 0.754
R13498 out_p.n474 out_p.n473 0.754
R13499 out_p.n472 out_p.n471 0.754
R13500 out_p.n471 out_p.n470 0.754
R13501 out_p.n470 out_p.n469 0.754
R13502 out_p.n469 out_p.n468 0.754
R13503 out_p.n489 out_p.n488 0.754
R13504 out_p.n488 out_p.n487 0.754
R13505 out_p.n487 out_p.n486 0.754
R13506 out_p.n486 out_p.n485 0.754
R13507 out_p.n484 out_p.n483 0.754
R13508 out_p.n483 out_p.n482 0.754
R13509 out_p.n482 out_p.n481 0.754
R13510 out_p.n481 out_p.n480 0.754
R13511 out_p.n501 out_p.n500 0.754
R13512 out_p.n500 out_p.n499 0.754
R13513 out_p.n499 out_p.n498 0.754
R13514 out_p.n498 out_p.n497 0.754
R13515 out_p.n496 out_p.n495 0.754
R13516 out_p.n495 out_p.n494 0.754
R13517 out_p.n494 out_p.n493 0.754
R13518 out_p.n493 out_p.n492 0.754
R13519 out_p.n513 out_p.n512 0.754
R13520 out_p.n512 out_p.n511 0.754
R13521 out_p.n511 out_p.n510 0.754
R13522 out_p.n510 out_p.n509 0.754
R13523 out_p.n508 out_p.n507 0.754
R13524 out_p.n507 out_p.n506 0.754
R13525 out_p.n506 out_p.n505 0.754
R13526 out_p.n505 out_p.n504 0.754
R13527 out_p.n525 out_p.n524 0.754
R13528 out_p.n524 out_p.n523 0.754
R13529 out_p.n523 out_p.n522 0.754
R13530 out_p.n522 out_p.n521 0.754
R13531 out_p.n520 out_p.n519 0.754
R13532 out_p.n519 out_p.n518 0.754
R13533 out_p.n518 out_p.n517 0.754
R13534 out_p.n517 out_p.n516 0.754
R13535 out_p.n537 out_p.n536 0.754
R13536 out_p.n536 out_p.n535 0.754
R13537 out_p.n535 out_p.n534 0.754
R13538 out_p.n534 out_p.n533 0.754
R13539 out_p.n532 out_p.n531 0.754
R13540 out_p.n531 out_p.n530 0.754
R13541 out_p.n530 out_p.n529 0.754
R13542 out_p.n529 out_p.n528 0.754
R13543 out_p.n549 out_p.n548 0.754
R13544 out_p.n548 out_p.n547 0.754
R13545 out_p.n547 out_p.n546 0.754
R13546 out_p.n546 out_p.n545 0.754
R13547 out_p.n544 out_p.n543 0.754
R13548 out_p.n543 out_p.n542 0.754
R13549 out_p.n542 out_p.n541 0.754
R13550 out_p.n541 out_p.n540 0.754
R13551 out_p.n561 out_p.n560 0.754
R13552 out_p.n560 out_p.n559 0.754
R13553 out_p.n559 out_p.n558 0.754
R13554 out_p.n558 out_p.n557 0.754
R13555 out_p.n556 out_p.n555 0.754
R13556 out_p.n555 out_p.n554 0.754
R13557 out_p.n554 out_p.n553 0.754
R13558 out_p.n553 out_p.n552 0.754
R13559 out_p.n573 out_p.n572 0.754
R13560 out_p.n572 out_p.n571 0.754
R13561 out_p.n571 out_p.n570 0.754
R13562 out_p.n570 out_p.n569 0.754
R13563 out_p.n568 out_p.n567 0.754
R13564 out_p.n567 out_p.n566 0.754
R13565 out_p.n566 out_p.n565 0.754
R13566 out_p.n565 out_p.n564 0.754
R13567 out_p.n585 out_p.n584 0.754
R13568 out_p.n584 out_p.n583 0.754
R13569 out_p.n583 out_p.n582 0.754
R13570 out_p.n582 out_p.n581 0.754
R13571 out_p.n580 out_p.n579 0.754
R13572 out_p.n579 out_p.n578 0.754
R13573 out_p.n578 out_p.n577 0.754
R13574 out_p.n577 out_p.n576 0.754
R13575 out_p.n597 out_p.n596 0.754
R13576 out_p.n596 out_p.n595 0.754
R13577 out_p.n595 out_p.n594 0.754
R13578 out_p.n594 out_p.n593 0.754
R13579 out_p.n592 out_p.n591 0.754
R13580 out_p.n591 out_p.n590 0.754
R13581 out_p.n590 out_p.n589 0.754
R13582 out_p.n589 out_p.n588 0.754
R13583 out_p.n609 out_p.n608 0.754
R13584 out_p.n608 out_p.n607 0.754
R13585 out_p.n607 out_p.n606 0.754
R13586 out_p.n606 out_p.n605 0.754
R13587 out_p.n604 out_p.n603 0.754
R13588 out_p.n603 out_p.n602 0.754
R13589 out_p.n602 out_p.n601 0.754
R13590 out_p.n601 out_p.n600 0.754
R13591 out_p.n621 out_p.n620 0.754
R13592 out_p.n620 out_p.n619 0.754
R13593 out_p.n619 out_p.n618 0.754
R13594 out_p.n618 out_p.n617 0.754
R13595 out_p.n616 out_p.n615 0.754
R13596 out_p.n615 out_p.n614 0.754
R13597 out_p.n614 out_p.n613 0.754
R13598 out_p.n613 out_p.n612 0.754
R13599 out_p.n633 out_p.n632 0.754
R13600 out_p.n632 out_p.n631 0.754
R13601 out_p.n631 out_p.n630 0.754
R13602 out_p.n630 out_p.n629 0.754
R13603 out_p.n628 out_p.n627 0.754
R13604 out_p.n627 out_p.n626 0.754
R13605 out_p.n626 out_p.n625 0.754
R13606 out_p.n625 out_p.n624 0.754
R13607 out_p.n645 out_p.n644 0.754
R13608 out_p.n644 out_p.n643 0.754
R13609 out_p.n643 out_p.n642 0.754
R13610 out_p.n642 out_p.n641 0.754
R13611 out_p.n640 out_p.n639 0.754
R13612 out_p.n639 out_p.n638 0.754
R13613 out_p.n638 out_p.n637 0.754
R13614 out_p.n637 out_p.n636 0.754
R13615 out_p.n657 out_p.n656 0.754
R13616 out_p.n656 out_p.n655 0.754
R13617 out_p.n655 out_p.n654 0.754
R13618 out_p.n654 out_p.n653 0.754
R13619 out_p.n652 out_p.n651 0.754
R13620 out_p.n651 out_p.n650 0.754
R13621 out_p.n650 out_p.n649 0.754
R13622 out_p.n649 out_p.n648 0.754
R13623 out_p.n669 out_p.n668 0.754
R13624 out_p.n668 out_p.n667 0.754
R13625 out_p.n667 out_p.n666 0.754
R13626 out_p.n666 out_p.n665 0.754
R13627 out_p.n664 out_p.n663 0.754
R13628 out_p.n663 out_p.n662 0.754
R13629 out_p.n662 out_p.n661 0.754
R13630 out_p.n661 out_p.n660 0.754
R13631 out_p.n681 out_p.n680 0.754
R13632 out_p.n680 out_p.n679 0.754
R13633 out_p.n679 out_p.n678 0.754
R13634 out_p.n678 out_p.n677 0.754
R13635 out_p.n676 out_p.n675 0.754
R13636 out_p.n675 out_p.n674 0.754
R13637 out_p.n674 out_p.n673 0.754
R13638 out_p.n673 out_p.n672 0.754
R13639 out_p.n693 out_p.n692 0.754
R13640 out_p.n692 out_p.n691 0.754
R13641 out_p.n691 out_p.n690 0.754
R13642 out_p.n690 out_p.n689 0.754
R13643 out_p.n688 out_p.n687 0.754
R13644 out_p.n687 out_p.n686 0.754
R13645 out_p.n686 out_p.n685 0.754
R13646 out_p.n685 out_p.n684 0.754
R13647 out_p.n705 out_p.n704 0.754
R13648 out_p.n704 out_p.n703 0.754
R13649 out_p.n703 out_p.n702 0.754
R13650 out_p.n702 out_p.n701 0.754
R13651 out_p.n700 out_p.n699 0.754
R13652 out_p.n699 out_p.n698 0.754
R13653 out_p.n698 out_p.n697 0.754
R13654 out_p.n697 out_p.n696 0.754
R13655 out_p.n717 out_p.n716 0.754
R13656 out_p.n716 out_p.n715 0.754
R13657 out_p.n715 out_p.n714 0.754
R13658 out_p.n714 out_p.n713 0.754
R13659 out_p.n712 out_p.n711 0.754
R13660 out_p.n711 out_p.n710 0.754
R13661 out_p.n710 out_p.n709 0.754
R13662 out_p.n709 out_p.n708 0.754
R13663 out_p.n729 out_p.n728 0.754
R13664 out_p.n728 out_p.n727 0.754
R13665 out_p.n727 out_p.n726 0.754
R13666 out_p.n726 out_p.n725 0.754
R13667 out_p.n724 out_p.n723 0.754
R13668 out_p.n723 out_p.n722 0.754
R13669 out_p.n722 out_p.n721 0.754
R13670 out_p.n721 out_p.n720 0.754
R13671 out_p.n9 out_p.n8 0.754
R13672 out_p.n8 out_p.n7 0.754
R13673 out_p.n7 out_p.n6 0.754
R13674 out_p.n6 out_p.n5 0.754
R13675 out_p.n4 out_p.n3 0.754
R13676 out_p.n3 out_p.n2 0.754
R13677 out_p.n2 out_p.n1 0.754
R13678 out_p.n1 out_p.n0 0.754
R13679 out_p.n742 out_p.n731 0.554
R13680 out_p.n743 out_p.n719 0.554
R13681 out_p.n744 out_p.n707 0.554
R13682 out_p.n745 out_p.n695 0.554
R13683 out_p.n746 out_p.n683 0.554
R13684 out_p.n747 out_p.n671 0.554
R13685 out_p.n748 out_p.n659 0.554
R13686 out_p.n749 out_p.n647 0.554
R13687 out_p.n750 out_p.n635 0.554
R13688 out_p.n751 out_p.n623 0.554
R13689 out_p.n752 out_p.n611 0.554
R13690 out_p.n753 out_p.n599 0.554
R13691 out_p.n754 out_p.n587 0.554
R13692 out_p.n755 out_p.n575 0.554
R13693 out_p.n756 out_p.n563 0.554
R13694 out_p.n757 out_p.n551 0.554
R13695 out_p.n758 out_p.n539 0.554
R13696 out_p.n759 out_p.n527 0.554
R13697 out_p.n760 out_p.n515 0.554
R13698 out_p.n761 out_p.n503 0.554
R13699 out_p.n762 out_p.n491 0.554
R13700 out_p.n763 out_p.n479 0.554
R13701 out_p.n764 out_p.n467 0.554
R13702 out_p.n765 out_p.n455 0.554
R13703 out_p.n766 out_p.n443 0.554
R13704 out_p.n767 out_p.n431 0.554
R13705 out_p.n768 out_p.n419 0.554
R13706 out_p.n769 out_p.n407 0.554
R13707 out_p.n770 out_p.n395 0.554
R13708 out_p.n771 out_p.n383 0.554
R13709 out_p.n772 out_p.n371 0.554
R13710 out_p.n773 out_p.n359 0.554
R13711 out_p.n774 out_p.n347 0.554
R13712 out_p.n775 out_p.n335 0.554
R13713 out_p.n776 out_p.n323 0.554
R13714 out_p.n777 out_p.n311 0.554
R13715 out_p.n778 out_p.n299 0.554
R13716 out_p.n779 out_p.n287 0.554
R13717 out_p.n780 out_p.n275 0.554
R13718 out_p.n781 out_p.n263 0.554
R13719 out_p.n782 out_p.n251 0.554
R13720 out_p.n783 out_p.n239 0.554
R13721 out_p.n784 out_p.n227 0.554
R13722 out_p.n785 out_p.n215 0.554
R13723 out_p.n786 out_p.n203 0.554
R13724 out_p.n787 out_p.n191 0.554
R13725 out_p.n788 out_p.n179 0.554
R13726 out_p.n789 out_p.n167 0.554
R13727 out_p.n790 out_p.n155 0.554
R13728 out_p.n791 out_p.n143 0.554
R13729 out_p.n792 out_p.n131 0.554
R13730 out_p.n793 out_p.n119 0.554
R13731 out_p.n794 out_p.n107 0.554
R13732 out_p.n795 out_p.n95 0.554
R13733 out_p.n796 out_p.n83 0.554
R13734 out_p.n797 out_p.n71 0.554
R13735 out_p.n798 out_p.n59 0.554
R13736 out_p.n799 out_p.n47 0.554
R13737 out_p.n800 out_p.n35 0.554
R13738 out_p.n801 out_p.n23 0.554
R13739 out_p out_p.n21 0.554
R13740 out_p.n970 out_p.n803 0.554
R13741 out_p.n959 out_p.n805 0.554
R13742 out_p.n948 out_p.n807 0.554
R13743 out_p.n937 out_p.n809 0.554
R13744 out_p.n926 out_p.n811 0.554
R13745 out_p.n915 out_p.n813 0.554
R13746 out_p.n904 out_p.n815 0.554
R13747 out_p.n893 out_p.n817 0.554
R13748 out_p.n882 out_p.n819 0.554
R13749 out_p.n871 out_p.n821 0.554
R13750 out_p.n860 out_p.n823 0.554
R13751 out_p.n849 out_p.n825 0.554
R13752 out_p.n838 out_p.n827 0.554
R13753 out_p.n973 out_p.n972 0.554
R13754 out_p.n742 out_p.n741 0.541
R13755 out_p.n838 out_p.n837 0.524
R13756 out_p.n849 out_p.n848 0.524
R13757 out_p.n860 out_p.n859 0.524
R13758 out_p.n871 out_p.n870 0.524
R13759 out_p.n882 out_p.n881 0.524
R13760 out_p.n893 out_p.n892 0.524
R13761 out_p.n904 out_p.n903 0.524
R13762 out_p.n915 out_p.n914 0.524
R13763 out_p.n926 out_p.n925 0.524
R13764 out_p.n937 out_p.n936 0.524
R13765 out_p.n948 out_p.n947 0.524
R13766 out_p.n959 out_p.n958 0.524
R13767 out_p.n970 out_p.n969 0.524
R13768 out_p out_p.n19 0.524
R13769 out_p.n801 out_p.n33 0.524
R13770 out_p.n800 out_p.n45 0.524
R13771 out_p.n799 out_p.n57 0.524
R13772 out_p.n798 out_p.n69 0.524
R13773 out_p.n797 out_p.n81 0.524
R13774 out_p.n796 out_p.n93 0.524
R13775 out_p.n795 out_p.n105 0.524
R13776 out_p.n794 out_p.n117 0.524
R13777 out_p.n793 out_p.n129 0.524
R13778 out_p.n792 out_p.n141 0.524
R13779 out_p.n791 out_p.n153 0.524
R13780 out_p.n790 out_p.n165 0.524
R13781 out_p.n789 out_p.n177 0.524
R13782 out_p.n788 out_p.n189 0.524
R13783 out_p.n787 out_p.n201 0.524
R13784 out_p.n786 out_p.n213 0.524
R13785 out_p.n785 out_p.n225 0.524
R13786 out_p.n784 out_p.n237 0.524
R13787 out_p.n783 out_p.n249 0.524
R13788 out_p.n782 out_p.n261 0.524
R13789 out_p.n781 out_p.n273 0.524
R13790 out_p.n780 out_p.n285 0.524
R13791 out_p.n779 out_p.n297 0.524
R13792 out_p.n778 out_p.n309 0.524
R13793 out_p.n777 out_p.n321 0.524
R13794 out_p.n776 out_p.n333 0.524
R13795 out_p.n775 out_p.n345 0.524
R13796 out_p.n774 out_p.n357 0.524
R13797 out_p.n773 out_p.n369 0.524
R13798 out_p.n772 out_p.n381 0.524
R13799 out_p.n771 out_p.n393 0.524
R13800 out_p.n770 out_p.n405 0.524
R13801 out_p.n769 out_p.n417 0.524
R13802 out_p.n768 out_p.n429 0.524
R13803 out_p.n767 out_p.n441 0.524
R13804 out_p.n766 out_p.n453 0.524
R13805 out_p.n765 out_p.n465 0.524
R13806 out_p.n764 out_p.n477 0.524
R13807 out_p.n763 out_p.n489 0.524
R13808 out_p.n762 out_p.n501 0.524
R13809 out_p.n761 out_p.n513 0.524
R13810 out_p.n760 out_p.n525 0.524
R13811 out_p.n759 out_p.n537 0.524
R13812 out_p.n758 out_p.n549 0.524
R13813 out_p.n757 out_p.n561 0.524
R13814 out_p.n756 out_p.n573 0.524
R13815 out_p.n755 out_p.n585 0.524
R13816 out_p.n754 out_p.n597 0.524
R13817 out_p.n753 out_p.n609 0.524
R13818 out_p.n752 out_p.n621 0.524
R13819 out_p.n751 out_p.n633 0.524
R13820 out_p.n750 out_p.n645 0.524
R13821 out_p.n749 out_p.n657 0.524
R13822 out_p.n748 out_p.n669 0.524
R13823 out_p.n747 out_p.n681 0.524
R13824 out_p.n746 out_p.n693 0.524
R13825 out_p.n745 out_p.n705 0.524
R13826 out_p.n744 out_p.n717 0.524
R13827 out_p.n743 out_p.n729 0.524
R13828 out_p.n973 out_p.n9 0.524
R13829 out_p.n849 out_p.n838 0.002
R13830 out_p.n860 out_p.n849 0.002
R13831 out_p.n871 out_p.n860 0.002
R13832 out_p.n882 out_p.n871 0.002
R13833 out_p.n893 out_p.n882 0.002
R13834 out_p.n904 out_p.n893 0.002
R13835 out_p.n915 out_p.n904 0.002
R13836 out_p.n926 out_p.n915 0.002
R13837 out_p.n937 out_p.n926 0.002
R13838 out_p.n948 out_p.n937 0.002
R13839 out_p.n959 out_p.n948 0.002
R13840 out_p.n970 out_p.n959 0.002
R13841 out_p.n973 out_p.n970 0.002
R13842 out_p.n973 out_p 0.002
R13843 out_p out_p.n801 0.002
R13844 out_p.n801 out_p.n800 0.002
R13845 out_p.n800 out_p.n799 0.002
R13846 out_p.n799 out_p.n798 0.002
R13847 out_p.n798 out_p.n797 0.002
R13848 out_p.n797 out_p.n796 0.002
R13849 out_p.n796 out_p.n795 0.002
R13850 out_p.n795 out_p.n794 0.002
R13851 out_p.n794 out_p.n793 0.002
R13852 out_p.n793 out_p.n792 0.002
R13853 out_p.n792 out_p.n791 0.002
R13854 out_p.n791 out_p.n790 0.002
R13855 out_p.n790 out_p.n789 0.002
R13856 out_p.n789 out_p.n788 0.002
R13857 out_p.n788 out_p.n787 0.002
R13858 out_p.n787 out_p.n786 0.002
R13859 out_p.n786 out_p.n785 0.002
R13860 out_p.n785 out_p.n784 0.002
R13861 out_p.n784 out_p.n783 0.002
R13862 out_p.n783 out_p.n782 0.002
R13863 out_p.n782 out_p.n781 0.002
R13864 out_p.n781 out_p.n780 0.002
R13865 out_p.n780 out_p.n779 0.002
R13866 out_p.n779 out_p.n778 0.002
R13867 out_p.n778 out_p.n777 0.002
R13868 out_p.n777 out_p.n776 0.002
R13869 out_p.n776 out_p.n775 0.002
R13870 out_p.n775 out_p.n774 0.002
R13871 out_p.n774 out_p.n773 0.002
R13872 out_p.n773 out_p.n772 0.002
R13873 out_p.n772 out_p.n771 0.002
R13874 out_p.n771 out_p.n770 0.002
R13875 out_p.n770 out_p.n769 0.002
R13876 out_p.n769 out_p.n768 0.002
R13877 out_p.n768 out_p.n767 0.002
R13878 out_p.n767 out_p.n766 0.002
R13879 out_p.n766 out_p.n765 0.002
R13880 out_p.n765 out_p.n764 0.002
R13881 out_p.n764 out_p.n763 0.002
R13882 out_p.n763 out_p.n762 0.002
R13883 out_p.n762 out_p.n761 0.002
R13884 out_p.n761 out_p.n760 0.002
R13885 out_p.n760 out_p.n759 0.002
R13886 out_p.n759 out_p.n758 0.002
R13887 out_p.n758 out_p.n757 0.002
R13888 out_p.n757 out_p.n756 0.002
R13889 out_p.n756 out_p.n755 0.002
R13890 out_p.n755 out_p.n754 0.002
R13891 out_p.n754 out_p.n753 0.002
R13892 out_p.n753 out_p.n752 0.002
R13893 out_p.n752 out_p.n751 0.002
R13894 out_p.n751 out_p.n750 0.002
R13895 out_p.n750 out_p.n749 0.002
R13896 out_p.n749 out_p.n748 0.002
R13897 out_p.n748 out_p.n747 0.002
R13898 out_p.n747 out_p.n746 0.002
R13899 out_p.n746 out_p.n745 0.002
R13900 out_p.n745 out_p.n744 0.002
R13901 out_p.n744 out_p.n743 0.002
R13902 out_p.n743 out_p.n742 0.002
R13903 vdd1.n17 vdd1.n16 9250.59
R13904 vdd1.n23 vdd1.n22 9250.59
R13905 vdd1.n15 vdd1.n14 2878.29
R13906 vdd1.n21 vdd1.n20 2869.55
R13907 vdd1.n24 vdd1.n17 2247.42
R13908 vdd1.n24 vdd1.n23 2247.42
R13909 vdd1.n21 vdd1.n18 940.477
R13910 vdd1.n15 vdd1.n12 940.476
R13911 vdd1.n23 vdd1.n21 940.476
R13912 vdd1.n17 vdd1.n15 940.476
R13913 vdd1.n491 vdd1.t1404 10.284
R13914 vdd1.n38 vdd1.t823 8.711
R13915 vdd1.n46 vdd1.t69 8.131
R13916 vdd1.n45 vdd1.t189 8.131
R13917 vdd1.n44 vdd1.t745 8.131
R13918 vdd1.n43 vdd1.t1394 8.131
R13919 vdd1.n42 vdd1.t451 8.131
R13920 vdd1.n41 vdd1.t860 8.131
R13921 vdd1.n40 vdd1.t1437 8.131
R13922 vdd1.n39 vdd1.t147 8.131
R13923 vdd1.n38 vdd1.t270 8.131
R13924 vdd1.n499 vdd1.t627 8.126
R13925 vdd1.n498 vdd1.t750 8.126
R13926 vdd1.n497 vdd1.t1322 8.126
R13927 vdd1.n496 vdd1.t457 8.126
R13928 vdd1.n495 vdd1.t1021 8.126
R13929 vdd1.n491 vdd1.t826 8.126
R13930 vdd1.n492 vdd1.t705 8.126
R13931 vdd1.n493 vdd1.t506 8.126
R13932 vdd1.n494 vdd1.t1445 8.126
R13933 vdd1.n933 vdd1.t1121 8.126
R13934 vdd1.n933 vdd1.t1335 8.126
R13935 vdd1.n934 vdd1.t563 8.126
R13936 vdd1.n934 vdd1.t759 8.126
R13937 vdd1.n935 vdd1.t434 8.126
R13938 vdd1.n935 vdd1.t639 8.126
R13939 vdd1.n936 vdd1.t225 8.126
R13940 vdd1.n936 vdd1.t422 8.126
R13941 vdd1.n937 vdd1.t1156 8.126
R13942 vdd1.n937 vdd1.t1368 8.126
R13943 vdd1.n938 vdd1.t743 8.126
R13944 vdd1.n938 vdd1.t950 8.126
R13945 vdd1.n939 vdd1.t188 8.126
R13946 vdd1.n939 vdd1.t388 8.126
R13947 vdd1.n940 vdd1.t1042 8.126
R13948 vdd1.n940 vdd1.t1254 8.126
R13949 vdd1.n941 vdd1.t475 8.126
R13950 vdd1.n941 vdd1.t674 8.126
R13951 vdd1.n942 vdd1.t361 8.126
R13952 vdd1.n942 vdd1.t564 8.126
R13953 vdd1.n921 vdd1.t709 8.126
R13954 vdd1.n921 vdd1.t919 8.126
R13955 vdd1.n922 vdd1.t156 8.126
R13956 vdd1.n922 vdd1.t360 8.126
R13957 vdd1.n923 vdd1.t31 8.126
R13958 vdd1.n923 vdd1.t234 8.126
R13959 vdd1.n924 vdd1.t1320 8.126
R13960 vdd1.n924 vdd1.t26 8.126
R13961 vdd1.n925 vdd1.t747 8.126
R13962 vdd1.n925 vdd1.t952 8.126
R13963 vdd1.n926 vdd1.t341 8.126
R13964 vdd1.n926 vdd1.t546 8.126
R13965 vdd1.n927 vdd1.t1278 8.126
R13966 vdd1.n927 vdd1.t1490 8.126
R13967 vdd1.n928 vdd1.t632 8.126
R13968 vdd1.n928 vdd1.t835 8.126
R13969 vdd1.n929 vdd1.t75 8.126
R13970 vdd1.n929 vdd1.t276 8.126
R13971 vdd1.n930 vdd1.t1456 8.126
R13972 vdd1.n930 vdd1.t157 8.126
R13973 vdd1.n905 vdd1.t948 8.126
R13974 vdd1.n905 vdd1.t511 8.126
R13975 vdd1.n906 vdd1.t386 8.126
R13976 vdd1.n906 vdd1.t1455 8.126
R13977 vdd1.n907 vdd1.t264 8.126
R13978 vdd1.n907 vdd1.t1325 8.126
R13979 vdd1.n908 vdd1.t55 8.126
R13980 vdd1.n908 vdd1.t1108 8.126
R13981 vdd1.n909 vdd1.t983 8.126
R13982 vdd1.n909 vdd1.t550 8.126
R13983 vdd1.n910 vdd1.t575 8.126
R13984 vdd1.n910 vdd1.t140 8.126
R13985 vdd1.n911 vdd1.t20 8.126
R13986 vdd1.n911 vdd1.t1066 8.126
R13987 vdd1.n912 vdd1.t869 8.126
R13988 vdd1.n912 vdd1.t424 8.126
R13989 vdd1.n913 vdd1.t302 8.126
R13990 vdd1.n913 vdd1.t1369 8.126
R13991 vdd1.n914 vdd1.t185 8.126
R13992 vdd1.n914 vdd1.t1244 8.126
R13993 vdd1.n893 vdd1.t543 8.126
R13994 vdd1.n893 vdd1.t739 8.126
R13995 vdd1.n894 vdd1.t1485 8.126
R13996 vdd1.n894 vdd1.t183 8.126
R13997 vdd1.n895 vdd1.t1354 8.126
R13998 vdd1.n895 vdd1.t61 8.126
R13999 vdd1.n896 vdd1.t1139 8.126
R14000 vdd1.n896 vdd1.t1348 8.126
R14001 vdd1.n897 vdd1.t579 8.126
R14002 vdd1.n897 vdd1.t778 8.126
R14003 vdd1.n898 vdd1.t168 8.126
R14004 vdd1.n898 vdd1.t370 8.126
R14005 vdd1.n899 vdd1.t1097 8.126
R14006 vdd1.n899 vdd1.t1311 8.126
R14007 vdd1.n900 vdd1.t462 8.126
R14008 vdd1.n900 vdd1.t665 8.126
R14009 vdd1.n901 vdd1.t1399 8.126
R14010 vdd1.n901 vdd1.t103 8.126
R14011 vdd1.n902 vdd1.t1274 8.126
R14012 vdd1.n902 vdd1.t1486 8.126
R14013 vdd1.n877 vdd1.t611 8.126
R14014 vdd1.n877 vdd1.t172 8.126
R14015 vdd1.n878 vdd1.t46 8.126
R14016 vdd1.n878 vdd1.t1102 8.126
R14017 vdd1.n879 vdd1.t1428 8.126
R14018 vdd1.n879 vdd1.t977 8.126
R14019 vdd1.n880 vdd1.t1207 8.126
R14020 vdd1.n880 vdd1.t764 8.126
R14021 vdd1.n881 vdd1.t643 8.126
R14022 vdd1.n881 vdd1.t215 8.126
R14023 vdd1.n882 vdd1.t239 8.126
R14024 vdd1.n882 vdd1.t1299 8.126
R14025 vdd1.n883 vdd1.t1164 8.126
R14026 vdd1.n883 vdd1.t728 8.126
R14027 vdd1.n884 vdd1.t536 8.126
R14028 vdd1.n884 vdd1.t95 8.126
R14029 vdd1.n885 vdd1.t1467 8.126
R14030 vdd1.n885 vdd1.t1015 8.126
R14031 vdd1.n886 vdd1.t1344 8.126
R14032 vdd1.n886 vdd1.t901 8.126
R14033 vdd1.n865 vdd1.t208 8.126
R14034 vdd1.n865 vdd1.t406 8.126
R14035 vdd1.n866 vdd1.t1133 8.126
R14036 vdd1.n866 vdd1.t1343 8.126
R14037 vdd1.n867 vdd1.t1005 8.126
R14038 vdd1.n867 vdd1.t1217 8.126
R14039 vdd1.n868 vdd1.t791 8.126
R14040 vdd1.n868 vdd1.t996 8.126
R14041 vdd1.n869 vdd1.t241 8.126
R14042 vdd1.n869 vdd1.t438 8.126
R14043 vdd1.n870 vdd1.t1329 8.126
R14044 vdd1.n870 vdd1.t34 8.126
R14045 vdd1.n871 vdd1.t756 8.126
R14046 vdd1.n871 vdd1.t959 8.126
R14047 vdd1.n872 vdd1.t128 8.126
R14048 vdd1.n872 vdd1.t330 8.126
R14049 vdd1.n873 vdd1.t1049 8.126
R14050 vdd1.n873 vdd1.t1257 8.126
R14051 vdd1.n874 vdd1.t933 8.126
R14052 vdd1.n874 vdd1.t1134 8.126
R14053 vdd1.n849 vdd1.t1294 8.126
R14054 vdd1.n849 vdd1.t8 8.126
R14055 vdd1.n850 vdd1.t721 8.126
R14056 vdd1.n850 vdd1.t932 8.126
R14057 vdd1.n851 vdd1.t598 8.126
R14058 vdd1.n851 vdd1.t796 8.126
R14059 vdd1.n852 vdd1.t391 8.126
R14060 vdd1.n852 vdd1.t593 8.126
R14061 vdd1.n853 vdd1.t1334 8.126
R14062 vdd1.n853 vdd1.t38 8.126
R14063 vdd1.n854 vdd1.t915 8.126
R14064 vdd1.n854 vdd1.t1115 8.126
R14065 vdd1.n855 vdd1.t356 8.126
R14066 vdd1.n855 vdd1.t559 8.126
R14067 vdd1.n856 vdd1.t1211 8.126
R14068 vdd1.n856 vdd1.t1421 8.126
R14069 vdd1.n857 vdd1.t644 8.126
R14070 vdd1.n857 vdd1.t843 8.126
R14071 vdd1.n858 vdd1.t525 8.126
R14072 vdd1.n858 vdd1.t722 8.126
R14073 vdd1.n837 vdd1.t33 8.126
R14074 vdd1.n837 vdd1.t238 8.126
R14075 vdd1.n838 vdd1.t957 8.126
R14076 vdd1.n838 vdd1.t1163 8.126
R14077 vdd1.n839 vdd1.t832 8.126
R14078 vdd1.n839 vdd1.t1038 8.126
R14079 vdd1.n840 vdd1.t626 8.126
R14080 vdd1.n840 vdd1.t825 8.126
R14081 vdd1.n841 vdd1.t72 8.126
R14082 vdd1.n841 vdd1.t274 8.126
R14083 vdd1.n842 vdd1.t1148 8.126
R14084 vdd1.n842 vdd1.t1363 8.126
R14085 vdd1.n843 vdd1.t588 8.126
R14086 vdd1.n843 vdd1.t784 8.126
R14087 vdd1.n844 vdd1.t1459 8.126
R14088 vdd1.n844 vdd1.t159 8.126
R14089 vdd1.n845 vdd1.t874 8.126
R14090 vdd1.n845 vdd1.t1076 8.126
R14091 vdd1.n846 vdd1.t754 8.126
R14092 vdd1.n846 vdd1.t958 8.126
R14093 vdd1.n821 vdd1.t1112 8.126
R14094 vdd1.n821 vdd1.t1327 8.126
R14095 vdd1.n822 vdd1.t556 8.126
R14096 vdd1.n822 vdd1.t753 8.126
R14097 vdd1.n823 vdd1.t423 8.126
R14098 vdd1.n823 vdd1.t631 8.126
R14099 vdd1.n824 vdd1.t223 8.126
R14100 vdd1.n824 vdd1.t420 8.126
R14101 vdd1.n825 vdd1.t1154 8.126
R14102 vdd1.n825 vdd1.t1365 8.126
R14103 vdd1.n826 vdd1.t736 8.126
R14104 vdd1.n826 vdd1.t944 8.126
R14105 vdd1.n827 vdd1.t181 8.126
R14106 vdd1.n827 vdd1.t384 8.126
R14107 vdd1.n828 vdd1.t1032 8.126
R14108 vdd1.n828 vdd1.t1245 8.126
R14109 vdd1.n829 vdd1.t473 8.126
R14110 vdd1.n829 vdd1.t673 8.126
R14111 vdd1.n830 vdd1.t353 8.126
R14112 vdd1.n830 vdd1.t557 8.126
R14113 vdd1.n809 vdd1.t1191 8.126
R14114 vdd1.n809 vdd1.t740 8.126
R14115 vdd1.n810 vdd1.t617 8.126
R14116 vdd1.n810 vdd1.t184 8.126
R14117 vdd1.n811 vdd1.t499 8.126
R14118 vdd1.n811 vdd1.t62 8.126
R14119 vdd1.n812 vdd1.t288 8.126
R14120 vdd1.n812 vdd1.t1349 8.126
R14121 vdd1.n813 vdd1.t1222 8.126
R14122 vdd1.n813 vdd1.t779 8.126
R14123 vdd1.n814 vdd1.t805 8.126
R14124 vdd1.n814 vdd1.t371 8.126
R14125 vdd1.n815 vdd1.t247 8.126
R14126 vdd1.n815 vdd1.t1312 8.126
R14127 vdd1.n816 vdd1.t1105 8.126
R14128 vdd1.n816 vdd1.t666 8.126
R14129 vdd1.n817 vdd1.t538 8.126
R14130 vdd1.n817 vdd1.t104 8.126
R14131 vdd1.n818 vdd1.t413 8.126
R14132 vdd1.n818 vdd1.t1487 8.126
R14133 vdd1.n793 vdd1.t773 8.126
R14134 vdd1.n793 vdd1.t980 8.126
R14135 vdd1.n794 vdd1.t218 8.126
R14136 vdd1.n794 vdd1.t412 8.126
R14137 vdd1.n795 vdd1.t91 8.126
R14138 vdd1.n795 vdd1.t294 8.126
R14139 vdd1.n796 vdd1.t1381 8.126
R14140 vdd1.n796 vdd1.t87 8.126
R14141 vdd1.n797 vdd1.t808 8.126
R14142 vdd1.n797 vdd1.t1012 8.126
R14143 vdd1.n798 vdd1.t399 8.126
R14144 vdd1.n798 vdd1.t605 8.126
R14145 vdd1.n799 vdd1.t1340 8.126
R14146 vdd1.n799 vdd1.t43 8.126
R14147 vdd1.n800 vdd1.t694 8.126
R14148 vdd1.n800 vdd1.t904 8.126
R14149 vdd1.n801 vdd1.t134 8.126
R14150 vdd1.n801 vdd1.t334 8.126
R14151 vdd1.n802 vdd1.t19 8.126
R14152 vdd1.n802 vdd1.t219 8.126
R14153 vdd1.n781 vdd1.t367 8.126
R14154 vdd1.n781 vdd1.t574 8.126
R14155 vdd1.n782 vdd1.t1307 8.126
R14156 vdd1.n782 vdd1.t18 8.126
R14157 vdd1.n783 vdd1.t1175 8.126
R14158 vdd1.n783 vdd1.t1383 8.126
R14159 vdd1.n784 vdd1.t964 8.126
R14160 vdd1.n784 vdd1.t1172 8.126
R14161 vdd1.n785 vdd1.t403 8.126
R14162 vdd1.n785 vdd1.t609 8.126
R14163 vdd1.n786 vdd1.t4 8.126
R14164 vdd1.n786 vdd1.t204 8.126
R14165 vdd1.n787 vdd1.t929 8.126
R14166 vdd1.n787 vdd1.t1130 8.126
R14167 vdd1.n788 vdd1.t289 8.126
R14168 vdd1.n788 vdd1.t495 8.126
R14169 vdd1.n789 vdd1.t1223 8.126
R14170 vdd1.n789 vdd1.t1432 8.126
R14171 vdd1.n790 vdd1.t1094 8.126
R14172 vdd1.n790 vdd1.t1308 8.126
R14173 vdd1.n765 vdd1.t601 8.126
R14174 vdd1.n765 vdd1.t801 8.126
R14175 vdd1.n766 vdd1.t41 8.126
R14176 vdd1.n766 vdd1.t244 8.126
R14177 vdd1.n767 vdd1.t1420 8.126
R14178 vdd1.n767 vdd1.t125 8.126
R14179 vdd1.n768 vdd1.t1205 8.126
R14180 vdd1.n768 vdd1.t1415 8.126
R14181 vdd1.n769 vdd1.t642 8.126
R14182 vdd1.n769 vdd1.t842 8.126
R14183 vdd1.n770 vdd1.t231 8.126
R14184 vdd1.n770 vdd1.t430 8.126
R14185 vdd1.n771 vdd1.t1159 8.126
R14186 vdd1.n771 vdd1.t1370 8.126
R14187 vdd1.n772 vdd1.t529 8.126
R14188 vdd1.n772 vdd1.t725 8.126
R14189 vdd1.n773 vdd1.t1466 8.126
R14190 vdd1.n773 vdd1.t163 8.126
R14191 vdd1.n774 vdd1.t1338 8.126
R14192 vdd1.n774 vdd1.t42 8.126
R14193 vdd1.n753 vdd1.t199 8.126
R14194 vdd1.n753 vdd1.t395 8.126
R14195 vdd1.n754 vdd1.t1127 8.126
R14196 vdd1.n754 vdd1.t1337 8.126
R14197 vdd1.n755 vdd1.t997 8.126
R14198 vdd1.n755 vdd1.t1208 8.126
R14199 vdd1.n756 vdd1.t790 8.126
R14200 vdd1.n756 vdd1.t995 8.126
R14201 vdd1.n757 vdd1.t236 8.126
R14202 vdd1.n757 vdd1.t436 8.126
R14203 vdd1.n758 vdd1.t1324 8.126
R14204 vdd1.n758 vdd1.t30 8.126
R14205 vdd1.n759 vdd1.t751 8.126
R14206 vdd1.n759 vdd1.t955 8.126
R14207 vdd1.n760 vdd1.t121 8.126
R14208 vdd1.n760 vdd1.t321 8.126
R14209 vdd1.n761 vdd1.t1048 8.126
R14210 vdd1.n761 vdd1.t1256 8.126
R14211 vdd1.n762 vdd1.t926 8.126
R14212 vdd1.n762 vdd1.t1128 8.126
R14213 vdd1.n737 vdd1.t271 8.126
R14214 vdd1.n737 vdd1.t470 8.126
R14215 vdd1.n738 vdd1.t1196 8.126
R14216 vdd1.n738 vdd1.t1403 8.126
R14217 vdd1.n739 vdd1.t1070 8.126
R14218 vdd1.n739 vdd1.t1287 8.126
R14219 vdd1.n740 vdd1.t858 8.126
R14220 vdd1.n740 vdd1.t1062 8.126
R14221 vdd1.n741 vdd1.t300 8.126
R14222 vdd1.n741 vdd1.t504 8.126
R14223 vdd1.n742 vdd1.t1395 8.126
R14224 vdd1.n742 vdd1.t100 8.126
R14225 vdd1.n743 vdd1.t812 8.126
R14226 vdd1.n743 vdd1.t1017 8.126
R14227 vdd1.n744 vdd1.t190 8.126
R14228 vdd1.n744 vdd1.t387 8.126
R14229 vdd1.n745 vdd1.t1107 8.126
R14230 vdd1.n745 vdd1.t1319 8.126
R14231 vdd1.n746 vdd1.t986 8.126
R14232 vdd1.n746 vdd1.t1197 8.126
R14233 vdd1.n725 vdd1.t1357 8.126
R14234 vdd1.n725 vdd1.t65 8.126
R14235 vdd1.n726 vdd1.t781 8.126
R14236 vdd1.n726 vdd1.t985 8.126
R14237 vdd1.n727 vdd1.t662 8.126
R14238 vdd1.n727 vdd1.t867 8.126
R14239 vdd1.n728 vdd1.t454 8.126
R14240 vdd1.n728 vdd1.t657 8.126
R14241 vdd1.n729 vdd1.t1397 8.126
R14242 vdd1.n729 vdd1.t102 8.126
R14243 vdd1.n730 vdd1.t973 8.126
R14244 vdd1.n730 vdd1.t1181 8.126
R14245 vdd1.n731 vdd1.t410 8.126
R14246 vdd1.n731 vdd1.t614 8.126
R14247 vdd1.n732 vdd1.t1277 8.126
R14248 vdd1.n732 vdd1.t1492 8.126
R14249 vdd1.n733 vdd1.t701 8.126
R14250 vdd1.n733 vdd1.t908 8.126
R14251 vdd1.n734 vdd1.t586 8.126
R14252 vdd1.n734 vdd1.t782 8.126
R14253 vdd1.n709 vdd1.t1379 8.126
R14254 vdd1.n709 vdd1.t1144 8.126
R14255 vdd1.n710 vdd1.t800 8.126
R14256 vdd1.n710 vdd1.t585 8.126
R14257 vdd1.n711 vdd1.t681 8.126
R14258 vdd1.n711 vdd1.t458 8.126
R14259 vdd1.n712 vdd1.t477 8.126
R14260 vdd1.n712 vdd1.t257 8.126
R14261 vdd1.n713 vdd1.t1414 8.126
R14262 vdd1.n713 vdd1.t1190 8.126
R14263 vdd1.n714 vdd1.t992 8.126
R14264 vdd1.n714 vdd1.t770 8.126
R14265 vdd1.n715 vdd1.t429 8.126
R14266 vdd1.n715 vdd1.t217 8.126
R14267 vdd1.n716 vdd1.t1297 8.126
R14268 vdd1.n716 vdd1.t1065 8.126
R14269 vdd1.n717 vdd1.t724 8.126
R14270 vdd1.n717 vdd1.t505 8.126
R14271 vdd1.n718 vdd1.t602 8.126
R14272 vdd1.n718 vdd1.t382 8.126
R14273 vdd1.n697 vdd1.t963 8.126
R14274 vdd1.n697 vdd1.t1169 8.126
R14275 vdd1.n698 vdd1.t394 8.126
R14276 vdd1.n698 vdd1.t600 8.126
R14277 vdd1.n699 vdd1.t279 8.126
R14278 vdd1.n699 vdd1.t481 8.126
R14279 vdd1.n700 vdd1.t77 8.126
R14280 vdd1.n700 vdd1.t277 8.126
R14281 vdd1.n701 vdd1.t994 8.126
R14282 vdd1.n701 vdd1.t1204 8.126
R14283 vdd1.n702 vdd1.t591 8.126
R14284 vdd1.n702 vdd1.t787 8.126
R14285 vdd1.n703 vdd1.t29 8.126
R14286 vdd1.n703 vdd1.t230 8.126
R14287 vdd1.n704 vdd1.t882 8.126
R14288 vdd1.n704 vdd1.t1084 8.126
R14289 vdd1.n705 vdd1.t320 8.126
R14290 vdd1.n705 vdd1.t528 8.126
R14291 vdd1.n706 vdd1.t200 8.126
R14292 vdd1.n706 vdd1.t396 8.126
R14293 vdd1.n681 vdd1.t566 8.126
R14294 vdd1.n681 vdd1.t761 8.126
R14295 vdd1.n682 vdd1.t0 8.126
R14296 vdd1.n682 vdd1.t198 8.126
R14297 vdd1.n683 vdd1.t1374 8.126
R14298 vdd1.n683 vdd1.t78 8.126
R14299 vdd1.n684 vdd1.t1162 8.126
R14300 vdd1.n684 vdd1.t1373 8.126
R14301 vdd1.n685 vdd1.t592 8.126
R14302 vdd1.n685 vdd1.t789 8.126
R14303 vdd1.n686 vdd1.t193 8.126
R14304 vdd1.n686 vdd1.t390 8.126
R14305 vdd1.n687 vdd1.t1110 8.126
R14306 vdd1.n687 vdd1.t1323 8.126
R14307 vdd1.n688 vdd1.t479 8.126
R14308 vdd1.n688 vdd1.t679 8.126
R14309 vdd1.n689 vdd1.t1417 8.126
R14310 vdd1.n689 vdd1.t120 8.126
R14311 vdd1.n690 vdd1.t1289 8.126
R14312 vdd1.n690 vdd1.t1 8.126
R14313 vdd1.n669 vdd1.t623 8.126
R14314 vdd1.n669 vdd1.t822 8.126
R14315 vdd1.n670 vdd1.t64 8.126
R14316 vdd1.n670 vdd1.t268 8.126
R14317 vdd1.n671 vdd1.t1443 8.126
R14318 vdd1.n671 vdd1.t144 8.126
R14319 vdd1.n672 vdd1.t1227 8.126
R14320 vdd1.n672 vdd1.t1436 8.126
R14321 vdd1.n673 vdd1.t656 8.126
R14322 vdd1.n673 vdd1.t857 8.126
R14323 vdd1.n674 vdd1.t253 8.126
R14324 vdd1.n674 vdd1.t449 8.126
R14325 vdd1.n675 vdd1.t1180 8.126
R14326 vdd1.n675 vdd1.t1390 8.126
R14327 vdd1.n676 vdd1.t545 8.126
R14328 vdd1.n676 vdd1.t742 8.126
R14329 vdd1.n677 vdd1.t1489 8.126
R14330 vdd1.n677 vdd1.t187 8.126
R14331 vdd1.n678 vdd1.t1358 8.126
R14332 vdd1.n678 vdd1.t66 8.126
R14333 vdd1.n653 vdd1.t222 8.126
R14334 vdd1.n653 vdd1.t417 8.126
R14335 vdd1.n654 vdd1.t1143 8.126
R14336 vdd1.n654 vdd1.t1356 8.126
R14337 vdd1.n655 vdd1.t1022 8.126
R14338 vdd1.n655 vdd1.t1232 8.126
R14339 vdd1.n656 vdd1.t814 8.126
R14340 vdd1.n656 vdd1.t1018 8.126
R14341 vdd1.n657 vdd1.t256 8.126
R14342 vdd1.n657 vdd1.t453 8.126
R14343 vdd1.n658 vdd1.t1347 8.126
R14344 vdd1.n658 vdd1.t50 8.126
R14345 vdd1.n659 vdd1.t769 8.126
R14346 vdd1.n659 vdd1.t972 8.126
R14347 vdd1.n660 vdd1.t139 8.126
R14348 vdd1.n660 vdd1.t340 8.126
R14349 vdd1.n661 vdd1.t1064 8.126
R14350 vdd1.n661 vdd1.t1276 8.126
R14351 vdd1.n662 vdd1.t942 8.126
R14352 vdd1.n662 vdd1.t1145 8.126
R14353 vdd1.n641 vdd1.t447 8.126
R14354 vdd1.n641 vdd1.t24 8.126
R14355 vdd1.n642 vdd1.t1387 8.126
R14356 vdd1.n642 vdd1.t941 8.126
R14357 vdd1.n643 vdd1.t1262 8.126
R14358 vdd1.n643 vdd1.t815 8.126
R14359 vdd1.n644 vdd1.t1050 8.126
R14360 vdd1.n644 vdd1.t618 8.126
R14361 vdd1.n645 vdd1.t487 8.126
R14362 vdd1.n645 vdd1.t53 8.126
R14363 vdd1.n646 vdd1.t81 8.126
R14364 vdd1.n646 vdd1.t1138 8.126
R14365 vdd1.n647 vdd1.t1003 8.126
R14366 vdd1.n647 vdd1.t572 8.126
R14367 vdd1.n648 vdd1.t369 8.126
R14368 vdd1.n648 vdd1.t1440 8.126
R14369 vdd1.n649 vdd1.t1310 8.126
R14370 vdd1.n649 vdd1.t862 8.126
R14371 vdd1.n650 vdd1.t1178 8.126
R14372 vdd1.n650 vdd1.t733 8.126
R14373 vdd1.n625 vdd1.t48 8.126
R14374 vdd1.n625 vdd1.t251 8.126
R14375 vdd1.n626 vdd1.t968 8.126
R14376 vdd1.n626 vdd1.t1177 8.126
R14377 vdd1.n627 vdd1.t847 8.126
R14378 vdd1.n627 vdd1.t1054 8.126
R14379 vdd1.n628 vdd1.t646 8.126
R14380 vdd1.n628 vdd1.t845 8.126
R14381 vdd1.n629 vdd1.t83 8.126
R14382 vdd1.n629 vdd1.t284 8.126
R14383 vdd1.n630 vdd1.t1166 8.126
R14384 vdd1.n630 vdd1.t1376 8.126
R14385 vdd1.n631 vdd1.t595 8.126
R14386 vdd1.n631 vdd1.t795 8.126
R14387 vdd1.n632 vdd1.t1470 8.126
R14388 vdd1.n632 vdd1.t167 8.126
R14389 vdd1.n633 vdd1.t894 8.126
R14390 vdd1.n633 vdd1.t1096 8.126
R14391 vdd1.n634 vdd1.t766 8.126
R14392 vdd1.n634 vdd1.t969 8.126
R14393 vdd1.n613 vdd1.t1137 8.126
R14394 vdd1.n613 vdd1.t1346 8.126
R14395 vdd1.n614 vdd1.t569 8.126
R14396 vdd1.n614 vdd1.t765 8.126
R14397 vdd1.n615 vdd1.t443 8.126
R14398 vdd1.n615 vdd1.t648 8.126
R14399 vdd1.n616 vdd1.t246 8.126
R14400 vdd1.n616 vdd1.t442 8.126
R14401 vdd1.n617 vdd1.t1168 8.126
R14402 vdd1.n617 vdd1.t1377 8.126
R14403 vdd1.n618 vdd1.t760 8.126
R14404 vdd1.n618 vdd1.t962 8.126
R14405 vdd1.n619 vdd1.t194 8.126
R14406 vdd1.n619 vdd1.t392 8.126
R14407 vdd1.n620 vdd1.t1053 8.126
R14408 vdd1.n620 vdd1.t1259 8.126
R14409 vdd1.n621 vdd1.t491 8.126
R14410 vdd1.n621 vdd1.t688 8.126
R14411 vdd1.n622 vdd1.t364 8.126
R14412 vdd1.n622 vdd1.t570 8.126
R14413 vdd1.n597 vdd1.t1200 8.126
R14414 vdd1.n597 vdd1.t1410 8.126
R14415 vdd1.n598 vdd1.t633 8.126
R14416 vdd1.n598 vdd1.t836 8.126
R14417 vdd1.n599 vdd1.t512 8.126
R14418 vdd1.n599 vdd1.t710 8.126
R14419 vdd1.n600 vdd1.t303 8.126
R14420 vdd1.n600 vdd1.t508 8.126
R14421 vdd1.n601 vdd1.t1240 8.126
R14422 vdd1.n601 vdd1.t1452 8.126
R14423 vdd1.n602 vdd1.t818 8.126
R14424 vdd1.n602 vdd1.t1026 8.126
R14425 vdd1.n603 vdd1.t262 8.126
R14426 vdd1.n603 vdd1.t465 8.126
R14427 vdd1.n604 vdd1.t1114 8.126
R14428 vdd1.n604 vdd1.t1328 8.126
R14429 vdd1.n605 vdd1.t558 8.126
R14430 vdd1.n605 vdd1.t755 8.126
R14431 vdd1.n606 vdd1.t426 8.126
R14432 vdd1.n606 vdd1.t634 8.126
R14433 vdd1.n585 vdd1.t786 8.126
R14434 vdd1.n585 vdd1.t990 8.126
R14435 vdd1.n586 vdd1.t226 8.126
R14436 vdd1.n586 vdd1.t425 8.126
R14437 vdd1.n587 vdd1.t108 8.126
R14438 vdd1.n587 vdd1.t307 8.126
R14439 vdd1.n588 vdd1.t1402 8.126
R14440 vdd1.n588 vdd1.t106 8.126
R14441 vdd1.n589 vdd1.t820 8.126
R14442 vdd1.n589 vdd1.t1028 8.126
R14443 vdd1.n590 vdd1.t416 8.126
R14444 vdd1.n590 vdd1.t621 8.126
R14445 vdd1.n591 vdd1.t1352 8.126
R14446 vdd1.n591 vdd1.t59 8.126
R14447 vdd1.n592 vdd1.t707 8.126
R14448 vdd1.n592 vdd1.t914 8.126
R14449 vdd1.n593 vdd1.t154 8.126
R14450 vdd1.n593 vdd1.t355 8.126
R14451 vdd1.n594 vdd1.t27 8.126
R14452 vdd1.n594 vdd1.t227 8.126
R14453 vdd1.n569 vdd1.t1024 8.126
R14454 vdd1.n569 vdd1.t1235 8.126
R14455 vdd1.n570 vdd1.t460 8.126
R14456 vdd1.n570 vdd1.t664 8.126
R14457 vdd1.n571 vdd1.t338 8.126
R14458 vdd1.n571 vdd1.t542 8.126
R14459 vdd1.n572 vdd1.t135 8.126
R14460 vdd1.n572 vdd1.t335 8.126
R14461 vdd1.n573 vdd1.t1058 8.126
R14462 vdd1.n573 vdd1.t1269 8.126
R14463 vdd1.n574 vdd1.t650 8.126
R14464 vdd1.n574 vdd1.t850 8.126
R14465 vdd1.n575 vdd1.t90 8.126
R14466 vdd1.n575 vdd1.t291 8.126
R14467 vdd1.n576 vdd1.t943 8.126
R14468 vdd1.n576 vdd1.t1147 8.126
R14469 vdd1.n577 vdd1.t383 8.126
R14470 vdd1.n577 vdd1.t587 8.126
R14471 vdd1.n578 vdd1.t259 8.126
R14472 vdd1.n578 vdd1.t461 8.126
R14473 vdd1.n557 vdd1.t620 8.126
R14474 vdd1.n557 vdd1.t816 8.126
R14475 vdd1.n558 vdd1.t56 8.126
R14476 vdd1.n558 vdd1.t258 8.126
R14477 vdd1.n559 vdd1.t1438 8.126
R14478 vdd1.n559 vdd1.t137 8.126
R14479 vdd1.n560 vdd1.t1226 8.126
R14480 vdd1.n560 vdd1.t1434 8.126
R14481 vdd1.n561 vdd1.t652 8.126
R14482 vdd1.n561 vdd1.t852 8.126
R14483 vdd1.n562 vdd1.t250 8.126
R14484 vdd1.n562 vdd1.t444 8.126
R14485 vdd1.n563 vdd1.t1174 8.126
R14486 vdd1.n563 vdd1.t1382 8.126
R14487 vdd1.n564 vdd1.t541 8.126
R14488 vdd1.n564 vdd1.t735 8.126
R14489 vdd1.n565 vdd1.t1484 8.126
R14490 vdd1.n565 vdd1.t180 8.126
R14491 vdd1.n566 vdd1.t1351 8.126
R14492 vdd1.n566 vdd1.t57 8.126
R14493 vdd1.n541 vdd1.t849 8.126
R14494 vdd1.n541 vdd1.t415 8.126
R14495 vdd1.n542 vdd1.t290 8.126
R14496 vdd1.n542 vdd1.t1350 8.126
R14497 vdd1.n543 vdd1.t166 8.126
R14498 vdd1.n543 vdd1.t1229 8.126
R14499 vdd1.n544 vdd1.t1468 8.126
R14500 vdd1.n544 vdd1.t1016 8.126
R14501 vdd1.n545 vdd1.t888 8.126
R14502 vdd1.n545 vdd1.t446 8.126
R14503 vdd1.n546 vdd1.t480 8.126
R14504 vdd1.n546 vdd1.t47 8.126
R14505 vdd1.n547 vdd1.t1419 8.126
R14506 vdd1.n547 vdd1.t966 8.126
R14507 vdd1.n548 vdd1.t768 8.126
R14508 vdd1.n548 vdd1.t337 8.126
R14509 vdd1.n549 vdd1.t216 8.126
R14510 vdd1.n549 vdd1.t1273 8.126
R14511 vdd1.n550 vdd1.t89 8.126
R14512 vdd1.n550 vdd1.t1140 8.126
R14513 vdd1.n529 vdd1.t280 8.126
R14514 vdd1.n529 vdd1.t483 8.126
R14515 vdd1.n530 vdd1.t1209 8.126
R14516 vdd1.n530 vdd1.t1422 8.126
R14517 vdd1.n531 vdd1.t1081 8.126
R14518 vdd1.n531 vdd1.t1293 8.126
R14519 vdd1.n532 vdd1.t875 8.126
R14520 vdd1.n532 vdd1.t1077 8.126
R14521 vdd1.n533 vdd1.t313 8.126
R14522 vdd1.n533 vdd1.t521 8.126
R14523 vdd1.n534 vdd1.t1405 8.126
R14524 vdd1.n534 vdd1.t111 8.126
R14525 vdd1.n535 vdd1.t828 8.126
R14526 vdd1.n535 vdd1.t1037 8.126
R14527 vdd1.n536 vdd1.t203 8.126
R14528 vdd1.n536 vdd1.t398 8.126
R14529 vdd1.n537 vdd1.t1129 8.126
R14530 vdd1.n537 vdd1.t1339 8.126
R14531 vdd1.n538 vdd1.t999 8.126
R14532 vdd1.n538 vdd1.t1210 8.126
R14533 vdd1.n513 vdd1.t1375 8.126
R14534 vdd1.n513 vdd1.t79 8.126
R14535 vdd1.n514 vdd1.t792 8.126
R14536 vdd1.n514 vdd1.t998 8.126
R14537 vdd1.n515 vdd1.t678 8.126
R14538 vdd1.n515 vdd1.t879 8.126
R14539 vdd1.n516 vdd1.t476 8.126
R14540 vdd1.n516 vdd1.t675 8.126
R14541 vdd1.n517 vdd1.t1409 8.126
R14542 vdd1.n517 vdd1.t113 8.126
R14543 vdd1.n518 vdd1.t989 8.126
R14544 vdd1.n518 vdd1.t1198 8.126
R14545 vdd1.n519 vdd1.t421 8.126
R14546 vdd1.n519 vdd1.t628 8.126
R14547 vdd1.n520 vdd1.t1292 8.126
R14548 vdd1.n520 vdd1.t3 8.126
R14549 vdd1.n521 vdd1.t719 8.126
R14550 vdd1.n521 vdd1.t928 8.126
R14551 vdd1.n522 vdd1.t594 8.126
R14552 vdd1.n522 vdd1.t793 8.126
R14553 vdd1.n501 vdd1.t109 8.126
R14554 vdd1.n501 vdd1.t309 8.126
R14555 vdd1.n502 vdd1.t1033 8.126
R14556 vdd1.n502 vdd1.t1247 8.126
R14557 vdd1.n503 vdd1.t912 8.126
R14558 vdd1.n503 vdd1.t1113 8.126
R14559 vdd1.n504 vdd1.t702 8.126
R14560 vdd1.n504 vdd1.t909 8.126
R14561 vdd1.n505 vdd1.t146 8.126
R14562 vdd1.n505 vdd1.t349 8.126
R14563 vdd1.n506 vdd1.t1231 8.126
R14564 vdd1.n506 vdd1.t1441 8.126
R14565 vdd1.n507 vdd1.t660 8.126
R14566 vdd1.n507 vdd1.t863 8.126
R14567 vdd1.n508 vdd1.t28 8.126
R14568 vdd1.n508 vdd1.t229 8.126
R14569 vdd1.n509 vdd1.t954 8.126
R14570 vdd1.n509 vdd1.t1158 8.126
R14571 vdd1.n510 vdd1.t827 8.126
R14572 vdd1.n510 vdd1.t1034 8.126
R14573 vdd1.n47 vdd1.t418 8.126
R14574 vdd1.n47 vdd1.t624 8.126
R14575 vdd1.n48 vdd1.t1359 8.126
R14576 vdd1.n48 vdd1.t68 8.126
R14577 vdd1.n49 vdd1.t1234 8.126
R14578 vdd1.n49 vdd1.t1446 8.126
R14579 vdd1.n50 vdd1.t1019 8.126
R14580 vdd1.n50 vdd1.t1228 8.126
R14581 vdd1.n51 vdd1.t455 8.126
R14582 vdd1.n51 vdd1.t658 8.126
R14583 vdd1.n52 vdd1.t51 8.126
R14584 vdd1.n52 vdd1.t254 8.126
R14585 vdd1.n53 vdd1.t975 8.126
R14586 vdd1.n53 vdd1.t1185 8.126
R14587 vdd1.n54 vdd1.t343 8.126
R14588 vdd1.n54 vdd1.t548 8.126
R14589 vdd1.n55 vdd1.t1279 8.126
R14590 vdd1.n55 vdd1.t1491 8.126
R14591 vdd1.n56 vdd1.t1146 8.126
R14592 vdd1.n56 vdd1.t1360 8.126
R14593 vdd1.n58 vdd1.t492 8.126
R14594 vdd1.n58 vdd1.t54 8.126
R14595 vdd1.n59 vdd1.t1431 8.126
R14596 vdd1.n59 vdd1.t981 8.126
R14597 vdd1.n60 vdd1.t1304 8.126
R14598 vdd1.n60 vdd1.t853 8.126
R14599 vdd1.n61 vdd1.t1080 8.126
R14600 vdd1.n61 vdd1.t649 8.126
R14601 vdd1.n62 vdd1.t527 8.126
R14602 vdd1.n62 vdd1.t88 8.126
R14603 vdd1.n63 vdd1.t118 8.126
R14604 vdd1.n63 vdd1.t1171 8.126
R14605 vdd1.n64 vdd1.t1047 8.126
R14606 vdd1.n64 vdd1.t608 8.126
R14607 vdd1.n65 vdd1.t408 8.126
R14608 vdd1.n65 vdd1.t1480 8.126
R14609 vdd1.n66 vdd1.t1345 8.126
R14610 vdd1.n66 vdd1.t906 8.126
R14611 vdd1.n67 vdd1.t1221 8.126
R14612 vdd1.n67 vdd1.t774 8.126
R14613 vdd1.n69 vdd1.t86 8.126
R14614 vdd1.n69 vdd1.t287 8.126
R14615 vdd1.n70 vdd1.t1010 8.126
R14616 vdd1.n70 vdd1.t1220 8.126
R14617 vdd1.n71 vdd1.t889 8.126
R14618 vdd1.n71 vdd1.t1092 8.126
R14619 vdd1.n72 vdd1.t677 8.126
R14620 vdd1.n72 vdd1.t878 8.126
R14621 vdd1.n73 vdd1.t119 8.126
R14622 vdd1.n73 vdd1.t318 8.126
R14623 vdd1.n74 vdd1.t1203 8.126
R14624 vdd1.n74 vdd1.t1413 8.126
R14625 vdd1.n75 vdd1.t641 8.126
R14626 vdd1.n75 vdd1.t841 8.126
R14627 vdd1.n76 vdd1.t14 8.126
R14628 vdd1.n76 vdd1.t213 8.126
R14629 vdd1.n77 vdd1.t936 8.126
R14630 vdd1.n77 vdd1.t1136 8.126
R14631 vdd1.n78 vdd1.t804 8.126
R14632 vdd1.n78 vdd1.t1011 8.126
R14633 vdd1.n80 vdd1.t1170 8.126
R14634 vdd1.n80 vdd1.t1380 8.126
R14635 vdd1.n81 vdd1.t603 8.126
R14636 vdd1.n81 vdd1.t803 8.126
R14637 vdd1.n82 vdd1.t482 8.126
R14638 vdd1.n82 vdd1.t683 8.126
R14639 vdd1.n83 vdd1.t278 8.126
R14640 vdd1.n83 vdd1.t478 8.126
R14641 vdd1.n84 vdd1.t1206 8.126
R14642 vdd1.n84 vdd1.t1416 8.126
R14643 vdd1.n85 vdd1.t788 8.126
R14644 vdd1.n85 vdd1.t993 8.126
R14645 vdd1.n86 vdd1.t233 8.126
R14646 vdd1.n86 vdd1.t433 8.126
R14647 vdd1.n87 vdd1.t1087 8.126
R14648 vdd1.n87 vdd1.t1301 8.126
R14649 vdd1.n88 vdd1.t531 8.126
R14650 vdd1.n88 vdd1.t727 8.126
R14651 vdd1.n89 vdd1.t397 8.126
R14652 vdd1.n89 vdd1.t604 8.126
R14653 vdd1.n91 vdd1.t1411 8.126
R14654 vdd1.n91 vdd1.t116 8.126
R14655 vdd1.n92 vdd1.t837 8.126
R14656 vdd1.n92 vdd1.t1044 8.126
R14657 vdd1.n93 vdd1.t713 8.126
R14658 vdd1.n93 vdd1.t921 8.126
R14659 vdd1.n94 vdd1.t509 8.126
R14660 vdd1.n94 vdd1.t704 8.126
R14661 vdd1.n95 vdd1.t1453 8.126
R14662 vdd1.n95 vdd1.t152 8.126
R14663 vdd1.n96 vdd1.t1027 8.126
R14664 vdd1.n96 vdd1.t1238 8.126
R14665 vdd1.n97 vdd1.t466 8.126
R14666 vdd1.n97 vdd1.t669 8.126
R14667 vdd1.n98 vdd1.t1331 8.126
R14668 vdd1.n98 vdd1.t36 8.126
R14669 vdd1.n99 vdd1.t757 8.126
R14670 vdd1.n99 vdd1.t960 8.126
R14671 vdd1.n100 vdd1.t636 8.126
R14672 vdd1.n100 vdd1.t838 8.126
R14673 vdd1.n102 vdd1.t991 8.126
R14674 vdd1.n102 vdd1.t1201 8.126
R14675 vdd1.n103 vdd1.t427 8.126
R14676 vdd1.n103 vdd1.t635 8.126
R14677 vdd1.n104 vdd1.t306 8.126
R14678 vdd1.n104 vdd1.t515 8.126
R14679 vdd1.n105 vdd1.t107 8.126
R14680 vdd1.n105 vdd1.t304 8.126
R14681 vdd1.n106 vdd1.t1030 8.126
R14682 vdd1.n106 vdd1.t1241 8.126
R14683 vdd1.n107 vdd1.t622 8.126
R14684 vdd1.n107 vdd1.t819 8.126
R14685 vdd1.n108 vdd1.t60 8.126
R14686 vdd1.n108 vdd1.t263 8.126
R14687 vdd1.n109 vdd1.t917 8.126
R14688 vdd1.n109 vdd1.t1117 8.126
R14689 vdd1.n110 vdd1.t357 8.126
R14690 vdd1.n110 vdd1.t560 8.126
R14691 vdd1.n111 vdd1.t228 8.126
R14692 vdd1.n111 vdd1.t428 8.126
R14693 vdd1.n113 vdd1.t1061 8.126
R14694 vdd1.n113 vdd1.t1272 8.126
R14695 vdd1.n114 vdd1.t502 8.126
R14696 vdd1.n114 vdd1.t700 8.126
R14697 vdd1.n115 vdd1.t377 8.126
R14698 vdd1.n115 vdd1.t582 8.126
R14699 vdd1.n116 vdd1.t165 8.126
R14700 vdd1.n116 vdd1.t368 8.126
R14701 vdd1.n117 vdd1.t1095 8.126
R14702 vdd1.n117 vdd1.t1309 8.126
R14703 vdd1.n118 vdd1.t686 8.126
R14704 vdd1.n118 vdd1.t892 8.126
R14705 vdd1.n119 vdd1.t133 8.126
R14706 vdd1.n119 vdd1.t333 8.126
R14707 vdd1.n120 vdd1.t982 8.126
R14708 vdd1.n120 vdd1.t1192 8.126
R14709 vdd1.n121 vdd1.t414 8.126
R14710 vdd1.n121 vdd1.t619 8.126
R14711 vdd1.n122 vdd1.t298 8.126
R14712 vdd1.n122 vdd1.t503 8.126
R14713 vdd1.n124 vdd1.t653 8.126
R14714 vdd1.n124 vdd1.t855 8.126
R14715 vdd1.n125 vdd1.t96 8.126
R14716 vdd1.n125 vdd1.t297 8.126
R14717 vdd1.n126 vdd1.t1477 8.126
R14718 vdd1.n126 vdd1.t174 8.126
R14719 vdd1.n127 vdd1.t1258 8.126
R14720 vdd1.n127 vdd1.t1469 8.126
R14721 vdd1.n128 vdd1.t687 8.126
R14722 vdd1.n128 vdd1.t893 8.126
R14723 vdd1.n129 vdd1.t283 8.126
R14724 vdd1.n129 vdd1.t486 8.126
R14725 vdd1.n130 vdd1.t1216 8.126
R14726 vdd1.n130 vdd1.t1427 8.126
R14727 vdd1.n131 vdd1.t578 8.126
R14728 vdd1.n131 vdd1.t776 8.126
R14729 vdd1.n132 vdd1.t21 8.126
R14730 vdd1.n132 vdd1.t220 8.126
R14731 vdd1.n133 vdd1.t1389 8.126
R14732 vdd1.n133 vdd1.t97 8.126
R14733 vdd1.n135 vdd1.t890 8.126
R14734 vdd1.n135 vdd1.t448 8.126
R14735 vdd1.n136 vdd1.t331 8.126
R14736 vdd1.n136 vdd1.t1388 8.126
R14737 vdd1.n137 vdd1.t210 8.126
R14738 vdd1.n137 vdd1.t1264 8.126
R14739 vdd1.n138 vdd1.t2 8.126
R14740 vdd1.n138 vdd1.t1051 8.126
R14741 vdd1.n139 vdd1.t927 8.126
R14742 vdd1.n139 vdd1.t489 8.126
R14743 vdd1.n140 vdd1.t520 8.126
R14744 vdd1.n140 vdd1.t82 8.126
R14745 vdd1.n141 vdd1.t1464 8.126
R14746 vdd1.n141 vdd1.t1004 8.126
R14747 vdd1.n142 vdd1.t807 8.126
R14748 vdd1.n142 vdd1.t373 8.126
R14749 vdd1.n143 vdd1.t248 8.126
R14750 vdd1.n143 vdd1.t1313 8.126
R14751 vdd1.n144 vdd1.t130 8.126
R14752 vdd1.n144 vdd1.t1179 8.126
R14753 vdd1.n146 vdd1.t484 8.126
R14754 vdd1.n146 vdd1.t684 8.126
R14755 vdd1.n147 vdd1.t1423 8.126
R14756 vdd1.n147 vdd1.t129 8.126
R14757 vdd1.n148 vdd1.t1296 8.126
R14758 vdd1.n148 vdd1.t9 8.126
R14759 vdd1.n149 vdd1.t1078 8.126
R14760 vdd1.n149 vdd1.t1290 8.126
R14761 vdd1.n150 vdd1.t523 8.126
R14762 vdd1.n150 vdd1.t718 8.126
R14763 vdd1.n151 vdd1.t112 8.126
R14764 vdd1.n151 vdd1.t312 8.126
R14765 vdd1.n152 vdd1.t1041 8.126
R14766 vdd1.n152 vdd1.t1252 8.126
R14767 vdd1.n153 vdd1.t402 8.126
R14768 vdd1.n153 vdd1.t607 8.126
R14769 vdd1.n154 vdd1.t1341 8.126
R14770 vdd1.n154 vdd1.t44 8.126
R14771 vdd1.n155 vdd1.t1213 8.126
R14772 vdd1.n155 vdd1.t1424 8.126
R14773 vdd1.n157 vdd1.t80 8.126
R14774 vdd1.n157 vdd1.t281 8.126
R14775 vdd1.n158 vdd1.t1000 8.126
R14776 vdd1.n158 vdd1.t1212 8.126
R14777 vdd1.n159 vdd1.t881 8.126
R14778 vdd1.n159 vdd1.t1083 8.126
R14779 vdd1.n160 vdd1.t676 8.126
R14780 vdd1.n160 vdd1.t876 8.126
R14781 vdd1.n161 vdd1.t115 8.126
R14782 vdd1.n161 vdd1.t315 8.126
R14783 vdd1.n162 vdd1.t1199 8.126
R14784 vdd1.n162 vdd1.t1407 8.126
R14785 vdd1.n163 vdd1.t630 8.126
R14786 vdd1.n163 vdd1.t831 8.126
R14787 vdd1.n164 vdd1.t7 8.126
R14788 vdd1.n164 vdd1.t202 8.126
R14789 vdd1.n165 vdd1.t931 8.126
R14790 vdd1.n165 vdd1.t1131 8.126
R14791 vdd1.n166 vdd1.t794 8.126
R14792 vdd1.n166 vdd1.t1001 8.126
R14793 vdd1.n168 vdd1.t1031 8.126
R14794 vdd1.n168 vdd1.t1243 8.126
R14795 vdd1.n169 vdd1.t471 8.126
R14796 vdd1.n169 vdd1.t672 8.126
R14797 vdd1.n170 vdd1.t350 8.126
R14798 vdd1.n170 vdd1.t553 8.126
R14799 vdd1.n171 vdd1.t138 8.126
R14800 vdd1.n171 vdd1.t339 8.126
R14801 vdd1.n172 vdd1.t1063 8.126
R14802 vdd1.n172 vdd1.t1275 8.126
R14803 vdd1.n173 vdd1.t655 8.126
R14804 vdd1.n173 vdd1.t859 8.126
R14805 vdd1.n174 vdd1.t101 8.126
R14806 vdd1.n174 vdd1.t301 8.126
R14807 vdd1.n175 vdd1.t953 8.126
R14808 vdd1.n175 vdd1.t1157 8.126
R14809 vdd1.n176 vdd1.t389 8.126
R14810 vdd1.n176 vdd1.t590 8.126
R14811 vdd1.n177 vdd1.t273 8.126
R14812 vdd1.n177 vdd1.t472 8.126
R14813 vdd1.n179 vdd1.t625 8.126
R14814 vdd1.n179 vdd1.t824 8.126
R14815 vdd1.n180 vdd1.t70 8.126
R14816 vdd1.n180 vdd1.t272 8.126
R14817 vdd1.n181 vdd1.t1448 8.126
R14818 vdd1.n181 vdd1.t149 8.126
R14819 vdd1.n182 vdd1.t1230 8.126
R14820 vdd1.n182 vdd1.t1439 8.126
R14821 vdd1.n183 vdd1.t659 8.126
R14822 vdd1.n183 vdd1.t861 8.126
R14823 vdd1.n184 vdd1.t255 8.126
R14824 vdd1.n184 vdd1.t452 8.126
R14825 vdd1.n185 vdd1.t1189 8.126
R14826 vdd1.n185 vdd1.t1396 8.126
R14827 vdd1.n186 vdd1.t549 8.126
R14828 vdd1.n186 vdd1.t746 8.126
R14829 vdd1.n187 vdd1.t1493 8.126
R14830 vdd1.n187 vdd1.t191 8.126
R14831 vdd1.n188 vdd1.t1362 8.126
R14832 vdd1.n188 vdd1.t71 8.126
R14833 vdd1.n190 vdd1.t856 8.126
R14834 vdd1.n190 vdd1.t419 8.126
R14835 vdd1.n191 vdd1.t299 8.126
R14836 vdd1.n191 vdd1.t1361 8.126
R14837 vdd1.n192 vdd1.t176 8.126
R14838 vdd1.n192 vdd1.t1236 8.126
R14839 vdd1.n193 vdd1.t1471 8.126
R14840 vdd1.n193 vdd1.t1020 8.126
R14841 vdd1.n194 vdd1.t895 8.126
R14842 vdd1.n194 vdd1.t456 8.126
R14843 vdd1.n195 vdd1.t488 8.126
R14844 vdd1.n195 vdd1.t52 8.126
R14845 vdd1.n196 vdd1.t1430 8.126
R14846 vdd1.n196 vdd1.t979 8.126
R14847 vdd1.n197 vdd1.t777 8.126
R14848 vdd1.n197 vdd1.t344 8.126
R14849 vdd1.n198 vdd1.t221 8.126
R14850 vdd1.n198 vdd1.t1280 8.126
R14851 vdd1.n199 vdd1.t99 8.126
R14852 vdd1.n199 vdd1.t1150 8.126
R14853 vdd1.n201 vdd1.t450 8.126
R14854 vdd1.n201 vdd1.t654 8.126
R14855 vdd1.n202 vdd1.t1392 8.126
R14856 vdd1.n202 vdd1.t98 8.126
R14857 vdd1.n203 vdd1.t1265 8.126
R14858 vdd1.n203 vdd1.t1479 8.126
R14859 vdd1.n204 vdd1.t1052 8.126
R14860 vdd1.n204 vdd1.t1260 8.126
R14861 vdd1.n205 vdd1.t490 8.126
R14862 vdd1.n205 vdd1.t689 8.126
R14863 vdd1.n206 vdd1.t84 8.126
R14864 vdd1.n206 vdd1.t285 8.126
R14865 vdd1.n207 vdd1.t1007 8.126
R14866 vdd1.n207 vdd1.t1219 8.126
R14867 vdd1.n208 vdd1.t374 8.126
R14868 vdd1.n208 vdd1.t580 8.126
R14869 vdd1.n209 vdd1.t1314 8.126
R14870 vdd1.n209 vdd1.t22 8.126
R14871 vdd1.n210 vdd1.t1184 8.126
R14872 vdd1.n210 vdd1.t1393 8.126
R14873 vdd1.n212 vdd1.t49 8.126
R14874 vdd1.n212 vdd1.t252 8.126
R14875 vdd1.n213 vdd1.t970 8.126
R14876 vdd1.n213 vdd1.t1183 8.126
R14877 vdd1.n214 vdd1.t848 8.126
R14878 vdd1.n214 vdd1.t1056 8.126
R14879 vdd1.n215 vdd1.t647 8.126
R14880 vdd1.n215 vdd1.t846 8.126
R14881 vdd1.n216 vdd1.t85 8.126
R14882 vdd1.n216 vdd1.t286 8.126
R14883 vdd1.n217 vdd1.t1167 8.126
R14884 vdd1.n217 vdd1.t1378 8.126
R14885 vdd1.n218 vdd1.t597 8.126
R14886 vdd1.n218 vdd1.t799 8.126
R14887 vdd1.n219 vdd1.t1472 8.126
R14888 vdd1.n219 vdd1.t170 8.126
R14889 vdd1.n220 vdd1.t898 8.126
R14890 vdd1.n220 vdd1.t1100 8.126
R14891 vdd1.n221 vdd1.t767 8.126
R14892 vdd1.n221 vdd1.t971 8.126
R14893 vdd1.n223 vdd1.t117 8.126
R14894 vdd1.n223 vdd1.t317 8.126
R14895 vdd1.n224 vdd1.t1045 8.126
R14896 vdd1.n224 vdd1.t1255 8.126
R14897 vdd1.n225 vdd1.t923 8.126
R14898 vdd1.n225 vdd1.t1123 8.126
R14899 vdd1.n226 vdd1.t706 8.126
R14900 vdd1.n226 vdd1.t913 8.126
R14901 vdd1.n227 vdd1.t153 8.126
R14902 vdd1.n227 vdd1.t354 8.126
R14903 vdd1.n228 vdd1.t1239 8.126
R14904 vdd1.n228 vdd1.t1451 8.126
R14905 vdd1.n229 vdd1.t670 8.126
R14906 vdd1.n229 vdd1.t873 8.126
R14907 vdd1.n230 vdd1.t37 8.126
R14908 vdd1.n230 vdd1.t240 8.126
R14909 vdd1.n231 vdd1.t961 8.126
R14910 vdd1.n231 vdd1.t1165 8.126
R14911 vdd1.n232 vdd1.t840 8.126
R14912 vdd1.n232 vdd1.t1046 8.126
R14913 vdd1.n234 vdd1.t1202 8.126
R14914 vdd1.n234 vdd1.t1412 8.126
R14915 vdd1.n235 vdd1.t637 8.126
R14916 vdd1.n235 vdd1.t839 8.126
R14917 vdd1.n236 vdd1.t517 8.126
R14918 vdd1.n236 vdd1.t716 8.126
R14919 vdd1.n237 vdd1.t305 8.126
R14920 vdd1.n237 vdd1.t510 8.126
R14921 vdd1.n238 vdd1.t1242 8.126
R14922 vdd1.n238 vdd1.t1454 8.126
R14923 vdd1.n239 vdd1.t821 8.126
R14924 vdd1.n239 vdd1.t1029 8.126
R14925 vdd1.n240 vdd1.t267 8.126
R14926 vdd1.n240 vdd1.t468 8.126
R14927 vdd1.n241 vdd1.t1120 8.126
R14928 vdd1.n241 vdd1.t1333 8.126
R14929 vdd1.n242 vdd1.t562 8.126
R14930 vdd1.n242 vdd1.t758 8.126
R14931 vdd1.n243 vdd1.t432 8.126
R14932 vdd1.n243 vdd1.t638 8.126
R14933 vdd1.n245 vdd1.t1450 8.126
R14934 vdd1.n245 vdd1.t151 8.126
R14935 vdd1.n246 vdd1.t871 8.126
R14936 vdd1.n246 vdd1.t1075 8.126
R14937 vdd1.n247 vdd1.t744 8.126
R14938 vdd1.n247 vdd1.t949 8.126
R14939 vdd1.n248 vdd1.t540 8.126
R14940 vdd1.n248 vdd1.t734 8.126
R14941 vdd1.n249 vdd1.t1483 8.126
R14942 vdd1.n249 vdd1.t179 8.126
R14943 vdd1.n250 vdd1.t1059 8.126
R14944 vdd1.n250 vdd1.t1270 8.126
R14945 vdd1.n251 vdd1.t501 8.126
R14946 vdd1.n251 vdd1.t699 8.126
R14947 vdd1.n252 vdd1.t1367 8.126
R14948 vdd1.n252 vdd1.t74 8.126
R14949 vdd1.n253 vdd1.t785 8.126
R14950 vdd1.n253 vdd1.t988 8.126
R14951 vdd1.n254 vdd1.t668 8.126
R14952 vdd1.n254 vdd1.t872 8.126
R14953 vdd1.n256 vdd1.t1025 8.126
R14954 vdd1.n256 vdd1.t1237 8.126
R14955 vdd1.n257 vdd1.t463 8.126
R14956 vdd1.n257 vdd1.t667 8.126
R14957 vdd1.n258 vdd1.t342 8.126
R14958 vdd1.n258 vdd1.t547 8.126
R14959 vdd1.n259 vdd1.t136 8.126
R14960 vdd1.n259 vdd1.t336 8.126
R14961 vdd1.n260 vdd1.t1060 8.126
R14962 vdd1.n260 vdd1.t1271 8.126
R14963 vdd1.n261 vdd1.t651 8.126
R14964 vdd1.n261 vdd1.t851 8.126
R14965 vdd1.n262 vdd1.t93 8.126
R14966 vdd1.n262 vdd1.t293 8.126
R14967 vdd1.n263 vdd1.t947 8.126
R14968 vdd1.n263 vdd1.t1153 8.126
R14969 vdd1.n264 vdd1.t385 8.126
R14970 vdd1.n264 vdd1.t589 8.126
R14971 vdd1.n265 vdd1.t261 8.126
R14972 vdd1.n265 vdd1.t464 8.126
R14973 vdd1.n267 vdd1.t1267 8.126
R14974 vdd1.n267 vdd1.t817 8.126
R14975 vdd1.n268 vdd1.t696 8.126
R14976 vdd1.n268 vdd1.t260 8.126
R14977 vdd1.n269 vdd1.t576 8.126
R14978 vdd1.n269 vdd1.t141 8.126
R14979 vdd1.n270 vdd1.t365 8.126
R14980 vdd1.n270 vdd1.t1435 8.126
R14981 vdd1.n271 vdd1.t1305 8.126
R14982 vdd1.n271 vdd1.t854 8.126
R14983 vdd1.n272 vdd1.t886 8.126
R14984 vdd1.n272 vdd1.t445 8.126
R14985 vdd1.n273 vdd1.t328 8.126
R14986 vdd1.n273 vdd1.t1385 8.126
R14987 vdd1.n274 vdd1.t1187 8.126
R14988 vdd1.n274 vdd1.t738 8.126
R14989 vdd1.n275 vdd1.t615 8.126
R14990 vdd1.n275 vdd1.t182 8.126
R14991 vdd1.n276 vdd1.t497 8.126
R14992 vdd1.n276 vdd1.t58 8.126
R14993 vdd1.n278 vdd1.t685 8.126
R14994 vdd1.n278 vdd1.t891 8.126
R14995 vdd1.n279 vdd1.t131 8.126
R14996 vdd1.n279 vdd1.t332 8.126
R14997 vdd1.n280 vdd1.t13 8.126
R14998 vdd1.n280 vdd1.t212 8.126
R14999 vdd1.n281 vdd1.t1291 8.126
R15000 vdd1.n281 vdd1.t5 8.126
R15001 vdd1.n282 vdd1.t720 8.126
R15002 vdd1.n282 vdd1.t930 8.126
R15003 vdd1.n283 vdd1.t314 8.126
R15004 vdd1.n283 vdd1.t522 8.126
R15005 vdd1.n284 vdd1.t1253 8.126
R15006 vdd1.n284 vdd1.t1465 8.126
R15007 vdd1.n285 vdd1.t610 8.126
R15008 vdd1.n285 vdd1.t809 8.126
R15009 vdd1.n286 vdd1.t45 8.126
R15010 vdd1.n286 vdd1.t249 8.126
R15011 vdd1.n287 vdd1.t1426 8.126
R15012 vdd1.n287 vdd1.t132 8.126
R15013 vdd1.n289 vdd1.t282 8.126
R15014 vdd1.n289 vdd1.t485 8.126
R15015 vdd1.n290 vdd1.t1214 8.126
R15016 vdd1.n290 vdd1.t1425 8.126
R15017 vdd1.n291 vdd1.t1086 8.126
R15018 vdd1.n291 vdd1.t1300 8.126
R15019 vdd1.n292 vdd1.t877 8.126
R15020 vdd1.n292 vdd1.t1079 8.126
R15021 vdd1.n293 vdd1.t316 8.126
R15022 vdd1.n293 vdd1.t524 8.126
R15023 vdd1.n294 vdd1.t1408 8.126
R15024 vdd1.n294 vdd1.t114 8.126
R15025 vdd1.n295 vdd1.t834 8.126
R15026 vdd1.n295 vdd1.t1043 8.126
R15027 vdd1.n296 vdd1.t207 8.126
R15028 vdd1.n296 vdd1.t405 8.126
R15029 vdd1.n297 vdd1.t1132 8.126
R15030 vdd1.n297 vdd1.t1342 8.126
R15031 vdd1.n298 vdd1.t1002 8.126
R15032 vdd1.n298 vdd1.t1215 8.126
R15033 vdd1.n300 vdd1.t518 8.126
R15034 vdd1.n300 vdd1.t717 8.126
R15035 vdd1.n301 vdd1.t1461 8.126
R15036 vdd1.n301 vdd1.t162 8.126
R15037 vdd1.n302 vdd1.t1330 8.126
R15038 vdd1.n302 vdd1.t35 8.126
R15039 vdd1.n303 vdd1.t1109 8.126
R15040 vdd1.n303 vdd1.t1321 8.126
R15041 vdd1.n304 vdd1.t554 8.126
R15042 vdd1.n304 vdd1.t749 8.126
R15043 vdd1.n305 vdd1.t145 8.126
R15044 vdd1.n305 vdd1.t348 8.126
R15045 vdd1.n306 vdd1.t1073 8.126
R15046 vdd1.n306 vdd1.t1286 8.126
R15047 vdd1.n307 vdd1.t435 8.126
R15048 vdd1.n307 vdd1.t640 8.126
R15049 vdd1.n308 vdd1.t1371 8.126
R15050 vdd1.n308 vdd1.t76 8.126
R15051 vdd1.n309 vdd1.t1249 8.126
R15052 vdd1.n309 vdd1.t1462 8.126
R15053 vdd1.n311 vdd1.t110 8.126
R15054 vdd1.n311 vdd1.t310 8.126
R15055 vdd1.n312 vdd1.t1035 8.126
R15056 vdd1.n312 vdd1.t1248 8.126
R15057 vdd1.n313 vdd1.t916 8.126
R15058 vdd1.n313 vdd1.t1116 8.126
R15059 vdd1.n314 vdd1.t703 8.126
R15060 vdd1.n314 vdd1.t910 8.126
R15061 vdd1.n315 vdd1.t150 8.126
R15062 vdd1.n315 vdd1.t351 8.126
R15063 vdd1.n316 vdd1.t1233 8.126
R15064 vdd1.n316 vdd1.t1444 8.126
R15065 vdd1.n317 vdd1.t663 8.126
R15066 vdd1.n317 vdd1.t868 8.126
R15067 vdd1.n318 vdd1.t32 8.126
R15068 vdd1.n318 vdd1.t235 8.126
R15069 vdd1.n319 vdd1.t956 8.126
R15070 vdd1.n319 vdd1.t1160 8.126
R15071 vdd1.n320 vdd1.t830 8.126
R15072 vdd1.n320 vdd1.t1036 8.126
R15073 vdd1.n27 vdd1.t345 8.126
R15074 vdd1.n27 vdd1.t1406 8.126
R15075 vdd1.n28 vdd1.t1281 8.126
R15076 vdd1.n28 vdd1.t829 8.126
R15077 vdd1.n29 vdd1.t1149 8.126
R15078 vdd1.n29 vdd1.t708 8.126
R15079 vdd1.n30 vdd1.t938 8.126
R15080 vdd1.n30 vdd1.t507 8.126
R15081 vdd1.n31 vdd1.t379 8.126
R15082 vdd1.n31 vdd1.t1449 8.126
R15083 vdd1.n32 vdd1.t1475 8.126
R15084 vdd1.n32 vdd1.t1023 8.126
R15085 vdd1.n33 vdd1.t902 8.126
R15086 vdd1.n33 vdd1.t459 8.126
R15087 vdd1.n34 vdd1.t265 8.126
R15088 vdd1.n34 vdd1.t1326 8.126
R15089 vdd1.n35 vdd1.t1193 8.126
R15090 vdd1.n35 vdd1.t752 8.126
R15091 vdd1.n36 vdd1.t1068 8.126
R15092 vdd1.n36 vdd1.t629 8.126
R15093 vdd1.n323 vdd1.t1268 8.126
R15094 vdd1.n323 vdd1.t1482 8.126
R15095 vdd1.n324 vdd1.t697 8.126
R15096 vdd1.n324 vdd1.t907 8.126
R15097 vdd1.n325 vdd1.t577 8.126
R15098 vdd1.n325 vdd1.t775 8.126
R15099 vdd1.n326 vdd1.t366 8.126
R15100 vdd1.n326 vdd1.t571 8.126
R15101 vdd1.n327 vdd1.t1306 8.126
R15102 vdd1.n327 vdd1.t17 8.126
R15103 vdd1.n328 vdd1.t887 8.126
R15104 vdd1.n328 vdd1.t1091 8.126
R15105 vdd1.n329 vdd1.t329 8.126
R15106 vdd1.n329 vdd1.t537 8.126
R15107 vdd1.n330 vdd1.t1188 8.126
R15108 vdd1.n330 vdd1.t1398 8.126
R15109 vdd1.n331 vdd1.t616 8.126
R15110 vdd1.n331 vdd1.t813 8.126
R15111 vdd1.n332 vdd1.t498 8.126
R15112 vdd1.n332 vdd1.t698 8.126
R15113 vdd1.n334 vdd1.t16 8.126
R15114 vdd1.n334 vdd1.t1057 8.126
R15115 vdd1.n335 vdd1.t937 8.126
R15116 vdd1.n335 vdd1.t496 8.126
R15117 vdd1.n336 vdd1.t806 8.126
R15118 vdd1.n336 vdd1.t372 8.126
R15119 vdd1.n337 vdd1.t596 8.126
R15120 vdd1.n337 vdd1.t164 8.126
R15121 vdd1.n338 vdd1.t39 8.126
R15122 vdd1.n338 vdd1.t1093 8.126
R15123 vdd1.n339 vdd1.t1122 8.126
R15124 vdd1.n339 vdd1.t682 8.126
R15125 vdd1.n340 vdd1.t565 8.126
R15126 vdd1.n340 vdd1.t127 8.126
R15127 vdd1.n341 vdd1.t1429 8.126
R15128 vdd1.n341 vdd1.t978 8.126
R15129 vdd1.n342 vdd1.t844 8.126
R15130 vdd1.n342 vdd1.t411 8.126
R15131 vdd1.n343 vdd1.t730 8.126
R15132 vdd1.n343 vdd1.t292 8.126
R15133 vdd1.n345 vdd1.t1088 8.126
R15134 vdd1.n345 vdd1.t1303 8.126
R15135 vdd1.n346 vdd1.t532 8.126
R15136 vdd1.n346 vdd1.t729 8.126
R15137 vdd1.n347 vdd1.t400 8.126
R15138 vdd1.n347 vdd1.t606 8.126
R15139 vdd1.n348 vdd1.t195 8.126
R15140 vdd1.n348 vdd1.t393 8.126
R15141 vdd1.n349 vdd1.t1124 8.126
R15142 vdd1.n349 vdd1.t1336 8.126
R15143 vdd1.n350 vdd1.t711 8.126
R15144 vdd1.n350 vdd1.t920 8.126
R15145 vdd1.n351 vdd1.t158 8.126
R15146 vdd1.n351 vdd1.t362 8.126
R15147 vdd1.n352 vdd1.t1006 8.126
R15148 vdd1.n352 vdd1.t1218 8.126
R15149 vdd1.n353 vdd1.t439 8.126
R15150 vdd1.n353 vdd1.t645 8.126
R15151 vdd1.n354 vdd1.t324 8.126
R15152 vdd1.n354 vdd1.t534 8.126
R15153 vdd1.n356 vdd1.t680 8.126
R15154 vdd1.n356 vdd1.t883 8.126
R15155 vdd1.n357 vdd1.t122 8.126
R15156 vdd1.n357 vdd1.t322 8.126
R15157 vdd1.n358 vdd1.t6 8.126
R15158 vdd1.n358 vdd1.t201 8.126
R15159 vdd1.n359 vdd1.t1288 8.126
R15160 vdd1.n359 vdd1.t1497 8.126
R15161 vdd1.n360 vdd1.t715 8.126
R15162 vdd1.n360 vdd1.t922 8.126
R15163 vdd1.n361 vdd1.t308 8.126
R15164 vdd1.n361 vdd1.t513 8.126
R15165 vdd1.n362 vdd1.t1246 8.126
R15166 vdd1.n362 vdd1.t1457 8.126
R15167 vdd1.n363 vdd1.t599 8.126
R15168 vdd1.n363 vdd1.t797 8.126
R15169 vdd1.n364 vdd1.t40 8.126
R15170 vdd1.n364 vdd1.t242 8.126
R15171 vdd1.n365 vdd1.t1418 8.126
R15172 vdd1.n365 vdd1.t123 8.126
R15173 vdd1.n367 vdd1.t918 8.126
R15174 vdd1.n367 vdd1.t1119 8.126
R15175 vdd1.n368 vdd1.t358 8.126
R15176 vdd1.n368 vdd1.t561 8.126
R15177 vdd1.n369 vdd1.t232 8.126
R15178 vdd1.n369 vdd1.t431 8.126
R15179 vdd1.n370 vdd1.t25 8.126
R15180 vdd1.n370 vdd1.t224 8.126
R15181 vdd1.n371 vdd1.t951 8.126
R15182 vdd1.n371 vdd1.t1155 8.126
R15183 vdd1.n372 vdd1.t544 8.126
R15184 vdd1.n372 vdd1.t741 8.126
R15185 vdd1.n373 vdd1.t1488 8.126
R15186 vdd1.n373 vdd1.t186 8.126
R15187 vdd1.n374 vdd1.t833 8.126
R15188 vdd1.n374 vdd1.t1040 8.126
R15189 vdd1.n375 vdd1.t275 8.126
R15190 vdd1.n375 vdd1.t474 8.126
R15191 vdd1.n376 vdd1.t155 8.126
R15192 vdd1.n376 vdd1.t359 8.126
R15193 vdd1.n378 vdd1.t346 8.126
R15194 vdd1.n378 vdd1.t551 8.126
R15195 vdd1.n379 vdd1.t1282 8.126
R15196 vdd1.n379 vdd1.t1494 8.126
R15197 vdd1.n380 vdd1.t1151 8.126
R15198 vdd1.n380 vdd1.t1364 8.126
R15199 vdd1.n381 vdd1.t939 8.126
R15200 vdd1.n381 vdd1.t1141 8.126
R15201 vdd1.n382 vdd1.t380 8.126
R15202 vdd1.n382 vdd1.t583 8.126
R15203 vdd1.n383 vdd1.t1476 8.126
R15204 vdd1.n383 vdd1.t173 8.126
R15205 vdd1.n384 vdd1.t903 8.126
R15206 vdd1.n384 vdd1.t1104 8.126
R15207 vdd1.n385 vdd1.t266 8.126
R15208 vdd1.n385 vdd1.t467 8.126
R15209 vdd1.n386 vdd1.t1194 8.126
R15210 vdd1.n386 vdd1.t1400 8.126
R15211 vdd1.n387 vdd1.t1069 8.126
R15212 vdd1.n387 vdd1.t1283 8.126
R15213 vdd1.n389 vdd1.t581 8.126
R15214 vdd1.n389 vdd1.t142 8.126
R15215 vdd1.n390 vdd1.t23 8.126
R15216 vdd1.n390 vdd1.t1067 8.126
R15217 vdd1.n391 vdd1.t1391 8.126
R15218 vdd1.n391 vdd1.t945 8.126
R15219 vdd1.n392 vdd1.t1173 8.126
R15220 vdd1.n392 vdd1.t731 8.126
R15221 vdd1.n393 vdd1.t612 8.126
R15222 vdd1.n393 vdd1.t177 8.126
R15223 vdd1.n394 vdd1.t209 8.126
R15224 vdd1.n394 vdd1.t1263 8.126
R15225 vdd1.n395 vdd1.t1135 8.126
R15226 vdd1.n395 vdd1.t693 8.126
R15227 vdd1.n396 vdd1.t500 8.126
R15228 vdd1.n396 vdd1.t63 8.126
R15229 vdd1.n397 vdd1.t1433 8.126
R15230 vdd1.n397 vdd1.t984 8.126
R15231 vdd1.n398 vdd1.t1317 8.126
R15232 vdd1.n398 vdd1.t865 8.126
R15233 vdd1.n400 vdd1.t169 8.126
R15234 vdd1.n400 vdd1.t375 8.126
R15235 vdd1.n401 vdd1.t1098 8.126
R15236 vdd1.n401 vdd1.t1315 8.126
R15237 vdd1.n402 vdd1.t974 8.126
R15238 vdd1.n402 vdd1.t1182 8.126
R15239 vdd1.n403 vdd1.t762 8.126
R15240 vdd1.n403 vdd1.t965 8.126
R15241 vdd1.n404 vdd1.t211 8.126
R15242 vdd1.n404 vdd1.t407 8.126
R15243 vdd1.n405 vdd1.t1295 8.126
R15244 vdd1.n405 vdd1.t10 8.126
R15245 vdd1.n406 vdd1.t723 8.126
R15246 vdd1.n406 vdd1.t934 8.126
R15247 vdd1.n407 vdd1.t92 8.126
R15248 vdd1.n407 vdd1.t295 8.126
R15249 vdd1.n408 vdd1.t1013 8.126
R15250 vdd1.n408 vdd1.t1224 8.126
R15251 vdd1.n409 vdd1.t897 8.126
R15252 vdd1.n409 vdd1.t1099 8.126
R15253 vdd1.n411 vdd1.t1261 8.126
R15254 vdd1.n411 vdd1.t1473 8.126
R15255 vdd1.n412 vdd1.t690 8.126
R15256 vdd1.n412 vdd1.t896 8.126
R15257 vdd1.n413 vdd1.t573 8.126
R15258 vdd1.n413 vdd1.t771 8.126
R15259 vdd1.n414 vdd1.t363 8.126
R15260 vdd1.n414 vdd1.t567 8.126
R15261 vdd1.n415 vdd1.t1302 8.126
R15262 vdd1.n415 vdd1.t12 8.126
R15263 vdd1.n416 vdd1.t880 8.126
R15264 vdd1.n416 vdd1.t1082 8.126
R15265 vdd1.n417 vdd1.t319 8.126
R15266 vdd1.n417 vdd1.t526 8.126
R15267 vdd1.n418 vdd1.t1176 8.126
R15268 vdd1.n418 vdd1.t1384 8.126
R15269 vdd1.n419 vdd1.t613 8.126
R15270 vdd1.n419 vdd1.t810 8.126
R15271 vdd1.n420 vdd1.t493 8.126
R15272 vdd1.n420 vdd1.t691 8.126
R15273 vdd1.n422 vdd1.t884 8.126
R15274 vdd1.n422 vdd1.t1089 8.126
R15275 vdd1.n423 vdd1.t323 8.126
R15276 vdd1.n423 vdd1.t533 8.126
R15277 vdd1.n424 vdd1.t205 8.126
R15278 vdd1.n424 vdd1.t401 8.126
R15279 vdd1.n425 vdd1.t1498 8.126
R15280 vdd1.n425 vdd1.t196 8.126
R15281 vdd1.n426 vdd1.t924 8.126
R15282 vdd1.n426 vdd1.t1125 8.126
R15283 vdd1.n427 vdd1.t514 8.126
R15284 vdd1.n427 vdd1.t712 8.126
R15285 vdd1.n428 vdd1.t1458 8.126
R15286 vdd1.n428 vdd1.t160 8.126
R15287 vdd1.n429 vdd1.t798 8.126
R15288 vdd1.n429 vdd1.t1008 8.126
R15289 vdd1.n430 vdd1.t243 8.126
R15290 vdd1.n430 vdd1.t440 8.126
R15291 vdd1.n431 vdd1.t124 8.126
R15292 vdd1.n431 vdd1.t325 8.126
R15293 vdd1.n433 vdd1.t311 8.126
R15294 vdd1.n433 vdd1.t519 8.126
R15295 vdd1.n434 vdd1.t1250 8.126
R15296 vdd1.n434 vdd1.t1463 8.126
R15297 vdd1.n435 vdd1.t1118 8.126
R15298 vdd1.n435 vdd1.t1332 8.126
R15299 vdd1.n436 vdd1.t911 8.126
R15300 vdd1.n436 vdd1.t1111 8.126
R15301 vdd1.n437 vdd1.t352 8.126
R15302 vdd1.n437 vdd1.t555 8.126
R15303 vdd1.n438 vdd1.t1447 8.126
R15304 vdd1.n438 vdd1.t148 8.126
R15305 vdd1.n439 vdd1.t870 8.126
R15306 vdd1.n439 vdd1.t1074 8.126
R15307 vdd1.n440 vdd1.t237 8.126
R15308 vdd1.n440 vdd1.t437 8.126
R15309 vdd1.n441 vdd1.t1161 8.126
R15310 vdd1.n441 vdd1.t1372 8.126
R15311 vdd1.n442 vdd1.t1039 8.126
R15312 vdd1.n442 vdd1.t1251 8.126
R15313 vdd1.n445 vdd1.t552 8.126
R15314 vdd1.n445 vdd1.t748 8.126
R15315 vdd1.n446 vdd1.t1495 8.126
R15316 vdd1.n446 vdd1.t192 8.126
R15317 vdd1.n447 vdd1.t1366 8.126
R15318 vdd1.n447 vdd1.t73 8.126
R15319 vdd1.n448 vdd1.t1142 8.126
R15320 vdd1.n448 vdd1.t1353 8.126
R15321 vdd1.n449 vdd1.t584 8.126
R15322 vdd1.n449 vdd1.t780 8.126
R15323 vdd1.n450 vdd1.t175 8.126
R15324 vdd1.n450 vdd1.t378 8.126
R15325 vdd1.n451 vdd1.t1106 8.126
R15326 vdd1.n451 vdd1.t1318 8.126
R15327 vdd1.n452 vdd1.t469 8.126
R15328 vdd1.n452 vdd1.t671 8.126
R15329 vdd1.n453 vdd1.t1401 8.126
R15330 vdd1.n453 vdd1.t105 8.126
R15331 vdd1.n454 vdd1.t1285 8.126
R15332 vdd1.n454 vdd1.t1496 8.126
R15333 vdd1.n457 vdd1.t143 8.126
R15334 vdd1.n457 vdd1.t347 8.126
R15335 vdd1.n458 vdd1.t1071 8.126
R15336 vdd1.n458 vdd1.t1284 8.126
R15337 vdd1.n459 vdd1.t946 8.126
R15338 vdd1.n459 vdd1.t1152 8.126
R15339 vdd1.n460 vdd1.t732 8.126
R15340 vdd1.n460 vdd1.t940 8.126
R15341 vdd1.n461 vdd1.t178 8.126
R15342 vdd1.n461 vdd1.t381 8.126
R15343 vdd1.n462 vdd1.t1266 8.126
R15344 vdd1.n462 vdd1.t1478 8.126
R15345 vdd1.n463 vdd1.t695 8.126
R15346 vdd1.n463 vdd1.t905 8.126
R15347 vdd1.n464 vdd1.t67 8.126
R15348 vdd1.n464 vdd1.t269 8.126
R15349 vdd1.n465 vdd1.t987 8.126
R15350 vdd1.n465 vdd1.t1195 8.126
R15351 vdd1.n466 vdd1.t866 8.126
R15352 vdd1.n466 vdd1.t1072 8.126
R15353 vdd1.n468 vdd1.t376 8.126
R15354 vdd1.n468 vdd1.t1442 8.126
R15355 vdd1.n469 vdd1.t1316 8.126
R15356 vdd1.n469 vdd1.t864 8.126
R15357 vdd1.n470 vdd1.t1186 8.126
R15358 vdd1.n470 vdd1.t737 8.126
R15359 vdd1.n471 vdd1.t967 8.126
R15360 vdd1.n471 vdd1.t539 8.126
R15361 vdd1.n472 vdd1.t409 8.126
R15362 vdd1.n472 vdd1.t1481 8.126
R15363 vdd1.n473 vdd1.t11 8.126
R15364 vdd1.n473 vdd1.t1055 8.126
R15365 vdd1.n474 vdd1.t935 8.126
R15366 vdd1.n474 vdd1.t494 8.126
R15367 vdd1.n475 vdd1.t296 8.126
R15368 vdd1.n475 vdd1.t1355 8.126
R15369 vdd1.n476 vdd1.t1225 8.126
R15370 vdd1.n476 vdd1.t783 8.126
R15371 vdd1.n477 vdd1.t1103 8.126
R15372 vdd1.n477 vdd1.t661 8.126
R15373 vdd1.n479 vdd1.t1474 8.126
R15374 vdd1.n479 vdd1.t171 8.126
R15375 vdd1.n480 vdd1.t899 8.126
R15376 vdd1.n480 vdd1.t1101 8.126
R15377 vdd1.n481 vdd1.t772 8.126
R15378 vdd1.n481 vdd1.t976 8.126
R15379 vdd1.n482 vdd1.t568 8.126
R15380 vdd1.n482 vdd1.t763 8.126
R15381 vdd1.n483 vdd1.t15 8.126
R15382 vdd1.n483 vdd1.t214 8.126
R15383 vdd1.n484 vdd1.t1085 8.126
R15384 vdd1.n484 vdd1.t1298 8.126
R15385 vdd1.n485 vdd1.t530 8.126
R15386 vdd1.n485 vdd1.t726 8.126
R15387 vdd1.n486 vdd1.t1386 8.126
R15388 vdd1.n486 vdd1.t94 8.126
R15389 vdd1.n487 vdd1.t811 8.126
R15390 vdd1.n487 vdd1.t1014 8.126
R15391 vdd1.n488 vdd1.t692 8.126
R15392 vdd1.n488 vdd1.t900 8.126
R15393 vdd1.n0 vdd1.t885 8.126
R15394 vdd1.n0 vdd1.t1090 8.126
R15395 vdd1.n1 vdd1.t326 8.126
R15396 vdd1.n1 vdd1.t535 8.126
R15397 vdd1.n2 vdd1.t206 8.126
R15398 vdd1.n2 vdd1.t404 8.126
R15399 vdd1.n3 vdd1.t1499 8.126
R15400 vdd1.n3 vdd1.t197 8.126
R15401 vdd1.n4 vdd1.t925 8.126
R15402 vdd1.n4 vdd1.t1126 8.126
R15403 vdd1.n5 vdd1.t516 8.126
R15404 vdd1.n5 vdd1.t714 8.126
R15405 vdd1.n6 vdd1.t1460 8.126
R15406 vdd1.n6 vdd1.t161 8.126
R15407 vdd1.n7 vdd1.t802 8.126
R15408 vdd1.n7 vdd1.t1009 8.126
R15409 vdd1.n8 vdd1.t245 8.126
R15410 vdd1.n8 vdd1.t441 8.126
R15411 vdd1.n9 vdd1.t126 8.126
R15412 vdd1.n9 vdd1.t327 8.126
R15413 vdd1.n20 vdd1.n19 7.5
R15414 vdd1.n14 vdd1.n13 3.75
R15415 vdd1.n495 vdd1.n494 2.427
R15416 vdd1.n492 vdd1.n491 2.158
R15417 vdd1.n493 vdd1.n492 2.158
R15418 vdd1.n494 vdd1.n493 2.158
R15419 vdd1.n496 vdd1.n495 2.158
R15420 vdd1.n497 vdd1.n496 2.158
R15421 vdd1.n498 vdd1.n497 2.158
R15422 vdd1.n499 vdd1.n498 2.158
R15423 vdd1.n500 vdd1.n499 1.211
R15424 vdd1.n506 vdd1.n505 0.866
R15425 vdd1.n938 vdd1.n937 0.85
R15426 vdd1.n926 vdd1.n925 0.85
R15427 vdd1.n910 vdd1.n909 0.85
R15428 vdd1.n898 vdd1.n897 0.85
R15429 vdd1.n882 vdd1.n881 0.85
R15430 vdd1.n870 vdd1.n869 0.85
R15431 vdd1.n854 vdd1.n853 0.85
R15432 vdd1.n842 vdd1.n841 0.85
R15433 vdd1.n826 vdd1.n825 0.85
R15434 vdd1.n814 vdd1.n813 0.85
R15435 vdd1.n798 vdd1.n797 0.85
R15436 vdd1.n786 vdd1.n785 0.85
R15437 vdd1.n770 vdd1.n769 0.85
R15438 vdd1.n758 vdd1.n757 0.85
R15439 vdd1.n742 vdd1.n741 0.85
R15440 vdd1.n730 vdd1.n729 0.85
R15441 vdd1.n714 vdd1.n713 0.85
R15442 vdd1.n702 vdd1.n701 0.85
R15443 vdd1.n686 vdd1.n685 0.85
R15444 vdd1.n674 vdd1.n673 0.85
R15445 vdd1.n658 vdd1.n657 0.85
R15446 vdd1.n646 vdd1.n645 0.85
R15447 vdd1.n630 vdd1.n629 0.85
R15448 vdd1.n618 vdd1.n617 0.85
R15449 vdd1.n602 vdd1.n601 0.85
R15450 vdd1.n590 vdd1.n589 0.85
R15451 vdd1.n574 vdd1.n573 0.85
R15452 vdd1.n562 vdd1.n561 0.85
R15453 vdd1.n546 vdd1.n545 0.85
R15454 vdd1.n534 vdd1.n533 0.85
R15455 vdd1.n518 vdd1.n517 0.85
R15456 vdd1.n52 vdd1.n51 0.85
R15457 vdd1.n63 vdd1.n62 0.85
R15458 vdd1.n74 vdd1.n73 0.85
R15459 vdd1.n85 vdd1.n84 0.85
R15460 vdd1.n96 vdd1.n95 0.85
R15461 vdd1.n107 vdd1.n106 0.85
R15462 vdd1.n118 vdd1.n117 0.85
R15463 vdd1.n129 vdd1.n128 0.85
R15464 vdd1.n140 vdd1.n139 0.85
R15465 vdd1.n151 vdd1.n150 0.85
R15466 vdd1.n162 vdd1.n161 0.85
R15467 vdd1.n173 vdd1.n172 0.85
R15468 vdd1.n184 vdd1.n183 0.85
R15469 vdd1.n195 vdd1.n194 0.85
R15470 vdd1.n206 vdd1.n205 0.85
R15471 vdd1.n217 vdd1.n216 0.85
R15472 vdd1.n228 vdd1.n227 0.85
R15473 vdd1.n239 vdd1.n238 0.85
R15474 vdd1.n250 vdd1.n249 0.85
R15475 vdd1.n261 vdd1.n260 0.85
R15476 vdd1.n272 vdd1.n271 0.85
R15477 vdd1.n283 vdd1.n282 0.85
R15478 vdd1.n294 vdd1.n293 0.85
R15479 vdd1.n305 vdd1.n304 0.85
R15480 vdd1.n316 vdd1.n315 0.85
R15481 vdd1.n32 vdd1.n31 0.85
R15482 vdd1.n328 vdd1.n327 0.85
R15483 vdd1.n339 vdd1.n338 0.85
R15484 vdd1.n350 vdd1.n349 0.85
R15485 vdd1.n361 vdd1.n360 0.85
R15486 vdd1.n372 vdd1.n371 0.85
R15487 vdd1.n383 vdd1.n382 0.85
R15488 vdd1.n394 vdd1.n393 0.85
R15489 vdd1.n405 vdd1.n404 0.85
R15490 vdd1.n416 vdd1.n415 0.85
R15491 vdd1.n427 vdd1.n426 0.85
R15492 vdd1.n438 vdd1.n437 0.85
R15493 vdd1.n450 vdd1.n449 0.85
R15494 vdd1.n462 vdd1.n461 0.85
R15495 vdd1.n473 vdd1.n472 0.85
R15496 vdd1.n484 vdd1.n483 0.85
R15497 vdd1.n5 vdd1.n4 0.85
R15498 vdd1.n502 vdd1.n501 0.77
R15499 vdd1.n503 vdd1.n502 0.77
R15500 vdd1.n504 vdd1.n503 0.77
R15501 vdd1.n505 vdd1.n504 0.77
R15502 vdd1.n507 vdd1.n506 0.77
R15503 vdd1.n508 vdd1.n507 0.77
R15504 vdd1.n509 vdd1.n508 0.77
R15505 vdd1.n510 vdd1.n509 0.77
R15506 vdd1.n942 vdd1.n941 0.754
R15507 vdd1.n941 vdd1.n940 0.754
R15508 vdd1.n940 vdd1.n939 0.754
R15509 vdd1.n939 vdd1.n938 0.754
R15510 vdd1.n937 vdd1.n936 0.754
R15511 vdd1.n936 vdd1.n935 0.754
R15512 vdd1.n935 vdd1.n934 0.754
R15513 vdd1.n934 vdd1.n933 0.754
R15514 vdd1.n930 vdd1.n929 0.754
R15515 vdd1.n929 vdd1.n928 0.754
R15516 vdd1.n928 vdd1.n927 0.754
R15517 vdd1.n927 vdd1.n926 0.754
R15518 vdd1.n925 vdd1.n924 0.754
R15519 vdd1.n924 vdd1.n923 0.754
R15520 vdd1.n923 vdd1.n922 0.754
R15521 vdd1.n922 vdd1.n921 0.754
R15522 vdd1.n914 vdd1.n913 0.754
R15523 vdd1.n913 vdd1.n912 0.754
R15524 vdd1.n912 vdd1.n911 0.754
R15525 vdd1.n911 vdd1.n910 0.754
R15526 vdd1.n909 vdd1.n908 0.754
R15527 vdd1.n908 vdd1.n907 0.754
R15528 vdd1.n907 vdd1.n906 0.754
R15529 vdd1.n906 vdd1.n905 0.754
R15530 vdd1.n902 vdd1.n901 0.754
R15531 vdd1.n901 vdd1.n900 0.754
R15532 vdd1.n900 vdd1.n899 0.754
R15533 vdd1.n899 vdd1.n898 0.754
R15534 vdd1.n897 vdd1.n896 0.754
R15535 vdd1.n896 vdd1.n895 0.754
R15536 vdd1.n895 vdd1.n894 0.754
R15537 vdd1.n894 vdd1.n893 0.754
R15538 vdd1.n886 vdd1.n885 0.754
R15539 vdd1.n885 vdd1.n884 0.754
R15540 vdd1.n884 vdd1.n883 0.754
R15541 vdd1.n883 vdd1.n882 0.754
R15542 vdd1.n881 vdd1.n880 0.754
R15543 vdd1.n880 vdd1.n879 0.754
R15544 vdd1.n879 vdd1.n878 0.754
R15545 vdd1.n878 vdd1.n877 0.754
R15546 vdd1.n874 vdd1.n873 0.754
R15547 vdd1.n873 vdd1.n872 0.754
R15548 vdd1.n872 vdd1.n871 0.754
R15549 vdd1.n871 vdd1.n870 0.754
R15550 vdd1.n869 vdd1.n868 0.754
R15551 vdd1.n868 vdd1.n867 0.754
R15552 vdd1.n867 vdd1.n866 0.754
R15553 vdd1.n866 vdd1.n865 0.754
R15554 vdd1.n858 vdd1.n857 0.754
R15555 vdd1.n857 vdd1.n856 0.754
R15556 vdd1.n856 vdd1.n855 0.754
R15557 vdd1.n855 vdd1.n854 0.754
R15558 vdd1.n853 vdd1.n852 0.754
R15559 vdd1.n852 vdd1.n851 0.754
R15560 vdd1.n851 vdd1.n850 0.754
R15561 vdd1.n850 vdd1.n849 0.754
R15562 vdd1.n846 vdd1.n845 0.754
R15563 vdd1.n845 vdd1.n844 0.754
R15564 vdd1.n844 vdd1.n843 0.754
R15565 vdd1.n843 vdd1.n842 0.754
R15566 vdd1.n841 vdd1.n840 0.754
R15567 vdd1.n840 vdd1.n839 0.754
R15568 vdd1.n839 vdd1.n838 0.754
R15569 vdd1.n838 vdd1.n837 0.754
R15570 vdd1.n830 vdd1.n829 0.754
R15571 vdd1.n829 vdd1.n828 0.754
R15572 vdd1.n828 vdd1.n827 0.754
R15573 vdd1.n827 vdd1.n826 0.754
R15574 vdd1.n825 vdd1.n824 0.754
R15575 vdd1.n824 vdd1.n823 0.754
R15576 vdd1.n823 vdd1.n822 0.754
R15577 vdd1.n822 vdd1.n821 0.754
R15578 vdd1.n818 vdd1.n817 0.754
R15579 vdd1.n817 vdd1.n816 0.754
R15580 vdd1.n816 vdd1.n815 0.754
R15581 vdd1.n815 vdd1.n814 0.754
R15582 vdd1.n813 vdd1.n812 0.754
R15583 vdd1.n812 vdd1.n811 0.754
R15584 vdd1.n811 vdd1.n810 0.754
R15585 vdd1.n810 vdd1.n809 0.754
R15586 vdd1.n802 vdd1.n801 0.754
R15587 vdd1.n801 vdd1.n800 0.754
R15588 vdd1.n800 vdd1.n799 0.754
R15589 vdd1.n799 vdd1.n798 0.754
R15590 vdd1.n797 vdd1.n796 0.754
R15591 vdd1.n796 vdd1.n795 0.754
R15592 vdd1.n795 vdd1.n794 0.754
R15593 vdd1.n794 vdd1.n793 0.754
R15594 vdd1.n790 vdd1.n789 0.754
R15595 vdd1.n789 vdd1.n788 0.754
R15596 vdd1.n788 vdd1.n787 0.754
R15597 vdd1.n787 vdd1.n786 0.754
R15598 vdd1.n785 vdd1.n784 0.754
R15599 vdd1.n784 vdd1.n783 0.754
R15600 vdd1.n783 vdd1.n782 0.754
R15601 vdd1.n782 vdd1.n781 0.754
R15602 vdd1.n774 vdd1.n773 0.754
R15603 vdd1.n773 vdd1.n772 0.754
R15604 vdd1.n772 vdd1.n771 0.754
R15605 vdd1.n771 vdd1.n770 0.754
R15606 vdd1.n769 vdd1.n768 0.754
R15607 vdd1.n768 vdd1.n767 0.754
R15608 vdd1.n767 vdd1.n766 0.754
R15609 vdd1.n766 vdd1.n765 0.754
R15610 vdd1.n762 vdd1.n761 0.754
R15611 vdd1.n761 vdd1.n760 0.754
R15612 vdd1.n760 vdd1.n759 0.754
R15613 vdd1.n759 vdd1.n758 0.754
R15614 vdd1.n757 vdd1.n756 0.754
R15615 vdd1.n756 vdd1.n755 0.754
R15616 vdd1.n755 vdd1.n754 0.754
R15617 vdd1.n754 vdd1.n753 0.754
R15618 vdd1.n746 vdd1.n745 0.754
R15619 vdd1.n745 vdd1.n744 0.754
R15620 vdd1.n744 vdd1.n743 0.754
R15621 vdd1.n743 vdd1.n742 0.754
R15622 vdd1.n741 vdd1.n740 0.754
R15623 vdd1.n740 vdd1.n739 0.754
R15624 vdd1.n739 vdd1.n738 0.754
R15625 vdd1.n738 vdd1.n737 0.754
R15626 vdd1.n734 vdd1.n733 0.754
R15627 vdd1.n733 vdd1.n732 0.754
R15628 vdd1.n732 vdd1.n731 0.754
R15629 vdd1.n731 vdd1.n730 0.754
R15630 vdd1.n729 vdd1.n728 0.754
R15631 vdd1.n728 vdd1.n727 0.754
R15632 vdd1.n727 vdd1.n726 0.754
R15633 vdd1.n726 vdd1.n725 0.754
R15634 vdd1.n718 vdd1.n717 0.754
R15635 vdd1.n717 vdd1.n716 0.754
R15636 vdd1.n716 vdd1.n715 0.754
R15637 vdd1.n715 vdd1.n714 0.754
R15638 vdd1.n713 vdd1.n712 0.754
R15639 vdd1.n712 vdd1.n711 0.754
R15640 vdd1.n711 vdd1.n710 0.754
R15641 vdd1.n710 vdd1.n709 0.754
R15642 vdd1.n706 vdd1.n705 0.754
R15643 vdd1.n705 vdd1.n704 0.754
R15644 vdd1.n704 vdd1.n703 0.754
R15645 vdd1.n703 vdd1.n702 0.754
R15646 vdd1.n701 vdd1.n700 0.754
R15647 vdd1.n700 vdd1.n699 0.754
R15648 vdd1.n699 vdd1.n698 0.754
R15649 vdd1.n698 vdd1.n697 0.754
R15650 vdd1.n690 vdd1.n689 0.754
R15651 vdd1.n689 vdd1.n688 0.754
R15652 vdd1.n688 vdd1.n687 0.754
R15653 vdd1.n687 vdd1.n686 0.754
R15654 vdd1.n685 vdd1.n684 0.754
R15655 vdd1.n684 vdd1.n683 0.754
R15656 vdd1.n683 vdd1.n682 0.754
R15657 vdd1.n682 vdd1.n681 0.754
R15658 vdd1.n678 vdd1.n677 0.754
R15659 vdd1.n677 vdd1.n676 0.754
R15660 vdd1.n676 vdd1.n675 0.754
R15661 vdd1.n675 vdd1.n674 0.754
R15662 vdd1.n673 vdd1.n672 0.754
R15663 vdd1.n672 vdd1.n671 0.754
R15664 vdd1.n671 vdd1.n670 0.754
R15665 vdd1.n670 vdd1.n669 0.754
R15666 vdd1.n662 vdd1.n661 0.754
R15667 vdd1.n661 vdd1.n660 0.754
R15668 vdd1.n660 vdd1.n659 0.754
R15669 vdd1.n659 vdd1.n658 0.754
R15670 vdd1.n657 vdd1.n656 0.754
R15671 vdd1.n656 vdd1.n655 0.754
R15672 vdd1.n655 vdd1.n654 0.754
R15673 vdd1.n654 vdd1.n653 0.754
R15674 vdd1.n650 vdd1.n649 0.754
R15675 vdd1.n649 vdd1.n648 0.754
R15676 vdd1.n648 vdd1.n647 0.754
R15677 vdd1.n647 vdd1.n646 0.754
R15678 vdd1.n645 vdd1.n644 0.754
R15679 vdd1.n644 vdd1.n643 0.754
R15680 vdd1.n643 vdd1.n642 0.754
R15681 vdd1.n642 vdd1.n641 0.754
R15682 vdd1.n634 vdd1.n633 0.754
R15683 vdd1.n633 vdd1.n632 0.754
R15684 vdd1.n632 vdd1.n631 0.754
R15685 vdd1.n631 vdd1.n630 0.754
R15686 vdd1.n629 vdd1.n628 0.754
R15687 vdd1.n628 vdd1.n627 0.754
R15688 vdd1.n627 vdd1.n626 0.754
R15689 vdd1.n626 vdd1.n625 0.754
R15690 vdd1.n622 vdd1.n621 0.754
R15691 vdd1.n621 vdd1.n620 0.754
R15692 vdd1.n620 vdd1.n619 0.754
R15693 vdd1.n619 vdd1.n618 0.754
R15694 vdd1.n617 vdd1.n616 0.754
R15695 vdd1.n616 vdd1.n615 0.754
R15696 vdd1.n615 vdd1.n614 0.754
R15697 vdd1.n614 vdd1.n613 0.754
R15698 vdd1.n606 vdd1.n605 0.754
R15699 vdd1.n605 vdd1.n604 0.754
R15700 vdd1.n604 vdd1.n603 0.754
R15701 vdd1.n603 vdd1.n602 0.754
R15702 vdd1.n601 vdd1.n600 0.754
R15703 vdd1.n600 vdd1.n599 0.754
R15704 vdd1.n599 vdd1.n598 0.754
R15705 vdd1.n598 vdd1.n597 0.754
R15706 vdd1.n594 vdd1.n593 0.754
R15707 vdd1.n593 vdd1.n592 0.754
R15708 vdd1.n592 vdd1.n591 0.754
R15709 vdd1.n591 vdd1.n590 0.754
R15710 vdd1.n589 vdd1.n588 0.754
R15711 vdd1.n588 vdd1.n587 0.754
R15712 vdd1.n587 vdd1.n586 0.754
R15713 vdd1.n586 vdd1.n585 0.754
R15714 vdd1.n578 vdd1.n577 0.754
R15715 vdd1.n577 vdd1.n576 0.754
R15716 vdd1.n576 vdd1.n575 0.754
R15717 vdd1.n575 vdd1.n574 0.754
R15718 vdd1.n573 vdd1.n572 0.754
R15719 vdd1.n572 vdd1.n571 0.754
R15720 vdd1.n571 vdd1.n570 0.754
R15721 vdd1.n570 vdd1.n569 0.754
R15722 vdd1.n566 vdd1.n565 0.754
R15723 vdd1.n565 vdd1.n564 0.754
R15724 vdd1.n564 vdd1.n563 0.754
R15725 vdd1.n563 vdd1.n562 0.754
R15726 vdd1.n561 vdd1.n560 0.754
R15727 vdd1.n560 vdd1.n559 0.754
R15728 vdd1.n559 vdd1.n558 0.754
R15729 vdd1.n558 vdd1.n557 0.754
R15730 vdd1.n550 vdd1.n549 0.754
R15731 vdd1.n549 vdd1.n548 0.754
R15732 vdd1.n548 vdd1.n547 0.754
R15733 vdd1.n547 vdd1.n546 0.754
R15734 vdd1.n545 vdd1.n544 0.754
R15735 vdd1.n544 vdd1.n543 0.754
R15736 vdd1.n543 vdd1.n542 0.754
R15737 vdd1.n542 vdd1.n541 0.754
R15738 vdd1.n538 vdd1.n537 0.754
R15739 vdd1.n537 vdd1.n536 0.754
R15740 vdd1.n536 vdd1.n535 0.754
R15741 vdd1.n535 vdd1.n534 0.754
R15742 vdd1.n533 vdd1.n532 0.754
R15743 vdd1.n532 vdd1.n531 0.754
R15744 vdd1.n531 vdd1.n530 0.754
R15745 vdd1.n530 vdd1.n529 0.754
R15746 vdd1.n522 vdd1.n521 0.754
R15747 vdd1.n521 vdd1.n520 0.754
R15748 vdd1.n520 vdd1.n519 0.754
R15749 vdd1.n519 vdd1.n518 0.754
R15750 vdd1.n517 vdd1.n516 0.754
R15751 vdd1.n516 vdd1.n515 0.754
R15752 vdd1.n515 vdd1.n514 0.754
R15753 vdd1.n514 vdd1.n513 0.754
R15754 vdd1.n56 vdd1.n55 0.754
R15755 vdd1.n55 vdd1.n54 0.754
R15756 vdd1.n54 vdd1.n53 0.754
R15757 vdd1.n53 vdd1.n52 0.754
R15758 vdd1.n51 vdd1.n50 0.754
R15759 vdd1.n50 vdd1.n49 0.754
R15760 vdd1.n49 vdd1.n48 0.754
R15761 vdd1.n48 vdd1.n47 0.754
R15762 vdd1.n67 vdd1.n66 0.754
R15763 vdd1.n66 vdd1.n65 0.754
R15764 vdd1.n65 vdd1.n64 0.754
R15765 vdd1.n64 vdd1.n63 0.754
R15766 vdd1.n62 vdd1.n61 0.754
R15767 vdd1.n61 vdd1.n60 0.754
R15768 vdd1.n60 vdd1.n59 0.754
R15769 vdd1.n59 vdd1.n58 0.754
R15770 vdd1.n78 vdd1.n77 0.754
R15771 vdd1.n77 vdd1.n76 0.754
R15772 vdd1.n76 vdd1.n75 0.754
R15773 vdd1.n75 vdd1.n74 0.754
R15774 vdd1.n73 vdd1.n72 0.754
R15775 vdd1.n72 vdd1.n71 0.754
R15776 vdd1.n71 vdd1.n70 0.754
R15777 vdd1.n70 vdd1.n69 0.754
R15778 vdd1.n89 vdd1.n88 0.754
R15779 vdd1.n88 vdd1.n87 0.754
R15780 vdd1.n87 vdd1.n86 0.754
R15781 vdd1.n86 vdd1.n85 0.754
R15782 vdd1.n84 vdd1.n83 0.754
R15783 vdd1.n83 vdd1.n82 0.754
R15784 vdd1.n82 vdd1.n81 0.754
R15785 vdd1.n81 vdd1.n80 0.754
R15786 vdd1.n100 vdd1.n99 0.754
R15787 vdd1.n99 vdd1.n98 0.754
R15788 vdd1.n98 vdd1.n97 0.754
R15789 vdd1.n97 vdd1.n96 0.754
R15790 vdd1.n95 vdd1.n94 0.754
R15791 vdd1.n94 vdd1.n93 0.754
R15792 vdd1.n93 vdd1.n92 0.754
R15793 vdd1.n92 vdd1.n91 0.754
R15794 vdd1.n111 vdd1.n110 0.754
R15795 vdd1.n110 vdd1.n109 0.754
R15796 vdd1.n109 vdd1.n108 0.754
R15797 vdd1.n108 vdd1.n107 0.754
R15798 vdd1.n106 vdd1.n105 0.754
R15799 vdd1.n105 vdd1.n104 0.754
R15800 vdd1.n104 vdd1.n103 0.754
R15801 vdd1.n103 vdd1.n102 0.754
R15802 vdd1.n122 vdd1.n121 0.754
R15803 vdd1.n121 vdd1.n120 0.754
R15804 vdd1.n120 vdd1.n119 0.754
R15805 vdd1.n119 vdd1.n118 0.754
R15806 vdd1.n117 vdd1.n116 0.754
R15807 vdd1.n116 vdd1.n115 0.754
R15808 vdd1.n115 vdd1.n114 0.754
R15809 vdd1.n114 vdd1.n113 0.754
R15810 vdd1.n133 vdd1.n132 0.754
R15811 vdd1.n132 vdd1.n131 0.754
R15812 vdd1.n131 vdd1.n130 0.754
R15813 vdd1.n130 vdd1.n129 0.754
R15814 vdd1.n128 vdd1.n127 0.754
R15815 vdd1.n127 vdd1.n126 0.754
R15816 vdd1.n126 vdd1.n125 0.754
R15817 vdd1.n125 vdd1.n124 0.754
R15818 vdd1.n144 vdd1.n143 0.754
R15819 vdd1.n143 vdd1.n142 0.754
R15820 vdd1.n142 vdd1.n141 0.754
R15821 vdd1.n141 vdd1.n140 0.754
R15822 vdd1.n139 vdd1.n138 0.754
R15823 vdd1.n138 vdd1.n137 0.754
R15824 vdd1.n137 vdd1.n136 0.754
R15825 vdd1.n136 vdd1.n135 0.754
R15826 vdd1.n155 vdd1.n154 0.754
R15827 vdd1.n154 vdd1.n153 0.754
R15828 vdd1.n153 vdd1.n152 0.754
R15829 vdd1.n152 vdd1.n151 0.754
R15830 vdd1.n150 vdd1.n149 0.754
R15831 vdd1.n149 vdd1.n148 0.754
R15832 vdd1.n148 vdd1.n147 0.754
R15833 vdd1.n147 vdd1.n146 0.754
R15834 vdd1.n166 vdd1.n165 0.754
R15835 vdd1.n165 vdd1.n164 0.754
R15836 vdd1.n164 vdd1.n163 0.754
R15837 vdd1.n163 vdd1.n162 0.754
R15838 vdd1.n161 vdd1.n160 0.754
R15839 vdd1.n160 vdd1.n159 0.754
R15840 vdd1.n159 vdd1.n158 0.754
R15841 vdd1.n158 vdd1.n157 0.754
R15842 vdd1.n177 vdd1.n176 0.754
R15843 vdd1.n176 vdd1.n175 0.754
R15844 vdd1.n175 vdd1.n174 0.754
R15845 vdd1.n174 vdd1.n173 0.754
R15846 vdd1.n172 vdd1.n171 0.754
R15847 vdd1.n171 vdd1.n170 0.754
R15848 vdd1.n170 vdd1.n169 0.754
R15849 vdd1.n169 vdd1.n168 0.754
R15850 vdd1.n188 vdd1.n187 0.754
R15851 vdd1.n187 vdd1.n186 0.754
R15852 vdd1.n186 vdd1.n185 0.754
R15853 vdd1.n185 vdd1.n184 0.754
R15854 vdd1.n183 vdd1.n182 0.754
R15855 vdd1.n182 vdd1.n181 0.754
R15856 vdd1.n181 vdd1.n180 0.754
R15857 vdd1.n180 vdd1.n179 0.754
R15858 vdd1.n199 vdd1.n198 0.754
R15859 vdd1.n198 vdd1.n197 0.754
R15860 vdd1.n197 vdd1.n196 0.754
R15861 vdd1.n196 vdd1.n195 0.754
R15862 vdd1.n194 vdd1.n193 0.754
R15863 vdd1.n193 vdd1.n192 0.754
R15864 vdd1.n192 vdd1.n191 0.754
R15865 vdd1.n191 vdd1.n190 0.754
R15866 vdd1.n210 vdd1.n209 0.754
R15867 vdd1.n209 vdd1.n208 0.754
R15868 vdd1.n208 vdd1.n207 0.754
R15869 vdd1.n207 vdd1.n206 0.754
R15870 vdd1.n205 vdd1.n204 0.754
R15871 vdd1.n204 vdd1.n203 0.754
R15872 vdd1.n203 vdd1.n202 0.754
R15873 vdd1.n202 vdd1.n201 0.754
R15874 vdd1.n221 vdd1.n220 0.754
R15875 vdd1.n220 vdd1.n219 0.754
R15876 vdd1.n219 vdd1.n218 0.754
R15877 vdd1.n218 vdd1.n217 0.754
R15878 vdd1.n216 vdd1.n215 0.754
R15879 vdd1.n215 vdd1.n214 0.754
R15880 vdd1.n214 vdd1.n213 0.754
R15881 vdd1.n213 vdd1.n212 0.754
R15882 vdd1.n232 vdd1.n231 0.754
R15883 vdd1.n231 vdd1.n230 0.754
R15884 vdd1.n230 vdd1.n229 0.754
R15885 vdd1.n229 vdd1.n228 0.754
R15886 vdd1.n227 vdd1.n226 0.754
R15887 vdd1.n226 vdd1.n225 0.754
R15888 vdd1.n225 vdd1.n224 0.754
R15889 vdd1.n224 vdd1.n223 0.754
R15890 vdd1.n243 vdd1.n242 0.754
R15891 vdd1.n242 vdd1.n241 0.754
R15892 vdd1.n241 vdd1.n240 0.754
R15893 vdd1.n240 vdd1.n239 0.754
R15894 vdd1.n238 vdd1.n237 0.754
R15895 vdd1.n237 vdd1.n236 0.754
R15896 vdd1.n236 vdd1.n235 0.754
R15897 vdd1.n235 vdd1.n234 0.754
R15898 vdd1.n254 vdd1.n253 0.754
R15899 vdd1.n253 vdd1.n252 0.754
R15900 vdd1.n252 vdd1.n251 0.754
R15901 vdd1.n251 vdd1.n250 0.754
R15902 vdd1.n249 vdd1.n248 0.754
R15903 vdd1.n248 vdd1.n247 0.754
R15904 vdd1.n247 vdd1.n246 0.754
R15905 vdd1.n246 vdd1.n245 0.754
R15906 vdd1.n265 vdd1.n264 0.754
R15907 vdd1.n264 vdd1.n263 0.754
R15908 vdd1.n263 vdd1.n262 0.754
R15909 vdd1.n262 vdd1.n261 0.754
R15910 vdd1.n260 vdd1.n259 0.754
R15911 vdd1.n259 vdd1.n258 0.754
R15912 vdd1.n258 vdd1.n257 0.754
R15913 vdd1.n257 vdd1.n256 0.754
R15914 vdd1.n276 vdd1.n275 0.754
R15915 vdd1.n275 vdd1.n274 0.754
R15916 vdd1.n274 vdd1.n273 0.754
R15917 vdd1.n273 vdd1.n272 0.754
R15918 vdd1.n271 vdd1.n270 0.754
R15919 vdd1.n270 vdd1.n269 0.754
R15920 vdd1.n269 vdd1.n268 0.754
R15921 vdd1.n268 vdd1.n267 0.754
R15922 vdd1.n287 vdd1.n286 0.754
R15923 vdd1.n286 vdd1.n285 0.754
R15924 vdd1.n285 vdd1.n284 0.754
R15925 vdd1.n284 vdd1.n283 0.754
R15926 vdd1.n282 vdd1.n281 0.754
R15927 vdd1.n281 vdd1.n280 0.754
R15928 vdd1.n280 vdd1.n279 0.754
R15929 vdd1.n279 vdd1.n278 0.754
R15930 vdd1.n298 vdd1.n297 0.754
R15931 vdd1.n297 vdd1.n296 0.754
R15932 vdd1.n296 vdd1.n295 0.754
R15933 vdd1.n295 vdd1.n294 0.754
R15934 vdd1.n293 vdd1.n292 0.754
R15935 vdd1.n292 vdd1.n291 0.754
R15936 vdd1.n291 vdd1.n290 0.754
R15937 vdd1.n290 vdd1.n289 0.754
R15938 vdd1.n309 vdd1.n308 0.754
R15939 vdd1.n308 vdd1.n307 0.754
R15940 vdd1.n307 vdd1.n306 0.754
R15941 vdd1.n306 vdd1.n305 0.754
R15942 vdd1.n304 vdd1.n303 0.754
R15943 vdd1.n303 vdd1.n302 0.754
R15944 vdd1.n302 vdd1.n301 0.754
R15945 vdd1.n301 vdd1.n300 0.754
R15946 vdd1.n320 vdd1.n319 0.754
R15947 vdd1.n319 vdd1.n318 0.754
R15948 vdd1.n318 vdd1.n317 0.754
R15949 vdd1.n317 vdd1.n316 0.754
R15950 vdd1.n315 vdd1.n314 0.754
R15951 vdd1.n314 vdd1.n313 0.754
R15952 vdd1.n313 vdd1.n312 0.754
R15953 vdd1.n312 vdd1.n311 0.754
R15954 vdd1.n36 vdd1.n35 0.754
R15955 vdd1.n35 vdd1.n34 0.754
R15956 vdd1.n34 vdd1.n33 0.754
R15957 vdd1.n33 vdd1.n32 0.754
R15958 vdd1.n31 vdd1.n30 0.754
R15959 vdd1.n30 vdd1.n29 0.754
R15960 vdd1.n29 vdd1.n28 0.754
R15961 vdd1.n28 vdd1.n27 0.754
R15962 vdd1.n332 vdd1.n331 0.754
R15963 vdd1.n331 vdd1.n330 0.754
R15964 vdd1.n330 vdd1.n329 0.754
R15965 vdd1.n329 vdd1.n328 0.754
R15966 vdd1.n327 vdd1.n326 0.754
R15967 vdd1.n326 vdd1.n325 0.754
R15968 vdd1.n325 vdd1.n324 0.754
R15969 vdd1.n324 vdd1.n323 0.754
R15970 vdd1.n343 vdd1.n342 0.754
R15971 vdd1.n342 vdd1.n341 0.754
R15972 vdd1.n341 vdd1.n340 0.754
R15973 vdd1.n340 vdd1.n339 0.754
R15974 vdd1.n338 vdd1.n337 0.754
R15975 vdd1.n337 vdd1.n336 0.754
R15976 vdd1.n336 vdd1.n335 0.754
R15977 vdd1.n335 vdd1.n334 0.754
R15978 vdd1.n354 vdd1.n353 0.754
R15979 vdd1.n353 vdd1.n352 0.754
R15980 vdd1.n352 vdd1.n351 0.754
R15981 vdd1.n351 vdd1.n350 0.754
R15982 vdd1.n349 vdd1.n348 0.754
R15983 vdd1.n348 vdd1.n347 0.754
R15984 vdd1.n347 vdd1.n346 0.754
R15985 vdd1.n346 vdd1.n345 0.754
R15986 vdd1.n365 vdd1.n364 0.754
R15987 vdd1.n364 vdd1.n363 0.754
R15988 vdd1.n363 vdd1.n362 0.754
R15989 vdd1.n362 vdd1.n361 0.754
R15990 vdd1.n360 vdd1.n359 0.754
R15991 vdd1.n359 vdd1.n358 0.754
R15992 vdd1.n358 vdd1.n357 0.754
R15993 vdd1.n357 vdd1.n356 0.754
R15994 vdd1.n376 vdd1.n375 0.754
R15995 vdd1.n375 vdd1.n374 0.754
R15996 vdd1.n374 vdd1.n373 0.754
R15997 vdd1.n373 vdd1.n372 0.754
R15998 vdd1.n371 vdd1.n370 0.754
R15999 vdd1.n370 vdd1.n369 0.754
R16000 vdd1.n369 vdd1.n368 0.754
R16001 vdd1.n368 vdd1.n367 0.754
R16002 vdd1.n387 vdd1.n386 0.754
R16003 vdd1.n386 vdd1.n385 0.754
R16004 vdd1.n385 vdd1.n384 0.754
R16005 vdd1.n384 vdd1.n383 0.754
R16006 vdd1.n382 vdd1.n381 0.754
R16007 vdd1.n381 vdd1.n380 0.754
R16008 vdd1.n380 vdd1.n379 0.754
R16009 vdd1.n379 vdd1.n378 0.754
R16010 vdd1.n398 vdd1.n397 0.754
R16011 vdd1.n397 vdd1.n396 0.754
R16012 vdd1.n396 vdd1.n395 0.754
R16013 vdd1.n395 vdd1.n394 0.754
R16014 vdd1.n393 vdd1.n392 0.754
R16015 vdd1.n392 vdd1.n391 0.754
R16016 vdd1.n391 vdd1.n390 0.754
R16017 vdd1.n390 vdd1.n389 0.754
R16018 vdd1.n409 vdd1.n408 0.754
R16019 vdd1.n408 vdd1.n407 0.754
R16020 vdd1.n407 vdd1.n406 0.754
R16021 vdd1.n406 vdd1.n405 0.754
R16022 vdd1.n404 vdd1.n403 0.754
R16023 vdd1.n403 vdd1.n402 0.754
R16024 vdd1.n402 vdd1.n401 0.754
R16025 vdd1.n401 vdd1.n400 0.754
R16026 vdd1.n420 vdd1.n419 0.754
R16027 vdd1.n419 vdd1.n418 0.754
R16028 vdd1.n418 vdd1.n417 0.754
R16029 vdd1.n417 vdd1.n416 0.754
R16030 vdd1.n415 vdd1.n414 0.754
R16031 vdd1.n414 vdd1.n413 0.754
R16032 vdd1.n413 vdd1.n412 0.754
R16033 vdd1.n412 vdd1.n411 0.754
R16034 vdd1.n431 vdd1.n430 0.754
R16035 vdd1.n430 vdd1.n429 0.754
R16036 vdd1.n429 vdd1.n428 0.754
R16037 vdd1.n428 vdd1.n427 0.754
R16038 vdd1.n426 vdd1.n425 0.754
R16039 vdd1.n425 vdd1.n424 0.754
R16040 vdd1.n424 vdd1.n423 0.754
R16041 vdd1.n423 vdd1.n422 0.754
R16042 vdd1.n442 vdd1.n441 0.754
R16043 vdd1.n441 vdd1.n440 0.754
R16044 vdd1.n440 vdd1.n439 0.754
R16045 vdd1.n439 vdd1.n438 0.754
R16046 vdd1.n437 vdd1.n436 0.754
R16047 vdd1.n436 vdd1.n435 0.754
R16048 vdd1.n435 vdd1.n434 0.754
R16049 vdd1.n434 vdd1.n433 0.754
R16050 vdd1.n454 vdd1.n453 0.754
R16051 vdd1.n453 vdd1.n452 0.754
R16052 vdd1.n452 vdd1.n451 0.754
R16053 vdd1.n451 vdd1.n450 0.754
R16054 vdd1.n449 vdd1.n448 0.754
R16055 vdd1.n448 vdd1.n447 0.754
R16056 vdd1.n447 vdd1.n446 0.754
R16057 vdd1.n446 vdd1.n445 0.754
R16058 vdd1.n466 vdd1.n465 0.754
R16059 vdd1.n465 vdd1.n464 0.754
R16060 vdd1.n464 vdd1.n463 0.754
R16061 vdd1.n463 vdd1.n462 0.754
R16062 vdd1.n461 vdd1.n460 0.754
R16063 vdd1.n460 vdd1.n459 0.754
R16064 vdd1.n459 vdd1.n458 0.754
R16065 vdd1.n458 vdd1.n457 0.754
R16066 vdd1.n477 vdd1.n476 0.754
R16067 vdd1.n476 vdd1.n475 0.754
R16068 vdd1.n475 vdd1.n474 0.754
R16069 vdd1.n474 vdd1.n473 0.754
R16070 vdd1.n472 vdd1.n471 0.754
R16071 vdd1.n471 vdd1.n470 0.754
R16072 vdd1.n470 vdd1.n469 0.754
R16073 vdd1.n469 vdd1.n468 0.754
R16074 vdd1.n488 vdd1.n487 0.754
R16075 vdd1.n487 vdd1.n486 0.754
R16076 vdd1.n486 vdd1.n485 0.754
R16077 vdd1.n485 vdd1.n484 0.754
R16078 vdd1.n483 vdd1.n482 0.754
R16079 vdd1.n482 vdd1.n481 0.754
R16080 vdd1.n481 vdd1.n480 0.754
R16081 vdd1.n480 vdd1.n479 0.754
R16082 vdd1.n9 vdd1.n8 0.754
R16083 vdd1.n8 vdd1.n7 0.754
R16084 vdd1.n7 vdd1.n6 0.754
R16085 vdd1.n6 vdd1.n5 0.754
R16086 vdd1.n4 vdd1.n3 0.754
R16087 vdd1.n3 vdd1.n2 0.754
R16088 vdd1.n2 vdd1.n1 0.754
R16089 vdd1.n1 vdd1.n0 0.754
R16090 vdd1.n42 vdd1.n41 0.726
R16091 vdd1.n39 vdd1.n38 0.58
R16092 vdd1.n40 vdd1.n39 0.58
R16093 vdd1.n41 vdd1.n40 0.58
R16094 vdd1.n43 vdd1.n42 0.58
R16095 vdd1.n44 vdd1.n43 0.58
R16096 vdd1.n45 vdd1.n44 0.58
R16097 vdd1.n46 vdd1.n45 0.58
R16098 vdd1.n57 vdd1.n46 0.516
R16099 vdd1.n68 vdd1.n67 0.427
R16100 vdd1.n79 vdd1.n78 0.427
R16101 vdd1.n90 vdd1.n89 0.427
R16102 vdd1.n101 vdd1.n100 0.427
R16103 vdd1.n112 vdd1.n111 0.427
R16104 vdd1.n123 vdd1.n122 0.427
R16105 vdd1.n134 vdd1.n133 0.427
R16106 vdd1.n145 vdd1.n144 0.427
R16107 vdd1.n156 vdd1.n155 0.427
R16108 vdd1.n167 vdd1.n166 0.427
R16109 vdd1.n178 vdd1.n177 0.427
R16110 vdd1.n189 vdd1.n188 0.427
R16111 vdd1.n200 vdd1.n199 0.427
R16112 vdd1.n211 vdd1.n210 0.427
R16113 vdd1.n222 vdd1.n221 0.427
R16114 vdd1.n233 vdd1.n232 0.427
R16115 vdd1.n244 vdd1.n243 0.427
R16116 vdd1.n255 vdd1.n254 0.427
R16117 vdd1.n266 vdd1.n265 0.427
R16118 vdd1.n277 vdd1.n276 0.427
R16119 vdd1.n288 vdd1.n287 0.427
R16120 vdd1.n299 vdd1.n298 0.427
R16121 vdd1.n310 vdd1.n309 0.427
R16122 vdd1.n321 vdd1.n320 0.427
R16123 vdd1.n333 vdd1.n332 0.427
R16124 vdd1.n344 vdd1.n343 0.427
R16125 vdd1.n355 vdd1.n354 0.427
R16126 vdd1.n366 vdd1.n365 0.427
R16127 vdd1.n377 vdd1.n376 0.427
R16128 vdd1.n388 vdd1.n387 0.427
R16129 vdd1.n399 vdd1.n398 0.427
R16130 vdd1.n410 vdd1.n409 0.427
R16131 vdd1.n421 vdd1.n420 0.427
R16132 vdd1.n432 vdd1.n431 0.427
R16133 vdd1.n443 vdd1.n442 0.427
R16134 vdd1.n467 vdd1.n466 0.427
R16135 vdd1.n478 vdd1.n477 0.427
R16136 vdd1.n489 vdd1.n488 0.427
R16137 vdd1.n57 vdd1.n56 0.427
R16138 vdd1.n455 vdd1.n454 0.427
R16139 vdd1.n943 vdd1.n942 0.426
R16140 vdd1.n931 vdd1.n930 0.426
R16141 vdd1.n915 vdd1.n914 0.426
R16142 vdd1.n903 vdd1.n902 0.426
R16143 vdd1.n887 vdd1.n886 0.426
R16144 vdd1.n875 vdd1.n874 0.426
R16145 vdd1.n859 vdd1.n858 0.426
R16146 vdd1.n847 vdd1.n846 0.426
R16147 vdd1.n831 vdd1.n830 0.426
R16148 vdd1.n819 vdd1.n818 0.426
R16149 vdd1.n803 vdd1.n802 0.426
R16150 vdd1.n791 vdd1.n790 0.426
R16151 vdd1.n775 vdd1.n774 0.426
R16152 vdd1.n763 vdd1.n762 0.426
R16153 vdd1.n747 vdd1.n746 0.426
R16154 vdd1.n735 vdd1.n734 0.426
R16155 vdd1.n719 vdd1.n718 0.426
R16156 vdd1.n707 vdd1.n706 0.426
R16157 vdd1.n691 vdd1.n690 0.426
R16158 vdd1.n679 vdd1.n678 0.426
R16159 vdd1.n663 vdd1.n662 0.426
R16160 vdd1.n651 vdd1.n650 0.426
R16161 vdd1.n635 vdd1.n634 0.426
R16162 vdd1.n623 vdd1.n622 0.426
R16163 vdd1.n607 vdd1.n606 0.426
R16164 vdd1.n595 vdd1.n594 0.426
R16165 vdd1.n579 vdd1.n578 0.426
R16166 vdd1.n567 vdd1.n566 0.426
R16167 vdd1.n551 vdd1.n550 0.426
R16168 vdd1.n539 vdd1.n538 0.426
R16169 vdd1.n523 vdd1.n522 0.426
R16170 vdd1.n511 vdd1.n510 0.426
R16171 vdd1.n37 vdd1.n36 0.426
R16172 vdd1.n10 vdd1.n9 0.426
R16173 vdd1 vdd1.n26 0.224
R16174 vdd1.n37 vdd1.n26 0.16
R16175 vdd1.n949 vdd1.n948 0.094
R16176 vdd1.n945 vdd1.n944 0.094
R16177 vdd1.n920 vdd1.n919 0.094
R16178 vdd1.n917 vdd1.n916 0.094
R16179 vdd1.n892 vdd1.n891 0.094
R16180 vdd1.n889 vdd1.n888 0.094
R16181 vdd1.n864 vdd1.n863 0.094
R16182 vdd1.n861 vdd1.n860 0.094
R16183 vdd1.n836 vdd1.n835 0.094
R16184 vdd1.n833 vdd1.n832 0.094
R16185 vdd1.n808 vdd1.n807 0.094
R16186 vdd1.n805 vdd1.n804 0.094
R16187 vdd1.n780 vdd1.n779 0.094
R16188 vdd1.n777 vdd1.n776 0.094
R16189 vdd1.n752 vdd1.n751 0.094
R16190 vdd1.n749 vdd1.n748 0.094
R16191 vdd1.n724 vdd1.n723 0.094
R16192 vdd1.n721 vdd1.n720 0.094
R16193 vdd1.n696 vdd1.n695 0.094
R16194 vdd1.n693 vdd1.n692 0.094
R16195 vdd1.n668 vdd1.n667 0.094
R16196 vdd1.n665 vdd1.n664 0.094
R16197 vdd1.n640 vdd1.n639 0.094
R16198 vdd1.n637 vdd1.n636 0.094
R16199 vdd1.n612 vdd1.n611 0.094
R16200 vdd1.n609 vdd1.n608 0.094
R16201 vdd1.n584 vdd1.n583 0.094
R16202 vdd1.n581 vdd1.n580 0.094
R16203 vdd1.n556 vdd1.n555 0.094
R16204 vdd1.n553 vdd1.n552 0.094
R16205 vdd1.n528 vdd1.n527 0.094
R16206 vdd1.n525 vdd1.n524 0.094
R16207 vdd1.n322 vdd1.n26 0.094
R16208 vdd1.n490 vdd1.n11 0.094
R16209 vdd1.n444 vdd1.n25 0.093
R16210 vdd1.n68 vdd1.n57 0.004
R16211 vdd1.n90 vdd1.n79 0.004
R16212 vdd1.n112 vdd1.n101 0.004
R16213 vdd1.n134 vdd1.n123 0.004
R16214 vdd1.n156 vdd1.n145 0.004
R16215 vdd1.n178 vdd1.n167 0.004
R16216 vdd1.n200 vdd1.n189 0.004
R16217 vdd1.n222 vdd1.n211 0.004
R16218 vdd1.n244 vdd1.n233 0.004
R16219 vdd1.n266 vdd1.n255 0.004
R16220 vdd1.n288 vdd1.n277 0.004
R16221 vdd1.n310 vdd1.n299 0.004
R16222 vdd1.n344 vdd1.n333 0.004
R16223 vdd1.n366 vdd1.n355 0.004
R16224 vdd1.n388 vdd1.n377 0.004
R16225 vdd1.n410 vdd1.n399 0.004
R16226 vdd1.n432 vdd1.n421 0.004
R16227 vdd1.n478 vdd1.n467 0.004
R16228 vdd1.n79 vdd1.n68 0.004
R16229 vdd1.n101 vdd1.n90 0.004
R16230 vdd1.n123 vdd1.n112 0.004
R16231 vdd1.n145 vdd1.n134 0.004
R16232 vdd1.n167 vdd1.n156 0.004
R16233 vdd1.n189 vdd1.n178 0.004
R16234 vdd1.n211 vdd1.n200 0.004
R16235 vdd1.n233 vdd1.n222 0.004
R16236 vdd1.n255 vdd1.n244 0.004
R16237 vdd1.n277 vdd1.n266 0.004
R16238 vdd1.n299 vdd1.n288 0.004
R16239 vdd1.n321 vdd1.n310 0.004
R16240 vdd1.n355 vdd1.n344 0.004
R16241 vdd1.n377 vdd1.n366 0.004
R16242 vdd1.n399 vdd1.n388 0.004
R16243 vdd1.n421 vdd1.n410 0.004
R16244 vdd1.n443 vdd1.n432 0.004
R16245 vdd1.n489 vdd1.n478 0.004
R16246 vdd1.n333 vdd1 0.003
R16247 vdd1.n467 vdd1.n456 0.003
R16248 vdd1 vdd1.n322 0.002
R16249 vdd1.n456 vdd1.n444 0.002
R16250 vdd1.n947 vdd1.n490 0.002
R16251 vdd1.n947 vdd1.n946 0.002
R16252 vdd1.n946 vdd1.n932 0.002
R16253 vdd1.n932 vdd1.n918 0.002
R16254 vdd1.n918 vdd1.n904 0.002
R16255 vdd1.n904 vdd1.n890 0.002
R16256 vdd1.n890 vdd1.n876 0.002
R16257 vdd1.n876 vdd1.n862 0.002
R16258 vdd1.n862 vdd1.n848 0.002
R16259 vdd1.n848 vdd1.n834 0.002
R16260 vdd1.n834 vdd1.n820 0.002
R16261 vdd1.n820 vdd1.n806 0.002
R16262 vdd1.n806 vdd1.n792 0.002
R16263 vdd1.n792 vdd1.n778 0.002
R16264 vdd1.n778 vdd1.n764 0.002
R16265 vdd1.n764 vdd1.n750 0.002
R16266 vdd1.n750 vdd1.n736 0.002
R16267 vdd1.n736 vdd1.n722 0.002
R16268 vdd1.n722 vdd1.n708 0.002
R16269 vdd1.n708 vdd1.n694 0.002
R16270 vdd1.n694 vdd1.n680 0.002
R16271 vdd1.n680 vdd1.n666 0.002
R16272 vdd1.n666 vdd1.n652 0.002
R16273 vdd1.n652 vdd1.n638 0.002
R16274 vdd1.n638 vdd1.n624 0.002
R16275 vdd1.n624 vdd1.n610 0.002
R16276 vdd1.n610 vdd1.n596 0.002
R16277 vdd1.n596 vdd1.n582 0.002
R16278 vdd1.n582 vdd1.n568 0.002
R16279 vdd1.n568 vdd1.n554 0.002
R16280 vdd1.n554 vdd1.n540 0.002
R16281 vdd1.n540 vdd1.n526 0.002
R16282 vdd1.n526 vdd1.n512 0.002
R16283 vdd1.n456 vdd1.n455 0.001
R16284 vdd1.n946 vdd1.n943 0.001
R16285 vdd1.n932 vdd1.n931 0.001
R16286 vdd1.n918 vdd1.n915 0.001
R16287 vdd1.n904 vdd1.n903 0.001
R16288 vdd1.n890 vdd1.n887 0.001
R16289 vdd1.n876 vdd1.n875 0.001
R16290 vdd1.n862 vdd1.n859 0.001
R16291 vdd1.n848 vdd1.n847 0.001
R16292 vdd1.n834 vdd1.n831 0.001
R16293 vdd1.n820 vdd1.n819 0.001
R16294 vdd1.n806 vdd1.n803 0.001
R16295 vdd1.n792 vdd1.n791 0.001
R16296 vdd1.n778 vdd1.n775 0.001
R16297 vdd1.n764 vdd1.n763 0.001
R16298 vdd1.n750 vdd1.n747 0.001
R16299 vdd1.n736 vdd1.n735 0.001
R16300 vdd1.n722 vdd1.n719 0.001
R16301 vdd1.n708 vdd1.n707 0.001
R16302 vdd1.n694 vdd1.n691 0.001
R16303 vdd1.n680 vdd1.n679 0.001
R16304 vdd1.n666 vdd1.n663 0.001
R16305 vdd1.n652 vdd1.n651 0.001
R16306 vdd1.n638 vdd1.n635 0.001
R16307 vdd1.n624 vdd1.n623 0.001
R16308 vdd1.n610 vdd1.n607 0.001
R16309 vdd1.n596 vdd1.n595 0.001
R16310 vdd1.n582 vdd1.n579 0.001
R16311 vdd1.n568 vdd1.n567 0.001
R16312 vdd1.n554 vdd1.n551 0.001
R16313 vdd1.n540 vdd1.n539 0.001
R16314 vdd1.n526 vdd1.n523 0.001
R16315 vdd1.n512 vdd1.n511 0.001
R16316 vdd1 vdd1.n37 0.001
R16317 vdd1.n947 vdd1.n10 0.001
R16318 vdd1.n25 vdd1.n24 0.001
R16319 vdd1.n512 vdd1.n500 0.001
R16320 vdd1.n322 vdd1.n321 0.001
R16321 vdd1.n444 vdd1.n443 0.001
R16322 vdd1.n490 vdd1.n489 0.001
R16323 vdd1.n526 vdd1.n525 0.001
R16324 vdd1.n540 vdd1.n528 0.001
R16325 vdd1.n554 vdd1.n553 0.001
R16326 vdd1.n568 vdd1.n556 0.001
R16327 vdd1.n582 vdd1.n581 0.001
R16328 vdd1.n596 vdd1.n584 0.001
R16329 vdd1.n610 vdd1.n609 0.001
R16330 vdd1.n624 vdd1.n612 0.001
R16331 vdd1.n638 vdd1.n637 0.001
R16332 vdd1.n652 vdd1.n640 0.001
R16333 vdd1.n666 vdd1.n665 0.001
R16334 vdd1.n680 vdd1.n668 0.001
R16335 vdd1.n694 vdd1.n693 0.001
R16336 vdd1.n708 vdd1.n696 0.001
R16337 vdd1.n722 vdd1.n721 0.001
R16338 vdd1.n736 vdd1.n724 0.001
R16339 vdd1.n750 vdd1.n749 0.001
R16340 vdd1.n764 vdd1.n752 0.001
R16341 vdd1.n778 vdd1.n777 0.001
R16342 vdd1.n792 vdd1.n780 0.001
R16343 vdd1.n806 vdd1.n805 0.001
R16344 vdd1.n820 vdd1.n808 0.001
R16345 vdd1.n834 vdd1.n833 0.001
R16346 vdd1.n848 vdd1.n836 0.001
R16347 vdd1.n862 vdd1.n861 0.001
R16348 vdd1.n876 vdd1.n864 0.001
R16349 vdd1.n890 vdd1.n889 0.001
R16350 vdd1.n904 vdd1.n892 0.001
R16351 vdd1.n918 vdd1.n917 0.001
R16352 vdd1.n932 vdd1.n920 0.001
R16353 vdd1.n946 vdd1.n945 0.001
R16354 vdd1.n949 vdd1.n947 0.001
R16355 vp_n.n221 vp_n.t280 721.861
R16356 vp_n.n219 vp_n.t27 721.861
R16357 vp_n.n217 vp_n.t244 721.861
R16358 vp_n.n215 vp_n.t123 721.861
R16359 vp_n.n213 vp_n.t168 721.861
R16360 vp_n.n211 vp_n.t93 721.861
R16361 vp_n.n209 vp_n.t133 721.861
R16362 vp_n.n207 vp_n.t60 721.861
R16363 vp_n.n205 vp_n.t69 721.861
R16364 vp_n.n203 vp_n.t291 721.861
R16365 vp_n.n201 vp_n.t203 721.861
R16366 vp_n.n199 vp_n.t254 721.861
R16367 vp_n.n197 vp_n.t167 721.861
R16368 vp_n.n195 vp_n.t178 721.861
R16369 vp_n.n193 vp_n.t102 721.861
R16370 vp_n.n191 vp_n.t26 721.861
R16371 vp_n.n189 vp_n.t30 721.861
R16372 vp_n.n187 vp_n.t247 721.861
R16373 vp_n.n185 vp_n.t259 721.861
R16374 vp_n.n183 vp_n.t173 721.861
R16375 vp_n.n181 vp_n.t221 721.861
R16376 vp_n.n179 vp_n.t136 721.861
R16377 vp_n.n177 vp_n.t63 721.861
R16378 vp_n.n175 vp_n.t76 721.861
R16379 vp_n.n173 vp_n.t295 721.861
R16380 vp_n.n171 vp_n.t40 721.861
R16381 vp_n.n169 vp_n.t258 721.861
R16382 vp_n.n167 vp_n.t172 721.861
R16383 vp_n.n165 vp_n.t184 721.861
R16384 vp_n.n163 vp_n.t106 721.861
R16385 vp_n.n161 vp_n.t150 721.861
R16386 vp_n.n159 vp_n.t74 721.861
R16387 vp_n.n157 vp_n.t116 721.861
R16388 vp_n.n155 vp_n.t7 721.861
R16389 vp_n.n153 vp_n.t219 721.861
R16390 vp_n.n151 vp_n.t272 721.861
R16391 vp_n.n149 vp_n.t182 721.861
R16392 vp_n.n147 vp_n.t234 721.861
R16393 vp_n.n145 vp_n.t117 721.861
R16394 vp_n.n143 vp_n.t49 721.861
R16395 vp_n.n141 vp_n.t266 721.861
R16396 vp_n.n139 vp_n.t176 721.861
R16397 vp_n.n137 vp_n.t227 721.861
R16398 vp_n.n135 vp_n.t110 721.861
R16399 vp_n.n133 vp_n.t158 721.861
R16400 vp_n.n131 vp_n.t82 721.861
R16401 vp_n.n129 vp_n.t0 721.861
R16402 vp_n.n127 vp_n.t47 721.861
R16403 vp_n.n125 vp_n.t228 721.861
R16404 vp_n.n123 vp_n.t279 721.861
R16405 vp_n.n121 vp_n.t188 721.861
R16406 vp_n.n119 vp_n.t242 721.861
R16407 vp_n.n117 vp_n.t156 721.861
R16408 vp_n.n115 vp_n.t48 721.861
R16409 vp_n.n113 vp_n.t92 721.861
R16410 vp_n.n111 vp_n.t12 721.861
R16411 vp_n.n109 vp_n.t58 721.861
R16412 vp_n.n107 vp_n.t277 721.861
R16413 vp_n.n105 vp_n.t290 721.861
R16414 vp_n.n103 vp_n.t201 721.861
R16415 vp_n.n101 vp_n.t121 721.861
R16416 vp_n.n99 vp_n.t165 721.861
R16417 vp_n.n97 vp_n.t91 721.861
R16418 vp_n.n95 vp_n.t284 721.861
R16419 vp_n.n93 vp_n.t196 721.861
R16420 vp_n.n91 vp_n.t115 721.861
R16421 vp_n.n89 vp_n.t162 721.861
R16422 vp_n.n87 vp_n.t86 721.861
R16423 vp_n.n85 vp_n.t96 721.861
R16424 vp_n.n83 vp_n.t19 721.861
R16425 vp_n.n81 vp_n.t64 721.861
R16426 vp_n.n79 vp_n.t283 721.861
R16427 vp_n.n77 vp_n.t194 721.861
R16428 vp_n.n75 vp_n.t208 721.861
R16429 vp_n.n74 vp_n.t127 721.861
R16430 vp_n.n221 vp_n.t5 721.861
R16431 vp_n.n219 vp_n.t52 721.861
R16432 vp_n.n217 vp_n.t270 721.861
R16433 vp_n.n215 vp_n.t148 721.861
R16434 vp_n.n213 vp_n.t193 721.861
R16435 vp_n.n211 vp_n.t113 721.861
R16436 vp_n.n209 vp_n.t160 721.861
R16437 vp_n.n207 vp_n.t85 721.861
R16438 vp_n.n205 vp_n.t95 721.861
R16439 vp_n.n203 vp_n.t17 721.861
R16440 vp_n.n201 vp_n.t232 721.861
R16441 vp_n.n199 vp_n.t282 721.861
R16442 vp_n.n197 vp_n.t192 721.861
R16443 vp_n.n195 vp_n.t206 721.861
R16444 vp_n.n193 vp_n.t125 721.861
R16445 vp_n.n191 vp_n.t51 721.861
R16446 vp_n.n189 vp_n.t56 721.861
R16447 vp_n.n187 vp_n.t274 721.861
R16448 vp_n.n185 vp_n.t287 721.861
R16449 vp_n.n183 vp_n.t199 721.861
R16450 vp_n.n181 vp_n.t252 721.861
R16451 vp_n.n179 vp_n.t163 721.861
R16452 vp_n.n177 vp_n.t88 721.861
R16453 vp_n.n175 vp_n.t100 721.861
R16454 vp_n.n173 vp_n.t23 721.861
R16455 vp_n.n171 vp_n.t67 721.861
R16456 vp_n.n169 vp_n.t286 721.861
R16457 vp_n.n167 vp_n.t198 721.861
R16458 vp_n.n165 vp_n.t213 721.861
R16459 vp_n.n163 vp_n.t131 721.861
R16460 vp_n.n161 vp_n.t175 721.861
R16461 vp_n.n159 vp_n.t98 721.861
R16462 vp_n.n157 vp_n.t140 721.861
R16463 vp_n.n155 vp_n.t33 721.861
R16464 vp_n.n153 vp_n.t250 721.861
R16465 vp_n.n151 vp_n.t298 721.861
R16466 vp_n.n149 vp_n.t211 721.861
R16467 vp_n.n147 vp_n.t261 721.861
R16468 vp_n.n145 vp_n.t141 721.861
R16469 vp_n.n143 vp_n.t73 721.861
R16470 vp_n.n141 vp_n.t294 721.861
R16471 vp_n.n139 vp_n.t204 721.861
R16472 vp_n.n137 vp_n.t256 721.861
R16473 vp_n.n135 vp_n.t135 721.861
R16474 vp_n.n133 vp_n.t181 721.861
R16475 vp_n.n131 vp_n.t105 721.861
R16476 vp_n.n129 vp_n.t28 721.861
R16477 vp_n.n127 vp_n.t71 721.861
R16478 vp_n.n125 vp_n.t257 721.861
R16479 vp_n.n123 vp_n.t4 721.861
R16480 vp_n.n121 vp_n.t217 721.861
R16481 vp_n.n119 vp_n.t268 721.861
R16482 vp_n.n117 vp_n.t179 721.861
R16483 vp_n.n115 vp_n.t72 721.861
R16484 vp_n.n113 vp_n.t112 721.861
R16485 vp_n.n111 vp_n.t37 721.861
R16486 vp_n.n109 vp_n.t83 721.861
R16487 vp_n.n107 vp_n.t2 721.861
R16488 vp_n.n105 vp_n.t16 721.861
R16489 vp_n.n103 vp_n.t230 721.861
R16490 vp_n.n101 vp_n.t146 721.861
R16491 vp_n.n99 vp_n.t190 721.861
R16492 vp_n.n97 vp_n.t111 721.861
R16493 vp_n.n95 vp_n.t10 721.861
R16494 vp_n.n93 vp_n.t224 721.861
R16495 vp_n.n91 vp_n.t139 721.861
R16496 vp_n.n89 vp_n.t186 721.861
R16497 vp_n.n87 vp_n.t107 721.861
R16498 vp_n.n85 vp_n.t119 721.861
R16499 vp_n.n83 vp_n.t42 721.861
R16500 vp_n.n81 vp_n.t89 721.861
R16501 vp_n.n79 vp_n.t9 721.861
R16502 vp_n.n77 vp_n.t222 721.861
R16503 vp_n.n75 vp_n.t238 721.861
R16504 vp_n.n74 vp_n.t152 721.861
R16505 vp_n.n0 vp_n.t166 691.553
R16506 vp_n.n223 vp_n.t191 691.553
R16507 vp_n.n73 vp_n.t22 690.412
R16508 vp_n.n72 vp_n.t236 690.412
R16509 vp_n.n71 vp_n.t285 690.412
R16510 vp_n.n70 vp_n.t197 690.412
R16511 vp_n.n69 vp_n.t210 690.412
R16512 vp_n.n68 vp_n.t130 690.412
R16513 vp_n.n67 vp_n.t55 690.412
R16514 vp_n.n66 vp_n.t97 690.412
R16515 vp_n.n65 vp_n.t20 690.412
R16516 vp_n.n64 vp_n.t31 690.412
R16517 vp_n.n63 vp_n.t249 690.412
R16518 vp_n.n62 vp_n.t296 690.412
R16519 vp_n.n61 vp_n.t209 690.412
R16520 vp_n.n60 vp_n.t128 690.412
R16521 vp_n.n59 vp_n.t137 690.412
R16522 vp_n.n58 vp_n.t65 690.412
R16523 vp_n.n57 vp_n.t68 690.412
R16524 vp_n.n56 vp_n.t288 690.412
R16525 vp_n.n55 vp_n.t200 690.412
R16526 vp_n.n54 vp_n.t215 690.412
R16527 vp_n.n53 vp_n.t132 690.412
R16528 vp_n.n52 vp_n.t177 690.412
R16529 vp_n.n51 vp_n.t101 690.412
R16530 vp_n.n50 vp_n.t144 690.412
R16531 vp_n.n49 vp_n.t36 690.412
R16532 vp_n.n48 vp_n.t253 690.412
R16533 vp_n.n47 vp_n.t1 690.412
R16534 vp_n.n46 vp_n.t214 690.412
R16535 vp_n.n45 vp_n.t264 690.412
R16536 vp_n.n44 vp_n.t145 690.412
R16537 vp_n.n43 vp_n.t189 690.412
R16538 vp_n.n42 vp_n.t109 690.412
R16539 vp_n.n41 vp_n.t35 690.412
R16540 vp_n.n40 vp_n.t80 690.412
R16541 vp_n.n39 vp_n.t265 690.412
R16542 vp_n.n38 vp_n.t13 690.412
R16543 vp_n.n37 vp_n.t226 690.412
R16544 vp_n.n36 vp_n.t143 690.412
R16545 vp_n.n35 vp_n.t187 690.412
R16546 vp_n.n34 vp_n.t81 690.412
R16547 vp_n.n33 vp_n.t8 690.412
R16548 vp_n.n32 vp_n.t220 690.412
R16549 vp_n.n31 vp_n.t273 690.412
R16550 vp_n.n30 vp_n.t183 690.412
R16551 vp_n.n29 vp_n.t75 690.412
R16552 vp_n.n28 vp_n.t118 690.412
R16553 vp_n.n27 vp_n.t39 690.412
R16554 vp_n.n26 vp_n.t87 690.412
R16555 vp_n.n25 vp_n.t6 690.412
R16556 vp_n.n24 vp_n.t21 690.412
R16557 vp_n.n23 vp_n.t235 690.412
R16558 vp_n.n22 vp_n.t149 690.412
R16559 vp_n.n21 vp_n.t195 690.412
R16560 vp_n.n20 vp_n.t114 690.412
R16561 vp_n.n19 vp_n.t129 690.412
R16562 vp_n.n18 vp_n.t54 690.412
R16563 vp_n.n17 vp_n.t271 690.412
R16564 vp_n.n16 vp_n.t18 690.412
R16565 vp_n.n15 vp_n.t233 690.412
R16566 vp_n.n14 vp_n.t248 690.412
R16567 vp_n.n13 vp_n.t161 690.412
R16568 vp_n.n12 vp_n.t207 690.412
R16569 vp_n.n11 vp_n.t126 690.412
R16570 vp_n.n10 vp_n.t53 690.412
R16571 vp_n.n9 vp_n.t243 690.412
R16572 vp_n.n8 vp_n.t157 690.412
R16573 vp_n.n7 vp_n.t202 690.412
R16574 vp_n.n6 vp_n.t122 690.412
R16575 vp_n.n5 vp_n.t46 690.412
R16576 vp_n.n4 vp_n.t59 690.412
R16577 vp_n.n3 vp_n.t278 690.412
R16578 vp_n.n2 vp_n.t25 690.412
R16579 vp_n.n1 vp_n.t241 690.412
R16580 vp_n.n0 vp_n.t289 690.412
R16581 vp_n.n223 vp_n.t15 690.412
R16582 vp_n.n224 vp_n.t267 690.412
R16583 vp_n.n225 vp_n.t50 690.412
R16584 vp_n.n226 vp_n.t3 690.412
R16585 vp_n.n227 vp_n.t84 690.412
R16586 vp_n.n228 vp_n.t70 690.412
R16587 vp_n.n229 vp_n.t147 690.412
R16588 vp_n.n230 vp_n.t231 690.412
R16589 vp_n.n231 vp_n.t180 690.412
R16590 vp_n.n232 vp_n.t269 690.412
R16591 vp_n.n233 vp_n.t77 690.412
R16592 vp_n.n234 vp_n.t151 690.412
R16593 vp_n.n235 vp_n.t237 690.412
R16594 vp_n.n236 vp_n.t185 690.412
R16595 vp_n.n237 vp_n.t275 690.412
R16596 vp_n.n238 vp_n.t260 690.412
R16597 vp_n.n239 vp_n.t41 690.412
R16598 vp_n.n240 vp_n.t297 690.412
R16599 vp_n.n241 vp_n.t78 690.412
R16600 vp_n.n242 vp_n.t154 690.412
R16601 vp_n.n243 vp_n.t138 690.412
R16602 vp_n.n244 vp_n.t223 690.412
R16603 vp_n.n245 vp_n.t174 690.412
R16604 vp_n.n246 vp_n.t262 690.412
R16605 vp_n.n247 vp_n.t44 690.412
R16606 vp_n.n248 vp_n.t32 690.412
R16607 vp_n.n249 vp_n.t108 690.412
R16608 vp_n.n250 vp_n.t66 690.412
R16609 vp_n.n251 vp_n.t142 690.412
R16610 vp_n.n252 vp_n.t99 690.412
R16611 vp_n.n253 vp_n.t212 690.412
R16612 vp_n.n254 vp_n.t299 690.412
R16613 vp_n.n255 vp_n.t251 690.412
R16614 vp_n.n256 vp_n.t34 690.412
R16615 vp_n.n257 vp_n.t104 690.412
R16616 vp_n.n258 vp_n.t216 690.412
R16617 vp_n.n259 vp_n.t169 690.412
R16618 vp_n.n260 vp_n.t255 690.412
R16619 vp_n.n261 vp_n.t38 690.412
R16620 vp_n.n262 vp_n.t293 690.412
R16621 vp_n.n263 vp_n.t103 690.412
R16622 vp_n.n264 vp_n.t61 690.412
R16623 vp_n.n265 vp_n.t134 690.412
R16624 vp_n.n266 vp_n.t218 690.412
R16625 vp_n.n267 vp_n.t171 690.412
R16626 vp_n.n268 vp_n.t292 690.412
R16627 vp_n.n269 vp_n.t245 690.412
R16628 vp_n.n270 vp_n.t29 690.412
R16629 vp_n.n271 vp_n.t281 690.412
R16630 vp_n.n272 vp_n.t62 690.412
R16631 vp_n.n273 vp_n.t170 690.412
R16632 vp_n.n274 vp_n.t124 690.412
R16633 vp_n.n275 vp_n.t205 690.412
R16634 vp_n.n276 vp_n.t159 690.412
R16635 vp_n.n277 vp_n.t246 690.412
R16636 vp_n.n278 vp_n.t229 690.412
R16637 vp_n.n279 vp_n.t14 690.412
R16638 vp_n.n280 vp_n.t94 690.412
R16639 vp_n.n281 vp_n.t90 690.412
R16640 vp_n.n282 vp_n.t164 690.412
R16641 vp_n.n283 vp_n.t153 690.412
R16642 vp_n.n284 vp_n.t239 690.412
R16643 vp_n.n285 vp_n.t24 690.412
R16644 vp_n.n286 vp_n.t276 690.412
R16645 vp_n.n287 vp_n.t57 690.412
R16646 vp_n.n288 vp_n.t43 690.412
R16647 vp_n.n289 vp_n.t120 690.412
R16648 vp_n.n290 vp_n.t79 690.412
R16649 vp_n.n291 vp_n.t155 690.412
R16650 vp_n.n292 vp_n.t240 690.412
R16651 vp_n.n293 vp_n.t225 690.412
R16652 vp_n.n294 vp_n.t11 690.412
R16653 vp_n.n295 vp_n.t263 690.412
R16654 vp_n.n296 vp_n.t45 690.412
R16655 vp_n.n76 vp_n.n74 6.382
R16656 vp_n.n76 vp_n.n75 6.013
R16657 vp_n.n78 vp_n.n77 6.013
R16658 vp_n.n80 vp_n.n79 6.013
R16659 vp_n.n82 vp_n.n81 6.013
R16660 vp_n.n84 vp_n.n83 6.013
R16661 vp_n.n86 vp_n.n85 6.013
R16662 vp_n.n88 vp_n.n87 6.013
R16663 vp_n.n90 vp_n.n89 6.013
R16664 vp_n.n92 vp_n.n91 6.013
R16665 vp_n.n94 vp_n.n93 6.013
R16666 vp_n.n96 vp_n.n95 6.013
R16667 vp_n.n98 vp_n.n97 6.013
R16668 vp_n.n100 vp_n.n99 6.013
R16669 vp_n.n102 vp_n.n101 6.013
R16670 vp_n.n104 vp_n.n103 6.013
R16671 vp_n.n106 vp_n.n105 6.013
R16672 vp_n.n108 vp_n.n107 6.013
R16673 vp_n.n110 vp_n.n109 6.013
R16674 vp_n.n112 vp_n.n111 6.013
R16675 vp_n.n114 vp_n.n113 6.013
R16676 vp_n.n116 vp_n.n115 6.013
R16677 vp_n.n118 vp_n.n117 6.013
R16678 vp_n.n120 vp_n.n119 6.013
R16679 vp_n.n122 vp_n.n121 6.013
R16680 vp_n.n124 vp_n.n123 6.013
R16681 vp_n.n126 vp_n.n125 6.013
R16682 vp_n.n128 vp_n.n127 6.013
R16683 vp_n.n130 vp_n.n129 6.013
R16684 vp_n.n132 vp_n.n131 6.013
R16685 vp_n.n134 vp_n.n133 6.013
R16686 vp_n.n136 vp_n.n135 6.013
R16687 vp_n.n138 vp_n.n137 6.013
R16688 vp_n.n140 vp_n.n139 6.013
R16689 vp_n.n142 vp_n.n141 6.013
R16690 vp_n.n144 vp_n.n143 6.013
R16691 vp_n.n146 vp_n.n145 6.013
R16692 vp_n.n148 vp_n.n147 6.013
R16693 vp_n.n150 vp_n.n149 6.013
R16694 vp_n.n152 vp_n.n151 6.013
R16695 vp_n.n154 vp_n.n153 6.013
R16696 vp_n.n156 vp_n.n155 6.013
R16697 vp_n.n158 vp_n.n157 6.013
R16698 vp_n.n160 vp_n.n159 6.013
R16699 vp_n.n162 vp_n.n161 6.013
R16700 vp_n.n164 vp_n.n163 6.013
R16701 vp_n.n166 vp_n.n165 6.013
R16702 vp_n.n168 vp_n.n167 6.013
R16703 vp_n.n170 vp_n.n169 6.013
R16704 vp_n.n172 vp_n.n171 6.013
R16705 vp_n.n174 vp_n.n173 6.013
R16706 vp_n.n176 vp_n.n175 6.013
R16707 vp_n.n178 vp_n.n177 6.013
R16708 vp_n.n180 vp_n.n179 6.013
R16709 vp_n.n182 vp_n.n181 6.013
R16710 vp_n.n184 vp_n.n183 6.013
R16711 vp_n.n186 vp_n.n185 6.013
R16712 vp_n.n188 vp_n.n187 6.013
R16713 vp_n.n190 vp_n.n189 6.013
R16714 vp_n.n192 vp_n.n191 6.013
R16715 vp_n.n194 vp_n.n193 6.013
R16716 vp_n.n196 vp_n.n195 6.013
R16717 vp_n.n198 vp_n.n197 6.013
R16718 vp_n.n200 vp_n.n199 6.013
R16719 vp_n.n202 vp_n.n201 6.013
R16720 vp_n.n204 vp_n.n203 6.013
R16721 vp_n.n206 vp_n.n205 6.013
R16722 vp_n.n208 vp_n.n207 6.013
R16723 vp_n.n210 vp_n.n209 6.013
R16724 vp_n.n212 vp_n.n211 6.013
R16725 vp_n.n214 vp_n.n213 6.013
R16726 vp_n.n216 vp_n.n215 6.013
R16727 vp_n.n218 vp_n.n217 6.013
R16728 vp_n.n220 vp_n.n219 6.013
R16729 vp_n.n222 vp_n.n221 6.013
R16730 vp_n.n1 vp_n.n0 1.141
R16731 vp_n.n2 vp_n.n1 1.141
R16732 vp_n.n3 vp_n.n2 1.141
R16733 vp_n.n4 vp_n.n3 1.141
R16734 vp_n.n5 vp_n.n4 1.141
R16735 vp_n.n6 vp_n.n5 1.141
R16736 vp_n.n7 vp_n.n6 1.141
R16737 vp_n.n8 vp_n.n7 1.141
R16738 vp_n.n9 vp_n.n8 1.141
R16739 vp_n.n10 vp_n.n9 1.141
R16740 vp_n.n11 vp_n.n10 1.141
R16741 vp_n.n12 vp_n.n11 1.141
R16742 vp_n.n13 vp_n.n12 1.141
R16743 vp_n.n14 vp_n.n13 1.141
R16744 vp_n.n15 vp_n.n14 1.141
R16745 vp_n.n16 vp_n.n15 1.141
R16746 vp_n.n17 vp_n.n16 1.141
R16747 vp_n.n18 vp_n.n17 1.141
R16748 vp_n.n19 vp_n.n18 1.141
R16749 vp_n.n20 vp_n.n19 1.141
R16750 vp_n.n21 vp_n.n20 1.141
R16751 vp_n.n22 vp_n.n21 1.141
R16752 vp_n.n23 vp_n.n22 1.141
R16753 vp_n.n24 vp_n.n23 1.141
R16754 vp_n.n25 vp_n.n24 1.141
R16755 vp_n.n26 vp_n.n25 1.141
R16756 vp_n.n27 vp_n.n26 1.141
R16757 vp_n.n28 vp_n.n27 1.141
R16758 vp_n.n29 vp_n.n28 1.141
R16759 vp_n.n30 vp_n.n29 1.141
R16760 vp_n.n31 vp_n.n30 1.141
R16761 vp_n.n32 vp_n.n31 1.141
R16762 vp_n.n33 vp_n.n32 1.141
R16763 vp_n.n34 vp_n.n33 1.141
R16764 vp_n.n35 vp_n.n34 1.141
R16765 vp_n.n36 vp_n.n35 1.141
R16766 vp_n.n37 vp_n.n36 1.141
R16767 vp_n.n38 vp_n.n37 1.141
R16768 vp_n.n39 vp_n.n38 1.141
R16769 vp_n.n40 vp_n.n39 1.141
R16770 vp_n.n41 vp_n.n40 1.141
R16771 vp_n.n42 vp_n.n41 1.141
R16772 vp_n.n43 vp_n.n42 1.141
R16773 vp_n.n44 vp_n.n43 1.141
R16774 vp_n.n45 vp_n.n44 1.141
R16775 vp_n.n46 vp_n.n45 1.141
R16776 vp_n.n47 vp_n.n46 1.141
R16777 vp_n.n48 vp_n.n47 1.141
R16778 vp_n.n49 vp_n.n48 1.141
R16779 vp_n.n50 vp_n.n49 1.141
R16780 vp_n.n51 vp_n.n50 1.141
R16781 vp_n.n52 vp_n.n51 1.141
R16782 vp_n.n53 vp_n.n52 1.141
R16783 vp_n.n54 vp_n.n53 1.141
R16784 vp_n.n55 vp_n.n54 1.141
R16785 vp_n.n56 vp_n.n55 1.141
R16786 vp_n.n57 vp_n.n56 1.141
R16787 vp_n.n58 vp_n.n57 1.141
R16788 vp_n.n59 vp_n.n58 1.141
R16789 vp_n.n60 vp_n.n59 1.141
R16790 vp_n.n61 vp_n.n60 1.141
R16791 vp_n.n62 vp_n.n61 1.141
R16792 vp_n.n63 vp_n.n62 1.141
R16793 vp_n.n64 vp_n.n63 1.141
R16794 vp_n.n65 vp_n.n64 1.141
R16795 vp_n.n66 vp_n.n65 1.141
R16796 vp_n.n67 vp_n.n66 1.141
R16797 vp_n.n68 vp_n.n67 1.141
R16798 vp_n.n69 vp_n.n68 1.141
R16799 vp_n.n70 vp_n.n69 1.141
R16800 vp_n.n71 vp_n.n70 1.141
R16801 vp_n.n72 vp_n.n71 1.141
R16802 vp_n.n73 vp_n.n72 1.141
R16803 vp_n.n224 vp_n.n223 1.141
R16804 vp_n.n225 vp_n.n224 1.141
R16805 vp_n.n226 vp_n.n225 1.141
R16806 vp_n.n227 vp_n.n226 1.141
R16807 vp_n.n228 vp_n.n227 1.141
R16808 vp_n.n229 vp_n.n228 1.141
R16809 vp_n.n230 vp_n.n229 1.141
R16810 vp_n.n231 vp_n.n230 1.141
R16811 vp_n.n232 vp_n.n231 1.141
R16812 vp_n.n233 vp_n.n232 1.141
R16813 vp_n.n234 vp_n.n233 1.141
R16814 vp_n.n235 vp_n.n234 1.141
R16815 vp_n.n236 vp_n.n235 1.141
R16816 vp_n.n237 vp_n.n236 1.141
R16817 vp_n.n238 vp_n.n237 1.141
R16818 vp_n.n239 vp_n.n238 1.141
R16819 vp_n.n240 vp_n.n239 1.141
R16820 vp_n.n241 vp_n.n240 1.141
R16821 vp_n.n242 vp_n.n241 1.141
R16822 vp_n.n243 vp_n.n242 1.141
R16823 vp_n.n244 vp_n.n243 1.141
R16824 vp_n.n245 vp_n.n244 1.141
R16825 vp_n.n246 vp_n.n245 1.141
R16826 vp_n.n247 vp_n.n246 1.141
R16827 vp_n.n248 vp_n.n247 1.141
R16828 vp_n.n249 vp_n.n248 1.141
R16829 vp_n.n250 vp_n.n249 1.141
R16830 vp_n.n251 vp_n.n250 1.141
R16831 vp_n.n252 vp_n.n251 1.141
R16832 vp_n.n253 vp_n.n252 1.141
R16833 vp_n.n254 vp_n.n253 1.141
R16834 vp_n.n255 vp_n.n254 1.141
R16835 vp_n.n256 vp_n.n255 1.141
R16836 vp_n.n257 vp_n.n256 1.141
R16837 vp_n.n258 vp_n.n257 1.141
R16838 vp_n.n259 vp_n.n258 1.141
R16839 vp_n.n260 vp_n.n259 1.141
R16840 vp_n.n261 vp_n.n260 1.141
R16841 vp_n.n262 vp_n.n261 1.141
R16842 vp_n.n263 vp_n.n262 1.141
R16843 vp_n.n264 vp_n.n263 1.141
R16844 vp_n.n265 vp_n.n264 1.141
R16845 vp_n.n266 vp_n.n265 1.141
R16846 vp_n.n267 vp_n.n266 1.141
R16847 vp_n.n268 vp_n.n267 1.141
R16848 vp_n.n269 vp_n.n268 1.141
R16849 vp_n.n270 vp_n.n269 1.141
R16850 vp_n.n271 vp_n.n270 1.141
R16851 vp_n.n272 vp_n.n271 1.141
R16852 vp_n.n273 vp_n.n272 1.141
R16853 vp_n.n274 vp_n.n273 1.141
R16854 vp_n.n275 vp_n.n274 1.141
R16855 vp_n.n276 vp_n.n275 1.141
R16856 vp_n.n277 vp_n.n276 1.141
R16857 vp_n.n278 vp_n.n277 1.141
R16858 vp_n.n279 vp_n.n278 1.141
R16859 vp_n.n280 vp_n.n279 1.141
R16860 vp_n.n281 vp_n.n280 1.141
R16861 vp_n.n282 vp_n.n281 1.141
R16862 vp_n.n283 vp_n.n282 1.141
R16863 vp_n.n284 vp_n.n283 1.141
R16864 vp_n.n285 vp_n.n284 1.141
R16865 vp_n.n286 vp_n.n285 1.141
R16866 vp_n.n287 vp_n.n286 1.141
R16867 vp_n.n288 vp_n.n287 1.141
R16868 vp_n.n289 vp_n.n288 1.141
R16869 vp_n.n290 vp_n.n289 1.141
R16870 vp_n.n291 vp_n.n290 1.141
R16871 vp_n.n292 vp_n.n291 1.141
R16872 vp_n.n293 vp_n.n292 1.141
R16873 vp_n.n294 vp_n.n293 1.141
R16874 vp_n.n295 vp_n.n294 1.141
R16875 vp_n.n296 vp_n.n295 1.141
R16876 vp_n.n297 vp_n.n296 0.948
R16877 vp_n vp_n.n73 0.872
R16878 vp_n.n297 vp_n.n222 0.413
R16879 vp_n.n78 vp_n.n76 0.369
R16880 vp_n.n80 vp_n.n78 0.369
R16881 vp_n.n82 vp_n.n80 0.369
R16882 vp_n.n84 vp_n.n82 0.369
R16883 vp_n.n86 vp_n.n84 0.369
R16884 vp_n.n88 vp_n.n86 0.369
R16885 vp_n.n90 vp_n.n88 0.369
R16886 vp_n.n92 vp_n.n90 0.369
R16887 vp_n.n94 vp_n.n92 0.369
R16888 vp_n.n96 vp_n.n94 0.369
R16889 vp_n.n98 vp_n.n96 0.369
R16890 vp_n.n100 vp_n.n98 0.369
R16891 vp_n.n102 vp_n.n100 0.369
R16892 vp_n.n104 vp_n.n102 0.369
R16893 vp_n.n106 vp_n.n104 0.369
R16894 vp_n.n108 vp_n.n106 0.369
R16895 vp_n.n110 vp_n.n108 0.369
R16896 vp_n.n112 vp_n.n110 0.369
R16897 vp_n.n114 vp_n.n112 0.369
R16898 vp_n.n116 vp_n.n114 0.369
R16899 vp_n.n118 vp_n.n116 0.369
R16900 vp_n.n120 vp_n.n118 0.369
R16901 vp_n.n122 vp_n.n120 0.369
R16902 vp_n.n124 vp_n.n122 0.369
R16903 vp_n.n126 vp_n.n124 0.369
R16904 vp_n.n128 vp_n.n126 0.369
R16905 vp_n.n130 vp_n.n128 0.369
R16906 vp_n.n132 vp_n.n130 0.369
R16907 vp_n.n134 vp_n.n132 0.369
R16908 vp_n.n136 vp_n.n134 0.369
R16909 vp_n.n138 vp_n.n136 0.369
R16910 vp_n.n140 vp_n.n138 0.369
R16911 vp_n.n142 vp_n.n140 0.369
R16912 vp_n.n144 vp_n.n142 0.369
R16913 vp_n.n146 vp_n.n144 0.369
R16914 vp_n.n148 vp_n.n146 0.369
R16915 vp_n.n150 vp_n.n148 0.369
R16916 vp_n.n152 vp_n.n150 0.369
R16917 vp_n.n154 vp_n.n152 0.369
R16918 vp_n.n156 vp_n.n154 0.369
R16919 vp_n.n158 vp_n.n156 0.369
R16920 vp_n.n160 vp_n.n158 0.369
R16921 vp_n.n162 vp_n.n160 0.369
R16922 vp_n.n164 vp_n.n162 0.369
R16923 vp_n.n166 vp_n.n164 0.369
R16924 vp_n.n168 vp_n.n166 0.369
R16925 vp_n.n170 vp_n.n168 0.369
R16926 vp_n.n172 vp_n.n170 0.369
R16927 vp_n.n174 vp_n.n172 0.369
R16928 vp_n.n176 vp_n.n174 0.369
R16929 vp_n.n178 vp_n.n176 0.369
R16930 vp_n.n180 vp_n.n178 0.369
R16931 vp_n.n182 vp_n.n180 0.369
R16932 vp_n.n184 vp_n.n182 0.369
R16933 vp_n.n186 vp_n.n184 0.369
R16934 vp_n.n188 vp_n.n186 0.369
R16935 vp_n.n190 vp_n.n188 0.369
R16936 vp_n.n192 vp_n.n190 0.369
R16937 vp_n.n194 vp_n.n192 0.369
R16938 vp_n.n196 vp_n.n194 0.369
R16939 vp_n.n198 vp_n.n196 0.369
R16940 vp_n.n200 vp_n.n198 0.369
R16941 vp_n.n202 vp_n.n200 0.369
R16942 vp_n.n204 vp_n.n202 0.369
R16943 vp_n.n206 vp_n.n204 0.369
R16944 vp_n.n208 vp_n.n206 0.369
R16945 vp_n.n210 vp_n.n208 0.369
R16946 vp_n.n212 vp_n.n210 0.369
R16947 vp_n.n214 vp_n.n212 0.369
R16948 vp_n.n216 vp_n.n214 0.369
R16949 vp_n.n218 vp_n.n216 0.369
R16950 vp_n.n220 vp_n.n218 0.369
R16951 vp_n.n222 vp_n.n220 0.369
R16952 vp_n vp_n.n297 0.03
R16953 vss.n194 vss.t516 7.272
R16954 vss.n491 vss.t41 7.272
R16955 vss.n411 vss.t409 6.619
R16956 vss.n2 vss.t256 6.619
R16957 vss.n411 vss.t434 4.955
R16958 vss.n2 vss.t57 4.955
R16959 vss.n194 vss.t539 4.95
R16960 vss.n191 vss.t556 4.95
R16961 vss.n191 vss.t298 4.95
R16962 vss.n192 vss.t281 4.95
R16963 vss.n192 vss.t325 4.95
R16964 vss.n195 vss.t509 4.95
R16965 vss.n195 vss.t550 4.95
R16966 vss.n196 vss.t534 4.95
R16967 vss.n196 vss.t276 4.95
R16968 vss.n198 vss.t291 4.95
R16969 vss.n198 vss.t336 4.95
R16970 vss.n199 vss.t317 4.95
R16971 vss.n199 vss.t364 4.95
R16972 vss.n201 vss.t413 4.95
R16973 vss.n201 vss.t321 4.95
R16974 vss.n202 vss.t438 4.95
R16975 vss.n202 vss.t351 4.95
R16976 vss.n204 vss.t368 4.95
R16977 vss.n204 vss.t406 4.95
R16978 vss.n205 vss.t393 4.95
R16979 vss.n205 vss.t431 4.95
R16980 vss.n207 vss.t448 4.95
R16981 vss.n207 vss.t482 4.95
R16982 vss.n208 vss.t468 4.95
R16983 vss.n208 vss.t506 4.95
R16984 vss.n210 vss.t401 4.95
R16985 vss.n210 vss.t441 4.95
R16986 vss.n211 vss.t428 4.95
R16987 vss.n211 vss.t464 4.95
R16988 vss.n213 vss.t476 4.95
R16989 vss.n213 vss.t518 4.95
R16990 vss.n214 vss.t501 4.95
R16991 vss.n214 vss.t541 4.95
R16992 vss.n216 vss.t466 4.95
R16993 vss.n216 vss.t504 4.95
R16994 vss.n217 vss.t492 4.95
R16995 vss.n217 vss.t530 4.95
R16996 vss.n219 vss.t544 4.95
R16997 vss.n219 vss.t285 4.95
R16998 vss.n220 vss.t270 4.95
R16999 vss.n220 vss.t312 4.95
R17000 vss.n222 vss.t329 4.95
R17001 vss.n222 vss.t537 4.95
R17002 vss.n223 vss.t358 4.95
R17003 vss.n223 vss.t265 4.95
R17004 vss.n225 vss.t279 4.95
R17005 vss.n225 vss.t322 4.95
R17006 vss.n226 vss.t307 4.95
R17007 vss.n226 vss.t352 4.95
R17008 vss.n228 vss.t369 4.95
R17009 vss.n228 vss.t408 4.95
R17010 vss.n229 vss.t394 4.95
R17011 vss.n229 vss.t433 4.95
R17012 vss.n231 vss.t355 4.95
R17013 vss.n231 vss.t397 4.95
R17014 vss.n232 vss.t383 4.95
R17015 vss.n232 vss.t424 4.95
R17016 vss.n234 vss.t436 4.95
R17017 vss.n234 vss.t471 4.95
R17018 vss.n235 vss.t459 4.95
R17019 vss.n235 vss.t496 4.95
R17020 vss.n237 vss.t510 4.95
R17021 vss.n237 vss.t467 4.95
R17022 vss.n238 vss.t535 4.95
R17023 vss.n238 vss.t493 4.95
R17024 vss.n240 vss.t505 4.95
R17025 vss.n240 vss.t547 4.95
R17026 vss.n241 vss.t531 4.95
R17027 vss.n241 vss.t273 4.95
R17028 vss.n243 vss.t287 4.95
R17029 vss.n243 vss.t332 4.95
R17030 vss.n244 vss.t314 4.95
R17031 vss.n244 vss.t361 4.95
R17032 vss.n246 vss.t274 4.95
R17033 vss.n246 vss.t315 4.95
R17034 vss.n247 vss.t302 4.95
R17035 vss.n247 vss.t346 4.95
R17036 vss.n249 vss.t362 4.95
R17037 vss.n249 vss.t402 4.95
R17038 vss.n250 vss.t388 4.95
R17039 vss.n250 vss.t429 4.95
R17040 vss.n252 vss.t309 4.95
R17041 vss.n252 vss.t356 4.95
R17042 vss.n253 vss.t340 4.95
R17043 vss.n253 vss.t384 4.95
R17044 vss.n255 vss.t398 4.95
R17045 vss.n255 vss.t437 4.95
R17046 vss.n256 vss.t425 4.95
R17047 vss.n256 vss.t460 4.95
R17048 vss.n258 vss.t473 4.95
R17049 vss.n258 vss.t391 4.95
R17050 vss.n259 vss.t498 4.95
R17051 vss.n259 vss.t417 4.95
R17052 vss.n261 vss.t461 4.95
R17053 vss.n261 vss.t499 4.95
R17054 vss.n262 vss.t485 4.95
R17055 vss.n262 vss.t525 4.95
R17056 vss.n264 vss.t538 4.95
R17057 vss.n264 vss.t280 4.95
R17058 vss.n265 vss.t266 4.95
R17059 vss.n265 vss.t308 4.95
R17060 vss.n267 vss.t494 4.95
R17061 vss.n267 vss.t532 4.95
R17062 vss.n268 vss.t521 4.95
R17063 vss.n268 vss.t560 4.95
R17064 vss.n412 vss.t323 4.95
R17065 vss.n412 vss.t370 4.95
R17066 vss.n413 vss.t353 4.95
R17067 vss.n413 vss.t395 4.95
R17068 vss.n408 vss.t339 4.95
R17069 vss.n408 vss.t546 4.95
R17070 vss.n409 vss.t367 4.95
R17071 vss.n409 vss.t272 4.95
R17072 vss.n405 vss.t552 4.95
R17073 vss.n405 vss.t294 4.95
R17074 vss.n406 vss.t278 4.95
R17075 vss.n406 vss.t320 4.95
R17076 vss.n402 vss.t472 4.95
R17077 vss.n402 vss.t511 4.95
R17078 vss.n403 vss.t497 4.95
R17079 vss.n403 vss.t536 4.95
R17080 vss.n399 vss.t519 4.95
R17081 vss.n399 vss.t558 4.95
R17082 vss.n400 vss.t542 4.95
R17083 vss.n400 vss.t283 4.95
R17084 vss.n396 vss.t442 4.95
R17085 vss.n396 vss.t477 4.95
R17086 vss.n397 vss.t465 4.95
R17087 vss.n397 vss.t502 4.95
R17088 vss.n393 vss.t454 4.95
R17089 vss.n393 vss.t491 4.95
R17090 vss.n394 vss.t475 4.95
R17091 vss.n394 vss.t515 4.95
R17092 vss.n390 vss.t375 4.95
R17093 vss.n390 vss.t414 4.95
R17094 vss.n391 vss.t399 4.95
R17095 vss.n391 vss.t439 4.95
R17096 vss.n387 vss.t422 4.95
R17097 vss.n387 vss.t330 4.95
R17098 vss.n388 vss.t446 4.95
R17099 vss.n388 vss.t359 4.95
R17100 vss.n384 vss.t337 4.95
R17101 vss.n384 vss.t381 4.95
R17102 vss.n385 vss.t365 4.95
R17103 vss.n385 vss.t404 4.95
R17104 vss.n381 vss.t551 4.95
R17105 vss.n381 vss.t292 4.95
R17106 vss.n382 vss.t277 4.95
R17107 vss.n382 vss.t318 4.95
R17108 vss.n378 vss.t450 4.95
R17109 vss.n378 vss.t484 4.95
R17110 vss.n379 vss.t470 4.95
R17111 vss.n379 vss.t508 4.95
R17112 vss.n375 vss.t371 4.95
R17113 vss.n375 vss.t410 4.95
R17114 vss.n376 vss.t396 4.95
R17115 vss.n376 vss.t435 4.95
R17116 vss.n372 vss.t415 4.95
R17117 vss.n372 vss.t324 4.95
R17118 vss.n373 vss.t440 4.95
R17119 vss.n373 vss.t354 4.95
R17120 vss.n369 vss.t331 4.95
R17121 vss.n369 vss.t376 4.95
R17122 vss.n370 vss.t360 4.95
R17123 vss.n370 vss.t400 4.95
R17124 vss.n366 vss.t545 4.95
R17125 vss.n366 vss.t286 4.95
R17126 vss.n367 vss.t271 4.95
R17127 vss.n367 vss.t313 4.95
R17128 vss.n363 vss.t559 4.95
R17129 vss.n363 vss.t301 4.95
R17130 vss.n364 vss.t284 4.95
R17131 vss.n364 vss.t328 4.95
R17132 vss.n360 vss.t478 4.95
R17133 vss.n360 vss.t520 4.95
R17134 vss.n361 vss.t503 4.95
R17135 vss.n361 vss.t543 4.95
R17136 vss.n357 vss.t524 4.95
R17137 vss.n357 vss.t264 4.95
R17138 vss.n358 vss.t549 4.95
R17139 vss.n358 vss.t290 4.95
R17140 vss.n354 vss.t449 4.95
R17141 vss.n354 vss.t483 4.95
R17142 vss.n355 vss.t469 4.95
R17143 vss.n355 vss.t507 4.95
R17144 vss.n351 vss.t489 4.95
R17145 vss.n351 vss.t407 4.95
R17146 vss.n352 vss.t513 4.95
R17147 vss.n352 vss.t432 4.95
R17148 vss.n348 vss.t382 4.95
R17149 vss.n348 vss.t423 4.95
R17150 vss.n349 vss.t405 4.95
R17151 vss.n349 vss.t447 4.95
R17152 vss.n345 vss.t293 4.95
R17153 vss.n345 vss.t338 4.95
R17154 vss.n346 vss.t319 4.95
R17155 vss.n346 vss.t366 4.95
R17156 vss.n342 vss.t344 4.95
R17157 vss.n342 vss.t387 4.95
R17158 vss.n343 vss.t373 4.95
R17159 vss.n343 vss.t412 4.95
R17160 vss.n339 vss.t557 4.95
R17161 vss.n339 vss.t299 4.95
R17162 vss.n340 vss.t282 4.95
R17163 vss.n340 vss.t326 4.95
R17164 vss.n336 vss.t304 4.95
R17165 vss.n336 vss.t517 4.95
R17166 vss.n337 vss.t333 4.95
R17167 vss.n337 vss.t540 4.95
R17168 vss.n333 vss.t490 4.95
R17169 vss.n333 vss.t529 4.95
R17170 vss.n334 vss.t514 4.95
R17171 vss.n334 vss.t555 4.95
R17172 vss.n330 vss.t533 4.95
R17173 vss.n330 vss.t453 4.95
R17174 vss.n331 vss.t561 4.95
R17175 vss.n331 vss.t474 4.95
R17176 vss.n327 vss.t456 4.95
R17177 vss.n327 vss.t495 4.95
R17178 vss.n328 vss.t479 4.95
R17179 vss.n328 vss.t522 4.95
R17180 vss.n324 vss.t380 4.95
R17181 vss.n324 vss.t419 4.95
R17182 vss.n325 vss.t403 4.95
R17183 vss.n325 vss.t443 4.95
R17184 vss.n321 vss.t426 4.95
R17185 vss.n321 vss.t462 4.95
R17186 vss.n322 vss.t451 4.95
R17187 vss.n322 vss.t486 4.95
R17188 vss.n318 vss.t305 4.95
R17189 vss.n318 vss.t349 4.95
R17190 vss.n319 vss.t334 4.95
R17191 vss.n319 vss.t378 4.95
R17192 vss.n315 vss.t357 4.95
R17193 vss.n315 vss.t262 4.95
R17194 vss.n316 vss.t385 4.95
R17195 vss.n316 vss.t288 4.95
R17196 vss.n312 vss.t267 4.95
R17197 vss.n312 vss.t310 4.95
R17198 vss.n313 vss.t295 4.95
R17199 vss.n313 vss.t341 4.95
R17200 vss.n309 vss.t488 4.95
R17201 vss.n309 vss.t527 4.95
R17202 vss.n310 vss.t512 4.95
R17203 vss.n310 vss.t553 4.95
R17204 vss.n306 vss.t420 4.95
R17205 vss.n306 vss.t457 4.95
R17206 vss.n307 vss.t444 4.95
R17207 vss.n307 vss.t480 4.95
R17208 vss.n303 vss.t300 4.95
R17209 vss.n303 vss.t345 4.95
R17210 vss.n304 vss.t327 4.95
R17211 vss.n304 vss.t374 4.95
R17212 vss.n300 vss.t350 4.95
R17213 vss.n300 vss.t392 4.95
R17214 vss.n301 vss.t379 4.95
R17215 vss.n301 vss.t418 4.95
R17216 vss.n297 vss.t263 4.95
R17217 vss.n297 vss.t306 4.95
R17218 vss.n298 vss.t289 4.95
R17219 vss.n298 vss.t335 4.95
R17220 vss.n294 vss.t311 4.95
R17221 vss.n294 vss.t523 4.95
R17222 vss.n295 vss.t342 4.95
R17223 vss.n295 vss.t548 4.95
R17224 vss.n291 vss.t528 4.95
R17225 vss.n291 vss.t268 4.95
R17226 vss.n292 vss.t554 4.95
R17227 vss.n292 vss.t296 4.95
R17228 vss.n288 vss.t421 4.95
R17229 vss.n288 vss.t458 4.95
R17230 vss.n289 vss.t445 4.95
R17231 vss.n289 vss.t481 4.95
R17232 vss.n285 vss.t463 4.95
R17233 vss.n285 vss.t500 4.95
R17234 vss.n286 vss.t487 4.95
R17235 vss.n286 vss.t526 4.95
R17236 vss.n282 vss.t386 4.95
R17237 vss.n282 vss.t427 4.95
R17238 vss.n283 vss.t411 4.95
R17239 vss.n283 vss.t452 4.95
R17240 vss.n279 vss.t430 4.95
R17241 vss.n279 vss.t343 4.95
R17242 vss.n280 vss.t455 4.95
R17243 vss.n280 vss.t372 4.95
R17244 vss.n276 vss.t348 4.95
R17245 vss.n276 vss.t390 4.95
R17246 vss.n277 vss.t377 4.95
R17247 vss.n277 vss.t416 4.95
R17248 vss.n273 vss.t363 4.95
R17249 vss.n273 vss.t269 4.95
R17250 vss.n274 vss.t389 4.95
R17251 vss.n274 vss.t297 4.95
R17252 vss.n270 vss.t275 4.95
R17253 vss.n270 vss.t316 4.95
R17254 vss.n271 vss.t303 4.95
R17255 vss.n271 vss.t347 4.95
R17256 vss.n594 vss.t40 4.95
R17257 vss.n594 vss.t197 4.95
R17258 vss.n595 vss.t37 4.95
R17259 vss.n595 vss.t44 4.95
R17260 vss.n590 vss.t98 4.95
R17261 vss.n590 vss.t171 4.95
R17262 vss.n591 vss.t62 4.95
R17263 vss.n591 vss.t125 4.95
R17264 vss.n586 vss.t569 4.95
R17265 vss.n586 vss.t101 4.95
R17266 vss.n587 vss.t594 4.95
R17267 vss.n587 vss.t120 4.95
R17268 vss.n582 vss.t186 4.95
R17269 vss.n582 vss.t126 4.95
R17270 vss.n583 vss.t158 4.95
R17271 vss.n583 vss.t15 4.95
R17272 vss.n578 vss.t225 4.95
R17273 vss.n578 vss.t32 4.95
R17274 vss.n579 vss.t199 4.95
R17275 vss.n579 vss.t581 4.95
R17276 vss.n574 vss.t570 4.95
R17277 vss.n574 vss.t246 4.95
R17278 vss.n575 vss.t24 4.95
R17279 vss.n575 vss.t51 4.95
R17280 vss.n570 vss.t160 4.95
R17281 vss.n570 vss.t130 4.95
R17282 vss.n571 vss.t91 4.95
R17283 vss.n571 vss.t146 4.95
R17284 vss.n566 vss.t210 4.95
R17285 vss.n566 vss.t21 4.95
R17286 vss.n567 vss.t248 4.95
R17287 vss.n567 vss.t82 4.95
R17288 vss.n562 vss.t582 4.95
R17289 vss.n562 vss.t205 4.95
R17290 vss.n563 vss.t179 4.95
R17291 vss.n563 vss.t36 4.95
R17292 vss.n558 vss.t563 4.95
R17293 vss.n558 vss.t139 4.95
R17294 vss.n559 vss.t589 4.95
R17295 vss.n559 vss.t103 4.95
R17296 vss.n554 vss.t20 4.95
R17297 vss.n554 vss.t154 4.95
R17298 vss.n555 vss.t81 4.95
R17299 vss.n555 vss.t67 4.95
R17300 vss.n550 vss.t170 4.95
R17301 vss.n550 vss.t209 4.95
R17302 vss.n551 vss.t142 4.95
R17303 vss.n551 vss.t247 4.95
R17304 vss.n546 vss.t100 4.95
R17305 vss.n546 vss.t96 4.95
R17306 vss.n547 vss.t109 4.95
R17307 vss.n547 vss.t60 4.95
R17308 vss.n542 vss.t153 4.95
R17309 vss.n542 vss.t562 4.95
R17310 vss.n543 vss.t66 4.95
R17311 vss.n543 vss.t588 4.95
R17312 vss.n538 vss.t31 4.95
R17313 vss.n538 vss.t185 4.95
R17314 vss.n539 vss.t580 4.95
R17315 vss.n539 vss.t157 4.95
R17316 vss.n534 vss.t213 4.95
R17317 vss.n534 vss.t224 4.95
R17318 vss.n535 vss.t189 4.95
R17319 vss.n535 vss.t217 4.95
R17320 vss.n530 vss.t129 4.95
R17321 vss.n530 vss.t260 4.95
R17322 vss.n531 vss.t145 4.95
R17323 vss.n531 vss.t119 4.95
R17324 vss.n526 vss.t19 4.95
R17325 vss.n526 vss.t159 4.95
R17326 vss.n527 vss.t11 4.95
R17327 vss.n527 vss.t89 4.95
R17328 vss.n522 vss.t204 4.95
R17329 vss.n522 vss.t194 4.95
R17330 vss.n523 vss.t173 4.95
R17331 vss.n523 vss.t212 4.95
R17332 vss.n518 vss.t138 4.95
R17333 vss.n518 vss.t115 4.95
R17334 vss.n519 vss.t102 4.95
R17335 vss.n519 vss.t99 4.95
R17336 vss.n514 vss.t567 4.95
R17337 vss.n514 vss.t177 4.95
R17338 vss.n515 vss.t593 4.95
R17339 vss.n515 vss.t108 4.95
R17340 vss.n510 vss.t239 4.95
R17341 vss.n510 vss.t167 4.95
R17342 vss.n511 vss.t237 4.95
R17343 vss.n511 vss.t71 4.95
R17344 vss.n506 vss.t252 4.95
R17345 vss.n506 vss.t576 4.95
R17346 vss.n507 vss.t55 4.95
R17347 vss.n507 vss.t254 4.95
R17348 vss.n502 vss.t2 4.95
R17349 vss.n502 vss.t242 4.95
R17350 vss.n503 vss.t132 4.95
R17351 vss.n503 vss.t49 4.95
R17352 vss.n498 vss.t56 4.95
R17353 vss.n498 vss.t221 4.95
R17354 vss.n499 vss.t22 4.95
R17355 vss.n499 vss.t161 4.95
R17356 vss.n494 vss.t198 4.95
R17357 vss.n494 vss.t17 4.95
R17358 vss.n495 vss.t47 4.95
R17359 vss.n495 vss.t10 4.95
R17360 vss.n491 vss.t140 4.95
R17361 vss.n4 vss.t118 4.95
R17362 vss.n4 vss.t203 4.95
R17363 vss.n5 vss.t207 4.95
R17364 vss.n5 vss.t195 4.95
R17365 vss.n7 vss.t163 4.95
R17366 vss.n7 vss.t74 4.95
R17367 vss.n8 vss.t92 4.95
R17368 vss.n8 vss.t229 4.95
R17369 vss.n11 vss.t211 4.95
R17370 vss.n11 vss.t23 4.95
R17371 vss.n12 vss.t249 4.95
R17372 vss.n12 vss.t83 4.95
R17373 vss.n15 vss.t97 4.95
R17374 vss.n15 vss.t172 4.95
R17375 vss.n16 vss.t61 4.95
R17376 vss.n16 vss.t143 4.95
R17377 vss.n19 vss.t107 4.95
R17378 vss.n19 vss.t183 4.95
R17379 vss.n20 vss.t124 4.95
R17380 vss.n20 vss.t30 4.95
R17381 vss.n23 vss.t70 4.95
R17382 vss.n23 vss.t592 4.95
R17383 vss.n24 vss.t4 4.95
R17384 vss.n24 vss.t244 4.95
R17385 vss.n27 vss.t577 4.95
R17386 vss.n27 vss.t155 4.95
R17387 vss.n28 vss.t257 4.95
R17388 vss.n28 vss.t218 4.95
R17389 vss.n31 vss.t261 4.95
R17390 vss.n31 vss.t214 4.95
R17391 vss.n32 vss.t77 4.95
R17392 vss.n32 vss.t190 4.95
R17393 vss.n35 vss.t29 4.95
R17394 vss.n35 vss.t131 4.95
R17395 vss.n36 vss.t114 4.95
R17396 vss.n36 vss.t147 4.95
R17397 vss.n39 vss.t9 4.95
R17398 vss.n39 vss.t232 4.95
R17399 vss.n40 vss.t88 4.95
R17400 vss.n40 vss.t137 4.95
R17401 vss.n43 vss.t39 4.95
R17402 vss.n43 vss.t46 4.95
R17403 vss.n44 vss.t598 4.95
R17404 vss.n44 vss.t151 4.95
R17405 vss.n47 vss.t12 4.95
R17406 vss.n47 vss.t90 4.95
R17407 vss.n48 vss.t564 4.95
R17408 vss.n48 vss.t174 4.95
R17409 vss.n51 vss.t141 4.95
R17410 vss.n51 vss.t48 4.95
R17411 vss.n52 vss.t187 4.95
R17412 vss.n52 vss.t164 4.95
R17413 vss.n55 vss.t65 4.95
R17414 vss.n55 vss.t184 4.95
R17415 vss.n56 vss.t578 4.95
R17416 vss.n56 vss.t33 4.95
R17417 vss.n59 vss.t243 4.95
R17418 vss.n59 vss.t123 4.95
R17419 vss.n60 vss.t50 4.95
R17420 vss.n60 vss.t215 4.95
R17421 vss.n63 vss.t222 4.95
R17422 vss.n63 vss.t3 4.95
R17423 vss.n64 vss.t162 4.95
R17424 vss.n64 vss.t133 4.95
R17425 vss.n67 vss.t202 4.95
R17426 vss.n67 vss.t255 4.95
R17427 vss.n68 vss.t196 4.95
R17428 vss.n68 vss.t58 4.95
R17429 vss.n71 vss.t144 4.95
R17430 vss.n71 vss.t117 4.95
R17431 vss.n72 vss.t583 4.95
R17432 vss.n72 vss.t206 4.95
R17433 vss.n75 vss.t136 4.95
R17434 vss.n75 vss.t112 4.95
R17435 vss.n76 vss.t178 4.95
R17436 vss.n76 vss.t95 4.95
R17437 vss.n79 vss.t150 4.95
R17438 vss.n79 vss.t86 4.95
R17439 vss.n80 vss.t168 4.95
R17440 vss.n80 vss.t568 4.95
R17441 vss.n83 vss.t14 4.95
R17442 vss.n83 vss.t597 4.95
R17443 vss.n84 vss.t234 4.95
R17444 vss.n84 vss.t240 4.95
R17445 vss.n87 vss.t591 4.95
R17446 vss.n87 vss.t106 4.95
R17447 vss.n88 vss.t245 4.95
R17448 vss.n88 vss.t223 4.95
R17449 vss.n91 vss.t236 4.95
R17450 vss.n91 vss.t69 4.95
R17451 vss.n92 vss.t72 4.95
R17452 vss.n92 vss.t5 4.95
R17453 vss.n95 vss.t54 4.95
R17454 vss.n95 vss.t220 4.95
R17455 vss.n96 vss.t18 4.95
R17456 vss.n96 vss.t76 4.95
R17457 vss.n99 vss.t79 4.95
R17458 vss.n99 vss.t192 4.95
R17459 vss.n100 vss.t43 4.95
R17460 vss.n100 vss.t208 4.95
R17461 vss.n103 vss.t585 4.95
R17462 vss.n103 vss.t111 4.95
R17463 vss.n104 vss.t181 4.95
R17464 vss.n104 vss.t587 4.95
R17465 vss.n107 vss.t45 4.95
R17466 vss.n107 vss.t8 4.95
R17467 vss.n108 vss.t152 4.95
R17468 vss.n108 vss.t87 4.95
R17469 vss.n111 vss.t128 4.95
R17470 vss.n111 vss.t38 4.95
R17471 vss.n112 vss.t238 4.95
R17472 vss.n112 vss.t599 4.95
R17473 vss.n115 vss.t121 4.95
R17474 vss.n115 vss.t63 4.95
R17475 vss.n116 vss.t227 4.95
R17476 vss.n116 vss.t35 4.95
R17477 vss.n119 vss.t1 4.95
R17478 vss.n119 vss.t595 4.95
R17479 vss.n120 vss.t574 4.95
R17480 vss.n120 vss.t259 4.95
R17481 vss.n123 vss.t75 4.95
R17482 vss.n123 vss.t572 4.95
R17483 vss.n124 vss.t230 4.95
R17484 vss.n124 vss.t25 4.95
R17485 vss.n127 vss.t52 4.95
R17486 vss.n127 vss.t200 4.95
R17487 vss.n128 vss.t80 4.95
R17488 vss.n128 vss.t193 4.95
R17489 vss.n131 vss.t148 4.95
R17490 vss.n131 vss.t27 4.95
R17491 vss.n132 vss.t586 4.95
R17492 vss.n132 vss.t113 4.95
R17493 vss.n135 vss.t84 4.95
R17494 vss.n135 vss.t93 4.95
R17495 vss.n136 vss.t566 4.95
R17496 vss.n136 vss.t176 4.95
R17497 vss.n139 vss.t127 4.95
R17498 vss.n139 vss.t250 4.95
R17499 vss.n140 vss.t16 4.95
R17500 vss.n140 vss.t166 4.95
R17501 vss.n143 vss.t104 4.95
R17502 vss.n143 vss.t180 4.95
R17503 vss.n144 vss.t122 4.95
R17504 vss.n144 vss.t64 4.95
R17505 vss.n147 vss.t596 4.95
R17506 vss.n147 vss.t251 4.95
R17507 vss.n148 vss.t241 4.95
R17508 vss.n148 vss.t169 4.95
R17509 vss.n151 vss.t34 4.95
R17510 vss.n151 vss.t13 4.95
R17511 vss.n152 vss.t253 4.95
R17512 vss.n152 vss.t235 4.95
R17513 vss.n155 vss.t258 4.95
R17514 vss.n155 vss.t226 4.95
R17515 vss.n156 vss.t116 4.95
R17516 vss.n156 vss.t201 4.95
R17517 vss.n159 vss.t134 4.95
R17518 vss.n159 vss.t573 4.95
R17519 vss.n160 vss.t149 4.95
R17520 vss.n160 vss.t28 4.95
R17521 vss.n163 vss.t6 4.95
R17522 vss.n163 vss.t228 4.95
R17523 vss.n164 vss.t85 4.95
R17524 vss.n164 vss.t135 4.95
R17525 vss.n167 vss.t110 4.95
R17526 vss.n167 vss.t78 4.95
R17527 vss.n168 vss.t94 4.95
R17528 vss.n168 vss.t42 4.95
R17529 vss.n171 vss.t175 4.95
R17530 vss.n171 vss.t584 4.95
R17531 vss.n172 vss.t105 4.95
R17532 vss.n172 vss.t182 4.95
R17533 vss.n175 vss.t165 4.95
R17534 vss.n175 vss.t565 4.95
R17535 vss.n176 vss.t68 4.95
R17536 vss.n176 vss.t590 4.95
R17537 vss.n179 vss.t156 4.95
R17538 vss.n179 vss.t188 4.95
R17539 vss.n180 vss.t219 4.95
R17540 vss.n180 vss.t233 4.95
R17541 vss.n183 vss.t216 4.95
R17542 vss.n183 vss.t579 4.95
R17543 vss.n184 vss.t191 4.95
R17544 vss.n184 vss.t53 4.95
R17545 vss.n187 vss.t571 4.95
R17546 vss.n187 vss.t0 4.95
R17547 vss.n188 vss.t26 4.95
R17548 vss.n188 vss.t575 4.95
R17549 vss.n0 vss.t59 4.95
R17550 vss.n0 vss.t73 4.95
R17551 vss.n1 vss.t7 4.95
R17552 vss.n1 vss.t231 4.95
R17553 vss.n493 vss 1.679
R17554 vss.n489 vss.n194 1.287
R17555 vss.n492 vss.n491 1.287
R17556 vss.n415 vss.n411 0.989
R17557 vss.n3 vss.n2 0.989
R17558 vss.n192 vss.n191 0.76
R17559 vss.n196 vss.n195 0.76
R17560 vss.n199 vss.n198 0.76
R17561 vss.n202 vss.n201 0.76
R17562 vss.n205 vss.n204 0.76
R17563 vss.n208 vss.n207 0.76
R17564 vss.n211 vss.n210 0.76
R17565 vss.n214 vss.n213 0.76
R17566 vss.n217 vss.n216 0.76
R17567 vss.n220 vss.n219 0.76
R17568 vss.n223 vss.n222 0.76
R17569 vss.n226 vss.n225 0.76
R17570 vss.n229 vss.n228 0.76
R17571 vss.n232 vss.n231 0.76
R17572 vss.n235 vss.n234 0.76
R17573 vss.n238 vss.n237 0.76
R17574 vss.n241 vss.n240 0.76
R17575 vss.n244 vss.n243 0.76
R17576 vss.n247 vss.n246 0.76
R17577 vss.n250 vss.n249 0.76
R17578 vss.n253 vss.n252 0.76
R17579 vss.n256 vss.n255 0.76
R17580 vss.n259 vss.n258 0.76
R17581 vss.n262 vss.n261 0.76
R17582 vss.n265 vss.n264 0.76
R17583 vss.n268 vss.n267 0.76
R17584 vss.n413 vss.n412 0.76
R17585 vss.n409 vss.n408 0.76
R17586 vss.n406 vss.n405 0.76
R17587 vss.n403 vss.n402 0.76
R17588 vss.n400 vss.n399 0.76
R17589 vss.n397 vss.n396 0.76
R17590 vss.n394 vss.n393 0.76
R17591 vss.n391 vss.n390 0.76
R17592 vss.n388 vss.n387 0.76
R17593 vss.n385 vss.n384 0.76
R17594 vss.n382 vss.n381 0.76
R17595 vss.n379 vss.n378 0.76
R17596 vss.n376 vss.n375 0.76
R17597 vss.n373 vss.n372 0.76
R17598 vss.n370 vss.n369 0.76
R17599 vss.n367 vss.n366 0.76
R17600 vss.n364 vss.n363 0.76
R17601 vss.n361 vss.n360 0.76
R17602 vss.n358 vss.n357 0.76
R17603 vss.n355 vss.n354 0.76
R17604 vss.n352 vss.n351 0.76
R17605 vss.n349 vss.n348 0.76
R17606 vss.n346 vss.n345 0.76
R17607 vss.n343 vss.n342 0.76
R17608 vss.n340 vss.n339 0.76
R17609 vss.n337 vss.n336 0.76
R17610 vss.n334 vss.n333 0.76
R17611 vss.n331 vss.n330 0.76
R17612 vss.n328 vss.n327 0.76
R17613 vss.n325 vss.n324 0.76
R17614 vss.n322 vss.n321 0.76
R17615 vss.n319 vss.n318 0.76
R17616 vss.n316 vss.n315 0.76
R17617 vss.n313 vss.n312 0.76
R17618 vss.n310 vss.n309 0.76
R17619 vss.n307 vss.n306 0.76
R17620 vss.n304 vss.n303 0.76
R17621 vss.n301 vss.n300 0.76
R17622 vss.n298 vss.n297 0.76
R17623 vss.n295 vss.n294 0.76
R17624 vss.n292 vss.n291 0.76
R17625 vss.n289 vss.n288 0.76
R17626 vss.n286 vss.n285 0.76
R17627 vss.n283 vss.n282 0.76
R17628 vss.n280 vss.n279 0.76
R17629 vss.n277 vss.n276 0.76
R17630 vss.n274 vss.n273 0.76
R17631 vss.n271 vss.n270 0.76
R17632 vss.n595 vss.n594 0.76
R17633 vss.n591 vss.n590 0.76
R17634 vss.n587 vss.n586 0.76
R17635 vss.n583 vss.n582 0.76
R17636 vss.n579 vss.n578 0.76
R17637 vss.n575 vss.n574 0.76
R17638 vss.n571 vss.n570 0.76
R17639 vss.n567 vss.n566 0.76
R17640 vss.n563 vss.n562 0.76
R17641 vss.n559 vss.n558 0.76
R17642 vss.n555 vss.n554 0.76
R17643 vss.n551 vss.n550 0.76
R17644 vss.n547 vss.n546 0.76
R17645 vss.n543 vss.n542 0.76
R17646 vss.n539 vss.n538 0.76
R17647 vss.n535 vss.n534 0.76
R17648 vss.n531 vss.n530 0.76
R17649 vss.n527 vss.n526 0.76
R17650 vss.n523 vss.n522 0.76
R17651 vss.n519 vss.n518 0.76
R17652 vss.n515 vss.n514 0.76
R17653 vss.n511 vss.n510 0.76
R17654 vss.n507 vss.n506 0.76
R17655 vss.n503 vss.n502 0.76
R17656 vss.n499 vss.n498 0.76
R17657 vss.n495 vss.n494 0.76
R17658 vss.n5 vss.n4 0.76
R17659 vss.n8 vss.n7 0.76
R17660 vss.n12 vss.n11 0.76
R17661 vss.n16 vss.n15 0.76
R17662 vss.n20 vss.n19 0.76
R17663 vss.n24 vss.n23 0.76
R17664 vss.n28 vss.n27 0.76
R17665 vss.n32 vss.n31 0.76
R17666 vss.n36 vss.n35 0.76
R17667 vss.n40 vss.n39 0.76
R17668 vss.n44 vss.n43 0.76
R17669 vss.n48 vss.n47 0.76
R17670 vss.n52 vss.n51 0.76
R17671 vss.n56 vss.n55 0.76
R17672 vss.n60 vss.n59 0.76
R17673 vss.n64 vss.n63 0.76
R17674 vss.n68 vss.n67 0.76
R17675 vss.n72 vss.n71 0.76
R17676 vss.n76 vss.n75 0.76
R17677 vss.n80 vss.n79 0.76
R17678 vss.n84 vss.n83 0.76
R17679 vss.n88 vss.n87 0.76
R17680 vss.n92 vss.n91 0.76
R17681 vss.n96 vss.n95 0.76
R17682 vss.n100 vss.n99 0.76
R17683 vss.n104 vss.n103 0.76
R17684 vss.n108 vss.n107 0.76
R17685 vss.n112 vss.n111 0.76
R17686 vss.n116 vss.n115 0.76
R17687 vss.n120 vss.n119 0.76
R17688 vss.n124 vss.n123 0.76
R17689 vss.n128 vss.n127 0.76
R17690 vss.n132 vss.n131 0.76
R17691 vss.n136 vss.n135 0.76
R17692 vss.n140 vss.n139 0.76
R17693 vss.n144 vss.n143 0.76
R17694 vss.n148 vss.n147 0.76
R17695 vss.n152 vss.n151 0.76
R17696 vss.n156 vss.n155 0.76
R17697 vss.n160 vss.n159 0.76
R17698 vss.n164 vss.n163 0.76
R17699 vss.n168 vss.n167 0.76
R17700 vss.n172 vss.n171 0.76
R17701 vss.n176 vss.n175 0.76
R17702 vss.n180 vss.n179 0.76
R17703 vss.n184 vss.n183 0.76
R17704 vss.n188 vss.n187 0.76
R17705 vss.n1 vss.n0 0.76
R17706 vss.n193 vss.n192 0.419
R17707 vss.n197 vss.n196 0.419
R17708 vss.n200 vss.n199 0.419
R17709 vss.n203 vss.n202 0.419
R17710 vss.n206 vss.n205 0.419
R17711 vss.n209 vss.n208 0.419
R17712 vss.n212 vss.n211 0.419
R17713 vss.n215 vss.n214 0.419
R17714 vss.n218 vss.n217 0.419
R17715 vss.n221 vss.n220 0.419
R17716 vss.n224 vss.n223 0.419
R17717 vss.n227 vss.n226 0.419
R17718 vss.n230 vss.n229 0.419
R17719 vss.n233 vss.n232 0.419
R17720 vss.n236 vss.n235 0.419
R17721 vss.n239 vss.n238 0.419
R17722 vss.n242 vss.n241 0.419
R17723 vss.n245 vss.n244 0.419
R17724 vss.n248 vss.n247 0.419
R17725 vss.n251 vss.n250 0.419
R17726 vss.n254 vss.n253 0.419
R17727 vss.n257 vss.n256 0.419
R17728 vss.n260 vss.n259 0.419
R17729 vss.n263 vss.n262 0.419
R17730 vss.n266 vss.n265 0.419
R17731 vss.n269 vss.n268 0.419
R17732 vss.n414 vss.n413 0.419
R17733 vss.n410 vss.n409 0.419
R17734 vss.n407 vss.n406 0.419
R17735 vss.n404 vss.n403 0.419
R17736 vss.n401 vss.n400 0.419
R17737 vss.n398 vss.n397 0.419
R17738 vss.n395 vss.n394 0.419
R17739 vss.n392 vss.n391 0.419
R17740 vss.n389 vss.n388 0.419
R17741 vss.n386 vss.n385 0.419
R17742 vss.n383 vss.n382 0.419
R17743 vss.n380 vss.n379 0.419
R17744 vss.n377 vss.n376 0.419
R17745 vss.n374 vss.n373 0.419
R17746 vss.n371 vss.n370 0.419
R17747 vss.n368 vss.n367 0.419
R17748 vss.n365 vss.n364 0.419
R17749 vss.n362 vss.n361 0.419
R17750 vss.n359 vss.n358 0.419
R17751 vss.n356 vss.n355 0.419
R17752 vss.n353 vss.n352 0.419
R17753 vss.n350 vss.n349 0.419
R17754 vss.n347 vss.n346 0.419
R17755 vss.n344 vss.n343 0.419
R17756 vss.n341 vss.n340 0.419
R17757 vss.n338 vss.n337 0.419
R17758 vss.n335 vss.n334 0.419
R17759 vss.n332 vss.n331 0.419
R17760 vss.n329 vss.n328 0.419
R17761 vss.n326 vss.n325 0.419
R17762 vss.n323 vss.n322 0.419
R17763 vss.n320 vss.n319 0.419
R17764 vss.n317 vss.n316 0.419
R17765 vss.n314 vss.n313 0.419
R17766 vss.n311 vss.n310 0.419
R17767 vss.n308 vss.n307 0.419
R17768 vss.n305 vss.n304 0.419
R17769 vss.n302 vss.n301 0.419
R17770 vss.n299 vss.n298 0.419
R17771 vss.n296 vss.n295 0.419
R17772 vss.n293 vss.n292 0.419
R17773 vss.n290 vss.n289 0.419
R17774 vss.n287 vss.n286 0.419
R17775 vss.n284 vss.n283 0.419
R17776 vss.n281 vss.n280 0.419
R17777 vss.n278 vss.n277 0.419
R17778 vss.n275 vss.n274 0.419
R17779 vss.n272 vss.n271 0.419
R17780 vss.n597 vss.n595 0.419
R17781 vss.n593 vss.n591 0.419
R17782 vss.n589 vss.n587 0.419
R17783 vss.n585 vss.n583 0.419
R17784 vss.n581 vss.n579 0.419
R17785 vss.n577 vss.n575 0.419
R17786 vss.n573 vss.n571 0.419
R17787 vss.n569 vss.n567 0.419
R17788 vss.n565 vss.n563 0.419
R17789 vss.n561 vss.n559 0.419
R17790 vss.n557 vss.n555 0.419
R17791 vss.n553 vss.n551 0.419
R17792 vss.n549 vss.n547 0.419
R17793 vss.n545 vss.n543 0.419
R17794 vss.n541 vss.n539 0.419
R17795 vss.n537 vss.n535 0.419
R17796 vss.n533 vss.n531 0.419
R17797 vss.n529 vss.n527 0.419
R17798 vss.n525 vss.n523 0.419
R17799 vss.n521 vss.n519 0.419
R17800 vss.n517 vss.n515 0.419
R17801 vss.n513 vss.n511 0.419
R17802 vss.n509 vss.n507 0.419
R17803 vss.n505 vss.n503 0.419
R17804 vss.n501 vss.n499 0.419
R17805 vss.n497 vss.n495 0.419
R17806 vss.n6 vss.n5 0.419
R17807 vss.n10 vss.n8 0.419
R17808 vss.n14 vss.n12 0.419
R17809 vss.n18 vss.n16 0.419
R17810 vss.n22 vss.n20 0.419
R17811 vss.n26 vss.n24 0.419
R17812 vss.n30 vss.n28 0.419
R17813 vss.n34 vss.n32 0.419
R17814 vss.n38 vss.n36 0.419
R17815 vss.n42 vss.n40 0.419
R17816 vss.n46 vss.n44 0.419
R17817 vss.n50 vss.n48 0.419
R17818 vss.n54 vss.n52 0.419
R17819 vss.n58 vss.n56 0.419
R17820 vss.n62 vss.n60 0.419
R17821 vss.n66 vss.n64 0.419
R17822 vss.n70 vss.n68 0.419
R17823 vss.n74 vss.n72 0.419
R17824 vss.n78 vss.n76 0.419
R17825 vss.n82 vss.n80 0.419
R17826 vss.n86 vss.n84 0.419
R17827 vss.n90 vss.n88 0.419
R17828 vss.n94 vss.n92 0.419
R17829 vss.n98 vss.n96 0.419
R17830 vss.n102 vss.n100 0.419
R17831 vss.n106 vss.n104 0.419
R17832 vss.n110 vss.n108 0.419
R17833 vss.n114 vss.n112 0.419
R17834 vss.n118 vss.n116 0.419
R17835 vss.n122 vss.n120 0.419
R17836 vss.n126 vss.n124 0.419
R17837 vss.n130 vss.n128 0.419
R17838 vss.n134 vss.n132 0.419
R17839 vss.n138 vss.n136 0.419
R17840 vss.n142 vss.n140 0.419
R17841 vss.n146 vss.n144 0.419
R17842 vss.n150 vss.n148 0.419
R17843 vss.n154 vss.n152 0.419
R17844 vss.n158 vss.n156 0.419
R17845 vss.n162 vss.n160 0.419
R17846 vss.n166 vss.n164 0.419
R17847 vss.n170 vss.n168 0.419
R17848 vss.n174 vss.n172 0.419
R17849 vss.n178 vss.n176 0.419
R17850 vss.n182 vss.n180 0.419
R17851 vss.n186 vss.n184 0.419
R17852 vss.n190 vss.n188 0.419
R17853 vss.n598 vss.n1 0.419
R17854 vss vss.n490 0.226
R17855 vss.n416 vss.n415 0.191
R17856 vss.n452 vss.n451 0.19
R17857 vss.n488 vss.n487 0.189
R17858 vss.n451 vss.n450 0.189
R17859 vss.n417 vss.n416 0.189
R17860 vss.n418 vss.n417 0.189
R17861 vss.n419 vss.n418 0.189
R17862 vss.n420 vss.n419 0.189
R17863 vss.n421 vss.n420 0.189
R17864 vss.n422 vss.n421 0.189
R17865 vss.n423 vss.n422 0.189
R17866 vss.n424 vss.n423 0.189
R17867 vss.n425 vss.n424 0.189
R17868 vss.n426 vss.n425 0.189
R17869 vss.n427 vss.n426 0.189
R17870 vss.n428 vss.n427 0.189
R17871 vss.n429 vss.n428 0.189
R17872 vss.n430 vss.n429 0.189
R17873 vss.n431 vss.n430 0.189
R17874 vss.n432 vss.n431 0.189
R17875 vss.n433 vss.n432 0.189
R17876 vss.n434 vss.n433 0.189
R17877 vss.n435 vss.n434 0.189
R17878 vss.n436 vss.n435 0.189
R17879 vss.n437 vss.n436 0.189
R17880 vss.n438 vss.n437 0.189
R17881 vss.n439 vss.n438 0.189
R17882 vss.n440 vss.n439 0.189
R17883 vss.n441 vss.n440 0.189
R17884 vss.n442 vss.n441 0.189
R17885 vss.n443 vss.n442 0.189
R17886 vss.n444 vss.n443 0.189
R17887 vss.n445 vss.n444 0.189
R17888 vss.n446 vss.n445 0.189
R17889 vss.n447 vss.n446 0.189
R17890 vss.n448 vss.n447 0.189
R17891 vss.n449 vss.n448 0.189
R17892 vss.n450 vss.n449 0.189
R17893 vss.n453 vss.n452 0.189
R17894 vss.n454 vss.n453 0.189
R17895 vss.n455 vss.n454 0.189
R17896 vss.n456 vss.n455 0.189
R17897 vss.n457 vss.n456 0.189
R17898 vss.n458 vss.n457 0.189
R17899 vss.n459 vss.n458 0.189
R17900 vss.n460 vss.n459 0.189
R17901 vss.n461 vss.n460 0.189
R17902 vss.n464 vss.n463 0.189
R17903 vss.n465 vss.n464 0.189
R17904 vss.n466 vss.n465 0.189
R17905 vss.n467 vss.n466 0.189
R17906 vss.n468 vss.n467 0.189
R17907 vss.n469 vss.n468 0.189
R17908 vss.n470 vss.n469 0.189
R17909 vss.n471 vss.n470 0.189
R17910 vss.n472 vss.n471 0.189
R17911 vss.n473 vss.n472 0.189
R17912 vss.n474 vss.n473 0.189
R17913 vss.n475 vss.n474 0.189
R17914 vss.n476 vss.n475 0.189
R17915 vss.n477 vss.n476 0.189
R17916 vss.n478 vss.n477 0.189
R17917 vss.n479 vss.n478 0.189
R17918 vss.n480 vss.n479 0.189
R17919 vss.n481 vss.n480 0.189
R17920 vss.n482 vss.n481 0.189
R17921 vss.n483 vss.n482 0.189
R17922 vss.n484 vss.n483 0.189
R17923 vss.n485 vss.n484 0.189
R17924 vss.n486 vss.n485 0.189
R17925 vss.n487 vss.n486 0.189
R17926 vss.n462 vss.n461 0.189
R17927 vss.n463 vss.n462 0.189
R17928 vss.n489 vss.n488 0.172
R17929 vss.n490 vss.n489 0.012
R17930 vss.n493 vss.n492 0.012
R17931 vss.n414 vss.n410 0.002
R17932 vss.n410 vss.n407 0.002
R17933 vss.n407 vss.n404 0.002
R17934 vss.n404 vss.n401 0.002
R17935 vss.n401 vss.n398 0.002
R17936 vss.n398 vss.n395 0.002
R17937 vss.n395 vss.n392 0.002
R17938 vss.n392 vss.n389 0.002
R17939 vss.n389 vss.n386 0.002
R17940 vss.n386 vss.n383 0.002
R17941 vss.n383 vss.n380 0.002
R17942 vss.n380 vss.n377 0.002
R17943 vss.n377 vss.n374 0.002
R17944 vss.n374 vss.n371 0.002
R17945 vss.n371 vss.n368 0.002
R17946 vss.n368 vss.n365 0.002
R17947 vss.n365 vss.n362 0.002
R17948 vss.n362 vss.n359 0.002
R17949 vss.n359 vss.n356 0.002
R17950 vss.n356 vss.n353 0.002
R17951 vss.n353 vss.n350 0.002
R17952 vss.n350 vss.n347 0.002
R17953 vss.n347 vss.n344 0.002
R17954 vss.n344 vss.n341 0.002
R17955 vss.n341 vss.n338 0.002
R17956 vss.n338 vss.n335 0.002
R17957 vss.n335 vss.n332 0.002
R17958 vss.n332 vss.n329 0.002
R17959 vss.n329 vss.n326 0.002
R17960 vss.n326 vss.n323 0.002
R17961 vss.n323 vss.n320 0.002
R17962 vss.n320 vss.n317 0.002
R17963 vss.n317 vss.n314 0.002
R17964 vss.n314 vss.n311 0.002
R17965 vss.n311 vss.n308 0.002
R17966 vss.n308 vss.n305 0.002
R17967 vss.n305 vss.n302 0.002
R17968 vss.n302 vss.n299 0.002
R17969 vss.n299 vss.n296 0.002
R17970 vss.n296 vss.n293 0.002
R17971 vss.n293 vss.n290 0.002
R17972 vss.n290 vss.n287 0.002
R17973 vss.n287 vss.n284 0.002
R17974 vss.n284 vss.n281 0.002
R17975 vss.n281 vss.n278 0.002
R17976 vss.n278 vss.n275 0.002
R17977 vss.n275 vss.n272 0.002
R17978 vss.n272 vss.n269 0.002
R17979 vss.n269 vss.n266 0.002
R17980 vss.n266 vss.n263 0.002
R17981 vss.n263 vss.n260 0.002
R17982 vss.n260 vss.n257 0.002
R17983 vss.n257 vss.n254 0.002
R17984 vss.n254 vss.n251 0.002
R17985 vss.n251 vss.n248 0.002
R17986 vss.n248 vss.n245 0.002
R17987 vss.n245 vss.n242 0.002
R17988 vss.n242 vss.n239 0.002
R17989 vss.n239 vss.n236 0.002
R17990 vss.n236 vss.n233 0.002
R17991 vss.n233 vss.n230 0.002
R17992 vss.n230 vss.n227 0.002
R17993 vss.n227 vss.n224 0.002
R17994 vss.n224 vss.n221 0.002
R17995 vss.n221 vss.n218 0.002
R17996 vss.n218 vss.n215 0.002
R17997 vss.n215 vss.n212 0.002
R17998 vss.n212 vss.n209 0.002
R17999 vss.n209 vss.n206 0.002
R18000 vss.n206 vss.n203 0.002
R18001 vss.n203 vss.n200 0.002
R18002 vss.n200 vss.n197 0.002
R18003 vss.n197 vss.n193 0.002
R18004 vss.n490 vss.n193 0.002
R18005 vss.n10 vss.n6 0.002
R18006 vss.n14 vss.n10 0.002
R18007 vss.n18 vss.n14 0.002
R18008 vss.n22 vss.n18 0.002
R18009 vss.n26 vss.n22 0.002
R18010 vss.n30 vss.n26 0.002
R18011 vss.n34 vss.n30 0.002
R18012 vss.n38 vss.n34 0.002
R18013 vss.n42 vss.n38 0.002
R18014 vss.n46 vss.n42 0.002
R18015 vss.n50 vss.n46 0.002
R18016 vss.n54 vss.n50 0.002
R18017 vss.n58 vss.n54 0.002
R18018 vss.n62 vss.n58 0.002
R18019 vss.n66 vss.n62 0.002
R18020 vss.n70 vss.n66 0.002
R18021 vss.n74 vss.n70 0.002
R18022 vss.n78 vss.n74 0.002
R18023 vss.n82 vss.n78 0.002
R18024 vss.n86 vss.n82 0.002
R18025 vss.n90 vss.n86 0.002
R18026 vss.n94 vss.n90 0.002
R18027 vss.n98 vss.n94 0.002
R18028 vss.n102 vss.n98 0.002
R18029 vss.n106 vss.n102 0.002
R18030 vss.n110 vss.n106 0.002
R18031 vss.n114 vss.n110 0.002
R18032 vss.n118 vss.n114 0.002
R18033 vss.n122 vss.n118 0.002
R18034 vss.n126 vss.n122 0.002
R18035 vss.n130 vss.n126 0.002
R18036 vss.n134 vss.n130 0.002
R18037 vss.n138 vss.n134 0.002
R18038 vss.n142 vss.n138 0.002
R18039 vss.n146 vss.n142 0.002
R18040 vss.n150 vss.n146 0.002
R18041 vss.n154 vss.n150 0.002
R18042 vss.n158 vss.n154 0.002
R18043 vss.n162 vss.n158 0.002
R18044 vss.n166 vss.n162 0.002
R18045 vss.n170 vss.n166 0.002
R18046 vss.n174 vss.n170 0.002
R18047 vss.n178 vss.n174 0.002
R18048 vss.n182 vss.n178 0.002
R18049 vss.n186 vss.n182 0.002
R18050 vss.n190 vss.n186 0.002
R18051 vss.n598 vss.n190 0.002
R18052 vss.n598 vss.n597 0.002
R18053 vss.n597 vss.n593 0.002
R18054 vss.n593 vss.n589 0.002
R18055 vss.n589 vss.n585 0.002
R18056 vss.n585 vss.n581 0.002
R18057 vss.n581 vss.n577 0.002
R18058 vss.n577 vss.n573 0.002
R18059 vss.n573 vss.n569 0.002
R18060 vss.n569 vss.n565 0.002
R18061 vss.n565 vss.n561 0.002
R18062 vss.n561 vss.n557 0.002
R18063 vss.n557 vss.n553 0.002
R18064 vss.n553 vss.n549 0.002
R18065 vss.n549 vss.n545 0.002
R18066 vss.n545 vss.n541 0.002
R18067 vss.n541 vss.n537 0.002
R18068 vss.n537 vss.n533 0.002
R18069 vss.n533 vss.n529 0.002
R18070 vss.n529 vss.n525 0.002
R18071 vss.n525 vss.n521 0.002
R18072 vss.n521 vss.n517 0.002
R18073 vss.n517 vss.n513 0.002
R18074 vss.n513 vss.n509 0.002
R18075 vss.n509 vss.n505 0.002
R18076 vss.n505 vss.n501 0.002
R18077 vss.n501 vss.n497 0.002
R18078 vss.n497 vss.n493 0.002
R18079 vss.n462 vss.n272 0.001
R18080 vss.n463 vss.n269 0.001
R18081 vss.n464 vss.n266 0.001
R18082 vss.n465 vss.n263 0.001
R18083 vss.n466 vss.n260 0.001
R18084 vss.n467 vss.n257 0.001
R18085 vss.n468 vss.n254 0.001
R18086 vss.n469 vss.n251 0.001
R18087 vss.n470 vss.n248 0.001
R18088 vss.n471 vss.n245 0.001
R18089 vss.n472 vss.n242 0.001
R18090 vss.n473 vss.n239 0.001
R18091 vss.n474 vss.n236 0.001
R18092 vss.n475 vss.n233 0.001
R18093 vss.n476 vss.n230 0.001
R18094 vss.n477 vss.n227 0.001
R18095 vss.n478 vss.n224 0.001
R18096 vss.n479 vss.n221 0.001
R18097 vss.n480 vss.n218 0.001
R18098 vss.n481 vss.n215 0.001
R18099 vss.n482 vss.n212 0.001
R18100 vss.n483 vss.n209 0.001
R18101 vss.n484 vss.n206 0.001
R18102 vss.n485 vss.n203 0.001
R18103 vss.n486 vss.n200 0.001
R18104 vss.n487 vss.n197 0.001
R18105 vss.n416 vss.n410 0.001
R18106 vss.n417 vss.n407 0.001
R18107 vss.n418 vss.n404 0.001
R18108 vss.n419 vss.n401 0.001
R18109 vss.n420 vss.n398 0.001
R18110 vss.n421 vss.n395 0.001
R18111 vss.n422 vss.n392 0.001
R18112 vss.n423 vss.n389 0.001
R18113 vss.n424 vss.n386 0.001
R18114 vss.n425 vss.n383 0.001
R18115 vss.n426 vss.n380 0.001
R18116 vss.n427 vss.n377 0.001
R18117 vss.n428 vss.n374 0.001
R18118 vss.n429 vss.n371 0.001
R18119 vss.n430 vss.n368 0.001
R18120 vss.n431 vss.n365 0.001
R18121 vss.n432 vss.n362 0.001
R18122 vss.n433 vss.n359 0.001
R18123 vss.n434 vss.n356 0.001
R18124 vss.n435 vss.n353 0.001
R18125 vss.n436 vss.n350 0.001
R18126 vss.n437 vss.n347 0.001
R18127 vss.n438 vss.n344 0.001
R18128 vss.n439 vss.n341 0.001
R18129 vss.n440 vss.n338 0.001
R18130 vss.n441 vss.n335 0.001
R18131 vss.n442 vss.n332 0.001
R18132 vss.n443 vss.n329 0.001
R18133 vss.n444 vss.n326 0.001
R18134 vss.n445 vss.n323 0.001
R18135 vss.n446 vss.n320 0.001
R18136 vss.n447 vss.n317 0.001
R18137 vss.n448 vss.n314 0.001
R18138 vss.n449 vss.n311 0.001
R18139 vss.n450 vss.n308 0.001
R18140 vss.n452 vss.n302 0.001
R18141 vss.n453 vss.n299 0.001
R18142 vss.n454 vss.n296 0.001
R18143 vss.n455 vss.n293 0.001
R18144 vss.n456 vss.n290 0.001
R18145 vss.n457 vss.n287 0.001
R18146 vss.n458 vss.n284 0.001
R18147 vss.n459 vss.n281 0.001
R18148 vss.n460 vss.n278 0.001
R18149 vss.n461 vss.n275 0.001
R18150 vss.n599 vss.n598 0.001
R18151 vss.n10 vss.n9 0.001
R18152 vss.n14 vss.n13 0.001
R18153 vss.n18 vss.n17 0.001
R18154 vss.n22 vss.n21 0.001
R18155 vss.n26 vss.n25 0.001
R18156 vss.n30 vss.n29 0.001
R18157 vss.n34 vss.n33 0.001
R18158 vss.n38 vss.n37 0.001
R18159 vss.n42 vss.n41 0.001
R18160 vss.n46 vss.n45 0.001
R18161 vss.n50 vss.n49 0.001
R18162 vss.n54 vss.n53 0.001
R18163 vss.n58 vss.n57 0.001
R18164 vss.n62 vss.n61 0.001
R18165 vss.n66 vss.n65 0.001
R18166 vss.n70 vss.n69 0.001
R18167 vss.n74 vss.n73 0.001
R18168 vss.n78 vss.n77 0.001
R18169 vss.n82 vss.n81 0.001
R18170 vss.n86 vss.n85 0.001
R18171 vss.n90 vss.n89 0.001
R18172 vss.n94 vss.n93 0.001
R18173 vss.n98 vss.n97 0.001
R18174 vss.n102 vss.n101 0.001
R18175 vss.n106 vss.n105 0.001
R18176 vss.n110 vss.n109 0.001
R18177 vss.n114 vss.n113 0.001
R18178 vss.n118 vss.n117 0.001
R18179 vss.n122 vss.n121 0.001
R18180 vss.n126 vss.n125 0.001
R18181 vss.n130 vss.n129 0.001
R18182 vss.n134 vss.n133 0.001
R18183 vss.n138 vss.n137 0.001
R18184 vss.n142 vss.n141 0.001
R18185 vss.n146 vss.n145 0.001
R18186 vss.n154 vss.n153 0.001
R18187 vss.n158 vss.n157 0.001
R18188 vss.n162 vss.n161 0.001
R18189 vss.n166 vss.n165 0.001
R18190 vss.n170 vss.n169 0.001
R18191 vss.n174 vss.n173 0.001
R18192 vss.n178 vss.n177 0.001
R18193 vss.n182 vss.n181 0.001
R18194 vss.n186 vss.n185 0.001
R18195 vss.n190 vss.n189 0.001
R18196 vss.n451 vss.n305 0.001
R18197 vss.n150 vss.n149 0.001
R18198 vss.n497 vss.n496 0.001
R18199 vss.n501 vss.n500 0.001
R18200 vss.n505 vss.n504 0.001
R18201 vss.n509 vss.n508 0.001
R18202 vss.n513 vss.n512 0.001
R18203 vss.n517 vss.n516 0.001
R18204 vss.n521 vss.n520 0.001
R18205 vss.n525 vss.n524 0.001
R18206 vss.n529 vss.n528 0.001
R18207 vss.n533 vss.n532 0.001
R18208 vss.n537 vss.n536 0.001
R18209 vss.n541 vss.n540 0.001
R18210 vss.n545 vss.n544 0.001
R18211 vss.n549 vss.n548 0.001
R18212 vss.n553 vss.n552 0.001
R18213 vss.n557 vss.n556 0.001
R18214 vss.n561 vss.n560 0.001
R18215 vss.n565 vss.n564 0.001
R18216 vss.n569 vss.n568 0.001
R18217 vss.n573 vss.n572 0.001
R18218 vss.n577 vss.n576 0.001
R18219 vss.n581 vss.n580 0.001
R18220 vss.n585 vss.n584 0.001
R18221 vss.n589 vss.n588 0.001
R18222 vss.n593 vss.n592 0.001
R18223 vss.n597 vss.n596 0.001
R18224 vss.n488 vss.n193 0.001
R18225 vss.n415 vss.n414 0.001
R18226 vss.n6 vss.n3 0.001
R18227 vn_n.n147 vn_n.t139 721.861
R18228 vn_n.n145 vn_n.t253 721.861
R18229 vn_n.n143 vn_n.t174 721.861
R18230 vn_n.n141 vn_n.t244 721.861
R18231 vn_n.n139 vn_n.t53 721.861
R18232 vn_n.n137 vn_n.t284 721.861
R18233 vn_n.n135 vn_n.t93 721.861
R18234 vn_n.n133 vn_n.t16 721.861
R18235 vn_n.n131 vn_n.t259 721.861
R18236 vn_n.n129 vn_n.t184 721.861
R18237 vn_n.n127 vn_n.t120 721.861
R18238 vn_n.n125 vn_n.t233 721.861
R18239 vn_n.n123 vn_n.t158 721.861
R18240 vn_n.n121 vn_n.t100 721.861
R18241 vn_n.n119 vn_n.t24 721.861
R18242 vn_n.n117 vn_n.t260 721.861
R18243 vn_n.n115 vn_n.t280 721.861
R18244 vn_n.n113 vn_n.t208 721.861
R18245 vn_n.n111 vn_n.t142 721.861
R18246 vn_n.n109 vn_n.t76 721.861
R18247 vn_n.n107 vn_n.t178 721.861
R18248 vn_n.n105 vn_n.t117 721.861
R18249 vn_n.n103 vn_n.t45 721.861
R18250 vn_n.n101 vn_n.t286 721.861
R18251 vn_n.n99 vn_n.t218 721.861
R18252 vn_n.n97 vn_n.t20 721.861
R18253 vn_n.n95 vn_n.t256 721.861
R18254 vn_n.n93 vn_n.t179 721.861
R18255 vn_n.n91 vn_n.t123 721.861
R18256 vn_n.n89 vn_n.t57 721.861
R18257 vn_n.n87 vn_n.t161 721.861
R18258 vn_n.n85 vn_n.t96 721.861
R18259 vn_n.n83 vn_n.t202 721.861
R18260 vn_n.n81 vn_n.t264 721.861
R18261 vn_n.n79 vn_n.t189 721.861
R18262 vn_n.n77 vn_n.t0 721.861
R18263 vn_n.n75 vn_n.t236 721.861
R18264 vn_n.n73 vn_n.t40 721.861
R18265 vn_n.n71 vn_n.t104 721.861
R18266 vn_n.n69 vn_n.t38 721.861
R18267 vn_n.n67 vn_n.t274 721.861
R18268 vn_n.n65 vn_n.t200 721.861
R18269 vn_n.n63 vn_n.t7 721.861
R18270 vn_n.n61 vn_n.t73 721.861
R18271 vn_n.n59 vn_n.t173 721.861
R18272 vn_n.n57 vn_n.t111 721.861
R18273 vn_n.n55 vn_n.t39 721.861
R18274 vn_n.n53 vn_n.t146 721.861
R18275 vn_n.n51 vn_n.t211 721.861
R18276 vn_n.n49 vn_n.t14 721.861
R18277 vn_n.n47 vn_n.t251 721.861
R18278 vn_n.n45 vn_n.t63 721.861
R18279 vn_n.n43 vn_n.t290 721.861
R18280 vn_n.n41 vn_n.t49 721.861
R18281 vn_n.n39 vn_n.t155 721.861
R18282 vn_n.n37 vn_n.t91 721.861
R18283 vn_n.n35 vn_n.t196 721.861
R18284 vn_n.n33 vn_n.t128 721.861
R18285 vn_n.n31 vn_n.t69 721.861
R18286 vn_n.n29 vn_n.t296 721.861
R18287 vn_n.n27 vn_n.t231 721.861
R18288 vn_n.n25 vn_n.t33 721.861
R18289 vn_n.n23 vn_n.t270 721.861
R18290 vn_n.n21 vn_n.t31 721.861
R18291 vn_n.n19 vn_n.t267 721.861
R18292 vn_n.n17 vn_n.t195 721.861
R18293 vn_n.n15 vn_n.t3 721.861
R18294 vn_n.n13 vn_n.t239 721.861
R18295 vn_n.n11 vn_n.t170 721.861
R18296 vn_n.n9 vn_n.t107 721.861
R18297 vn_n.n7 vn_n.t217 721.861
R18298 vn_n.n5 vn_n.t143 721.861
R18299 vn_n.n3 vn_n.t79 721.861
R18300 vn_n.n1 vn_n.t10 721.861
R18301 vn_n.n0 vn_n.t248 721.861
R18302 vn_n.n147 vn_n.t148 721.861
R18303 vn_n.n145 vn_n.t262 721.861
R18304 vn_n.n143 vn_n.t187 721.861
R18305 vn_n.n141 vn_n.t252 721.861
R18306 vn_n.n139 vn_n.t64 721.861
R18307 vn_n.n137 vn_n.t292 721.861
R18308 vn_n.n135 vn_n.t102 721.861
R18309 vn_n.n133 vn_n.t27 721.861
R18310 vn_n.n131 vn_n.t269 721.861
R18311 vn_n.n129 vn_n.t197 721.861
R18312 vn_n.n127 vn_n.t130 721.861
R18313 vn_n.n125 vn_n.t242 721.861
R18314 vn_n.n123 vn_n.t166 721.861
R18315 vn_n.n121 vn_n.t109 721.861
R18316 vn_n.n119 vn_n.t34 721.861
R18317 vn_n.n117 vn_n.t271 721.861
R18318 vn_n.n115 vn_n.t288 721.861
R18319 vn_n.n113 vn_n.t220 721.861
R18320 vn_n.n111 vn_n.t151 721.861
R18321 vn_n.n109 vn_n.t87 721.861
R18322 vn_n.n107 vn_n.t190 721.861
R18323 vn_n.n105 vn_n.t125 721.861
R18324 vn_n.n103 vn_n.t59 721.861
R18325 vn_n.n101 vn_n.t293 721.861
R18326 vn_n.n99 vn_n.t228 721.861
R18327 vn_n.n97 vn_n.t29 721.861
R18328 vn_n.n95 vn_n.t265 721.861
R18329 vn_n.n93 vn_n.t192 721.861
R18330 vn_n.n91 vn_n.t132 721.861
R18331 vn_n.n89 vn_n.t66 721.861
R18332 vn_n.n87 vn_n.t168 721.861
R18333 vn_n.n85 vn_n.t105 721.861
R18334 vn_n.n83 vn_n.t214 721.861
R18335 vn_n.n81 vn_n.t275 721.861
R18336 vn_n.n79 vn_n.t201 721.861
R18337 vn_n.n77 vn_n.t8 721.861
R18338 vn_n.n75 vn_n.t245 721.861
R18339 vn_n.n73 vn_n.t55 721.861
R18340 vn_n.n71 vn_n.t112 721.861
R18341 vn_n.n69 vn_n.t51 721.861
R18342 vn_n.n67 vn_n.t283 721.861
R18343 vn_n.n65 vn_n.t212 721.861
R18344 vn_n.n63 vn_n.t15 721.861
R18345 vn_n.n61 vn_n.t82 721.861
R18346 vn_n.n59 vn_n.t182 721.861
R18347 vn_n.n57 vn_n.t119 721.861
R18348 vn_n.n55 vn_n.t52 721.861
R18349 vn_n.n53 vn_n.t157 721.861
R18350 vn_n.n51 vn_n.t222 721.861
R18351 vn_n.n49 vn_n.t23 721.861
R18352 vn_n.n47 vn_n.t258 721.861
R18353 vn_n.n45 vn_n.t70 721.861
R18354 vn_n.n43 vn_n.t298 721.861
R18355 vn_n.n41 vn_n.t61 721.861
R18356 vn_n.n39 vn_n.t164 721.861
R18357 vn_n.n37 vn_n.t99 721.861
R18358 vn_n.n35 vn_n.t209 721.861
R18359 vn_n.n33 vn_n.t137 721.861
R18360 vn_n.n31 vn_n.t78 721.861
R18361 vn_n.n29 vn_n.t5 721.861
R18362 vn_n.n27 vn_n.t240 721.861
R18363 vn_n.n25 vn_n.t46 721.861
R18364 vn_n.n23 vn_n.t281 721.861
R18365 vn_n.n21 vn_n.t42 721.861
R18366 vn_n.n19 vn_n.t278 721.861
R18367 vn_n.n17 vn_n.t206 721.861
R18368 vn_n.n15 vn_n.t12 721.861
R18369 vn_n.n13 vn_n.t249 721.861
R18370 vn_n.n11 vn_n.t176 721.861
R18371 vn_n.n9 vn_n.t114 721.861
R18372 vn_n.n7 vn_n.t227 721.861
R18373 vn_n.n5 vn_n.t152 721.861
R18374 vn_n.n3 vn_n.t88 721.861
R18375 vn_n.n1 vn_n.t19 721.861
R18376 vn_n.n0 vn_n.t254 721.861
R18377 vn_n.n149 vn_n.t129 691.553
R18378 vn_n.n224 vn_n.t136 691.553
R18379 vn_n.n222 vn_n.t21 690.412
R18380 vn_n.n221 vn_n.t257 690.412
R18381 vn_n.n220 vn_n.t68 690.412
R18382 vn_n.n219 vn_n.t295 690.412
R18383 vn_n.n218 vn_n.t238 690.412
R18384 vn_n.n217 vn_n.t163 690.412
R18385 vn_n.n216 vn_n.t98 690.412
R18386 vn_n.n215 vn_n.t207 690.412
R18387 vn_n.n214 vn_n.t135 690.412
R18388 vn_n.n213 vn_n.t75 690.412
R18389 vn_n.n212 vn_n.t2 690.412
R18390 vn_n.n211 vn_n.t116 690.412
R18391 vn_n.n210 vn_n.t44 690.412
R18392 vn_n.n209 vn_n.t279 690.412
R18393 vn_n.n208 vn_n.t216 690.412
R18394 vn_n.n207 vn_n.t141 690.412
R18395 vn_n.n206 vn_n.t159 690.412
R18396 vn_n.n205 vn_n.t94 690.412
R18397 vn_n.n204 vn_n.t17 690.412
R18398 vn_n.n203 vn_n.t261 690.412
R18399 vn_n.n202 vn_n.t185 690.412
R18400 vn_n.n201 vn_n.t299 690.412
R18401 vn_n.n200 vn_n.t234 690.412
R18402 vn_n.n199 vn_n.t37 690.412
R18403 vn_n.n198 vn_n.t101 690.412
R18404 vn_n.n197 vn_n.t25 690.412
R18405 vn_n.n196 vn_n.t138 690.412
R18406 vn_n.n195 vn_n.t71 690.412
R18407 vn_n.n194 vn_n.t172 690.412
R18408 vn_n.n193 vn_n.t241 690.412
R18409 vn_n.n192 vn_n.t47 690.412
R18410 vn_n.n191 vn_n.t282 690.412
R18411 vn_n.n190 vn_n.t210 690.412
R18412 vn_n.n189 vn_n.t13 690.412
R18413 vn_n.n188 vn_n.t80 690.412
R18414 vn_n.n187 vn_n.t181 690.412
R18415 vn_n.n186 vn_n.t118 690.412
R18416 vn_n.n185 vn_n.t48 690.412
R18417 vn_n.n184 vn_n.t154 690.412
R18418 vn_n.n183 vn_n.t221 690.412
R18419 vn_n.n182 vn_n.t153 690.412
R18420 vn_n.n181 vn_n.t89 690.412
R18421 vn_n.n180 vn_n.t193 690.412
R18422 vn_n.n179 vn_n.t126 690.412
R18423 vn_n.n178 vn_n.t180 690.412
R18424 vn_n.n177 vn_n.t294 690.412
R18425 vn_n.n176 vn_n.t229 690.412
R18426 vn_n.n175 vn_n.t30 690.412
R18427 vn_n.n174 vn_n.t266 690.412
R18428 vn_n.n173 vn_n.t203 690.412
R18429 vn_n.n172 vn_n.t133 690.412
R18430 vn_n.n171 vn_n.t67 690.412
R18431 vn_n.n170 vn_n.t169 690.412
R18432 vn_n.n169 vn_n.t106 690.412
R18433 vn_n.n168 vn_n.t41 690.412
R18434 vn_n.n167 vn_n.t276 690.412
R18435 vn_n.n166 vn_n.t204 690.412
R18436 vn_n.n165 vn_n.t9 690.412
R18437 vn_n.n164 vn_n.t247 690.412
R18438 vn_n.n163 vn_n.t175 690.412
R18439 vn_n.n162 vn_n.t113 690.412
R18440 vn_n.n161 vn_n.t225 690.412
R18441 vn_n.n160 vn_n.t149 690.412
R18442 vn_n.n159 vn_n.t86 690.412
R18443 vn_n.n158 vn_n.t147 690.412
R18444 vn_n.n157 vn_n.t84 690.412
R18445 vn_n.n156 vn_n.t186 690.412
R18446 vn_n.n155 vn_n.t121 690.412
R18447 vn_n.n154 vn_n.t56 690.412
R18448 vn_n.n153 vn_n.t291 690.412
R18449 vn_n.n152 vn_n.t224 690.412
R18450 vn_n.n151 vn_n.t26 690.412
R18451 vn_n.n150 vn_n.t263 690.412
R18452 vn_n.n149 vn_n.t72 690.412
R18453 vn_n.n224 vn_n.t81 690.412
R18454 vn_n.n225 vn_n.t273 690.412
R18455 vn_n.n226 vn_n.t35 690.412
R18456 vn_n.n227 vn_n.t232 690.412
R18457 vn_n.n228 vn_n.t297 690.412
R18458 vn_n.n229 vn_n.t65 690.412
R18459 vn_n.n230 vn_n.t131 690.412
R18460 vn_n.n231 vn_n.t199 690.412
R18461 vn_n.n232 vn_n.t92 690.412
R18462 vn_n.n233 vn_n.t156 690.412
R18463 vn_n.n234 vn_n.t95 690.412
R18464 vn_n.n235 vn_n.t160 690.412
R18465 vn_n.n236 vn_n.t235 690.412
R18466 vn_n.n237 vn_n.t122 690.412
R18467 vn_n.n238 vn_n.t188 690.412
R18468 vn_n.n239 vn_n.t255 690.412
R18469 vn_n.n240 vn_n.t18 690.412
R18470 vn_n.n241 vn_n.t215 690.412
R18471 vn_n.n242 vn_n.t285 690.412
R18472 vn_n.n243 vn_n.t54 690.412
R18473 vn_n.n244 vn_n.t115 690.412
R18474 vn_n.n245 vn_n.t177 690.412
R18475 vn_n.n246 vn_n.t74 690.412
R18476 vn_n.n247 vn_n.t140 690.412
R18477 vn_n.n248 vn_n.t213 690.412
R18478 vn_n.n249 vn_n.t277 690.412
R18479 vn_n.n250 vn_n.t43 690.412
R18480 vn_n.n251 vn_n.t237 690.412
R18481 vn_n.n252 vn_n.t1 690.412
R18482 vn_n.n253 vn_n.t191 690.412
R18483 vn_n.n254 vn_n.t134 690.412
R18484 vn_n.n255 vn_n.t205 690.412
R18485 vn_n.n256 vn_n.t97 690.412
R18486 vn_n.n257 vn_n.t162 690.412
R18487 vn_n.n258 vn_n.t230 690.412
R18488 vn_n.n259 vn_n.t165 690.412
R18489 vn_n.n260 vn_n.t62 690.412
R18490 vn_n.n261 vn_n.t127 690.412
R18491 vn_n.n262 vn_n.t194 690.412
R18492 vn_n.n263 vn_n.t90 690.412
R18493 vn_n.n264 vn_n.t22 690.412
R18494 vn_n.n265 vn_n.t223 690.412
R18495 vn_n.n266 vn_n.t289 690.412
R18496 vn_n.n267 vn_n.t60 690.412
R18497 vn_n.n268 vn_n.t250 690.412
R18498 vn_n.n269 vn_n.t183 690.412
R18499 vn_n.n270 vn_n.t83 690.412
R18500 vn_n.n271 vn_n.t145 690.412
R18501 vn_n.n272 vn_n.t36 690.412
R18502 vn_n.n273 vn_n.t110 690.412
R18503 vn_n.n274 vn_n.t50 690.412
R18504 vn_n.n275 vn_n.t243 690.412
R18505 vn_n.n276 vn_n.t6 690.412
R18506 vn_n.n277 vn_n.t198 690.412
R18507 vn_n.n278 vn_n.t272 690.412
R18508 vn_n.n279 vn_n.t28 690.412
R18509 vn_n.n280 vn_n.t103 690.412
R18510 vn_n.n281 vn_n.t167 690.412
R18511 vn_n.n282 vn_n.t150 690.412
R18512 vn_n.n283 vn_n.t226 690.412
R18513 vn_n.n284 vn_n.t287 690.412
R18514 vn_n.n285 vn_n.t58 690.412
R18515 vn_n.n286 vn_n.t124 690.412
R18516 vn_n.n287 vn_n.t11 690.412
R18517 vn_n.n288 vn_n.t85 690.412
R18518 vn_n.n289 vn_n.t144 690.412
R18519 vn_n.n290 vn_n.t219 690.412
R18520 vn_n.n291 vn_n.t108 690.412
R18521 vn_n.n292 vn_n.t171 690.412
R18522 vn_n.n293 vn_n.t246 690.412
R18523 vn_n.n294 vn_n.t4 690.412
R18524 vn_n.n295 vn_n.t77 690.412
R18525 vn_n.n296 vn_n.t268 690.412
R18526 vn_n.n297 vn_n.t32 690.412
R18527 vn_n.n2 vn_n.n0 6.382
R18528 vn_n.n2 vn_n.n1 6.013
R18529 vn_n.n4 vn_n.n3 6.013
R18530 vn_n.n6 vn_n.n5 6.013
R18531 vn_n.n8 vn_n.n7 6.013
R18532 vn_n.n10 vn_n.n9 6.013
R18533 vn_n.n12 vn_n.n11 6.013
R18534 vn_n.n14 vn_n.n13 6.013
R18535 vn_n.n16 vn_n.n15 6.013
R18536 vn_n.n18 vn_n.n17 6.013
R18537 vn_n.n20 vn_n.n19 6.013
R18538 vn_n.n22 vn_n.n21 6.013
R18539 vn_n.n24 vn_n.n23 6.013
R18540 vn_n.n26 vn_n.n25 6.013
R18541 vn_n.n28 vn_n.n27 6.013
R18542 vn_n.n30 vn_n.n29 6.013
R18543 vn_n.n32 vn_n.n31 6.013
R18544 vn_n.n34 vn_n.n33 6.013
R18545 vn_n.n36 vn_n.n35 6.013
R18546 vn_n.n38 vn_n.n37 6.013
R18547 vn_n.n40 vn_n.n39 6.013
R18548 vn_n.n42 vn_n.n41 6.013
R18549 vn_n.n44 vn_n.n43 6.013
R18550 vn_n.n46 vn_n.n45 6.013
R18551 vn_n.n48 vn_n.n47 6.013
R18552 vn_n.n50 vn_n.n49 6.013
R18553 vn_n.n52 vn_n.n51 6.013
R18554 vn_n.n54 vn_n.n53 6.013
R18555 vn_n.n56 vn_n.n55 6.013
R18556 vn_n.n58 vn_n.n57 6.013
R18557 vn_n.n60 vn_n.n59 6.013
R18558 vn_n.n62 vn_n.n61 6.013
R18559 vn_n.n64 vn_n.n63 6.013
R18560 vn_n.n66 vn_n.n65 6.013
R18561 vn_n.n68 vn_n.n67 6.013
R18562 vn_n.n70 vn_n.n69 6.013
R18563 vn_n.n72 vn_n.n71 6.013
R18564 vn_n.n74 vn_n.n73 6.013
R18565 vn_n.n76 vn_n.n75 6.013
R18566 vn_n.n78 vn_n.n77 6.013
R18567 vn_n.n80 vn_n.n79 6.013
R18568 vn_n.n82 vn_n.n81 6.013
R18569 vn_n.n84 vn_n.n83 6.013
R18570 vn_n.n86 vn_n.n85 6.013
R18571 vn_n.n88 vn_n.n87 6.013
R18572 vn_n.n90 vn_n.n89 6.013
R18573 vn_n.n92 vn_n.n91 6.013
R18574 vn_n.n94 vn_n.n93 6.013
R18575 vn_n.n96 vn_n.n95 6.013
R18576 vn_n.n98 vn_n.n97 6.013
R18577 vn_n.n100 vn_n.n99 6.013
R18578 vn_n.n102 vn_n.n101 6.013
R18579 vn_n.n104 vn_n.n103 6.013
R18580 vn_n.n106 vn_n.n105 6.013
R18581 vn_n.n108 vn_n.n107 6.013
R18582 vn_n.n110 vn_n.n109 6.013
R18583 vn_n.n112 vn_n.n111 6.013
R18584 vn_n.n114 vn_n.n113 6.013
R18585 vn_n.n116 vn_n.n115 6.013
R18586 vn_n.n118 vn_n.n117 6.013
R18587 vn_n.n120 vn_n.n119 6.013
R18588 vn_n.n122 vn_n.n121 6.013
R18589 vn_n.n124 vn_n.n123 6.013
R18590 vn_n.n126 vn_n.n125 6.013
R18591 vn_n.n128 vn_n.n127 6.013
R18592 vn_n.n130 vn_n.n129 6.013
R18593 vn_n.n132 vn_n.n131 6.013
R18594 vn_n.n134 vn_n.n133 6.013
R18595 vn_n.n136 vn_n.n135 6.013
R18596 vn_n.n138 vn_n.n137 6.013
R18597 vn_n.n140 vn_n.n139 6.013
R18598 vn_n.n142 vn_n.n141 6.013
R18599 vn_n.n144 vn_n.n143 6.013
R18600 vn_n.n146 vn_n.n145 6.013
R18601 vn_n.n148 vn_n.n147 6.013
R18602 vn_n vn_n.n297 1.227
R18603 vn_n.n150 vn_n.n149 1.141
R18604 vn_n.n151 vn_n.n150 1.141
R18605 vn_n.n152 vn_n.n151 1.141
R18606 vn_n.n153 vn_n.n152 1.141
R18607 vn_n.n154 vn_n.n153 1.141
R18608 vn_n.n155 vn_n.n154 1.141
R18609 vn_n.n156 vn_n.n155 1.141
R18610 vn_n.n157 vn_n.n156 1.141
R18611 vn_n.n158 vn_n.n157 1.141
R18612 vn_n.n159 vn_n.n158 1.141
R18613 vn_n.n160 vn_n.n159 1.141
R18614 vn_n.n161 vn_n.n160 1.141
R18615 vn_n.n162 vn_n.n161 1.141
R18616 vn_n.n163 vn_n.n162 1.141
R18617 vn_n.n164 vn_n.n163 1.141
R18618 vn_n.n165 vn_n.n164 1.141
R18619 vn_n.n166 vn_n.n165 1.141
R18620 vn_n.n167 vn_n.n166 1.141
R18621 vn_n.n168 vn_n.n167 1.141
R18622 vn_n.n169 vn_n.n168 1.141
R18623 vn_n.n170 vn_n.n169 1.141
R18624 vn_n.n171 vn_n.n170 1.141
R18625 vn_n.n172 vn_n.n171 1.141
R18626 vn_n.n173 vn_n.n172 1.141
R18627 vn_n.n174 vn_n.n173 1.141
R18628 vn_n.n175 vn_n.n174 1.141
R18629 vn_n.n176 vn_n.n175 1.141
R18630 vn_n.n177 vn_n.n176 1.141
R18631 vn_n.n178 vn_n.n177 1.141
R18632 vn_n.n179 vn_n.n178 1.141
R18633 vn_n.n180 vn_n.n179 1.141
R18634 vn_n.n181 vn_n.n180 1.141
R18635 vn_n.n182 vn_n.n181 1.141
R18636 vn_n.n183 vn_n.n182 1.141
R18637 vn_n.n184 vn_n.n183 1.141
R18638 vn_n.n185 vn_n.n184 1.141
R18639 vn_n.n186 vn_n.n185 1.141
R18640 vn_n.n187 vn_n.n186 1.141
R18641 vn_n.n188 vn_n.n187 1.141
R18642 vn_n.n189 vn_n.n188 1.141
R18643 vn_n.n190 vn_n.n189 1.141
R18644 vn_n.n191 vn_n.n190 1.141
R18645 vn_n.n192 vn_n.n191 1.141
R18646 vn_n.n193 vn_n.n192 1.141
R18647 vn_n.n194 vn_n.n193 1.141
R18648 vn_n.n195 vn_n.n194 1.141
R18649 vn_n.n196 vn_n.n195 1.141
R18650 vn_n.n197 vn_n.n196 1.141
R18651 vn_n.n198 vn_n.n197 1.141
R18652 vn_n.n199 vn_n.n198 1.141
R18653 vn_n.n200 vn_n.n199 1.141
R18654 vn_n.n201 vn_n.n200 1.141
R18655 vn_n.n202 vn_n.n201 1.141
R18656 vn_n.n203 vn_n.n202 1.141
R18657 vn_n.n204 vn_n.n203 1.141
R18658 vn_n.n205 vn_n.n204 1.141
R18659 vn_n.n206 vn_n.n205 1.141
R18660 vn_n.n207 vn_n.n206 1.141
R18661 vn_n.n208 vn_n.n207 1.141
R18662 vn_n.n209 vn_n.n208 1.141
R18663 vn_n.n210 vn_n.n209 1.141
R18664 vn_n.n211 vn_n.n210 1.141
R18665 vn_n.n212 vn_n.n211 1.141
R18666 vn_n.n213 vn_n.n212 1.141
R18667 vn_n.n214 vn_n.n213 1.141
R18668 vn_n.n215 vn_n.n214 1.141
R18669 vn_n.n216 vn_n.n215 1.141
R18670 vn_n.n217 vn_n.n216 1.141
R18671 vn_n.n218 vn_n.n217 1.141
R18672 vn_n.n219 vn_n.n218 1.141
R18673 vn_n.n220 vn_n.n219 1.141
R18674 vn_n.n221 vn_n.n220 1.141
R18675 vn_n.n222 vn_n.n221 1.141
R18676 vn_n.n225 vn_n.n224 1.141
R18677 vn_n.n226 vn_n.n225 1.141
R18678 vn_n.n227 vn_n.n226 1.141
R18679 vn_n.n228 vn_n.n227 1.141
R18680 vn_n.n229 vn_n.n228 1.141
R18681 vn_n.n230 vn_n.n229 1.141
R18682 vn_n.n231 vn_n.n230 1.141
R18683 vn_n.n232 vn_n.n231 1.141
R18684 vn_n.n233 vn_n.n232 1.141
R18685 vn_n.n234 vn_n.n233 1.141
R18686 vn_n.n235 vn_n.n234 1.141
R18687 vn_n.n236 vn_n.n235 1.141
R18688 vn_n.n237 vn_n.n236 1.141
R18689 vn_n.n238 vn_n.n237 1.141
R18690 vn_n.n239 vn_n.n238 1.141
R18691 vn_n.n240 vn_n.n239 1.141
R18692 vn_n.n241 vn_n.n240 1.141
R18693 vn_n.n242 vn_n.n241 1.141
R18694 vn_n.n243 vn_n.n242 1.141
R18695 vn_n.n244 vn_n.n243 1.141
R18696 vn_n.n245 vn_n.n244 1.141
R18697 vn_n.n246 vn_n.n245 1.141
R18698 vn_n.n247 vn_n.n246 1.141
R18699 vn_n.n248 vn_n.n247 1.141
R18700 vn_n.n249 vn_n.n248 1.141
R18701 vn_n.n250 vn_n.n249 1.141
R18702 vn_n.n251 vn_n.n250 1.141
R18703 vn_n.n252 vn_n.n251 1.141
R18704 vn_n.n253 vn_n.n252 1.141
R18705 vn_n.n254 vn_n.n253 1.141
R18706 vn_n.n255 vn_n.n254 1.141
R18707 vn_n.n256 vn_n.n255 1.141
R18708 vn_n.n257 vn_n.n256 1.141
R18709 vn_n.n258 vn_n.n257 1.141
R18710 vn_n.n259 vn_n.n258 1.141
R18711 vn_n.n260 vn_n.n259 1.141
R18712 vn_n.n261 vn_n.n260 1.141
R18713 vn_n.n262 vn_n.n261 1.141
R18714 vn_n.n263 vn_n.n262 1.141
R18715 vn_n.n264 vn_n.n263 1.141
R18716 vn_n.n265 vn_n.n264 1.141
R18717 vn_n.n266 vn_n.n265 1.141
R18718 vn_n.n267 vn_n.n266 1.141
R18719 vn_n.n268 vn_n.n267 1.141
R18720 vn_n.n269 vn_n.n268 1.141
R18721 vn_n.n270 vn_n.n269 1.141
R18722 vn_n.n271 vn_n.n270 1.141
R18723 vn_n.n272 vn_n.n271 1.141
R18724 vn_n.n273 vn_n.n272 1.141
R18725 vn_n.n274 vn_n.n273 1.141
R18726 vn_n.n275 vn_n.n274 1.141
R18727 vn_n.n276 vn_n.n275 1.141
R18728 vn_n.n277 vn_n.n276 1.141
R18729 vn_n.n278 vn_n.n277 1.141
R18730 vn_n.n279 vn_n.n278 1.141
R18731 vn_n.n280 vn_n.n279 1.141
R18732 vn_n.n281 vn_n.n280 1.141
R18733 vn_n.n282 vn_n.n281 1.141
R18734 vn_n.n283 vn_n.n282 1.141
R18735 vn_n.n284 vn_n.n283 1.141
R18736 vn_n.n285 vn_n.n284 1.141
R18737 vn_n.n286 vn_n.n285 1.141
R18738 vn_n.n287 vn_n.n286 1.141
R18739 vn_n.n288 vn_n.n287 1.141
R18740 vn_n.n289 vn_n.n288 1.141
R18741 vn_n.n290 vn_n.n289 1.141
R18742 vn_n.n291 vn_n.n290 1.141
R18743 vn_n.n292 vn_n.n291 1.141
R18744 vn_n.n293 vn_n.n292 1.141
R18745 vn_n.n294 vn_n.n293 1.141
R18746 vn_n.n295 vn_n.n294 1.141
R18747 vn_n.n296 vn_n.n295 1.141
R18748 vn_n.n297 vn_n.n296 1.141
R18749 vn_n.n223 vn_n.n222 0.946
R18750 vn_n.n223 vn_n.n148 0.397
R18751 vn_n.n4 vn_n.n2 0.369
R18752 vn_n.n6 vn_n.n4 0.369
R18753 vn_n.n8 vn_n.n6 0.369
R18754 vn_n.n10 vn_n.n8 0.369
R18755 vn_n.n12 vn_n.n10 0.369
R18756 vn_n.n14 vn_n.n12 0.369
R18757 vn_n.n16 vn_n.n14 0.369
R18758 vn_n.n18 vn_n.n16 0.369
R18759 vn_n.n20 vn_n.n18 0.369
R18760 vn_n.n22 vn_n.n20 0.369
R18761 vn_n.n24 vn_n.n22 0.369
R18762 vn_n.n26 vn_n.n24 0.369
R18763 vn_n.n28 vn_n.n26 0.369
R18764 vn_n.n30 vn_n.n28 0.369
R18765 vn_n.n32 vn_n.n30 0.369
R18766 vn_n.n34 vn_n.n32 0.369
R18767 vn_n.n36 vn_n.n34 0.369
R18768 vn_n.n38 vn_n.n36 0.369
R18769 vn_n.n40 vn_n.n38 0.369
R18770 vn_n.n42 vn_n.n40 0.369
R18771 vn_n.n44 vn_n.n42 0.369
R18772 vn_n.n46 vn_n.n44 0.369
R18773 vn_n.n48 vn_n.n46 0.369
R18774 vn_n.n50 vn_n.n48 0.369
R18775 vn_n.n52 vn_n.n50 0.369
R18776 vn_n.n54 vn_n.n52 0.369
R18777 vn_n.n56 vn_n.n54 0.369
R18778 vn_n.n58 vn_n.n56 0.369
R18779 vn_n.n60 vn_n.n58 0.369
R18780 vn_n.n62 vn_n.n60 0.369
R18781 vn_n.n64 vn_n.n62 0.369
R18782 vn_n.n66 vn_n.n64 0.369
R18783 vn_n.n68 vn_n.n66 0.369
R18784 vn_n.n70 vn_n.n68 0.369
R18785 vn_n.n72 vn_n.n70 0.369
R18786 vn_n.n74 vn_n.n72 0.369
R18787 vn_n.n76 vn_n.n74 0.369
R18788 vn_n.n78 vn_n.n76 0.369
R18789 vn_n.n80 vn_n.n78 0.369
R18790 vn_n.n82 vn_n.n80 0.369
R18791 vn_n.n84 vn_n.n82 0.369
R18792 vn_n.n86 vn_n.n84 0.369
R18793 vn_n.n88 vn_n.n86 0.369
R18794 vn_n.n90 vn_n.n88 0.369
R18795 vn_n.n92 vn_n.n90 0.369
R18796 vn_n.n94 vn_n.n92 0.369
R18797 vn_n.n96 vn_n.n94 0.369
R18798 vn_n.n98 vn_n.n96 0.369
R18799 vn_n.n100 vn_n.n98 0.369
R18800 vn_n.n102 vn_n.n100 0.369
R18801 vn_n.n104 vn_n.n102 0.369
R18802 vn_n.n106 vn_n.n104 0.369
R18803 vn_n.n108 vn_n.n106 0.369
R18804 vn_n.n110 vn_n.n108 0.369
R18805 vn_n.n112 vn_n.n110 0.369
R18806 vn_n.n114 vn_n.n112 0.369
R18807 vn_n.n116 vn_n.n114 0.369
R18808 vn_n.n118 vn_n.n116 0.369
R18809 vn_n.n120 vn_n.n118 0.369
R18810 vn_n.n122 vn_n.n120 0.369
R18811 vn_n.n124 vn_n.n122 0.369
R18812 vn_n.n126 vn_n.n124 0.369
R18813 vn_n.n128 vn_n.n126 0.369
R18814 vn_n.n130 vn_n.n128 0.369
R18815 vn_n.n132 vn_n.n130 0.369
R18816 vn_n.n134 vn_n.n132 0.369
R18817 vn_n.n136 vn_n.n134 0.369
R18818 vn_n.n138 vn_n.n136 0.369
R18819 vn_n.n140 vn_n.n138 0.369
R18820 vn_n.n142 vn_n.n140 0.369
R18821 vn_n.n144 vn_n.n142 0.369
R18822 vn_n.n146 vn_n.n144 0.369
R18823 vn_n.n148 vn_n.n146 0.369
R18824 vn_n vn_n.n223 0.03
C8 vn_n vss 211.75fF
C9 out_n vss 1049.19fF
C10 vn_p vss 351.92fF
C11 vp_p vss 351.92fF
C12 out_p vss 1048.31fF
C13 vp_n vss 211.49fF
C14 vdd2 vss 1217.91fF
C15 vdd1 vss 1213.72fF
C16 vn_n.n2 vss 1.56fF $ **FLOATING
C17 vn_n.n4 vss 1.00fF $ **FLOATING
C18 vn_n.n6 vss 1.00fF $ **FLOATING
C19 vn_n.n8 vss 1.00fF $ **FLOATING
C20 vn_n.n10 vss 1.00fF $ **FLOATING
C21 vn_n.n12 vss 1.00fF $ **FLOATING
C22 vn_n.n14 vss 1.00fF $ **FLOATING
C23 vn_n.n16 vss 1.00fF $ **FLOATING
C24 vn_n.n18 vss 1.00fF $ **FLOATING
C25 vn_n.n20 vss 1.00fF $ **FLOATING
C26 vn_n.n22 vss 1.00fF $ **FLOATING
C27 vn_n.n24 vss 1.00fF $ **FLOATING
C28 vn_n.n26 vss 1.00fF $ **FLOATING
C29 vn_n.n28 vss 1.00fF $ **FLOATING
C30 vn_n.n30 vss 1.00fF $ **FLOATING
C31 vn_n.n32 vss 1.00fF $ **FLOATING
C32 vn_n.n34 vss 1.00fF $ **FLOATING
C33 vn_n.n36 vss 1.00fF $ **FLOATING
C34 vn_n.n38 vss 1.00fF $ **FLOATING
C35 vn_n.n40 vss 1.00fF $ **FLOATING
C36 vn_n.n42 vss 1.00fF $ **FLOATING
C37 vn_n.n44 vss 1.00fF $ **FLOATING
C38 vn_n.n46 vss 1.00fF $ **FLOATING
C39 vn_n.n48 vss 1.00fF $ **FLOATING
C40 vn_n.n50 vss 1.00fF $ **FLOATING
C41 vn_n.n52 vss 1.00fF $ **FLOATING
C42 vn_n.n54 vss 1.00fF $ **FLOATING
C43 vn_n.n56 vss 1.00fF $ **FLOATING
C44 vn_n.n58 vss 1.00fF $ **FLOATING
C45 vn_n.n60 vss 1.00fF $ **FLOATING
C46 vn_n.n62 vss 1.00fF $ **FLOATING
C47 vn_n.n64 vss 1.00fF $ **FLOATING
C48 vn_n.n66 vss 1.00fF $ **FLOATING
C49 vn_n.n68 vss 1.00fF $ **FLOATING
C50 vn_n.n70 vss 1.00fF $ **FLOATING
C51 vn_n.n72 vss 1.00fF $ **FLOATING
C52 vn_n.n74 vss 1.00fF $ **FLOATING
C53 vn_n.n76 vss 1.00fF $ **FLOATING
C54 vn_n.n78 vss 1.00fF $ **FLOATING
C55 vn_n.n80 vss 1.00fF $ **FLOATING
C56 vn_n.n82 vss 1.00fF $ **FLOATING
C57 vn_n.n84 vss 1.00fF $ **FLOATING
C58 vn_n.n86 vss 1.00fF $ **FLOATING
C59 vn_n.n88 vss 1.00fF $ **FLOATING
C60 vn_n.n90 vss 1.00fF $ **FLOATING
C61 vn_n.n92 vss 1.00fF $ **FLOATING
C62 vn_n.n94 vss 1.00fF $ **FLOATING
C63 vn_n.n96 vss 1.00fF $ **FLOATING
C64 vn_n.n98 vss 1.00fF $ **FLOATING
C65 vn_n.n100 vss 1.00fF $ **FLOATING
C66 vn_n.n102 vss 1.00fF $ **FLOATING
C67 vn_n.n104 vss 1.00fF $ **FLOATING
C68 vn_n.n106 vss 1.00fF $ **FLOATING
C69 vn_n.n108 vss 1.00fF $ **FLOATING
C70 vn_n.n110 vss 1.00fF $ **FLOATING
C71 vn_n.n112 vss 1.00fF $ **FLOATING
C72 vn_n.n114 vss 1.00fF $ **FLOATING
C73 vn_n.n116 vss 1.00fF $ **FLOATING
C74 vn_n.n118 vss 1.00fF $ **FLOATING
C75 vn_n.n120 vss 1.00fF $ **FLOATING
C76 vn_n.n122 vss 1.00fF $ **FLOATING
C77 vn_n.n124 vss 1.00fF $ **FLOATING
C78 vn_n.n126 vss 1.00fF $ **FLOATING
C79 vn_n.n128 vss 1.00fF $ **FLOATING
C80 vn_n.n130 vss 1.00fF $ **FLOATING
C81 vn_n.n132 vss 1.00fF $ **FLOATING
C82 vn_n.n134 vss 1.00fF $ **FLOATING
C83 vn_n.n136 vss 1.00fF $ **FLOATING
C84 vn_n.n138 vss 1.00fF $ **FLOATING
C85 vn_n.n140 vss 1.00fF $ **FLOATING
C86 vn_n.n142 vss 1.00fF $ **FLOATING
C87 vn_n.n144 vss 1.00fF $ **FLOATING
C88 vn_n.n146 vss 1.00fF $ **FLOATING
C89 vn_n.n148 vss 1.04fF $ **FLOATING
C90 vn_n.n149 vss 1.16fF $ **FLOATING
C91 vn_n.n222 vss 1.56fF $ **FLOATING
C92 vn_n.n223 vss 12.59fF $ **FLOATING
C93 vn_n.n224 vss 1.09fF $ **FLOATING
C94 vp_n.n0 vss 1.10fF $ **FLOATING
C95 vp_n.n76 vss 1.56fF $ **FLOATING
C96 vp_n.n78 vss 1.00fF $ **FLOATING
C97 vp_n.n80 vss 1.00fF $ **FLOATING
C98 vp_n.n82 vss 1.00fF $ **FLOATING
C99 vp_n.n84 vss 1.00fF $ **FLOATING
C100 vp_n.n86 vss 1.00fF $ **FLOATING
C101 vp_n.n88 vss 1.00fF $ **FLOATING
C102 vp_n.n90 vss 1.00fF $ **FLOATING
C103 vp_n.n92 vss 1.00fF $ **FLOATING
C104 vp_n.n94 vss 1.00fF $ **FLOATING
C105 vp_n.n96 vss 1.00fF $ **FLOATING
C106 vp_n.n98 vss 1.00fF $ **FLOATING
C107 vp_n.n100 vss 1.00fF $ **FLOATING
C108 vp_n.n102 vss 1.00fF $ **FLOATING
C109 vp_n.n104 vss 1.00fF $ **FLOATING
C110 vp_n.n106 vss 1.00fF $ **FLOATING
C111 vp_n.n108 vss 1.00fF $ **FLOATING
C112 vp_n.n110 vss 1.00fF $ **FLOATING
C113 vp_n.n112 vss 1.00fF $ **FLOATING
C114 vp_n.n114 vss 1.00fF $ **FLOATING
C115 vp_n.n116 vss 1.00fF $ **FLOATING
C116 vp_n.n118 vss 1.00fF $ **FLOATING
C117 vp_n.n120 vss 1.00fF $ **FLOATING
C118 vp_n.n122 vss 1.00fF $ **FLOATING
C119 vp_n.n124 vss 1.00fF $ **FLOATING
C120 vp_n.n126 vss 1.00fF $ **FLOATING
C121 vp_n.n128 vss 1.00fF $ **FLOATING
C122 vp_n.n130 vss 1.00fF $ **FLOATING
C123 vp_n.n132 vss 1.00fF $ **FLOATING
C124 vp_n.n134 vss 1.00fF $ **FLOATING
C125 vp_n.n136 vss 1.00fF $ **FLOATING
C126 vp_n.n138 vss 1.00fF $ **FLOATING
C127 vp_n.n140 vss 1.00fF $ **FLOATING
C128 vp_n.n142 vss 1.00fF $ **FLOATING
C129 vp_n.n144 vss 1.00fF $ **FLOATING
C130 vp_n.n146 vss 1.00fF $ **FLOATING
C131 vp_n.n148 vss 1.00fF $ **FLOATING
C132 vp_n.n150 vss 1.00fF $ **FLOATING
C133 vp_n.n152 vss 1.00fF $ **FLOATING
C134 vp_n.n154 vss 1.00fF $ **FLOATING
C135 vp_n.n156 vss 1.00fF $ **FLOATING
C136 vp_n.n158 vss 1.00fF $ **FLOATING
C137 vp_n.n160 vss 1.00fF $ **FLOATING
C138 vp_n.n162 vss 1.00fF $ **FLOATING
C139 vp_n.n164 vss 1.00fF $ **FLOATING
C140 vp_n.n166 vss 1.00fF $ **FLOATING
C141 vp_n.n168 vss 1.00fF $ **FLOATING
C142 vp_n.n170 vss 1.00fF $ **FLOATING
C143 vp_n.n172 vss 1.00fF $ **FLOATING
C144 vp_n.n174 vss 1.00fF $ **FLOATING
C145 vp_n.n176 vss 1.00fF $ **FLOATING
C146 vp_n.n178 vss 1.00fF $ **FLOATING
C147 vp_n.n180 vss 1.00fF $ **FLOATING
C148 vp_n.n182 vss 1.00fF $ **FLOATING
C149 vp_n.n184 vss 1.00fF $ **FLOATING
C150 vp_n.n186 vss 1.00fF $ **FLOATING
C151 vp_n.n188 vss 1.00fF $ **FLOATING
C152 vp_n.n190 vss 1.00fF $ **FLOATING
C153 vp_n.n192 vss 1.00fF $ **FLOATING
C154 vp_n.n194 vss 1.00fF $ **FLOATING
C155 vp_n.n196 vss 1.00fF $ **FLOATING
C156 vp_n.n198 vss 1.00fF $ **FLOATING
C157 vp_n.n200 vss 1.00fF $ **FLOATING
C158 vp_n.n202 vss 1.00fF $ **FLOATING
C159 vp_n.n204 vss 1.00fF $ **FLOATING
C160 vp_n.n206 vss 1.00fF $ **FLOATING
C161 vp_n.n208 vss 1.00fF $ **FLOATING
C162 vp_n.n210 vss 1.00fF $ **FLOATING
C163 vp_n.n212 vss 1.00fF $ **FLOATING
C164 vp_n.n214 vss 1.00fF $ **FLOATING
C165 vp_n.n216 vss 1.00fF $ **FLOATING
C166 vp_n.n218 vss 1.00fF $ **FLOATING
C167 vp_n.n220 vss 1.00fF $ **FLOATING
C168 vp_n.n222 vss 1.06fF $ **FLOATING
C169 vp_n.n223 vss 1.16fF $ **FLOATING
C170 vp_n.n296 vss 1.58fF $ **FLOATING
C171 vp_n.n297 vss 12.55fF $ **FLOATING
C172 vdd1.n0 vss 4.27fF $ **FLOATING
C173 vdd1.n1 vss 4.48fF $ **FLOATING
C174 vdd1.n2 vss 4.48fF $ **FLOATING
C175 vdd1.n3 vss 4.48fF $ **FLOATING
C176 vdd1.n4 vss 4.59fF $ **FLOATING
C177 vdd1.n5 vss 4.60fF $ **FLOATING
C178 vdd1.n6 vss 4.48fF $ **FLOATING
C179 vdd1.n7 vss 4.48fF $ **FLOATING
C180 vdd1.n8 vss 4.48fF $ **FLOATING
C181 vdd1.n9 vss 4.08fF $ **FLOATING
C182 vdd1.n12 vss 13.99fF $ **FLOATING
C183 vdd1.n13 vss 5.53fF $ **FLOATING
C184 vdd1.n14 vss 5.53fF $ **FLOATING
C185 vdd1.n15 vss 6.46fF $ **FLOATING
C186 vdd1.n16 vss 6.46fF $ **FLOATING
C187 vdd1.n17 vss 11.77fF $ **FLOATING
C188 vdd1.n18 vss 13.99fF $ **FLOATING
C189 vdd1.n19 vss 5.52fF $ **FLOATING
C190 vdd1.n20 vss 5.52fF $ **FLOATING
C191 vdd1.n21 vss 6.44fF $ **FLOATING
C192 vdd1.n22 vss 6.44fF $ **FLOATING
C193 vdd1.n23 vss 11.77fF $ **FLOATING
C194 vdd1.n24 vss 6.53fF $ **FLOATING
C195 vdd1.n25 vss 33.04fF $ **FLOATING
C196 vdd1.n27 vss 4.27fF $ **FLOATING
C197 vdd1.n28 vss 4.48fF $ **FLOATING
C198 vdd1.n29 vss 4.48fF $ **FLOATING
C199 vdd1.n30 vss 4.48fF $ **FLOATING
C200 vdd1.n31 vss 4.59fF $ **FLOATING
C201 vdd1.n32 vss 4.60fF $ **FLOATING
C202 vdd1.n33 vss 4.48fF $ **FLOATING
C203 vdd1.n34 vss 4.48fF $ **FLOATING
C204 vdd1.n35 vss 4.48fF $ **FLOATING
C205 vdd1.n36 vss 4.08fF $ **FLOATING
C206 vdd1.n38 vss 5.75fF $ **FLOATING
C207 vdd1.n39 vss 3.09fF $ **FLOATING
C208 vdd1.n40 vss 3.09fF $ **FLOATING
C209 vdd1.n41 vss 3.13fF $ **FLOATING
C210 vdd1.n42 vss 3.19fF $ **FLOATING
C211 vdd1.n43 vss 3.09fF $ **FLOATING
C212 vdd1.n44 vss 3.09fF $ **FLOATING
C213 vdd1.n45 vss 3.09fF $ **FLOATING
C214 vdd1.n46 vss 2.61fF $ **FLOATING
C215 vdd1.n47 vss 4.27fF $ **FLOATING
C216 vdd1.n48 vss 4.48fF $ **FLOATING
C217 vdd1.n49 vss 4.48fF $ **FLOATING
C218 vdd1.n50 vss 4.48fF $ **FLOATING
C219 vdd1.n51 vss 4.59fF $ **FLOATING
C220 vdd1.n52 vss 4.60fF $ **FLOATING
C221 vdd1.n53 vss 4.48fF $ **FLOATING
C222 vdd1.n54 vss 4.48fF $ **FLOATING
C223 vdd1.n55 vss 4.48fF $ **FLOATING
C224 vdd1.n56 vss 4.08fF $ **FLOATING
C225 vdd1.n57 vss 11.29fF $ **FLOATING
C226 vdd1.n58 vss 4.27fF $ **FLOATING
C227 vdd1.n59 vss 4.48fF $ **FLOATING
C228 vdd1.n60 vss 4.48fF $ **FLOATING
C229 vdd1.n61 vss 4.48fF $ **FLOATING
C230 vdd1.n62 vss 4.59fF $ **FLOATING
C231 vdd1.n63 vss 4.60fF $ **FLOATING
C232 vdd1.n64 vss 4.48fF $ **FLOATING
C233 vdd1.n65 vss 4.48fF $ **FLOATING
C234 vdd1.n66 vss 4.48fF $ **FLOATING
C235 vdd1.n67 vss 4.08fF $ **FLOATING
C236 vdd1.n68 vss 32.35fF $ **FLOATING
C237 vdd1.n69 vss 4.27fF $ **FLOATING
C238 vdd1.n70 vss 4.48fF $ **FLOATING
C239 vdd1.n71 vss 4.48fF $ **FLOATING
C240 vdd1.n72 vss 4.48fF $ **FLOATING
C241 vdd1.n73 vss 4.59fF $ **FLOATING
C242 vdd1.n74 vss 4.60fF $ **FLOATING
C243 vdd1.n75 vss 4.48fF $ **FLOATING
C244 vdd1.n76 vss 4.48fF $ **FLOATING
C245 vdd1.n77 vss 4.48fF $ **FLOATING
C246 vdd1.n78 vss 4.08fF $ **FLOATING
C247 vdd1.n79 vss 34.58fF $ **FLOATING
C248 vdd1.n80 vss 4.27fF $ **FLOATING
C249 vdd1.n81 vss 4.48fF $ **FLOATING
C250 vdd1.n82 vss 4.48fF $ **FLOATING
C251 vdd1.n83 vss 4.48fF $ **FLOATING
C252 vdd1.n84 vss 4.59fF $ **FLOATING
C253 vdd1.n85 vss 4.60fF $ **FLOATING
C254 vdd1.n86 vss 4.48fF $ **FLOATING
C255 vdd1.n87 vss 4.48fF $ **FLOATING
C256 vdd1.n88 vss 4.48fF $ **FLOATING
C257 vdd1.n89 vss 4.08fF $ **FLOATING
C258 vdd1.n90 vss 34.58fF $ **FLOATING
C259 vdd1.n91 vss 4.27fF $ **FLOATING
C260 vdd1.n92 vss 4.48fF $ **FLOATING
C261 vdd1.n93 vss 4.48fF $ **FLOATING
C262 vdd1.n94 vss 4.48fF $ **FLOATING
C263 vdd1.n95 vss 4.59fF $ **FLOATING
C264 vdd1.n96 vss 4.60fF $ **FLOATING
C265 vdd1.n97 vss 4.48fF $ **FLOATING
C266 vdd1.n98 vss 4.48fF $ **FLOATING
C267 vdd1.n99 vss 4.48fF $ **FLOATING
C268 vdd1.n100 vss 4.08fF $ **FLOATING
C269 vdd1.n101 vss 34.58fF $ **FLOATING
C270 vdd1.n102 vss 4.27fF $ **FLOATING
C271 vdd1.n103 vss 4.48fF $ **FLOATING
C272 vdd1.n104 vss 4.48fF $ **FLOATING
C273 vdd1.n105 vss 4.48fF $ **FLOATING
C274 vdd1.n106 vss 4.59fF $ **FLOATING
C275 vdd1.n107 vss 4.60fF $ **FLOATING
C276 vdd1.n108 vss 4.48fF $ **FLOATING
C277 vdd1.n109 vss 4.48fF $ **FLOATING
C278 vdd1.n110 vss 4.48fF $ **FLOATING
C279 vdd1.n111 vss 4.08fF $ **FLOATING
C280 vdd1.n112 vss 34.58fF $ **FLOATING
C281 vdd1.n113 vss 4.27fF $ **FLOATING
C282 vdd1.n114 vss 4.48fF $ **FLOATING
C283 vdd1.n115 vss 4.48fF $ **FLOATING
C284 vdd1.n116 vss 4.48fF $ **FLOATING
C285 vdd1.n117 vss 4.59fF $ **FLOATING
C286 vdd1.n118 vss 4.60fF $ **FLOATING
C287 vdd1.n119 vss 4.48fF $ **FLOATING
C288 vdd1.n120 vss 4.48fF $ **FLOATING
C289 vdd1.n121 vss 4.48fF $ **FLOATING
C290 vdd1.n122 vss 4.08fF $ **FLOATING
C291 vdd1.n123 vss 34.58fF $ **FLOATING
C292 vdd1.n124 vss 4.27fF $ **FLOATING
C293 vdd1.n125 vss 4.48fF $ **FLOATING
C294 vdd1.n126 vss 4.48fF $ **FLOATING
C295 vdd1.n127 vss 4.48fF $ **FLOATING
C296 vdd1.n128 vss 4.59fF $ **FLOATING
C297 vdd1.n129 vss 4.60fF $ **FLOATING
C298 vdd1.n130 vss 4.48fF $ **FLOATING
C299 vdd1.n131 vss 4.48fF $ **FLOATING
C300 vdd1.n132 vss 4.48fF $ **FLOATING
C301 vdd1.n133 vss 4.08fF $ **FLOATING
C302 vdd1.n134 vss 34.58fF $ **FLOATING
C303 vdd1.n135 vss 4.27fF $ **FLOATING
C304 vdd1.n136 vss 4.48fF $ **FLOATING
C305 vdd1.n137 vss 4.48fF $ **FLOATING
C306 vdd1.n138 vss 4.48fF $ **FLOATING
C307 vdd1.n139 vss 4.59fF $ **FLOATING
C308 vdd1.n140 vss 4.60fF $ **FLOATING
C309 vdd1.n141 vss 4.48fF $ **FLOATING
C310 vdd1.n142 vss 4.48fF $ **FLOATING
C311 vdd1.n143 vss 4.48fF $ **FLOATING
C312 vdd1.n144 vss 4.08fF $ **FLOATING
C313 vdd1.n145 vss 34.58fF $ **FLOATING
C314 vdd1.n146 vss 4.27fF $ **FLOATING
C315 vdd1.n147 vss 4.48fF $ **FLOATING
C316 vdd1.n148 vss 4.48fF $ **FLOATING
C317 vdd1.n149 vss 4.48fF $ **FLOATING
C318 vdd1.n150 vss 4.59fF $ **FLOATING
C319 vdd1.n151 vss 4.60fF $ **FLOATING
C320 vdd1.n152 vss 4.48fF $ **FLOATING
C321 vdd1.n153 vss 4.48fF $ **FLOATING
C322 vdd1.n154 vss 4.48fF $ **FLOATING
C323 vdd1.n155 vss 4.08fF $ **FLOATING
C324 vdd1.n156 vss 34.58fF $ **FLOATING
C325 vdd1.n157 vss 4.27fF $ **FLOATING
C326 vdd1.n158 vss 4.48fF $ **FLOATING
C327 vdd1.n159 vss 4.48fF $ **FLOATING
C328 vdd1.n160 vss 4.48fF $ **FLOATING
C329 vdd1.n161 vss 4.59fF $ **FLOATING
C330 vdd1.n162 vss 4.60fF $ **FLOATING
C331 vdd1.n163 vss 4.48fF $ **FLOATING
C332 vdd1.n164 vss 4.48fF $ **FLOATING
C333 vdd1.n165 vss 4.48fF $ **FLOATING
C334 vdd1.n166 vss 4.08fF $ **FLOATING
C335 vdd1.n167 vss 34.58fF $ **FLOATING
C336 vdd1.n168 vss 4.27fF $ **FLOATING
C337 vdd1.n169 vss 4.48fF $ **FLOATING
C338 vdd1.n170 vss 4.48fF $ **FLOATING
C339 vdd1.n171 vss 4.48fF $ **FLOATING
C340 vdd1.n172 vss 4.59fF $ **FLOATING
C341 vdd1.n173 vss 4.60fF $ **FLOATING
C342 vdd1.n174 vss 4.48fF $ **FLOATING
C343 vdd1.n175 vss 4.48fF $ **FLOATING
C344 vdd1.n176 vss 4.48fF $ **FLOATING
C345 vdd1.n177 vss 4.08fF $ **FLOATING
C346 vdd1.n178 vss 34.58fF $ **FLOATING
C347 vdd1.n179 vss 4.27fF $ **FLOATING
C348 vdd1.n180 vss 4.48fF $ **FLOATING
C349 vdd1.n181 vss 4.48fF $ **FLOATING
C350 vdd1.n182 vss 4.48fF $ **FLOATING
C351 vdd1.n183 vss 4.59fF $ **FLOATING
C352 vdd1.n184 vss 4.60fF $ **FLOATING
C353 vdd1.n185 vss 4.48fF $ **FLOATING
C354 vdd1.n186 vss 4.48fF $ **FLOATING
C355 vdd1.n187 vss 4.48fF $ **FLOATING
C356 vdd1.n188 vss 4.08fF $ **FLOATING
C357 vdd1.n189 vss 34.58fF $ **FLOATING
C358 vdd1.n190 vss 4.27fF $ **FLOATING
C359 vdd1.n191 vss 4.48fF $ **FLOATING
C360 vdd1.n192 vss 4.48fF $ **FLOATING
C361 vdd1.n193 vss 4.48fF $ **FLOATING
C362 vdd1.n194 vss 4.59fF $ **FLOATING
C363 vdd1.n195 vss 4.60fF $ **FLOATING
C364 vdd1.n196 vss 4.48fF $ **FLOATING
C365 vdd1.n197 vss 4.48fF $ **FLOATING
C366 vdd1.n198 vss 4.48fF $ **FLOATING
C367 vdd1.n199 vss 4.08fF $ **FLOATING
C368 vdd1.n200 vss 34.58fF $ **FLOATING
C369 vdd1.n201 vss 4.27fF $ **FLOATING
C370 vdd1.n202 vss 4.48fF $ **FLOATING
C371 vdd1.n203 vss 4.48fF $ **FLOATING
C372 vdd1.n204 vss 4.48fF $ **FLOATING
C373 vdd1.n205 vss 4.59fF $ **FLOATING
C374 vdd1.n206 vss 4.60fF $ **FLOATING
C375 vdd1.n207 vss 4.48fF $ **FLOATING
C376 vdd1.n208 vss 4.48fF $ **FLOATING
C377 vdd1.n209 vss 4.48fF $ **FLOATING
C378 vdd1.n210 vss 4.08fF $ **FLOATING
C379 vdd1.n211 vss 34.58fF $ **FLOATING
C380 vdd1.n212 vss 4.27fF $ **FLOATING
C381 vdd1.n213 vss 4.48fF $ **FLOATING
C382 vdd1.n214 vss 4.48fF $ **FLOATING
C383 vdd1.n215 vss 4.48fF $ **FLOATING
C384 vdd1.n216 vss 4.59fF $ **FLOATING
C385 vdd1.n217 vss 4.60fF $ **FLOATING
C386 vdd1.n218 vss 4.48fF $ **FLOATING
C387 vdd1.n219 vss 4.48fF $ **FLOATING
C388 vdd1.n220 vss 4.48fF $ **FLOATING
C389 vdd1.n221 vss 4.08fF $ **FLOATING
C390 vdd1.n222 vss 34.58fF $ **FLOATING
C391 vdd1.n223 vss 4.27fF $ **FLOATING
C392 vdd1.n224 vss 4.48fF $ **FLOATING
C393 vdd1.n225 vss 4.48fF $ **FLOATING
C394 vdd1.n226 vss 4.48fF $ **FLOATING
C395 vdd1.n227 vss 4.59fF $ **FLOATING
C396 vdd1.n228 vss 4.60fF $ **FLOATING
C397 vdd1.n229 vss 4.48fF $ **FLOATING
C398 vdd1.n230 vss 4.48fF $ **FLOATING
C399 vdd1.n231 vss 4.48fF $ **FLOATING
C400 vdd1.n232 vss 4.08fF $ **FLOATING
C401 vdd1.n233 vss 34.58fF $ **FLOATING
C402 vdd1.n234 vss 4.27fF $ **FLOATING
C403 vdd1.n235 vss 4.48fF $ **FLOATING
C404 vdd1.n236 vss 4.48fF $ **FLOATING
C405 vdd1.n237 vss 4.48fF $ **FLOATING
C406 vdd1.n238 vss 4.59fF $ **FLOATING
C407 vdd1.n239 vss 4.60fF $ **FLOATING
C408 vdd1.n240 vss 4.48fF $ **FLOATING
C409 vdd1.n241 vss 4.48fF $ **FLOATING
C410 vdd1.n242 vss 4.48fF $ **FLOATING
C411 vdd1.n243 vss 4.08fF $ **FLOATING
C412 vdd1.n244 vss 34.58fF $ **FLOATING
C413 vdd1.n245 vss 4.27fF $ **FLOATING
C414 vdd1.n246 vss 4.48fF $ **FLOATING
C415 vdd1.n247 vss 4.48fF $ **FLOATING
C416 vdd1.n248 vss 4.48fF $ **FLOATING
C417 vdd1.n249 vss 4.59fF $ **FLOATING
C418 vdd1.n250 vss 4.60fF $ **FLOATING
C419 vdd1.n251 vss 4.48fF $ **FLOATING
C420 vdd1.n252 vss 4.48fF $ **FLOATING
C421 vdd1.n253 vss 4.48fF $ **FLOATING
C422 vdd1.n254 vss 4.08fF $ **FLOATING
C423 vdd1.n255 vss 34.58fF $ **FLOATING
C424 vdd1.n256 vss 4.27fF $ **FLOATING
C425 vdd1.n257 vss 4.48fF $ **FLOATING
C426 vdd1.n258 vss 4.48fF $ **FLOATING
C427 vdd1.n259 vss 4.48fF $ **FLOATING
C428 vdd1.n260 vss 4.59fF $ **FLOATING
C429 vdd1.n261 vss 4.60fF $ **FLOATING
C430 vdd1.n262 vss 4.48fF $ **FLOATING
C431 vdd1.n263 vss 4.48fF $ **FLOATING
C432 vdd1.n264 vss 4.48fF $ **FLOATING
C433 vdd1.n265 vss 4.08fF $ **FLOATING
C434 vdd1.n266 vss 34.58fF $ **FLOATING
C435 vdd1.n267 vss 4.27fF $ **FLOATING
C436 vdd1.n268 vss 4.48fF $ **FLOATING
C437 vdd1.n269 vss 4.48fF $ **FLOATING
C438 vdd1.n270 vss 4.48fF $ **FLOATING
C439 vdd1.n271 vss 4.59fF $ **FLOATING
C440 vdd1.n272 vss 4.60fF $ **FLOATING
C441 vdd1.n273 vss 4.48fF $ **FLOATING
C442 vdd1.n274 vss 4.48fF $ **FLOATING
C443 vdd1.n275 vss 4.48fF $ **FLOATING
C444 vdd1.n276 vss 4.08fF $ **FLOATING
C445 vdd1.n277 vss 34.58fF $ **FLOATING
C446 vdd1.n278 vss 4.27fF $ **FLOATING
C447 vdd1.n279 vss 4.48fF $ **FLOATING
C448 vdd1.n280 vss 4.48fF $ **FLOATING
C449 vdd1.n281 vss 4.48fF $ **FLOATING
C450 vdd1.n282 vss 4.59fF $ **FLOATING
C451 vdd1.n283 vss 4.60fF $ **FLOATING
C452 vdd1.n284 vss 4.48fF $ **FLOATING
C453 vdd1.n285 vss 4.48fF $ **FLOATING
C454 vdd1.n286 vss 4.48fF $ **FLOATING
C455 vdd1.n287 vss 4.08fF $ **FLOATING
C456 vdd1.n288 vss 34.58fF $ **FLOATING
C457 vdd1.n289 vss 4.27fF $ **FLOATING
C458 vdd1.n290 vss 4.48fF $ **FLOATING
C459 vdd1.n291 vss 4.48fF $ **FLOATING
C460 vdd1.n292 vss 4.48fF $ **FLOATING
C461 vdd1.n293 vss 4.59fF $ **FLOATING
C462 vdd1.n294 vss 4.60fF $ **FLOATING
C463 vdd1.n295 vss 4.48fF $ **FLOATING
C464 vdd1.n296 vss 4.48fF $ **FLOATING
C465 vdd1.n297 vss 4.48fF $ **FLOATING
C466 vdd1.n298 vss 4.08fF $ **FLOATING
C467 vdd1.n299 vss 34.58fF $ **FLOATING
C468 vdd1.n300 vss 4.27fF $ **FLOATING
C469 vdd1.n301 vss 4.48fF $ **FLOATING
C470 vdd1.n302 vss 4.48fF $ **FLOATING
C471 vdd1.n303 vss 4.48fF $ **FLOATING
C472 vdd1.n304 vss 4.59fF $ **FLOATING
C473 vdd1.n305 vss 4.60fF $ **FLOATING
C474 vdd1.n306 vss 4.48fF $ **FLOATING
C475 vdd1.n307 vss 4.48fF $ **FLOATING
C476 vdd1.n308 vss 4.48fF $ **FLOATING
C477 vdd1.n309 vss 4.08fF $ **FLOATING
C478 vdd1.n310 vss 34.58fF $ **FLOATING
C479 vdd1.n311 vss 4.27fF $ **FLOATING
C480 vdd1.n312 vss 4.48fF $ **FLOATING
C481 vdd1.n313 vss 4.48fF $ **FLOATING
C482 vdd1.n314 vss 4.48fF $ **FLOATING
C483 vdd1.n315 vss 4.59fF $ **FLOATING
C484 vdd1.n316 vss 4.60fF $ **FLOATING
C485 vdd1.n317 vss 4.48fF $ **FLOATING
C486 vdd1.n318 vss 4.48fF $ **FLOATING
C487 vdd1.n319 vss 4.48fF $ **FLOATING
C488 vdd1.n320 vss 4.08fF $ **FLOATING
C489 vdd1.n321 vss 5.32fF $ **FLOATING
C490 vdd1.n322 vss 33.29fF $ **FLOATING
C491 vdd1.n323 vss 4.27fF $ **FLOATING
C492 vdd1.n324 vss 4.48fF $ **FLOATING
C493 vdd1.n325 vss 4.48fF $ **FLOATING
C494 vdd1.n326 vss 4.48fF $ **FLOATING
C495 vdd1.n327 vss 4.59fF $ **FLOATING
C496 vdd1.n328 vss 4.60fF $ **FLOATING
C497 vdd1.n329 vss 4.48fF $ **FLOATING
C498 vdd1.n330 vss 4.48fF $ **FLOATING
C499 vdd1.n331 vss 4.48fF $ **FLOATING
C500 vdd1.n332 vss 4.08fF $ **FLOATING
C501 vdd1.n333 vss 28.31fF $ **FLOATING
C502 vdd1.n334 vss 4.27fF $ **FLOATING
C503 vdd1.n335 vss 4.48fF $ **FLOATING
C504 vdd1.n336 vss 4.48fF $ **FLOATING
C505 vdd1.n337 vss 4.48fF $ **FLOATING
C506 vdd1.n338 vss 4.59fF $ **FLOATING
C507 vdd1.n339 vss 4.60fF $ **FLOATING
C508 vdd1.n340 vss 4.48fF $ **FLOATING
C509 vdd1.n341 vss 4.48fF $ **FLOATING
C510 vdd1.n342 vss 4.48fF $ **FLOATING
C511 vdd1.n343 vss 4.08fF $ **FLOATING
C512 vdd1.n344 vss 34.29fF $ **FLOATING
C513 vdd1.n345 vss 4.27fF $ **FLOATING
C514 vdd1.n346 vss 4.48fF $ **FLOATING
C515 vdd1.n347 vss 4.48fF $ **FLOATING
C516 vdd1.n348 vss 4.48fF $ **FLOATING
C517 vdd1.n349 vss 4.59fF $ **FLOATING
C518 vdd1.n350 vss 4.60fF $ **FLOATING
C519 vdd1.n351 vss 4.48fF $ **FLOATING
C520 vdd1.n352 vss 4.48fF $ **FLOATING
C521 vdd1.n353 vss 4.48fF $ **FLOATING
C522 vdd1.n354 vss 4.08fF $ **FLOATING
C523 vdd1.n355 vss 34.58fF $ **FLOATING
C524 vdd1.n356 vss 4.27fF $ **FLOATING
C525 vdd1.n357 vss 4.48fF $ **FLOATING
C526 vdd1.n358 vss 4.48fF $ **FLOATING
C527 vdd1.n359 vss 4.48fF $ **FLOATING
C528 vdd1.n360 vss 4.59fF $ **FLOATING
C529 vdd1.n361 vss 4.60fF $ **FLOATING
C530 vdd1.n362 vss 4.48fF $ **FLOATING
C531 vdd1.n363 vss 4.48fF $ **FLOATING
C532 vdd1.n364 vss 4.48fF $ **FLOATING
C533 vdd1.n365 vss 4.08fF $ **FLOATING
C534 vdd1.n366 vss 34.58fF $ **FLOATING
C535 vdd1.n367 vss 4.27fF $ **FLOATING
C536 vdd1.n368 vss 4.48fF $ **FLOATING
C537 vdd1.n369 vss 4.48fF $ **FLOATING
C538 vdd1.n370 vss 4.48fF $ **FLOATING
C539 vdd1.n371 vss 4.59fF $ **FLOATING
C540 vdd1.n372 vss 4.60fF $ **FLOATING
C541 vdd1.n373 vss 4.48fF $ **FLOATING
C542 vdd1.n374 vss 4.48fF $ **FLOATING
C543 vdd1.n375 vss 4.48fF $ **FLOATING
C544 vdd1.n376 vss 4.08fF $ **FLOATING
C545 vdd1.n377 vss 34.58fF $ **FLOATING
C546 vdd1.n378 vss 4.27fF $ **FLOATING
C547 vdd1.n379 vss 4.48fF $ **FLOATING
C548 vdd1.n380 vss 4.48fF $ **FLOATING
C549 vdd1.n381 vss 4.48fF $ **FLOATING
C550 vdd1.n382 vss 4.59fF $ **FLOATING
C551 vdd1.n383 vss 4.60fF $ **FLOATING
C552 vdd1.n384 vss 4.48fF $ **FLOATING
C553 vdd1.n385 vss 4.48fF $ **FLOATING
C554 vdd1.n386 vss 4.48fF $ **FLOATING
C555 vdd1.n387 vss 4.08fF $ **FLOATING
C556 vdd1.n388 vss 34.58fF $ **FLOATING
C557 vdd1.n389 vss 4.27fF $ **FLOATING
C558 vdd1.n390 vss 4.48fF $ **FLOATING
C559 vdd1.n391 vss 4.48fF $ **FLOATING
C560 vdd1.n392 vss 4.48fF $ **FLOATING
C561 vdd1.n393 vss 4.59fF $ **FLOATING
C562 vdd1.n394 vss 4.60fF $ **FLOATING
C563 vdd1.n395 vss 4.48fF $ **FLOATING
C564 vdd1.n396 vss 4.48fF $ **FLOATING
C565 vdd1.n397 vss 4.48fF $ **FLOATING
C566 vdd1.n398 vss 4.08fF $ **FLOATING
C567 vdd1.n399 vss 34.58fF $ **FLOATING
C568 vdd1.n400 vss 4.27fF $ **FLOATING
C569 vdd1.n401 vss 4.48fF $ **FLOATING
C570 vdd1.n402 vss 4.48fF $ **FLOATING
C571 vdd1.n403 vss 4.48fF $ **FLOATING
C572 vdd1.n404 vss 4.59fF $ **FLOATING
C573 vdd1.n405 vss 4.60fF $ **FLOATING
C574 vdd1.n406 vss 4.48fF $ **FLOATING
C575 vdd1.n407 vss 4.48fF $ **FLOATING
C576 vdd1.n408 vss 4.48fF $ **FLOATING
C577 vdd1.n409 vss 4.08fF $ **FLOATING
C578 vdd1.n410 vss 34.58fF $ **FLOATING
C579 vdd1.n411 vss 4.27fF $ **FLOATING
C580 vdd1.n412 vss 4.48fF $ **FLOATING
C581 vdd1.n413 vss 4.48fF $ **FLOATING
C582 vdd1.n414 vss 4.48fF $ **FLOATING
C583 vdd1.n415 vss 4.59fF $ **FLOATING
C584 vdd1.n416 vss 4.60fF $ **FLOATING
C585 vdd1.n417 vss 4.48fF $ **FLOATING
C586 vdd1.n418 vss 4.48fF $ **FLOATING
C587 vdd1.n419 vss 4.48fF $ **FLOATING
C588 vdd1.n420 vss 4.08fF $ **FLOATING
C589 vdd1.n421 vss 34.58fF $ **FLOATING
C590 vdd1.n422 vss 4.27fF $ **FLOATING
C591 vdd1.n423 vss 4.48fF $ **FLOATING
C592 vdd1.n424 vss 4.48fF $ **FLOATING
C593 vdd1.n425 vss 4.48fF $ **FLOATING
C594 vdd1.n426 vss 4.59fF $ **FLOATING
C595 vdd1.n427 vss 4.60fF $ **FLOATING
C596 vdd1.n428 vss 4.48fF $ **FLOATING
C597 vdd1.n429 vss 4.48fF $ **FLOATING
C598 vdd1.n430 vss 4.48fF $ **FLOATING
C599 vdd1.n431 vss 4.08fF $ **FLOATING
C600 vdd1.n432 vss 34.58fF $ **FLOATING
C601 vdd1.n433 vss 4.27fF $ **FLOATING
C602 vdd1.n434 vss 4.48fF $ **FLOATING
C603 vdd1.n435 vss 4.48fF $ **FLOATING
C604 vdd1.n436 vss 4.48fF $ **FLOATING
C605 vdd1.n437 vss 4.59fF $ **FLOATING
C606 vdd1.n438 vss 4.60fF $ **FLOATING
C607 vdd1.n439 vss 4.48fF $ **FLOATING
C608 vdd1.n440 vss 4.48fF $ **FLOATING
C609 vdd1.n441 vss 4.48fF $ **FLOATING
C610 vdd1.n442 vss 4.08fF $ **FLOATING
C611 vdd1.n443 vss 5.32fF $ **FLOATING
C612 vdd1.n444 vss 33.29fF $ **FLOATING
C613 vdd1.n445 vss 4.27fF $ **FLOATING
C614 vdd1.n446 vss 4.48fF $ **FLOATING
C615 vdd1.n447 vss 4.48fF $ **FLOATING
C616 vdd1.n448 vss 4.48fF $ **FLOATING
C617 vdd1.n449 vss 4.59fF $ **FLOATING
C618 vdd1.n450 vss 4.60fF $ **FLOATING
C619 vdd1.n451 vss 4.48fF $ **FLOATING
C620 vdd1.n452 vss 4.48fF $ **FLOATING
C621 vdd1.n453 vss 4.48fF $ **FLOATING
C622 vdd1.n454 vss 4.08fF $ **FLOATING
C623 vdd1.n456 vss 33.55fF $ **FLOATING
C624 vdd1.n457 vss 4.27fF $ **FLOATING
C625 vdd1.n458 vss 4.48fF $ **FLOATING
C626 vdd1.n459 vss 4.48fF $ **FLOATING
C627 vdd1.n460 vss 4.48fF $ **FLOATING
C628 vdd1.n461 vss 4.59fF $ **FLOATING
C629 vdd1.n462 vss 4.60fF $ **FLOATING
C630 vdd1.n463 vss 4.48fF $ **FLOATING
C631 vdd1.n464 vss 4.48fF $ **FLOATING
C632 vdd1.n465 vss 4.48fF $ **FLOATING
C633 vdd1.n466 vss 4.08fF $ **FLOATING
C634 vdd1.n467 vss 30.28fF $ **FLOATING
C635 vdd1.n468 vss 4.27fF $ **FLOATING
C636 vdd1.n469 vss 4.48fF $ **FLOATING
C637 vdd1.n470 vss 4.48fF $ **FLOATING
C638 vdd1.n471 vss 4.48fF $ **FLOATING
C639 vdd1.n472 vss 4.59fF $ **FLOATING
C640 vdd1.n473 vss 4.60fF $ **FLOATING
C641 vdd1.n474 vss 4.48fF $ **FLOATING
C642 vdd1.n475 vss 4.48fF $ **FLOATING
C643 vdd1.n476 vss 4.48fF $ **FLOATING
C644 vdd1.n477 vss 4.08fF $ **FLOATING
C645 vdd1.n478 vss 34.58fF $ **FLOATING
C646 vdd1.n479 vss 4.27fF $ **FLOATING
C647 vdd1.n480 vss 4.48fF $ **FLOATING
C648 vdd1.n481 vss 4.48fF $ **FLOATING
C649 vdd1.n482 vss 4.48fF $ **FLOATING
C650 vdd1.n483 vss 4.59fF $ **FLOATING
C651 vdd1.n484 vss 4.60fF $ **FLOATING
C652 vdd1.n485 vss 4.48fF $ **FLOATING
C653 vdd1.n486 vss 4.48fF $ **FLOATING
C654 vdd1.n487 vss 4.48fF $ **FLOATING
C655 vdd1.n488 vss 4.08fF $ **FLOATING
C656 vdd1.n489 vss 5.32fF $ **FLOATING
C657 vdd1.n490 vss 33.29fF $ **FLOATING
C658 vdd1.n491 vss 3.34fF $ **FLOATING
C659 vdd1.n492 vss 1.90fF $ **FLOATING
C660 vdd1.n493 vss 1.90fF $ **FLOATING
C661 vdd1.n494 vss 1.94fF $ **FLOATING
C662 vdd1.n495 vss 1.99fF $ **FLOATING
C663 vdd1.n496 vss 1.95fF $ **FLOATING
C664 vdd1.n497 vss 1.95fF $ **FLOATING
C665 vdd1.n498 vss 1.95fF $ **FLOATING
C666 vdd1.n499 vss 1.80fF $ **FLOATING
C667 vdd1.n501 vss 4.27fF $ **FLOATING
C668 vdd1.n502 vss 4.48fF $ **FLOATING
C669 vdd1.n503 vss 4.48fF $ **FLOATING
C670 vdd1.n504 vss 4.48fF $ **FLOATING
C671 vdd1.n505 vss 4.59fF $ **FLOATING
C672 vdd1.n506 vss 4.59fF $ **FLOATING
C673 vdd1.n507 vss 4.48fF $ **FLOATING
C674 vdd1.n508 vss 4.48fF $ **FLOATING
C675 vdd1.n509 vss 4.48fF $ **FLOATING
C676 vdd1.n510 vss 4.07fF $ **FLOATING
C677 vdd1.n512 vss 28.05fF $ **FLOATING
C678 vdd1.n513 vss 4.27fF $ **FLOATING
C679 vdd1.n514 vss 4.48fF $ **FLOATING
C680 vdd1.n515 vss 4.48fF $ **FLOATING
C681 vdd1.n516 vss 4.48fF $ **FLOATING
C682 vdd1.n517 vss 4.59fF $ **FLOATING
C683 vdd1.n518 vss 4.60fF $ **FLOATING
C684 vdd1.n519 vss 4.48fF $ **FLOATING
C685 vdd1.n520 vss 4.48fF $ **FLOATING
C686 vdd1.n521 vss 4.48fF $ **FLOATING
C687 vdd1.n522 vss 4.08fF $ **FLOATING
C688 vdd1.n526 vss 33.04fF $ **FLOATING
C689 vdd1.n529 vss 4.27fF $ **FLOATING
C690 vdd1.n530 vss 4.48fF $ **FLOATING
C691 vdd1.n531 vss 4.48fF $ **FLOATING
C692 vdd1.n532 vss 4.48fF $ **FLOATING
C693 vdd1.n533 vss 4.59fF $ **FLOATING
C694 vdd1.n534 vss 4.60fF $ **FLOATING
C695 vdd1.n535 vss 4.48fF $ **FLOATING
C696 vdd1.n536 vss 4.48fF $ **FLOATING
C697 vdd1.n537 vss 4.48fF $ **FLOATING
C698 vdd1.n538 vss 4.08fF $ **FLOATING
C699 vdd1.n540 vss 33.04fF $ **FLOATING
C700 vdd1.n541 vss 4.27fF $ **FLOATING
C701 vdd1.n542 vss 4.48fF $ **FLOATING
C702 vdd1.n543 vss 4.48fF $ **FLOATING
C703 vdd1.n544 vss 4.48fF $ **FLOATING
C704 vdd1.n545 vss 4.59fF $ **FLOATING
C705 vdd1.n546 vss 4.60fF $ **FLOATING
C706 vdd1.n547 vss 4.48fF $ **FLOATING
C707 vdd1.n548 vss 4.48fF $ **FLOATING
C708 vdd1.n549 vss 4.48fF $ **FLOATING
C709 vdd1.n550 vss 4.08fF $ **FLOATING
C710 vdd1.n554 vss 33.04fF $ **FLOATING
C711 vdd1.n557 vss 4.27fF $ **FLOATING
C712 vdd1.n558 vss 4.48fF $ **FLOATING
C713 vdd1.n559 vss 4.48fF $ **FLOATING
C714 vdd1.n560 vss 4.48fF $ **FLOATING
C715 vdd1.n561 vss 4.59fF $ **FLOATING
C716 vdd1.n562 vss 4.60fF $ **FLOATING
C717 vdd1.n563 vss 4.48fF $ **FLOATING
C718 vdd1.n564 vss 4.48fF $ **FLOATING
C719 vdd1.n565 vss 4.48fF $ **FLOATING
C720 vdd1.n566 vss 4.08fF $ **FLOATING
C721 vdd1.n568 vss 33.04fF $ **FLOATING
C722 vdd1.n569 vss 4.27fF $ **FLOATING
C723 vdd1.n570 vss 4.48fF $ **FLOATING
C724 vdd1.n571 vss 4.48fF $ **FLOATING
C725 vdd1.n572 vss 4.48fF $ **FLOATING
C726 vdd1.n573 vss 4.59fF $ **FLOATING
C727 vdd1.n574 vss 4.60fF $ **FLOATING
C728 vdd1.n575 vss 4.48fF $ **FLOATING
C729 vdd1.n576 vss 4.48fF $ **FLOATING
C730 vdd1.n577 vss 4.48fF $ **FLOATING
C731 vdd1.n578 vss 4.08fF $ **FLOATING
C732 vdd1.n582 vss 33.04fF $ **FLOATING
C733 vdd1.n585 vss 4.27fF $ **FLOATING
C734 vdd1.n586 vss 4.48fF $ **FLOATING
C735 vdd1.n587 vss 4.48fF $ **FLOATING
C736 vdd1.n588 vss 4.48fF $ **FLOATING
C737 vdd1.n589 vss 4.59fF $ **FLOATING
C738 vdd1.n590 vss 4.60fF $ **FLOATING
C739 vdd1.n591 vss 4.48fF $ **FLOATING
C740 vdd1.n592 vss 4.48fF $ **FLOATING
C741 vdd1.n593 vss 4.48fF $ **FLOATING
C742 vdd1.n594 vss 4.08fF $ **FLOATING
C743 vdd1.n596 vss 33.04fF $ **FLOATING
C744 vdd1.n597 vss 4.27fF $ **FLOATING
C745 vdd1.n598 vss 4.48fF $ **FLOATING
C746 vdd1.n599 vss 4.48fF $ **FLOATING
C747 vdd1.n600 vss 4.48fF $ **FLOATING
C748 vdd1.n601 vss 4.59fF $ **FLOATING
C749 vdd1.n602 vss 4.60fF $ **FLOATING
C750 vdd1.n603 vss 4.48fF $ **FLOATING
C751 vdd1.n604 vss 4.48fF $ **FLOATING
C752 vdd1.n605 vss 4.48fF $ **FLOATING
C753 vdd1.n606 vss 4.08fF $ **FLOATING
C754 vdd1.n610 vss 33.04fF $ **FLOATING
C755 vdd1.n613 vss 4.27fF $ **FLOATING
C756 vdd1.n614 vss 4.48fF $ **FLOATING
C757 vdd1.n615 vss 4.48fF $ **FLOATING
C758 vdd1.n616 vss 4.48fF $ **FLOATING
C759 vdd1.n617 vss 4.59fF $ **FLOATING
C760 vdd1.n618 vss 4.60fF $ **FLOATING
C761 vdd1.n619 vss 4.48fF $ **FLOATING
C762 vdd1.n620 vss 4.48fF $ **FLOATING
C763 vdd1.n621 vss 4.48fF $ **FLOATING
C764 vdd1.n622 vss 4.08fF $ **FLOATING
C765 vdd1.n624 vss 33.04fF $ **FLOATING
C766 vdd1.n625 vss 4.27fF $ **FLOATING
C767 vdd1.n626 vss 4.48fF $ **FLOATING
C768 vdd1.n627 vss 4.48fF $ **FLOATING
C769 vdd1.n628 vss 4.48fF $ **FLOATING
C770 vdd1.n629 vss 4.59fF $ **FLOATING
C771 vdd1.n630 vss 4.60fF $ **FLOATING
C772 vdd1.n631 vss 4.48fF $ **FLOATING
C773 vdd1.n632 vss 4.48fF $ **FLOATING
C774 vdd1.n633 vss 4.48fF $ **FLOATING
C775 vdd1.n634 vss 4.08fF $ **FLOATING
C776 vdd1.n638 vss 33.04fF $ **FLOATING
C777 vdd1.n641 vss 4.27fF $ **FLOATING
C778 vdd1.n642 vss 4.48fF $ **FLOATING
C779 vdd1.n643 vss 4.48fF $ **FLOATING
C780 vdd1.n644 vss 4.48fF $ **FLOATING
C781 vdd1.n645 vss 4.59fF $ **FLOATING
C782 vdd1.n646 vss 4.60fF $ **FLOATING
C783 vdd1.n647 vss 4.48fF $ **FLOATING
C784 vdd1.n648 vss 4.48fF $ **FLOATING
C785 vdd1.n649 vss 4.48fF $ **FLOATING
C786 vdd1.n650 vss 4.08fF $ **FLOATING
C787 vdd1.n652 vss 33.04fF $ **FLOATING
C788 vdd1.n653 vss 4.27fF $ **FLOATING
C789 vdd1.n654 vss 4.48fF $ **FLOATING
C790 vdd1.n655 vss 4.48fF $ **FLOATING
C791 vdd1.n656 vss 4.48fF $ **FLOATING
C792 vdd1.n657 vss 4.59fF $ **FLOATING
C793 vdd1.n658 vss 4.60fF $ **FLOATING
C794 vdd1.n659 vss 4.48fF $ **FLOATING
C795 vdd1.n660 vss 4.48fF $ **FLOATING
C796 vdd1.n661 vss 4.48fF $ **FLOATING
C797 vdd1.n662 vss 4.08fF $ **FLOATING
C798 vdd1.n666 vss 33.04fF $ **FLOATING
C799 vdd1.n669 vss 4.27fF $ **FLOATING
C800 vdd1.n670 vss 4.48fF $ **FLOATING
C801 vdd1.n671 vss 4.48fF $ **FLOATING
C802 vdd1.n672 vss 4.48fF $ **FLOATING
C803 vdd1.n673 vss 4.59fF $ **FLOATING
C804 vdd1.n674 vss 4.60fF $ **FLOATING
C805 vdd1.n675 vss 4.48fF $ **FLOATING
C806 vdd1.n676 vss 4.48fF $ **FLOATING
C807 vdd1.n677 vss 4.48fF $ **FLOATING
C808 vdd1.n678 vss 4.08fF $ **FLOATING
C809 vdd1.n680 vss 33.04fF $ **FLOATING
C810 vdd1.n681 vss 4.27fF $ **FLOATING
C811 vdd1.n682 vss 4.48fF $ **FLOATING
C812 vdd1.n683 vss 4.48fF $ **FLOATING
C813 vdd1.n684 vss 4.48fF $ **FLOATING
C814 vdd1.n685 vss 4.59fF $ **FLOATING
C815 vdd1.n686 vss 4.60fF $ **FLOATING
C816 vdd1.n687 vss 4.48fF $ **FLOATING
C817 vdd1.n688 vss 4.48fF $ **FLOATING
C818 vdd1.n689 vss 4.48fF $ **FLOATING
C819 vdd1.n690 vss 4.08fF $ **FLOATING
C820 vdd1.n694 vss 33.04fF $ **FLOATING
C821 vdd1.n697 vss 4.27fF $ **FLOATING
C822 vdd1.n698 vss 4.48fF $ **FLOATING
C823 vdd1.n699 vss 4.48fF $ **FLOATING
C824 vdd1.n700 vss 4.48fF $ **FLOATING
C825 vdd1.n701 vss 4.59fF $ **FLOATING
C826 vdd1.n702 vss 4.60fF $ **FLOATING
C827 vdd1.n703 vss 4.48fF $ **FLOATING
C828 vdd1.n704 vss 4.48fF $ **FLOATING
C829 vdd1.n705 vss 4.48fF $ **FLOATING
C830 vdd1.n706 vss 4.08fF $ **FLOATING
C831 vdd1.n708 vss 33.04fF $ **FLOATING
C832 vdd1.n709 vss 4.27fF $ **FLOATING
C833 vdd1.n710 vss 4.48fF $ **FLOATING
C834 vdd1.n711 vss 4.48fF $ **FLOATING
C835 vdd1.n712 vss 4.48fF $ **FLOATING
C836 vdd1.n713 vss 4.59fF $ **FLOATING
C837 vdd1.n714 vss 4.60fF $ **FLOATING
C838 vdd1.n715 vss 4.48fF $ **FLOATING
C839 vdd1.n716 vss 4.48fF $ **FLOATING
C840 vdd1.n717 vss 4.48fF $ **FLOATING
C841 vdd1.n718 vss 4.08fF $ **FLOATING
C842 vdd1.n722 vss 33.04fF $ **FLOATING
C843 vdd1.n725 vss 4.27fF $ **FLOATING
C844 vdd1.n726 vss 4.48fF $ **FLOATING
C845 vdd1.n727 vss 4.48fF $ **FLOATING
C846 vdd1.n728 vss 4.48fF $ **FLOATING
C847 vdd1.n729 vss 4.59fF $ **FLOATING
C848 vdd1.n730 vss 4.60fF $ **FLOATING
C849 vdd1.n731 vss 4.48fF $ **FLOATING
C850 vdd1.n732 vss 4.48fF $ **FLOATING
C851 vdd1.n733 vss 4.48fF $ **FLOATING
C852 vdd1.n734 vss 4.08fF $ **FLOATING
C853 vdd1.n736 vss 33.04fF $ **FLOATING
C854 vdd1.n737 vss 4.27fF $ **FLOATING
C855 vdd1.n738 vss 4.48fF $ **FLOATING
C856 vdd1.n739 vss 4.48fF $ **FLOATING
C857 vdd1.n740 vss 4.48fF $ **FLOATING
C858 vdd1.n741 vss 4.59fF $ **FLOATING
C859 vdd1.n742 vss 4.60fF $ **FLOATING
C860 vdd1.n743 vss 4.48fF $ **FLOATING
C861 vdd1.n744 vss 4.48fF $ **FLOATING
C862 vdd1.n745 vss 4.48fF $ **FLOATING
C863 vdd1.n746 vss 4.08fF $ **FLOATING
C864 vdd1.n750 vss 33.04fF $ **FLOATING
C865 vdd1.n753 vss 4.27fF $ **FLOATING
C866 vdd1.n754 vss 4.48fF $ **FLOATING
C867 vdd1.n755 vss 4.48fF $ **FLOATING
C868 vdd1.n756 vss 4.48fF $ **FLOATING
C869 vdd1.n757 vss 4.59fF $ **FLOATING
C870 vdd1.n758 vss 4.60fF $ **FLOATING
C871 vdd1.n759 vss 4.48fF $ **FLOATING
C872 vdd1.n760 vss 4.48fF $ **FLOATING
C873 vdd1.n761 vss 4.48fF $ **FLOATING
C874 vdd1.n762 vss 4.08fF $ **FLOATING
C875 vdd1.n764 vss 33.04fF $ **FLOATING
C876 vdd1.n765 vss 4.27fF $ **FLOATING
C877 vdd1.n766 vss 4.48fF $ **FLOATING
C878 vdd1.n767 vss 4.48fF $ **FLOATING
C879 vdd1.n768 vss 4.48fF $ **FLOATING
C880 vdd1.n769 vss 4.59fF $ **FLOATING
C881 vdd1.n770 vss 4.60fF $ **FLOATING
C882 vdd1.n771 vss 4.48fF $ **FLOATING
C883 vdd1.n772 vss 4.48fF $ **FLOATING
C884 vdd1.n773 vss 4.48fF $ **FLOATING
C885 vdd1.n774 vss 4.08fF $ **FLOATING
C886 vdd1.n778 vss 33.04fF $ **FLOATING
C887 vdd1.n781 vss 4.27fF $ **FLOATING
C888 vdd1.n782 vss 4.48fF $ **FLOATING
C889 vdd1.n783 vss 4.48fF $ **FLOATING
C890 vdd1.n784 vss 4.48fF $ **FLOATING
C891 vdd1.n785 vss 4.59fF $ **FLOATING
C892 vdd1.n786 vss 4.60fF $ **FLOATING
C893 vdd1.n787 vss 4.48fF $ **FLOATING
C894 vdd1.n788 vss 4.48fF $ **FLOATING
C895 vdd1.n789 vss 4.48fF $ **FLOATING
C896 vdd1.n790 vss 4.08fF $ **FLOATING
C897 vdd1.n792 vss 33.04fF $ **FLOATING
C898 vdd1.n793 vss 4.27fF $ **FLOATING
C899 vdd1.n794 vss 4.48fF $ **FLOATING
C900 vdd1.n795 vss 4.48fF $ **FLOATING
C901 vdd1.n796 vss 4.48fF $ **FLOATING
C902 vdd1.n797 vss 4.59fF $ **FLOATING
C903 vdd1.n798 vss 4.60fF $ **FLOATING
C904 vdd1.n799 vss 4.48fF $ **FLOATING
C905 vdd1.n800 vss 4.48fF $ **FLOATING
C906 vdd1.n801 vss 4.48fF $ **FLOATING
C907 vdd1.n802 vss 4.08fF $ **FLOATING
C908 vdd1.n806 vss 33.04fF $ **FLOATING
C909 vdd1.n809 vss 4.27fF $ **FLOATING
C910 vdd1.n810 vss 4.48fF $ **FLOATING
C911 vdd1.n811 vss 4.48fF $ **FLOATING
C912 vdd1.n812 vss 4.48fF $ **FLOATING
C913 vdd1.n813 vss 4.59fF $ **FLOATING
C914 vdd1.n814 vss 4.60fF $ **FLOATING
C915 vdd1.n815 vss 4.48fF $ **FLOATING
C916 vdd1.n816 vss 4.48fF $ **FLOATING
C917 vdd1.n817 vss 4.48fF $ **FLOATING
C918 vdd1.n818 vss 4.08fF $ **FLOATING
C919 vdd1.n820 vss 33.04fF $ **FLOATING
C920 vdd1.n821 vss 4.27fF $ **FLOATING
C921 vdd1.n822 vss 4.48fF $ **FLOATING
C922 vdd1.n823 vss 4.48fF $ **FLOATING
C923 vdd1.n824 vss 4.48fF $ **FLOATING
C924 vdd1.n825 vss 4.59fF $ **FLOATING
C925 vdd1.n826 vss 4.60fF $ **FLOATING
C926 vdd1.n827 vss 4.48fF $ **FLOATING
C927 vdd1.n828 vss 4.48fF $ **FLOATING
C928 vdd1.n829 vss 4.48fF $ **FLOATING
C929 vdd1.n830 vss 4.08fF $ **FLOATING
C930 vdd1.n834 vss 33.04fF $ **FLOATING
C931 vdd1.n837 vss 4.27fF $ **FLOATING
C932 vdd1.n838 vss 4.48fF $ **FLOATING
C933 vdd1.n839 vss 4.48fF $ **FLOATING
C934 vdd1.n840 vss 4.48fF $ **FLOATING
C935 vdd1.n841 vss 4.59fF $ **FLOATING
C936 vdd1.n842 vss 4.60fF $ **FLOATING
C937 vdd1.n843 vss 4.48fF $ **FLOATING
C938 vdd1.n844 vss 4.48fF $ **FLOATING
C939 vdd1.n845 vss 4.48fF $ **FLOATING
C940 vdd1.n846 vss 4.08fF $ **FLOATING
C941 vdd1.n848 vss 33.04fF $ **FLOATING
C942 vdd1.n849 vss 4.27fF $ **FLOATING
C943 vdd1.n850 vss 4.48fF $ **FLOATING
C944 vdd1.n851 vss 4.48fF $ **FLOATING
C945 vdd1.n852 vss 4.48fF $ **FLOATING
C946 vdd1.n853 vss 4.59fF $ **FLOATING
C947 vdd1.n854 vss 4.60fF $ **FLOATING
C948 vdd1.n855 vss 4.48fF $ **FLOATING
C949 vdd1.n856 vss 4.48fF $ **FLOATING
C950 vdd1.n857 vss 4.48fF $ **FLOATING
C951 vdd1.n858 vss 4.08fF $ **FLOATING
C952 vdd1.n862 vss 33.04fF $ **FLOATING
C953 vdd1.n865 vss 4.27fF $ **FLOATING
C954 vdd1.n866 vss 4.48fF $ **FLOATING
C955 vdd1.n867 vss 4.48fF $ **FLOATING
C956 vdd1.n868 vss 4.48fF $ **FLOATING
C957 vdd1.n869 vss 4.59fF $ **FLOATING
C958 vdd1.n870 vss 4.60fF $ **FLOATING
C959 vdd1.n871 vss 4.48fF $ **FLOATING
C960 vdd1.n872 vss 4.48fF $ **FLOATING
C961 vdd1.n873 vss 4.48fF $ **FLOATING
C962 vdd1.n874 vss 4.08fF $ **FLOATING
C963 vdd1.n876 vss 33.04fF $ **FLOATING
C964 vdd1.n877 vss 4.27fF $ **FLOATING
C965 vdd1.n878 vss 4.48fF $ **FLOATING
C966 vdd1.n879 vss 4.48fF $ **FLOATING
C967 vdd1.n880 vss 4.48fF $ **FLOATING
C968 vdd1.n881 vss 4.59fF $ **FLOATING
C969 vdd1.n882 vss 4.60fF $ **FLOATING
C970 vdd1.n883 vss 4.48fF $ **FLOATING
C971 vdd1.n884 vss 4.48fF $ **FLOATING
C972 vdd1.n885 vss 4.48fF $ **FLOATING
C973 vdd1.n886 vss 4.08fF $ **FLOATING
C974 vdd1.n890 vss 33.04fF $ **FLOATING
C975 vdd1.n893 vss 4.27fF $ **FLOATING
C976 vdd1.n894 vss 4.48fF $ **FLOATING
C977 vdd1.n895 vss 4.48fF $ **FLOATING
C978 vdd1.n896 vss 4.48fF $ **FLOATING
C979 vdd1.n897 vss 4.59fF $ **FLOATING
C980 vdd1.n898 vss 4.60fF $ **FLOATING
C981 vdd1.n899 vss 4.48fF $ **FLOATING
C982 vdd1.n900 vss 4.48fF $ **FLOATING
C983 vdd1.n901 vss 4.48fF $ **FLOATING
C984 vdd1.n902 vss 4.08fF $ **FLOATING
C985 vdd1.n904 vss 33.04fF $ **FLOATING
C986 vdd1.n905 vss 4.27fF $ **FLOATING
C987 vdd1.n906 vss 4.48fF $ **FLOATING
C988 vdd1.n907 vss 4.48fF $ **FLOATING
C989 vdd1.n908 vss 4.48fF $ **FLOATING
C990 vdd1.n909 vss 4.59fF $ **FLOATING
C991 vdd1.n910 vss 4.60fF $ **FLOATING
C992 vdd1.n911 vss 4.48fF $ **FLOATING
C993 vdd1.n912 vss 4.48fF $ **FLOATING
C994 vdd1.n913 vss 4.48fF $ **FLOATING
C995 vdd1.n914 vss 4.08fF $ **FLOATING
C996 vdd1.n918 vss 33.04fF $ **FLOATING
C997 vdd1.n921 vss 4.27fF $ **FLOATING
C998 vdd1.n922 vss 4.48fF $ **FLOATING
C999 vdd1.n923 vss 4.48fF $ **FLOATING
C1000 vdd1.n924 vss 4.48fF $ **FLOATING
C1001 vdd1.n925 vss 4.59fF $ **FLOATING
C1002 vdd1.n926 vss 4.60fF $ **FLOATING
C1003 vdd1.n927 vss 4.48fF $ **FLOATING
C1004 vdd1.n928 vss 4.48fF $ **FLOATING
C1005 vdd1.n929 vss 4.48fF $ **FLOATING
C1006 vdd1.n930 vss 4.08fF $ **FLOATING
C1007 vdd1.n932 vss 33.04fF $ **FLOATING
C1008 vdd1.n933 vss 4.27fF $ **FLOATING
C1009 vdd1.n934 vss 4.48fF $ **FLOATING
C1010 vdd1.n935 vss 4.48fF $ **FLOATING
C1011 vdd1.n936 vss 4.48fF $ **FLOATING
C1012 vdd1.n937 vss 4.59fF $ **FLOATING
C1013 vdd1.n938 vss 4.60fF $ **FLOATING
C1014 vdd1.n939 vss 4.48fF $ **FLOATING
C1015 vdd1.n940 vss 4.48fF $ **FLOATING
C1016 vdd1.n941 vss 4.48fF $ **FLOATING
C1017 vdd1.n942 vss 4.08fF $ **FLOATING
C1018 vdd1.n946 vss 30.38fF $ **FLOATING
C1019 vdd1.n947 vss 35.69fF $ **FLOATING
C1020 out_p.n0 vss 3.87fF $ **FLOATING
C1021 out_p.n1 vss 4.05fF $ **FLOATING
C1022 out_p.n2 vss 4.05fF $ **FLOATING
C1023 out_p.n3 vss 4.05fF $ **FLOATING
C1024 out_p.n4 vss 4.15fF $ **FLOATING
C1025 out_p.n5 vss 4.15fF $ **FLOATING
C1026 out_p.n6 vss 4.05fF $ **FLOATING
C1027 out_p.n7 vss 4.05fF $ **FLOATING
C1028 out_p.n8 vss 4.05fF $ **FLOATING
C1029 out_p.n9 vss 3.80fF $ **FLOATING
C1030 out_p.n10 vss 3.87fF $ **FLOATING
C1031 out_p.n11 vss 4.05fF $ **FLOATING
C1032 out_p.n12 vss 4.05fF $ **FLOATING
C1033 out_p.n13 vss 4.05fF $ **FLOATING
C1034 out_p.n14 vss 4.15fF $ **FLOATING
C1035 out_p.n15 vss 4.15fF $ **FLOATING
C1036 out_p.n16 vss 4.05fF $ **FLOATING
C1037 out_p.n17 vss 4.05fF $ **FLOATING
C1038 out_p.n18 vss 4.05fF $ **FLOATING
C1039 out_p.n19 vss 3.80fF $ **FLOATING
C1040 out_p.n20 vss 3.85fF $ **FLOATING
C1041 out_p.n21 vss 3.81fF $ **FLOATING
C1042 out_p.n22 vss 3.85fF $ **FLOATING
C1043 out_p.n23 vss 3.81fF $ **FLOATING
C1044 out_p.n24 vss 3.87fF $ **FLOATING
C1045 out_p.n25 vss 4.05fF $ **FLOATING
C1046 out_p.n26 vss 4.05fF $ **FLOATING
C1047 out_p.n27 vss 4.05fF $ **FLOATING
C1048 out_p.n28 vss 4.15fF $ **FLOATING
C1049 out_p.n29 vss 4.15fF $ **FLOATING
C1050 out_p.n30 vss 4.05fF $ **FLOATING
C1051 out_p.n31 vss 4.05fF $ **FLOATING
C1052 out_p.n32 vss 4.05fF $ **FLOATING
C1053 out_p.n33 vss 3.80fF $ **FLOATING
C1054 out_p.n34 vss 3.85fF $ **FLOATING
C1055 out_p.n35 vss 3.81fF $ **FLOATING
C1056 out_p.n36 vss 3.87fF $ **FLOATING
C1057 out_p.n37 vss 4.05fF $ **FLOATING
C1058 out_p.n38 vss 4.05fF $ **FLOATING
C1059 out_p.n39 vss 4.05fF $ **FLOATING
C1060 out_p.n40 vss 4.15fF $ **FLOATING
C1061 out_p.n41 vss 4.15fF $ **FLOATING
C1062 out_p.n42 vss 4.05fF $ **FLOATING
C1063 out_p.n43 vss 4.05fF $ **FLOATING
C1064 out_p.n44 vss 4.05fF $ **FLOATING
C1065 out_p.n45 vss 3.80fF $ **FLOATING
C1066 out_p.n46 vss 3.85fF $ **FLOATING
C1067 out_p.n47 vss 3.81fF $ **FLOATING
C1068 out_p.n48 vss 3.87fF $ **FLOATING
C1069 out_p.n49 vss 4.05fF $ **FLOATING
C1070 out_p.n50 vss 4.05fF $ **FLOATING
C1071 out_p.n51 vss 4.05fF $ **FLOATING
C1072 out_p.n52 vss 4.15fF $ **FLOATING
C1073 out_p.n53 vss 4.15fF $ **FLOATING
C1074 out_p.n54 vss 4.05fF $ **FLOATING
C1075 out_p.n55 vss 4.05fF $ **FLOATING
C1076 out_p.n56 vss 4.05fF $ **FLOATING
C1077 out_p.n57 vss 3.80fF $ **FLOATING
C1078 out_p.n58 vss 3.85fF $ **FLOATING
C1079 out_p.n59 vss 3.81fF $ **FLOATING
C1080 out_p.n60 vss 3.87fF $ **FLOATING
C1081 out_p.n61 vss 4.05fF $ **FLOATING
C1082 out_p.n62 vss 4.05fF $ **FLOATING
C1083 out_p.n63 vss 4.05fF $ **FLOATING
C1084 out_p.n64 vss 4.15fF $ **FLOATING
C1085 out_p.n65 vss 4.15fF $ **FLOATING
C1086 out_p.n66 vss 4.05fF $ **FLOATING
C1087 out_p.n67 vss 4.05fF $ **FLOATING
C1088 out_p.n68 vss 4.05fF $ **FLOATING
C1089 out_p.n69 vss 3.80fF $ **FLOATING
C1090 out_p.n70 vss 3.85fF $ **FLOATING
C1091 out_p.n71 vss 3.81fF $ **FLOATING
C1092 out_p.n72 vss 3.87fF $ **FLOATING
C1093 out_p.n73 vss 4.05fF $ **FLOATING
C1094 out_p.n74 vss 4.05fF $ **FLOATING
C1095 out_p.n75 vss 4.05fF $ **FLOATING
C1096 out_p.n76 vss 4.15fF $ **FLOATING
C1097 out_p.n77 vss 4.15fF $ **FLOATING
C1098 out_p.n78 vss 4.05fF $ **FLOATING
C1099 out_p.n79 vss 4.05fF $ **FLOATING
C1100 out_p.n80 vss 4.05fF $ **FLOATING
C1101 out_p.n81 vss 3.80fF $ **FLOATING
C1102 out_p.n82 vss 3.85fF $ **FLOATING
C1103 out_p.n83 vss 3.81fF $ **FLOATING
C1104 out_p.n84 vss 3.87fF $ **FLOATING
C1105 out_p.n85 vss 4.05fF $ **FLOATING
C1106 out_p.n86 vss 4.05fF $ **FLOATING
C1107 out_p.n87 vss 4.05fF $ **FLOATING
C1108 out_p.n88 vss 4.15fF $ **FLOATING
C1109 out_p.n89 vss 4.15fF $ **FLOATING
C1110 out_p.n90 vss 4.05fF $ **FLOATING
C1111 out_p.n91 vss 4.05fF $ **FLOATING
C1112 out_p.n92 vss 4.05fF $ **FLOATING
C1113 out_p.n93 vss 3.80fF $ **FLOATING
C1114 out_p.n94 vss 3.85fF $ **FLOATING
C1115 out_p.n95 vss 3.81fF $ **FLOATING
C1116 out_p.n96 vss 3.87fF $ **FLOATING
C1117 out_p.n97 vss 4.05fF $ **FLOATING
C1118 out_p.n98 vss 4.05fF $ **FLOATING
C1119 out_p.n99 vss 4.05fF $ **FLOATING
C1120 out_p.n100 vss 4.15fF $ **FLOATING
C1121 out_p.n101 vss 4.15fF $ **FLOATING
C1122 out_p.n102 vss 4.05fF $ **FLOATING
C1123 out_p.n103 vss 4.05fF $ **FLOATING
C1124 out_p.n104 vss 4.05fF $ **FLOATING
C1125 out_p.n105 vss 3.80fF $ **FLOATING
C1126 out_p.n106 vss 3.85fF $ **FLOATING
C1127 out_p.n107 vss 3.81fF $ **FLOATING
C1128 out_p.n108 vss 3.87fF $ **FLOATING
C1129 out_p.n109 vss 4.05fF $ **FLOATING
C1130 out_p.n110 vss 4.05fF $ **FLOATING
C1131 out_p.n111 vss 4.05fF $ **FLOATING
C1132 out_p.n112 vss 4.15fF $ **FLOATING
C1133 out_p.n113 vss 4.15fF $ **FLOATING
C1134 out_p.n114 vss 4.05fF $ **FLOATING
C1135 out_p.n115 vss 4.05fF $ **FLOATING
C1136 out_p.n116 vss 4.05fF $ **FLOATING
C1137 out_p.n117 vss 3.80fF $ **FLOATING
C1138 out_p.n118 vss 3.85fF $ **FLOATING
C1139 out_p.n119 vss 3.81fF $ **FLOATING
C1140 out_p.n120 vss 3.87fF $ **FLOATING
C1141 out_p.n121 vss 4.05fF $ **FLOATING
C1142 out_p.n122 vss 4.05fF $ **FLOATING
C1143 out_p.n123 vss 4.05fF $ **FLOATING
C1144 out_p.n124 vss 4.15fF $ **FLOATING
C1145 out_p.n125 vss 4.15fF $ **FLOATING
C1146 out_p.n126 vss 4.05fF $ **FLOATING
C1147 out_p.n127 vss 4.05fF $ **FLOATING
C1148 out_p.n128 vss 4.05fF $ **FLOATING
C1149 out_p.n129 vss 3.80fF $ **FLOATING
C1150 out_p.n130 vss 3.85fF $ **FLOATING
C1151 out_p.n131 vss 3.81fF $ **FLOATING
C1152 out_p.n132 vss 3.87fF $ **FLOATING
C1153 out_p.n133 vss 4.05fF $ **FLOATING
C1154 out_p.n134 vss 4.05fF $ **FLOATING
C1155 out_p.n135 vss 4.05fF $ **FLOATING
C1156 out_p.n136 vss 4.15fF $ **FLOATING
C1157 out_p.n137 vss 4.15fF $ **FLOATING
C1158 out_p.n138 vss 4.05fF $ **FLOATING
C1159 out_p.n139 vss 4.05fF $ **FLOATING
C1160 out_p.n140 vss 4.05fF $ **FLOATING
C1161 out_p.n141 vss 3.80fF $ **FLOATING
C1162 out_p.n142 vss 3.85fF $ **FLOATING
C1163 out_p.n143 vss 3.81fF $ **FLOATING
C1164 out_p.n144 vss 3.87fF $ **FLOATING
C1165 out_p.n145 vss 4.05fF $ **FLOATING
C1166 out_p.n146 vss 4.05fF $ **FLOATING
C1167 out_p.n147 vss 4.05fF $ **FLOATING
C1168 out_p.n148 vss 4.15fF $ **FLOATING
C1169 out_p.n149 vss 4.15fF $ **FLOATING
C1170 out_p.n150 vss 4.05fF $ **FLOATING
C1171 out_p.n151 vss 4.05fF $ **FLOATING
C1172 out_p.n152 vss 4.05fF $ **FLOATING
C1173 out_p.n153 vss 3.80fF $ **FLOATING
C1174 out_p.n154 vss 3.85fF $ **FLOATING
C1175 out_p.n155 vss 3.81fF $ **FLOATING
C1176 out_p.n156 vss 3.87fF $ **FLOATING
C1177 out_p.n157 vss 4.05fF $ **FLOATING
C1178 out_p.n158 vss 4.05fF $ **FLOATING
C1179 out_p.n159 vss 4.05fF $ **FLOATING
C1180 out_p.n160 vss 4.15fF $ **FLOATING
C1181 out_p.n161 vss 4.15fF $ **FLOATING
C1182 out_p.n162 vss 4.05fF $ **FLOATING
C1183 out_p.n163 vss 4.05fF $ **FLOATING
C1184 out_p.n164 vss 4.05fF $ **FLOATING
C1185 out_p.n165 vss 3.80fF $ **FLOATING
C1186 out_p.n166 vss 3.85fF $ **FLOATING
C1187 out_p.n167 vss 3.81fF $ **FLOATING
C1188 out_p.n168 vss 3.87fF $ **FLOATING
C1189 out_p.n169 vss 4.05fF $ **FLOATING
C1190 out_p.n170 vss 4.05fF $ **FLOATING
C1191 out_p.n171 vss 4.05fF $ **FLOATING
C1192 out_p.n172 vss 4.15fF $ **FLOATING
C1193 out_p.n173 vss 4.15fF $ **FLOATING
C1194 out_p.n174 vss 4.05fF $ **FLOATING
C1195 out_p.n175 vss 4.05fF $ **FLOATING
C1196 out_p.n176 vss 4.05fF $ **FLOATING
C1197 out_p.n177 vss 3.80fF $ **FLOATING
C1198 out_p.n178 vss 3.85fF $ **FLOATING
C1199 out_p.n179 vss 3.81fF $ **FLOATING
C1200 out_p.n180 vss 3.87fF $ **FLOATING
C1201 out_p.n181 vss 4.05fF $ **FLOATING
C1202 out_p.n182 vss 4.05fF $ **FLOATING
C1203 out_p.n183 vss 4.05fF $ **FLOATING
C1204 out_p.n184 vss 4.15fF $ **FLOATING
C1205 out_p.n185 vss 4.15fF $ **FLOATING
C1206 out_p.n186 vss 4.05fF $ **FLOATING
C1207 out_p.n187 vss 4.05fF $ **FLOATING
C1208 out_p.n188 vss 4.05fF $ **FLOATING
C1209 out_p.n189 vss 3.80fF $ **FLOATING
C1210 out_p.n190 vss 3.85fF $ **FLOATING
C1211 out_p.n191 vss 3.81fF $ **FLOATING
C1212 out_p.n192 vss 3.87fF $ **FLOATING
C1213 out_p.n193 vss 4.05fF $ **FLOATING
C1214 out_p.n194 vss 4.05fF $ **FLOATING
C1215 out_p.n195 vss 4.05fF $ **FLOATING
C1216 out_p.n196 vss 4.15fF $ **FLOATING
C1217 out_p.n197 vss 4.15fF $ **FLOATING
C1218 out_p.n198 vss 4.05fF $ **FLOATING
C1219 out_p.n199 vss 4.05fF $ **FLOATING
C1220 out_p.n200 vss 4.05fF $ **FLOATING
C1221 out_p.n201 vss 3.80fF $ **FLOATING
C1222 out_p.n202 vss 3.85fF $ **FLOATING
C1223 out_p.n203 vss 3.81fF $ **FLOATING
C1224 out_p.n204 vss 3.87fF $ **FLOATING
C1225 out_p.n205 vss 4.05fF $ **FLOATING
C1226 out_p.n206 vss 4.05fF $ **FLOATING
C1227 out_p.n207 vss 4.05fF $ **FLOATING
C1228 out_p.n208 vss 4.15fF $ **FLOATING
C1229 out_p.n209 vss 4.15fF $ **FLOATING
C1230 out_p.n210 vss 4.05fF $ **FLOATING
C1231 out_p.n211 vss 4.05fF $ **FLOATING
C1232 out_p.n212 vss 4.05fF $ **FLOATING
C1233 out_p.n213 vss 3.80fF $ **FLOATING
C1234 out_p.n214 vss 3.85fF $ **FLOATING
C1235 out_p.n215 vss 3.81fF $ **FLOATING
C1236 out_p.n216 vss 3.87fF $ **FLOATING
C1237 out_p.n217 vss 4.05fF $ **FLOATING
C1238 out_p.n218 vss 4.05fF $ **FLOATING
C1239 out_p.n219 vss 4.05fF $ **FLOATING
C1240 out_p.n220 vss 4.15fF $ **FLOATING
C1241 out_p.n221 vss 4.15fF $ **FLOATING
C1242 out_p.n222 vss 4.05fF $ **FLOATING
C1243 out_p.n223 vss 4.05fF $ **FLOATING
C1244 out_p.n224 vss 4.05fF $ **FLOATING
C1245 out_p.n225 vss 3.80fF $ **FLOATING
C1246 out_p.n226 vss 3.85fF $ **FLOATING
C1247 out_p.n227 vss 3.81fF $ **FLOATING
C1248 out_p.n228 vss 3.87fF $ **FLOATING
C1249 out_p.n229 vss 4.05fF $ **FLOATING
C1250 out_p.n230 vss 4.05fF $ **FLOATING
C1251 out_p.n231 vss 4.05fF $ **FLOATING
C1252 out_p.n232 vss 4.15fF $ **FLOATING
C1253 out_p.n233 vss 4.15fF $ **FLOATING
C1254 out_p.n234 vss 4.05fF $ **FLOATING
C1255 out_p.n235 vss 4.05fF $ **FLOATING
C1256 out_p.n236 vss 4.05fF $ **FLOATING
C1257 out_p.n237 vss 3.80fF $ **FLOATING
C1258 out_p.n238 vss 3.85fF $ **FLOATING
C1259 out_p.n239 vss 3.81fF $ **FLOATING
C1260 out_p.n240 vss 3.87fF $ **FLOATING
C1261 out_p.n241 vss 4.05fF $ **FLOATING
C1262 out_p.n242 vss 4.05fF $ **FLOATING
C1263 out_p.n243 vss 4.05fF $ **FLOATING
C1264 out_p.n244 vss 4.15fF $ **FLOATING
C1265 out_p.n245 vss 4.15fF $ **FLOATING
C1266 out_p.n246 vss 4.05fF $ **FLOATING
C1267 out_p.n247 vss 4.05fF $ **FLOATING
C1268 out_p.n248 vss 4.05fF $ **FLOATING
C1269 out_p.n249 vss 3.80fF $ **FLOATING
C1270 out_p.n250 vss 3.85fF $ **FLOATING
C1271 out_p.n251 vss 3.81fF $ **FLOATING
C1272 out_p.n252 vss 3.87fF $ **FLOATING
C1273 out_p.n253 vss 4.05fF $ **FLOATING
C1274 out_p.n254 vss 4.05fF $ **FLOATING
C1275 out_p.n255 vss 4.05fF $ **FLOATING
C1276 out_p.n256 vss 4.15fF $ **FLOATING
C1277 out_p.n257 vss 4.15fF $ **FLOATING
C1278 out_p.n258 vss 4.05fF $ **FLOATING
C1279 out_p.n259 vss 4.05fF $ **FLOATING
C1280 out_p.n260 vss 4.05fF $ **FLOATING
C1281 out_p.n261 vss 3.80fF $ **FLOATING
C1282 out_p.n262 vss 3.85fF $ **FLOATING
C1283 out_p.n263 vss 3.81fF $ **FLOATING
C1284 out_p.n264 vss 3.87fF $ **FLOATING
C1285 out_p.n265 vss 4.05fF $ **FLOATING
C1286 out_p.n266 vss 4.05fF $ **FLOATING
C1287 out_p.n267 vss 4.05fF $ **FLOATING
C1288 out_p.n268 vss 4.15fF $ **FLOATING
C1289 out_p.n269 vss 4.15fF $ **FLOATING
C1290 out_p.n270 vss 4.05fF $ **FLOATING
C1291 out_p.n271 vss 4.05fF $ **FLOATING
C1292 out_p.n272 vss 4.05fF $ **FLOATING
C1293 out_p.n273 vss 3.80fF $ **FLOATING
C1294 out_p.n274 vss 3.85fF $ **FLOATING
C1295 out_p.n275 vss 3.81fF $ **FLOATING
C1296 out_p.n276 vss 3.87fF $ **FLOATING
C1297 out_p.n277 vss 4.05fF $ **FLOATING
C1298 out_p.n278 vss 4.05fF $ **FLOATING
C1299 out_p.n279 vss 4.05fF $ **FLOATING
C1300 out_p.n280 vss 4.15fF $ **FLOATING
C1301 out_p.n281 vss 4.15fF $ **FLOATING
C1302 out_p.n282 vss 4.05fF $ **FLOATING
C1303 out_p.n283 vss 4.05fF $ **FLOATING
C1304 out_p.n284 vss 4.05fF $ **FLOATING
C1305 out_p.n285 vss 3.80fF $ **FLOATING
C1306 out_p.n286 vss 3.85fF $ **FLOATING
C1307 out_p.n287 vss 3.81fF $ **FLOATING
C1308 out_p.n288 vss 3.87fF $ **FLOATING
C1309 out_p.n289 vss 4.05fF $ **FLOATING
C1310 out_p.n290 vss 4.05fF $ **FLOATING
C1311 out_p.n291 vss 4.05fF $ **FLOATING
C1312 out_p.n292 vss 4.15fF $ **FLOATING
C1313 out_p.n293 vss 4.15fF $ **FLOATING
C1314 out_p.n294 vss 4.05fF $ **FLOATING
C1315 out_p.n295 vss 4.05fF $ **FLOATING
C1316 out_p.n296 vss 4.05fF $ **FLOATING
C1317 out_p.n297 vss 3.80fF $ **FLOATING
C1318 out_p.n298 vss 3.85fF $ **FLOATING
C1319 out_p.n299 vss 3.81fF $ **FLOATING
C1320 out_p.n300 vss 3.87fF $ **FLOATING
C1321 out_p.n301 vss 4.05fF $ **FLOATING
C1322 out_p.n302 vss 4.05fF $ **FLOATING
C1323 out_p.n303 vss 4.05fF $ **FLOATING
C1324 out_p.n304 vss 4.15fF $ **FLOATING
C1325 out_p.n305 vss 4.15fF $ **FLOATING
C1326 out_p.n306 vss 4.05fF $ **FLOATING
C1327 out_p.n307 vss 4.05fF $ **FLOATING
C1328 out_p.n308 vss 4.05fF $ **FLOATING
C1329 out_p.n309 vss 3.80fF $ **FLOATING
C1330 out_p.n310 vss 3.85fF $ **FLOATING
C1331 out_p.n311 vss 3.81fF $ **FLOATING
C1332 out_p.n312 vss 3.87fF $ **FLOATING
C1333 out_p.n313 vss 4.05fF $ **FLOATING
C1334 out_p.n314 vss 4.05fF $ **FLOATING
C1335 out_p.n315 vss 4.05fF $ **FLOATING
C1336 out_p.n316 vss 4.15fF $ **FLOATING
C1337 out_p.n317 vss 4.15fF $ **FLOATING
C1338 out_p.n318 vss 4.05fF $ **FLOATING
C1339 out_p.n319 vss 4.05fF $ **FLOATING
C1340 out_p.n320 vss 4.05fF $ **FLOATING
C1341 out_p.n321 vss 3.80fF $ **FLOATING
C1342 out_p.n322 vss 3.85fF $ **FLOATING
C1343 out_p.n323 vss 3.81fF $ **FLOATING
C1344 out_p.n324 vss 3.87fF $ **FLOATING
C1345 out_p.n325 vss 4.05fF $ **FLOATING
C1346 out_p.n326 vss 4.05fF $ **FLOATING
C1347 out_p.n327 vss 4.05fF $ **FLOATING
C1348 out_p.n328 vss 4.15fF $ **FLOATING
C1349 out_p.n329 vss 4.15fF $ **FLOATING
C1350 out_p.n330 vss 4.05fF $ **FLOATING
C1351 out_p.n331 vss 4.05fF $ **FLOATING
C1352 out_p.n332 vss 4.05fF $ **FLOATING
C1353 out_p.n333 vss 3.80fF $ **FLOATING
C1354 out_p.n334 vss 3.85fF $ **FLOATING
C1355 out_p.n335 vss 3.81fF $ **FLOATING
C1356 out_p.n336 vss 3.87fF $ **FLOATING
C1357 out_p.n337 vss 4.05fF $ **FLOATING
C1358 out_p.n338 vss 4.05fF $ **FLOATING
C1359 out_p.n339 vss 4.05fF $ **FLOATING
C1360 out_p.n340 vss 4.15fF $ **FLOATING
C1361 out_p.n341 vss 4.15fF $ **FLOATING
C1362 out_p.n342 vss 4.05fF $ **FLOATING
C1363 out_p.n343 vss 4.05fF $ **FLOATING
C1364 out_p.n344 vss 4.05fF $ **FLOATING
C1365 out_p.n345 vss 3.80fF $ **FLOATING
C1366 out_p.n346 vss 3.85fF $ **FLOATING
C1367 out_p.n347 vss 3.81fF $ **FLOATING
C1368 out_p.n348 vss 3.87fF $ **FLOATING
C1369 out_p.n349 vss 4.05fF $ **FLOATING
C1370 out_p.n350 vss 4.05fF $ **FLOATING
C1371 out_p.n351 vss 4.05fF $ **FLOATING
C1372 out_p.n352 vss 4.15fF $ **FLOATING
C1373 out_p.n353 vss 4.15fF $ **FLOATING
C1374 out_p.n354 vss 4.05fF $ **FLOATING
C1375 out_p.n355 vss 4.05fF $ **FLOATING
C1376 out_p.n356 vss 4.05fF $ **FLOATING
C1377 out_p.n357 vss 3.80fF $ **FLOATING
C1378 out_p.n358 vss 3.85fF $ **FLOATING
C1379 out_p.n359 vss 3.81fF $ **FLOATING
C1380 out_p.n360 vss 3.87fF $ **FLOATING
C1381 out_p.n361 vss 4.05fF $ **FLOATING
C1382 out_p.n362 vss 4.05fF $ **FLOATING
C1383 out_p.n363 vss 4.05fF $ **FLOATING
C1384 out_p.n364 vss 4.15fF $ **FLOATING
C1385 out_p.n365 vss 4.15fF $ **FLOATING
C1386 out_p.n366 vss 4.05fF $ **FLOATING
C1387 out_p.n367 vss 4.05fF $ **FLOATING
C1388 out_p.n368 vss 4.05fF $ **FLOATING
C1389 out_p.n369 vss 3.80fF $ **FLOATING
C1390 out_p.n370 vss 3.85fF $ **FLOATING
C1391 out_p.n371 vss 3.81fF $ **FLOATING
C1392 out_p.n372 vss 3.87fF $ **FLOATING
C1393 out_p.n373 vss 4.05fF $ **FLOATING
C1394 out_p.n374 vss 4.05fF $ **FLOATING
C1395 out_p.n375 vss 4.05fF $ **FLOATING
C1396 out_p.n376 vss 4.15fF $ **FLOATING
C1397 out_p.n377 vss 4.15fF $ **FLOATING
C1398 out_p.n378 vss 4.05fF $ **FLOATING
C1399 out_p.n379 vss 4.05fF $ **FLOATING
C1400 out_p.n380 vss 4.05fF $ **FLOATING
C1401 out_p.n381 vss 3.80fF $ **FLOATING
C1402 out_p.n382 vss 3.85fF $ **FLOATING
C1403 out_p.n383 vss 3.81fF $ **FLOATING
C1404 out_p.n384 vss 3.87fF $ **FLOATING
C1405 out_p.n385 vss 4.05fF $ **FLOATING
C1406 out_p.n386 vss 4.05fF $ **FLOATING
C1407 out_p.n387 vss 4.05fF $ **FLOATING
C1408 out_p.n388 vss 4.15fF $ **FLOATING
C1409 out_p.n389 vss 4.15fF $ **FLOATING
C1410 out_p.n390 vss 4.05fF $ **FLOATING
C1411 out_p.n391 vss 4.05fF $ **FLOATING
C1412 out_p.n392 vss 4.05fF $ **FLOATING
C1413 out_p.n393 vss 3.80fF $ **FLOATING
C1414 out_p.n394 vss 3.85fF $ **FLOATING
C1415 out_p.n395 vss 3.81fF $ **FLOATING
C1416 out_p.n396 vss 3.87fF $ **FLOATING
C1417 out_p.n397 vss 4.05fF $ **FLOATING
C1418 out_p.n398 vss 4.05fF $ **FLOATING
C1419 out_p.n399 vss 4.05fF $ **FLOATING
C1420 out_p.n400 vss 4.15fF $ **FLOATING
C1421 out_p.n401 vss 4.15fF $ **FLOATING
C1422 out_p.n402 vss 4.05fF $ **FLOATING
C1423 out_p.n403 vss 4.05fF $ **FLOATING
C1424 out_p.n404 vss 4.05fF $ **FLOATING
C1425 out_p.n405 vss 3.80fF $ **FLOATING
C1426 out_p.n406 vss 3.85fF $ **FLOATING
C1427 out_p.n407 vss 3.81fF $ **FLOATING
C1428 out_p.n408 vss 3.87fF $ **FLOATING
C1429 out_p.n409 vss 4.05fF $ **FLOATING
C1430 out_p.n410 vss 4.05fF $ **FLOATING
C1431 out_p.n411 vss 4.05fF $ **FLOATING
C1432 out_p.n412 vss 4.15fF $ **FLOATING
C1433 out_p.n413 vss 4.15fF $ **FLOATING
C1434 out_p.n414 vss 4.05fF $ **FLOATING
C1435 out_p.n415 vss 4.05fF $ **FLOATING
C1436 out_p.n416 vss 4.05fF $ **FLOATING
C1437 out_p.n417 vss 3.80fF $ **FLOATING
C1438 out_p.n418 vss 3.85fF $ **FLOATING
C1439 out_p.n419 vss 3.81fF $ **FLOATING
C1440 out_p.n420 vss 3.87fF $ **FLOATING
C1441 out_p.n421 vss 4.05fF $ **FLOATING
C1442 out_p.n422 vss 4.05fF $ **FLOATING
C1443 out_p.n423 vss 4.05fF $ **FLOATING
C1444 out_p.n424 vss 4.15fF $ **FLOATING
C1445 out_p.n425 vss 4.15fF $ **FLOATING
C1446 out_p.n426 vss 4.05fF $ **FLOATING
C1447 out_p.n427 vss 4.05fF $ **FLOATING
C1448 out_p.n428 vss 4.05fF $ **FLOATING
C1449 out_p.n429 vss 3.80fF $ **FLOATING
C1450 out_p.n430 vss 3.85fF $ **FLOATING
C1451 out_p.n431 vss 3.81fF $ **FLOATING
C1452 out_p.n432 vss 3.87fF $ **FLOATING
C1453 out_p.n433 vss 4.05fF $ **FLOATING
C1454 out_p.n434 vss 4.05fF $ **FLOATING
C1455 out_p.n435 vss 4.05fF $ **FLOATING
C1456 out_p.n436 vss 4.15fF $ **FLOATING
C1457 out_p.n437 vss 4.15fF $ **FLOATING
C1458 out_p.n438 vss 4.05fF $ **FLOATING
C1459 out_p.n439 vss 4.05fF $ **FLOATING
C1460 out_p.n440 vss 4.05fF $ **FLOATING
C1461 out_p.n441 vss 3.80fF $ **FLOATING
C1462 out_p.n442 vss 3.85fF $ **FLOATING
C1463 out_p.n443 vss 3.81fF $ **FLOATING
C1464 out_p.n444 vss 3.87fF $ **FLOATING
C1465 out_p.n445 vss 4.05fF $ **FLOATING
C1466 out_p.n446 vss 4.05fF $ **FLOATING
C1467 out_p.n447 vss 4.05fF $ **FLOATING
C1468 out_p.n448 vss 4.15fF $ **FLOATING
C1469 out_p.n449 vss 4.15fF $ **FLOATING
C1470 out_p.n450 vss 4.05fF $ **FLOATING
C1471 out_p.n451 vss 4.05fF $ **FLOATING
C1472 out_p.n452 vss 4.05fF $ **FLOATING
C1473 out_p.n453 vss 3.80fF $ **FLOATING
C1474 out_p.n454 vss 3.85fF $ **FLOATING
C1475 out_p.n455 vss 3.81fF $ **FLOATING
C1476 out_p.n456 vss 3.87fF $ **FLOATING
C1477 out_p.n457 vss 4.05fF $ **FLOATING
C1478 out_p.n458 vss 4.05fF $ **FLOATING
C1479 out_p.n459 vss 4.05fF $ **FLOATING
C1480 out_p.n460 vss 4.15fF $ **FLOATING
C1481 out_p.n461 vss 4.15fF $ **FLOATING
C1482 out_p.n462 vss 4.05fF $ **FLOATING
C1483 out_p.n463 vss 4.05fF $ **FLOATING
C1484 out_p.n464 vss 4.05fF $ **FLOATING
C1485 out_p.n465 vss 3.80fF $ **FLOATING
C1486 out_p.n466 vss 3.85fF $ **FLOATING
C1487 out_p.n467 vss 3.81fF $ **FLOATING
C1488 out_p.n468 vss 3.87fF $ **FLOATING
C1489 out_p.n469 vss 4.05fF $ **FLOATING
C1490 out_p.n470 vss 4.05fF $ **FLOATING
C1491 out_p.n471 vss 4.05fF $ **FLOATING
C1492 out_p.n472 vss 4.15fF $ **FLOATING
C1493 out_p.n473 vss 4.15fF $ **FLOATING
C1494 out_p.n474 vss 4.05fF $ **FLOATING
C1495 out_p.n475 vss 4.05fF $ **FLOATING
C1496 out_p.n476 vss 4.05fF $ **FLOATING
C1497 out_p.n477 vss 3.80fF $ **FLOATING
C1498 out_p.n478 vss 3.85fF $ **FLOATING
C1499 out_p.n479 vss 3.81fF $ **FLOATING
C1500 out_p.n480 vss 3.87fF $ **FLOATING
C1501 out_p.n481 vss 4.05fF $ **FLOATING
C1502 out_p.n482 vss 4.05fF $ **FLOATING
C1503 out_p.n483 vss 4.05fF $ **FLOATING
C1504 out_p.n484 vss 4.15fF $ **FLOATING
C1505 out_p.n485 vss 4.15fF $ **FLOATING
C1506 out_p.n486 vss 4.05fF $ **FLOATING
C1507 out_p.n487 vss 4.05fF $ **FLOATING
C1508 out_p.n488 vss 4.05fF $ **FLOATING
C1509 out_p.n489 vss 3.80fF $ **FLOATING
C1510 out_p.n490 vss 3.85fF $ **FLOATING
C1511 out_p.n491 vss 3.81fF $ **FLOATING
C1512 out_p.n492 vss 3.87fF $ **FLOATING
C1513 out_p.n493 vss 4.05fF $ **FLOATING
C1514 out_p.n494 vss 4.05fF $ **FLOATING
C1515 out_p.n495 vss 4.05fF $ **FLOATING
C1516 out_p.n496 vss 4.15fF $ **FLOATING
C1517 out_p.n497 vss 4.15fF $ **FLOATING
C1518 out_p.n498 vss 4.05fF $ **FLOATING
C1519 out_p.n499 vss 4.05fF $ **FLOATING
C1520 out_p.n500 vss 4.05fF $ **FLOATING
C1521 out_p.n501 vss 3.80fF $ **FLOATING
C1522 out_p.n502 vss 3.85fF $ **FLOATING
C1523 out_p.n503 vss 3.81fF $ **FLOATING
C1524 out_p.n504 vss 3.87fF $ **FLOATING
C1525 out_p.n505 vss 4.05fF $ **FLOATING
C1526 out_p.n506 vss 4.05fF $ **FLOATING
C1527 out_p.n507 vss 4.05fF $ **FLOATING
C1528 out_p.n508 vss 4.15fF $ **FLOATING
C1529 out_p.n509 vss 4.15fF $ **FLOATING
C1530 out_p.n510 vss 4.05fF $ **FLOATING
C1531 out_p.n511 vss 4.05fF $ **FLOATING
C1532 out_p.n512 vss 4.05fF $ **FLOATING
C1533 out_p.n513 vss 3.80fF $ **FLOATING
C1534 out_p.n514 vss 3.85fF $ **FLOATING
C1535 out_p.n515 vss 3.81fF $ **FLOATING
C1536 out_p.n516 vss 3.87fF $ **FLOATING
C1537 out_p.n517 vss 4.05fF $ **FLOATING
C1538 out_p.n518 vss 4.05fF $ **FLOATING
C1539 out_p.n519 vss 4.05fF $ **FLOATING
C1540 out_p.n520 vss 4.15fF $ **FLOATING
C1541 out_p.n521 vss 4.15fF $ **FLOATING
C1542 out_p.n522 vss 4.05fF $ **FLOATING
C1543 out_p.n523 vss 4.05fF $ **FLOATING
C1544 out_p.n524 vss 4.05fF $ **FLOATING
C1545 out_p.n525 vss 3.80fF $ **FLOATING
C1546 out_p.n526 vss 3.85fF $ **FLOATING
C1547 out_p.n527 vss 3.81fF $ **FLOATING
C1548 out_p.n528 vss 3.87fF $ **FLOATING
C1549 out_p.n529 vss 4.05fF $ **FLOATING
C1550 out_p.n530 vss 4.05fF $ **FLOATING
C1551 out_p.n531 vss 4.05fF $ **FLOATING
C1552 out_p.n532 vss 4.15fF $ **FLOATING
C1553 out_p.n533 vss 4.15fF $ **FLOATING
C1554 out_p.n534 vss 4.05fF $ **FLOATING
C1555 out_p.n535 vss 4.05fF $ **FLOATING
C1556 out_p.n536 vss 4.05fF $ **FLOATING
C1557 out_p.n537 vss 3.80fF $ **FLOATING
C1558 out_p.n538 vss 3.85fF $ **FLOATING
C1559 out_p.n539 vss 3.81fF $ **FLOATING
C1560 out_p.n540 vss 3.87fF $ **FLOATING
C1561 out_p.n541 vss 4.05fF $ **FLOATING
C1562 out_p.n542 vss 4.05fF $ **FLOATING
C1563 out_p.n543 vss 4.05fF $ **FLOATING
C1564 out_p.n544 vss 4.15fF $ **FLOATING
C1565 out_p.n545 vss 4.15fF $ **FLOATING
C1566 out_p.n546 vss 4.05fF $ **FLOATING
C1567 out_p.n547 vss 4.05fF $ **FLOATING
C1568 out_p.n548 vss 4.05fF $ **FLOATING
C1569 out_p.n549 vss 3.80fF $ **FLOATING
C1570 out_p.n550 vss 3.85fF $ **FLOATING
C1571 out_p.n551 vss 3.81fF $ **FLOATING
C1572 out_p.n552 vss 3.87fF $ **FLOATING
C1573 out_p.n553 vss 4.05fF $ **FLOATING
C1574 out_p.n554 vss 4.05fF $ **FLOATING
C1575 out_p.n555 vss 4.05fF $ **FLOATING
C1576 out_p.n556 vss 4.15fF $ **FLOATING
C1577 out_p.n557 vss 4.15fF $ **FLOATING
C1578 out_p.n558 vss 4.05fF $ **FLOATING
C1579 out_p.n559 vss 4.05fF $ **FLOATING
C1580 out_p.n560 vss 4.05fF $ **FLOATING
C1581 out_p.n561 vss 3.80fF $ **FLOATING
C1582 out_p.n562 vss 3.85fF $ **FLOATING
C1583 out_p.n563 vss 3.81fF $ **FLOATING
C1584 out_p.n564 vss 3.87fF $ **FLOATING
C1585 out_p.n565 vss 4.05fF $ **FLOATING
C1586 out_p.n566 vss 4.05fF $ **FLOATING
C1587 out_p.n567 vss 4.05fF $ **FLOATING
C1588 out_p.n568 vss 4.15fF $ **FLOATING
C1589 out_p.n569 vss 4.15fF $ **FLOATING
C1590 out_p.n570 vss 4.05fF $ **FLOATING
C1591 out_p.n571 vss 4.05fF $ **FLOATING
C1592 out_p.n572 vss 4.05fF $ **FLOATING
C1593 out_p.n573 vss 3.80fF $ **FLOATING
C1594 out_p.n574 vss 3.85fF $ **FLOATING
C1595 out_p.n575 vss 3.81fF $ **FLOATING
C1596 out_p.n576 vss 3.87fF $ **FLOATING
C1597 out_p.n577 vss 4.05fF $ **FLOATING
C1598 out_p.n578 vss 4.05fF $ **FLOATING
C1599 out_p.n579 vss 4.05fF $ **FLOATING
C1600 out_p.n580 vss 4.15fF $ **FLOATING
C1601 out_p.n581 vss 4.15fF $ **FLOATING
C1602 out_p.n582 vss 4.05fF $ **FLOATING
C1603 out_p.n583 vss 4.05fF $ **FLOATING
C1604 out_p.n584 vss 4.05fF $ **FLOATING
C1605 out_p.n585 vss 3.80fF $ **FLOATING
C1606 out_p.n586 vss 3.85fF $ **FLOATING
C1607 out_p.n587 vss 3.81fF $ **FLOATING
C1608 out_p.n588 vss 3.87fF $ **FLOATING
C1609 out_p.n589 vss 4.05fF $ **FLOATING
C1610 out_p.n590 vss 4.05fF $ **FLOATING
C1611 out_p.n591 vss 4.05fF $ **FLOATING
C1612 out_p.n592 vss 4.15fF $ **FLOATING
C1613 out_p.n593 vss 4.15fF $ **FLOATING
C1614 out_p.n594 vss 4.05fF $ **FLOATING
C1615 out_p.n595 vss 4.05fF $ **FLOATING
C1616 out_p.n596 vss 4.05fF $ **FLOATING
C1617 out_p.n597 vss 3.80fF $ **FLOATING
C1618 out_p.n598 vss 3.85fF $ **FLOATING
C1619 out_p.n599 vss 3.81fF $ **FLOATING
C1620 out_p.n600 vss 3.87fF $ **FLOATING
C1621 out_p.n601 vss 4.05fF $ **FLOATING
C1622 out_p.n602 vss 4.05fF $ **FLOATING
C1623 out_p.n603 vss 4.05fF $ **FLOATING
C1624 out_p.n604 vss 4.15fF $ **FLOATING
C1625 out_p.n605 vss 4.15fF $ **FLOATING
C1626 out_p.n606 vss 4.05fF $ **FLOATING
C1627 out_p.n607 vss 4.05fF $ **FLOATING
C1628 out_p.n608 vss 4.05fF $ **FLOATING
C1629 out_p.n609 vss 3.80fF $ **FLOATING
C1630 out_p.n610 vss 3.85fF $ **FLOATING
C1631 out_p.n611 vss 3.81fF $ **FLOATING
C1632 out_p.n612 vss 3.87fF $ **FLOATING
C1633 out_p.n613 vss 4.05fF $ **FLOATING
C1634 out_p.n614 vss 4.05fF $ **FLOATING
C1635 out_p.n615 vss 4.05fF $ **FLOATING
C1636 out_p.n616 vss 4.15fF $ **FLOATING
C1637 out_p.n617 vss 4.15fF $ **FLOATING
C1638 out_p.n618 vss 4.05fF $ **FLOATING
C1639 out_p.n619 vss 4.05fF $ **FLOATING
C1640 out_p.n620 vss 4.05fF $ **FLOATING
C1641 out_p.n621 vss 3.80fF $ **FLOATING
C1642 out_p.n622 vss 3.85fF $ **FLOATING
C1643 out_p.n623 vss 3.81fF $ **FLOATING
C1644 out_p.n624 vss 3.87fF $ **FLOATING
C1645 out_p.n625 vss 4.05fF $ **FLOATING
C1646 out_p.n626 vss 4.05fF $ **FLOATING
C1647 out_p.n627 vss 4.05fF $ **FLOATING
C1648 out_p.n628 vss 4.15fF $ **FLOATING
C1649 out_p.n629 vss 4.15fF $ **FLOATING
C1650 out_p.n630 vss 4.05fF $ **FLOATING
C1651 out_p.n631 vss 4.05fF $ **FLOATING
C1652 out_p.n632 vss 4.05fF $ **FLOATING
C1653 out_p.n633 vss 3.80fF $ **FLOATING
C1654 out_p.n634 vss 3.85fF $ **FLOATING
C1655 out_p.n635 vss 3.81fF $ **FLOATING
C1656 out_p.n636 vss 3.87fF $ **FLOATING
C1657 out_p.n637 vss 4.05fF $ **FLOATING
C1658 out_p.n638 vss 4.05fF $ **FLOATING
C1659 out_p.n639 vss 4.05fF $ **FLOATING
C1660 out_p.n640 vss 4.15fF $ **FLOATING
C1661 out_p.n641 vss 4.15fF $ **FLOATING
C1662 out_p.n642 vss 4.05fF $ **FLOATING
C1663 out_p.n643 vss 4.05fF $ **FLOATING
C1664 out_p.n644 vss 4.05fF $ **FLOATING
C1665 out_p.n645 vss 3.80fF $ **FLOATING
C1666 out_p.n646 vss 3.85fF $ **FLOATING
C1667 out_p.n647 vss 3.81fF $ **FLOATING
C1668 out_p.n648 vss 3.87fF $ **FLOATING
C1669 out_p.n649 vss 4.05fF $ **FLOATING
C1670 out_p.n650 vss 4.05fF $ **FLOATING
C1671 out_p.n651 vss 4.05fF $ **FLOATING
C1672 out_p.n652 vss 4.15fF $ **FLOATING
C1673 out_p.n653 vss 4.15fF $ **FLOATING
C1674 out_p.n654 vss 4.05fF $ **FLOATING
C1675 out_p.n655 vss 4.05fF $ **FLOATING
C1676 out_p.n656 vss 4.05fF $ **FLOATING
C1677 out_p.n657 vss 3.80fF $ **FLOATING
C1678 out_p.n658 vss 3.85fF $ **FLOATING
C1679 out_p.n659 vss 3.81fF $ **FLOATING
C1680 out_p.n660 vss 3.87fF $ **FLOATING
C1681 out_p.n661 vss 4.05fF $ **FLOATING
C1682 out_p.n662 vss 4.05fF $ **FLOATING
C1683 out_p.n663 vss 4.05fF $ **FLOATING
C1684 out_p.n664 vss 4.15fF $ **FLOATING
C1685 out_p.n665 vss 4.15fF $ **FLOATING
C1686 out_p.n666 vss 4.05fF $ **FLOATING
C1687 out_p.n667 vss 4.05fF $ **FLOATING
C1688 out_p.n668 vss 4.05fF $ **FLOATING
C1689 out_p.n669 vss 3.80fF $ **FLOATING
C1690 out_p.n670 vss 3.85fF $ **FLOATING
C1691 out_p.n671 vss 3.81fF $ **FLOATING
C1692 out_p.n672 vss 3.87fF $ **FLOATING
C1693 out_p.n673 vss 4.05fF $ **FLOATING
C1694 out_p.n674 vss 4.05fF $ **FLOATING
C1695 out_p.n675 vss 4.05fF $ **FLOATING
C1696 out_p.n676 vss 4.15fF $ **FLOATING
C1697 out_p.n677 vss 4.15fF $ **FLOATING
C1698 out_p.n678 vss 4.05fF $ **FLOATING
C1699 out_p.n679 vss 4.05fF $ **FLOATING
C1700 out_p.n680 vss 4.05fF $ **FLOATING
C1701 out_p.n681 vss 3.80fF $ **FLOATING
C1702 out_p.n682 vss 3.85fF $ **FLOATING
C1703 out_p.n683 vss 3.81fF $ **FLOATING
C1704 out_p.n684 vss 3.87fF $ **FLOATING
C1705 out_p.n685 vss 4.05fF $ **FLOATING
C1706 out_p.n686 vss 4.05fF $ **FLOATING
C1707 out_p.n687 vss 4.05fF $ **FLOATING
C1708 out_p.n688 vss 4.15fF $ **FLOATING
C1709 out_p.n689 vss 4.15fF $ **FLOATING
C1710 out_p.n690 vss 4.05fF $ **FLOATING
C1711 out_p.n691 vss 4.05fF $ **FLOATING
C1712 out_p.n692 vss 4.05fF $ **FLOATING
C1713 out_p.n693 vss 3.80fF $ **FLOATING
C1714 out_p.n694 vss 3.85fF $ **FLOATING
C1715 out_p.n695 vss 3.81fF $ **FLOATING
C1716 out_p.n696 vss 3.87fF $ **FLOATING
C1717 out_p.n697 vss 4.05fF $ **FLOATING
C1718 out_p.n698 vss 4.05fF $ **FLOATING
C1719 out_p.n699 vss 4.05fF $ **FLOATING
C1720 out_p.n700 vss 4.15fF $ **FLOATING
C1721 out_p.n701 vss 4.15fF $ **FLOATING
C1722 out_p.n702 vss 4.05fF $ **FLOATING
C1723 out_p.n703 vss 4.05fF $ **FLOATING
C1724 out_p.n704 vss 4.05fF $ **FLOATING
C1725 out_p.n705 vss 3.80fF $ **FLOATING
C1726 out_p.n706 vss 3.85fF $ **FLOATING
C1727 out_p.n707 vss 3.81fF $ **FLOATING
C1728 out_p.n708 vss 3.87fF $ **FLOATING
C1729 out_p.n709 vss 4.05fF $ **FLOATING
C1730 out_p.n710 vss 4.05fF $ **FLOATING
C1731 out_p.n711 vss 4.05fF $ **FLOATING
C1732 out_p.n712 vss 4.15fF $ **FLOATING
C1733 out_p.n713 vss 4.15fF $ **FLOATING
C1734 out_p.n714 vss 4.05fF $ **FLOATING
C1735 out_p.n715 vss 4.05fF $ **FLOATING
C1736 out_p.n716 vss 4.05fF $ **FLOATING
C1737 out_p.n717 vss 3.80fF $ **FLOATING
C1738 out_p.n718 vss 3.85fF $ **FLOATING
C1739 out_p.n719 vss 3.81fF $ **FLOATING
C1740 out_p.n720 vss 3.87fF $ **FLOATING
C1741 out_p.n721 vss 4.05fF $ **FLOATING
C1742 out_p.n722 vss 4.05fF $ **FLOATING
C1743 out_p.n723 vss 4.05fF $ **FLOATING
C1744 out_p.n724 vss 4.15fF $ **FLOATING
C1745 out_p.n725 vss 4.15fF $ **FLOATING
C1746 out_p.n726 vss 4.05fF $ **FLOATING
C1747 out_p.n727 vss 4.05fF $ **FLOATING
C1748 out_p.n728 vss 4.05fF $ **FLOATING
C1749 out_p.n729 vss 3.80fF $ **FLOATING
C1750 out_p.n730 vss 3.85fF $ **FLOATING
C1751 out_p.n731 vss 3.81fF $ **FLOATING
C1752 out_p.n732 vss 3.86fF $ **FLOATING
C1753 out_p.n733 vss 4.05fF $ **FLOATING
C1754 out_p.n734 vss 4.05fF $ **FLOATING
C1755 out_p.n735 vss 4.05fF $ **FLOATING
C1756 out_p.n736 vss 4.15fF $ **FLOATING
C1757 out_p.n737 vss 4.15fF $ **FLOATING
C1758 out_p.n738 vss 4.05fF $ **FLOATING
C1759 out_p.n739 vss 4.05fF $ **FLOATING
C1760 out_p.n740 vss 4.05fF $ **FLOATING
C1761 out_p.n741 vss 3.81fF $ **FLOATING
C1762 out_p.n742 vss 23.47fF $ **FLOATING
C1763 out_p.n743 vss 30.23fF $ **FLOATING
C1764 out_p.n744 vss 30.23fF $ **FLOATING
C1765 out_p.n745 vss 30.23fF $ **FLOATING
C1766 out_p.n746 vss 30.23fF $ **FLOATING
C1767 out_p.n747 vss 30.23fF $ **FLOATING
C1768 out_p.n748 vss 30.23fF $ **FLOATING
C1769 out_p.n749 vss 30.23fF $ **FLOATING
C1770 out_p.n750 vss 30.23fF $ **FLOATING
C1771 out_p.n751 vss 30.23fF $ **FLOATING
C1772 out_p.n752 vss 30.23fF $ **FLOATING
C1773 out_p.n753 vss 30.23fF $ **FLOATING
C1774 out_p.n754 vss 30.23fF $ **FLOATING
C1775 out_p.n755 vss 30.23fF $ **FLOATING
C1776 out_p.n756 vss 30.23fF $ **FLOATING
C1777 out_p.n757 vss 30.23fF $ **FLOATING
C1778 out_p.n758 vss 30.23fF $ **FLOATING
C1779 out_p.n759 vss 30.23fF $ **FLOATING
C1780 out_p.n760 vss 30.23fF $ **FLOATING
C1781 out_p.n761 vss 30.23fF $ **FLOATING
C1782 out_p.n762 vss 30.23fF $ **FLOATING
C1783 out_p.n763 vss 30.23fF $ **FLOATING
C1784 out_p.n764 vss 30.23fF $ **FLOATING
C1785 out_p.n765 vss 30.23fF $ **FLOATING
C1786 out_p.n766 vss 30.23fF $ **FLOATING
C1787 out_p.n767 vss 30.23fF $ **FLOATING
C1788 out_p.n768 vss 30.23fF $ **FLOATING
C1789 out_p.n769 vss 30.23fF $ **FLOATING
C1790 out_p.n770 vss 30.23fF $ **FLOATING
C1791 out_p.n771 vss 30.23fF $ **FLOATING
C1792 out_p.n772 vss 30.23fF $ **FLOATING
C1793 out_p.n773 vss 30.23fF $ **FLOATING
C1794 out_p.n774 vss 30.23fF $ **FLOATING
C1795 out_p.n775 vss 30.23fF $ **FLOATING
C1796 out_p.n776 vss 30.23fF $ **FLOATING
C1797 out_p.n777 vss 30.23fF $ **FLOATING
C1798 out_p.n778 vss 30.23fF $ **FLOATING
C1799 out_p.n779 vss 30.23fF $ **FLOATING
C1800 out_p.n780 vss 30.23fF $ **FLOATING
C1801 out_p.n781 vss 30.23fF $ **FLOATING
C1802 out_p.n782 vss 30.23fF $ **FLOATING
C1803 out_p.n783 vss 30.23fF $ **FLOATING
C1804 out_p.n784 vss 30.23fF $ **FLOATING
C1805 out_p.n785 vss 30.23fF $ **FLOATING
C1806 out_p.n786 vss 30.23fF $ **FLOATING
C1807 out_p.n787 vss 30.23fF $ **FLOATING
C1808 out_p.n788 vss 30.23fF $ **FLOATING
C1809 out_p.n789 vss 30.23fF $ **FLOATING
C1810 out_p.n790 vss 30.23fF $ **FLOATING
C1811 out_p.n791 vss 30.23fF $ **FLOATING
C1812 out_p.n792 vss 30.23fF $ **FLOATING
C1813 out_p.n793 vss 30.23fF $ **FLOATING
C1814 out_p.n794 vss 30.23fF $ **FLOATING
C1815 out_p.n795 vss 30.23fF $ **FLOATING
C1816 out_p.n796 vss 30.23fF $ **FLOATING
C1817 out_p.n797 vss 30.23fF $ **FLOATING
C1818 out_p.n798 vss 30.23fF $ **FLOATING
C1819 out_p.n799 vss 30.23fF $ **FLOATING
C1820 out_p.n800 vss 30.23fF $ **FLOATING
C1821 out_p.n801 vss 28.94fF $ **FLOATING
C1822 out_p.n802 vss 3.85fF $ **FLOATING
C1823 out_p.n803 vss 3.81fF $ **FLOATING
C1824 out_p.n804 vss 3.85fF $ **FLOATING
C1825 out_p.n805 vss 3.81fF $ **FLOATING
C1826 out_p.n806 vss 3.85fF $ **FLOATING
C1827 out_p.n807 vss 3.81fF $ **FLOATING
C1828 out_p.n808 vss 3.85fF $ **FLOATING
C1829 out_p.n809 vss 3.81fF $ **FLOATING
C1830 out_p.n810 vss 3.85fF $ **FLOATING
C1831 out_p.n811 vss 3.81fF $ **FLOATING
C1832 out_p.n812 vss 3.85fF $ **FLOATING
C1833 out_p.n813 vss 3.81fF $ **FLOATING
C1834 out_p.n814 vss 3.85fF $ **FLOATING
C1835 out_p.n815 vss 3.81fF $ **FLOATING
C1836 out_p.n816 vss 3.85fF $ **FLOATING
C1837 out_p.n817 vss 3.81fF $ **FLOATING
C1838 out_p.n818 vss 3.85fF $ **FLOATING
C1839 out_p.n819 vss 3.81fF $ **FLOATING
C1840 out_p.n820 vss 3.85fF $ **FLOATING
C1841 out_p.n821 vss 3.81fF $ **FLOATING
C1842 out_p.n822 vss 3.85fF $ **FLOATING
C1843 out_p.n823 vss 3.81fF $ **FLOATING
C1844 out_p.n824 vss 3.85fF $ **FLOATING
C1845 out_p.n825 vss 3.81fF $ **FLOATING
C1846 out_p.n826 vss 3.85fF $ **FLOATING
C1847 out_p.n827 vss 3.81fF $ **FLOATING
C1848 out_p.n828 vss 3.87fF $ **FLOATING
C1849 out_p.n829 vss 4.05fF $ **FLOATING
C1850 out_p.n830 vss 4.05fF $ **FLOATING
C1851 out_p.n831 vss 4.05fF $ **FLOATING
C1852 out_p.n832 vss 4.15fF $ **FLOATING
C1853 out_p.n833 vss 4.15fF $ **FLOATING
C1854 out_p.n834 vss 4.05fF $ **FLOATING
C1855 out_p.n835 vss 4.05fF $ **FLOATING
C1856 out_p.n836 vss 4.05fF $ **FLOATING
C1857 out_p.n837 vss 3.80fF $ **FLOATING
C1858 out_p.n838 vss 33.39fF $ **FLOATING
C1859 out_p.n839 vss 3.87fF $ **FLOATING
C1860 out_p.n840 vss 4.05fF $ **FLOATING
C1861 out_p.n841 vss 4.05fF $ **FLOATING
C1862 out_p.n842 vss 4.05fF $ **FLOATING
C1863 out_p.n843 vss 4.15fF $ **FLOATING
C1864 out_p.n844 vss 4.15fF $ **FLOATING
C1865 out_p.n845 vss 4.05fF $ **FLOATING
C1866 out_p.n846 vss 4.05fF $ **FLOATING
C1867 out_p.n847 vss 4.05fF $ **FLOATING
C1868 out_p.n848 vss 3.80fF $ **FLOATING
C1869 out_p.n849 vss 30.23fF $ **FLOATING
C1870 out_p.n850 vss 3.87fF $ **FLOATING
C1871 out_p.n851 vss 4.05fF $ **FLOATING
C1872 out_p.n852 vss 4.05fF $ **FLOATING
C1873 out_p.n853 vss 4.05fF $ **FLOATING
C1874 out_p.n854 vss 4.15fF $ **FLOATING
C1875 out_p.n855 vss 4.15fF $ **FLOATING
C1876 out_p.n856 vss 4.05fF $ **FLOATING
C1877 out_p.n857 vss 4.05fF $ **FLOATING
C1878 out_p.n858 vss 4.05fF $ **FLOATING
C1879 out_p.n859 vss 3.80fF $ **FLOATING
C1880 out_p.n860 vss 30.23fF $ **FLOATING
C1881 out_p.n861 vss 3.87fF $ **FLOATING
C1882 out_p.n862 vss 4.05fF $ **FLOATING
C1883 out_p.n863 vss 4.05fF $ **FLOATING
C1884 out_p.n864 vss 4.05fF $ **FLOATING
C1885 out_p.n865 vss 4.15fF $ **FLOATING
C1886 out_p.n866 vss 4.15fF $ **FLOATING
C1887 out_p.n867 vss 4.05fF $ **FLOATING
C1888 out_p.n868 vss 4.05fF $ **FLOATING
C1889 out_p.n869 vss 4.05fF $ **FLOATING
C1890 out_p.n870 vss 3.80fF $ **FLOATING
C1891 out_p.n871 vss 30.23fF $ **FLOATING
C1892 out_p.n872 vss 3.87fF $ **FLOATING
C1893 out_p.n873 vss 4.05fF $ **FLOATING
C1894 out_p.n874 vss 4.05fF $ **FLOATING
C1895 out_p.n875 vss 4.05fF $ **FLOATING
C1896 out_p.n876 vss 4.15fF $ **FLOATING
C1897 out_p.n877 vss 4.15fF $ **FLOATING
C1898 out_p.n878 vss 4.05fF $ **FLOATING
C1899 out_p.n879 vss 4.05fF $ **FLOATING
C1900 out_p.n880 vss 4.05fF $ **FLOATING
C1901 out_p.n881 vss 3.80fF $ **FLOATING
C1902 out_p.n882 vss 30.23fF $ **FLOATING
C1903 out_p.n883 vss 3.87fF $ **FLOATING
C1904 out_p.n884 vss 4.05fF $ **FLOATING
C1905 out_p.n885 vss 4.05fF $ **FLOATING
C1906 out_p.n886 vss 4.05fF $ **FLOATING
C1907 out_p.n887 vss 4.15fF $ **FLOATING
C1908 out_p.n888 vss 4.15fF $ **FLOATING
C1909 out_p.n889 vss 4.05fF $ **FLOATING
C1910 out_p.n890 vss 4.05fF $ **FLOATING
C1911 out_p.n891 vss 4.05fF $ **FLOATING
C1912 out_p.n892 vss 3.80fF $ **FLOATING
C1913 out_p.n893 vss 30.23fF $ **FLOATING
C1914 out_p.n894 vss 3.87fF $ **FLOATING
C1915 out_p.n895 vss 4.05fF $ **FLOATING
C1916 out_p.n896 vss 4.05fF $ **FLOATING
C1917 out_p.n897 vss 4.05fF $ **FLOATING
C1918 out_p.n898 vss 4.15fF $ **FLOATING
C1919 out_p.n899 vss 4.15fF $ **FLOATING
C1920 out_p.n900 vss 4.05fF $ **FLOATING
C1921 out_p.n901 vss 4.05fF $ **FLOATING
C1922 out_p.n902 vss 4.05fF $ **FLOATING
C1923 out_p.n903 vss 3.80fF $ **FLOATING
C1924 out_p.n904 vss 30.23fF $ **FLOATING
C1925 out_p.n905 vss 3.87fF $ **FLOATING
C1926 out_p.n906 vss 4.05fF $ **FLOATING
C1927 out_p.n907 vss 4.05fF $ **FLOATING
C1928 out_p.n908 vss 4.05fF $ **FLOATING
C1929 out_p.n909 vss 4.15fF $ **FLOATING
C1930 out_p.n910 vss 4.15fF $ **FLOATING
C1931 out_p.n911 vss 4.05fF $ **FLOATING
C1932 out_p.n912 vss 4.05fF $ **FLOATING
C1933 out_p.n913 vss 4.05fF $ **FLOATING
C1934 out_p.n914 vss 3.80fF $ **FLOATING
C1935 out_p.n915 vss 30.23fF $ **FLOATING
C1936 out_p.n916 vss 3.87fF $ **FLOATING
C1937 out_p.n917 vss 4.05fF $ **FLOATING
C1938 out_p.n918 vss 4.05fF $ **FLOATING
C1939 out_p.n919 vss 4.05fF $ **FLOATING
C1940 out_p.n920 vss 4.15fF $ **FLOATING
C1941 out_p.n921 vss 4.15fF $ **FLOATING
C1942 out_p.n922 vss 4.05fF $ **FLOATING
C1943 out_p.n923 vss 4.05fF $ **FLOATING
C1944 out_p.n924 vss 4.05fF $ **FLOATING
C1945 out_p.n925 vss 3.80fF $ **FLOATING
C1946 out_p.n926 vss 30.23fF $ **FLOATING
C1947 out_p.n927 vss 3.87fF $ **FLOATING
C1948 out_p.n928 vss 4.05fF $ **FLOATING
C1949 out_p.n929 vss 4.05fF $ **FLOATING
C1950 out_p.n930 vss 4.05fF $ **FLOATING
C1951 out_p.n931 vss 4.15fF $ **FLOATING
C1952 out_p.n932 vss 4.15fF $ **FLOATING
C1953 out_p.n933 vss 4.05fF $ **FLOATING
C1954 out_p.n934 vss 4.05fF $ **FLOATING
C1955 out_p.n935 vss 4.05fF $ **FLOATING
C1956 out_p.n936 vss 3.80fF $ **FLOATING
C1957 out_p.n937 vss 30.23fF $ **FLOATING
C1958 out_p.n938 vss 3.87fF $ **FLOATING
C1959 out_p.n939 vss 4.05fF $ **FLOATING
C1960 out_p.n940 vss 4.05fF $ **FLOATING
C1961 out_p.n941 vss 4.05fF $ **FLOATING
C1962 out_p.n942 vss 4.15fF $ **FLOATING
C1963 out_p.n943 vss 4.15fF $ **FLOATING
C1964 out_p.n944 vss 4.05fF $ **FLOATING
C1965 out_p.n945 vss 4.05fF $ **FLOATING
C1966 out_p.n946 vss 4.05fF $ **FLOATING
C1967 out_p.n947 vss 3.80fF $ **FLOATING
C1968 out_p.n948 vss 30.23fF $ **FLOATING
C1969 out_p.n949 vss 3.87fF $ **FLOATING
C1970 out_p.n950 vss 4.05fF $ **FLOATING
C1971 out_p.n951 vss 4.05fF $ **FLOATING
C1972 out_p.n952 vss 4.05fF $ **FLOATING
C1973 out_p.n953 vss 4.15fF $ **FLOATING
C1974 out_p.n954 vss 4.15fF $ **FLOATING
C1975 out_p.n955 vss 4.05fF $ **FLOATING
C1976 out_p.n956 vss 4.05fF $ **FLOATING
C1977 out_p.n957 vss 4.05fF $ **FLOATING
C1978 out_p.n958 vss 3.80fF $ **FLOATING
C1979 out_p.n959 vss 30.23fF $ **FLOATING
C1980 out_p.n960 vss 3.87fF $ **FLOATING
C1981 out_p.n961 vss 4.05fF $ **FLOATING
C1982 out_p.n962 vss 4.05fF $ **FLOATING
C1983 out_p.n963 vss 4.05fF $ **FLOATING
C1984 out_p.n964 vss 4.15fF $ **FLOATING
C1985 out_p.n965 vss 4.15fF $ **FLOATING
C1986 out_p.n966 vss 4.05fF $ **FLOATING
C1987 out_p.n967 vss 4.05fF $ **FLOATING
C1988 out_p.n968 vss 4.05fF $ **FLOATING
C1989 out_p.n969 vss 3.80fF $ **FLOATING
C1990 out_p.n970 vss 30.23fF $ **FLOATING
C1991 out_p.n971 vss 3.85fF $ **FLOATING
C1992 out_p.n972 vss 3.81fF $ **FLOATING
C1993 out_p.n973 vss 30.94fF $ **FLOATING
C1994 vp_p.n0 vss 1.04fF $ **FLOATING
C1995 vp_p.n76 vss 1.09fF $ **FLOATING
C1996 vp_p.n78 vss 1.03fF $ **FLOATING
C1997 vp_p.n80 vss 1.03fF $ **FLOATING
C1998 vp_p.n82 vss 1.03fF $ **FLOATING
C1999 vp_p.n84 vss 1.03fF $ **FLOATING
C2000 vp_p.n86 vss 1.03fF $ **FLOATING
C2001 vp_p.n88 vss 1.03fF $ **FLOATING
C2002 vp_p.n90 vss 1.03fF $ **FLOATING
C2003 vp_p.n92 vss 1.03fF $ **FLOATING
C2004 vp_p.n94 vss 1.03fF $ **FLOATING
C2005 vp_p.n96 vss 1.03fF $ **FLOATING
C2006 vp_p.n98 vss 1.03fF $ **FLOATING
C2007 vp_p.n100 vss 1.03fF $ **FLOATING
C2008 vp_p.n102 vss 1.03fF $ **FLOATING
C2009 vp_p.n104 vss 1.03fF $ **FLOATING
C2010 vp_p.n106 vss 1.03fF $ **FLOATING
C2011 vp_p.n108 vss 1.03fF $ **FLOATING
C2012 vp_p.n110 vss 1.03fF $ **FLOATING
C2013 vp_p.n112 vss 1.03fF $ **FLOATING
C2014 vp_p.n114 vss 1.03fF $ **FLOATING
C2015 vp_p.n116 vss 1.03fF $ **FLOATING
C2016 vp_p.n118 vss 1.03fF $ **FLOATING
C2017 vp_p.n120 vss 1.03fF $ **FLOATING
C2018 vp_p.n122 vss 1.03fF $ **FLOATING
C2019 vp_p.n124 vss 1.03fF $ **FLOATING
C2020 vp_p.n126 vss 1.03fF $ **FLOATING
C2021 vp_p.n128 vss 1.03fF $ **FLOATING
C2022 vp_p.n130 vss 1.03fF $ **FLOATING
C2023 vp_p.n132 vss 1.03fF $ **FLOATING
C2024 vp_p.n134 vss 1.03fF $ **FLOATING
C2025 vp_p.n136 vss 1.03fF $ **FLOATING
C2026 vp_p.n138 vss 1.03fF $ **FLOATING
C2027 vp_p.n140 vss 1.03fF $ **FLOATING
C2028 vp_p.n142 vss 1.03fF $ **FLOATING
C2029 vp_p.n144 vss 1.03fF $ **FLOATING
C2030 vp_p.n146 vss 1.03fF $ **FLOATING
C2031 vp_p.n148 vss 1.03fF $ **FLOATING
C2032 vp_p.n150 vss 1.03fF $ **FLOATING
C2033 vp_p.n152 vss 1.03fF $ **FLOATING
C2034 vp_p.n154 vss 1.03fF $ **FLOATING
C2035 vp_p.n156 vss 1.03fF $ **FLOATING
C2036 vp_p.n158 vss 1.03fF $ **FLOATING
C2037 vp_p.n160 vss 1.03fF $ **FLOATING
C2038 vp_p.n162 vss 1.03fF $ **FLOATING
C2039 vp_p.n164 vss 1.03fF $ **FLOATING
C2040 vp_p.n166 vss 1.03fF $ **FLOATING
C2041 vp_p.n168 vss 1.03fF $ **FLOATING
C2042 vp_p.n170 vss 1.03fF $ **FLOATING
C2043 vp_p.n172 vss 1.03fF $ **FLOATING
C2044 vp_p.n174 vss 1.03fF $ **FLOATING
C2045 vp_p.n176 vss 1.03fF $ **FLOATING
C2046 vp_p.n178 vss 1.03fF $ **FLOATING
C2047 vp_p.n180 vss 1.03fF $ **FLOATING
C2048 vp_p.n182 vss 1.03fF $ **FLOATING
C2049 vp_p.n184 vss 1.03fF $ **FLOATING
C2050 vp_p.n186 vss 1.03fF $ **FLOATING
C2051 vp_p.n188 vss 1.03fF $ **FLOATING
C2052 vp_p.n190 vss 1.03fF $ **FLOATING
C2053 vp_p.n192 vss 1.03fF $ **FLOATING
C2054 vp_p.n194 vss 1.03fF $ **FLOATING
C2055 vp_p.n196 vss 1.03fF $ **FLOATING
C2056 vp_p.n198 vss 1.03fF $ **FLOATING
C2057 vp_p.n200 vss 1.03fF $ **FLOATING
C2058 vp_p.n202 vss 1.03fF $ **FLOATING
C2059 vp_p.n204 vss 1.03fF $ **FLOATING
C2060 vp_p.n206 vss 1.03fF $ **FLOATING
C2061 vp_p.n208 vss 1.03fF $ **FLOATING
C2062 vp_p.n210 vss 1.03fF $ **FLOATING
C2063 vp_p.n212 vss 1.03fF $ **FLOATING
C2064 vp_p.n214 vss 1.03fF $ **FLOATING
C2065 vp_p.n216 vss 1.03fF $ **FLOATING
C2066 vp_p.n218 vss 1.03fF $ **FLOATING
C2067 vp_p.n220 vss 1.03fF $ **FLOATING
C2068 vp_p.n225 vss 1.09fF $ **FLOATING
C2069 vp_p.n227 vss 1.03fF $ **FLOATING
C2070 vp_p.n229 vss 1.03fF $ **FLOATING
C2071 vp_p.n231 vss 1.03fF $ **FLOATING
C2072 vp_p.n233 vss 1.03fF $ **FLOATING
C2073 vp_p.n235 vss 1.03fF $ **FLOATING
C2074 vp_p.n237 vss 1.03fF $ **FLOATING
C2075 vp_p.n239 vss 1.03fF $ **FLOATING
C2076 vp_p.n241 vss 1.03fF $ **FLOATING
C2077 vp_p.n243 vss 1.03fF $ **FLOATING
C2078 vp_p.n245 vss 1.03fF $ **FLOATING
C2079 vp_p.n247 vss 1.03fF $ **FLOATING
C2080 vp_p.n249 vss 1.03fF $ **FLOATING
C2081 vp_p.n251 vss 1.03fF $ **FLOATING
C2082 vp_p.n253 vss 1.03fF $ **FLOATING
C2083 vp_p.n255 vss 1.03fF $ **FLOATING
C2084 vp_p.n257 vss 1.03fF $ **FLOATING
C2085 vp_p.n259 vss 1.03fF $ **FLOATING
C2086 vp_p.n261 vss 1.03fF $ **FLOATING
C2087 vp_p.n263 vss 1.03fF $ **FLOATING
C2088 vp_p.n265 vss 1.03fF $ **FLOATING
C2089 vp_p.n267 vss 1.03fF $ **FLOATING
C2090 vp_p.n269 vss 1.03fF $ **FLOATING
C2091 vp_p.n271 vss 1.03fF $ **FLOATING
C2092 vp_p.n273 vss 1.03fF $ **FLOATING
C2093 vp_p.n275 vss 1.03fF $ **FLOATING
C2094 vp_p.n277 vss 1.03fF $ **FLOATING
C2095 vp_p.n279 vss 1.03fF $ **FLOATING
C2096 vp_p.n281 vss 1.03fF $ **FLOATING
C2097 vp_p.n283 vss 1.03fF $ **FLOATING
C2098 vp_p.n285 vss 1.03fF $ **FLOATING
C2099 vp_p.n287 vss 1.03fF $ **FLOATING
C2100 vp_p.n289 vss 1.03fF $ **FLOATING
C2101 vp_p.n291 vss 1.03fF $ **FLOATING
C2102 vp_p.n293 vss 1.03fF $ **FLOATING
C2103 vp_p.n295 vss 1.03fF $ **FLOATING
C2104 vp_p.n297 vss 1.03fF $ **FLOATING
C2105 vp_p.n299 vss 1.03fF $ **FLOATING
C2106 vp_p.n301 vss 1.03fF $ **FLOATING
C2107 vp_p.n303 vss 1.03fF $ **FLOATING
C2108 vp_p.n305 vss 1.03fF $ **FLOATING
C2109 vp_p.n307 vss 1.03fF $ **FLOATING
C2110 vp_p.n309 vss 1.03fF $ **FLOATING
C2111 vp_p.n311 vss 1.03fF $ **FLOATING
C2112 vp_p.n313 vss 1.03fF $ **FLOATING
C2113 vp_p.n315 vss 1.03fF $ **FLOATING
C2114 vp_p.n317 vss 1.03fF $ **FLOATING
C2115 vp_p.n319 vss 1.03fF $ **FLOATING
C2116 vp_p.n321 vss 1.03fF $ **FLOATING
C2117 vp_p.n323 vss 1.03fF $ **FLOATING
C2118 vp_p.n325 vss 1.03fF $ **FLOATING
C2119 vp_p.n327 vss 1.03fF $ **FLOATING
C2120 vp_p.n329 vss 1.03fF $ **FLOATING
C2121 vp_p.n331 vss 1.03fF $ **FLOATING
C2122 vp_p.n333 vss 1.03fF $ **FLOATING
C2123 vp_p.n335 vss 1.03fF $ **FLOATING
C2124 vp_p.n337 vss 1.03fF $ **FLOATING
C2125 vp_p.n339 vss 1.03fF $ **FLOATING
C2126 vp_p.n341 vss 1.03fF $ **FLOATING
C2127 vp_p.n343 vss 1.03fF $ **FLOATING
C2128 vp_p.n345 vss 1.03fF $ **FLOATING
C2129 vp_p.n347 vss 1.03fF $ **FLOATING
C2130 vp_p.n349 vss 1.03fF $ **FLOATING
C2131 vp_p.n351 vss 1.03fF $ **FLOATING
C2132 vp_p.n353 vss 1.03fF $ **FLOATING
C2133 vp_p.n355 vss 1.03fF $ **FLOATING
C2134 vp_p.n357 vss 1.03fF $ **FLOATING
C2135 vp_p.n359 vss 1.03fF $ **FLOATING
C2136 vp_p.n361 vss 1.03fF $ **FLOATING
C2137 vp_p.n363 vss 1.03fF $ **FLOATING
C2138 vp_p.n365 vss 1.03fF $ **FLOATING
C2139 vp_p.n367 vss 1.03fF $ **FLOATING
C2140 vp_p.n369 vss 1.03fF $ **FLOATING
C2141 vp_p.n374 vss 1.09fF $ **FLOATING
C2142 vp_p.n376 vss 1.03fF $ **FLOATING
C2143 vp_p.n378 vss 1.03fF $ **FLOATING
C2144 vp_p.n380 vss 1.03fF $ **FLOATING
C2145 vp_p.n382 vss 1.03fF $ **FLOATING
C2146 vp_p.n384 vss 1.03fF $ **FLOATING
C2147 vp_p.n386 vss 1.03fF $ **FLOATING
C2148 vp_p.n388 vss 1.03fF $ **FLOATING
C2149 vp_p.n390 vss 1.03fF $ **FLOATING
C2150 vp_p.n392 vss 1.03fF $ **FLOATING
C2151 vp_p.n394 vss 1.03fF $ **FLOATING
C2152 vp_p.n396 vss 1.03fF $ **FLOATING
C2153 vp_p.n398 vss 1.03fF $ **FLOATING
C2154 vp_p.n400 vss 1.03fF $ **FLOATING
C2155 vp_p.n402 vss 1.03fF $ **FLOATING
C2156 vp_p.n404 vss 1.03fF $ **FLOATING
C2157 vp_p.n406 vss 1.03fF $ **FLOATING
C2158 vp_p.n408 vss 1.03fF $ **FLOATING
C2159 vp_p.n410 vss 1.03fF $ **FLOATING
C2160 vp_p.n412 vss 1.03fF $ **FLOATING
C2161 vp_p.n414 vss 1.03fF $ **FLOATING
C2162 vp_p.n416 vss 1.03fF $ **FLOATING
C2163 vp_p.n418 vss 1.03fF $ **FLOATING
C2164 vp_p.n420 vss 1.03fF $ **FLOATING
C2165 vp_p.n422 vss 1.03fF $ **FLOATING
C2166 vp_p.n424 vss 1.03fF $ **FLOATING
C2167 vp_p.n426 vss 1.03fF $ **FLOATING
C2168 vp_p.n428 vss 1.03fF $ **FLOATING
C2169 vp_p.n430 vss 1.03fF $ **FLOATING
C2170 vp_p.n432 vss 1.03fF $ **FLOATING
C2171 vp_p.n434 vss 1.03fF $ **FLOATING
C2172 vp_p.n436 vss 1.03fF $ **FLOATING
C2173 vp_p.n438 vss 1.03fF $ **FLOATING
C2174 vp_p.n440 vss 1.03fF $ **FLOATING
C2175 vp_p.n442 vss 1.03fF $ **FLOATING
C2176 vp_p.n444 vss 1.03fF $ **FLOATING
C2177 vp_p.n446 vss 1.03fF $ **FLOATING
C2178 vp_p.n448 vss 1.03fF $ **FLOATING
C2179 vp_p.n450 vss 1.03fF $ **FLOATING
C2180 vp_p.n452 vss 1.03fF $ **FLOATING
C2181 vp_p.n454 vss 1.03fF $ **FLOATING
C2182 vp_p.n456 vss 1.03fF $ **FLOATING
C2183 vp_p.n458 vss 1.03fF $ **FLOATING
C2184 vp_p.n460 vss 1.03fF $ **FLOATING
C2185 vp_p.n462 vss 1.03fF $ **FLOATING
C2186 vp_p.n464 vss 1.03fF $ **FLOATING
C2187 vp_p.n466 vss 1.03fF $ **FLOATING
C2188 vp_p.n468 vss 1.03fF $ **FLOATING
C2189 vp_p.n470 vss 1.03fF $ **FLOATING
C2190 vp_p.n472 vss 1.03fF $ **FLOATING
C2191 vp_p.n474 vss 1.03fF $ **FLOATING
C2192 vp_p.n476 vss 1.03fF $ **FLOATING
C2193 vp_p.n478 vss 1.03fF $ **FLOATING
C2194 vp_p.n480 vss 1.03fF $ **FLOATING
C2195 vp_p.n482 vss 1.03fF $ **FLOATING
C2196 vp_p.n484 vss 1.03fF $ **FLOATING
C2197 vp_p.n486 vss 1.03fF $ **FLOATING
C2198 vp_p.n488 vss 1.03fF $ **FLOATING
C2199 vp_p.n490 vss 1.03fF $ **FLOATING
C2200 vp_p.n492 vss 1.03fF $ **FLOATING
C2201 vp_p.n494 vss 1.03fF $ **FLOATING
C2202 vp_p.n496 vss 1.03fF $ **FLOATING
C2203 vp_p.n498 vss 1.03fF $ **FLOATING
C2204 vp_p.n500 vss 1.03fF $ **FLOATING
C2205 vp_p.n502 vss 1.03fF $ **FLOATING
C2206 vp_p.n504 vss 1.03fF $ **FLOATING
C2207 vp_p.n506 vss 1.03fF $ **FLOATING
C2208 vp_p.n508 vss 1.03fF $ **FLOATING
C2209 vp_p.n510 vss 1.03fF $ **FLOATING
C2210 vp_p.n512 vss 1.03fF $ **FLOATING
C2211 vp_p.n514 vss 1.03fF $ **FLOATING
C2212 vp_p.n516 vss 1.03fF $ **FLOATING
C2213 vp_p.n518 vss 1.03fF $ **FLOATING
C2214 vp_p.n523 vss 1.09fF $ **FLOATING
C2215 vp_p.n525 vss 1.03fF $ **FLOATING
C2216 vp_p.n527 vss 1.03fF $ **FLOATING
C2217 vp_p.n529 vss 1.03fF $ **FLOATING
C2218 vp_p.n531 vss 1.03fF $ **FLOATING
C2219 vp_p.n533 vss 1.03fF $ **FLOATING
C2220 vp_p.n535 vss 1.03fF $ **FLOATING
C2221 vp_p.n537 vss 1.03fF $ **FLOATING
C2222 vp_p.n539 vss 1.03fF $ **FLOATING
C2223 vp_p.n541 vss 1.03fF $ **FLOATING
C2224 vp_p.n543 vss 1.03fF $ **FLOATING
C2225 vp_p.n545 vss 1.03fF $ **FLOATING
C2226 vp_p.n547 vss 1.03fF $ **FLOATING
C2227 vp_p.n549 vss 1.03fF $ **FLOATING
C2228 vp_p.n551 vss 1.03fF $ **FLOATING
C2229 vp_p.n553 vss 1.03fF $ **FLOATING
C2230 vp_p.n555 vss 1.03fF $ **FLOATING
C2231 vp_p.n557 vss 1.03fF $ **FLOATING
C2232 vp_p.n559 vss 1.03fF $ **FLOATING
C2233 vp_p.n561 vss 1.03fF $ **FLOATING
C2234 vp_p.n563 vss 1.03fF $ **FLOATING
C2235 vp_p.n565 vss 1.03fF $ **FLOATING
C2236 vp_p.n567 vss 1.03fF $ **FLOATING
C2237 vp_p.n569 vss 1.03fF $ **FLOATING
C2238 vp_p.n571 vss 1.03fF $ **FLOATING
C2239 vp_p.n573 vss 1.03fF $ **FLOATING
C2240 vp_p.n575 vss 1.03fF $ **FLOATING
C2241 vp_p.n577 vss 1.03fF $ **FLOATING
C2242 vp_p.n579 vss 1.03fF $ **FLOATING
C2243 vp_p.n581 vss 1.03fF $ **FLOATING
C2244 vp_p.n583 vss 1.03fF $ **FLOATING
C2245 vp_p.n585 vss 1.03fF $ **FLOATING
C2246 vp_p.n587 vss 1.03fF $ **FLOATING
C2247 vp_p.n589 vss 1.03fF $ **FLOATING
C2248 vp_p.n591 vss 1.03fF $ **FLOATING
C2249 vp_p.n593 vss 1.03fF $ **FLOATING
C2250 vp_p.n595 vss 1.03fF $ **FLOATING
C2251 vp_p.n597 vss 1.03fF $ **FLOATING
C2252 vp_p.n599 vss 1.03fF $ **FLOATING
C2253 vp_p.n601 vss 1.03fF $ **FLOATING
C2254 vp_p.n603 vss 1.03fF $ **FLOATING
C2255 vp_p.n605 vss 1.03fF $ **FLOATING
C2256 vp_p.n607 vss 1.03fF $ **FLOATING
C2257 vp_p.n609 vss 1.03fF $ **FLOATING
C2258 vp_p.n611 vss 1.03fF $ **FLOATING
C2259 vp_p.n613 vss 1.03fF $ **FLOATING
C2260 vp_p.n615 vss 1.03fF $ **FLOATING
C2261 vp_p.n617 vss 1.03fF $ **FLOATING
C2262 vp_p.n619 vss 1.03fF $ **FLOATING
C2263 vp_p.n621 vss 1.03fF $ **FLOATING
C2264 vp_p.n623 vss 1.03fF $ **FLOATING
C2265 vp_p.n625 vss 1.03fF $ **FLOATING
C2266 vp_p.n627 vss 1.03fF $ **FLOATING
C2267 vp_p.n629 vss 1.03fF $ **FLOATING
C2268 vp_p.n631 vss 1.03fF $ **FLOATING
C2269 vp_p.n633 vss 1.03fF $ **FLOATING
C2270 vp_p.n635 vss 1.03fF $ **FLOATING
C2271 vp_p.n637 vss 1.03fF $ **FLOATING
C2272 vp_p.n639 vss 1.03fF $ **FLOATING
C2273 vp_p.n641 vss 1.03fF $ **FLOATING
C2274 vp_p.n643 vss 1.03fF $ **FLOATING
C2275 vp_p.n645 vss 1.03fF $ **FLOATING
C2276 vp_p.n647 vss 1.03fF $ **FLOATING
C2277 vp_p.n649 vss 1.03fF $ **FLOATING
C2278 vp_p.n651 vss 1.03fF $ **FLOATING
C2279 vp_p.n653 vss 1.03fF $ **FLOATING
C2280 vp_p.n655 vss 1.03fF $ **FLOATING
C2281 vp_p.n657 vss 1.03fF $ **FLOATING
C2282 vp_p.n659 vss 1.03fF $ **FLOATING
C2283 vp_p.n661 vss 1.03fF $ **FLOATING
C2284 vp_p.n663 vss 1.03fF $ **FLOATING
C2285 vp_p.n665 vss 1.03fF $ **FLOATING
C2286 vp_p.n667 vss 1.03fF $ **FLOATING
C2287 vp_p.n670 vss 1.10fF $ **FLOATING
C2288 vp_p.n743 vss 1.92fF $ **FLOATING
C2289 vp_p.n744 vss 18.53fF $ **FLOATING
C2290 vp_p.n745 vss 7.33fF $ **FLOATING
C2291 vp_p.n746 vss 13.12fF $ **FLOATING
C2292 vp_p.n747 vss 13.09fF $ **FLOATING
C2293 vp_p.n748 vss 7.69fF $ **FLOATING
C2294 vp_p.n749 vss 1.05fF $ **FLOATING
C2295 vp_p.n825 vss 1.09fF $ **FLOATING
C2296 vp_p.n827 vss 1.03fF $ **FLOATING
C2297 vp_p.n829 vss 1.03fF $ **FLOATING
C2298 vp_p.n831 vss 1.03fF $ **FLOATING
C2299 vp_p.n833 vss 1.03fF $ **FLOATING
C2300 vp_p.n835 vss 1.03fF $ **FLOATING
C2301 vp_p.n837 vss 1.03fF $ **FLOATING
C2302 vp_p.n839 vss 1.03fF $ **FLOATING
C2303 vp_p.n841 vss 1.03fF $ **FLOATING
C2304 vp_p.n843 vss 1.03fF $ **FLOATING
C2305 vp_p.n845 vss 1.03fF $ **FLOATING
C2306 vp_p.n847 vss 1.03fF $ **FLOATING
C2307 vp_p.n849 vss 1.03fF $ **FLOATING
C2308 vp_p.n851 vss 1.03fF $ **FLOATING
C2309 vp_p.n853 vss 1.03fF $ **FLOATING
C2310 vp_p.n855 vss 1.03fF $ **FLOATING
C2311 vp_p.n857 vss 1.03fF $ **FLOATING
C2312 vp_p.n859 vss 1.03fF $ **FLOATING
C2313 vp_p.n861 vss 1.03fF $ **FLOATING
C2314 vp_p.n863 vss 1.03fF $ **FLOATING
C2315 vp_p.n865 vss 1.03fF $ **FLOATING
C2316 vp_p.n867 vss 1.03fF $ **FLOATING
C2317 vp_p.n869 vss 1.03fF $ **FLOATING
C2318 vp_p.n871 vss 1.03fF $ **FLOATING
C2319 vp_p.n873 vss 1.03fF $ **FLOATING
C2320 vp_p.n875 vss 1.03fF $ **FLOATING
C2321 vp_p.n877 vss 1.03fF $ **FLOATING
C2322 vp_p.n879 vss 1.03fF $ **FLOATING
C2323 vp_p.n881 vss 1.03fF $ **FLOATING
C2324 vp_p.n883 vss 1.03fF $ **FLOATING
C2325 vp_p.n885 vss 1.03fF $ **FLOATING
C2326 vp_p.n887 vss 1.03fF $ **FLOATING
C2327 vp_p.n889 vss 1.03fF $ **FLOATING
C2328 vp_p.n891 vss 1.03fF $ **FLOATING
C2329 vp_p.n893 vss 1.03fF $ **FLOATING
C2330 vp_p.n895 vss 1.03fF $ **FLOATING
C2331 vp_p.n897 vss 1.03fF $ **FLOATING
C2332 vp_p.n899 vss 1.03fF $ **FLOATING
C2333 vp_p.n901 vss 1.03fF $ **FLOATING
C2334 vp_p.n903 vss 1.03fF $ **FLOATING
C2335 vp_p.n905 vss 1.03fF $ **FLOATING
C2336 vp_p.n907 vss 1.03fF $ **FLOATING
C2337 vp_p.n909 vss 1.03fF $ **FLOATING
C2338 vp_p.n911 vss 1.03fF $ **FLOATING
C2339 vp_p.n913 vss 1.03fF $ **FLOATING
C2340 vp_p.n915 vss 1.03fF $ **FLOATING
C2341 vp_p.n917 vss 1.03fF $ **FLOATING
C2342 vp_p.n919 vss 1.03fF $ **FLOATING
C2343 vp_p.n921 vss 1.03fF $ **FLOATING
C2344 vp_p.n923 vss 1.03fF $ **FLOATING
C2345 vp_p.n925 vss 1.03fF $ **FLOATING
C2346 vp_p.n927 vss 1.03fF $ **FLOATING
C2347 vp_p.n929 vss 1.03fF $ **FLOATING
C2348 vp_p.n931 vss 1.03fF $ **FLOATING
C2349 vp_p.n933 vss 1.03fF $ **FLOATING
C2350 vp_p.n935 vss 1.03fF $ **FLOATING
C2351 vp_p.n937 vss 1.03fF $ **FLOATING
C2352 vp_p.n939 vss 1.03fF $ **FLOATING
C2353 vp_p.n941 vss 1.03fF $ **FLOATING
C2354 vp_p.n943 vss 1.03fF $ **FLOATING
C2355 vp_p.n945 vss 1.03fF $ **FLOATING
C2356 vp_p.n947 vss 1.03fF $ **FLOATING
C2357 vp_p.n949 vss 1.03fF $ **FLOATING
C2358 vp_p.n951 vss 1.03fF $ **FLOATING
C2359 vp_p.n953 vss 1.03fF $ **FLOATING
C2360 vp_p.n955 vss 1.03fF $ **FLOATING
C2361 vp_p.n957 vss 1.03fF $ **FLOATING
C2362 vp_p.n959 vss 1.03fF $ **FLOATING
C2363 vp_p.n961 vss 1.03fF $ **FLOATING
C2364 vp_p.n963 vss 1.03fF $ **FLOATING
C2365 vp_p.n965 vss 1.03fF $ **FLOATING
C2366 vp_p.n967 vss 1.03fF $ **FLOATING
C2367 vp_p.n969 vss 1.03fF $ **FLOATING
C2368 vp_p.n974 vss 1.09fF $ **FLOATING
C2369 vp_p.n976 vss 1.03fF $ **FLOATING
C2370 vp_p.n978 vss 1.03fF $ **FLOATING
C2371 vp_p.n980 vss 1.03fF $ **FLOATING
C2372 vp_p.n982 vss 1.03fF $ **FLOATING
C2373 vp_p.n984 vss 1.03fF $ **FLOATING
C2374 vp_p.n986 vss 1.03fF $ **FLOATING
C2375 vp_p.n988 vss 1.03fF $ **FLOATING
C2376 vp_p.n990 vss 1.03fF $ **FLOATING
C2377 vp_p.n992 vss 1.03fF $ **FLOATING
C2378 vp_p.n994 vss 1.03fF $ **FLOATING
C2379 vp_p.n996 vss 1.03fF $ **FLOATING
C2380 vp_p.n998 vss 1.03fF $ **FLOATING
C2381 vp_p.n1000 vss 1.03fF $ **FLOATING
C2382 vp_p.n1002 vss 1.03fF $ **FLOATING
C2383 vp_p.n1004 vss 1.03fF $ **FLOATING
C2384 vp_p.n1006 vss 1.03fF $ **FLOATING
C2385 vp_p.n1008 vss 1.03fF $ **FLOATING
C2386 vp_p.n1010 vss 1.03fF $ **FLOATING
C2387 vp_p.n1012 vss 1.03fF $ **FLOATING
C2388 vp_p.n1014 vss 1.03fF $ **FLOATING
C2389 vp_p.n1016 vss 1.03fF $ **FLOATING
C2390 vp_p.n1018 vss 1.03fF $ **FLOATING
C2391 vp_p.n1020 vss 1.03fF $ **FLOATING
C2392 vp_p.n1022 vss 1.03fF $ **FLOATING
C2393 vp_p.n1024 vss 1.03fF $ **FLOATING
C2394 vp_p.n1026 vss 1.03fF $ **FLOATING
C2395 vp_p.n1028 vss 1.03fF $ **FLOATING
C2396 vp_p.n1030 vss 1.03fF $ **FLOATING
C2397 vp_p.n1032 vss 1.03fF $ **FLOATING
C2398 vp_p.n1034 vss 1.03fF $ **FLOATING
C2399 vp_p.n1036 vss 1.03fF $ **FLOATING
C2400 vp_p.n1038 vss 1.03fF $ **FLOATING
C2401 vp_p.n1040 vss 1.03fF $ **FLOATING
C2402 vp_p.n1042 vss 1.03fF $ **FLOATING
C2403 vp_p.n1044 vss 1.03fF $ **FLOATING
C2404 vp_p.n1046 vss 1.03fF $ **FLOATING
C2405 vp_p.n1048 vss 1.03fF $ **FLOATING
C2406 vp_p.n1050 vss 1.03fF $ **FLOATING
C2407 vp_p.n1052 vss 1.03fF $ **FLOATING
C2408 vp_p.n1054 vss 1.03fF $ **FLOATING
C2409 vp_p.n1056 vss 1.03fF $ **FLOATING
C2410 vp_p.n1058 vss 1.03fF $ **FLOATING
C2411 vp_p.n1060 vss 1.03fF $ **FLOATING
C2412 vp_p.n1062 vss 1.03fF $ **FLOATING
C2413 vp_p.n1064 vss 1.03fF $ **FLOATING
C2414 vp_p.n1066 vss 1.03fF $ **FLOATING
C2415 vp_p.n1068 vss 1.03fF $ **FLOATING
C2416 vp_p.n1070 vss 1.03fF $ **FLOATING
C2417 vp_p.n1072 vss 1.03fF $ **FLOATING
C2418 vp_p.n1074 vss 1.03fF $ **FLOATING
C2419 vp_p.n1076 vss 1.03fF $ **FLOATING
C2420 vp_p.n1078 vss 1.03fF $ **FLOATING
C2421 vp_p.n1080 vss 1.03fF $ **FLOATING
C2422 vp_p.n1082 vss 1.03fF $ **FLOATING
C2423 vp_p.n1084 vss 1.03fF $ **FLOATING
C2424 vp_p.n1086 vss 1.03fF $ **FLOATING
C2425 vp_p.n1088 vss 1.03fF $ **FLOATING
C2426 vp_p.n1090 vss 1.03fF $ **FLOATING
C2427 vp_p.n1092 vss 1.03fF $ **FLOATING
C2428 vp_p.n1094 vss 1.03fF $ **FLOATING
C2429 vp_p.n1096 vss 1.03fF $ **FLOATING
C2430 vp_p.n1098 vss 1.03fF $ **FLOATING
C2431 vp_p.n1100 vss 1.03fF $ **FLOATING
C2432 vp_p.n1102 vss 1.03fF $ **FLOATING
C2433 vp_p.n1104 vss 1.03fF $ **FLOATING
C2434 vp_p.n1106 vss 1.03fF $ **FLOATING
C2435 vp_p.n1108 vss 1.03fF $ **FLOATING
C2436 vp_p.n1110 vss 1.03fF $ **FLOATING
C2437 vp_p.n1112 vss 1.03fF $ **FLOATING
C2438 vp_p.n1114 vss 1.03fF $ **FLOATING
C2439 vp_p.n1116 vss 1.03fF $ **FLOATING
C2440 vp_p.n1118 vss 1.03fF $ **FLOATING
C2441 vp_p.n1123 vss 1.09fF $ **FLOATING
C2442 vp_p.n1125 vss 1.03fF $ **FLOATING
C2443 vp_p.n1127 vss 1.03fF $ **FLOATING
C2444 vp_p.n1129 vss 1.03fF $ **FLOATING
C2445 vp_p.n1131 vss 1.03fF $ **FLOATING
C2446 vp_p.n1133 vss 1.03fF $ **FLOATING
C2447 vp_p.n1135 vss 1.03fF $ **FLOATING
C2448 vp_p.n1137 vss 1.03fF $ **FLOATING
C2449 vp_p.n1139 vss 1.03fF $ **FLOATING
C2450 vp_p.n1141 vss 1.03fF $ **FLOATING
C2451 vp_p.n1143 vss 1.03fF $ **FLOATING
C2452 vp_p.n1145 vss 1.03fF $ **FLOATING
C2453 vp_p.n1147 vss 1.03fF $ **FLOATING
C2454 vp_p.n1149 vss 1.03fF $ **FLOATING
C2455 vp_p.n1151 vss 1.03fF $ **FLOATING
C2456 vp_p.n1153 vss 1.03fF $ **FLOATING
C2457 vp_p.n1155 vss 1.03fF $ **FLOATING
C2458 vp_p.n1157 vss 1.03fF $ **FLOATING
C2459 vp_p.n1159 vss 1.03fF $ **FLOATING
C2460 vp_p.n1161 vss 1.03fF $ **FLOATING
C2461 vp_p.n1163 vss 1.03fF $ **FLOATING
C2462 vp_p.n1165 vss 1.03fF $ **FLOATING
C2463 vp_p.n1167 vss 1.03fF $ **FLOATING
C2464 vp_p.n1169 vss 1.03fF $ **FLOATING
C2465 vp_p.n1171 vss 1.03fF $ **FLOATING
C2466 vp_p.n1173 vss 1.03fF $ **FLOATING
C2467 vp_p.n1175 vss 1.03fF $ **FLOATING
C2468 vp_p.n1177 vss 1.03fF $ **FLOATING
C2469 vp_p.n1179 vss 1.03fF $ **FLOATING
C2470 vp_p.n1181 vss 1.03fF $ **FLOATING
C2471 vp_p.n1183 vss 1.03fF $ **FLOATING
C2472 vp_p.n1185 vss 1.03fF $ **FLOATING
C2473 vp_p.n1187 vss 1.03fF $ **FLOATING
C2474 vp_p.n1189 vss 1.03fF $ **FLOATING
C2475 vp_p.n1191 vss 1.03fF $ **FLOATING
C2476 vp_p.n1193 vss 1.03fF $ **FLOATING
C2477 vp_p.n1195 vss 1.03fF $ **FLOATING
C2478 vp_p.n1197 vss 1.03fF $ **FLOATING
C2479 vp_p.n1199 vss 1.03fF $ **FLOATING
C2480 vp_p.n1201 vss 1.03fF $ **FLOATING
C2481 vp_p.n1203 vss 1.03fF $ **FLOATING
C2482 vp_p.n1205 vss 1.03fF $ **FLOATING
C2483 vp_p.n1207 vss 1.03fF $ **FLOATING
C2484 vp_p.n1209 vss 1.03fF $ **FLOATING
C2485 vp_p.n1211 vss 1.03fF $ **FLOATING
C2486 vp_p.n1213 vss 1.03fF $ **FLOATING
C2487 vp_p.n1215 vss 1.03fF $ **FLOATING
C2488 vp_p.n1217 vss 1.03fF $ **FLOATING
C2489 vp_p.n1219 vss 1.03fF $ **FLOATING
C2490 vp_p.n1221 vss 1.03fF $ **FLOATING
C2491 vp_p.n1223 vss 1.03fF $ **FLOATING
C2492 vp_p.n1225 vss 1.03fF $ **FLOATING
C2493 vp_p.n1227 vss 1.03fF $ **FLOATING
C2494 vp_p.n1229 vss 1.03fF $ **FLOATING
C2495 vp_p.n1231 vss 1.03fF $ **FLOATING
C2496 vp_p.n1233 vss 1.03fF $ **FLOATING
C2497 vp_p.n1235 vss 1.03fF $ **FLOATING
C2498 vp_p.n1237 vss 1.03fF $ **FLOATING
C2499 vp_p.n1239 vss 1.03fF $ **FLOATING
C2500 vp_p.n1241 vss 1.03fF $ **FLOATING
C2501 vp_p.n1243 vss 1.03fF $ **FLOATING
C2502 vp_p.n1245 vss 1.03fF $ **FLOATING
C2503 vp_p.n1247 vss 1.03fF $ **FLOATING
C2504 vp_p.n1249 vss 1.03fF $ **FLOATING
C2505 vp_p.n1251 vss 1.03fF $ **FLOATING
C2506 vp_p.n1253 vss 1.03fF $ **FLOATING
C2507 vp_p.n1255 vss 1.03fF $ **FLOATING
C2508 vp_p.n1257 vss 1.03fF $ **FLOATING
C2509 vp_p.n1259 vss 1.03fF $ **FLOATING
C2510 vp_p.n1261 vss 1.03fF $ **FLOATING
C2511 vp_p.n1263 vss 1.03fF $ **FLOATING
C2512 vp_p.n1265 vss 1.03fF $ **FLOATING
C2513 vp_p.n1267 vss 1.03fF $ **FLOATING
C2514 vp_p.n1272 vss 1.09fF $ **FLOATING
C2515 vp_p.n1274 vss 1.03fF $ **FLOATING
C2516 vp_p.n1276 vss 1.03fF $ **FLOATING
C2517 vp_p.n1278 vss 1.03fF $ **FLOATING
C2518 vp_p.n1280 vss 1.03fF $ **FLOATING
C2519 vp_p.n1282 vss 1.03fF $ **FLOATING
C2520 vp_p.n1284 vss 1.03fF $ **FLOATING
C2521 vp_p.n1286 vss 1.03fF $ **FLOATING
C2522 vp_p.n1288 vss 1.03fF $ **FLOATING
C2523 vp_p.n1290 vss 1.03fF $ **FLOATING
C2524 vp_p.n1292 vss 1.03fF $ **FLOATING
C2525 vp_p.n1294 vss 1.03fF $ **FLOATING
C2526 vp_p.n1296 vss 1.03fF $ **FLOATING
C2527 vp_p.n1298 vss 1.03fF $ **FLOATING
C2528 vp_p.n1300 vss 1.03fF $ **FLOATING
C2529 vp_p.n1302 vss 1.03fF $ **FLOATING
C2530 vp_p.n1304 vss 1.03fF $ **FLOATING
C2531 vp_p.n1306 vss 1.03fF $ **FLOATING
C2532 vp_p.n1308 vss 1.03fF $ **FLOATING
C2533 vp_p.n1310 vss 1.03fF $ **FLOATING
C2534 vp_p.n1312 vss 1.03fF $ **FLOATING
C2535 vp_p.n1314 vss 1.03fF $ **FLOATING
C2536 vp_p.n1316 vss 1.03fF $ **FLOATING
C2537 vp_p.n1318 vss 1.03fF $ **FLOATING
C2538 vp_p.n1320 vss 1.03fF $ **FLOATING
C2539 vp_p.n1322 vss 1.03fF $ **FLOATING
C2540 vp_p.n1324 vss 1.03fF $ **FLOATING
C2541 vp_p.n1326 vss 1.03fF $ **FLOATING
C2542 vp_p.n1328 vss 1.03fF $ **FLOATING
C2543 vp_p.n1330 vss 1.03fF $ **FLOATING
C2544 vp_p.n1332 vss 1.03fF $ **FLOATING
C2545 vp_p.n1334 vss 1.03fF $ **FLOATING
C2546 vp_p.n1336 vss 1.03fF $ **FLOATING
C2547 vp_p.n1338 vss 1.03fF $ **FLOATING
C2548 vp_p.n1340 vss 1.03fF $ **FLOATING
C2549 vp_p.n1342 vss 1.03fF $ **FLOATING
C2550 vp_p.n1344 vss 1.03fF $ **FLOATING
C2551 vp_p.n1346 vss 1.03fF $ **FLOATING
C2552 vp_p.n1348 vss 1.03fF $ **FLOATING
C2553 vp_p.n1350 vss 1.03fF $ **FLOATING
C2554 vp_p.n1352 vss 1.03fF $ **FLOATING
C2555 vp_p.n1354 vss 1.03fF $ **FLOATING
C2556 vp_p.n1356 vss 1.03fF $ **FLOATING
C2557 vp_p.n1358 vss 1.03fF $ **FLOATING
C2558 vp_p.n1360 vss 1.03fF $ **FLOATING
C2559 vp_p.n1362 vss 1.03fF $ **FLOATING
C2560 vp_p.n1364 vss 1.03fF $ **FLOATING
C2561 vp_p.n1366 vss 1.03fF $ **FLOATING
C2562 vp_p.n1368 vss 1.03fF $ **FLOATING
C2563 vp_p.n1370 vss 1.03fF $ **FLOATING
C2564 vp_p.n1372 vss 1.03fF $ **FLOATING
C2565 vp_p.n1374 vss 1.03fF $ **FLOATING
C2566 vp_p.n1376 vss 1.03fF $ **FLOATING
C2567 vp_p.n1378 vss 1.03fF $ **FLOATING
C2568 vp_p.n1380 vss 1.03fF $ **FLOATING
C2569 vp_p.n1382 vss 1.03fF $ **FLOATING
C2570 vp_p.n1384 vss 1.03fF $ **FLOATING
C2571 vp_p.n1386 vss 1.03fF $ **FLOATING
C2572 vp_p.n1388 vss 1.03fF $ **FLOATING
C2573 vp_p.n1390 vss 1.03fF $ **FLOATING
C2574 vp_p.n1392 vss 1.03fF $ **FLOATING
C2575 vp_p.n1394 vss 1.03fF $ **FLOATING
C2576 vp_p.n1396 vss 1.03fF $ **FLOATING
C2577 vp_p.n1398 vss 1.03fF $ **FLOATING
C2578 vp_p.n1400 vss 1.03fF $ **FLOATING
C2579 vp_p.n1402 vss 1.03fF $ **FLOATING
C2580 vp_p.n1404 vss 1.03fF $ **FLOATING
C2581 vp_p.n1406 vss 1.03fF $ **FLOATING
C2582 vp_p.n1408 vss 1.03fF $ **FLOATING
C2583 vp_p.n1410 vss 1.03fF $ **FLOATING
C2584 vp_p.n1412 vss 1.03fF $ **FLOATING
C2585 vp_p.n1414 vss 1.03fF $ **FLOATING
C2586 vp_p.n1416 vss 1.03fF $ **FLOATING
C2587 vp_p.n1419 vss 1.04fF $ **FLOATING
C2588 vp_p.n1492 vss 1.34fF $ **FLOATING
C2589 vp_p.n1493 vss 19.04fF $ **FLOATING
C2590 vp_p.n1494 vss 13.65fF $ **FLOATING
C2591 vp_p.n1495 vss 13.44fF $ **FLOATING
C2592 vp_p.n1496 vss 13.30fF $ **FLOATING
C2593 vp_p.n1497 vss 6.61fF $ **FLOATING
C2594 out_n.n0 vss 3.87fF $ **FLOATING
C2595 out_n.n1 vss 4.05fF $ **FLOATING
C2596 out_n.n2 vss 4.05fF $ **FLOATING
C2597 out_n.n3 vss 4.05fF $ **FLOATING
C2598 out_n.n4 vss 4.15fF $ **FLOATING
C2599 out_n.n5 vss 4.15fF $ **FLOATING
C2600 out_n.n6 vss 4.05fF $ **FLOATING
C2601 out_n.n7 vss 4.05fF $ **FLOATING
C2602 out_n.n8 vss 4.05fF $ **FLOATING
C2603 out_n.n9 vss 3.80fF $ **FLOATING
C2604 out_n.n10 vss 3.87fF $ **FLOATING
C2605 out_n.n11 vss 4.05fF $ **FLOATING
C2606 out_n.n12 vss 4.05fF $ **FLOATING
C2607 out_n.n13 vss 4.05fF $ **FLOATING
C2608 out_n.n14 vss 4.15fF $ **FLOATING
C2609 out_n.n15 vss 4.15fF $ **FLOATING
C2610 out_n.n16 vss 4.05fF $ **FLOATING
C2611 out_n.n17 vss 4.05fF $ **FLOATING
C2612 out_n.n18 vss 4.05fF $ **FLOATING
C2613 out_n.n19 vss 3.80fF $ **FLOATING
C2614 out_n.n20 vss 3.87fF $ **FLOATING
C2615 out_n.n21 vss 4.05fF $ **FLOATING
C2616 out_n.n22 vss 4.05fF $ **FLOATING
C2617 out_n.n23 vss 4.05fF $ **FLOATING
C2618 out_n.n24 vss 4.15fF $ **FLOATING
C2619 out_n.n25 vss 4.15fF $ **FLOATING
C2620 out_n.n26 vss 4.05fF $ **FLOATING
C2621 out_n.n27 vss 4.05fF $ **FLOATING
C2622 out_n.n28 vss 4.05fF $ **FLOATING
C2623 out_n.n29 vss 3.80fF $ **FLOATING
C2624 out_n.n30 vss 3.87fF $ **FLOATING
C2625 out_n.n31 vss 4.05fF $ **FLOATING
C2626 out_n.n32 vss 4.05fF $ **FLOATING
C2627 out_n.n33 vss 4.05fF $ **FLOATING
C2628 out_n.n34 vss 4.15fF $ **FLOATING
C2629 out_n.n35 vss 4.15fF $ **FLOATING
C2630 out_n.n36 vss 4.05fF $ **FLOATING
C2631 out_n.n37 vss 4.05fF $ **FLOATING
C2632 out_n.n38 vss 4.05fF $ **FLOATING
C2633 out_n.n39 vss 3.80fF $ **FLOATING
C2634 out_n.n40 vss 3.87fF $ **FLOATING
C2635 out_n.n41 vss 4.05fF $ **FLOATING
C2636 out_n.n42 vss 4.05fF $ **FLOATING
C2637 out_n.n43 vss 4.05fF $ **FLOATING
C2638 out_n.n44 vss 4.15fF $ **FLOATING
C2639 out_n.n45 vss 4.15fF $ **FLOATING
C2640 out_n.n46 vss 4.05fF $ **FLOATING
C2641 out_n.n47 vss 4.05fF $ **FLOATING
C2642 out_n.n48 vss 4.05fF $ **FLOATING
C2643 out_n.n49 vss 3.80fF $ **FLOATING
C2644 out_n.n50 vss 3.87fF $ **FLOATING
C2645 out_n.n51 vss 4.05fF $ **FLOATING
C2646 out_n.n52 vss 4.05fF $ **FLOATING
C2647 out_n.n53 vss 4.05fF $ **FLOATING
C2648 out_n.n54 vss 4.15fF $ **FLOATING
C2649 out_n.n55 vss 4.15fF $ **FLOATING
C2650 out_n.n56 vss 4.05fF $ **FLOATING
C2651 out_n.n57 vss 4.05fF $ **FLOATING
C2652 out_n.n58 vss 4.05fF $ **FLOATING
C2653 out_n.n59 vss 3.80fF $ **FLOATING
C2654 out_n.n60 vss 3.87fF $ **FLOATING
C2655 out_n.n61 vss 4.05fF $ **FLOATING
C2656 out_n.n62 vss 4.05fF $ **FLOATING
C2657 out_n.n63 vss 4.05fF $ **FLOATING
C2658 out_n.n64 vss 4.15fF $ **FLOATING
C2659 out_n.n65 vss 4.15fF $ **FLOATING
C2660 out_n.n66 vss 4.05fF $ **FLOATING
C2661 out_n.n67 vss 4.05fF $ **FLOATING
C2662 out_n.n68 vss 4.05fF $ **FLOATING
C2663 out_n.n69 vss 3.80fF $ **FLOATING
C2664 out_n.n70 vss 3.87fF $ **FLOATING
C2665 out_n.n71 vss 4.05fF $ **FLOATING
C2666 out_n.n72 vss 4.05fF $ **FLOATING
C2667 out_n.n73 vss 4.05fF $ **FLOATING
C2668 out_n.n74 vss 4.15fF $ **FLOATING
C2669 out_n.n75 vss 4.15fF $ **FLOATING
C2670 out_n.n76 vss 4.05fF $ **FLOATING
C2671 out_n.n77 vss 4.05fF $ **FLOATING
C2672 out_n.n78 vss 4.05fF $ **FLOATING
C2673 out_n.n79 vss 3.80fF $ **FLOATING
C2674 out_n.n80 vss 3.87fF $ **FLOATING
C2675 out_n.n81 vss 4.05fF $ **FLOATING
C2676 out_n.n82 vss 4.05fF $ **FLOATING
C2677 out_n.n83 vss 4.05fF $ **FLOATING
C2678 out_n.n84 vss 4.15fF $ **FLOATING
C2679 out_n.n85 vss 4.15fF $ **FLOATING
C2680 out_n.n86 vss 4.05fF $ **FLOATING
C2681 out_n.n87 vss 4.05fF $ **FLOATING
C2682 out_n.n88 vss 4.05fF $ **FLOATING
C2683 out_n.n89 vss 3.80fF $ **FLOATING
C2684 out_n.n90 vss 3.87fF $ **FLOATING
C2685 out_n.n91 vss 4.05fF $ **FLOATING
C2686 out_n.n92 vss 4.05fF $ **FLOATING
C2687 out_n.n93 vss 4.05fF $ **FLOATING
C2688 out_n.n94 vss 4.15fF $ **FLOATING
C2689 out_n.n95 vss 4.15fF $ **FLOATING
C2690 out_n.n96 vss 4.05fF $ **FLOATING
C2691 out_n.n97 vss 4.05fF $ **FLOATING
C2692 out_n.n98 vss 4.05fF $ **FLOATING
C2693 out_n.n99 vss 3.80fF $ **FLOATING
C2694 out_n.n100 vss 3.87fF $ **FLOATING
C2695 out_n.n101 vss 4.05fF $ **FLOATING
C2696 out_n.n102 vss 4.05fF $ **FLOATING
C2697 out_n.n103 vss 4.05fF $ **FLOATING
C2698 out_n.n104 vss 4.15fF $ **FLOATING
C2699 out_n.n105 vss 4.15fF $ **FLOATING
C2700 out_n.n106 vss 4.05fF $ **FLOATING
C2701 out_n.n107 vss 4.05fF $ **FLOATING
C2702 out_n.n108 vss 4.05fF $ **FLOATING
C2703 out_n.n109 vss 3.80fF $ **FLOATING
C2704 out_n.n110 vss 3.87fF $ **FLOATING
C2705 out_n.n111 vss 4.05fF $ **FLOATING
C2706 out_n.n112 vss 4.05fF $ **FLOATING
C2707 out_n.n113 vss 4.05fF $ **FLOATING
C2708 out_n.n114 vss 4.15fF $ **FLOATING
C2709 out_n.n115 vss 4.15fF $ **FLOATING
C2710 out_n.n116 vss 4.05fF $ **FLOATING
C2711 out_n.n117 vss 4.05fF $ **FLOATING
C2712 out_n.n118 vss 4.05fF $ **FLOATING
C2713 out_n.n119 vss 3.80fF $ **FLOATING
C2714 out_n.n120 vss 3.87fF $ **FLOATING
C2715 out_n.n121 vss 4.05fF $ **FLOATING
C2716 out_n.n122 vss 4.05fF $ **FLOATING
C2717 out_n.n123 vss 4.05fF $ **FLOATING
C2718 out_n.n124 vss 4.15fF $ **FLOATING
C2719 out_n.n125 vss 4.15fF $ **FLOATING
C2720 out_n.n126 vss 4.05fF $ **FLOATING
C2721 out_n.n127 vss 4.05fF $ **FLOATING
C2722 out_n.n128 vss 4.05fF $ **FLOATING
C2723 out_n.n129 vss 3.80fF $ **FLOATING
C2724 out_n.n130 vss 3.87fF $ **FLOATING
C2725 out_n.n131 vss 4.05fF $ **FLOATING
C2726 out_n.n132 vss 4.05fF $ **FLOATING
C2727 out_n.n133 vss 4.05fF $ **FLOATING
C2728 out_n.n134 vss 4.15fF $ **FLOATING
C2729 out_n.n135 vss 4.15fF $ **FLOATING
C2730 out_n.n136 vss 4.05fF $ **FLOATING
C2731 out_n.n137 vss 4.05fF $ **FLOATING
C2732 out_n.n138 vss 4.05fF $ **FLOATING
C2733 out_n.n139 vss 3.80fF $ **FLOATING
C2734 out_n.n140 vss 3.87fF $ **FLOATING
C2735 out_n.n141 vss 4.05fF $ **FLOATING
C2736 out_n.n142 vss 4.05fF $ **FLOATING
C2737 out_n.n143 vss 4.05fF $ **FLOATING
C2738 out_n.n144 vss 4.15fF $ **FLOATING
C2739 out_n.n145 vss 4.15fF $ **FLOATING
C2740 out_n.n146 vss 4.05fF $ **FLOATING
C2741 out_n.n147 vss 4.05fF $ **FLOATING
C2742 out_n.n148 vss 4.05fF $ **FLOATING
C2743 out_n.n149 vss 3.80fF $ **FLOATING
C2744 out_n.n150 vss 3.87fF $ **FLOATING
C2745 out_n.n151 vss 4.05fF $ **FLOATING
C2746 out_n.n152 vss 4.05fF $ **FLOATING
C2747 out_n.n153 vss 4.05fF $ **FLOATING
C2748 out_n.n154 vss 4.15fF $ **FLOATING
C2749 out_n.n155 vss 4.15fF $ **FLOATING
C2750 out_n.n156 vss 4.05fF $ **FLOATING
C2751 out_n.n157 vss 4.05fF $ **FLOATING
C2752 out_n.n158 vss 4.05fF $ **FLOATING
C2753 out_n.n159 vss 3.80fF $ **FLOATING
C2754 out_n.n160 vss 3.87fF $ **FLOATING
C2755 out_n.n161 vss 4.05fF $ **FLOATING
C2756 out_n.n162 vss 4.05fF $ **FLOATING
C2757 out_n.n163 vss 4.05fF $ **FLOATING
C2758 out_n.n164 vss 4.15fF $ **FLOATING
C2759 out_n.n165 vss 4.15fF $ **FLOATING
C2760 out_n.n166 vss 4.05fF $ **FLOATING
C2761 out_n.n167 vss 4.05fF $ **FLOATING
C2762 out_n.n168 vss 4.05fF $ **FLOATING
C2763 out_n.n169 vss 3.80fF $ **FLOATING
C2764 out_n.n170 vss 3.87fF $ **FLOATING
C2765 out_n.n171 vss 4.05fF $ **FLOATING
C2766 out_n.n172 vss 4.05fF $ **FLOATING
C2767 out_n.n173 vss 4.05fF $ **FLOATING
C2768 out_n.n174 vss 4.15fF $ **FLOATING
C2769 out_n.n175 vss 4.15fF $ **FLOATING
C2770 out_n.n176 vss 4.05fF $ **FLOATING
C2771 out_n.n177 vss 4.05fF $ **FLOATING
C2772 out_n.n178 vss 4.05fF $ **FLOATING
C2773 out_n.n179 vss 3.80fF $ **FLOATING
C2774 out_n.n180 vss 3.87fF $ **FLOATING
C2775 out_n.n181 vss 4.05fF $ **FLOATING
C2776 out_n.n182 vss 4.05fF $ **FLOATING
C2777 out_n.n183 vss 4.05fF $ **FLOATING
C2778 out_n.n184 vss 4.15fF $ **FLOATING
C2779 out_n.n185 vss 4.15fF $ **FLOATING
C2780 out_n.n186 vss 4.05fF $ **FLOATING
C2781 out_n.n187 vss 4.05fF $ **FLOATING
C2782 out_n.n188 vss 4.05fF $ **FLOATING
C2783 out_n.n189 vss 3.80fF $ **FLOATING
C2784 out_n.n190 vss 3.87fF $ **FLOATING
C2785 out_n.n191 vss 4.05fF $ **FLOATING
C2786 out_n.n192 vss 4.05fF $ **FLOATING
C2787 out_n.n193 vss 4.05fF $ **FLOATING
C2788 out_n.n194 vss 4.15fF $ **FLOATING
C2789 out_n.n195 vss 4.15fF $ **FLOATING
C2790 out_n.n196 vss 4.05fF $ **FLOATING
C2791 out_n.n197 vss 4.05fF $ **FLOATING
C2792 out_n.n198 vss 4.05fF $ **FLOATING
C2793 out_n.n199 vss 3.80fF $ **FLOATING
C2794 out_n.n200 vss 3.87fF $ **FLOATING
C2795 out_n.n201 vss 4.05fF $ **FLOATING
C2796 out_n.n202 vss 4.05fF $ **FLOATING
C2797 out_n.n203 vss 4.05fF $ **FLOATING
C2798 out_n.n204 vss 4.15fF $ **FLOATING
C2799 out_n.n205 vss 4.15fF $ **FLOATING
C2800 out_n.n206 vss 4.05fF $ **FLOATING
C2801 out_n.n207 vss 4.05fF $ **FLOATING
C2802 out_n.n208 vss 4.05fF $ **FLOATING
C2803 out_n.n209 vss 3.80fF $ **FLOATING
C2804 out_n.n210 vss 3.87fF $ **FLOATING
C2805 out_n.n211 vss 4.05fF $ **FLOATING
C2806 out_n.n212 vss 4.05fF $ **FLOATING
C2807 out_n.n213 vss 4.05fF $ **FLOATING
C2808 out_n.n214 vss 4.15fF $ **FLOATING
C2809 out_n.n215 vss 4.15fF $ **FLOATING
C2810 out_n.n216 vss 4.05fF $ **FLOATING
C2811 out_n.n217 vss 4.05fF $ **FLOATING
C2812 out_n.n218 vss 4.05fF $ **FLOATING
C2813 out_n.n219 vss 3.80fF $ **FLOATING
C2814 out_n.n220 vss 3.87fF $ **FLOATING
C2815 out_n.n221 vss 4.05fF $ **FLOATING
C2816 out_n.n222 vss 4.05fF $ **FLOATING
C2817 out_n.n223 vss 4.05fF $ **FLOATING
C2818 out_n.n224 vss 4.15fF $ **FLOATING
C2819 out_n.n225 vss 4.15fF $ **FLOATING
C2820 out_n.n226 vss 4.05fF $ **FLOATING
C2821 out_n.n227 vss 4.05fF $ **FLOATING
C2822 out_n.n228 vss 4.05fF $ **FLOATING
C2823 out_n.n229 vss 3.80fF $ **FLOATING
C2824 out_n.n230 vss 3.87fF $ **FLOATING
C2825 out_n.n231 vss 4.05fF $ **FLOATING
C2826 out_n.n232 vss 4.05fF $ **FLOATING
C2827 out_n.n233 vss 4.05fF $ **FLOATING
C2828 out_n.n234 vss 4.15fF $ **FLOATING
C2829 out_n.n235 vss 4.15fF $ **FLOATING
C2830 out_n.n236 vss 4.05fF $ **FLOATING
C2831 out_n.n237 vss 4.05fF $ **FLOATING
C2832 out_n.n238 vss 4.05fF $ **FLOATING
C2833 out_n.n239 vss 3.80fF $ **FLOATING
C2834 out_n.n240 vss 3.87fF $ **FLOATING
C2835 out_n.n241 vss 4.05fF $ **FLOATING
C2836 out_n.n242 vss 4.05fF $ **FLOATING
C2837 out_n.n243 vss 4.05fF $ **FLOATING
C2838 out_n.n244 vss 4.15fF $ **FLOATING
C2839 out_n.n245 vss 4.15fF $ **FLOATING
C2840 out_n.n246 vss 4.05fF $ **FLOATING
C2841 out_n.n247 vss 4.05fF $ **FLOATING
C2842 out_n.n248 vss 4.05fF $ **FLOATING
C2843 out_n.n249 vss 3.80fF $ **FLOATING
C2844 out_n.n250 vss 3.87fF $ **FLOATING
C2845 out_n.n251 vss 4.05fF $ **FLOATING
C2846 out_n.n252 vss 4.05fF $ **FLOATING
C2847 out_n.n253 vss 4.05fF $ **FLOATING
C2848 out_n.n254 vss 4.15fF $ **FLOATING
C2849 out_n.n255 vss 4.15fF $ **FLOATING
C2850 out_n.n256 vss 4.05fF $ **FLOATING
C2851 out_n.n257 vss 4.05fF $ **FLOATING
C2852 out_n.n258 vss 4.05fF $ **FLOATING
C2853 out_n.n259 vss 3.80fF $ **FLOATING
C2854 out_n.n260 vss 3.87fF $ **FLOATING
C2855 out_n.n261 vss 4.05fF $ **FLOATING
C2856 out_n.n262 vss 4.05fF $ **FLOATING
C2857 out_n.n263 vss 4.05fF $ **FLOATING
C2858 out_n.n264 vss 4.15fF $ **FLOATING
C2859 out_n.n265 vss 4.15fF $ **FLOATING
C2860 out_n.n266 vss 4.05fF $ **FLOATING
C2861 out_n.n267 vss 4.05fF $ **FLOATING
C2862 out_n.n268 vss 4.05fF $ **FLOATING
C2863 out_n.n269 vss 3.80fF $ **FLOATING
C2864 out_n.n270 vss 3.87fF $ **FLOATING
C2865 out_n.n271 vss 4.05fF $ **FLOATING
C2866 out_n.n272 vss 4.05fF $ **FLOATING
C2867 out_n.n273 vss 4.05fF $ **FLOATING
C2868 out_n.n274 vss 4.15fF $ **FLOATING
C2869 out_n.n275 vss 4.15fF $ **FLOATING
C2870 out_n.n276 vss 4.05fF $ **FLOATING
C2871 out_n.n277 vss 4.05fF $ **FLOATING
C2872 out_n.n278 vss 4.05fF $ **FLOATING
C2873 out_n.n279 vss 3.80fF $ **FLOATING
C2874 out_n.n280 vss 3.87fF $ **FLOATING
C2875 out_n.n281 vss 4.05fF $ **FLOATING
C2876 out_n.n282 vss 4.05fF $ **FLOATING
C2877 out_n.n283 vss 4.05fF $ **FLOATING
C2878 out_n.n284 vss 4.15fF $ **FLOATING
C2879 out_n.n285 vss 4.15fF $ **FLOATING
C2880 out_n.n286 vss 4.05fF $ **FLOATING
C2881 out_n.n287 vss 4.05fF $ **FLOATING
C2882 out_n.n288 vss 4.05fF $ **FLOATING
C2883 out_n.n289 vss 3.80fF $ **FLOATING
C2884 out_n.n290 vss 3.87fF $ **FLOATING
C2885 out_n.n291 vss 4.05fF $ **FLOATING
C2886 out_n.n292 vss 4.05fF $ **FLOATING
C2887 out_n.n293 vss 4.05fF $ **FLOATING
C2888 out_n.n294 vss 4.15fF $ **FLOATING
C2889 out_n.n295 vss 4.15fF $ **FLOATING
C2890 out_n.n296 vss 4.05fF $ **FLOATING
C2891 out_n.n297 vss 4.05fF $ **FLOATING
C2892 out_n.n298 vss 4.05fF $ **FLOATING
C2893 out_n.n299 vss 3.80fF $ **FLOATING
C2894 out_n.n300 vss 3.87fF $ **FLOATING
C2895 out_n.n301 vss 4.05fF $ **FLOATING
C2896 out_n.n302 vss 4.05fF $ **FLOATING
C2897 out_n.n303 vss 4.05fF $ **FLOATING
C2898 out_n.n304 vss 4.15fF $ **FLOATING
C2899 out_n.n305 vss 4.15fF $ **FLOATING
C2900 out_n.n306 vss 4.05fF $ **FLOATING
C2901 out_n.n307 vss 4.05fF $ **FLOATING
C2902 out_n.n308 vss 4.05fF $ **FLOATING
C2903 out_n.n309 vss 3.80fF $ **FLOATING
C2904 out_n.n310 vss 3.87fF $ **FLOATING
C2905 out_n.n311 vss 4.05fF $ **FLOATING
C2906 out_n.n312 vss 4.05fF $ **FLOATING
C2907 out_n.n313 vss 4.05fF $ **FLOATING
C2908 out_n.n314 vss 4.15fF $ **FLOATING
C2909 out_n.n315 vss 4.15fF $ **FLOATING
C2910 out_n.n316 vss 4.05fF $ **FLOATING
C2911 out_n.n317 vss 4.05fF $ **FLOATING
C2912 out_n.n318 vss 4.05fF $ **FLOATING
C2913 out_n.n319 vss 3.80fF $ **FLOATING
C2914 out_n.n320 vss 3.87fF $ **FLOATING
C2915 out_n.n321 vss 4.05fF $ **FLOATING
C2916 out_n.n322 vss 4.05fF $ **FLOATING
C2917 out_n.n323 vss 4.05fF $ **FLOATING
C2918 out_n.n324 vss 4.15fF $ **FLOATING
C2919 out_n.n325 vss 4.15fF $ **FLOATING
C2920 out_n.n326 vss 4.05fF $ **FLOATING
C2921 out_n.n327 vss 4.05fF $ **FLOATING
C2922 out_n.n328 vss 4.05fF $ **FLOATING
C2923 out_n.n329 vss 3.80fF $ **FLOATING
C2924 out_n.n330 vss 3.87fF $ **FLOATING
C2925 out_n.n331 vss 4.05fF $ **FLOATING
C2926 out_n.n332 vss 4.05fF $ **FLOATING
C2927 out_n.n333 vss 4.05fF $ **FLOATING
C2928 out_n.n334 vss 4.15fF $ **FLOATING
C2929 out_n.n335 vss 4.15fF $ **FLOATING
C2930 out_n.n336 vss 4.05fF $ **FLOATING
C2931 out_n.n337 vss 4.05fF $ **FLOATING
C2932 out_n.n338 vss 4.05fF $ **FLOATING
C2933 out_n.n339 vss 3.80fF $ **FLOATING
C2934 out_n.n340 vss 3.87fF $ **FLOATING
C2935 out_n.n341 vss 4.05fF $ **FLOATING
C2936 out_n.n342 vss 4.05fF $ **FLOATING
C2937 out_n.n343 vss 4.05fF $ **FLOATING
C2938 out_n.n344 vss 4.15fF $ **FLOATING
C2939 out_n.n345 vss 4.15fF $ **FLOATING
C2940 out_n.n346 vss 4.05fF $ **FLOATING
C2941 out_n.n347 vss 4.05fF $ **FLOATING
C2942 out_n.n348 vss 4.05fF $ **FLOATING
C2943 out_n.n349 vss 3.80fF $ **FLOATING
C2944 out_n.n350 vss 3.87fF $ **FLOATING
C2945 out_n.n351 vss 4.05fF $ **FLOATING
C2946 out_n.n352 vss 4.05fF $ **FLOATING
C2947 out_n.n353 vss 4.05fF $ **FLOATING
C2948 out_n.n354 vss 4.15fF $ **FLOATING
C2949 out_n.n355 vss 4.15fF $ **FLOATING
C2950 out_n.n356 vss 4.05fF $ **FLOATING
C2951 out_n.n357 vss 4.05fF $ **FLOATING
C2952 out_n.n358 vss 4.05fF $ **FLOATING
C2953 out_n.n359 vss 3.80fF $ **FLOATING
C2954 out_n.n360 vss 3.87fF $ **FLOATING
C2955 out_n.n361 vss 4.05fF $ **FLOATING
C2956 out_n.n362 vss 4.05fF $ **FLOATING
C2957 out_n.n363 vss 4.05fF $ **FLOATING
C2958 out_n.n364 vss 4.15fF $ **FLOATING
C2959 out_n.n365 vss 4.15fF $ **FLOATING
C2960 out_n.n366 vss 4.05fF $ **FLOATING
C2961 out_n.n367 vss 4.05fF $ **FLOATING
C2962 out_n.n368 vss 4.05fF $ **FLOATING
C2963 out_n.n369 vss 3.80fF $ **FLOATING
C2964 out_n.n370 vss 3.87fF $ **FLOATING
C2965 out_n.n371 vss 4.05fF $ **FLOATING
C2966 out_n.n372 vss 4.05fF $ **FLOATING
C2967 out_n.n373 vss 4.05fF $ **FLOATING
C2968 out_n.n374 vss 4.15fF $ **FLOATING
C2969 out_n.n375 vss 4.15fF $ **FLOATING
C2970 out_n.n376 vss 4.05fF $ **FLOATING
C2971 out_n.n377 vss 4.05fF $ **FLOATING
C2972 out_n.n378 vss 4.05fF $ **FLOATING
C2973 out_n.n379 vss 3.80fF $ **FLOATING
C2974 out_n.n380 vss 3.87fF $ **FLOATING
C2975 out_n.n381 vss 4.05fF $ **FLOATING
C2976 out_n.n382 vss 4.05fF $ **FLOATING
C2977 out_n.n383 vss 4.05fF $ **FLOATING
C2978 out_n.n384 vss 4.15fF $ **FLOATING
C2979 out_n.n385 vss 4.15fF $ **FLOATING
C2980 out_n.n386 vss 4.05fF $ **FLOATING
C2981 out_n.n387 vss 4.05fF $ **FLOATING
C2982 out_n.n388 vss 4.05fF $ **FLOATING
C2983 out_n.n389 vss 3.80fF $ **FLOATING
C2984 out_n.n390 vss 3.87fF $ **FLOATING
C2985 out_n.n391 vss 4.05fF $ **FLOATING
C2986 out_n.n392 vss 4.05fF $ **FLOATING
C2987 out_n.n393 vss 4.05fF $ **FLOATING
C2988 out_n.n394 vss 4.15fF $ **FLOATING
C2989 out_n.n395 vss 4.15fF $ **FLOATING
C2990 out_n.n396 vss 4.05fF $ **FLOATING
C2991 out_n.n397 vss 4.05fF $ **FLOATING
C2992 out_n.n398 vss 4.05fF $ **FLOATING
C2993 out_n.n399 vss 3.80fF $ **FLOATING
C2994 out_n.n400 vss 3.87fF $ **FLOATING
C2995 out_n.n401 vss 4.05fF $ **FLOATING
C2996 out_n.n402 vss 4.05fF $ **FLOATING
C2997 out_n.n403 vss 4.05fF $ **FLOATING
C2998 out_n.n404 vss 4.15fF $ **FLOATING
C2999 out_n.n405 vss 4.15fF $ **FLOATING
C3000 out_n.n406 vss 4.05fF $ **FLOATING
C3001 out_n.n407 vss 4.05fF $ **FLOATING
C3002 out_n.n408 vss 4.05fF $ **FLOATING
C3003 out_n.n409 vss 3.80fF $ **FLOATING
C3004 out_n.n410 vss 3.87fF $ **FLOATING
C3005 out_n.n411 vss 4.05fF $ **FLOATING
C3006 out_n.n412 vss 4.05fF $ **FLOATING
C3007 out_n.n413 vss 4.05fF $ **FLOATING
C3008 out_n.n414 vss 4.15fF $ **FLOATING
C3009 out_n.n415 vss 4.15fF $ **FLOATING
C3010 out_n.n416 vss 4.05fF $ **FLOATING
C3011 out_n.n417 vss 4.05fF $ **FLOATING
C3012 out_n.n418 vss 4.05fF $ **FLOATING
C3013 out_n.n419 vss 3.80fF $ **FLOATING
C3014 out_n.n420 vss 3.87fF $ **FLOATING
C3015 out_n.n421 vss 4.05fF $ **FLOATING
C3016 out_n.n422 vss 4.05fF $ **FLOATING
C3017 out_n.n423 vss 4.05fF $ **FLOATING
C3018 out_n.n424 vss 4.15fF $ **FLOATING
C3019 out_n.n425 vss 4.15fF $ **FLOATING
C3020 out_n.n426 vss 4.05fF $ **FLOATING
C3021 out_n.n427 vss 4.05fF $ **FLOATING
C3022 out_n.n428 vss 4.05fF $ **FLOATING
C3023 out_n.n429 vss 3.80fF $ **FLOATING
C3024 out_n.n430 vss 3.87fF $ **FLOATING
C3025 out_n.n431 vss 4.05fF $ **FLOATING
C3026 out_n.n432 vss 4.05fF $ **FLOATING
C3027 out_n.n433 vss 4.05fF $ **FLOATING
C3028 out_n.n434 vss 4.15fF $ **FLOATING
C3029 out_n.n435 vss 4.15fF $ **FLOATING
C3030 out_n.n436 vss 4.05fF $ **FLOATING
C3031 out_n.n437 vss 4.05fF $ **FLOATING
C3032 out_n.n438 vss 4.05fF $ **FLOATING
C3033 out_n.n439 vss 3.80fF $ **FLOATING
C3034 out_n.n440 vss 3.87fF $ **FLOATING
C3035 out_n.n441 vss 4.05fF $ **FLOATING
C3036 out_n.n442 vss 4.05fF $ **FLOATING
C3037 out_n.n443 vss 4.05fF $ **FLOATING
C3038 out_n.n444 vss 4.15fF $ **FLOATING
C3039 out_n.n445 vss 4.15fF $ **FLOATING
C3040 out_n.n446 vss 4.05fF $ **FLOATING
C3041 out_n.n447 vss 4.05fF $ **FLOATING
C3042 out_n.n448 vss 4.05fF $ **FLOATING
C3043 out_n.n449 vss 3.80fF $ **FLOATING
C3044 out_n.n450 vss 3.87fF $ **FLOATING
C3045 out_n.n451 vss 4.05fF $ **FLOATING
C3046 out_n.n452 vss 4.05fF $ **FLOATING
C3047 out_n.n453 vss 4.05fF $ **FLOATING
C3048 out_n.n454 vss 4.15fF $ **FLOATING
C3049 out_n.n455 vss 4.15fF $ **FLOATING
C3050 out_n.n456 vss 4.05fF $ **FLOATING
C3051 out_n.n457 vss 4.05fF $ **FLOATING
C3052 out_n.n458 vss 4.05fF $ **FLOATING
C3053 out_n.n459 vss 3.80fF $ **FLOATING
C3054 out_n.n460 vss 3.87fF $ **FLOATING
C3055 out_n.n461 vss 4.05fF $ **FLOATING
C3056 out_n.n462 vss 4.05fF $ **FLOATING
C3057 out_n.n463 vss 4.05fF $ **FLOATING
C3058 out_n.n464 vss 4.15fF $ **FLOATING
C3059 out_n.n465 vss 4.15fF $ **FLOATING
C3060 out_n.n466 vss 4.05fF $ **FLOATING
C3061 out_n.n467 vss 4.05fF $ **FLOATING
C3062 out_n.n468 vss 4.05fF $ **FLOATING
C3063 out_n.n469 vss 3.80fF $ **FLOATING
C3064 out_n.n470 vss 3.87fF $ **FLOATING
C3065 out_n.n471 vss 4.05fF $ **FLOATING
C3066 out_n.n472 vss 4.05fF $ **FLOATING
C3067 out_n.n473 vss 4.05fF $ **FLOATING
C3068 out_n.n474 vss 4.15fF $ **FLOATING
C3069 out_n.n475 vss 4.15fF $ **FLOATING
C3070 out_n.n476 vss 4.05fF $ **FLOATING
C3071 out_n.n477 vss 4.05fF $ **FLOATING
C3072 out_n.n478 vss 4.05fF $ **FLOATING
C3073 out_n.n479 vss 3.80fF $ **FLOATING
C3074 out_n.n480 vss 3.87fF $ **FLOATING
C3075 out_n.n481 vss 4.05fF $ **FLOATING
C3076 out_n.n482 vss 4.05fF $ **FLOATING
C3077 out_n.n483 vss 4.05fF $ **FLOATING
C3078 out_n.n484 vss 4.15fF $ **FLOATING
C3079 out_n.n485 vss 4.15fF $ **FLOATING
C3080 out_n.n486 vss 4.05fF $ **FLOATING
C3081 out_n.n487 vss 4.05fF $ **FLOATING
C3082 out_n.n488 vss 4.05fF $ **FLOATING
C3083 out_n.n489 vss 3.80fF $ **FLOATING
C3084 out_n.n490 vss 3.87fF $ **FLOATING
C3085 out_n.n491 vss 4.05fF $ **FLOATING
C3086 out_n.n492 vss 4.05fF $ **FLOATING
C3087 out_n.n493 vss 4.05fF $ **FLOATING
C3088 out_n.n494 vss 4.15fF $ **FLOATING
C3089 out_n.n495 vss 4.15fF $ **FLOATING
C3090 out_n.n496 vss 4.05fF $ **FLOATING
C3091 out_n.n497 vss 4.05fF $ **FLOATING
C3092 out_n.n498 vss 4.05fF $ **FLOATING
C3093 out_n.n499 vss 3.80fF $ **FLOATING
C3094 out_n.n500 vss 3.87fF $ **FLOATING
C3095 out_n.n501 vss 4.05fF $ **FLOATING
C3096 out_n.n502 vss 4.05fF $ **FLOATING
C3097 out_n.n503 vss 4.05fF $ **FLOATING
C3098 out_n.n504 vss 4.15fF $ **FLOATING
C3099 out_n.n505 vss 4.15fF $ **FLOATING
C3100 out_n.n506 vss 4.05fF $ **FLOATING
C3101 out_n.n507 vss 4.05fF $ **FLOATING
C3102 out_n.n508 vss 4.05fF $ **FLOATING
C3103 out_n.n509 vss 3.80fF $ **FLOATING
C3104 out_n.n510 vss 3.87fF $ **FLOATING
C3105 out_n.n511 vss 4.05fF $ **FLOATING
C3106 out_n.n512 vss 4.05fF $ **FLOATING
C3107 out_n.n513 vss 4.05fF $ **FLOATING
C3108 out_n.n514 vss 4.15fF $ **FLOATING
C3109 out_n.n515 vss 4.15fF $ **FLOATING
C3110 out_n.n516 vss 4.05fF $ **FLOATING
C3111 out_n.n517 vss 4.05fF $ **FLOATING
C3112 out_n.n518 vss 4.05fF $ **FLOATING
C3113 out_n.n519 vss 3.80fF $ **FLOATING
C3114 out_n.n520 vss 3.87fF $ **FLOATING
C3115 out_n.n521 vss 4.05fF $ **FLOATING
C3116 out_n.n522 vss 4.05fF $ **FLOATING
C3117 out_n.n523 vss 4.05fF $ **FLOATING
C3118 out_n.n524 vss 4.15fF $ **FLOATING
C3119 out_n.n525 vss 4.15fF $ **FLOATING
C3120 out_n.n526 vss 4.05fF $ **FLOATING
C3121 out_n.n527 vss 4.05fF $ **FLOATING
C3122 out_n.n528 vss 4.05fF $ **FLOATING
C3123 out_n.n529 vss 3.80fF $ **FLOATING
C3124 out_n.n530 vss 3.87fF $ **FLOATING
C3125 out_n.n531 vss 4.05fF $ **FLOATING
C3126 out_n.n532 vss 4.05fF $ **FLOATING
C3127 out_n.n533 vss 4.05fF $ **FLOATING
C3128 out_n.n534 vss 4.15fF $ **FLOATING
C3129 out_n.n535 vss 4.15fF $ **FLOATING
C3130 out_n.n536 vss 4.05fF $ **FLOATING
C3131 out_n.n537 vss 4.05fF $ **FLOATING
C3132 out_n.n538 vss 4.05fF $ **FLOATING
C3133 out_n.n539 vss 3.80fF $ **FLOATING
C3134 out_n.n540 vss 3.87fF $ **FLOATING
C3135 out_n.n541 vss 4.05fF $ **FLOATING
C3136 out_n.n542 vss 4.05fF $ **FLOATING
C3137 out_n.n543 vss 4.05fF $ **FLOATING
C3138 out_n.n544 vss 4.15fF $ **FLOATING
C3139 out_n.n545 vss 4.15fF $ **FLOATING
C3140 out_n.n546 vss 4.05fF $ **FLOATING
C3141 out_n.n547 vss 4.05fF $ **FLOATING
C3142 out_n.n548 vss 4.05fF $ **FLOATING
C3143 out_n.n549 vss 3.80fF $ **FLOATING
C3144 out_n.n550 vss 3.87fF $ **FLOATING
C3145 out_n.n551 vss 4.05fF $ **FLOATING
C3146 out_n.n552 vss 4.05fF $ **FLOATING
C3147 out_n.n553 vss 4.05fF $ **FLOATING
C3148 out_n.n554 vss 4.15fF $ **FLOATING
C3149 out_n.n555 vss 4.15fF $ **FLOATING
C3150 out_n.n556 vss 4.05fF $ **FLOATING
C3151 out_n.n557 vss 4.05fF $ **FLOATING
C3152 out_n.n558 vss 4.05fF $ **FLOATING
C3153 out_n.n559 vss 3.80fF $ **FLOATING
C3154 out_n.n560 vss 3.87fF $ **FLOATING
C3155 out_n.n561 vss 4.05fF $ **FLOATING
C3156 out_n.n562 vss 4.05fF $ **FLOATING
C3157 out_n.n563 vss 4.05fF $ **FLOATING
C3158 out_n.n564 vss 4.15fF $ **FLOATING
C3159 out_n.n565 vss 4.15fF $ **FLOATING
C3160 out_n.n566 vss 4.05fF $ **FLOATING
C3161 out_n.n567 vss 4.05fF $ **FLOATING
C3162 out_n.n568 vss 4.05fF $ **FLOATING
C3163 out_n.n569 vss 3.80fF $ **FLOATING
C3164 out_n.n570 vss 3.87fF $ **FLOATING
C3165 out_n.n571 vss 4.05fF $ **FLOATING
C3166 out_n.n572 vss 4.05fF $ **FLOATING
C3167 out_n.n573 vss 4.05fF $ **FLOATING
C3168 out_n.n574 vss 4.15fF $ **FLOATING
C3169 out_n.n575 vss 4.15fF $ **FLOATING
C3170 out_n.n576 vss 4.05fF $ **FLOATING
C3171 out_n.n577 vss 4.05fF $ **FLOATING
C3172 out_n.n578 vss 4.05fF $ **FLOATING
C3173 out_n.n579 vss 3.80fF $ **FLOATING
C3174 out_n.n580 vss 3.87fF $ **FLOATING
C3175 out_n.n581 vss 4.05fF $ **FLOATING
C3176 out_n.n582 vss 4.05fF $ **FLOATING
C3177 out_n.n583 vss 4.05fF $ **FLOATING
C3178 out_n.n584 vss 4.15fF $ **FLOATING
C3179 out_n.n585 vss 4.15fF $ **FLOATING
C3180 out_n.n586 vss 4.05fF $ **FLOATING
C3181 out_n.n587 vss 4.05fF $ **FLOATING
C3182 out_n.n588 vss 4.05fF $ **FLOATING
C3183 out_n.n589 vss 3.80fF $ **FLOATING
C3184 out_n.n590 vss 3.87fF $ **FLOATING
C3185 out_n.n591 vss 4.05fF $ **FLOATING
C3186 out_n.n592 vss 4.05fF $ **FLOATING
C3187 out_n.n593 vss 4.05fF $ **FLOATING
C3188 out_n.n594 vss 4.15fF $ **FLOATING
C3189 out_n.n595 vss 4.15fF $ **FLOATING
C3190 out_n.n596 vss 4.05fF $ **FLOATING
C3191 out_n.n597 vss 4.05fF $ **FLOATING
C3192 out_n.n598 vss 4.05fF $ **FLOATING
C3193 out_n.n599 vss 3.80fF $ **FLOATING
C3194 out_n.n600 vss 3.87fF $ **FLOATING
C3195 out_n.n601 vss 4.05fF $ **FLOATING
C3196 out_n.n602 vss 4.05fF $ **FLOATING
C3197 out_n.n603 vss 4.05fF $ **FLOATING
C3198 out_n.n604 vss 4.15fF $ **FLOATING
C3199 out_n.n605 vss 4.15fF $ **FLOATING
C3200 out_n.n606 vss 4.05fF $ **FLOATING
C3201 out_n.n607 vss 4.05fF $ **FLOATING
C3202 out_n.n608 vss 4.05fF $ **FLOATING
C3203 out_n.n609 vss 3.80fF $ **FLOATING
C3204 out_n.n610 vss 3.86fF $ **FLOATING
C3205 out_n.n611 vss 4.05fF $ **FLOATING
C3206 out_n.n612 vss 4.05fF $ **FLOATING
C3207 out_n.n613 vss 4.05fF $ **FLOATING
C3208 out_n.n614 vss 4.15fF $ **FLOATING
C3209 out_n.n615 vss 4.15fF $ **FLOATING
C3210 out_n.n616 vss 4.05fF $ **FLOATING
C3211 out_n.n617 vss 4.05fF $ **FLOATING
C3212 out_n.n618 vss 4.05fF $ **FLOATING
C3213 out_n.n619 vss 3.81fF $ **FLOATING
C3214 out_n.n620 vss 3.85fF $ **FLOATING
C3215 out_n.n621 vss 3.81fF $ **FLOATING
C3216 out_n.n622 vss 23.47fF $ **FLOATING
C3217 out_n.n623 vss 3.85fF $ **FLOATING
C3218 out_n.n624 vss 3.81fF $ **FLOATING
C3219 out_n.n625 vss 30.23fF $ **FLOATING
C3220 out_n.n626 vss 3.85fF $ **FLOATING
C3221 out_n.n627 vss 3.81fF $ **FLOATING
C3222 out_n.n628 vss 30.23fF $ **FLOATING
C3223 out_n.n629 vss 3.85fF $ **FLOATING
C3224 out_n.n630 vss 3.81fF $ **FLOATING
C3225 out_n.n631 vss 30.23fF $ **FLOATING
C3226 out_n.n632 vss 3.85fF $ **FLOATING
C3227 out_n.n633 vss 3.81fF $ **FLOATING
C3228 out_n.n634 vss 30.23fF $ **FLOATING
C3229 out_n.n635 vss 3.85fF $ **FLOATING
C3230 out_n.n636 vss 3.81fF $ **FLOATING
C3231 out_n.n637 vss 30.23fF $ **FLOATING
C3232 out_n.n638 vss 3.85fF $ **FLOATING
C3233 out_n.n639 vss 3.81fF $ **FLOATING
C3234 out_n.n640 vss 30.23fF $ **FLOATING
C3235 out_n.n641 vss 3.85fF $ **FLOATING
C3236 out_n.n642 vss 3.81fF $ **FLOATING
C3237 out_n.n643 vss 30.23fF $ **FLOATING
C3238 out_n.n644 vss 3.85fF $ **FLOATING
C3239 out_n.n645 vss 3.81fF $ **FLOATING
C3240 out_n.n646 vss 30.23fF $ **FLOATING
C3241 out_n.n647 vss 3.85fF $ **FLOATING
C3242 out_n.n648 vss 3.81fF $ **FLOATING
C3243 out_n.n649 vss 30.23fF $ **FLOATING
C3244 out_n.n650 vss 3.85fF $ **FLOATING
C3245 out_n.n651 vss 3.81fF $ **FLOATING
C3246 out_n.n652 vss 30.23fF $ **FLOATING
C3247 out_n.n653 vss 3.85fF $ **FLOATING
C3248 out_n.n654 vss 3.81fF $ **FLOATING
C3249 out_n.n655 vss 30.23fF $ **FLOATING
C3250 out_n.n656 vss 3.85fF $ **FLOATING
C3251 out_n.n657 vss 3.81fF $ **FLOATING
C3252 out_n.n658 vss 30.23fF $ **FLOATING
C3253 out_n.n659 vss 3.85fF $ **FLOATING
C3254 out_n.n660 vss 3.81fF $ **FLOATING
C3255 out_n.n661 vss 30.23fF $ **FLOATING
C3256 out_n.n662 vss 3.85fF $ **FLOATING
C3257 out_n.n663 vss 3.81fF $ **FLOATING
C3258 out_n.n664 vss 30.23fF $ **FLOATING
C3259 out_n.n665 vss 3.85fF $ **FLOATING
C3260 out_n.n666 vss 3.81fF $ **FLOATING
C3261 out_n.n667 vss 30.23fF $ **FLOATING
C3262 out_n.n668 vss 3.85fF $ **FLOATING
C3263 out_n.n669 vss 3.81fF $ **FLOATING
C3264 out_n.n670 vss 30.23fF $ **FLOATING
C3265 out_n.n671 vss 3.85fF $ **FLOATING
C3266 out_n.n672 vss 3.81fF $ **FLOATING
C3267 out_n.n673 vss 30.23fF $ **FLOATING
C3268 out_n.n674 vss 3.85fF $ **FLOATING
C3269 out_n.n675 vss 3.81fF $ **FLOATING
C3270 out_n.n676 vss 30.23fF $ **FLOATING
C3271 out_n.n677 vss 3.85fF $ **FLOATING
C3272 out_n.n678 vss 3.81fF $ **FLOATING
C3273 out_n.n679 vss 30.23fF $ **FLOATING
C3274 out_n.n680 vss 3.85fF $ **FLOATING
C3275 out_n.n681 vss 3.81fF $ **FLOATING
C3276 out_n.n682 vss 30.23fF $ **FLOATING
C3277 out_n.n683 vss 3.85fF $ **FLOATING
C3278 out_n.n684 vss 3.81fF $ **FLOATING
C3279 out_n.n685 vss 30.23fF $ **FLOATING
C3280 out_n.n686 vss 3.85fF $ **FLOATING
C3281 out_n.n687 vss 3.81fF $ **FLOATING
C3282 out_n.n688 vss 30.23fF $ **FLOATING
C3283 out_n.n689 vss 3.85fF $ **FLOATING
C3284 out_n.n690 vss 3.81fF $ **FLOATING
C3285 out_n.n691 vss 30.23fF $ **FLOATING
C3286 out_n.n692 vss 3.85fF $ **FLOATING
C3287 out_n.n693 vss 3.81fF $ **FLOATING
C3288 out_n.n694 vss 30.23fF $ **FLOATING
C3289 out_n.n695 vss 3.85fF $ **FLOATING
C3290 out_n.n696 vss 3.81fF $ **FLOATING
C3291 out_n.n697 vss 30.23fF $ **FLOATING
C3292 out_n.n698 vss 3.85fF $ **FLOATING
C3293 out_n.n699 vss 3.81fF $ **FLOATING
C3294 out_n.n700 vss 30.23fF $ **FLOATING
C3295 out_n.n701 vss 3.85fF $ **FLOATING
C3296 out_n.n702 vss 3.81fF $ **FLOATING
C3297 out_n.n703 vss 30.23fF $ **FLOATING
C3298 out_n.n704 vss 3.85fF $ **FLOATING
C3299 out_n.n705 vss 3.81fF $ **FLOATING
C3300 out_n.n706 vss 30.23fF $ **FLOATING
C3301 out_n.n707 vss 3.85fF $ **FLOATING
C3302 out_n.n708 vss 3.81fF $ **FLOATING
C3303 out_n.n709 vss 30.23fF $ **FLOATING
C3304 out_n.n710 vss 3.85fF $ **FLOATING
C3305 out_n.n711 vss 3.81fF $ **FLOATING
C3306 out_n.n712 vss 30.23fF $ **FLOATING
C3307 out_n.n713 vss 3.85fF $ **FLOATING
C3308 out_n.n714 vss 3.81fF $ **FLOATING
C3309 out_n.n715 vss 30.23fF $ **FLOATING
C3310 out_n.n716 vss 3.85fF $ **FLOATING
C3311 out_n.n717 vss 3.81fF $ **FLOATING
C3312 out_n.n718 vss 30.23fF $ **FLOATING
C3313 out_n.n719 vss 3.85fF $ **FLOATING
C3314 out_n.n720 vss 3.81fF $ **FLOATING
C3315 out_n.n721 vss 30.23fF $ **FLOATING
C3316 out_n.n722 vss 3.85fF $ **FLOATING
C3317 out_n.n723 vss 3.81fF $ **FLOATING
C3318 out_n.n724 vss 30.23fF $ **FLOATING
C3319 out_n.n725 vss 3.85fF $ **FLOATING
C3320 out_n.n726 vss 3.81fF $ **FLOATING
C3321 out_n.n727 vss 30.23fF $ **FLOATING
C3322 out_n.n728 vss 3.85fF $ **FLOATING
C3323 out_n.n729 vss 3.81fF $ **FLOATING
C3324 out_n.n730 vss 30.23fF $ **FLOATING
C3325 out_n.n731 vss 3.85fF $ **FLOATING
C3326 out_n.n732 vss 3.81fF $ **FLOATING
C3327 out_n.n733 vss 30.23fF $ **FLOATING
C3328 out_n.n734 vss 3.85fF $ **FLOATING
C3329 out_n.n735 vss 3.81fF $ **FLOATING
C3330 out_n.n736 vss 30.23fF $ **FLOATING
C3331 out_n.n737 vss 3.85fF $ **FLOATING
C3332 out_n.n738 vss 3.81fF $ **FLOATING
C3333 out_n.n739 vss 30.23fF $ **FLOATING
C3334 out_n.n740 vss 3.85fF $ **FLOATING
C3335 out_n.n741 vss 3.81fF $ **FLOATING
C3336 out_n.n742 vss 30.23fF $ **FLOATING
C3337 out_n.n743 vss 3.85fF $ **FLOATING
C3338 out_n.n744 vss 3.81fF $ **FLOATING
C3339 out_n.n745 vss 30.23fF $ **FLOATING
C3340 out_n.n746 vss 3.85fF $ **FLOATING
C3341 out_n.n747 vss 3.81fF $ **FLOATING
C3342 out_n.n748 vss 30.23fF $ **FLOATING
C3343 out_n.n749 vss 3.85fF $ **FLOATING
C3344 out_n.n750 vss 3.81fF $ **FLOATING
C3345 out_n.n751 vss 30.23fF $ **FLOATING
C3346 out_n.n752 vss 3.85fF $ **FLOATING
C3347 out_n.n753 vss 3.81fF $ **FLOATING
C3348 out_n.n754 vss 30.23fF $ **FLOATING
C3349 out_n.n755 vss 3.85fF $ **FLOATING
C3350 out_n.n756 vss 3.81fF $ **FLOATING
C3351 out_n.n757 vss 30.23fF $ **FLOATING
C3352 out_n.n758 vss 3.85fF $ **FLOATING
C3353 out_n.n759 vss 3.81fF $ **FLOATING
C3354 out_n.n760 vss 30.23fF $ **FLOATING
C3355 out_n.n761 vss 3.85fF $ **FLOATING
C3356 out_n.n762 vss 3.81fF $ **FLOATING
C3357 out_n.n763 vss 30.23fF $ **FLOATING
C3358 out_n.n764 vss 3.85fF $ **FLOATING
C3359 out_n.n765 vss 3.81fF $ **FLOATING
C3360 out_n.n766 vss 30.23fF $ **FLOATING
C3361 out_n.n767 vss 3.85fF $ **FLOATING
C3362 out_n.n768 vss 3.81fF $ **FLOATING
C3363 out_n.n769 vss 30.23fF $ **FLOATING
C3364 out_n.n770 vss 3.85fF $ **FLOATING
C3365 out_n.n771 vss 3.81fF $ **FLOATING
C3366 out_n.n772 vss 30.23fF $ **FLOATING
C3367 out_n.n773 vss 3.85fF $ **FLOATING
C3368 out_n.n774 vss 3.81fF $ **FLOATING
C3369 out_n.n775 vss 30.23fF $ **FLOATING
C3370 out_n.n776 vss 3.85fF $ **FLOATING
C3371 out_n.n777 vss 3.81fF $ **FLOATING
C3372 out_n.n778 vss 30.23fF $ **FLOATING
C3373 out_n.n779 vss 3.85fF $ **FLOATING
C3374 out_n.n780 vss 3.81fF $ **FLOATING
C3375 out_n.n781 vss 30.23fF $ **FLOATING
C3376 out_n.n782 vss 3.85fF $ **FLOATING
C3377 out_n.n783 vss 3.81fF $ **FLOATING
C3378 out_n.n784 vss 30.23fF $ **FLOATING
C3379 out_n.n785 vss 3.85fF $ **FLOATING
C3380 out_n.n786 vss 3.81fF $ **FLOATING
C3381 out_n.n787 vss 30.23fF $ **FLOATING
C3382 out_n.n788 vss 3.85fF $ **FLOATING
C3383 out_n.n789 vss 3.81fF $ **FLOATING
C3384 out_n.n790 vss 30.23fF $ **FLOATING
C3385 out_n.n791 vss 3.85fF $ **FLOATING
C3386 out_n.n792 vss 3.81fF $ **FLOATING
C3387 out_n.n793 vss 30.23fF $ **FLOATING
C3388 out_n.n794 vss 3.85fF $ **FLOATING
C3389 out_n.n795 vss 3.81fF $ **FLOATING
C3390 out_n.n796 vss 30.23fF $ **FLOATING
C3391 out_n.n797 vss 3.85fF $ **FLOATING
C3392 out_n.n798 vss 3.81fF $ **FLOATING
C3393 out_n.n799 vss 30.23fF $ **FLOATING
C3394 out_n.n800 vss 3.85fF $ **FLOATING
C3395 out_n.n801 vss 3.81fF $ **FLOATING
C3396 out_n.n802 vss 29.51fF $ **FLOATING
C3397 out_n.n803 vss 3.85fF $ **FLOATING
C3398 out_n.n804 vss 3.81fF $ **FLOATING
C3399 out_n.n805 vss 3.87fF $ **FLOATING
C3400 out_n.n806 vss 4.05fF $ **FLOATING
C3401 out_n.n807 vss 4.05fF $ **FLOATING
C3402 out_n.n808 vss 4.05fF $ **FLOATING
C3403 out_n.n809 vss 4.15fF $ **FLOATING
C3404 out_n.n810 vss 4.15fF $ **FLOATING
C3405 out_n.n811 vss 4.05fF $ **FLOATING
C3406 out_n.n812 vss 4.05fF $ **FLOATING
C3407 out_n.n813 vss 4.05fF $ **FLOATING
C3408 out_n.n814 vss 3.80fF $ **FLOATING
C3409 out_n.n815 vss 3.87fF $ **FLOATING
C3410 out_n.n816 vss 4.05fF $ **FLOATING
C3411 out_n.n817 vss 4.05fF $ **FLOATING
C3412 out_n.n818 vss 4.05fF $ **FLOATING
C3413 out_n.n819 vss 4.15fF $ **FLOATING
C3414 out_n.n820 vss 4.15fF $ **FLOATING
C3415 out_n.n821 vss 4.05fF $ **FLOATING
C3416 out_n.n822 vss 4.05fF $ **FLOATING
C3417 out_n.n823 vss 4.05fF $ **FLOATING
C3418 out_n.n824 vss 3.80fF $ **FLOATING
C3419 out_n.n825 vss 3.85fF $ **FLOATING
C3420 out_n.n826 vss 3.81fF $ **FLOATING
C3421 out_n.n827 vss 3.87fF $ **FLOATING
C3422 out_n.n828 vss 4.05fF $ **FLOATING
C3423 out_n.n829 vss 4.05fF $ **FLOATING
C3424 out_n.n830 vss 4.05fF $ **FLOATING
C3425 out_n.n831 vss 4.15fF $ **FLOATING
C3426 out_n.n832 vss 4.15fF $ **FLOATING
C3427 out_n.n833 vss 4.05fF $ **FLOATING
C3428 out_n.n834 vss 4.05fF $ **FLOATING
C3429 out_n.n835 vss 4.05fF $ **FLOATING
C3430 out_n.n836 vss 3.80fF $ **FLOATING
C3431 out_n.n837 vss 3.85fF $ **FLOATING
C3432 out_n.n838 vss 3.81fF $ **FLOATING
C3433 out_n.n839 vss 3.87fF $ **FLOATING
C3434 out_n.n840 vss 4.05fF $ **FLOATING
C3435 out_n.n841 vss 4.05fF $ **FLOATING
C3436 out_n.n842 vss 4.05fF $ **FLOATING
C3437 out_n.n843 vss 4.15fF $ **FLOATING
C3438 out_n.n844 vss 4.15fF $ **FLOATING
C3439 out_n.n845 vss 4.05fF $ **FLOATING
C3440 out_n.n846 vss 4.05fF $ **FLOATING
C3441 out_n.n847 vss 4.05fF $ **FLOATING
C3442 out_n.n848 vss 3.80fF $ **FLOATING
C3443 out_n.n849 vss 3.85fF $ **FLOATING
C3444 out_n.n850 vss 3.81fF $ **FLOATING
C3445 out_n.n851 vss 3.87fF $ **FLOATING
C3446 out_n.n852 vss 4.05fF $ **FLOATING
C3447 out_n.n853 vss 4.05fF $ **FLOATING
C3448 out_n.n854 vss 4.05fF $ **FLOATING
C3449 out_n.n855 vss 4.15fF $ **FLOATING
C3450 out_n.n856 vss 4.15fF $ **FLOATING
C3451 out_n.n857 vss 4.05fF $ **FLOATING
C3452 out_n.n858 vss 4.05fF $ **FLOATING
C3453 out_n.n859 vss 4.05fF $ **FLOATING
C3454 out_n.n860 vss 3.80fF $ **FLOATING
C3455 out_n.n861 vss 3.85fF $ **FLOATING
C3456 out_n.n862 vss 3.81fF $ **FLOATING
C3457 out_n.n863 vss 3.87fF $ **FLOATING
C3458 out_n.n864 vss 4.05fF $ **FLOATING
C3459 out_n.n865 vss 4.05fF $ **FLOATING
C3460 out_n.n866 vss 4.05fF $ **FLOATING
C3461 out_n.n867 vss 4.15fF $ **FLOATING
C3462 out_n.n868 vss 4.15fF $ **FLOATING
C3463 out_n.n869 vss 4.05fF $ **FLOATING
C3464 out_n.n870 vss 4.05fF $ **FLOATING
C3465 out_n.n871 vss 4.05fF $ **FLOATING
C3466 out_n.n872 vss 3.80fF $ **FLOATING
C3467 out_n.n873 vss 3.85fF $ **FLOATING
C3468 out_n.n874 vss 3.81fF $ **FLOATING
C3469 out_n.n875 vss 3.87fF $ **FLOATING
C3470 out_n.n876 vss 4.05fF $ **FLOATING
C3471 out_n.n877 vss 4.05fF $ **FLOATING
C3472 out_n.n878 vss 4.05fF $ **FLOATING
C3473 out_n.n879 vss 4.15fF $ **FLOATING
C3474 out_n.n880 vss 4.15fF $ **FLOATING
C3475 out_n.n881 vss 4.05fF $ **FLOATING
C3476 out_n.n882 vss 4.05fF $ **FLOATING
C3477 out_n.n883 vss 4.05fF $ **FLOATING
C3478 out_n.n884 vss 3.80fF $ **FLOATING
C3479 out_n.n885 vss 3.85fF $ **FLOATING
C3480 out_n.n886 vss 3.81fF $ **FLOATING
C3481 out_n.n887 vss 3.87fF $ **FLOATING
C3482 out_n.n888 vss 4.05fF $ **FLOATING
C3483 out_n.n889 vss 4.05fF $ **FLOATING
C3484 out_n.n890 vss 4.05fF $ **FLOATING
C3485 out_n.n891 vss 4.15fF $ **FLOATING
C3486 out_n.n892 vss 4.15fF $ **FLOATING
C3487 out_n.n893 vss 4.05fF $ **FLOATING
C3488 out_n.n894 vss 4.05fF $ **FLOATING
C3489 out_n.n895 vss 4.05fF $ **FLOATING
C3490 out_n.n896 vss 3.80fF $ **FLOATING
C3491 out_n.n897 vss 3.85fF $ **FLOATING
C3492 out_n.n898 vss 3.81fF $ **FLOATING
C3493 out_n.n899 vss 3.87fF $ **FLOATING
C3494 out_n.n900 vss 4.05fF $ **FLOATING
C3495 out_n.n901 vss 4.05fF $ **FLOATING
C3496 out_n.n902 vss 4.05fF $ **FLOATING
C3497 out_n.n903 vss 4.15fF $ **FLOATING
C3498 out_n.n904 vss 4.15fF $ **FLOATING
C3499 out_n.n905 vss 4.05fF $ **FLOATING
C3500 out_n.n906 vss 4.05fF $ **FLOATING
C3501 out_n.n907 vss 4.05fF $ **FLOATING
C3502 out_n.n908 vss 3.80fF $ **FLOATING
C3503 out_n.n909 vss 3.85fF $ **FLOATING
C3504 out_n.n910 vss 3.81fF $ **FLOATING
C3505 out_n.n911 vss 3.87fF $ **FLOATING
C3506 out_n.n912 vss 4.05fF $ **FLOATING
C3507 out_n.n913 vss 4.05fF $ **FLOATING
C3508 out_n.n914 vss 4.05fF $ **FLOATING
C3509 out_n.n915 vss 4.15fF $ **FLOATING
C3510 out_n.n916 vss 4.15fF $ **FLOATING
C3511 out_n.n917 vss 4.05fF $ **FLOATING
C3512 out_n.n918 vss 4.05fF $ **FLOATING
C3513 out_n.n919 vss 4.05fF $ **FLOATING
C3514 out_n.n920 vss 3.80fF $ **FLOATING
C3515 out_n.n921 vss 3.85fF $ **FLOATING
C3516 out_n.n922 vss 3.81fF $ **FLOATING
C3517 out_n.n923 vss 3.87fF $ **FLOATING
C3518 out_n.n924 vss 4.05fF $ **FLOATING
C3519 out_n.n925 vss 4.05fF $ **FLOATING
C3520 out_n.n926 vss 4.05fF $ **FLOATING
C3521 out_n.n927 vss 4.15fF $ **FLOATING
C3522 out_n.n928 vss 4.15fF $ **FLOATING
C3523 out_n.n929 vss 4.05fF $ **FLOATING
C3524 out_n.n930 vss 4.05fF $ **FLOATING
C3525 out_n.n931 vss 4.05fF $ **FLOATING
C3526 out_n.n932 vss 3.80fF $ **FLOATING
C3527 out_n.n933 vss 3.85fF $ **FLOATING
C3528 out_n.n934 vss 3.81fF $ **FLOATING
C3529 out_n.n935 vss 3.87fF $ **FLOATING
C3530 out_n.n936 vss 4.05fF $ **FLOATING
C3531 out_n.n937 vss 4.05fF $ **FLOATING
C3532 out_n.n938 vss 4.05fF $ **FLOATING
C3533 out_n.n939 vss 4.15fF $ **FLOATING
C3534 out_n.n940 vss 4.15fF $ **FLOATING
C3535 out_n.n941 vss 4.05fF $ **FLOATING
C3536 out_n.n942 vss 4.05fF $ **FLOATING
C3537 out_n.n943 vss 4.05fF $ **FLOATING
C3538 out_n.n944 vss 3.80fF $ **FLOATING
C3539 out_n.n945 vss 3.85fF $ **FLOATING
C3540 out_n.n946 vss 3.81fF $ **FLOATING
C3541 out_n.n947 vss 3.87fF $ **FLOATING
C3542 out_n.n948 vss 4.05fF $ **FLOATING
C3543 out_n.n949 vss 4.05fF $ **FLOATING
C3544 out_n.n950 vss 4.05fF $ **FLOATING
C3545 out_n.n951 vss 4.15fF $ **FLOATING
C3546 out_n.n952 vss 4.15fF $ **FLOATING
C3547 out_n.n953 vss 4.05fF $ **FLOATING
C3548 out_n.n954 vss 4.05fF $ **FLOATING
C3549 out_n.n955 vss 4.05fF $ **FLOATING
C3550 out_n.n956 vss 3.80fF $ **FLOATING
C3551 out_n.n957 vss 3.85fF $ **FLOATING
C3552 out_n.n958 vss 3.81fF $ **FLOATING
C3553 out_n.n959 vss 33.39fF $ **FLOATING
C3554 out_n.n960 vss 30.23fF $ **FLOATING
C3555 out_n.n961 vss 30.23fF $ **FLOATING
C3556 out_n.n962 vss 30.23fF $ **FLOATING
C3557 out_n.n963 vss 30.23fF $ **FLOATING
C3558 out_n.n964 vss 30.23fF $ **FLOATING
C3559 out_n.n965 vss 30.23fF $ **FLOATING
C3560 out_n.n966 vss 30.23fF $ **FLOATING
C3561 out_n.n967 vss 30.23fF $ **FLOATING
C3562 out_n.n968 vss 30.23fF $ **FLOATING
C3563 out_n.n969 vss 30.23fF $ **FLOATING
C3564 out_n.n970 vss 28.77fF $ **FLOATING
C3565 out_n.n971 vss 3.85fF $ **FLOATING
C3566 out_n.n972 vss 3.81fF $ **FLOATING
C3567 out_n.n973 vss 30.94fF $ **FLOATING
C3568 vdd2.n0 vss 4.18fF $ **FLOATING
C3569 vdd2.n1 vss 4.39fF $ **FLOATING
C3570 vdd2.n2 vss 4.39fF $ **FLOATING
C3571 vdd2.n3 vss 4.39fF $ **FLOATING
C3572 vdd2.n4 vss 4.50fF $ **FLOATING
C3573 vdd2.n5 vss 4.50fF $ **FLOATING
C3574 vdd2.n6 vss 4.39fF $ **FLOATING
C3575 vdd2.n7 vss 4.39fF $ **FLOATING
C3576 vdd2.n8 vss 4.39fF $ **FLOATING
C3577 vdd2.n9 vss 4.00fF $ **FLOATING
C3578 vdd2.n12 vss 4.18fF $ **FLOATING
C3579 vdd2.n13 vss 4.39fF $ **FLOATING
C3580 vdd2.n14 vss 4.39fF $ **FLOATING
C3581 vdd2.n15 vss 4.39fF $ **FLOATING
C3582 vdd2.n16 vss 4.50fF $ **FLOATING
C3583 vdd2.n17 vss 4.50fF $ **FLOATING
C3584 vdd2.n18 vss 4.39fF $ **FLOATING
C3585 vdd2.n19 vss 4.39fF $ **FLOATING
C3586 vdd2.n20 vss 4.39fF $ **FLOATING
C3587 vdd2.n21 vss 4.00fF $ **FLOATING
C3588 vdd2.n23 vss 5.63fF $ **FLOATING
C3589 vdd2.n24 vss 3.02fF $ **FLOATING
C3590 vdd2.n25 vss 3.02fF $ **FLOATING
C3591 vdd2.n26 vss 3.06fF $ **FLOATING
C3592 vdd2.n27 vss 3.12fF $ **FLOATING
C3593 vdd2.n28 vss 3.02fF $ **FLOATING
C3594 vdd2.n29 vss 3.02fF $ **FLOATING
C3595 vdd2.n30 vss 3.02fF $ **FLOATING
C3596 vdd2.n31 vss 2.58fF $ **FLOATING
C3597 vdd2.n32 vss 4.18fF $ **FLOATING
C3598 vdd2.n33 vss 4.39fF $ **FLOATING
C3599 vdd2.n34 vss 4.39fF $ **FLOATING
C3600 vdd2.n35 vss 4.39fF $ **FLOATING
C3601 vdd2.n36 vss 4.50fF $ **FLOATING
C3602 vdd2.n37 vss 4.50fF $ **FLOATING
C3603 vdd2.n38 vss 4.39fF $ **FLOATING
C3604 vdd2.n39 vss 4.39fF $ **FLOATING
C3605 vdd2.n40 vss 4.39fF $ **FLOATING
C3606 vdd2.n41 vss 4.00fF $ **FLOATING
C3607 vdd2.n42 vss 15.93fF $ **FLOATING
C3608 vdd2.n43 vss 4.18fF $ **FLOATING
C3609 vdd2.n44 vss 4.39fF $ **FLOATING
C3610 vdd2.n45 vss 4.39fF $ **FLOATING
C3611 vdd2.n46 vss 4.39fF $ **FLOATING
C3612 vdd2.n47 vss 4.50fF $ **FLOATING
C3613 vdd2.n48 vss 4.50fF $ **FLOATING
C3614 vdd2.n49 vss 4.39fF $ **FLOATING
C3615 vdd2.n50 vss 4.39fF $ **FLOATING
C3616 vdd2.n51 vss 4.39fF $ **FLOATING
C3617 vdd2.n52 vss 4.00fF $ **FLOATING
C3618 vdd2.n53 vss 33.85fF $ **FLOATING
C3619 vdd2.n54 vss 4.18fF $ **FLOATING
C3620 vdd2.n55 vss 4.39fF $ **FLOATING
C3621 vdd2.n56 vss 4.39fF $ **FLOATING
C3622 vdd2.n57 vss 4.39fF $ **FLOATING
C3623 vdd2.n58 vss 4.50fF $ **FLOATING
C3624 vdd2.n59 vss 4.50fF $ **FLOATING
C3625 vdd2.n60 vss 4.39fF $ **FLOATING
C3626 vdd2.n61 vss 4.39fF $ **FLOATING
C3627 vdd2.n62 vss 4.39fF $ **FLOATING
C3628 vdd2.n63 vss 4.00fF $ **FLOATING
C3629 vdd2.n64 vss 35.61fF $ **FLOATING
C3630 vdd2.n65 vss 4.18fF $ **FLOATING
C3631 vdd2.n66 vss 4.39fF $ **FLOATING
C3632 vdd2.n67 vss 4.39fF $ **FLOATING
C3633 vdd2.n68 vss 4.39fF $ **FLOATING
C3634 vdd2.n69 vss 4.50fF $ **FLOATING
C3635 vdd2.n70 vss 4.50fF $ **FLOATING
C3636 vdd2.n71 vss 4.39fF $ **FLOATING
C3637 vdd2.n72 vss 4.39fF $ **FLOATING
C3638 vdd2.n73 vss 4.39fF $ **FLOATING
C3639 vdd2.n74 vss 4.00fF $ **FLOATING
C3640 vdd2.n75 vss 35.61fF $ **FLOATING
C3641 vdd2.n76 vss 4.18fF $ **FLOATING
C3642 vdd2.n77 vss 4.39fF $ **FLOATING
C3643 vdd2.n78 vss 4.39fF $ **FLOATING
C3644 vdd2.n79 vss 4.39fF $ **FLOATING
C3645 vdd2.n80 vss 4.50fF $ **FLOATING
C3646 vdd2.n81 vss 4.50fF $ **FLOATING
C3647 vdd2.n82 vss 4.39fF $ **FLOATING
C3648 vdd2.n83 vss 4.39fF $ **FLOATING
C3649 vdd2.n84 vss 4.39fF $ **FLOATING
C3650 vdd2.n85 vss 4.00fF $ **FLOATING
C3651 vdd2.n86 vss 35.61fF $ **FLOATING
C3652 vdd2.n87 vss 4.18fF $ **FLOATING
C3653 vdd2.n88 vss 4.39fF $ **FLOATING
C3654 vdd2.n89 vss 4.39fF $ **FLOATING
C3655 vdd2.n90 vss 4.39fF $ **FLOATING
C3656 vdd2.n91 vss 4.50fF $ **FLOATING
C3657 vdd2.n92 vss 4.50fF $ **FLOATING
C3658 vdd2.n93 vss 4.39fF $ **FLOATING
C3659 vdd2.n94 vss 4.39fF $ **FLOATING
C3660 vdd2.n95 vss 4.39fF $ **FLOATING
C3661 vdd2.n96 vss 4.00fF $ **FLOATING
C3662 vdd2.n97 vss 35.61fF $ **FLOATING
C3663 vdd2.n98 vss 4.18fF $ **FLOATING
C3664 vdd2.n99 vss 4.39fF $ **FLOATING
C3665 vdd2.n100 vss 4.39fF $ **FLOATING
C3666 vdd2.n101 vss 4.39fF $ **FLOATING
C3667 vdd2.n102 vss 4.50fF $ **FLOATING
C3668 vdd2.n103 vss 4.50fF $ **FLOATING
C3669 vdd2.n104 vss 4.39fF $ **FLOATING
C3670 vdd2.n105 vss 4.39fF $ **FLOATING
C3671 vdd2.n106 vss 4.39fF $ **FLOATING
C3672 vdd2.n107 vss 4.00fF $ **FLOATING
C3673 vdd2.n108 vss 35.61fF $ **FLOATING
C3674 vdd2.n109 vss 4.18fF $ **FLOATING
C3675 vdd2.n110 vss 4.39fF $ **FLOATING
C3676 vdd2.n111 vss 4.39fF $ **FLOATING
C3677 vdd2.n112 vss 4.39fF $ **FLOATING
C3678 vdd2.n113 vss 4.50fF $ **FLOATING
C3679 vdd2.n114 vss 4.50fF $ **FLOATING
C3680 vdd2.n115 vss 4.39fF $ **FLOATING
C3681 vdd2.n116 vss 4.39fF $ **FLOATING
C3682 vdd2.n117 vss 4.39fF $ **FLOATING
C3683 vdd2.n118 vss 4.00fF $ **FLOATING
C3684 vdd2.n119 vss 35.61fF $ **FLOATING
C3685 vdd2.n120 vss 4.18fF $ **FLOATING
C3686 vdd2.n121 vss 4.39fF $ **FLOATING
C3687 vdd2.n122 vss 4.39fF $ **FLOATING
C3688 vdd2.n123 vss 4.39fF $ **FLOATING
C3689 vdd2.n124 vss 4.50fF $ **FLOATING
C3690 vdd2.n125 vss 4.50fF $ **FLOATING
C3691 vdd2.n126 vss 4.39fF $ **FLOATING
C3692 vdd2.n127 vss 4.39fF $ **FLOATING
C3693 vdd2.n128 vss 4.39fF $ **FLOATING
C3694 vdd2.n129 vss 4.00fF $ **FLOATING
C3695 vdd2.n130 vss 35.61fF $ **FLOATING
C3696 vdd2.n131 vss 4.18fF $ **FLOATING
C3697 vdd2.n132 vss 4.39fF $ **FLOATING
C3698 vdd2.n133 vss 4.39fF $ **FLOATING
C3699 vdd2.n134 vss 4.39fF $ **FLOATING
C3700 vdd2.n135 vss 4.50fF $ **FLOATING
C3701 vdd2.n136 vss 4.50fF $ **FLOATING
C3702 vdd2.n137 vss 4.39fF $ **FLOATING
C3703 vdd2.n138 vss 4.39fF $ **FLOATING
C3704 vdd2.n139 vss 4.39fF $ **FLOATING
C3705 vdd2.n140 vss 4.00fF $ **FLOATING
C3706 vdd2.n141 vss 35.61fF $ **FLOATING
C3707 vdd2.n142 vss 4.18fF $ **FLOATING
C3708 vdd2.n143 vss 4.39fF $ **FLOATING
C3709 vdd2.n144 vss 4.39fF $ **FLOATING
C3710 vdd2.n145 vss 4.39fF $ **FLOATING
C3711 vdd2.n146 vss 4.50fF $ **FLOATING
C3712 vdd2.n147 vss 4.50fF $ **FLOATING
C3713 vdd2.n148 vss 4.39fF $ **FLOATING
C3714 vdd2.n149 vss 4.39fF $ **FLOATING
C3715 vdd2.n150 vss 4.39fF $ **FLOATING
C3716 vdd2.n151 vss 4.00fF $ **FLOATING
C3717 vdd2.n152 vss 35.61fF $ **FLOATING
C3718 vdd2.n153 vss 4.18fF $ **FLOATING
C3719 vdd2.n154 vss 4.39fF $ **FLOATING
C3720 vdd2.n155 vss 4.39fF $ **FLOATING
C3721 vdd2.n156 vss 4.39fF $ **FLOATING
C3722 vdd2.n157 vss 4.50fF $ **FLOATING
C3723 vdd2.n158 vss 4.50fF $ **FLOATING
C3724 vdd2.n159 vss 4.39fF $ **FLOATING
C3725 vdd2.n160 vss 4.39fF $ **FLOATING
C3726 vdd2.n161 vss 4.39fF $ **FLOATING
C3727 vdd2.n162 vss 4.00fF $ **FLOATING
C3728 vdd2.n163 vss 35.61fF $ **FLOATING
C3729 vdd2.n164 vss 4.18fF $ **FLOATING
C3730 vdd2.n165 vss 4.39fF $ **FLOATING
C3731 vdd2.n166 vss 4.39fF $ **FLOATING
C3732 vdd2.n167 vss 4.39fF $ **FLOATING
C3733 vdd2.n168 vss 4.50fF $ **FLOATING
C3734 vdd2.n169 vss 4.50fF $ **FLOATING
C3735 vdd2.n170 vss 4.39fF $ **FLOATING
C3736 vdd2.n171 vss 4.39fF $ **FLOATING
C3737 vdd2.n172 vss 4.39fF $ **FLOATING
C3738 vdd2.n173 vss 4.00fF $ **FLOATING
C3739 vdd2.n174 vss 35.61fF $ **FLOATING
C3740 vdd2.n175 vss 4.18fF $ **FLOATING
C3741 vdd2.n176 vss 4.39fF $ **FLOATING
C3742 vdd2.n177 vss 4.39fF $ **FLOATING
C3743 vdd2.n178 vss 4.39fF $ **FLOATING
C3744 vdd2.n179 vss 4.50fF $ **FLOATING
C3745 vdd2.n180 vss 4.50fF $ **FLOATING
C3746 vdd2.n181 vss 4.39fF $ **FLOATING
C3747 vdd2.n182 vss 4.39fF $ **FLOATING
C3748 vdd2.n183 vss 4.39fF $ **FLOATING
C3749 vdd2.n184 vss 4.00fF $ **FLOATING
C3750 vdd2.n185 vss 35.61fF $ **FLOATING
C3751 vdd2.n186 vss 4.18fF $ **FLOATING
C3752 vdd2.n187 vss 4.39fF $ **FLOATING
C3753 vdd2.n188 vss 4.39fF $ **FLOATING
C3754 vdd2.n189 vss 4.39fF $ **FLOATING
C3755 vdd2.n190 vss 4.50fF $ **FLOATING
C3756 vdd2.n191 vss 4.50fF $ **FLOATING
C3757 vdd2.n192 vss 4.39fF $ **FLOATING
C3758 vdd2.n193 vss 4.39fF $ **FLOATING
C3759 vdd2.n194 vss 4.39fF $ **FLOATING
C3760 vdd2.n195 vss 4.00fF $ **FLOATING
C3761 vdd2.n196 vss 35.61fF $ **FLOATING
C3762 vdd2.n197 vss 4.18fF $ **FLOATING
C3763 vdd2.n198 vss 4.39fF $ **FLOATING
C3764 vdd2.n199 vss 4.39fF $ **FLOATING
C3765 vdd2.n200 vss 4.39fF $ **FLOATING
C3766 vdd2.n201 vss 4.50fF $ **FLOATING
C3767 vdd2.n202 vss 4.50fF $ **FLOATING
C3768 vdd2.n203 vss 4.39fF $ **FLOATING
C3769 vdd2.n204 vss 4.39fF $ **FLOATING
C3770 vdd2.n205 vss 4.39fF $ **FLOATING
C3771 vdd2.n206 vss 4.00fF $ **FLOATING
C3772 vdd2.n207 vss 35.61fF $ **FLOATING
C3773 vdd2.n208 vss 4.18fF $ **FLOATING
C3774 vdd2.n209 vss 4.39fF $ **FLOATING
C3775 vdd2.n210 vss 4.39fF $ **FLOATING
C3776 vdd2.n211 vss 4.39fF $ **FLOATING
C3777 vdd2.n212 vss 4.50fF $ **FLOATING
C3778 vdd2.n213 vss 4.50fF $ **FLOATING
C3779 vdd2.n214 vss 4.39fF $ **FLOATING
C3780 vdd2.n215 vss 4.39fF $ **FLOATING
C3781 vdd2.n216 vss 4.39fF $ **FLOATING
C3782 vdd2.n217 vss 4.00fF $ **FLOATING
C3783 vdd2.n218 vss 35.61fF $ **FLOATING
C3784 vdd2.n219 vss 4.18fF $ **FLOATING
C3785 vdd2.n220 vss 4.39fF $ **FLOATING
C3786 vdd2.n221 vss 4.39fF $ **FLOATING
C3787 vdd2.n222 vss 4.39fF $ **FLOATING
C3788 vdd2.n223 vss 4.50fF $ **FLOATING
C3789 vdd2.n224 vss 4.50fF $ **FLOATING
C3790 vdd2.n225 vss 4.39fF $ **FLOATING
C3791 vdd2.n226 vss 4.39fF $ **FLOATING
C3792 vdd2.n227 vss 4.39fF $ **FLOATING
C3793 vdd2.n228 vss 4.00fF $ **FLOATING
C3794 vdd2.n229 vss 35.61fF $ **FLOATING
C3795 vdd2.n230 vss 4.18fF $ **FLOATING
C3796 vdd2.n231 vss 4.39fF $ **FLOATING
C3797 vdd2.n232 vss 4.39fF $ **FLOATING
C3798 vdd2.n233 vss 4.39fF $ **FLOATING
C3799 vdd2.n234 vss 4.50fF $ **FLOATING
C3800 vdd2.n235 vss 4.50fF $ **FLOATING
C3801 vdd2.n236 vss 4.39fF $ **FLOATING
C3802 vdd2.n237 vss 4.39fF $ **FLOATING
C3803 vdd2.n238 vss 4.39fF $ **FLOATING
C3804 vdd2.n239 vss 4.00fF $ **FLOATING
C3805 vdd2.n240 vss 35.61fF $ **FLOATING
C3806 vdd2.n241 vss 4.18fF $ **FLOATING
C3807 vdd2.n242 vss 4.39fF $ **FLOATING
C3808 vdd2.n243 vss 4.39fF $ **FLOATING
C3809 vdd2.n244 vss 4.39fF $ **FLOATING
C3810 vdd2.n245 vss 4.50fF $ **FLOATING
C3811 vdd2.n246 vss 4.50fF $ **FLOATING
C3812 vdd2.n247 vss 4.39fF $ **FLOATING
C3813 vdd2.n248 vss 4.39fF $ **FLOATING
C3814 vdd2.n249 vss 4.39fF $ **FLOATING
C3815 vdd2.n250 vss 4.00fF $ **FLOATING
C3816 vdd2.n251 vss 35.61fF $ **FLOATING
C3817 vdd2.n252 vss 4.18fF $ **FLOATING
C3818 vdd2.n253 vss 4.39fF $ **FLOATING
C3819 vdd2.n254 vss 4.39fF $ **FLOATING
C3820 vdd2.n255 vss 4.39fF $ **FLOATING
C3821 vdd2.n256 vss 4.50fF $ **FLOATING
C3822 vdd2.n257 vss 4.50fF $ **FLOATING
C3823 vdd2.n258 vss 4.39fF $ **FLOATING
C3824 vdd2.n259 vss 4.39fF $ **FLOATING
C3825 vdd2.n260 vss 4.39fF $ **FLOATING
C3826 vdd2.n261 vss 4.00fF $ **FLOATING
C3827 vdd2.n262 vss 35.61fF $ **FLOATING
C3828 vdd2.n263 vss 4.18fF $ **FLOATING
C3829 vdd2.n264 vss 4.39fF $ **FLOATING
C3830 vdd2.n265 vss 4.39fF $ **FLOATING
C3831 vdd2.n266 vss 4.39fF $ **FLOATING
C3832 vdd2.n267 vss 4.50fF $ **FLOATING
C3833 vdd2.n268 vss 4.50fF $ **FLOATING
C3834 vdd2.n269 vss 4.39fF $ **FLOATING
C3835 vdd2.n270 vss 4.39fF $ **FLOATING
C3836 vdd2.n271 vss 4.39fF $ **FLOATING
C3837 vdd2.n272 vss 4.00fF $ **FLOATING
C3838 vdd2.n273 vss 35.61fF $ **FLOATING
C3839 vdd2.n274 vss 4.18fF $ **FLOATING
C3840 vdd2.n275 vss 4.39fF $ **FLOATING
C3841 vdd2.n276 vss 4.39fF $ **FLOATING
C3842 vdd2.n277 vss 4.39fF $ **FLOATING
C3843 vdd2.n278 vss 4.50fF $ **FLOATING
C3844 vdd2.n279 vss 4.50fF $ **FLOATING
C3845 vdd2.n280 vss 4.39fF $ **FLOATING
C3846 vdd2.n281 vss 4.39fF $ **FLOATING
C3847 vdd2.n282 vss 4.39fF $ **FLOATING
C3848 vdd2.n283 vss 4.00fF $ **FLOATING
C3849 vdd2.n284 vss 35.61fF $ **FLOATING
C3850 vdd2.n285 vss 4.18fF $ **FLOATING
C3851 vdd2.n286 vss 4.39fF $ **FLOATING
C3852 vdd2.n287 vss 4.39fF $ **FLOATING
C3853 vdd2.n288 vss 4.39fF $ **FLOATING
C3854 vdd2.n289 vss 4.50fF $ **FLOATING
C3855 vdd2.n290 vss 4.50fF $ **FLOATING
C3856 vdd2.n291 vss 4.39fF $ **FLOATING
C3857 vdd2.n292 vss 4.39fF $ **FLOATING
C3858 vdd2.n293 vss 4.39fF $ **FLOATING
C3859 vdd2.n294 vss 4.00fF $ **FLOATING
C3860 vdd2.n295 vss 35.61fF $ **FLOATING
C3861 vdd2.n296 vss 4.18fF $ **FLOATING
C3862 vdd2.n297 vss 4.39fF $ **FLOATING
C3863 vdd2.n298 vss 4.39fF $ **FLOATING
C3864 vdd2.n299 vss 4.39fF $ **FLOATING
C3865 vdd2.n300 vss 4.50fF $ **FLOATING
C3866 vdd2.n301 vss 4.50fF $ **FLOATING
C3867 vdd2.n302 vss 4.39fF $ **FLOATING
C3868 vdd2.n303 vss 4.39fF $ **FLOATING
C3869 vdd2.n304 vss 4.39fF $ **FLOATING
C3870 vdd2.n305 vss 4.00fF $ **FLOATING
C3871 vdd2.n306 vss 35.61fF $ **FLOATING
C3872 vdd2.n307 vss 4.18fF $ **FLOATING
C3873 vdd2.n308 vss 4.39fF $ **FLOATING
C3874 vdd2.n309 vss 4.39fF $ **FLOATING
C3875 vdd2.n310 vss 4.39fF $ **FLOATING
C3876 vdd2.n311 vss 4.50fF $ **FLOATING
C3877 vdd2.n312 vss 4.50fF $ **FLOATING
C3878 vdd2.n313 vss 4.39fF $ **FLOATING
C3879 vdd2.n314 vss 4.39fF $ **FLOATING
C3880 vdd2.n315 vss 4.39fF $ **FLOATING
C3881 vdd2.n316 vss 4.00fF $ **FLOATING
C3882 vdd2.n317 vss 35.61fF $ **FLOATING
C3883 vdd2.n318 vss 4.18fF $ **FLOATING
C3884 vdd2.n319 vss 4.39fF $ **FLOATING
C3885 vdd2.n320 vss 4.39fF $ **FLOATING
C3886 vdd2.n321 vss 4.39fF $ **FLOATING
C3887 vdd2.n322 vss 4.50fF $ **FLOATING
C3888 vdd2.n323 vss 4.50fF $ **FLOATING
C3889 vdd2.n324 vss 4.39fF $ **FLOATING
C3890 vdd2.n325 vss 4.39fF $ **FLOATING
C3891 vdd2.n326 vss 4.39fF $ **FLOATING
C3892 vdd2.n327 vss 4.00fF $ **FLOATING
C3893 vdd2.n328 vss 35.61fF $ **FLOATING
C3894 vdd2.n329 vss 4.18fF $ **FLOATING
C3895 vdd2.n330 vss 4.39fF $ **FLOATING
C3896 vdd2.n331 vss 4.39fF $ **FLOATING
C3897 vdd2.n332 vss 4.39fF $ **FLOATING
C3898 vdd2.n333 vss 4.50fF $ **FLOATING
C3899 vdd2.n334 vss 4.50fF $ **FLOATING
C3900 vdd2.n335 vss 4.39fF $ **FLOATING
C3901 vdd2.n336 vss 4.39fF $ **FLOATING
C3902 vdd2.n337 vss 4.39fF $ **FLOATING
C3903 vdd2.n338 vss 4.00fF $ **FLOATING
C3904 vdd2.n339 vss 35.61fF $ **FLOATING
C3905 vdd2.n340 vss 4.18fF $ **FLOATING
C3906 vdd2.n341 vss 4.39fF $ **FLOATING
C3907 vdd2.n342 vss 4.39fF $ **FLOATING
C3908 vdd2.n343 vss 4.39fF $ **FLOATING
C3909 vdd2.n344 vss 4.50fF $ **FLOATING
C3910 vdd2.n345 vss 4.50fF $ **FLOATING
C3911 vdd2.n346 vss 4.39fF $ **FLOATING
C3912 vdd2.n347 vss 4.39fF $ **FLOATING
C3913 vdd2.n348 vss 4.39fF $ **FLOATING
C3914 vdd2.n349 vss 4.00fF $ **FLOATING
C3915 vdd2.n350 vss 35.61fF $ **FLOATING
C3916 vdd2.n351 vss 4.18fF $ **FLOATING
C3917 vdd2.n352 vss 4.39fF $ **FLOATING
C3918 vdd2.n353 vss 4.39fF $ **FLOATING
C3919 vdd2.n354 vss 4.39fF $ **FLOATING
C3920 vdd2.n355 vss 4.50fF $ **FLOATING
C3921 vdd2.n356 vss 4.50fF $ **FLOATING
C3922 vdd2.n357 vss 4.39fF $ **FLOATING
C3923 vdd2.n358 vss 4.39fF $ **FLOATING
C3924 vdd2.n359 vss 4.39fF $ **FLOATING
C3925 vdd2.n360 vss 4.00fF $ **FLOATING
C3926 vdd2.n361 vss 35.61fF $ **FLOATING
C3927 vdd2.n362 vss 4.18fF $ **FLOATING
C3928 vdd2.n363 vss 4.39fF $ **FLOATING
C3929 vdd2.n364 vss 4.39fF $ **FLOATING
C3930 vdd2.n365 vss 4.39fF $ **FLOATING
C3931 vdd2.n366 vss 4.50fF $ **FLOATING
C3932 vdd2.n367 vss 4.50fF $ **FLOATING
C3933 vdd2.n368 vss 4.39fF $ **FLOATING
C3934 vdd2.n369 vss 4.39fF $ **FLOATING
C3935 vdd2.n370 vss 4.39fF $ **FLOATING
C3936 vdd2.n371 vss 4.00fF $ **FLOATING
C3937 vdd2.n372 vss 35.61fF $ **FLOATING
C3938 vdd2.n373 vss 4.18fF $ **FLOATING
C3939 vdd2.n374 vss 4.39fF $ **FLOATING
C3940 vdd2.n375 vss 4.39fF $ **FLOATING
C3941 vdd2.n376 vss 4.39fF $ **FLOATING
C3942 vdd2.n377 vss 4.50fF $ **FLOATING
C3943 vdd2.n378 vss 4.50fF $ **FLOATING
C3944 vdd2.n379 vss 4.39fF $ **FLOATING
C3945 vdd2.n380 vss 4.39fF $ **FLOATING
C3946 vdd2.n381 vss 4.39fF $ **FLOATING
C3947 vdd2.n382 vss 4.00fF $ **FLOATING
C3948 vdd2.n383 vss 35.61fF $ **FLOATING
C3949 vdd2.n384 vss 4.18fF $ **FLOATING
C3950 vdd2.n385 vss 4.39fF $ **FLOATING
C3951 vdd2.n386 vss 4.39fF $ **FLOATING
C3952 vdd2.n387 vss 4.39fF $ **FLOATING
C3953 vdd2.n388 vss 4.50fF $ **FLOATING
C3954 vdd2.n389 vss 4.50fF $ **FLOATING
C3955 vdd2.n390 vss 4.39fF $ **FLOATING
C3956 vdd2.n391 vss 4.39fF $ **FLOATING
C3957 vdd2.n392 vss 4.39fF $ **FLOATING
C3958 vdd2.n393 vss 4.00fF $ **FLOATING
C3959 vdd2.n394 vss 5.44fF $ **FLOATING
C3960 vdd2.n395 vss 34.35fF $ **FLOATING
C3961 vdd2.n396 vss 4.18fF $ **FLOATING
C3962 vdd2.n397 vss 4.39fF $ **FLOATING
C3963 vdd2.n398 vss 4.39fF $ **FLOATING
C3964 vdd2.n399 vss 4.39fF $ **FLOATING
C3965 vdd2.n400 vss 4.50fF $ **FLOATING
C3966 vdd2.n401 vss 4.50fF $ **FLOATING
C3967 vdd2.n402 vss 4.39fF $ **FLOATING
C3968 vdd2.n403 vss 4.39fF $ **FLOATING
C3969 vdd2.n404 vss 4.39fF $ **FLOATING
C3970 vdd2.n405 vss 4.00fF $ **FLOATING
C3971 vdd2.n406 vss 28.86fF $ **FLOATING
C3972 vdd2.n407 vss 4.18fF $ **FLOATING
C3973 vdd2.n408 vss 4.39fF $ **FLOATING
C3974 vdd2.n409 vss 4.39fF $ **FLOATING
C3975 vdd2.n410 vss 4.39fF $ **FLOATING
C3976 vdd2.n411 vss 4.50fF $ **FLOATING
C3977 vdd2.n412 vss 4.50fF $ **FLOATING
C3978 vdd2.n413 vss 4.39fF $ **FLOATING
C3979 vdd2.n414 vss 4.39fF $ **FLOATING
C3980 vdd2.n415 vss 4.39fF $ **FLOATING
C3981 vdd2.n416 vss 4.00fF $ **FLOATING
C3982 vdd2.n417 vss 35.26fF $ **FLOATING
C3983 vdd2.n418 vss 4.18fF $ **FLOATING
C3984 vdd2.n419 vss 4.39fF $ **FLOATING
C3985 vdd2.n420 vss 4.39fF $ **FLOATING
C3986 vdd2.n421 vss 4.39fF $ **FLOATING
C3987 vdd2.n422 vss 4.50fF $ **FLOATING
C3988 vdd2.n423 vss 4.50fF $ **FLOATING
C3989 vdd2.n424 vss 4.39fF $ **FLOATING
C3990 vdd2.n425 vss 4.39fF $ **FLOATING
C3991 vdd2.n426 vss 4.39fF $ **FLOATING
C3992 vdd2.n427 vss 4.00fF $ **FLOATING
C3993 vdd2.n428 vss 5.44fF $ **FLOATING
C3994 vdd2.n429 vss 6.32fF $ **FLOATING
C3995 vdd2.n430 vss 13.70fF $ **FLOATING
C3996 vdd2.n431 vss 5.42fF $ **FLOATING
C3997 vdd2.n432 vss 5.42fF $ **FLOATING
C3998 vdd2.n433 vss 6.32fF $ **FLOATING
C3999 vdd2.n434 vss 11.52fF $ **FLOATING
C4000 vdd2.n435 vss 13.70fF $ **FLOATING
C4001 vdd2.n436 vss 5.40fF $ **FLOATING
C4002 vdd2.n437 vss 5.40fF $ **FLOATING
C4003 vdd2.n438 vss 6.30fF $ **FLOATING
C4004 vdd2.n439 vss 6.30fF $ **FLOATING
C4005 vdd2.n440 vss 11.52fF $ **FLOATING
C4006 vdd2.n441 vss 6.39fF $ **FLOATING
C4007 vdd2.n442 vss 32.35fF $ **FLOATING
C4008 vdd2.n443 vss 34.35fF $ **FLOATING
C4009 vdd2.n444 vss 4.18fF $ **FLOATING
C4010 vdd2.n445 vss 4.39fF $ **FLOATING
C4011 vdd2.n446 vss 4.39fF $ **FLOATING
C4012 vdd2.n447 vss 4.39fF $ **FLOATING
C4013 vdd2.n448 vss 4.50fF $ **FLOATING
C4014 vdd2.n449 vss 4.50fF $ **FLOATING
C4015 vdd2.n450 vss 4.39fF $ **FLOATING
C4016 vdd2.n451 vss 4.39fF $ **FLOATING
C4017 vdd2.n452 vss 4.39fF $ **FLOATING
C4018 vdd2.n453 vss 4.00fF $ **FLOATING
C4019 vdd2.n455 vss 34.60fF $ **FLOATING
C4020 vdd2.n456 vss 4.18fF $ **FLOATING
C4021 vdd2.n457 vss 4.39fF $ **FLOATING
C4022 vdd2.n458 vss 4.39fF $ **FLOATING
C4023 vdd2.n459 vss 4.39fF $ **FLOATING
C4024 vdd2.n460 vss 4.50fF $ **FLOATING
C4025 vdd2.n461 vss 4.50fF $ **FLOATING
C4026 vdd2.n462 vss 4.39fF $ **FLOATING
C4027 vdd2.n463 vss 4.39fF $ **FLOATING
C4028 vdd2.n464 vss 4.39fF $ **FLOATING
C4029 vdd2.n465 vss 4.00fF $ **FLOATING
C4030 vdd2.n466 vss 31.18fF $ **FLOATING
C4031 vdd2.n467 vss 4.18fF $ **FLOATING
C4032 vdd2.n468 vss 4.39fF $ **FLOATING
C4033 vdd2.n469 vss 4.39fF $ **FLOATING
C4034 vdd2.n470 vss 4.39fF $ **FLOATING
C4035 vdd2.n471 vss 4.50fF $ **FLOATING
C4036 vdd2.n472 vss 4.50fF $ **FLOATING
C4037 vdd2.n473 vss 4.39fF $ **FLOATING
C4038 vdd2.n474 vss 4.39fF $ **FLOATING
C4039 vdd2.n475 vss 4.39fF $ **FLOATING
C4040 vdd2.n476 vss 4.00fF $ **FLOATING
C4041 vdd2.n477 vss 35.61fF $ **FLOATING
C4042 vdd2.n478 vss 4.18fF $ **FLOATING
C4043 vdd2.n479 vss 4.39fF $ **FLOATING
C4044 vdd2.n480 vss 4.39fF $ **FLOATING
C4045 vdd2.n481 vss 4.39fF $ **FLOATING
C4046 vdd2.n482 vss 4.50fF $ **FLOATING
C4047 vdd2.n483 vss 4.50fF $ **FLOATING
C4048 vdd2.n484 vss 4.39fF $ **FLOATING
C4049 vdd2.n485 vss 4.39fF $ **FLOATING
C4050 vdd2.n486 vss 4.39fF $ **FLOATING
C4051 vdd2.n487 vss 4.00fF $ **FLOATING
C4052 vdd2.n488 vss 5.44fF $ **FLOATING
C4053 vdd2.n490 vss 34.35fF $ **FLOATING
C4054 vdd2.n491 vss 4.18fF $ **FLOATING
C4055 vdd2.n492 vss 4.39fF $ **FLOATING
C4056 vdd2.n493 vss 4.39fF $ **FLOATING
C4057 vdd2.n494 vss 4.39fF $ **FLOATING
C4058 vdd2.n495 vss 4.50fF $ **FLOATING
C4059 vdd2.n496 vss 4.50fF $ **FLOATING
C4060 vdd2.n497 vss 4.39fF $ **FLOATING
C4061 vdd2.n498 vss 4.39fF $ **FLOATING
C4062 vdd2.n499 vss 4.39fF $ **FLOATING
C4063 vdd2.n500 vss 4.00fF $ **FLOATING
C4064 vdd2.n501 vss 1.00fF $ **FLOATING
C4065 vdd2.n502 vss 3.27fF $ **FLOATING
C4066 vdd2.n503 vss 1.86fF $ **FLOATING
C4067 vdd2.n504 vss 1.86fF $ **FLOATING
C4068 vdd2.n505 vss 1.90fF $ **FLOATING
C4069 vdd2.n506 vss 1.95fF $ **FLOATING
C4070 vdd2.n507 vss 1.91fF $ **FLOATING
C4071 vdd2.n508 vss 1.91fF $ **FLOATING
C4072 vdd2.n509 vss 1.91fF $ **FLOATING
C4073 vdd2.n510 vss 1.78fF $ **FLOATING
C4074 vdd2.n511 vss 4.18fF $ **FLOATING
C4075 vdd2.n512 vss 4.38fF $ **FLOATING
C4076 vdd2.n513 vss 4.38fF $ **FLOATING
C4077 vdd2.n514 vss 4.38fF $ **FLOATING
C4078 vdd2.n515 vss 4.49fF $ **FLOATING
C4079 vdd2.n516 vss 4.49fF $ **FLOATING
C4080 vdd2.n517 vss 4.38fF $ **FLOATING
C4081 vdd2.n518 vss 4.38fF $ **FLOATING
C4082 vdd2.n519 vss 4.38fF $ **FLOATING
C4083 vdd2.n520 vss 3.99fF $ **FLOATING
C4084 vdd2.n521 vss 34.31fF $ **FLOATING
C4085 vdd2.n522 vss 4.18fF $ **FLOATING
C4086 vdd2.n523 vss 4.39fF $ **FLOATING
C4087 vdd2.n524 vss 4.39fF $ **FLOATING
C4088 vdd2.n525 vss 4.39fF $ **FLOATING
C4089 vdd2.n526 vss 4.50fF $ **FLOATING
C4090 vdd2.n527 vss 4.50fF $ **FLOATING
C4091 vdd2.n528 vss 4.39fF $ **FLOATING
C4092 vdd2.n529 vss 4.39fF $ **FLOATING
C4093 vdd2.n530 vss 4.39fF $ **FLOATING
C4094 vdd2.n531 vss 4.00fF $ **FLOATING
C4095 vdd2.n532 vss 35.61fF $ **FLOATING
C4096 vdd2.n533 vss 4.18fF $ **FLOATING
C4097 vdd2.n534 vss 4.39fF $ **FLOATING
C4098 vdd2.n535 vss 4.39fF $ **FLOATING
C4099 vdd2.n536 vss 4.39fF $ **FLOATING
C4100 vdd2.n537 vss 4.50fF $ **FLOATING
C4101 vdd2.n538 vss 4.50fF $ **FLOATING
C4102 vdd2.n539 vss 4.39fF $ **FLOATING
C4103 vdd2.n540 vss 4.39fF $ **FLOATING
C4104 vdd2.n541 vss 4.39fF $ **FLOATING
C4105 vdd2.n542 vss 4.00fF $ **FLOATING
C4106 vdd2.n543 vss 35.61fF $ **FLOATING
C4107 vdd2.n544 vss 4.18fF $ **FLOATING
C4108 vdd2.n545 vss 4.39fF $ **FLOATING
C4109 vdd2.n546 vss 4.39fF $ **FLOATING
C4110 vdd2.n547 vss 4.39fF $ **FLOATING
C4111 vdd2.n548 vss 4.50fF $ **FLOATING
C4112 vdd2.n549 vss 4.50fF $ **FLOATING
C4113 vdd2.n550 vss 4.39fF $ **FLOATING
C4114 vdd2.n551 vss 4.39fF $ **FLOATING
C4115 vdd2.n552 vss 4.39fF $ **FLOATING
C4116 vdd2.n553 vss 4.00fF $ **FLOATING
C4117 vdd2.n554 vss 35.61fF $ **FLOATING
C4118 vdd2.n555 vss 4.18fF $ **FLOATING
C4119 vdd2.n556 vss 4.39fF $ **FLOATING
C4120 vdd2.n557 vss 4.39fF $ **FLOATING
C4121 vdd2.n558 vss 4.39fF $ **FLOATING
C4122 vdd2.n559 vss 4.50fF $ **FLOATING
C4123 vdd2.n560 vss 4.50fF $ **FLOATING
C4124 vdd2.n561 vss 4.39fF $ **FLOATING
C4125 vdd2.n562 vss 4.39fF $ **FLOATING
C4126 vdd2.n563 vss 4.39fF $ **FLOATING
C4127 vdd2.n564 vss 4.00fF $ **FLOATING
C4128 vdd2.n565 vss 35.61fF $ **FLOATING
C4129 vdd2.n566 vss 4.18fF $ **FLOATING
C4130 vdd2.n567 vss 4.39fF $ **FLOATING
C4131 vdd2.n568 vss 4.39fF $ **FLOATING
C4132 vdd2.n569 vss 4.39fF $ **FLOATING
C4133 vdd2.n570 vss 4.50fF $ **FLOATING
C4134 vdd2.n571 vss 4.50fF $ **FLOATING
C4135 vdd2.n572 vss 4.39fF $ **FLOATING
C4136 vdd2.n573 vss 4.39fF $ **FLOATING
C4137 vdd2.n574 vss 4.39fF $ **FLOATING
C4138 vdd2.n575 vss 4.00fF $ **FLOATING
C4139 vdd2.n576 vss 35.61fF $ **FLOATING
C4140 vdd2.n577 vss 4.18fF $ **FLOATING
C4141 vdd2.n578 vss 4.39fF $ **FLOATING
C4142 vdd2.n579 vss 4.39fF $ **FLOATING
C4143 vdd2.n580 vss 4.39fF $ **FLOATING
C4144 vdd2.n581 vss 4.50fF $ **FLOATING
C4145 vdd2.n582 vss 4.50fF $ **FLOATING
C4146 vdd2.n583 vss 4.39fF $ **FLOATING
C4147 vdd2.n584 vss 4.39fF $ **FLOATING
C4148 vdd2.n585 vss 4.39fF $ **FLOATING
C4149 vdd2.n586 vss 4.00fF $ **FLOATING
C4150 vdd2.n587 vss 35.61fF $ **FLOATING
C4151 vdd2.n588 vss 4.18fF $ **FLOATING
C4152 vdd2.n589 vss 4.39fF $ **FLOATING
C4153 vdd2.n590 vss 4.39fF $ **FLOATING
C4154 vdd2.n591 vss 4.39fF $ **FLOATING
C4155 vdd2.n592 vss 4.50fF $ **FLOATING
C4156 vdd2.n593 vss 4.50fF $ **FLOATING
C4157 vdd2.n594 vss 4.39fF $ **FLOATING
C4158 vdd2.n595 vss 4.39fF $ **FLOATING
C4159 vdd2.n596 vss 4.39fF $ **FLOATING
C4160 vdd2.n597 vss 4.00fF $ **FLOATING
C4161 vdd2.n598 vss 35.61fF $ **FLOATING
C4162 vdd2.n599 vss 4.18fF $ **FLOATING
C4163 vdd2.n600 vss 4.39fF $ **FLOATING
C4164 vdd2.n601 vss 4.39fF $ **FLOATING
C4165 vdd2.n602 vss 4.39fF $ **FLOATING
C4166 vdd2.n603 vss 4.50fF $ **FLOATING
C4167 vdd2.n604 vss 4.50fF $ **FLOATING
C4168 vdd2.n605 vss 4.39fF $ **FLOATING
C4169 vdd2.n606 vss 4.39fF $ **FLOATING
C4170 vdd2.n607 vss 4.39fF $ **FLOATING
C4171 vdd2.n608 vss 4.00fF $ **FLOATING
C4172 vdd2.n609 vss 35.61fF $ **FLOATING
C4173 vdd2.n610 vss 4.18fF $ **FLOATING
C4174 vdd2.n611 vss 4.39fF $ **FLOATING
C4175 vdd2.n612 vss 4.39fF $ **FLOATING
C4176 vdd2.n613 vss 4.39fF $ **FLOATING
C4177 vdd2.n614 vss 4.50fF $ **FLOATING
C4178 vdd2.n615 vss 4.50fF $ **FLOATING
C4179 vdd2.n616 vss 4.39fF $ **FLOATING
C4180 vdd2.n617 vss 4.39fF $ **FLOATING
C4181 vdd2.n618 vss 4.39fF $ **FLOATING
C4182 vdd2.n619 vss 4.00fF $ **FLOATING
C4183 vdd2.n620 vss 35.61fF $ **FLOATING
C4184 vdd2.n621 vss 4.18fF $ **FLOATING
C4185 vdd2.n622 vss 4.39fF $ **FLOATING
C4186 vdd2.n623 vss 4.39fF $ **FLOATING
C4187 vdd2.n624 vss 4.39fF $ **FLOATING
C4188 vdd2.n625 vss 4.50fF $ **FLOATING
C4189 vdd2.n626 vss 4.50fF $ **FLOATING
C4190 vdd2.n627 vss 4.39fF $ **FLOATING
C4191 vdd2.n628 vss 4.39fF $ **FLOATING
C4192 vdd2.n629 vss 4.39fF $ **FLOATING
C4193 vdd2.n630 vss 4.00fF $ **FLOATING
C4194 vdd2.n631 vss 35.61fF $ **FLOATING
C4195 vdd2.n632 vss 4.18fF $ **FLOATING
C4196 vdd2.n633 vss 4.39fF $ **FLOATING
C4197 vdd2.n634 vss 4.39fF $ **FLOATING
C4198 vdd2.n635 vss 4.39fF $ **FLOATING
C4199 vdd2.n636 vss 4.50fF $ **FLOATING
C4200 vdd2.n637 vss 4.50fF $ **FLOATING
C4201 vdd2.n638 vss 4.39fF $ **FLOATING
C4202 vdd2.n639 vss 4.39fF $ **FLOATING
C4203 vdd2.n640 vss 4.39fF $ **FLOATING
C4204 vdd2.n641 vss 4.00fF $ **FLOATING
C4205 vdd2.n642 vss 35.61fF $ **FLOATING
C4206 vdd2.n643 vss 4.18fF $ **FLOATING
C4207 vdd2.n644 vss 4.39fF $ **FLOATING
C4208 vdd2.n645 vss 4.39fF $ **FLOATING
C4209 vdd2.n646 vss 4.39fF $ **FLOATING
C4210 vdd2.n647 vss 4.50fF $ **FLOATING
C4211 vdd2.n648 vss 4.50fF $ **FLOATING
C4212 vdd2.n649 vss 4.39fF $ **FLOATING
C4213 vdd2.n650 vss 4.39fF $ **FLOATING
C4214 vdd2.n651 vss 4.39fF $ **FLOATING
C4215 vdd2.n652 vss 4.00fF $ **FLOATING
C4216 vdd2.n653 vss 35.61fF $ **FLOATING
C4217 vdd2.n654 vss 4.18fF $ **FLOATING
C4218 vdd2.n655 vss 4.39fF $ **FLOATING
C4219 vdd2.n656 vss 4.39fF $ **FLOATING
C4220 vdd2.n657 vss 4.39fF $ **FLOATING
C4221 vdd2.n658 vss 4.50fF $ **FLOATING
C4222 vdd2.n659 vss 4.50fF $ **FLOATING
C4223 vdd2.n660 vss 4.39fF $ **FLOATING
C4224 vdd2.n661 vss 4.39fF $ **FLOATING
C4225 vdd2.n662 vss 4.39fF $ **FLOATING
C4226 vdd2.n663 vss 4.00fF $ **FLOATING
C4227 vdd2.n664 vss 35.61fF $ **FLOATING
C4228 vdd2.n665 vss 4.18fF $ **FLOATING
C4229 vdd2.n666 vss 4.39fF $ **FLOATING
C4230 vdd2.n667 vss 4.39fF $ **FLOATING
C4231 vdd2.n668 vss 4.39fF $ **FLOATING
C4232 vdd2.n669 vss 4.50fF $ **FLOATING
C4233 vdd2.n670 vss 4.50fF $ **FLOATING
C4234 vdd2.n671 vss 4.39fF $ **FLOATING
C4235 vdd2.n672 vss 4.39fF $ **FLOATING
C4236 vdd2.n673 vss 4.39fF $ **FLOATING
C4237 vdd2.n674 vss 4.00fF $ **FLOATING
C4238 vdd2.n675 vss 35.61fF $ **FLOATING
C4239 vdd2.n676 vss 4.18fF $ **FLOATING
C4240 vdd2.n677 vss 4.39fF $ **FLOATING
C4241 vdd2.n678 vss 4.39fF $ **FLOATING
C4242 vdd2.n679 vss 4.39fF $ **FLOATING
C4243 vdd2.n680 vss 4.50fF $ **FLOATING
C4244 vdd2.n681 vss 4.50fF $ **FLOATING
C4245 vdd2.n682 vss 4.39fF $ **FLOATING
C4246 vdd2.n683 vss 4.39fF $ **FLOATING
C4247 vdd2.n684 vss 4.39fF $ **FLOATING
C4248 vdd2.n685 vss 4.00fF $ **FLOATING
C4249 vdd2.n686 vss 35.61fF $ **FLOATING
C4250 vdd2.n687 vss 4.18fF $ **FLOATING
C4251 vdd2.n688 vss 4.39fF $ **FLOATING
C4252 vdd2.n689 vss 4.39fF $ **FLOATING
C4253 vdd2.n690 vss 4.39fF $ **FLOATING
C4254 vdd2.n691 vss 4.50fF $ **FLOATING
C4255 vdd2.n692 vss 4.50fF $ **FLOATING
C4256 vdd2.n693 vss 4.39fF $ **FLOATING
C4257 vdd2.n694 vss 4.39fF $ **FLOATING
C4258 vdd2.n695 vss 4.39fF $ **FLOATING
C4259 vdd2.n696 vss 4.00fF $ **FLOATING
C4260 vdd2.n697 vss 35.61fF $ **FLOATING
C4261 vdd2.n698 vss 4.18fF $ **FLOATING
C4262 vdd2.n699 vss 4.39fF $ **FLOATING
C4263 vdd2.n700 vss 4.39fF $ **FLOATING
C4264 vdd2.n701 vss 4.39fF $ **FLOATING
C4265 vdd2.n702 vss 4.50fF $ **FLOATING
C4266 vdd2.n703 vss 4.50fF $ **FLOATING
C4267 vdd2.n704 vss 4.39fF $ **FLOATING
C4268 vdd2.n705 vss 4.39fF $ **FLOATING
C4269 vdd2.n706 vss 4.39fF $ **FLOATING
C4270 vdd2.n707 vss 4.00fF $ **FLOATING
C4271 vdd2.n708 vss 35.61fF $ **FLOATING
C4272 vdd2.n709 vss 4.18fF $ **FLOATING
C4273 vdd2.n710 vss 4.39fF $ **FLOATING
C4274 vdd2.n711 vss 4.39fF $ **FLOATING
C4275 vdd2.n712 vss 4.39fF $ **FLOATING
C4276 vdd2.n713 vss 4.50fF $ **FLOATING
C4277 vdd2.n714 vss 4.50fF $ **FLOATING
C4278 vdd2.n715 vss 4.39fF $ **FLOATING
C4279 vdd2.n716 vss 4.39fF $ **FLOATING
C4280 vdd2.n717 vss 4.39fF $ **FLOATING
C4281 vdd2.n718 vss 4.00fF $ **FLOATING
C4282 vdd2.n719 vss 35.61fF $ **FLOATING
C4283 vdd2.n720 vss 4.18fF $ **FLOATING
C4284 vdd2.n721 vss 4.39fF $ **FLOATING
C4285 vdd2.n722 vss 4.39fF $ **FLOATING
C4286 vdd2.n723 vss 4.39fF $ **FLOATING
C4287 vdd2.n724 vss 4.50fF $ **FLOATING
C4288 vdd2.n725 vss 4.50fF $ **FLOATING
C4289 vdd2.n726 vss 4.39fF $ **FLOATING
C4290 vdd2.n727 vss 4.39fF $ **FLOATING
C4291 vdd2.n728 vss 4.39fF $ **FLOATING
C4292 vdd2.n729 vss 4.00fF $ **FLOATING
C4293 vdd2.n730 vss 35.61fF $ **FLOATING
C4294 vdd2.n731 vss 4.18fF $ **FLOATING
C4295 vdd2.n732 vss 4.39fF $ **FLOATING
C4296 vdd2.n733 vss 4.39fF $ **FLOATING
C4297 vdd2.n734 vss 4.39fF $ **FLOATING
C4298 vdd2.n735 vss 4.50fF $ **FLOATING
C4299 vdd2.n736 vss 4.50fF $ **FLOATING
C4300 vdd2.n737 vss 4.39fF $ **FLOATING
C4301 vdd2.n738 vss 4.39fF $ **FLOATING
C4302 vdd2.n739 vss 4.39fF $ **FLOATING
C4303 vdd2.n740 vss 4.00fF $ **FLOATING
C4304 vdd2.n741 vss 35.61fF $ **FLOATING
C4305 vdd2.n742 vss 4.18fF $ **FLOATING
C4306 vdd2.n743 vss 4.39fF $ **FLOATING
C4307 vdd2.n744 vss 4.39fF $ **FLOATING
C4308 vdd2.n745 vss 4.39fF $ **FLOATING
C4309 vdd2.n746 vss 4.50fF $ **FLOATING
C4310 vdd2.n747 vss 4.50fF $ **FLOATING
C4311 vdd2.n748 vss 4.39fF $ **FLOATING
C4312 vdd2.n749 vss 4.39fF $ **FLOATING
C4313 vdd2.n750 vss 4.39fF $ **FLOATING
C4314 vdd2.n751 vss 4.00fF $ **FLOATING
C4315 vdd2.n752 vss 35.61fF $ **FLOATING
C4316 vdd2.n753 vss 4.18fF $ **FLOATING
C4317 vdd2.n754 vss 4.39fF $ **FLOATING
C4318 vdd2.n755 vss 4.39fF $ **FLOATING
C4319 vdd2.n756 vss 4.39fF $ **FLOATING
C4320 vdd2.n757 vss 4.50fF $ **FLOATING
C4321 vdd2.n758 vss 4.50fF $ **FLOATING
C4322 vdd2.n759 vss 4.39fF $ **FLOATING
C4323 vdd2.n760 vss 4.39fF $ **FLOATING
C4324 vdd2.n761 vss 4.39fF $ **FLOATING
C4325 vdd2.n762 vss 4.00fF $ **FLOATING
C4326 vdd2.n763 vss 35.61fF $ **FLOATING
C4327 vdd2.n764 vss 4.18fF $ **FLOATING
C4328 vdd2.n765 vss 4.39fF $ **FLOATING
C4329 vdd2.n766 vss 4.39fF $ **FLOATING
C4330 vdd2.n767 vss 4.39fF $ **FLOATING
C4331 vdd2.n768 vss 4.50fF $ **FLOATING
C4332 vdd2.n769 vss 4.50fF $ **FLOATING
C4333 vdd2.n770 vss 4.39fF $ **FLOATING
C4334 vdd2.n771 vss 4.39fF $ **FLOATING
C4335 vdd2.n772 vss 4.39fF $ **FLOATING
C4336 vdd2.n773 vss 4.00fF $ **FLOATING
C4337 vdd2.n774 vss 35.61fF $ **FLOATING
C4338 vdd2.n775 vss 4.18fF $ **FLOATING
C4339 vdd2.n776 vss 4.39fF $ **FLOATING
C4340 vdd2.n777 vss 4.39fF $ **FLOATING
C4341 vdd2.n778 vss 4.39fF $ **FLOATING
C4342 vdd2.n779 vss 4.50fF $ **FLOATING
C4343 vdd2.n780 vss 4.50fF $ **FLOATING
C4344 vdd2.n781 vss 4.39fF $ **FLOATING
C4345 vdd2.n782 vss 4.39fF $ **FLOATING
C4346 vdd2.n783 vss 4.39fF $ **FLOATING
C4347 vdd2.n784 vss 4.00fF $ **FLOATING
C4348 vdd2.n785 vss 35.61fF $ **FLOATING
C4349 vdd2.n786 vss 4.18fF $ **FLOATING
C4350 vdd2.n787 vss 4.39fF $ **FLOATING
C4351 vdd2.n788 vss 4.39fF $ **FLOATING
C4352 vdd2.n789 vss 4.39fF $ **FLOATING
C4353 vdd2.n790 vss 4.50fF $ **FLOATING
C4354 vdd2.n791 vss 4.50fF $ **FLOATING
C4355 vdd2.n792 vss 4.39fF $ **FLOATING
C4356 vdd2.n793 vss 4.39fF $ **FLOATING
C4357 vdd2.n794 vss 4.39fF $ **FLOATING
C4358 vdd2.n795 vss 4.00fF $ **FLOATING
C4359 vdd2.n796 vss 35.61fF $ **FLOATING
C4360 vdd2.n797 vss 4.18fF $ **FLOATING
C4361 vdd2.n798 vss 4.39fF $ **FLOATING
C4362 vdd2.n799 vss 4.39fF $ **FLOATING
C4363 vdd2.n800 vss 4.39fF $ **FLOATING
C4364 vdd2.n801 vss 4.50fF $ **FLOATING
C4365 vdd2.n802 vss 4.50fF $ **FLOATING
C4366 vdd2.n803 vss 4.39fF $ **FLOATING
C4367 vdd2.n804 vss 4.39fF $ **FLOATING
C4368 vdd2.n805 vss 4.39fF $ **FLOATING
C4369 vdd2.n806 vss 4.00fF $ **FLOATING
C4370 vdd2.n807 vss 35.61fF $ **FLOATING
C4371 vdd2.n808 vss 4.18fF $ **FLOATING
C4372 vdd2.n809 vss 4.39fF $ **FLOATING
C4373 vdd2.n810 vss 4.39fF $ **FLOATING
C4374 vdd2.n811 vss 4.39fF $ **FLOATING
C4375 vdd2.n812 vss 4.50fF $ **FLOATING
C4376 vdd2.n813 vss 4.50fF $ **FLOATING
C4377 vdd2.n814 vss 4.39fF $ **FLOATING
C4378 vdd2.n815 vss 4.39fF $ **FLOATING
C4379 vdd2.n816 vss 4.39fF $ **FLOATING
C4380 vdd2.n817 vss 4.00fF $ **FLOATING
C4381 vdd2.n818 vss 35.61fF $ **FLOATING
C4382 vdd2.n819 vss 4.18fF $ **FLOATING
C4383 vdd2.n820 vss 4.39fF $ **FLOATING
C4384 vdd2.n821 vss 4.39fF $ **FLOATING
C4385 vdd2.n822 vss 4.39fF $ **FLOATING
C4386 vdd2.n823 vss 4.50fF $ **FLOATING
C4387 vdd2.n824 vss 4.50fF $ **FLOATING
C4388 vdd2.n825 vss 4.39fF $ **FLOATING
C4389 vdd2.n826 vss 4.39fF $ **FLOATING
C4390 vdd2.n827 vss 4.39fF $ **FLOATING
C4391 vdd2.n828 vss 4.00fF $ **FLOATING
C4392 vdd2.n829 vss 35.61fF $ **FLOATING
C4393 vdd2.n830 vss 4.18fF $ **FLOATING
C4394 vdd2.n831 vss 4.39fF $ **FLOATING
C4395 vdd2.n832 vss 4.39fF $ **FLOATING
C4396 vdd2.n833 vss 4.39fF $ **FLOATING
C4397 vdd2.n834 vss 4.50fF $ **FLOATING
C4398 vdd2.n835 vss 4.50fF $ **FLOATING
C4399 vdd2.n836 vss 4.39fF $ **FLOATING
C4400 vdd2.n837 vss 4.39fF $ **FLOATING
C4401 vdd2.n838 vss 4.39fF $ **FLOATING
C4402 vdd2.n839 vss 4.00fF $ **FLOATING
C4403 vdd2.n840 vss 35.61fF $ **FLOATING
C4404 vdd2.n841 vss 4.18fF $ **FLOATING
C4405 vdd2.n842 vss 4.39fF $ **FLOATING
C4406 vdd2.n843 vss 4.39fF $ **FLOATING
C4407 vdd2.n844 vss 4.39fF $ **FLOATING
C4408 vdd2.n845 vss 4.50fF $ **FLOATING
C4409 vdd2.n846 vss 4.50fF $ **FLOATING
C4410 vdd2.n847 vss 4.39fF $ **FLOATING
C4411 vdd2.n848 vss 4.39fF $ **FLOATING
C4412 vdd2.n849 vss 4.39fF $ **FLOATING
C4413 vdd2.n850 vss 4.00fF $ **FLOATING
C4414 vdd2.n851 vss 31.18fF $ **FLOATING
C4415 vdd2.n852 vss 31.86fF $ **FLOATING
C4416 vdd2.n853 vss 36.84fF $ **FLOATING
C4417 vn_p.n0 vss 1.05fF $ **FLOATING
C4418 vn_p.n76 vss 1.09fF $ **FLOATING
C4419 vn_p.n78 vss 1.03fF $ **FLOATING
C4420 vn_p.n80 vss 1.03fF $ **FLOATING
C4421 vn_p.n82 vss 1.03fF $ **FLOATING
C4422 vn_p.n84 vss 1.03fF $ **FLOATING
C4423 vn_p.n86 vss 1.03fF $ **FLOATING
C4424 vn_p.n88 vss 1.03fF $ **FLOATING
C4425 vn_p.n90 vss 1.03fF $ **FLOATING
C4426 vn_p.n92 vss 1.03fF $ **FLOATING
C4427 vn_p.n94 vss 1.03fF $ **FLOATING
C4428 vn_p.n96 vss 1.03fF $ **FLOATING
C4429 vn_p.n98 vss 1.03fF $ **FLOATING
C4430 vn_p.n100 vss 1.03fF $ **FLOATING
C4431 vn_p.n102 vss 1.03fF $ **FLOATING
C4432 vn_p.n104 vss 1.03fF $ **FLOATING
C4433 vn_p.n106 vss 1.03fF $ **FLOATING
C4434 vn_p.n108 vss 1.03fF $ **FLOATING
C4435 vn_p.n110 vss 1.03fF $ **FLOATING
C4436 vn_p.n112 vss 1.03fF $ **FLOATING
C4437 vn_p.n114 vss 1.03fF $ **FLOATING
C4438 vn_p.n116 vss 1.03fF $ **FLOATING
C4439 vn_p.n118 vss 1.03fF $ **FLOATING
C4440 vn_p.n120 vss 1.03fF $ **FLOATING
C4441 vn_p.n122 vss 1.03fF $ **FLOATING
C4442 vn_p.n124 vss 1.03fF $ **FLOATING
C4443 vn_p.n126 vss 1.03fF $ **FLOATING
C4444 vn_p.n128 vss 1.03fF $ **FLOATING
C4445 vn_p.n130 vss 1.03fF $ **FLOATING
C4446 vn_p.n132 vss 1.03fF $ **FLOATING
C4447 vn_p.n134 vss 1.03fF $ **FLOATING
C4448 vn_p.n136 vss 1.03fF $ **FLOATING
C4449 vn_p.n138 vss 1.03fF $ **FLOATING
C4450 vn_p.n140 vss 1.03fF $ **FLOATING
C4451 vn_p.n142 vss 1.03fF $ **FLOATING
C4452 vn_p.n144 vss 1.03fF $ **FLOATING
C4453 vn_p.n146 vss 1.03fF $ **FLOATING
C4454 vn_p.n148 vss 1.03fF $ **FLOATING
C4455 vn_p.n150 vss 1.03fF $ **FLOATING
C4456 vn_p.n152 vss 1.03fF $ **FLOATING
C4457 vn_p.n154 vss 1.03fF $ **FLOATING
C4458 vn_p.n156 vss 1.03fF $ **FLOATING
C4459 vn_p.n158 vss 1.03fF $ **FLOATING
C4460 vn_p.n160 vss 1.03fF $ **FLOATING
C4461 vn_p.n162 vss 1.03fF $ **FLOATING
C4462 vn_p.n164 vss 1.03fF $ **FLOATING
C4463 vn_p.n166 vss 1.03fF $ **FLOATING
C4464 vn_p.n168 vss 1.03fF $ **FLOATING
C4465 vn_p.n170 vss 1.03fF $ **FLOATING
C4466 vn_p.n172 vss 1.03fF $ **FLOATING
C4467 vn_p.n174 vss 1.03fF $ **FLOATING
C4468 vn_p.n176 vss 1.03fF $ **FLOATING
C4469 vn_p.n178 vss 1.03fF $ **FLOATING
C4470 vn_p.n180 vss 1.03fF $ **FLOATING
C4471 vn_p.n182 vss 1.03fF $ **FLOATING
C4472 vn_p.n184 vss 1.03fF $ **FLOATING
C4473 vn_p.n186 vss 1.03fF $ **FLOATING
C4474 vn_p.n188 vss 1.03fF $ **FLOATING
C4475 vn_p.n190 vss 1.03fF $ **FLOATING
C4476 vn_p.n192 vss 1.03fF $ **FLOATING
C4477 vn_p.n194 vss 1.03fF $ **FLOATING
C4478 vn_p.n196 vss 1.03fF $ **FLOATING
C4479 vn_p.n198 vss 1.03fF $ **FLOATING
C4480 vn_p.n200 vss 1.03fF $ **FLOATING
C4481 vn_p.n202 vss 1.03fF $ **FLOATING
C4482 vn_p.n204 vss 1.03fF $ **FLOATING
C4483 vn_p.n206 vss 1.03fF $ **FLOATING
C4484 vn_p.n208 vss 1.03fF $ **FLOATING
C4485 vn_p.n210 vss 1.03fF $ **FLOATING
C4486 vn_p.n212 vss 1.03fF $ **FLOATING
C4487 vn_p.n214 vss 1.03fF $ **FLOATING
C4488 vn_p.n216 vss 1.03fF $ **FLOATING
C4489 vn_p.n218 vss 1.03fF $ **FLOATING
C4490 vn_p.n220 vss 1.03fF $ **FLOATING
C4491 vn_p.n225 vss 1.09fF $ **FLOATING
C4492 vn_p.n227 vss 1.03fF $ **FLOATING
C4493 vn_p.n229 vss 1.03fF $ **FLOATING
C4494 vn_p.n231 vss 1.03fF $ **FLOATING
C4495 vn_p.n233 vss 1.03fF $ **FLOATING
C4496 vn_p.n235 vss 1.03fF $ **FLOATING
C4497 vn_p.n237 vss 1.03fF $ **FLOATING
C4498 vn_p.n239 vss 1.03fF $ **FLOATING
C4499 vn_p.n241 vss 1.03fF $ **FLOATING
C4500 vn_p.n243 vss 1.03fF $ **FLOATING
C4501 vn_p.n245 vss 1.03fF $ **FLOATING
C4502 vn_p.n247 vss 1.03fF $ **FLOATING
C4503 vn_p.n249 vss 1.03fF $ **FLOATING
C4504 vn_p.n251 vss 1.03fF $ **FLOATING
C4505 vn_p.n253 vss 1.03fF $ **FLOATING
C4506 vn_p.n255 vss 1.03fF $ **FLOATING
C4507 vn_p.n257 vss 1.03fF $ **FLOATING
C4508 vn_p.n259 vss 1.03fF $ **FLOATING
C4509 vn_p.n261 vss 1.03fF $ **FLOATING
C4510 vn_p.n263 vss 1.03fF $ **FLOATING
C4511 vn_p.n265 vss 1.03fF $ **FLOATING
C4512 vn_p.n267 vss 1.03fF $ **FLOATING
C4513 vn_p.n269 vss 1.03fF $ **FLOATING
C4514 vn_p.n271 vss 1.03fF $ **FLOATING
C4515 vn_p.n273 vss 1.03fF $ **FLOATING
C4516 vn_p.n275 vss 1.03fF $ **FLOATING
C4517 vn_p.n277 vss 1.03fF $ **FLOATING
C4518 vn_p.n279 vss 1.03fF $ **FLOATING
C4519 vn_p.n281 vss 1.03fF $ **FLOATING
C4520 vn_p.n283 vss 1.03fF $ **FLOATING
C4521 vn_p.n285 vss 1.03fF $ **FLOATING
C4522 vn_p.n287 vss 1.03fF $ **FLOATING
C4523 vn_p.n289 vss 1.03fF $ **FLOATING
C4524 vn_p.n291 vss 1.03fF $ **FLOATING
C4525 vn_p.n293 vss 1.03fF $ **FLOATING
C4526 vn_p.n295 vss 1.03fF $ **FLOATING
C4527 vn_p.n297 vss 1.03fF $ **FLOATING
C4528 vn_p.n299 vss 1.03fF $ **FLOATING
C4529 vn_p.n301 vss 1.03fF $ **FLOATING
C4530 vn_p.n303 vss 1.03fF $ **FLOATING
C4531 vn_p.n305 vss 1.03fF $ **FLOATING
C4532 vn_p.n307 vss 1.03fF $ **FLOATING
C4533 vn_p.n309 vss 1.03fF $ **FLOATING
C4534 vn_p.n311 vss 1.03fF $ **FLOATING
C4535 vn_p.n313 vss 1.03fF $ **FLOATING
C4536 vn_p.n315 vss 1.03fF $ **FLOATING
C4537 vn_p.n317 vss 1.03fF $ **FLOATING
C4538 vn_p.n319 vss 1.03fF $ **FLOATING
C4539 vn_p.n321 vss 1.03fF $ **FLOATING
C4540 vn_p.n323 vss 1.03fF $ **FLOATING
C4541 vn_p.n325 vss 1.03fF $ **FLOATING
C4542 vn_p.n327 vss 1.03fF $ **FLOATING
C4543 vn_p.n329 vss 1.03fF $ **FLOATING
C4544 vn_p.n331 vss 1.03fF $ **FLOATING
C4545 vn_p.n333 vss 1.03fF $ **FLOATING
C4546 vn_p.n335 vss 1.03fF $ **FLOATING
C4547 vn_p.n337 vss 1.03fF $ **FLOATING
C4548 vn_p.n339 vss 1.03fF $ **FLOATING
C4549 vn_p.n341 vss 1.03fF $ **FLOATING
C4550 vn_p.n343 vss 1.03fF $ **FLOATING
C4551 vn_p.n345 vss 1.03fF $ **FLOATING
C4552 vn_p.n347 vss 1.03fF $ **FLOATING
C4553 vn_p.n349 vss 1.03fF $ **FLOATING
C4554 vn_p.n351 vss 1.03fF $ **FLOATING
C4555 vn_p.n353 vss 1.03fF $ **FLOATING
C4556 vn_p.n355 vss 1.03fF $ **FLOATING
C4557 vn_p.n357 vss 1.03fF $ **FLOATING
C4558 vn_p.n359 vss 1.03fF $ **FLOATING
C4559 vn_p.n361 vss 1.03fF $ **FLOATING
C4560 vn_p.n363 vss 1.03fF $ **FLOATING
C4561 vn_p.n365 vss 1.03fF $ **FLOATING
C4562 vn_p.n367 vss 1.03fF $ **FLOATING
C4563 vn_p.n369 vss 1.03fF $ **FLOATING
C4564 vn_p.n374 vss 1.09fF $ **FLOATING
C4565 vn_p.n376 vss 1.03fF $ **FLOATING
C4566 vn_p.n378 vss 1.03fF $ **FLOATING
C4567 vn_p.n380 vss 1.03fF $ **FLOATING
C4568 vn_p.n382 vss 1.03fF $ **FLOATING
C4569 vn_p.n384 vss 1.03fF $ **FLOATING
C4570 vn_p.n386 vss 1.03fF $ **FLOATING
C4571 vn_p.n388 vss 1.03fF $ **FLOATING
C4572 vn_p.n390 vss 1.03fF $ **FLOATING
C4573 vn_p.n392 vss 1.03fF $ **FLOATING
C4574 vn_p.n394 vss 1.03fF $ **FLOATING
C4575 vn_p.n396 vss 1.03fF $ **FLOATING
C4576 vn_p.n398 vss 1.03fF $ **FLOATING
C4577 vn_p.n400 vss 1.03fF $ **FLOATING
C4578 vn_p.n402 vss 1.03fF $ **FLOATING
C4579 vn_p.n404 vss 1.03fF $ **FLOATING
C4580 vn_p.n406 vss 1.03fF $ **FLOATING
C4581 vn_p.n408 vss 1.03fF $ **FLOATING
C4582 vn_p.n410 vss 1.03fF $ **FLOATING
C4583 vn_p.n412 vss 1.03fF $ **FLOATING
C4584 vn_p.n414 vss 1.03fF $ **FLOATING
C4585 vn_p.n416 vss 1.03fF $ **FLOATING
C4586 vn_p.n418 vss 1.03fF $ **FLOATING
C4587 vn_p.n420 vss 1.03fF $ **FLOATING
C4588 vn_p.n422 vss 1.03fF $ **FLOATING
C4589 vn_p.n424 vss 1.03fF $ **FLOATING
C4590 vn_p.n426 vss 1.03fF $ **FLOATING
C4591 vn_p.n428 vss 1.03fF $ **FLOATING
C4592 vn_p.n430 vss 1.03fF $ **FLOATING
C4593 vn_p.n432 vss 1.03fF $ **FLOATING
C4594 vn_p.n434 vss 1.03fF $ **FLOATING
C4595 vn_p.n436 vss 1.03fF $ **FLOATING
C4596 vn_p.n438 vss 1.03fF $ **FLOATING
C4597 vn_p.n440 vss 1.03fF $ **FLOATING
C4598 vn_p.n442 vss 1.03fF $ **FLOATING
C4599 vn_p.n444 vss 1.03fF $ **FLOATING
C4600 vn_p.n446 vss 1.03fF $ **FLOATING
C4601 vn_p.n448 vss 1.03fF $ **FLOATING
C4602 vn_p.n450 vss 1.03fF $ **FLOATING
C4603 vn_p.n452 vss 1.03fF $ **FLOATING
C4604 vn_p.n454 vss 1.03fF $ **FLOATING
C4605 vn_p.n456 vss 1.03fF $ **FLOATING
C4606 vn_p.n458 vss 1.03fF $ **FLOATING
C4607 vn_p.n460 vss 1.03fF $ **FLOATING
C4608 vn_p.n462 vss 1.03fF $ **FLOATING
C4609 vn_p.n464 vss 1.03fF $ **FLOATING
C4610 vn_p.n466 vss 1.03fF $ **FLOATING
C4611 vn_p.n468 vss 1.03fF $ **FLOATING
C4612 vn_p.n470 vss 1.03fF $ **FLOATING
C4613 vn_p.n472 vss 1.03fF $ **FLOATING
C4614 vn_p.n474 vss 1.03fF $ **FLOATING
C4615 vn_p.n476 vss 1.03fF $ **FLOATING
C4616 vn_p.n478 vss 1.03fF $ **FLOATING
C4617 vn_p.n480 vss 1.03fF $ **FLOATING
C4618 vn_p.n482 vss 1.03fF $ **FLOATING
C4619 vn_p.n484 vss 1.03fF $ **FLOATING
C4620 vn_p.n486 vss 1.03fF $ **FLOATING
C4621 vn_p.n488 vss 1.03fF $ **FLOATING
C4622 vn_p.n490 vss 1.03fF $ **FLOATING
C4623 vn_p.n492 vss 1.03fF $ **FLOATING
C4624 vn_p.n494 vss 1.03fF $ **FLOATING
C4625 vn_p.n496 vss 1.03fF $ **FLOATING
C4626 vn_p.n498 vss 1.03fF $ **FLOATING
C4627 vn_p.n500 vss 1.03fF $ **FLOATING
C4628 vn_p.n502 vss 1.03fF $ **FLOATING
C4629 vn_p.n504 vss 1.03fF $ **FLOATING
C4630 vn_p.n506 vss 1.03fF $ **FLOATING
C4631 vn_p.n508 vss 1.03fF $ **FLOATING
C4632 vn_p.n510 vss 1.03fF $ **FLOATING
C4633 vn_p.n512 vss 1.03fF $ **FLOATING
C4634 vn_p.n514 vss 1.03fF $ **FLOATING
C4635 vn_p.n516 vss 1.03fF $ **FLOATING
C4636 vn_p.n518 vss 1.03fF $ **FLOATING
C4637 vn_p.n523 vss 1.09fF $ **FLOATING
C4638 vn_p.n525 vss 1.03fF $ **FLOATING
C4639 vn_p.n527 vss 1.03fF $ **FLOATING
C4640 vn_p.n529 vss 1.03fF $ **FLOATING
C4641 vn_p.n531 vss 1.03fF $ **FLOATING
C4642 vn_p.n533 vss 1.03fF $ **FLOATING
C4643 vn_p.n535 vss 1.03fF $ **FLOATING
C4644 vn_p.n537 vss 1.03fF $ **FLOATING
C4645 vn_p.n539 vss 1.03fF $ **FLOATING
C4646 vn_p.n541 vss 1.03fF $ **FLOATING
C4647 vn_p.n543 vss 1.03fF $ **FLOATING
C4648 vn_p.n545 vss 1.03fF $ **FLOATING
C4649 vn_p.n547 vss 1.03fF $ **FLOATING
C4650 vn_p.n549 vss 1.03fF $ **FLOATING
C4651 vn_p.n551 vss 1.03fF $ **FLOATING
C4652 vn_p.n553 vss 1.03fF $ **FLOATING
C4653 vn_p.n555 vss 1.03fF $ **FLOATING
C4654 vn_p.n557 vss 1.03fF $ **FLOATING
C4655 vn_p.n559 vss 1.03fF $ **FLOATING
C4656 vn_p.n561 vss 1.03fF $ **FLOATING
C4657 vn_p.n563 vss 1.03fF $ **FLOATING
C4658 vn_p.n565 vss 1.03fF $ **FLOATING
C4659 vn_p.n567 vss 1.03fF $ **FLOATING
C4660 vn_p.n569 vss 1.03fF $ **FLOATING
C4661 vn_p.n571 vss 1.03fF $ **FLOATING
C4662 vn_p.n573 vss 1.03fF $ **FLOATING
C4663 vn_p.n575 vss 1.03fF $ **FLOATING
C4664 vn_p.n577 vss 1.03fF $ **FLOATING
C4665 vn_p.n579 vss 1.03fF $ **FLOATING
C4666 vn_p.n581 vss 1.03fF $ **FLOATING
C4667 vn_p.n583 vss 1.03fF $ **FLOATING
C4668 vn_p.n585 vss 1.03fF $ **FLOATING
C4669 vn_p.n587 vss 1.03fF $ **FLOATING
C4670 vn_p.n589 vss 1.03fF $ **FLOATING
C4671 vn_p.n591 vss 1.03fF $ **FLOATING
C4672 vn_p.n593 vss 1.03fF $ **FLOATING
C4673 vn_p.n595 vss 1.03fF $ **FLOATING
C4674 vn_p.n597 vss 1.03fF $ **FLOATING
C4675 vn_p.n599 vss 1.03fF $ **FLOATING
C4676 vn_p.n601 vss 1.03fF $ **FLOATING
C4677 vn_p.n603 vss 1.03fF $ **FLOATING
C4678 vn_p.n605 vss 1.03fF $ **FLOATING
C4679 vn_p.n607 vss 1.03fF $ **FLOATING
C4680 vn_p.n609 vss 1.03fF $ **FLOATING
C4681 vn_p.n611 vss 1.03fF $ **FLOATING
C4682 vn_p.n613 vss 1.03fF $ **FLOATING
C4683 vn_p.n615 vss 1.03fF $ **FLOATING
C4684 vn_p.n617 vss 1.03fF $ **FLOATING
C4685 vn_p.n619 vss 1.03fF $ **FLOATING
C4686 vn_p.n621 vss 1.03fF $ **FLOATING
C4687 vn_p.n623 vss 1.03fF $ **FLOATING
C4688 vn_p.n625 vss 1.03fF $ **FLOATING
C4689 vn_p.n627 vss 1.03fF $ **FLOATING
C4690 vn_p.n629 vss 1.03fF $ **FLOATING
C4691 vn_p.n631 vss 1.03fF $ **FLOATING
C4692 vn_p.n633 vss 1.03fF $ **FLOATING
C4693 vn_p.n635 vss 1.03fF $ **FLOATING
C4694 vn_p.n637 vss 1.03fF $ **FLOATING
C4695 vn_p.n639 vss 1.03fF $ **FLOATING
C4696 vn_p.n641 vss 1.03fF $ **FLOATING
C4697 vn_p.n643 vss 1.03fF $ **FLOATING
C4698 vn_p.n645 vss 1.03fF $ **FLOATING
C4699 vn_p.n647 vss 1.03fF $ **FLOATING
C4700 vn_p.n649 vss 1.03fF $ **FLOATING
C4701 vn_p.n651 vss 1.03fF $ **FLOATING
C4702 vn_p.n653 vss 1.03fF $ **FLOATING
C4703 vn_p.n655 vss 1.03fF $ **FLOATING
C4704 vn_p.n657 vss 1.03fF $ **FLOATING
C4705 vn_p.n659 vss 1.03fF $ **FLOATING
C4706 vn_p.n661 vss 1.03fF $ **FLOATING
C4707 vn_p.n663 vss 1.03fF $ **FLOATING
C4708 vn_p.n665 vss 1.03fF $ **FLOATING
C4709 vn_p.n667 vss 1.03fF $ **FLOATING
C4710 vn_p.n670 vss 1.04fF $ **FLOATING
C4711 vn_p.n743 vss 1.34fF $ **FLOATING
C4712 vn_p.n744 vss 19.04fF $ **FLOATING
C4713 vn_p.n745 vss 13.65fF $ **FLOATING
C4714 vn_p.n746 vss 13.44fF $ **FLOATING
C4715 vn_p.n747 vss 13.30fF $ **FLOATING
C4716 vn_p.n748 vss 6.61fF $ **FLOATING
C4717 vn_p.n749 vss 1.04fF $ **FLOATING
C4718 vn_p.n825 vss 1.09fF $ **FLOATING
C4719 vn_p.n827 vss 1.03fF $ **FLOATING
C4720 vn_p.n829 vss 1.03fF $ **FLOATING
C4721 vn_p.n831 vss 1.03fF $ **FLOATING
C4722 vn_p.n833 vss 1.03fF $ **FLOATING
C4723 vn_p.n835 vss 1.03fF $ **FLOATING
C4724 vn_p.n837 vss 1.03fF $ **FLOATING
C4725 vn_p.n839 vss 1.03fF $ **FLOATING
C4726 vn_p.n841 vss 1.03fF $ **FLOATING
C4727 vn_p.n843 vss 1.03fF $ **FLOATING
C4728 vn_p.n845 vss 1.03fF $ **FLOATING
C4729 vn_p.n847 vss 1.03fF $ **FLOATING
C4730 vn_p.n849 vss 1.03fF $ **FLOATING
C4731 vn_p.n851 vss 1.03fF $ **FLOATING
C4732 vn_p.n853 vss 1.03fF $ **FLOATING
C4733 vn_p.n855 vss 1.03fF $ **FLOATING
C4734 vn_p.n857 vss 1.03fF $ **FLOATING
C4735 vn_p.n859 vss 1.03fF $ **FLOATING
C4736 vn_p.n861 vss 1.03fF $ **FLOATING
C4737 vn_p.n863 vss 1.03fF $ **FLOATING
C4738 vn_p.n865 vss 1.03fF $ **FLOATING
C4739 vn_p.n867 vss 1.03fF $ **FLOATING
C4740 vn_p.n869 vss 1.03fF $ **FLOATING
C4741 vn_p.n871 vss 1.03fF $ **FLOATING
C4742 vn_p.n873 vss 1.03fF $ **FLOATING
C4743 vn_p.n875 vss 1.03fF $ **FLOATING
C4744 vn_p.n877 vss 1.03fF $ **FLOATING
C4745 vn_p.n879 vss 1.03fF $ **FLOATING
C4746 vn_p.n881 vss 1.03fF $ **FLOATING
C4747 vn_p.n883 vss 1.03fF $ **FLOATING
C4748 vn_p.n885 vss 1.03fF $ **FLOATING
C4749 vn_p.n887 vss 1.03fF $ **FLOATING
C4750 vn_p.n889 vss 1.03fF $ **FLOATING
C4751 vn_p.n891 vss 1.03fF $ **FLOATING
C4752 vn_p.n893 vss 1.03fF $ **FLOATING
C4753 vn_p.n895 vss 1.03fF $ **FLOATING
C4754 vn_p.n897 vss 1.03fF $ **FLOATING
C4755 vn_p.n899 vss 1.03fF $ **FLOATING
C4756 vn_p.n901 vss 1.03fF $ **FLOATING
C4757 vn_p.n903 vss 1.03fF $ **FLOATING
C4758 vn_p.n905 vss 1.03fF $ **FLOATING
C4759 vn_p.n907 vss 1.03fF $ **FLOATING
C4760 vn_p.n909 vss 1.03fF $ **FLOATING
C4761 vn_p.n911 vss 1.03fF $ **FLOATING
C4762 vn_p.n913 vss 1.03fF $ **FLOATING
C4763 vn_p.n915 vss 1.03fF $ **FLOATING
C4764 vn_p.n917 vss 1.03fF $ **FLOATING
C4765 vn_p.n919 vss 1.03fF $ **FLOATING
C4766 vn_p.n921 vss 1.03fF $ **FLOATING
C4767 vn_p.n923 vss 1.03fF $ **FLOATING
C4768 vn_p.n925 vss 1.03fF $ **FLOATING
C4769 vn_p.n927 vss 1.03fF $ **FLOATING
C4770 vn_p.n929 vss 1.03fF $ **FLOATING
C4771 vn_p.n931 vss 1.03fF $ **FLOATING
C4772 vn_p.n933 vss 1.03fF $ **FLOATING
C4773 vn_p.n935 vss 1.03fF $ **FLOATING
C4774 vn_p.n937 vss 1.03fF $ **FLOATING
C4775 vn_p.n939 vss 1.03fF $ **FLOATING
C4776 vn_p.n941 vss 1.03fF $ **FLOATING
C4777 vn_p.n943 vss 1.03fF $ **FLOATING
C4778 vn_p.n945 vss 1.03fF $ **FLOATING
C4779 vn_p.n947 vss 1.03fF $ **FLOATING
C4780 vn_p.n949 vss 1.03fF $ **FLOATING
C4781 vn_p.n951 vss 1.03fF $ **FLOATING
C4782 vn_p.n953 vss 1.03fF $ **FLOATING
C4783 vn_p.n955 vss 1.03fF $ **FLOATING
C4784 vn_p.n957 vss 1.03fF $ **FLOATING
C4785 vn_p.n959 vss 1.03fF $ **FLOATING
C4786 vn_p.n961 vss 1.03fF $ **FLOATING
C4787 vn_p.n963 vss 1.03fF $ **FLOATING
C4788 vn_p.n965 vss 1.03fF $ **FLOATING
C4789 vn_p.n967 vss 1.03fF $ **FLOATING
C4790 vn_p.n969 vss 1.03fF $ **FLOATING
C4791 vn_p.n974 vss 1.09fF $ **FLOATING
C4792 vn_p.n976 vss 1.03fF $ **FLOATING
C4793 vn_p.n978 vss 1.03fF $ **FLOATING
C4794 vn_p.n980 vss 1.03fF $ **FLOATING
C4795 vn_p.n982 vss 1.03fF $ **FLOATING
C4796 vn_p.n984 vss 1.03fF $ **FLOATING
C4797 vn_p.n986 vss 1.03fF $ **FLOATING
C4798 vn_p.n988 vss 1.03fF $ **FLOATING
C4799 vn_p.n990 vss 1.03fF $ **FLOATING
C4800 vn_p.n992 vss 1.03fF $ **FLOATING
C4801 vn_p.n994 vss 1.03fF $ **FLOATING
C4802 vn_p.n996 vss 1.03fF $ **FLOATING
C4803 vn_p.n998 vss 1.03fF $ **FLOATING
C4804 vn_p.n1000 vss 1.03fF $ **FLOATING
C4805 vn_p.n1002 vss 1.03fF $ **FLOATING
C4806 vn_p.n1004 vss 1.03fF $ **FLOATING
C4807 vn_p.n1006 vss 1.03fF $ **FLOATING
C4808 vn_p.n1008 vss 1.03fF $ **FLOATING
C4809 vn_p.n1010 vss 1.03fF $ **FLOATING
C4810 vn_p.n1012 vss 1.03fF $ **FLOATING
C4811 vn_p.n1014 vss 1.03fF $ **FLOATING
C4812 vn_p.n1016 vss 1.03fF $ **FLOATING
C4813 vn_p.n1018 vss 1.03fF $ **FLOATING
C4814 vn_p.n1020 vss 1.03fF $ **FLOATING
C4815 vn_p.n1022 vss 1.03fF $ **FLOATING
C4816 vn_p.n1024 vss 1.03fF $ **FLOATING
C4817 vn_p.n1026 vss 1.03fF $ **FLOATING
C4818 vn_p.n1028 vss 1.03fF $ **FLOATING
C4819 vn_p.n1030 vss 1.03fF $ **FLOATING
C4820 vn_p.n1032 vss 1.03fF $ **FLOATING
C4821 vn_p.n1034 vss 1.03fF $ **FLOATING
C4822 vn_p.n1036 vss 1.03fF $ **FLOATING
C4823 vn_p.n1038 vss 1.03fF $ **FLOATING
C4824 vn_p.n1040 vss 1.03fF $ **FLOATING
C4825 vn_p.n1042 vss 1.03fF $ **FLOATING
C4826 vn_p.n1044 vss 1.03fF $ **FLOATING
C4827 vn_p.n1046 vss 1.03fF $ **FLOATING
C4828 vn_p.n1048 vss 1.03fF $ **FLOATING
C4829 vn_p.n1050 vss 1.03fF $ **FLOATING
C4830 vn_p.n1052 vss 1.03fF $ **FLOATING
C4831 vn_p.n1054 vss 1.03fF $ **FLOATING
C4832 vn_p.n1056 vss 1.03fF $ **FLOATING
C4833 vn_p.n1058 vss 1.03fF $ **FLOATING
C4834 vn_p.n1060 vss 1.03fF $ **FLOATING
C4835 vn_p.n1062 vss 1.03fF $ **FLOATING
C4836 vn_p.n1064 vss 1.03fF $ **FLOATING
C4837 vn_p.n1066 vss 1.03fF $ **FLOATING
C4838 vn_p.n1068 vss 1.03fF $ **FLOATING
C4839 vn_p.n1070 vss 1.03fF $ **FLOATING
C4840 vn_p.n1072 vss 1.03fF $ **FLOATING
C4841 vn_p.n1074 vss 1.03fF $ **FLOATING
C4842 vn_p.n1076 vss 1.03fF $ **FLOATING
C4843 vn_p.n1078 vss 1.03fF $ **FLOATING
C4844 vn_p.n1080 vss 1.03fF $ **FLOATING
C4845 vn_p.n1082 vss 1.03fF $ **FLOATING
C4846 vn_p.n1084 vss 1.03fF $ **FLOATING
C4847 vn_p.n1086 vss 1.03fF $ **FLOATING
C4848 vn_p.n1088 vss 1.03fF $ **FLOATING
C4849 vn_p.n1090 vss 1.03fF $ **FLOATING
C4850 vn_p.n1092 vss 1.03fF $ **FLOATING
C4851 vn_p.n1094 vss 1.03fF $ **FLOATING
C4852 vn_p.n1096 vss 1.03fF $ **FLOATING
C4853 vn_p.n1098 vss 1.03fF $ **FLOATING
C4854 vn_p.n1100 vss 1.03fF $ **FLOATING
C4855 vn_p.n1102 vss 1.03fF $ **FLOATING
C4856 vn_p.n1104 vss 1.03fF $ **FLOATING
C4857 vn_p.n1106 vss 1.03fF $ **FLOATING
C4858 vn_p.n1108 vss 1.03fF $ **FLOATING
C4859 vn_p.n1110 vss 1.03fF $ **FLOATING
C4860 vn_p.n1112 vss 1.03fF $ **FLOATING
C4861 vn_p.n1114 vss 1.03fF $ **FLOATING
C4862 vn_p.n1116 vss 1.03fF $ **FLOATING
C4863 vn_p.n1118 vss 1.03fF $ **FLOATING
C4864 vn_p.n1123 vss 1.09fF $ **FLOATING
C4865 vn_p.n1125 vss 1.03fF $ **FLOATING
C4866 vn_p.n1127 vss 1.03fF $ **FLOATING
C4867 vn_p.n1129 vss 1.03fF $ **FLOATING
C4868 vn_p.n1131 vss 1.03fF $ **FLOATING
C4869 vn_p.n1133 vss 1.03fF $ **FLOATING
C4870 vn_p.n1135 vss 1.03fF $ **FLOATING
C4871 vn_p.n1137 vss 1.03fF $ **FLOATING
C4872 vn_p.n1139 vss 1.03fF $ **FLOATING
C4873 vn_p.n1141 vss 1.03fF $ **FLOATING
C4874 vn_p.n1143 vss 1.03fF $ **FLOATING
C4875 vn_p.n1145 vss 1.03fF $ **FLOATING
C4876 vn_p.n1147 vss 1.03fF $ **FLOATING
C4877 vn_p.n1149 vss 1.03fF $ **FLOATING
C4878 vn_p.n1151 vss 1.03fF $ **FLOATING
C4879 vn_p.n1153 vss 1.03fF $ **FLOATING
C4880 vn_p.n1155 vss 1.03fF $ **FLOATING
C4881 vn_p.n1157 vss 1.03fF $ **FLOATING
C4882 vn_p.n1159 vss 1.03fF $ **FLOATING
C4883 vn_p.n1161 vss 1.03fF $ **FLOATING
C4884 vn_p.n1163 vss 1.03fF $ **FLOATING
C4885 vn_p.n1165 vss 1.03fF $ **FLOATING
C4886 vn_p.n1167 vss 1.03fF $ **FLOATING
C4887 vn_p.n1169 vss 1.03fF $ **FLOATING
C4888 vn_p.n1171 vss 1.03fF $ **FLOATING
C4889 vn_p.n1173 vss 1.03fF $ **FLOATING
C4890 vn_p.n1175 vss 1.03fF $ **FLOATING
C4891 vn_p.n1177 vss 1.03fF $ **FLOATING
C4892 vn_p.n1179 vss 1.03fF $ **FLOATING
C4893 vn_p.n1181 vss 1.03fF $ **FLOATING
C4894 vn_p.n1183 vss 1.03fF $ **FLOATING
C4895 vn_p.n1185 vss 1.03fF $ **FLOATING
C4896 vn_p.n1187 vss 1.03fF $ **FLOATING
C4897 vn_p.n1189 vss 1.03fF $ **FLOATING
C4898 vn_p.n1191 vss 1.03fF $ **FLOATING
C4899 vn_p.n1193 vss 1.03fF $ **FLOATING
C4900 vn_p.n1195 vss 1.03fF $ **FLOATING
C4901 vn_p.n1197 vss 1.03fF $ **FLOATING
C4902 vn_p.n1199 vss 1.03fF $ **FLOATING
C4903 vn_p.n1201 vss 1.03fF $ **FLOATING
C4904 vn_p.n1203 vss 1.03fF $ **FLOATING
C4905 vn_p.n1205 vss 1.03fF $ **FLOATING
C4906 vn_p.n1207 vss 1.03fF $ **FLOATING
C4907 vn_p.n1209 vss 1.03fF $ **FLOATING
C4908 vn_p.n1211 vss 1.03fF $ **FLOATING
C4909 vn_p.n1213 vss 1.03fF $ **FLOATING
C4910 vn_p.n1215 vss 1.03fF $ **FLOATING
C4911 vn_p.n1217 vss 1.03fF $ **FLOATING
C4912 vn_p.n1219 vss 1.03fF $ **FLOATING
C4913 vn_p.n1221 vss 1.03fF $ **FLOATING
C4914 vn_p.n1223 vss 1.03fF $ **FLOATING
C4915 vn_p.n1225 vss 1.03fF $ **FLOATING
C4916 vn_p.n1227 vss 1.03fF $ **FLOATING
C4917 vn_p.n1229 vss 1.03fF $ **FLOATING
C4918 vn_p.n1231 vss 1.03fF $ **FLOATING
C4919 vn_p.n1233 vss 1.03fF $ **FLOATING
C4920 vn_p.n1235 vss 1.03fF $ **FLOATING
C4921 vn_p.n1237 vss 1.03fF $ **FLOATING
C4922 vn_p.n1239 vss 1.03fF $ **FLOATING
C4923 vn_p.n1241 vss 1.03fF $ **FLOATING
C4924 vn_p.n1243 vss 1.03fF $ **FLOATING
C4925 vn_p.n1245 vss 1.03fF $ **FLOATING
C4926 vn_p.n1247 vss 1.03fF $ **FLOATING
C4927 vn_p.n1249 vss 1.03fF $ **FLOATING
C4928 vn_p.n1251 vss 1.03fF $ **FLOATING
C4929 vn_p.n1253 vss 1.03fF $ **FLOATING
C4930 vn_p.n1255 vss 1.03fF $ **FLOATING
C4931 vn_p.n1257 vss 1.03fF $ **FLOATING
C4932 vn_p.n1259 vss 1.03fF $ **FLOATING
C4933 vn_p.n1261 vss 1.03fF $ **FLOATING
C4934 vn_p.n1263 vss 1.03fF $ **FLOATING
C4935 vn_p.n1265 vss 1.03fF $ **FLOATING
C4936 vn_p.n1267 vss 1.03fF $ **FLOATING
C4937 vn_p.n1272 vss 1.09fF $ **FLOATING
C4938 vn_p.n1274 vss 1.03fF $ **FLOATING
C4939 vn_p.n1276 vss 1.03fF $ **FLOATING
C4940 vn_p.n1278 vss 1.03fF $ **FLOATING
C4941 vn_p.n1280 vss 1.03fF $ **FLOATING
C4942 vn_p.n1282 vss 1.03fF $ **FLOATING
C4943 vn_p.n1284 vss 1.03fF $ **FLOATING
C4944 vn_p.n1286 vss 1.03fF $ **FLOATING
C4945 vn_p.n1288 vss 1.03fF $ **FLOATING
C4946 vn_p.n1290 vss 1.03fF $ **FLOATING
C4947 vn_p.n1292 vss 1.03fF $ **FLOATING
C4948 vn_p.n1294 vss 1.03fF $ **FLOATING
C4949 vn_p.n1296 vss 1.03fF $ **FLOATING
C4950 vn_p.n1298 vss 1.03fF $ **FLOATING
C4951 vn_p.n1300 vss 1.03fF $ **FLOATING
C4952 vn_p.n1302 vss 1.03fF $ **FLOATING
C4953 vn_p.n1304 vss 1.03fF $ **FLOATING
C4954 vn_p.n1306 vss 1.03fF $ **FLOATING
C4955 vn_p.n1308 vss 1.03fF $ **FLOATING
C4956 vn_p.n1310 vss 1.03fF $ **FLOATING
C4957 vn_p.n1312 vss 1.03fF $ **FLOATING
C4958 vn_p.n1314 vss 1.03fF $ **FLOATING
C4959 vn_p.n1316 vss 1.03fF $ **FLOATING
C4960 vn_p.n1318 vss 1.03fF $ **FLOATING
C4961 vn_p.n1320 vss 1.03fF $ **FLOATING
C4962 vn_p.n1322 vss 1.03fF $ **FLOATING
C4963 vn_p.n1324 vss 1.03fF $ **FLOATING
C4964 vn_p.n1326 vss 1.03fF $ **FLOATING
C4965 vn_p.n1328 vss 1.03fF $ **FLOATING
C4966 vn_p.n1330 vss 1.03fF $ **FLOATING
C4967 vn_p.n1332 vss 1.03fF $ **FLOATING
C4968 vn_p.n1334 vss 1.03fF $ **FLOATING
C4969 vn_p.n1336 vss 1.03fF $ **FLOATING
C4970 vn_p.n1338 vss 1.03fF $ **FLOATING
C4971 vn_p.n1340 vss 1.03fF $ **FLOATING
C4972 vn_p.n1342 vss 1.03fF $ **FLOATING
C4973 vn_p.n1344 vss 1.03fF $ **FLOATING
C4974 vn_p.n1346 vss 1.03fF $ **FLOATING
C4975 vn_p.n1348 vss 1.03fF $ **FLOATING
C4976 vn_p.n1350 vss 1.03fF $ **FLOATING
C4977 vn_p.n1352 vss 1.03fF $ **FLOATING
C4978 vn_p.n1354 vss 1.03fF $ **FLOATING
C4979 vn_p.n1356 vss 1.03fF $ **FLOATING
C4980 vn_p.n1358 vss 1.03fF $ **FLOATING
C4981 vn_p.n1360 vss 1.03fF $ **FLOATING
C4982 vn_p.n1362 vss 1.03fF $ **FLOATING
C4983 vn_p.n1364 vss 1.03fF $ **FLOATING
C4984 vn_p.n1366 vss 1.03fF $ **FLOATING
C4985 vn_p.n1368 vss 1.03fF $ **FLOATING
C4986 vn_p.n1370 vss 1.03fF $ **FLOATING
C4987 vn_p.n1372 vss 1.03fF $ **FLOATING
C4988 vn_p.n1374 vss 1.03fF $ **FLOATING
C4989 vn_p.n1376 vss 1.03fF $ **FLOATING
C4990 vn_p.n1378 vss 1.03fF $ **FLOATING
C4991 vn_p.n1380 vss 1.03fF $ **FLOATING
C4992 vn_p.n1382 vss 1.03fF $ **FLOATING
C4993 vn_p.n1384 vss 1.03fF $ **FLOATING
C4994 vn_p.n1386 vss 1.03fF $ **FLOATING
C4995 vn_p.n1388 vss 1.03fF $ **FLOATING
C4996 vn_p.n1390 vss 1.03fF $ **FLOATING
C4997 vn_p.n1392 vss 1.03fF $ **FLOATING
C4998 vn_p.n1394 vss 1.03fF $ **FLOATING
C4999 vn_p.n1396 vss 1.03fF $ **FLOATING
C5000 vn_p.n1398 vss 1.03fF $ **FLOATING
C5001 vn_p.n1400 vss 1.03fF $ **FLOATING
C5002 vn_p.n1402 vss 1.03fF $ **FLOATING
C5003 vn_p.n1404 vss 1.03fF $ **FLOATING
C5004 vn_p.n1406 vss 1.03fF $ **FLOATING
C5005 vn_p.n1408 vss 1.03fF $ **FLOATING
C5006 vn_p.n1410 vss 1.03fF $ **FLOATING
C5007 vn_p.n1412 vss 1.03fF $ **FLOATING
C5008 vn_p.n1414 vss 1.03fF $ **FLOATING
C5009 vn_p.n1416 vss 1.03fF $ **FLOATING
C5010 vn_p.n1419 vss 1.10fF $ **FLOATING
C5011 vn_p.n1492 vss 1.92fF $ **FLOATING
C5012 vn_p.n1493 vss 18.52fF $ **FLOATING
C5013 vn_p.n1494 vss 8.04fF $ **FLOATING
C5014 vn_p.n1495 vss 12.42fF $ **FLOATING
C5015 vn_p.n1496 vss 13.09fF $ **FLOATING
C5016 vn_p.n1497 vss 7.69fF $ **FLOATING
.ends
