* NGSPICE file created from triangle_post.ext - technology: sky130A

.subckt triangle_post vdd vbias1 vbias2 vref vss vsquare vt
X1 vt.t200 a_19926_13536.t17 vss.t142 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X2 vss.t170 a_19926_29936.t17 vsquare.t146 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X3 vdd.t143 vbias2.t24 vsquare.t148 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4 a_23370_8306.t11 vref.t0 a_19926_13536.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X5 vt.t46 vbias1.t24 vdd.t196 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6 vss.t145 a_19926_29936.t18 vsquare.t145 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X7 vss.t146 a_19926_29936.t19 vsquare.t144 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X8 vdd.t197 vbias1.t25 vt.t47 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X9 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X10 vt.t48 vbias1.t26 vdd.t198 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X11 a_23370_24650.t11 vref.t1 a_23744_20184.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X12 vss.t9 a_23744_20184.t18 a_23744_20184.t19 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X13 vt.t49 vbias1.t27 vdd.t199 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X14 a_23744_20184.t8 vref.t2 a_23370_24650.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X15 vsquare.t149 vbias2.t25 vdd.t142 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X16 vdd.t141 vbias2.t26 vsquare.t150 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X17 vdd.t200 vbias1.t28 vt.t50 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X18 a_19926_29936.t9 OTA_0/vp a_23370_24650.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X19 vdd.t140 vbias2.t20 vbias2.t21 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X20 vdd.t139 vbias2.t27 vsquare.t151 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X21 vss.t147 a_19926_29936.t20 vsquare.t143 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X22 vsquare.t152 vbias2.t28 vdd.t138 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X23 vt.t51 vbias1.t29 vdd.t201 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X24 vt.t199 a_19926_13536.t18 vss.t141 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X25 vdd.t137 vbias2.t29 vsquare.t153 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X26 vdd.t202 vbias1.t30 vt.t52 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X27 vdd.t136 vbias2.t30 vsquare.t154 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X28 vdd.t203 vbias1.t31 a_23370_8306.t27 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X29 vss.t148 a_19926_29936.t21 vsquare.t142 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X30 vss.t149 a_19926_29936.t22 vsquare.t141 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X31 vt.t198 a_19926_13536.t19 vss.t140 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X32 vss.t139 a_19926_13536.t20 vt.t197 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X33 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X34 vt.t196 a_19926_13536.t21 vss.t138 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X35 vss.t8 a_23744_20184.t20 a_19926_29936.t2 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X36 vdd.t204 vbias1.t32 vt.t53 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X37 vss.t150 a_19926_29936.t23 vsquare.t140 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X38 a_23370_8306.t12 OTA_tri_0/vn a_23744_3840.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X39 vdd.t135 vbias2.t31 vsquare.t155 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X40 vdd.t134 vbias2.t22 vbias2.t23 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X41 vsquare.t156 vbias2.t32 vdd.t133 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X42 vdd.t205 vbias1.t33 vt.t54 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X43 vdd.t132 vbias2.t33 vsquare.t157 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X44 vdd.t131 vbias2.t34 vsquare.t158 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X45 vss.t151 a_19926_29936.t24 vsquare.t139 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X46 vsquare.t138 a_19926_29936.t25 vss.t152 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X47 vdd.t130 vbias2.t35 vsquare.t159 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X48 vsquare.t160 vbias2.t36 vdd.t129 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X49 vsquare.t161 vbias2.t37 vdd.t128 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X50 vss.t137 a_19926_13536.t22 vt.t195 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X51 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X52 vdd.t206 vbias1.t34 a_23370_8306.t28 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X53 vt.t194 a_19926_13536.t23 vss.t136 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X54 vss.t135 a_19926_13536.t24 vt.t193 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X55 vt.t55 vbias1.t35 vdd.t207 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X56 a_23370_24650.t9 vref.t3 a_23744_20184.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X57 a_19926_13536.t6 vref.t4 a_23370_8306.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X58 vss.t134 a_19926_13536.t25 vt.t192 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X59 a_19926_29936.t10 OTA_0/vp a_23370_24650.t34 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X60 vdd.t127 vbias2.t0 vbias2.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X61 vsquare.t162 vbias2.t38 vdd.t126 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X62 vsquare.t163 vbias2.t39 vdd.t125 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X63 vdd.t124 vbias2.t40 vsquare.t164 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X64 vss.t153 a_19926_29936.t26 vsquare.t137 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X65 vsquare.t136 a_19926_29936.t27 vss.t154 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X66 a_23370_24650.t23 vbias2.t41 vdd.t123 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X67 vsquare.t165 vbias2.t42 vdd.t122 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X68 vsquare.t166 vbias2.t43 vdd.t121 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X69 vdd.t120 vbias2.t44 vsquare.t167 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X70 vss.t133 a_19926_13536.t26 vt.t191 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X71 vt.t190 a_19926_13536.t27 vss.t132 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X73 a_23370_24650.t33 OTA_0/vp a_19926_29936.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X74 vsquare.t135 a_19926_29936.t28 vss.t155 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X75 a_23744_3840.t10 OTA_tri_0/vn a_23370_8306.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X77 vss.t131 a_19926_13536.t28 vt.t189 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X78 vsquare.t168 vbias2.t45 vdd.t119 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X79 vdd.t118 vbias2.t46 vsquare.t169 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X80 vbias1.t23 vbias1.t22 vdd.t195 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X81 vt.t56 vbias1.t36 vdd.t208 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X82 vsquare.t170 vbias2.t47 vdd.t117 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X83 vss.t130 a_19926_13536.t29 vt.t188 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X84 vsquare.t134 a_19926_29936.t29 vss.t156 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X85 a_23370_24650.t22 vbias2.t48 vdd.t116 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X86 vss.t129 a_19926_13536.t30 vt.t187 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X87 vsquare.t171 vbias2.t49 vdd.t115 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X88 OTA_0/vp vsquare.t147 vss sky130_fd_pr__res_xhigh_po w=350000u l=9e+06u
X89 vsquare.t172 vbias2.t50 vdd.t114 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X90 vdd.t113 vbias2.t51 vsquare.t173 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X91 vss.t128 a_19926_13536.t31 vt.t186 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X92 a_19926_13536.t13 vref.t5 a_23370_8306.t9 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X93 vsquare.t133 a_19926_29936.t30 vss.t157 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X94 vdd.t112 vbias2.t52 vsquare.t174 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X95 vsquare.t175 vbias2.t53 vdd.t111 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X96 a_19926_13536.t15 a_23744_3840.t20 vss.t62 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X97 vt.t57 vbias1.t37 vdd.t209 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X98 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X99 vsquare.t132 a_19926_29936.t31 vss.t158 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X100 a_23370_8306.t22 OTA_tri_0/vn a_23744_3840.t9 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X101 vsquare.t176 vbias2.t54 vdd.t110 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X102 vss.t127 a_19926_13536.t32 vt.t185 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X103 vdd.t109 vbias2.t55 vsquare.t177 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X104 vt.t58 vbias1.t38 vdd.t210 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X105 vsquare.t131 a_19926_29936.t32 vss.t159 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X106 vsquare.t178 vbias2.t56 vdd.t108 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X107 vss.t126 a_19926_13536.t33 vt.t184 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X108 vsquare.t179 vbias2.t57 vdd.t107 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X109 a_23370_24650.t21 vbias2.t58 vdd.t106 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X110 vdd.t105 vbias2.t59 vsquare.t180 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X111 vdd.t211 vbias1.t39 vt.t59 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X112 vsquare.t181 vbias2.t60 vdd.t104 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X113 vsquare.t130 a_19926_29936.t33 vss.t160 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X114 vt.t60 vbias1.t40 vdd.t212 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X115 a_23370_24650.t32 OTA_0/vp a_19926_29936.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X116 vss.t125 a_19926_13536.t34 vt.t183 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X117 vdd.t103 vbias2.t61 vsquare.t182 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X118 vsquare.t183 vbias2.t62 vdd.t102 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X119 vss.t124 a_19926_13536.t35 vt.t182 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X120 vdd.t213 vbias1.t41 vt.t61 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X121 vsquare.t129 a_19926_29936.t34 vss.t161 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X122 a_23370_24650.t20 vbias2.t63 vdd.t101 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X123 vdd.t214 vbias1.t42 vt.t62 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X124 vdd.t215 vbias1.t43 vt.t63 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X125 vdd.t216 vbias1.t44 vt.t64 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X126 vsquare.t128 a_19926_29936.t35 vss.t162 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X127 vsquare.t184 vbias2.t64 vdd.t100 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X128 a_23370_8306.t8 vref.t6 a_19926_13536.t2 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X129 a_23370_24650.t31 OTA_0/vp a_19926_29936.t8 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X130 vss.t175 a_23744_3840.t21 a_19926_13536.t16 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X131 vsquare.t127 a_19926_29936.t36 vss.t163 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X132 vdd.t217 vbias1.t45 vt.t65 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X133 vsquare.t185 vbias2.t65 vdd.t99 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X134 vdd.t98 vbias2.t66 vsquare.t186 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X135 OTA_tri_0/vn vsquare.t66 vss sky130_fd_pr__res_xhigh_po w=350000u l=1.7e+07u
X136 vt.t66 vbias1.t46 vdd.t218 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X137 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X138 vss.t123 a_19926_13536.t36 vt.t181 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X139 vdd.t97 vbias2.t67 vsquare.t187 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X140 vdd.t219 vbias1.t47 vt.t67 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X141 vt.t68 vbias1.t48 vdd.t220 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X142 vdd.t221 vbias1.t49 vt.t69 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X143 a_19926_29936.t4 a_30831_20339# vss sky130_fd_pr__res_xhigh_po w=350000u l=500000u
X144 a_23370_24650.t19 vbias2.t68 vdd.t96 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X145 vdd.t222 vbias1.t50 vt.t70 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X146 vdd.t223 vbias1.t51 vt.t71 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X147 vt.t72 vbias1.t52 vdd.t224 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X148 vdd.t225 vbias1.t53 vt.t73 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X149 vss.t122 a_19926_13536.t37 vt.t180 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X150 vdd.t226 vbias1.t54 vt.t74 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X151 vt.t179 a_19926_13536.t38 vss.t121 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X152 vss.t120 a_19926_13536.t39 vt.t178 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X153 vsquare.t188 vbias2.t69 vdd.t95 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X154 vsquare.t126 a_19926_29936.t37 vss.t164 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X155 vdd.t94 vbias2.t70 vsquare.t189 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X156 vbias1.t21 vbias1.t20 vdd.t194 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X157 vsquare.t125 a_19926_29936.t38 vss.t165 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X158 vdd.t93 vbias2.t71 vsquare.t190 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X159 vt.t75 vbias1.t55 vdd.t227 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X160 vdd.t228 vbias1.t56 vt.t76 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X161 vss.t119 a_19926_13536.t40 vt.t177 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X163 vsquare.t124 a_19926_29936.t39 vss.t166 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X164 vt.t77 vbias1.t57 vdd.t229 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X165 a_23370_24650.t18 vbias2.t72 vdd.t92 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X166 vt.t176 a_19926_13536.t41 vss.t118 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X167 vdd.t230 vbias1.t58 vt.t78 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X168 vss.t117 a_19926_13536.t42 vt.t175 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X169 vt.t79 vbias1.t59 vdd.t231 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X170 vdd.t232 vbias1.t60 vt.t80 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X171 vdd.t91 vbias2.t73 vsquare.t191 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X172 a_23744_3840.t19 a_23744_3840.t18 vss.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X173 a_23370_8306.t29 vbias1.t61 vdd.t233 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X174 vdd.t234 vbias1.t62 vt.t81 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X175 vsquare.t123 a_19926_29936.t40 vss.t167 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X176 vdd.t90 vbias2.t74 vsquare.t192 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X177 vdd.t235 vbias1.t63 vt.t82 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X178 vt.t174 a_19926_13536.t43 vss.t116 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X179 vdd.t89 vbias2.t75 vsquare.t193 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X180 vsquare.t122 a_19926_29936.t41 vss.t168 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X181 vsquare.t121 a_19926_29936.t42 vss.t169 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X182 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X183 a_23744_3840.t8 OTA_tri_0/vn a_23370_8306.t21 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X184 vdd.t236 vbias1.t64 vt.t83 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X185 vt.t84 vbias1.t65 vdd.t237 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X186 vdd.t88 vbias2.t76 vsquare.t194 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X187 vss.t115 a_19926_13536.t44 vt.t173 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X188 vdd.t238 vbias1.t66 vt.t85 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X189 a_23370_8306.t30 vbias1.t67 vdd.t239 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X190 vt.t172 a_19926_13536.t45 vss.t114 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X191 vdd.t87 vbias2.t77 vsquare.t195 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X192 vsquare.t196 vbias2.t78 vdd.t86 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X193 vdd.t146 vbias1.t68 vt.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X194 a_23370_8306.t7 vref.t7 a_19926_13536.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X196 vsquare.t120 a_19926_29936.t43 vss.t36 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X197 vss.t37 a_19926_29936.t44 vsquare.t119 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X198 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X199 vdd.t247 vbias1.t18 vbias1.t19 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X200 vt.t171 a_19926_13536.t46 vss.t113 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X201 vss.t112 a_19926_13536.t47 vt.t170 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X202 vt.t169 a_19926_13536.t48 vss.t111 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X203 vdd.t85 vbias2.t79 vsquare.t197 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X204 vsquare.t118 a_19926_29936.t45 vss.t38 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X205 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X206 vss.t39 a_19926_29936.t46 vsquare.t117 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X207 a_23744_20184.t9 vref.t8 a_23370_24650.t8 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X208 vsquare.t198 vbias2.t80 vdd.t84 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X209 a_23370_8306.t15 OTA_tri_0/vn a_23744_3840.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X210 vdd.t147 vbias1.t69 vt.t2 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X211 vsquare.t116 a_19926_29936.t47 vss.t40 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X213 vss.t41 a_19926_29936.t48 vsquare.t115 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X214 vdd.t148 vbias1.t70 vt.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X215 vt.t4 vbias1.t71 vdd.t149 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X216 vt.t168 a_19926_13536.t49 vss.t110 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X217 vt.t167 a_19926_13536.t50 vss.t109 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X218 vsquare.t199 vbias2.t81 vdd.t83 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X219 vss.t42 a_19926_29936.t49 vsquare.t114 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X220 vss.t43 a_19926_29936.t50 vsquare.t113 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X221 vsquare.t200 vbias2.t82 vdd.t82 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X222 vbias1.t17 vbias1.t16 vdd.t246 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X223 vdd.t150 vbias1.t72 vt.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X226 vsquare.t201 vbias2.t83 vdd.t81 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X227 vdd.t151 vbias1.t73 vt.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X228 vt.t7 vbias1.t74 vdd.t152 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X229 vss.t44 a_19926_29936.t51 vsquare.t112 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X230 vt.t166 a_19926_13536.t51 vss.t108 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X231 a_19926_13536.t0 vref.t9 a_23370_8306.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X232 a_23744_20184.t5 vref.t10 a_23370_24650.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X233 vt.t165 a_19926_13536.t52 vss.t107 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X234 a_23370_24650.t6 vref.t11 a_23744_20184.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X235 vss.t45 a_19926_29936.t52 vsquare.t111 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X236 a_23744_3840.t6 OTA_tri_0/vn a_23370_8306.t20 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X237 vt.t8 vbias1.t75 vdd.t153 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X238 vt.t9 vbias1.t76 vdd.t154 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X239 vsquare.t0 vbias2.t84 vdd.t80 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X240 vbias1.t15 vbias1.t14 vdd.t245 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X241 vt.t164 a_19926_13536.t53 vss.t106 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X242 vss.t46 a_19926_29936.t53 vsquare.t110 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X243 vdd.t155 vbias1.t77 vt.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X244 vt.t163 a_19926_13536.t54 vss.t105 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X245 a_19926_29936.t1 a_23744_20184.t21 vss.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X246 vsquare.t1 vbias2.t85 vdd.t79 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X247 vss.t47 a_19926_29936.t54 vsquare.t109 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X248 a_23370_8306.t24 vbias1.t78 vdd.t156 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X249 vdd.t157 vbias1.t79 vt.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X250 a_19926_29936.t12 OTA_0/vp a_23370_24650.t30 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X251 vss.t48 a_19926_29936.t55 vsquare.t108 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X252 vsquare.t2 vbias2.t86 vdd.t78 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X253 a_19926_13536.t12 vref.t12 a_23370_8306.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X254 vdd.t77 vbias2.t87 vsquare.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X255 vt.t12 vbias1.t80 vdd.t158 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X256 vdd.t159 vbias1.t81 vt.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X257 vss.t49 a_19926_29936.t56 vsquare.t107 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X258 vt.t162 a_19926_13536.t55 vss.t104 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X259 vt.t14 vbias1.t82 vdd.t160 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X260 vss.t103 a_19926_13536.t56 vt.t161 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X261 vt.t160 a_19926_13536.t57 vss.t102 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X262 vsquare.t4 vbias2.t88 vdd.t76 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X263 a_23744_20184.t17 a_23744_20184.t16 vss.t3 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X264 vss.t50 a_19926_29936.t57 vsquare.t106 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X265 vsquare.t5 vbias2.t89 vdd.t75 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X266 vss.t51 a_19926_29936.t58 vsquare.t105 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X267 vdd.t161 vbias1.t83 vt.t15 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X268 a_23370_8306.t25 vbias1.t84 vdd.t162 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X269 vsquare.t6 vbias2.t90 vdd.t74 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X270 vdd.t163 vbias1.t85 vt.t16 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X271 vbias1.t13 vbias1.t12 vdd.t244 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X273 vdd.t73 vbias2.t91 a_23370_24650.t17 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X274 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X275 vsquare.t7 vbias2.t92 vdd.t72 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X276 a_23370_8306.t23 OTA_tri_0/vn a_23744_3840.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X277 vdd.t164 vbias1.t86 vt.t17 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X278 vt.t159 a_19926_13536.t58 vss.t101 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X279 vss.t52 a_19926_29936.t59 vsquare.t104 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X280 vdd.t71 vbias2.t93 vsquare.t8 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X282 vss.t53 a_19926_29936.t60 vsquare.t103 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X283 vdd.t165 vbias1.t87 vt.t18 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X284 vt.t158 a_19926_13536.t59 vss.t100 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X285 vsquare.t9 vbias2.t94 vdd.t70 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X286 vdd.t166 vbias1.t88 vt.t19 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X287 vbias1.t11 vbias1.t10 vdd.t243 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X288 a_23744_20184.t7 vref.t13 a_23370_24650.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X289 vss.t54 a_19926_29936.t61 vsquare.t102 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X290 vdd.t167 vbias1.t89 vt.t20 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X291 a_23370_8306.t4 vref.t14 a_19926_13536.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X292 a_23744_3840.t17 a_23744_3840.t16 vss.t144 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X293 vt.t157 a_19926_13536.t60 vss.t99 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X294 vdd.t69 vbias2.t95 a_23370_24650.t16 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X295 vsquare.t10 vbias2.t96 vdd.t68 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X296 vdd.t168 vbias1.t90 vt.t21 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X297 vdd.t169 vbias1.t91 vt.t22 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X298 vdd.t170 vbias1.t92 vt.t23 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X299 vt.t24 vbias1.t93 vdd.t171 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X300 vdd.t67 vbias2.t97 a_23370_24650.t15 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X301 vss.t55 a_19926_29936.t62 vsquare.t101 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X302 vdd.t66 vbias2.t98 vsquare.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X304 vsquare.t12 vbias2.t99 vdd.t65 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X305 vss.t98 a_19926_13536.t61 vt.t156 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X306 vt.t25 vbias1.t94 vdd.t172 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X307 vdd.t242 vbias1.t8 vbias1.t9 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X308 vt.t26 vbias1.t95 vdd.t173 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X309 vt.t155 a_19926_13536.t62 vss.t97 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X310 vss.t56 a_19926_29936.t63 vsquare.t100 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X311 a_23370_24650.t29 OTA_0/vp a_19926_29936.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X312 vsquare.t99 a_19926_29936.t64 vss.t57 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X313 vsquare.t13 vbias2.t100 vdd.t64 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X315 vdd.t174 vbias1.t96 vt.t27 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X316 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X317 vdd.t63 vbias2.t101 a_23370_24650.t14 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X318 vdd.t175 vbias1.t97 vt.t28 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X319 vt.t29 vbias1.t98 vdd.t176 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X320 vdd.t177 vbias1.t99 vt.t30 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X321 vdd.t62 vbias2.t102 a_23370_24650.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X322 vsquare a_30831_20339# sky130_fd_pr__cap_mim_m3_1 l=1.35e+07u w=1.35e+07u
X323 vss.t58 a_19926_29936.t65 vsquare.t98 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X324 vdd.t178 vbias1.t100 vt.t31 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X325 vss.t143 a_23744_3840.t14 a_23744_3840.t15 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X326 vt.t32 vbias1.t101 vdd.t179 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X327 vt.t154 a_19926_13536.t63 vss.t96 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X328 vsquare.t14 vbias2.t103 vdd.t61 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X329 vt.t33 vbias1.t102 vdd.t180 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X330 vsquare.t97 a_19926_29936.t66 vss.t59 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X331 vbias2.t13 vbias2.t12 vdd.t60 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X332 vsquare.t15 vbias2.t104 vdd.t59 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X333 vt.t34 vbias1.t103 vdd.t181 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X334 vss.t95 a_19926_13536.t64 vt.t153 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X335 vt.t35 vbias1.t104 vdd.t182 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X336 vt.t36 vbias1.t105 vdd.t183 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X337 vdd.t184 vbias1.t106 vt.t37 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X338 vss.t7 a_23744_20184.t14 a_23744_20184.t15 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X339 vsquare.t96 a_19926_29936.t67 vss.t60 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X340 vss.t11 a_19926_29936.t68 vsquare.t95 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X341 vdd.t58 vbias2.t105 a_23370_24650.t12 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X342 vsquare.t94 a_19926_29936.t69 vss.t12 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X343 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X344 vdd.t185 vbias1.t107 vt.t38 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X345 vsquare.t16 vbias2.t106 vdd.t57 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X346 vt.t39 vbias1.t108 vdd.t186 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X347 vsquare.t17 vbias2.t107 vdd.t56 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X348 a_23744_3840.t4 OTA_tri_0/vn a_23370_8306.t14 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X349 vsquare.t18 vbias2.t108 vdd.t55 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X350 vsquare.t19 vbias2.t109 vdd.t54 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X351 vbias2.t17 vbias2.t16 vdd.t53 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X352 vt.t40 vbias1.t109 vdd.t187 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X353 vt.t41 vbias1.t110 vdd.t188 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X354 vss.t94 a_19926_13536.t65 vt.t152 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X355 vt.t151 a_19926_13536.t66 vss.t93 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X356 a_23370_24650.t28 OTA_0/vp a_19926_29936.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X357 vss.t92 a_19926_13536.t67 vt.t150 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X358 vdd.t189 vbias1.t111 vt.t42 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X359 vss.t0 a_23744_20184.t22 a_19926_29936.t0 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X360 vsquare.t93 a_19926_29936.t70 vss.t13 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X361 vt.t43 vbias1.t112 vdd.t190 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X362 a_23370_8306.t26 vbias1.t113 vdd.t191 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X363 vss.t91 a_19926_13536.t68 vt.t149 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X364 vsquare.t20 vbias2.t110 vdd.t52 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X365 vdd.t192 vbias1.t114 vt.t44 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X366 vt.t45 vbias1.t115 vdd.t193 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X367 vsquare.t92 a_19926_29936.t71 vss.t14 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X368 vsquare.t21 vbias2.t111 vdd.t51 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X369 vbias2.t11 vbias2.t10 vdd.t50 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X370 vsquare.t91 a_19926_29936.t72 vss.t15 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X371 a_23370_24650.t4 vref.t15 a_23744_20184.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X372 vsquare.t22 vbias2.t112 vdd.t49 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X373 vss.t90 a_19926_13536.t69 vt.t148 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X374 vdd.t248 vbias1.t116 vt.t86 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X375 vss.t89 a_19926_13536.t70 vt.t147 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X376 vdd.t48 vbias2.t113 vsquare.t23 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X377 vdd.t47 vbias2.t114 vsquare.t24 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X378 vdd.t249 vbias1.t117 vt.t87 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X379 a_19926_29936.t16 OTA_0/vp a_23370_24650.t27 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X380 vt.t88 vbias1.t118 vdd.t250 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X381 vt.t89 vbias1.t119 vdd.t251 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X382 a_23370_8306.t3 vref.t16 a_19926_13536.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X383 vt.t90 vbias1.t120 vdd.t252 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X384 vdd.t253 vbias1.t121 vt.t91 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X385 vss.t88 a_19926_13536.t71 vt.t146 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X387 vss.t87 a_19926_13536.t72 vt.t145 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X388 vsquare.t25 vbias2.t115 vdd.t46 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X390 vsquare.t90 a_19926_29936.t73 vss.t16 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X391 vsquare.t26 vbias2.t116 vdd.t45 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X392 vss.t86 a_19926_13536.t73 vt.t144 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X393 vdd.t44 vbias2.t117 vsquare.t27 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X394 vdd.t43 vbias2.t118 vsquare.t28 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X395 vdd.t42 vbias2.t119 vsquare.t29 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X396 vdd.t254 vbias1.t122 vt.t92 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X397 vt.t93 vbias1.t123 vdd.t255 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X398 vsquare.t89 a_19926_29936.t74 vss.t17 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X399 vt.t94 vbias1.t124 vdd.t256 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X400 a_23370_8306.t19 OTA_tri_0/vn a_23744_3840.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X401 vsquare.t88 a_19926_29936.t75 vss.t18 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X402 vss.t85 a_19926_13536.t74 vt.t143 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X403 vt.t95 vbias1.t125 vdd.t257 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X404 vdd.t258 vbias1.t126 a_23370_8306.t31 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X405 vss.t84 a_19926_13536.t75 vt.t142 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X406 vbias2.t9 vbias2.t8 vdd.t41 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X407 vss.t83 a_19926_13536.t76 vt.t141 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X408 a_23370_8306.t32 vbias1.t127 vdd.t259 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X409 vss.t82 a_19926_13536.t77 vt.t140 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X410 vt a_30793_4721# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X411 vsquare.t87 a_19926_29936.t76 vss.t19 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X412 vdd.t40 vbias2.t120 vsquare.t30 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X413 vdd.t39 vbias2.t121 vsquare.t31 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X414 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X415 vdd.t38 vbias2.t122 vsquare.t32 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X416 vsquare.t86 a_19926_29936.t77 vss.t20 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X417 vss.t81 a_19926_13536.t78 vt.t139 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X418 vt.t138 a_19926_13536.t79 vss.t80 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X419 vdd.t260 vbias1.t128 a_23370_8306.t33 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X420 vss.t79 a_19926_13536.t80 vt.t137 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X421 vdd.t37 vbias2.t123 vsquare.t33 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X422 vt.t96 vbias1.t129 vdd.t261 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X423 vbias2.t5 vbias2.t4 vdd.t36 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X424 vsquare.t85 a_19926_29936.t78 vss.t21 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X425 vdd.t262 vbias1.t130 vt.t97 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X426 vt.t98 vbias1.t131 vdd.t263 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X427 vt.t99 vbias1.t132 vdd.t264 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X428 vdd.t241 vbias1.t6 vbias1.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X429 vsquare.t84 a_19926_29936.t79 vss.t22 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X430 vss.t78 a_19926_13536.t81 vt.t136 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X431 a_19926_13536.t8 vref.t17 a_23370_8306.t2 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X432 a_23370_24650.t26 OTA_0/vp a_19926_29936.t14 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X433 vdd.t35 vbias2.t124 vsquare.t34 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X434 a_23370_24650.t3 vref.t18 a_23744_20184.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X435 a_23744_3840.t2 OTA_tri_0/vn a_23370_8306.t18 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X436 vdd.t34 vbias2.t125 vsquare.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X437 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X438 vdd.t265 vbias1.t133 vt.t100 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X439 vss.t77 a_19926_13536.t82 vt.t135 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X440 vsquare.t83 a_19926_29936.t80 vss.t23 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X441 vss.t24 a_19926_29936.t81 vsquare.t82 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X442 vbias2.t15 vbias2.t14 vdd.t33 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X443 vdd.t32 vbias2.t126 vsquare.t36 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X444 vsquare.t81 a_19926_29936.t82 vss.t25 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X445 a_19926_29936.t15 OTA_0/vp a_23370_24650.t25 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X446 vt.t101 vbias1.t134 vdd.t266 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X447 vdd.t240 vbias1.t4 vbias1.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X448 vdd.t31 vbias2.t127 vsquare.t37 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X449 vt.t102 vbias1.t135 vdd.t267 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X450 a_19926_13536.t14 vref.t19 a_23370_8306.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X451 vt.t134 a_19926_13536.t83 vss.t76 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X452 vt.t103 vbias1.t136 vdd.t268 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X453 vdd.t269 vbias1.t137 a_23370_8306.t34 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X454 vdd.t30 vbias2.t128 vsquare.t38 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X456 vdd.t29 vbias2.t2 vbias2.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X457 vdd.t270 vbias1.t138 vt.t104 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X458 vsquare.t80 a_19926_29936.t83 vss.t26 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X459 a_23370_8306.t16 OTA_tri_0/vn a_23744_3840.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X460 a_19926_13536.t3 a_30793_4721# vss sky130_fd_pr__res_xhigh_po w=350000u l=2.8e+06u
X461 vdd.t28 vbias2.t129 vsquare.t39 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X462 vsquare.t79 a_19926_29936.t84 vss.t27 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X463 vss.t4 a_23744_3840.t12 a_23744_3840.t13 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X464 vt.t133 a_19926_13536.t84 vss.t75 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X465 vdd.t27 vbias2.t130 vsquare.t40 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X466 vdd.t26 vbias2.t131 vsquare.t41 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X467 vss.t74 a_19926_13536.t85 vt.t132 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X468 vt.t131 a_19926_13536.t86 vss.t73 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X470 vt.t105 vbias1.t139 vdd.t271 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X471 vdd.t272 vbias1.t140 a_23370_8306.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X472 vsquare.t78 a_19926_29936.t85 vss.t28 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X473 vdd.t25 vbias2.t6 vbias2.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X474 vdd.t24 vbias2.t132 vsquare.t42 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X475 a_23370_24650.t2 vref.t20 a_23744_20184.t2 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X476 vsquare.t43 vbias2.t133 vdd.t23 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X477 vdd.t22 vbias2.t134 vsquare.t44 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X478 vdd.t273 vbias1.t141 vt.t106 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X479 vt.t130 a_19926_13536.t87 vss.t72 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X480 a_19926_29936.t3 a_23744_20184.t23 vss.t61 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X481 vss.t29 a_19926_29936.t86 vsquare.t77 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X482 vt.t107 vbias1.t142 vdd.t274 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X483 vt.t129 a_19926_13536.t88 vss.t71 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X484 a_23744_20184.t4 vref.t21 a_23370_24650.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X485 vdd.t21 vbias2.t135 vsquare.t45 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X486 a_23370_8306.t0 vref.t22 a_19926_13536.t9 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X487 vdd.t20 vbias2.t136 vsquare.t46 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X488 a_19926_29936.t7 OTA_0/vp a_23370_24650.t24 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X489 vt.t0 OTA_0/vp vss sky130_fd_pr__res_xhigh_po w=350000u l=4e+06u
X490 vdd.t19 vbias2.t18 vbias2.t19 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X491 vt.t128 a_19926_13536.t89 vss.t70 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X492 vsquare.t47 vbias2.t137 vdd.t18 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X493 vdd.t275 vbias1.t143 vt.t108 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X494 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X495 a_23744_20184.t13 a_23744_20184.t12 vss.t1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X496 vdd.t17 vbias2.t138 vsquare.t48 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X497 vsquare.t49 vbias2.t139 vdd.t16 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X498 vdd.t15 vbias2.t140 vsquare.t50 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X499 vt.t127 a_19926_13536.t90 vss.t69 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X500 vt.t109 vbias1.t144 vdd.t276 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X501 vsquare.t76 a_19926_29936.t87 vss.t30 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X502 vss.t31 a_19926_29936.t88 vsquare.t75 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X503 a_19926_13536.t1 a_23744_3840.t22 vss.t2 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X504 vsquare.t51 vbias2.t141 vdd.t14 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X505 vt.t126 a_19926_13536.t91 vss.t68 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X507 vdd.t13 vbias2.t142 vsquare.t52 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X508 vss.t32 a_19926_29936.t89 vsquare.t74 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X509 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X510 vt.t125 a_19926_13536.t92 vss.t67 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X512 vsquare.t53 vbias2.t143 vdd.t12 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X513 vt OTA_tri_0/vn sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X514 vdd.t11 vbias2.t144 vsquare.t54 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X515 vsquare.t55 vbias2.t145 vdd.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X516 vdd.t9 vbias2.t146 vsquare.t56 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X517 vss.t33 a_19926_29936.t90 vsquare.t73 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X518 vt.t110 vbias1.t145 vdd.t277 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X519 vt.t111 vbias1.t146 vdd.t278 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X520 vdd.t144 vbias1.t2 vbias1.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X521 vt.t124 a_19926_13536.t93 vss.t66 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X522 vsquare.t57 vbias2.t147 vdd.t8 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X523 vt.t123 a_19926_13536.t94 vss.t65 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X524 vsquare.t58 vbias2.t148 vdd.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X525 vdd.t6 vbias2.t149 vsquare.t59 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X526 vt.t112 vbias1.t147 vdd.t279 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X527 a_23744_20184.t3 vref.t23 a_23370_24650.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X528 vss.t34 a_19926_29936.t91 vsquare.t72 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X529 vdd.t280 vbias1.t148 vt.t113 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X530 vt.t114 vbias1.t149 vdd.t281 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X531 vss.t35 a_19926_29936.t92 vsquare.t71 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X532 vt.t115 vbias1.t150 vdd.t282 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X533 vt.t122 a_19926_13536.t95 vss.t64 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X534 vdd.t5 vbias2.t150 vsquare.t60 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X535 vsquare.t61 vbias2.t151 vdd.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X536 vss.t171 a_19926_29936.t93 vsquare.t70 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X537 a_23744_3840.t0 OTA_tri_0/vn a_23370_8306.t17 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X538 vt.t116 vbias1.t151 vdd.t283 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X539 vss.t10 a_23744_3840.t23 a_19926_13536.t10 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X540 vss.t172 a_19926_29936.t94 vsquare.t69 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X541 vdd.t145 vbias1.t0 vbias1.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X542 vt.t117 vbias1.t152 vdd.t284 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X543 vsquare.t62 vbias2.t152 vdd.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X544 vsquare.t63 vbias2.t153 vdd.t2 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X545 vdd.t1 vbias2.t154 vsquare.t64 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X546 vt.t118 vbias1.t153 vdd.t285 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X547 vss.t173 a_19926_29936.t95 vsquare.t68 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X548 vt.t119 vbias1.t154 vdd.t286 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X549 vdd.t0 vbias2.t155 vsquare.t65 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X550 vdd.t287 vbias1.t155 vt.t120 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X551 vss.t174 a_19926_29936.t96 vsquare.t67 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
X552 vt.t121 a_19926_13536.t96 vss.t63 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=350000u
C0 OTA_0/vp vref 3.40fF
C1 OTA_tri_0/vn vt 362.14fF
C2 vsquare vbias2 45.21fF
C3 vt a_30793_4721# 22.30fF
C4 vref vt 2.50fF
C5 vsquare OTA_0/vp 2.21fF
C6 vdd vbias1 72.50fF
C7 vsquare a_30831_20339# 18.79fF
C8 vdd vbias2 68.14fF
C9 vdd OTA_tri_0/vn 1.14fF
C10 vdd vref 2.82fF
C11 vdd OTA_0/vp 1.23fF
C12 vdd vt 18.79fF
C13 OTA_tri_0/vn vref 3.40fF
C14 vdd vsquare 18.69fF
C15 vt vbias1 48.47fF
R0 a_19926_13536.n9 a_19926_13536.t29 278.38
R1 a_19926_13536.n9 a_19926_13536.t43 278.184
R2 a_19926_13536.n6 a_19926_13536.t59 278.184
R3 a_19926_13536.n9 a_19926_13536.t45 278.183
R4 a_19926_13536.n9 a_19926_13536.t38 278.183
R5 a_19926_13536.n8 a_19926_13536.t41 278.183
R6 a_19926_13536.n8 a_19926_13536.t87 278.183
R7 a_19926_13536.n8 a_19926_13536.t89 278.183
R8 a_19926_13536.n8 a_19926_13536.t83 278.183
R9 a_19926_13536.n7 a_19926_13536.t84 278.183
R10 a_19926_13536.n7 a_19926_13536.t79 278.183
R11 a_19926_13536.n7 a_19926_13536.t53 278.183
R12 a_19926_13536.n7 a_19926_13536.t55 278.183
R13 a_19926_13536.n5 a_19926_13536.t49 278.183
R14 a_19926_13536.n5 a_19926_13536.t51 278.183
R15 a_19926_13536.n5 a_19926_13536.t46 278.183
R16 a_19926_13536.n5 a_19926_13536.t19 278.183
R17 a_19926_13536.n6 a_19926_13536.t95 278.183
R18 a_19926_13536.n6 a_19926_13536.t96 278.183
R19 a_19926_13536.n6 a_19926_13536.t91 278.183
R20 a_19926_13536.n6 a_19926_13536.t93 278.183
R21 a_19926_13536.n14 a_19926_13536.t90 278.182
R22 a_19926_13536.n9 a_19926_13536.t56 278.182
R23 a_19926_13536.n14 a_19926_13536.t24 278.182
R24 a_19926_13536.n14 a_19926_13536.t92 278.182
R25 a_19926_13536.n9 a_19926_13536.t33 278.182
R26 a_19926_13536.n14 a_19926_13536.t81 278.182
R27 a_19926_13536.n14 a_19926_13536.t86 278.182
R28 a_19926_13536.n8 a_19926_13536.t25 278.182
R29 a_19926_13536.n13 a_19926_13536.t72 278.182
R30 a_19926_13536.n13 a_19926_13536.t88 278.182
R31 a_19926_13536.n8 a_19926_13536.t28 278.182
R32 a_19926_13536.n13 a_19926_13536.t74 278.182
R33 a_19926_13536.n13 a_19926_13536.t54 278.182
R34 a_19926_13536.n8 a_19926_13536.t20 278.182
R35 a_19926_13536.n13 a_19926_13536.t67 278.182
R36 a_19926_13536.n13 a_19926_13536.t57 278.182
R37 a_19926_13536.n8 a_19926_13536.t22 278.182
R38 a_19926_13536.n13 a_19926_13536.t69 278.182
R39 a_19926_13536.n13 a_19926_13536.t50 278.182
R40 a_19926_13536.n7 a_19926_13536.t68 278.182
R41 a_19926_13536.n12 a_19926_13536.t39 278.182
R42 a_19926_13536.n12 a_19926_13536.t52 278.182
R43 a_19926_13536.n7 a_19926_13536.t71 278.182
R44 a_19926_13536.n12 a_19926_13536.t42 278.182
R45 a_19926_13536.n12 a_19926_13536.t48 278.182
R46 a_19926_13536.n7 a_19926_13536.t64 278.182
R47 a_19926_13536.n12 a_19926_13536.t35 278.182
R48 a_19926_13536.n12 a_19926_13536.t21 278.182
R49 a_19926_13536.n7 a_19926_13536.t65 278.182
R50 a_19926_13536.n12 a_19926_13536.t36 278.182
R51 a_19926_13536.n12 a_19926_13536.t23 278.182
R52 a_19926_13536.n5 a_19926_13536.t61 278.182
R53 a_19926_13536.n10 a_19926_13536.t31 278.182
R54 a_19926_13536.n10 a_19926_13536.t17 278.182
R55 a_19926_13536.n5 a_19926_13536.t37 278.182
R56 a_19926_13536.n10 a_19926_13536.t85 278.182
R57 a_19926_13536.n10 a_19926_13536.t18 278.182
R58 a_19926_13536.n5 a_19926_13536.t32 278.182
R59 a_19926_13536.n10 a_19926_13536.t80 278.182
R60 a_19926_13536.n10 a_19926_13536.t94 278.182
R61 a_19926_13536.n5 a_19926_13536.t34 278.182
R62 a_19926_13536.n10 a_19926_13536.t82 278.182
R63 a_19926_13536.n10 a_19926_13536.t66 278.182
R64 a_19926_13536.n6 a_19926_13536.t26 278.182
R65 a_19926_13536.n11 a_19926_13536.t73 278.182
R66 a_19926_13536.n11 a_19926_13536.t62 278.182
R67 a_19926_13536.n6 a_19926_13536.t30 278.182
R68 a_19926_13536.n11 a_19926_13536.t77 278.182
R69 a_19926_13536.n11 a_19926_13536.t63 278.182
R70 a_19926_13536.n6 a_19926_13536.t75 278.182
R71 a_19926_13536.n11 a_19926_13536.t44 278.182
R72 a_19926_13536.n11 a_19926_13536.t58 278.182
R73 a_19926_13536.n6 a_19926_13536.t78 278.182
R74 a_19926_13536.n11 a_19926_13536.t47 278.182
R75 a_19926_13536.n11 a_19926_13536.t60 278.182
R76 a_19926_13536.n6 a_19926_13536.t70 278.182
R77 a_19926_13536.n11 a_19926_13536.t40 278.182
R78 a_19926_13536.n11 a_19926_13536.t27 278.182
R79 a_19926_13536.n14 a_19926_13536.t76 278.182
R80 a_19926_13536.n17 a_19926_13536.t3 153.424
R81 a_19926_13536.n4 a_19926_13536.t9 7.146
R82 a_19926_13536.n3 a_19926_13536.t6 7.146
R83 a_19926_13536.n3 a_19926_13536.t7 7.146
R84 a_19926_13536.n4 a_19926_13536.t8 7.146
R85 a_19926_13536.n4 a_19926_13536.t2 7.146
R86 a_19926_13536.n2 a_19926_13536.t13 7.146
R87 a_19926_13536.n2 a_19926_13536.t5 7.146
R88 a_19926_13536.n2 a_19926_13536.t14 7.146
R89 a_19926_13536.n2 a_19926_13536.t11 7.146
R90 a_19926_13536.n1 a_19926_13536.t12 7.146
R91 a_19926_13536.n1 a_19926_13536.t4 7.146
R92 a_19926_13536.t0 a_19926_13536.n4 7.146
R93 a_19926_13536.n0 a_19926_13536.t16 5.807
R94 a_19926_13536.n0 a_19926_13536.t15 5.807
R95 a_19926_13536.n0 a_19926_13536.t10 5.807
R96 a_19926_13536.n0 a_19926_13536.t1 5.807
R97 a_19926_13536.n16 a_19926_13536.n17 4.373
R98 a_19926_13536.n16 a_19926_13536.n0 2.553
R99 a_19926_13536.n15 a_19926_13536.n11 2.073
R100 a_19926_13536.n15 a_19926_13536.n6 1.962
R101 a_19926_13536.n4 a_19926_13536.n3 1.654
R102 a_19926_13536.n2 a_19926_13536.n1 1.654
R103 a_19926_13536.n7 a_19926_13536.n8 1.571
R104 a_19926_13536.n5 a_19926_13536.n7 1.571
R105 a_19926_13536.n6 a_19926_13536.n5 1.571
R106 a_19926_13536.n12 a_19926_13536.n13 1.566
R107 a_19926_13536.n10 a_19926_13536.n12 1.566
R108 a_19926_13536.n11 a_19926_13536.n10 1.566
R109 a_19926_13536.n13 a_19926_13536.n14 1.566
R110 a_19926_13536.n17 a_19926_13536.n15 1.489
R111 a_19926_13536.n8 a_19926_13536.n9 1.375
R112 a_19926_13536.n4 a_19926_13536.n16 1.314
R113 a_19926_13536.n16 a_19926_13536.n2 1.313
R114 vss.n292 vss.n219 5703.2
R115 vss.n292 vss.n291 1390.68
R116 vss.n267 vss.n266 1390.68
R117 vss.n265 vss.n264 1390.68
R118 vss.n240 vss.n219 1390.68
R119 vss.n291 vss.n290 1390.59
R120 vss.n290 vss.n220 1390.59
R121 vss.n286 vss.n220 1390.59
R122 vss.n286 vss.n285 1390.59
R123 vss.n285 vss.n284 1390.59
R124 vss.n284 vss.n222 1390.59
R125 vss.n280 vss.n222 1390.59
R126 vss.n280 vss.n279 1390.59
R127 vss.n279 vss.n278 1390.59
R128 vss.n278 vss.n224 1390.59
R129 vss.n274 vss.n224 1390.59
R130 vss.n274 vss.n273 1390.59
R131 vss.n273 vss.n272 1390.59
R132 vss.n272 vss.n226 1390.59
R133 vss.n268 vss.n226 1390.59
R134 vss.n268 vss.n267 1390.59
R135 vss.n264 vss.n230 1390.59
R136 vss.n260 vss.n230 1390.59
R137 vss.n260 vss.n259 1390.59
R138 vss.n259 vss.n258 1390.59
R139 vss.n258 vss.n232 1390.59
R140 vss.n254 vss.n232 1390.59
R141 vss.n254 vss.n253 1390.59
R142 vss.n253 vss.n252 1390.59
R143 vss.n252 vss.n234 1390.59
R144 vss.n248 vss.n234 1390.59
R145 vss.n248 vss.n247 1390.59
R146 vss.n247 vss.n246 1390.59
R147 vss.n246 vss.n236 1390.59
R148 vss.n242 vss.n236 1390.59
R149 vss.n242 vss.n241 1390.59
R150 vss.n241 vss.n240 1390.59
R151 vss.n266 vss.n265 143.577
R152 vss.n132 vss.n130 75.701
R153 vss.n125 vss.n123 75.701
R154 vss.n118 vss.n116 75.701
R155 vss.n111 vss.n109 75.701
R156 vss.n104 vss.n102 75.701
R157 vss.n97 vss.n95 75.701
R158 vss.n90 vss.n88 75.701
R159 vss.n83 vss.n81 75.701
R160 vss.n76 vss.n74 75.701
R161 vss.n59 vss.n57 75.701
R162 vss.n52 vss.n50 75.701
R163 vss.n45 vss.n43 75.701
R164 vss.n38 vss.n36 75.701
R165 vss.n31 vss.n29 75.701
R166 vss.n24 vss.n22 75.701
R167 vss.n17 vss.n15 75.701
R168 vss.n10 vss.n8 75.701
R169 vss.n158 vss.n1 75.701
R170 vss.n293 vss.n218 75.701
R171 vss.n289 vss.n218 75.701
R172 vss.n289 vss.n288 75.701
R173 vss.n288 vss.n287 75.701
R174 vss.n287 vss.n221 75.701
R175 vss.n283 vss.n221 75.701
R176 vss.n283 vss.n282 75.701
R177 vss.n282 vss.n281 75.701
R178 vss.n281 vss.n223 75.701
R179 vss.n277 vss.n223 75.701
R180 vss.n277 vss.n276 75.701
R181 vss.n276 vss.n275 75.701
R182 vss.n275 vss.n225 75.701
R183 vss.n271 vss.n225 75.701
R184 vss.n271 vss.n270 75.701
R185 vss.n270 vss.n269 75.701
R186 vss.n269 vss.n227 75.701
R187 vss.n228 vss.n227 75.701
R188 vss.n263 vss.n229 75.701
R189 vss.n263 vss.n262 75.701
R190 vss.n262 vss.n261 75.701
R191 vss.n261 vss.n231 75.701
R192 vss.n257 vss.n231 75.701
R193 vss.n257 vss.n256 75.701
R194 vss.n256 vss.n255 75.701
R195 vss.n255 vss.n233 75.701
R196 vss.n251 vss.n233 75.701
R197 vss.n251 vss.n250 75.701
R198 vss.n250 vss.n249 75.701
R199 vss.n249 vss.n235 75.701
R200 vss.n245 vss.n235 75.701
R201 vss.n245 vss.n244 75.701
R202 vss.n244 vss.n243 75.701
R203 vss.n243 vss.n237 75.701
R204 vss.n239 vss.n237 75.701
R205 vss.n239 vss.n238 75.701
R206 vss.n6 vss.t67 5.807
R207 vss.n6 vss.t135 5.807
R208 vss.n5 vss.t114 5.807
R209 vss.n5 vss.t103 5.807
R210 vss.n13 vss.t73 5.807
R211 vss.n13 vss.t78 5.807
R212 vss.n12 vss.t121 5.807
R213 vss.n12 vss.t126 5.807
R214 vss.n20 vss.t71 5.807
R215 vss.n20 vss.t87 5.807
R216 vss.n19 vss.t118 5.807
R217 vss.n19 vss.t134 5.807
R218 vss.n27 vss.t105 5.807
R219 vss.n27 vss.t85 5.807
R220 vss.n26 vss.t72 5.807
R221 vss.n26 vss.t131 5.807
R222 vss.n34 vss.t102 5.807
R223 vss.n34 vss.t92 5.807
R224 vss.n33 vss.t70 5.807
R225 vss.n33 vss.t139 5.807
R226 vss.n41 vss.t109 5.807
R227 vss.n41 vss.t90 5.807
R228 vss.n40 vss.t76 5.807
R229 vss.n40 vss.t137 5.807
R230 vss.n48 vss.t107 5.807
R231 vss.n48 vss.t120 5.807
R232 vss.n47 vss.t75 5.807
R233 vss.n47 vss.t91 5.807
R234 vss.n55 vss.t111 5.807
R235 vss.n55 vss.t117 5.807
R236 vss.n54 vss.t80 5.807
R237 vss.n54 vss.t88 5.807
R238 vss.n62 vss.t138 5.807
R239 vss.n62 vss.t124 5.807
R240 vss.n61 vss.t106 5.807
R241 vss.n61 vss.t95 5.807
R242 vss.n72 vss.t136 5.807
R243 vss.n72 vss.t123 5.807
R244 vss.n71 vss.t104 5.807
R245 vss.n71 vss.t94 5.807
R246 vss.n79 vss.t142 5.807
R247 vss.n79 vss.t128 5.807
R248 vss.n78 vss.t110 5.807
R249 vss.n78 vss.t98 5.807
R250 vss.n86 vss.t141 5.807
R251 vss.n86 vss.t74 5.807
R252 vss.n85 vss.t108 5.807
R253 vss.n85 vss.t122 5.807
R254 vss.n93 vss.t65 5.807
R255 vss.n93 vss.t79 5.807
R256 vss.n92 vss.t113 5.807
R257 vss.n92 vss.t127 5.807
R258 vss.n100 vss.t93 5.807
R259 vss.n100 vss.t77 5.807
R260 vss.n99 vss.t140 5.807
R261 vss.n99 vss.t125 5.807
R262 vss.n107 vss.t97 5.807
R263 vss.n107 vss.t86 5.807
R264 vss.n106 vss.t64 5.807
R265 vss.n106 vss.t133 5.807
R266 vss.n114 vss.t96 5.807
R267 vss.n114 vss.t82 5.807
R268 vss.n113 vss.t63 5.807
R269 vss.n113 vss.t129 5.807
R270 vss.n121 vss.t101 5.807
R271 vss.n121 vss.t115 5.807
R272 vss.n120 vss.t68 5.807
R273 vss.n120 vss.t84 5.807
R274 vss.n128 vss.t99 5.807
R275 vss.n128 vss.t112 5.807
R276 vss.n127 vss.t66 5.807
R277 vss.n127 vss.t81 5.807
R278 vss.n137 vss.t132 5.807
R279 vss.n137 vss.t119 5.807
R280 vss.n136 vss.t100 5.807
R281 vss.n136 vss.t89 5.807
R282 vss.n4 vss.t69 5.807
R283 vss.n4 vss.t83 5.807
R284 vss.n3 vss.t116 5.807
R285 vss.n3 vss.t130 5.807
R286 vss.n69 vss.t8 5.807
R287 vss.n69 vss.t1 5.807
R288 vss.n68 vss.t0 5.807
R289 vss.n68 vss.t3 5.807
R290 vss.n67 vss.t9 5.807
R291 vss.n67 vss.t61 5.807
R292 vss.n66 vss.t7 5.807
R293 vss.n66 vss.t5 5.807
R294 vss.n160 vss.t158 5.807
R295 vss.n160 vss.t170 5.807
R296 vss.n159 vss.t60 5.807
R297 vss.n159 vss.t46 5.807
R298 vss.n163 vss.t160 5.807
R299 vss.n163 vss.t37 5.807
R300 vss.n162 vss.t13 5.807
R301 vss.n162 vss.t24 5.807
R302 vss.n166 vss.t154 5.807
R303 vss.n166 vss.t148 5.807
R304 vss.n165 vss.t57 5.807
R305 vss.n165 vss.t50 5.807
R306 vss.n169 vss.t156 5.807
R307 vss.n169 vss.t35 5.807
R308 vss.n168 vss.t59 5.807
R309 vss.n168 vss.t42 5.807
R310 vss.n172 vss.t18 5.807
R311 vss.n172 vss.t173 5.807
R312 vss.n171 vss.t159 5.807
R313 vss.n171 vss.t45 5.807
R314 vss.n175 vss.t20 5.807
R315 vss.n175 vss.t31 5.807
R316 vss.n174 vss.t161 5.807
R317 vss.n174 vss.t39 5.807
R318 vss.n178 vss.t15 5.807
R319 vss.n178 vss.t33 5.807
R320 vss.n177 vss.t155 5.807
R321 vss.n177 vss.t41 5.807
R322 vss.n181 vss.t16 5.807
R323 vss.n181 vss.t53 5.807
R324 vss.n180 vss.t157 5.807
R325 vss.n180 vss.t171 5.807
R326 vss.n184 vss.t12 5.807
R327 vss.n184 vss.t55 5.807
R328 vss.n183 vss.t152 5.807
R329 vss.n183 vss.t145 5.807
R330 vss.n187 vss.t169 5.807
R331 vss.n187 vss.t48 5.807
R332 vss.n186 vss.t21 5.807
R333 vss.n186 vss.t32 5.807
R334 vss.n190 vss.t36 5.807
R335 vss.n190 vss.t51 5.807
R336 vss.n189 vss.t23 5.807
R337 vss.n189 vss.t34 5.807
R338 vss.n193 vss.t165 5.807
R339 vss.n193 vss.t43 5.807
R340 vss.n192 vss.t17 5.807
R341 vss.n192 vss.t29 5.807
R342 vss.n196 vss.t167 5.807
R343 vss.n196 vss.t153 5.807
R344 vss.n195 vss.t19 5.807
R345 vss.n195 vss.t56 5.807
R346 vss.n199 vss.t162 5.807
R347 vss.n199 vss.t147 5.807
R348 vss.n198 vss.t14 5.807
R349 vss.n198 vss.t49 5.807
R350 vss.n202 vss.t30 5.807
R351 vss.n202 vss.t150 5.807
R352 vss.n201 vss.t38 5.807
R353 vss.n201 vss.t52 5.807
R354 vss.n205 vss.t26 5.807
R355 vss.n205 vss.t172 5.807
R356 vss.n204 vss.t166 5.807
R357 vss.n204 vss.t44 5.807
R358 vss.n208 vss.t28 5.807
R359 vss.n208 vss.t146 5.807
R360 vss.n207 vss.t168 5.807
R361 vss.n207 vss.t47 5.807
R362 vss.n211 vss.t22 5.807
R363 vss.n211 vss.t58 5.807
R364 vss.n210 vss.t163 5.807
R365 vss.n210 vss.t149 5.807
R366 vss.n214 vss.t25 5.807
R367 vss.n214 vss.t11 5.807
R368 vss.n213 vss.t164 5.807
R369 vss.n213 vss.t151 5.807
R370 vss.n217 vss.t40 5.807
R371 vss.n217 vss.t54 5.807
R372 vss.n216 vss.t27 5.807
R373 vss.n216 vss.t174 5.807
R374 vss.n316 vss.t10 5.807
R375 vss.n316 vss.t6 5.807
R376 vss.n315 vss.t175 5.807
R377 vss.n315 vss.t144 5.807
R378 vss.n314 vss.t143 5.807
R379 vss.n314 vss.t2 5.807
R380 vss.n313 vss.t4 5.807
R381 vss.n313 vss.t62 5.807
R382 vss.n70 vss.n69 1.455
R383 vss.n317 vss.n316 1.455
R384 vss.n70 vss.n67 1.429
R385 vss.n317 vss.n314 1.429
R386 vss.n138 vss.n137 1.271
R387 vss.n164 vss.n163 1.271
R388 vss.n170 vss.n169 1.271
R389 vss.n176 vss.n175 1.271
R390 vss.n182 vss.n181 1.271
R391 vss.n188 vss.n187 1.271
R392 vss.n194 vss.n193 1.271
R393 vss.n200 vss.n199 1.271
R394 vss.n206 vss.n205 1.271
R395 vss.n212 vss.n211 1.271
R396 vss.n133 vss.n128 1.271
R397 vss.n126 vss.n121 1.271
R398 vss.n119 vss.n114 1.271
R399 vss.n112 vss.n107 1.271
R400 vss.n105 vss.n100 1.271
R401 vss.n98 vss.n93 1.271
R402 vss.n91 vss.n86 1.271
R403 vss.n84 vss.n79 1.271
R404 vss.n77 vss.n72 1.271
R405 vss.n65 vss.n62 1.271
R406 vss.n60 vss.n55 1.271
R407 vss.n53 vss.n48 1.271
R408 vss.n46 vss.n41 1.271
R409 vss.n39 vss.n34 1.271
R410 vss.n32 vss.n27 1.271
R411 vss.n25 vss.n20 1.271
R412 vss.n18 vss.n13 1.271
R413 vss.n11 vss.n6 1.271
R414 vss.n215 vss.n214 1.271
R415 vss.n209 vss.n208 1.271
R416 vss.n203 vss.n202 1.271
R417 vss.n197 vss.n196 1.271
R418 vss.n191 vss.n190 1.271
R419 vss.n185 vss.n184 1.271
R420 vss.n179 vss.n178 1.271
R421 vss.n173 vss.n172 1.271
R422 vss.n167 vss.n166 1.271
R423 vss.n161 vss.n160 1.271
R424 vss.n158 vss.n4 1.27
R425 vss.n293 vss.n217 1.27
R426 vss.n318 vss.n312 0.906
R427 vss.n6 vss.n5 0.867
R428 vss.n13 vss.n12 0.867
R429 vss.n20 vss.n19 0.867
R430 vss.n27 vss.n26 0.867
R431 vss.n34 vss.n33 0.867
R432 vss.n41 vss.n40 0.867
R433 vss.n48 vss.n47 0.867
R434 vss.n55 vss.n54 0.867
R435 vss.n62 vss.n61 0.867
R436 vss.n72 vss.n71 0.867
R437 vss.n79 vss.n78 0.867
R438 vss.n86 vss.n85 0.867
R439 vss.n93 vss.n92 0.867
R440 vss.n100 vss.n99 0.867
R441 vss.n107 vss.n106 0.867
R442 vss.n114 vss.n113 0.867
R443 vss.n121 vss.n120 0.867
R444 vss.n128 vss.n127 0.867
R445 vss.n137 vss.n136 0.867
R446 vss.n4 vss.n3 0.867
R447 vss.n69 vss.n68 0.867
R448 vss.n67 vss.n66 0.867
R449 vss.n160 vss.n159 0.867
R450 vss.n163 vss.n162 0.867
R451 vss.n166 vss.n165 0.867
R452 vss.n169 vss.n168 0.867
R453 vss.n172 vss.n171 0.867
R454 vss.n175 vss.n174 0.867
R455 vss.n178 vss.n177 0.867
R456 vss.n181 vss.n180 0.867
R457 vss.n184 vss.n183 0.867
R458 vss.n187 vss.n186 0.867
R459 vss.n190 vss.n189 0.867
R460 vss.n193 vss.n192 0.867
R461 vss.n196 vss.n195 0.867
R462 vss.n199 vss.n198 0.867
R463 vss.n202 vss.n201 0.867
R464 vss.n205 vss.n204 0.867
R465 vss.n208 vss.n207 0.867
R466 vss.n211 vss.n210 0.867
R467 vss.n214 vss.n213 0.867
R468 vss.n217 vss.n216 0.867
R469 vss.n316 vss.n315 0.867
R470 vss.n314 vss.n313 0.867
R471 vss.n318 vss 0.545
R472 vss vss.n317 0.46
R473 vss vss.n158 0.174
R474 vss.n132 vss.n131 0.092
R475 vss.n125 vss.n124 0.092
R476 vss.n118 vss.n117 0.092
R477 vss.n111 vss.n110 0.092
R478 vss.n104 vss.n103 0.092
R479 vss.n97 vss.n96 0.092
R480 vss.n90 vss.n89 0.092
R481 vss.n83 vss.n82 0.092
R482 vss.n59 vss.n58 0.092
R483 vss.n52 vss.n51 0.092
R484 vss.n45 vss.n44 0.092
R485 vss.n38 vss.n37 0.092
R486 vss.n31 vss.n30 0.092
R487 vss.n24 vss.n23 0.092
R488 vss.n17 vss.n16 0.092
R489 vss.n10 vss.n9 0.092
R490 vss.n290 vss.n289 0.092
R491 vss.n287 vss.n286 0.092
R492 vss.n284 vss.n283 0.092
R493 vss.n281 vss.n280 0.092
R494 vss.n278 vss.n277 0.092
R495 vss.n275 vss.n274 0.092
R496 vss.n272 vss.n271 0.092
R497 vss.n269 vss.n268 0.092
R498 vss.n262 vss.n230 0.092
R499 vss.n259 vss.n231 0.092
R500 vss.n256 vss.n232 0.092
R501 vss.n253 vss.n233 0.092
R502 vss.n250 vss.n234 0.092
R503 vss.n247 vss.n235 0.092
R504 vss.n244 vss.n236 0.092
R505 vss.n241 vss.n237 0.092
R506 vss.n294 vss.n293 0.017
R507 vss.n295 vss.n294 0.017
R508 vss.n296 vss.n295 0.017
R509 vss.n297 vss.n296 0.017
R510 vss.n298 vss.n297 0.017
R511 vss.n299 vss.n298 0.017
R512 vss.n300 vss.n299 0.017
R513 vss.n301 vss.n300 0.017
R514 vss.n302 vss.n301 0.017
R515 vss.n303 vss.n302 0.017
R516 vss.n304 vss.n303 0.017
R517 vss.n305 vss.n304 0.017
R518 vss.n306 vss.n305 0.017
R519 vss.n307 vss.n306 0.017
R520 vss.n308 vss.n307 0.017
R521 vss.n309 vss.n308 0.017
R522 vss.n310 vss.n309 0.017
R523 vss.n311 vss.n310 0.017
R524 vss.n312 vss.n311 0.017
R525 vss vss.n318 0.011
R526 vss.n139 vss.n138 0.009
R527 vss.n140 vss.n139 0.008
R528 vss.n141 vss.n140 0.008
R529 vss.n142 vss.n141 0.008
R530 vss.n143 vss.n142 0.008
R531 vss.n144 vss.n143 0.008
R532 vss.n145 vss.n144 0.008
R533 vss.n146 vss.n145 0.008
R534 vss.n147 vss.n146 0.008
R535 vss.n150 vss.n149 0.008
R536 vss.n151 vss.n150 0.008
R537 vss.n152 vss.n151 0.008
R538 vss.n153 vss.n152 0.008
R539 vss.n154 vss.n153 0.008
R540 vss.n155 vss.n154 0.008
R541 vss.n156 vss.n155 0.008
R542 vss.n157 vss.n156 0.008
R543 vss.n158 vss.n157 0.008
R544 vss.n135 vss.n134 0.005
R545 vss.n158 vss.n2 0.005
R546 vss.n238 vss.n219 0.005
R547 vss.n293 vss.n292 0.005
R548 vss.n76 vss.n75 0.005
R549 vss.n64 vss.n63 0.005
R550 vss.n266 vss.n228 0.005
R551 vss.n265 vss.n229 0.005
R552 vss.n148 vss.n147 0.004
R553 vss.n149 vss.n148 0.003
R554 vss.n130 vss.n129 0.002
R555 vss.n123 vss.n122 0.002
R556 vss.n116 vss.n115 0.002
R557 vss.n109 vss.n108 0.002
R558 vss.n102 vss.n101 0.002
R559 vss.n95 vss.n94 0.002
R560 vss.n88 vss.n87 0.002
R561 vss.n81 vss.n80 0.002
R562 vss.n74 vss.n73 0.002
R563 vss.n57 vss.n56 0.002
R564 vss.n50 vss.n49 0.002
R565 vss.n43 vss.n42 0.002
R566 vss.n36 vss.n35 0.002
R567 vss.n29 vss.n28 0.002
R568 vss.n22 vss.n21 0.002
R569 vss.n15 vss.n14 0.002
R570 vss.n8 vss.n7 0.002
R571 vss.n1 vss.n0 0.002
R572 vss.n291 vss.n218 0.002
R573 vss.n288 vss.n220 0.002
R574 vss.n285 vss.n221 0.002
R575 vss.n282 vss.n222 0.002
R576 vss.n279 vss.n223 0.002
R577 vss.n276 vss.n224 0.002
R578 vss.n273 vss.n225 0.002
R579 vss.n270 vss.n226 0.002
R580 vss.n267 vss.n227 0.002
R581 vss.n264 vss.n263 0.002
R582 vss.n261 vss.n260 0.002
R583 vss.n258 vss.n257 0.002
R584 vss.n255 vss.n254 0.002
R585 vss.n252 vss.n251 0.002
R586 vss.n249 vss.n248 0.002
R587 vss.n246 vss.n245 0.002
R588 vss.n243 vss.n242 0.002
R589 vss.n240 vss.n239 0.002
R590 vss.n157 vss.n11 0.001
R591 vss.n156 vss.n18 0.001
R592 vss.n155 vss.n25 0.001
R593 vss.n154 vss.n32 0.001
R594 vss.n153 vss.n39 0.001
R595 vss.n152 vss.n46 0.001
R596 vss.n151 vss.n53 0.001
R597 vss.n150 vss.n60 0.001
R598 vss.n149 vss.n65 0.001
R599 vss.n147 vss.n77 0.001
R600 vss.n146 vss.n84 0.001
R601 vss.n145 vss.n91 0.001
R602 vss.n144 vss.n98 0.001
R603 vss.n143 vss.n105 0.001
R604 vss.n142 vss.n112 0.001
R605 vss.n141 vss.n119 0.001
R606 vss.n140 vss.n126 0.001
R607 vss.n139 vss.n133 0.001
R608 vss.n133 vss.n132 0.001
R609 vss.n126 vss.n125 0.001
R610 vss.n119 vss.n118 0.001
R611 vss.n112 vss.n111 0.001
R612 vss.n105 vss.n104 0.001
R613 vss.n98 vss.n97 0.001
R614 vss.n91 vss.n90 0.001
R615 vss.n84 vss.n83 0.001
R616 vss.n77 vss.n76 0.001
R617 vss.n65 vss.n64 0.001
R618 vss.n60 vss.n59 0.001
R619 vss.n53 vss.n52 0.001
R620 vss.n46 vss.n45 0.001
R621 vss.n39 vss.n38 0.001
R622 vss.n32 vss.n31 0.001
R623 vss.n25 vss.n24 0.001
R624 vss.n18 vss.n17 0.001
R625 vss.n11 vss.n10 0.001
R626 vss.n312 vss.n161 0.001
R627 vss.n310 vss.n167 0.001
R628 vss.n308 vss.n173 0.001
R629 vss.n306 vss.n179 0.001
R630 vss.n304 vss.n185 0.001
R631 vss.n302 vss.n191 0.001
R632 vss.n300 vss.n197 0.001
R633 vss.n298 vss.n203 0.001
R634 vss.n296 vss.n209 0.001
R635 vss.n294 vss.n215 0.001
R636 vss.n289 vss.n215 0.001
R637 vss.n283 vss.n209 0.001
R638 vss.n277 vss.n203 0.001
R639 vss.n271 vss.n197 0.001
R640 vss.n228 vss.n191 0.001
R641 vss.n262 vss.n185 0.001
R642 vss.n256 vss.n179 0.001
R643 vss.n250 vss.n173 0.001
R644 vss.n244 vss.n167 0.001
R645 vss.n238 vss.n161 0.001
R646 vss.n148 vss.n70 0.001
R647 vss.n138 vss.n135 0.001
R648 vss.n287 vss.n212 0.001
R649 vss.n295 vss.n212 0.001
R650 vss.n281 vss.n206 0.001
R651 vss.n297 vss.n206 0.001
R652 vss.n275 vss.n200 0.001
R653 vss.n299 vss.n200 0.001
R654 vss.n269 vss.n194 0.001
R655 vss.n301 vss.n194 0.001
R656 vss.n229 vss.n188 0.001
R657 vss.n303 vss.n188 0.001
R658 vss.n231 vss.n182 0.001
R659 vss.n305 vss.n182 0.001
R660 vss.n233 vss.n176 0.001
R661 vss.n307 vss.n176 0.001
R662 vss.n235 vss.n170 0.001
R663 vss.n309 vss.n170 0.001
R664 vss.n237 vss.n164 0.001
R665 vss.n311 vss.n164 0.001
R666 vt vt.t0 166.887
R667 vt.n42 vt.t65 8.632
R668 vt.n62 vt.t79 8.597
R669 vt.n102 vt.t70 8.211
R670 vt.n3 vt.t48 8.211
R671 vt.n103 vt.t2 7.146
R672 vt.n102 vt.t63 7.146
R673 vt.n101 vt.t97 7.146
R674 vt.n101 vt.t26 7.146
R675 vt.n100 vt.t73 7.146
R676 vt.n100 vt.t109 7.146
R677 vt.n99 vt.t78 7.146
R678 vt.n99 vt.t110 7.146
R679 vt.n98 vt.t71 7.146
R680 vt.n98 vt.t112 7.146
R681 vt.n97 vt.t81 7.146
R682 vt.n97 vt.t111 7.146
R683 vt.n96 vt.t85 7.146
R684 vt.n96 vt.t116 7.146
R685 vt.n95 vt.t37 7.146
R686 vt.n95 vt.t7 7.146
R687 vt.n94 vt.t86 7.146
R688 vt.n94 vt.t118 7.146
R689 vt.n93 vt.t92 7.146
R690 vt.n93 vt.t49 7.146
R691 vt.n92 vt.t1 7.146
R692 vt.n92 vt.t57 7.146
R693 vt.n91 vt.t11 7.146
R694 vt.n91 vt.t98 7.146
R695 vt.n90 vt.t15 7.146
R696 vt.n90 vt.t101 7.146
R697 vt.n89 vt.t104 7.146
R698 vt.n89 vt.t41 7.146
R699 vt.n88 vt.t17 7.146
R700 vt.n88 vt.t103 7.146
R701 vt.n87 vt.t21 7.146
R702 vt.n87 vt.t105 7.146
R703 vt.n86 vt.t62 7.146
R704 vt.n86 vt.t45 7.146
R705 vt.n85 vt.t22 7.146
R706 vt.n85 vt.t9 7.146
R707 vt.n84 vt.t28 7.146
R708 vt.n84 vt.t14 7.146
R709 vt.n83 vt.t91 7.146
R710 vt.n83 vt.t4 7.146
R711 vt.n82 vt.t31 7.146
R712 vt.n82 vt.t68 7.146
R713 vt.n81 vt.t38 7.146
R714 vt.n81 vt.t75 7.146
R715 vt.n79 vt.t13 7.146
R716 vt.n79 vt.t107 7.146
R717 vt.n78 vt.t106 7.146
R718 vt.n78 vt.t77 7.146
R719 vt.n77 vt.t108 7.146
R720 vt.n77 vt.t84 7.146
R721 vt.n72 vt.t64 7.146
R722 vt.n72 vt.t51 7.146
R723 vt.n71 vt.t42 7.146
R724 vt.n71 vt.t114 7.146
R725 vt.n70 vt.t87 7.146
R726 vt.n70 vt.t119 7.146
R727 vt.n63 vt.t58 7.146
R728 vt.n62 vt.t72 7.146
R729 vt.n43 vt.t83 7.146
R730 vt.n42 vt.t59 7.146
R731 vt.n35 vt.t100 7.146
R732 vt.n35 vt.t35 7.146
R733 vt.n34 vt.t67 7.146
R734 vt.n34 vt.t24 7.146
R735 vt.n33 vt.t76 7.146
R736 vt.n33 vt.t29 7.146
R737 vt.n28 vt.t18 7.146
R738 vt.n28 vt.t55 7.146
R739 vt.n27 vt.t50 7.146
R740 vt.n27 vt.t32 7.146
R741 vt.n26 vt.t53 7.146
R742 vt.n26 vt.t39 7.146
R743 vt.n24 vt.t6 7.146
R744 vt.n24 vt.t56 7.146
R745 vt.n23 vt.t113 7.146
R746 vt.n23 vt.t34 7.146
R747 vt.n22 vt.t120 7.146
R748 vt.n22 vt.t40 7.146
R749 vt.n21 vt.t27 7.146
R750 vt.n21 vt.t36 7.146
R751 vt.n20 vt.t74 7.146
R752 vt.n20 vt.t43 7.146
R753 vt.n19 vt.t80 7.146
R754 vt.n19 vt.t88 7.146
R755 vt.n18 vt.t82 7.146
R756 vt.n18 vt.t46 7.146
R757 vt.n17 vt.t52 7.146
R758 vt.n17 vt.t89 7.146
R759 vt.n16 vt.t54 7.146
R760 vt.n16 vt.t94 7.146
R761 vt.n15 vt.t44 7.146
R762 vt.n15 vt.t12 7.146
R763 vt.n14 vt.t5 7.146
R764 vt.n14 vt.t95 7.146
R765 vt.n13 vt.t10 7.146
R766 vt.n13 vt.t96 7.146
R767 vt.n12 vt.t3 7.146
R768 vt.n12 vt.t115 7.146
R769 vt.n11 vt.t61 7.146
R770 vt.n11 vt.t99 7.146
R771 vt.n10 vt.t69 7.146
R772 vt.n10 vt.t102 7.146
R773 vt.n9 vt.t19 7.146
R774 vt.n9 vt.t90 7.146
R775 vt.n8 vt.t16 7.146
R776 vt.n8 vt.t25 7.146
R777 vt.n7 vt.t20 7.146
R778 vt.n7 vt.t33 7.146
R779 vt.n2 vt.t47 7.146
R780 vt.n2 vt.t93 7.146
R781 vt.n1 vt.t23 7.146
R782 vt.n1 vt.t60 7.146
R783 vt.n0 vt.t30 7.146
R784 vt.n0 vt.t66 7.146
R785 vt.n4 vt.t8 7.146
R786 vt.n3 vt.t117 7.146
R787 vt.n25 vt.t190 6.774
R788 vt.n80 vt.t141 6.774
R789 vt.n25 vt.t158 5.807
R790 vt.n30 vt.t124 5.807
R791 vt.n30 vt.t147 5.807
R792 vt.n29 vt.t157 5.807
R793 vt.n29 vt.t177 5.807
R794 vt.n32 vt.t126 5.807
R795 vt.n32 vt.t139 5.807
R796 vt.n31 vt.t159 5.807
R797 vt.n31 vt.t170 5.807
R798 vt.n37 vt.t121 5.807
R799 vt.n37 vt.t142 5.807
R800 vt.n36 vt.t154 5.807
R801 vt.n36 vt.t173 5.807
R802 vt.n39 vt.t122 5.807
R803 vt.n39 vt.t187 5.807
R804 vt.n38 vt.t155 5.807
R805 vt.n38 vt.t140 5.807
R806 vt.n41 vt.t198 5.807
R807 vt.n41 vt.t191 5.807
R808 vt.n40 vt.t151 5.807
R809 vt.n40 vt.t144 5.807
R810 vt.n45 vt.t171 5.807
R811 vt.n45 vt.t183 5.807
R812 vt.n44 vt.t123 5.807
R813 vt.n44 vt.t135 5.807
R814 vt.n47 vt.t166 5.807
R815 vt.n47 vt.t185 5.807
R816 vt.n46 vt.t199 5.807
R817 vt.n46 vt.t137 5.807
R818 vt.n49 vt.t168 5.807
R819 vt.n49 vt.t180 5.807
R820 vt.n48 vt.t200 5.807
R821 vt.n48 vt.t132 5.807
R822 vt.n51 vt.t162 5.807
R823 vt.n51 vt.t156 5.807
R824 vt.n50 vt.t194 5.807
R825 vt.n50 vt.t186 5.807
R826 vt.n53 vt.t164 5.807
R827 vt.n53 vt.t152 5.807
R828 vt.n52 vt.t196 5.807
R829 vt.n52 vt.t181 5.807
R830 vt.n55 vt.t138 5.807
R831 vt.n55 vt.t153 5.807
R832 vt.n54 vt.t169 5.807
R833 vt.n54 vt.t182 5.807
R834 vt.n57 vt.t133 5.807
R835 vt.n57 vt.t146 5.807
R836 vt.n56 vt.t165 5.807
R837 vt.n56 vt.t175 5.807
R838 vt.n59 vt.t134 5.807
R839 vt.n59 vt.t149 5.807
R840 vt.n58 vt.t167 5.807
R841 vt.n58 vt.t178 5.807
R842 vt.n61 vt.t128 5.807
R843 vt.n61 vt.t195 5.807
R844 vt.n60 vt.t160 5.807
R845 vt.n60 vt.t148 5.807
R846 vt.n65 vt.t130 5.807
R847 vt.n65 vt.t197 5.807
R848 vt.n64 vt.t163 5.807
R849 vt.n64 vt.t150 5.807
R850 vt.n67 vt.t176 5.807
R851 vt.n67 vt.t189 5.807
R852 vt.n66 vt.t129 5.807
R853 vt.n66 vt.t143 5.807
R854 vt.n69 vt.t179 5.807
R855 vt.n69 vt.t192 5.807
R856 vt.n68 vt.t131 5.807
R857 vt.n68 vt.t145 5.807
R858 vt.n74 vt.t172 5.807
R859 vt.n74 vt.t184 5.807
R860 vt.n73 vt.t125 5.807
R861 vt.n73 vt.t136 5.807
R862 vt.n76 vt.t174 5.807
R863 vt.n76 vt.t161 5.807
R864 vt.n75 vt.t127 5.807
R865 vt.n75 vt.t193 5.807
R866 vt.n80 vt.t188 5.807
R867 vt.n135 vt.n30 2.241
R868 vt.n134 vt.n32 2.241
R869 vt.n132 vt.n37 2.241
R870 vt.n131 vt.n39 2.241
R871 vt.n130 vt.n41 2.241
R872 vt.n128 vt.n45 2.241
R873 vt.n127 vt.n47 2.241
R874 vt.n126 vt.n49 2.241
R875 vt.n125 vt.n51 2.241
R876 vt.n124 vt.n53 2.241
R877 vt.n123 vt.n55 2.241
R878 vt.n122 vt.n57 2.241
R879 vt.n121 vt.n59 2.241
R880 vt.n120 vt.n61 2.241
R881 vt.n118 vt.n65 2.241
R882 vt.n117 vt.n67 2.241
R883 vt.n116 vt.n69 2.241
R884 vt.n114 vt.n74 2.241
R885 vt.n113 vt.n76 2.241
R886 vt.n119 vt.n63 2.148
R887 vt.n129 vt.n43 2.148
R888 vt.n104 vt.n103 2.066
R889 vt.n137 vt.n25 1.957
R890 vt.n111 vt.n80 1.957
R891 vt.n104 vt.n101 1.912
R892 vt.n105 vt.n98 1.912
R893 vt.n106 vt.n95 1.912
R894 vt.n107 vt.n92 1.912
R895 vt.n108 vt.n89 1.912
R896 vt.n109 vt.n86 1.912
R897 vt.n110 vt.n83 1.912
R898 vt.n112 vt.n79 1.912
R899 vt.n115 vt.n72 1.912
R900 vt.n133 vt.n35 1.912
R901 vt.n136 vt.n28 1.912
R902 vt.n138 vt.n24 1.912
R903 vt.n139 vt.n21 1.912
R904 vt.n140 vt.n18 1.912
R905 vt.n141 vt.n15 1.912
R906 vt.n142 vt.n12 1.912
R907 vt.n143 vt.n9 1.912
R908 vt.n6 vt.n2 1.912
R909 vt.n5 vt.n4 1.887
R910 vt.n43 vt.n42 1.486
R911 vt.n63 vt.n62 1.459
R912 vt.n103 vt.n102 1.065
R913 vt.n4 vt.n3 1.065
R914 vt.n30 vt.n29 0.867
R915 vt.n37 vt.n36 0.867
R916 vt.n41 vt.n40 0.867
R917 vt.n47 vt.n46 0.867
R918 vt.n51 vt.n50 0.867
R919 vt.n55 vt.n54 0.867
R920 vt.n59 vt.n58 0.867
R921 vt.n65 vt.n64 0.867
R922 vt.n69 vt.n68 0.867
R923 vt.n76 vt.n75 0.867
R924 vt.n100 vt.n99 0.865
R925 vt.n101 vt.n100 0.865
R926 vt.n97 vt.n96 0.865
R927 vt.n98 vt.n97 0.865
R928 vt.n94 vt.n93 0.865
R929 vt.n95 vt.n94 0.865
R930 vt.n91 vt.n90 0.865
R931 vt.n92 vt.n91 0.865
R932 vt.n88 vt.n87 0.865
R933 vt.n89 vt.n88 0.865
R934 vt.n85 vt.n84 0.865
R935 vt.n86 vt.n85 0.865
R936 vt.n82 vt.n81 0.865
R937 vt.n83 vt.n82 0.865
R938 vt.n78 vt.n77 0.865
R939 vt.n79 vt.n78 0.865
R940 vt.n71 vt.n70 0.865
R941 vt.n72 vt.n71 0.865
R942 vt.n34 vt.n33 0.865
R943 vt.n35 vt.n34 0.865
R944 vt.n27 vt.n26 0.865
R945 vt.n28 vt.n27 0.865
R946 vt.n23 vt.n22 0.865
R947 vt.n24 vt.n23 0.865
R948 vt.n20 vt.n19 0.865
R949 vt.n21 vt.n20 0.865
R950 vt.n17 vt.n16 0.865
R951 vt.n18 vt.n17 0.865
R952 vt.n14 vt.n13 0.865
R953 vt.n15 vt.n14 0.865
R954 vt.n11 vt.n10 0.865
R955 vt.n12 vt.n11 0.865
R956 vt.n8 vt.n7 0.865
R957 vt.n9 vt.n8 0.865
R958 vt.n1 vt.n0 0.865
R959 vt.n2 vt.n1 0.865
R960 vt.n32 vt.n31 0.807
R961 vt.n39 vt.n38 0.807
R962 vt.n45 vt.n44 0.807
R963 vt.n49 vt.n48 0.807
R964 vt.n53 vt.n52 0.807
R965 vt.n57 vt.n56 0.807
R966 vt.n61 vt.n60 0.807
R967 vt.n67 vt.n66 0.807
R968 vt.n74 vt.n73 0.807
R969 vt.n6 vt.n5 0.182
R970 vt.n143 vt.n142 0.182
R971 vt.n141 vt.n140 0.182
R972 vt.n140 vt.n139 0.182
R973 vt.n139 vt.n138 0.182
R974 vt.n110 vt.n109 0.182
R975 vt.n109 vt.n108 0.182
R976 vt.n108 vt.n107 0.182
R977 vt.n107 vt.n106 0.182
R978 vt.n106 vt.n105 0.182
R979 vt.n105 vt.n104 0.182
R980 vt.n142 vt.n141 0.181
R981 vt.n138 vt.n137 0.166
R982 vt.n111 vt.n110 0.166
R983 vt vt.n143 0.135
R984 vt.n135 vt.n134 0.074
R985 vt.n132 vt.n131 0.074
R986 vt.n131 vt.n130 0.074
R987 vt.n128 vt.n127 0.074
R988 vt.n127 vt.n126 0.074
R989 vt.n126 vt.n125 0.074
R990 vt.n125 vt.n124 0.074
R991 vt.n124 vt.n123 0.074
R992 vt.n123 vt.n122 0.074
R993 vt.n122 vt.n121 0.074
R994 vt.n121 vt.n120 0.074
R995 vt.n118 vt.n117 0.074
R996 vt.n117 vt.n116 0.074
R997 vt.n114 vt.n113 0.074
R998 vt.n129 vt.n128 0.071
R999 vt.n120 vt.n119 0.071
R1000 vt.n136 vt.n135 0.059
R1001 vt.n113 vt.n112 0.059
R1002 vt.n134 vt.n133 0.048
R1003 vt.n115 vt.n114 0.048
R1004 vt vt.n6 0.047
R1005 vt.n5 vt 0.034
R1006 vt.n116 vt.n115 0.026
R1007 vt.n133 vt.n132 0.025
R1008 vt.n137 vt.n136 0.015
R1009 vt.n112 vt.n111 0.015
R1010 vt.n130 vt.n129 0.003
R1011 vt.n119 vt.n118 0.002
R1012 a_19926_29936.n9 a_19926_29936.t53 278.38
R1013 a_19926_29936.n9 a_19926_29936.t67 278.184
R1014 a_19926_29936.n6 a_19926_29936.t84 278.184
R1015 a_19926_29936.n9 a_19926_29936.t70 278.183
R1016 a_19926_29936.n9 a_19926_29936.t64 278.183
R1017 a_19926_29936.n8 a_19926_29936.t66 278.183
R1018 a_19926_29936.n8 a_19926_29936.t32 278.183
R1019 a_19926_29936.n8 a_19926_29936.t34 278.183
R1020 a_19926_29936.n8 a_19926_29936.t28 278.183
R1021 a_19926_29936.n7 a_19926_29936.t30 278.183
R1022 a_19926_29936.n7 a_19926_29936.t25 278.183
R1023 a_19926_29936.n7 a_19926_29936.t78 278.183
R1024 a_19926_29936.n7 a_19926_29936.t80 278.183
R1025 a_19926_29936.n5 a_19926_29936.t74 278.183
R1026 a_19926_29936.n5 a_19926_29936.t76 278.183
R1027 a_19926_29936.n5 a_19926_29936.t71 278.183
R1028 a_19926_29936.n5 a_19926_29936.t45 278.183
R1029 a_19926_29936.n6 a_19926_29936.t39 278.183
R1030 a_19926_29936.n6 a_19926_29936.t41 278.183
R1031 a_19926_29936.n6 a_19926_29936.t36 278.183
R1032 a_19926_29936.n6 a_19926_29936.t37 278.183
R1033 a_19926_29936.n14 a_19926_29936.t31 278.182
R1034 a_19926_29936.n9 a_19926_29936.t81 278.182
R1035 a_19926_29936.n14 a_19926_29936.t44 278.182
R1036 a_19926_29936.n14 a_19926_29936.t33 278.182
R1037 a_19926_29936.n9 a_19926_29936.t57 278.182
R1038 a_19926_29936.n14 a_19926_29936.t21 278.182
R1039 a_19926_29936.n14 a_19926_29936.t27 278.182
R1040 a_19926_29936.n8 a_19926_29936.t49 278.182
R1041 a_19926_29936.n13 a_19926_29936.t92 278.182
R1042 a_19926_29936.n13 a_19926_29936.t29 278.182
R1043 a_19926_29936.n8 a_19926_29936.t52 278.182
R1044 a_19926_29936.n13 a_19926_29936.t95 278.182
R1045 a_19926_29936.n13 a_19926_29936.t75 278.182
R1046 a_19926_29936.n8 a_19926_29936.t46 278.182
R1047 a_19926_29936.n13 a_19926_29936.t88 278.182
R1048 a_19926_29936.n13 a_19926_29936.t77 278.182
R1049 a_19926_29936.n8 a_19926_29936.t48 278.182
R1050 a_19926_29936.n13 a_19926_29936.t90 278.182
R1051 a_19926_29936.n13 a_19926_29936.t72 278.182
R1052 a_19926_29936.n7 a_19926_29936.t93 278.182
R1053 a_19926_29936.n12 a_19926_29936.t60 278.182
R1054 a_19926_29936.n12 a_19926_29936.t73 278.182
R1055 a_19926_29936.n7 a_19926_29936.t18 278.182
R1056 a_19926_29936.n12 a_19926_29936.t62 278.182
R1057 a_19926_29936.n12 a_19926_29936.t69 278.182
R1058 a_19926_29936.n7 a_19926_29936.t89 278.182
R1059 a_19926_29936.n12 a_19926_29936.t55 278.182
R1060 a_19926_29936.n12 a_19926_29936.t42 278.182
R1061 a_19926_29936.n7 a_19926_29936.t91 278.182
R1062 a_19926_29936.n12 a_19926_29936.t58 278.182
R1063 a_19926_29936.n12 a_19926_29936.t43 278.182
R1064 a_19926_29936.n5 a_19926_29936.t86 278.182
R1065 a_19926_29936.n10 a_19926_29936.t50 278.182
R1066 a_19926_29936.n10 a_19926_29936.t38 278.182
R1067 a_19926_29936.n5 a_19926_29936.t63 278.182
R1068 a_19926_29936.n10 a_19926_29936.t26 278.182
R1069 a_19926_29936.n10 a_19926_29936.t40 278.182
R1070 a_19926_29936.n5 a_19926_29936.t56 278.182
R1071 a_19926_29936.n10 a_19926_29936.t20 278.182
R1072 a_19926_29936.n10 a_19926_29936.t35 278.182
R1073 a_19926_29936.n5 a_19926_29936.t59 278.182
R1074 a_19926_29936.n10 a_19926_29936.t23 278.182
R1075 a_19926_29936.n10 a_19926_29936.t87 278.182
R1076 a_19926_29936.n6 a_19926_29936.t51 278.182
R1077 a_19926_29936.n11 a_19926_29936.t94 278.182
R1078 a_19926_29936.n11 a_19926_29936.t83 278.182
R1079 a_19926_29936.n6 a_19926_29936.t54 278.182
R1080 a_19926_29936.n11 a_19926_29936.t19 278.182
R1081 a_19926_29936.n11 a_19926_29936.t85 278.182
R1082 a_19926_29936.n6 a_19926_29936.t22 278.182
R1083 a_19926_29936.n11 a_19926_29936.t65 278.182
R1084 a_19926_29936.n11 a_19926_29936.t79 278.182
R1085 a_19926_29936.n6 a_19926_29936.t24 278.182
R1086 a_19926_29936.n11 a_19926_29936.t68 278.182
R1087 a_19926_29936.n11 a_19926_29936.t82 278.182
R1088 a_19926_29936.n6 a_19926_29936.t96 278.182
R1089 a_19926_29936.n11 a_19926_29936.t61 278.182
R1090 a_19926_29936.n11 a_19926_29936.t47 278.182
R1091 a_19926_29936.n14 a_19926_29936.t17 278.182
R1092 a_19926_29936.n17 a_19926_29936.t4 153.363
R1093 a_19926_29936.n2 a_19926_29936.t15 7.146
R1094 a_19926_29936.n2 a_19926_29936.t12 7.146
R1095 a_19926_29936.n2 a_19926_29936.t14 7.146
R1096 a_19926_29936.n1 a_19926_29936.t7 7.146
R1097 a_19926_29936.n1 a_19926_29936.t6 7.146
R1098 a_19926_29936.n4 a_19926_29936.t9 7.146
R1099 a_19926_29936.n4 a_19926_29936.t13 7.146
R1100 a_19926_29936.n4 a_19926_29936.t16 7.146
R1101 a_19926_29936.n4 a_19926_29936.t8 7.146
R1102 a_19926_29936.n3 a_19926_29936.t10 7.146
R1103 a_19926_29936.n3 a_19926_29936.t11 7.146
R1104 a_19926_29936.t5 a_19926_29936.n2 7.146
R1105 a_19926_29936.n0 a_19926_29936.t0 5.807
R1106 a_19926_29936.n0 a_19926_29936.t1 5.807
R1107 a_19926_29936.n0 a_19926_29936.t2 5.807
R1108 a_19926_29936.n0 a_19926_29936.t3 5.807
R1109 a_19926_29936.n16 a_19926_29936.n17 4.574
R1110 a_19926_29936.n16 a_19926_29936.n0 2.553
R1111 a_19926_29936.n15 a_19926_29936.n11 2.073
R1112 a_19926_29936.n15 a_19926_29936.n6 1.962
R1113 a_19926_29936.n4 a_19926_29936.n3 1.654
R1114 a_19926_29936.n2 a_19926_29936.n1 1.654
R1115 a_19926_29936.n7 a_19926_29936.n8 1.571
R1116 a_19926_29936.n5 a_19926_29936.n7 1.571
R1117 a_19926_29936.n6 a_19926_29936.n5 1.571
R1118 a_19926_29936.n12 a_19926_29936.n13 1.566
R1119 a_19926_29936.n10 a_19926_29936.n12 1.566
R1120 a_19926_29936.n11 a_19926_29936.n10 1.566
R1121 a_19926_29936.n13 a_19926_29936.n14 1.566
R1122 a_19926_29936.n17 a_19926_29936.n15 1.538
R1123 a_19926_29936.n8 a_19926_29936.n9 1.375
R1124 a_19926_29936.n2 a_19926_29936.n16 1.314
R1125 a_19926_29936.n16 a_19926_29936.n4 1.313
R1126 vsquare.n5 vsquare.t147 156.081
R1127 vsquare.n104 vsquare.t66 153.023
R1128 vsquare.n42 vsquare.t42 8.632
R1129 vsquare.n62 vsquare.t26 8.597
R1130 vsquare.n102 vsquare.t52 8.211
R1131 vsquare.n3 vsquare.t62 8.211
R1132 vsquare.n103 vsquare.t40 7.146
R1133 vsquare.n102 vsquare.t45 7.146
R1134 vsquare.n101 vsquare.t187 7.146
R1135 vsquare.n101 vsquare.t152 7.146
R1136 vsquare.n100 vsquare.t190 7.146
R1137 vsquare.n100 vsquare.t156 7.146
R1138 vsquare.n99 vsquare.t193 7.146
R1139 vsquare.n99 vsquare.t162 7.146
R1140 vsquare.n98 vsquare.t27 7.146
R1141 vsquare.n98 vsquare.t200 7.146
R1142 vsquare.n97 vsquare.t30 7.146
R1143 vsquare.n97 vsquare.t0 7.146
R1144 vsquare.n96 vsquare.t35 7.146
R1145 vsquare.n96 vsquare.t4 7.146
R1146 vsquare.n95 vsquare.t159 7.146
R1147 vsquare.n95 vsquare.t49 7.146
R1148 vsquare.n94 vsquare.t167 7.146
R1149 vsquare.n94 vsquare.t53 7.146
R1150 vsquare.n93 vsquare.t173 7.146
R1151 vsquare.n93 vsquare.t61 7.146
R1152 vsquare.n92 vsquare.t37 7.146
R1153 vsquare.n92 vsquare.t16 7.146
R1154 vsquare.n91 vsquare.t41 7.146
R1155 vsquare.n91 vsquare.t20 7.146
R1156 vsquare.n90 vsquare.t46 7.146
R1157 vsquare.n90 vsquare.t25 7.146
R1158 vsquare.n89 vsquare.t191 7.146
R1159 vsquare.n89 vsquare.t163 7.146
R1160 vsquare.n88 vsquare.t194 7.146
R1161 vsquare.n88 vsquare.t170 7.146
R1162 vsquare.n87 vsquare.t197 7.146
R1163 vsquare.n87 vsquare.t178 7.146
R1164 vsquare.n86 vsquare.t23 7.146
R1165 vsquare.n86 vsquare.t168 7.146
R1166 vsquare.n85 vsquare.t28 7.146
R1167 vsquare.n85 vsquare.t176 7.146
R1168 vsquare.n84 vsquare.t31 7.146
R1169 vsquare.n84 vsquare.t183 7.146
R1170 vsquare.n83 vsquare.t174 7.146
R1171 vsquare.n83 vsquare.t43 7.146
R1172 vsquare.n82 vsquare.t180 7.146
R1173 vsquare.n82 vsquare.t47 7.146
R1174 vsquare.n81 vsquare.t186 7.146
R1175 vsquare.n81 vsquare.t55 7.146
R1176 vsquare.n79 vsquare.t59 7.146
R1177 vsquare.n79 vsquare.t196 7.146
R1178 vsquare.n78 vsquare.t64 7.146
R1179 vsquare.n78 vsquare.t198 7.146
R1180 vsquare.n77 vsquare.t150 7.146
R1181 vsquare.n77 vsquare.t199 7.146
R1182 vsquare.n72 vsquare.t24 7.146
R1183 vsquare.n72 vsquare.t5 7.146
R1184 vsquare.n71 vsquare.t29 7.146
R1185 vsquare.n71 vsquare.t9 7.146
R1186 vsquare.n70 vsquare.t32 7.146
R1187 vsquare.n70 vsquare.t13 7.146
R1188 vsquare.n63 vsquare.t18 7.146
R1189 vsquare.n62 vsquare.t21 7.146
R1190 vsquare.n43 vsquare.t34 7.146
R1191 vsquare.n42 vsquare.t38 7.146
R1192 vsquare.n35 vsquare.t189 7.146
R1193 vsquare.n35 vsquare.t160 7.146
R1194 vsquare.n34 vsquare.t192 7.146
R1195 vsquare.n34 vsquare.t166 7.146
R1196 vsquare.n33 vsquare.t195 7.146
R1197 vsquare.n33 vsquare.t171 7.146
R1198 vsquare.n28 vsquare.t65 7.146
R1199 vsquare.n28 vsquare.t12 7.146
R1200 vsquare.n27 vsquare.t151 7.146
R1201 vsquare.n27 vsquare.t14 7.146
R1202 vsquare.n26 vsquare.t155 7.146
R1203 vsquare.n26 vsquare.t17 7.146
R1204 vsquare.n24 vsquare.t50 7.146
R1205 vsquare.n24 vsquare.t15 7.146
R1206 vsquare.n23 vsquare.t56 7.146
R1207 vsquare.n23 vsquare.t19 7.146
R1208 vsquare.n22 vsquare.t60 7.146
R1209 vsquare.n22 vsquare.t22 7.146
R1210 vsquare.n21 vsquare.t153 7.146
R1211 vsquare.n21 vsquare.t161 7.146
R1212 vsquare.n20 vsquare.t158 7.146
R1213 vsquare.n20 vsquare.t165 7.146
R1214 vsquare.n19 vsquare.t164 7.146
R1215 vsquare.n19 vsquare.t172 7.146
R1216 vsquare.n18 vsquare.t33 7.146
R1217 vsquare.n18 vsquare.t2 7.146
R1218 vsquare.n17 vsquare.t36 7.146
R1219 vsquare.n17 vsquare.t7 7.146
R1220 vsquare.n16 vsquare.t39 7.146
R1221 vsquare.n16 vsquare.t10 7.146
R1222 vsquare.n15 vsquare.t169 7.146
R1223 vsquare.n15 vsquare.t57 7.146
R1224 vsquare.n14 vsquare.t177 7.146
R1225 vsquare.n14 vsquare.t63 7.146
R1226 vsquare.n13 vsquare.t182 7.146
R1227 vsquare.n13 vsquare.t149 7.146
R1228 vsquare.n12 vsquare.t44 7.146
R1229 vsquare.n12 vsquare.t201 7.146
R1230 vsquare.n11 vsquare.t48 7.146
R1231 vsquare.n11 vsquare.t1 7.146
R1232 vsquare.n10 vsquare.t54 7.146
R1233 vsquare.n10 vsquare.t6 7.146
R1234 vsquare.n9 vsquare.t148 7.146
R1235 vsquare.n9 vsquare.t175 7.146
R1236 vsquare.n8 vsquare.t154 7.146
R1237 vsquare.n8 vsquare.t181 7.146
R1238 vsquare.n7 vsquare.t157 7.146
R1239 vsquare.n7 vsquare.t185 7.146
R1240 vsquare.n2 vsquare.t3 7.146
R1241 vsquare.n2 vsquare.t179 7.146
R1242 vsquare.n1 vsquare.t8 7.146
R1243 vsquare.n1 vsquare.t184 7.146
R1244 vsquare.n0 vsquare.t11 7.146
R1245 vsquare.n0 vsquare.t188 7.146
R1246 vsquare.n4 vsquare.t51 7.146
R1247 vsquare.n3 vsquare.t58 7.146
R1248 vsquare.n25 vsquare.t116 6.774
R1249 vsquare.n80 vsquare.t146 6.774
R1250 vsquare.n25 vsquare.t79 5.807
R1251 vsquare.n30 vsquare.t126 5.807
R1252 vsquare.n30 vsquare.t67 5.807
R1253 vsquare.n29 vsquare.t81 5.807
R1254 vsquare.n29 vsquare.t102 5.807
R1255 vsquare.n32 vsquare.t127 5.807
R1256 vsquare.n32 vsquare.t139 5.807
R1257 vsquare.n31 vsquare.t84 5.807
R1258 vsquare.n31 vsquare.t95 5.807
R1259 vsquare.n37 vsquare.t122 5.807
R1260 vsquare.n37 vsquare.t141 5.807
R1261 vsquare.n36 vsquare.t78 5.807
R1262 vsquare.n36 vsquare.t98 5.807
R1263 vsquare.n39 vsquare.t124 5.807
R1264 vsquare.n39 vsquare.t109 5.807
R1265 vsquare.n38 vsquare.t80 5.807
R1266 vsquare.n38 vsquare.t144 5.807
R1267 vsquare.n41 vsquare.t118 5.807
R1268 vsquare.n41 vsquare.t112 5.807
R1269 vsquare.n40 vsquare.t76 5.807
R1270 vsquare.n40 vsquare.t69 5.807
R1271 vsquare.n45 vsquare.t92 5.807
R1272 vsquare.n45 vsquare.t104 5.807
R1273 vsquare.n44 vsquare.t128 5.807
R1274 vsquare.n44 vsquare.t140 5.807
R1275 vsquare.n47 vsquare.t87 5.807
R1276 vsquare.n47 vsquare.t107 5.807
R1277 vsquare.n46 vsquare.t123 5.807
R1278 vsquare.n46 vsquare.t143 5.807
R1279 vsquare.n49 vsquare.t89 5.807
R1280 vsquare.n49 vsquare.t100 5.807
R1281 vsquare.n48 vsquare.t125 5.807
R1282 vsquare.n48 vsquare.t137 5.807
R1283 vsquare.n51 vsquare.t83 5.807
R1284 vsquare.n51 vsquare.t77 5.807
R1285 vsquare.n50 vsquare.t120 5.807
R1286 vsquare.n50 vsquare.t113 5.807
R1287 vsquare.n53 vsquare.t85 5.807
R1288 vsquare.n53 vsquare.t72 5.807
R1289 vsquare.n52 vsquare.t121 5.807
R1290 vsquare.n52 vsquare.t105 5.807
R1291 vsquare.n55 vsquare.t138 5.807
R1292 vsquare.n55 vsquare.t74 5.807
R1293 vsquare.n54 vsquare.t94 5.807
R1294 vsquare.n54 vsquare.t108 5.807
R1295 vsquare.n57 vsquare.t133 5.807
R1296 vsquare.n57 vsquare.t145 5.807
R1297 vsquare.n56 vsquare.t90 5.807
R1298 vsquare.n56 vsquare.t101 5.807
R1299 vsquare.n59 vsquare.t135 5.807
R1300 vsquare.n59 vsquare.t70 5.807
R1301 vsquare.n58 vsquare.t91 5.807
R1302 vsquare.n58 vsquare.t103 5.807
R1303 vsquare.n61 vsquare.t129 5.807
R1304 vsquare.n61 vsquare.t115 5.807
R1305 vsquare.n60 vsquare.t86 5.807
R1306 vsquare.n60 vsquare.t73 5.807
R1307 vsquare.n65 vsquare.t131 5.807
R1308 vsquare.n65 vsquare.t117 5.807
R1309 vsquare.n64 vsquare.t88 5.807
R1310 vsquare.n64 vsquare.t75 5.807
R1311 vsquare.n67 vsquare.t97 5.807
R1312 vsquare.n67 vsquare.t111 5.807
R1313 vsquare.n66 vsquare.t134 5.807
R1314 vsquare.n66 vsquare.t68 5.807
R1315 vsquare.n69 vsquare.t99 5.807
R1316 vsquare.n69 vsquare.t114 5.807
R1317 vsquare.n68 vsquare.t136 5.807
R1318 vsquare.n68 vsquare.t71 5.807
R1319 vsquare.n74 vsquare.t93 5.807
R1320 vsquare.n74 vsquare.t106 5.807
R1321 vsquare.n73 vsquare.t130 5.807
R1322 vsquare.n73 vsquare.t142 5.807
R1323 vsquare.n76 vsquare.t96 5.807
R1324 vsquare.n76 vsquare.t82 5.807
R1325 vsquare.n75 vsquare.t132 5.807
R1326 vsquare.n75 vsquare.t119 5.807
R1327 vsquare.n80 vsquare.t110 5.807
R1328 vsquare.n136 vsquare.n30 2.241
R1329 vsquare.n135 vsquare.n32 2.241
R1330 vsquare.n133 vsquare.n37 2.241
R1331 vsquare.n132 vsquare.n39 2.241
R1332 vsquare.n131 vsquare.n41 2.241
R1333 vsquare.n129 vsquare.n45 2.241
R1334 vsquare.n128 vsquare.n47 2.241
R1335 vsquare.n127 vsquare.n49 2.241
R1336 vsquare.n126 vsquare.n51 2.241
R1337 vsquare.n125 vsquare.n53 2.241
R1338 vsquare.n124 vsquare.n55 2.241
R1339 vsquare.n123 vsquare.n57 2.241
R1340 vsquare.n122 vsquare.n59 2.241
R1341 vsquare.n121 vsquare.n61 2.241
R1342 vsquare.n119 vsquare.n65 2.241
R1343 vsquare.n118 vsquare.n67 2.241
R1344 vsquare.n117 vsquare.n69 2.241
R1345 vsquare.n115 vsquare.n74 2.241
R1346 vsquare.n114 vsquare.n76 2.241
R1347 vsquare.n120 vsquare.n63 2.148
R1348 vsquare.n130 vsquare.n43 2.148
R1349 vsquare.n138 vsquare.n25 1.957
R1350 vsquare.n112 vsquare.n80 1.957
R1351 vsquare.n105 vsquare.n101 1.912
R1352 vsquare.n106 vsquare.n98 1.912
R1353 vsquare.n107 vsquare.n95 1.912
R1354 vsquare.n108 vsquare.n92 1.912
R1355 vsquare.n109 vsquare.n89 1.912
R1356 vsquare.n110 vsquare.n86 1.912
R1357 vsquare.n111 vsquare.n83 1.912
R1358 vsquare.n113 vsquare.n79 1.912
R1359 vsquare.n116 vsquare.n72 1.912
R1360 vsquare.n134 vsquare.n35 1.912
R1361 vsquare.n137 vsquare.n28 1.912
R1362 vsquare.n139 vsquare.n24 1.912
R1363 vsquare.n140 vsquare.n21 1.912
R1364 vsquare.n141 vsquare.n18 1.912
R1365 vsquare.n142 vsquare.n15 1.912
R1366 vsquare.n143 vsquare.n12 1.912
R1367 vsquare.n144 vsquare.n9 1.912
R1368 vsquare.n6 vsquare.n2 1.912
R1369 vsquare.n104 vsquare.n103 1.887
R1370 vsquare.n5 vsquare.n4 1.887
R1371 vsquare.n43 vsquare.n42 1.486
R1372 vsquare.n63 vsquare.n62 1.459
R1373 vsquare.n103 vsquare.n102 1.065
R1374 vsquare.n4 vsquare.n3 1.065
R1375 vsquare.n30 vsquare.n29 0.867
R1376 vsquare.n37 vsquare.n36 0.867
R1377 vsquare.n41 vsquare.n40 0.867
R1378 vsquare.n47 vsquare.n46 0.867
R1379 vsquare.n51 vsquare.n50 0.867
R1380 vsquare.n55 vsquare.n54 0.867
R1381 vsquare.n59 vsquare.n58 0.867
R1382 vsquare.n65 vsquare.n64 0.867
R1383 vsquare.n69 vsquare.n68 0.867
R1384 vsquare.n76 vsquare.n75 0.867
R1385 vsquare.n100 vsquare.n99 0.865
R1386 vsquare.n101 vsquare.n100 0.865
R1387 vsquare.n97 vsquare.n96 0.865
R1388 vsquare.n98 vsquare.n97 0.865
R1389 vsquare.n94 vsquare.n93 0.865
R1390 vsquare.n95 vsquare.n94 0.865
R1391 vsquare.n91 vsquare.n90 0.865
R1392 vsquare.n92 vsquare.n91 0.865
R1393 vsquare.n88 vsquare.n87 0.865
R1394 vsquare.n89 vsquare.n88 0.865
R1395 vsquare.n85 vsquare.n84 0.865
R1396 vsquare.n86 vsquare.n85 0.865
R1397 vsquare.n82 vsquare.n81 0.865
R1398 vsquare.n83 vsquare.n82 0.865
R1399 vsquare.n78 vsquare.n77 0.865
R1400 vsquare.n79 vsquare.n78 0.865
R1401 vsquare.n71 vsquare.n70 0.865
R1402 vsquare.n72 vsquare.n71 0.865
R1403 vsquare.n34 vsquare.n33 0.865
R1404 vsquare.n35 vsquare.n34 0.865
R1405 vsquare.n27 vsquare.n26 0.865
R1406 vsquare.n28 vsquare.n27 0.865
R1407 vsquare.n23 vsquare.n22 0.865
R1408 vsquare.n24 vsquare.n23 0.865
R1409 vsquare.n20 vsquare.n19 0.865
R1410 vsquare.n21 vsquare.n20 0.865
R1411 vsquare.n17 vsquare.n16 0.865
R1412 vsquare.n18 vsquare.n17 0.865
R1413 vsquare.n14 vsquare.n13 0.865
R1414 vsquare.n15 vsquare.n14 0.865
R1415 vsquare.n11 vsquare.n10 0.865
R1416 vsquare.n12 vsquare.n11 0.865
R1417 vsquare.n8 vsquare.n7 0.865
R1418 vsquare.n9 vsquare.n8 0.865
R1419 vsquare.n1 vsquare.n0 0.865
R1420 vsquare.n2 vsquare.n1 0.865
R1421 vsquare.n32 vsquare.n31 0.807
R1422 vsquare.n39 vsquare.n38 0.807
R1423 vsquare.n45 vsquare.n44 0.807
R1424 vsquare.n49 vsquare.n48 0.807
R1425 vsquare.n53 vsquare.n52 0.807
R1426 vsquare.n57 vsquare.n56 0.807
R1427 vsquare.n61 vsquare.n60 0.807
R1428 vsquare.n67 vsquare.n66 0.807
R1429 vsquare.n74 vsquare.n73 0.807
R1430 vsquare.n6 vsquare.n5 0.17
R1431 vsquare.n144 vsquare.n143 0.17
R1432 vsquare.n143 vsquare.n142 0.17
R1433 vsquare.n142 vsquare.n141 0.17
R1434 vsquare.n141 vsquare.n140 0.17
R1435 vsquare.n140 vsquare.n139 0.17
R1436 vsquare.n111 vsquare.n110 0.17
R1437 vsquare.n110 vsquare.n109 0.17
R1438 vsquare.n109 vsquare.n108 0.17
R1439 vsquare.n108 vsquare.n107 0.17
R1440 vsquare.n107 vsquare.n106 0.17
R1441 vsquare.n106 vsquare.n105 0.17
R1442 vsquare.n105 vsquare.n104 0.17
R1443 vsquare.n139 vsquare.n138 0.155
R1444 vsquare.n112 vsquare.n111 0.155
R1445 vsquare vsquare.n144 0.12
R1446 vsquare.n136 vsquare.n135 0.069
R1447 vsquare.n133 vsquare.n132 0.069
R1448 vsquare.n132 vsquare.n131 0.069
R1449 vsquare.n129 vsquare.n128 0.069
R1450 vsquare.n128 vsquare.n127 0.069
R1451 vsquare.n127 vsquare.n126 0.069
R1452 vsquare.n126 vsquare.n125 0.069
R1453 vsquare.n125 vsquare.n124 0.069
R1454 vsquare.n124 vsquare.n123 0.069
R1455 vsquare.n123 vsquare.n122 0.069
R1456 vsquare.n122 vsquare.n121 0.069
R1457 vsquare.n119 vsquare.n118 0.069
R1458 vsquare.n118 vsquare.n117 0.069
R1459 vsquare.n115 vsquare.n114 0.069
R1460 vsquare.n130 vsquare.n129 0.066
R1461 vsquare.n121 vsquare.n120 0.066
R1462 vsquare.n137 vsquare.n136 0.055
R1463 vsquare.n114 vsquare.n113 0.055
R1464 vsquare.n135 vsquare.n134 0.045
R1465 vsquare.n116 vsquare.n115 0.045
R1466 vsquare vsquare.n6 0.044
R1467 vsquare.n134 vsquare.n133 0.024
R1468 vsquare.n117 vsquare.n116 0.024
R1469 vsquare.n138 vsquare.n137 0.014
R1470 vsquare.n113 vsquare.n112 0.014
R1471 vsquare.n131 vsquare.n130 0.003
R1472 vsquare.n120 vsquare.n119 0.002
R1473 vbias2.n315 vbias2.n314 160.035
R1474 vbias2.n231 vbias2.n230 160.035
R1475 vbias2.n499 vbias2.n498 160.035
R1476 vbias2.n315 vbias2.n313 160.035
R1477 vbias2.n239 vbias2.n238 160.035
R1478 vbias2.n231 vbias2.n229 160.035
R1479 vbias2.n495 vbias2.n494 71.764
R1480 vbias2.n309 vbias2.n307 59.923
R1481 vbias2.n305 vbias2.n298 59.923
R1482 vbias2.n242 vbias2.n241 57.119
R1483 vbias2.n64 vbias2.t148 55.915
R1484 vbias2.n468 vbias2.t32 55.915
R1485 vbias2.n460 vbias2.t75 55.915
R1486 vbias2.n444 vbias2.t125 55.915
R1487 vbias2.n428 vbias2.t51 55.915
R1488 vbias2.n412 vbias2.t136 55.915
R1489 vbias2.n396 vbias2.t79 55.915
R1490 vbias2.n380 vbias2.t121 55.915
R1491 vbias2.n364 vbias2.t66 55.915
R1492 vbias2.n348 vbias2.t26 55.915
R1493 vbias2.n332 vbias2.t122 55.915
R1494 vbias2.n340 vbias2.t94 55.915
R1495 vbias2.n356 vbias2.t80 55.915
R1496 vbias2.n372 vbias2.t137 55.915
R1497 vbias2.n388 vbias2.t54 55.915
R1498 vbias2.n404 vbias2.t47 55.915
R1499 vbias2.n420 vbias2.t110 55.915
R1500 vbias2.n436 vbias2.t143 55.915
R1501 vbias2.n452 vbias2.t84 55.915
R1502 vbias2.n522 vbias2.t142 55.915
R1503 vbias2.n226 vbias2.t132 55.915
R1504 vbias2.n217 vbias2.t43 55.915
R1505 vbias2.n208 vbias2.t77 55.915
R1506 vbias2.n199 vbias2.t103 55.915
R1507 vbias2.n190 vbias2.t31 55.915
R1508 vbias2.n181 vbias2.t109 55.915
R1509 vbias2.n172 vbias2.t150 55.915
R1510 vbias2.n163 vbias2.t42 55.915
R1511 vbias2.n154 vbias2.t40 55.915
R1512 vbias2.n145 vbias2.t92 55.915
R1513 vbias2.n136 vbias2.t129 55.915
R1514 vbias2.n127 vbias2.t153 55.915
R1515 vbias2.n118 vbias2.t61 55.915
R1516 vbias2.n109 vbias2.t85 55.915
R1517 vbias2.n100 vbias2.t144 55.915
R1518 vbias2.n91 vbias2.t60 55.915
R1519 vbias2.n82 vbias2.t33 55.915
R1520 vbias2.n73 vbias2.t64 55.915
R1521 vbias2.n62 vbias2.t98 55.915
R1522 vbias2.n324 vbias2.t111 55.915
R1523 vbias2.t111 vbias2.n319 55.915
R1524 vbias2.n327 vbias2.t114 55.915
R1525 vbias2.n335 vbias2.t89 55.915
R1526 vbias2.n343 vbias2.t149 55.915
R1527 vbias2.n351 vbias2.t78 55.915
R1528 vbias2.n359 vbias2.t52 55.915
R1529 vbias2.n367 vbias2.t133 55.915
R1530 vbias2.n375 vbias2.t113 55.915
R1531 vbias2.n383 vbias2.t45 55.915
R1532 vbias2.n391 vbias2.t73 55.915
R1533 vbias2.n399 vbias2.t39 55.915
R1534 vbias2.n407 vbias2.t127 55.915
R1535 vbias2.n415 vbias2.t106 55.915
R1536 vbias2.n423 vbias2.t35 55.915
R1537 vbias2.n431 vbias2.t139 55.915
R1538 vbias2.n439 vbias2.t117 55.915
R1539 vbias2.n447 vbias2.t82 55.915
R1540 vbias2.n455 vbias2.t67 55.915
R1541 vbias2.n463 vbias2.t28 55.915
R1542 vbias2.n521 vbias2.t130 55.915
R1543 vbias2.t128 vbias2.n221 55.915
R1544 vbias2.t43 vbias2.n212 55.915
R1545 vbias2.t74 vbias2.n203 55.915
R1546 vbias2.t103 vbias2.n194 55.915
R1547 vbias2.t27 vbias2.n185 55.915
R1548 vbias2.t109 vbias2.n176 55.915
R1549 vbias2.t146 vbias2.n167 55.915
R1550 vbias2.t42 vbias2.n158 55.915
R1551 vbias2.t34 vbias2.n149 55.915
R1552 vbias2.t92 vbias2.n140 55.915
R1553 vbias2.t126 vbias2.n131 55.915
R1554 vbias2.t153 vbias2.n122 55.915
R1555 vbias2.t55 vbias2.n113 55.915
R1556 vbias2.t85 vbias2.n104 55.915
R1557 vbias2.t138 vbias2.n95 55.915
R1558 vbias2.t60 vbias2.n86 55.915
R1559 vbias2.t30 vbias2.n77 55.915
R1560 vbias2.t64 vbias2.n68 55.915
R1561 vbias2.t93 vbias2.n57 55.915
R1562 vbias2.t148 vbias2.n63 55.915
R1563 vbias2.t87 vbias2.n55 55.915
R1564 vbias2.n63 vbias2.t141 55.915
R1565 vbias2.n57 vbias2.t87 55.915
R1566 vbias2.n62 vbias2.t93 55.915
R1567 vbias2.n68 vbias2.t57 55.915
R1568 vbias2.n73 vbias2.t69 55.915
R1569 vbias2.n77 vbias2.t24 55.915
R1570 vbias2.n82 vbias2.t30 55.915
R1571 vbias2.n86 vbias2.t53 55.915
R1572 vbias2.n91 vbias2.t65 55.915
R1573 vbias2.n95 vbias2.t134 55.915
R1574 vbias2.n100 vbias2.t138 55.915
R1575 vbias2.n104 vbias2.t83 55.915
R1576 vbias2.n109 vbias2.t90 55.915
R1577 vbias2.n113 vbias2.t46 55.915
R1578 vbias2.n118 vbias2.t55 55.915
R1579 vbias2.n122 vbias2.t147 55.915
R1580 vbias2.n127 vbias2.t25 55.915
R1581 vbias2.n131 vbias2.t123 55.915
R1582 vbias2.n136 vbias2.t126 55.915
R1583 vbias2.n140 vbias2.t86 55.915
R1584 vbias2.n145 vbias2.t96 55.915
R1585 vbias2.n149 vbias2.t29 55.915
R1586 vbias2.n154 vbias2.t34 55.915
R1587 vbias2.n158 vbias2.t37 55.915
R1588 vbias2.n163 vbias2.t50 55.915
R1589 vbias2.n167 vbias2.t140 55.915
R1590 vbias2.n172 vbias2.t146 55.915
R1591 vbias2.n176 vbias2.t104 55.915
R1592 vbias2.n181 vbias2.t112 55.915
R1593 vbias2.n185 vbias2.t155 55.915
R1594 vbias2.n190 vbias2.t27 55.915
R1595 vbias2.n194 vbias2.t99 55.915
R1596 vbias2.n199 vbias2.t107 55.915
R1597 vbias2.n203 vbias2.t70 55.915
R1598 vbias2.n208 vbias2.t74 55.915
R1599 vbias2.n212 vbias2.t36 55.915
R1600 vbias2.n217 vbias2.t49 55.915
R1601 vbias2.n221 vbias2.t124 55.915
R1602 vbias2.n226 vbias2.t128 55.915
R1603 vbias2.n460 vbias2.t71 55.915
R1604 vbias2.n444 vbias2.t120 55.915
R1605 vbias2.n428 vbias2.t44 55.915
R1606 vbias2.n412 vbias2.t131 55.915
R1607 vbias2.n396 vbias2.t76 55.915
R1608 vbias2.n380 vbias2.t118 55.915
R1609 vbias2.n364 vbias2.t59 55.915
R1610 vbias2.n348 vbias2.t154 55.915
R1611 vbias2.n332 vbias2.t119 55.915
R1612 vbias2.n522 vbias2.t135 55.915
R1613 vbias2.n468 vbias2.t38 55.915
R1614 vbias2.n452 vbias2.t88 55.915
R1615 vbias2.n436 vbias2.t151 55.915
R1616 vbias2.n420 vbias2.t115 55.915
R1617 vbias2.n404 vbias2.t56 55.915
R1618 vbias2.n388 vbias2.t62 55.915
R1619 vbias2.n372 vbias2.t145 55.915
R1620 vbias2.n356 vbias2.t81 55.915
R1621 vbias2.n340 vbias2.t100 55.915
R1622 vbias2.n324 vbias2.t116 55.915
R1623 vbias2.n319 vbias2.t108 55.915
R1624 vbias2.t32 vbias2.n463 55.915
R1625 vbias2.t71 vbias2.n455 55.915
R1626 vbias2.t84 vbias2.n447 55.915
R1627 vbias2.t120 vbias2.n439 55.915
R1628 vbias2.t143 vbias2.n431 55.915
R1629 vbias2.t44 vbias2.n423 55.915
R1630 vbias2.t110 vbias2.n415 55.915
R1631 vbias2.t131 vbias2.n407 55.915
R1632 vbias2.t47 vbias2.n399 55.915
R1633 vbias2.t76 vbias2.n391 55.915
R1634 vbias2.t54 vbias2.n383 55.915
R1635 vbias2.t118 vbias2.n375 55.915
R1636 vbias2.t137 vbias2.n367 55.915
R1637 vbias2.t59 vbias2.n359 55.915
R1638 vbias2.t80 vbias2.n351 55.915
R1639 vbias2.t154 vbias2.n343 55.915
R1640 vbias2.t94 vbias2.n335 55.915
R1641 vbias2.t119 vbias2.n327 55.915
R1642 vbias2.t135 vbias2.n521 55.915
R1643 vbias2.n476 vbias2.t63 55.914
R1644 vbias2.n491 vbias2.t97 55.914
R1645 vbias2.n474 vbias2.t8 55.914
R1646 vbias2.n471 vbias2.t41 55.914
R1647 vbias2.n496 vbias2.t2 55.914
R1648 vbias2.n486 vbias2.t20 55.914
R1649 vbias2.n243 vbias2.t12 55.914
R1650 vbias2.t16 vbias2.n243 55.914
R1651 vbias2.n64 vbias2.t152 55.914
R1652 vbias2.t98 vbias2.n61 55.914
R1653 vbias2.t57 vbias2.n66 55.914
R1654 vbias2.t69 vbias2.n72 55.914
R1655 vbias2.t24 vbias2.n75 55.914
R1656 vbias2.t33 vbias2.n81 55.914
R1657 vbias2.t53 vbias2.n84 55.914
R1658 vbias2.t65 vbias2.n90 55.914
R1659 vbias2.t134 vbias2.n93 55.914
R1660 vbias2.t144 vbias2.n99 55.914
R1661 vbias2.t83 vbias2.n102 55.914
R1662 vbias2.t90 vbias2.n108 55.914
R1663 vbias2.t46 vbias2.n111 55.914
R1664 vbias2.t61 vbias2.n117 55.914
R1665 vbias2.t147 vbias2.n120 55.914
R1666 vbias2.t25 vbias2.n126 55.914
R1667 vbias2.t123 vbias2.n129 55.914
R1668 vbias2.t129 vbias2.n135 55.914
R1669 vbias2.t86 vbias2.n138 55.914
R1670 vbias2.t96 vbias2.n144 55.914
R1671 vbias2.t29 vbias2.n147 55.914
R1672 vbias2.t40 vbias2.n153 55.914
R1673 vbias2.t37 vbias2.n156 55.914
R1674 vbias2.t50 vbias2.n162 55.914
R1675 vbias2.t140 vbias2.n165 55.914
R1676 vbias2.t150 vbias2.n171 55.914
R1677 vbias2.t104 vbias2.n174 55.914
R1678 vbias2.t112 vbias2.n180 55.914
R1679 vbias2.t155 vbias2.n183 55.914
R1680 vbias2.t31 vbias2.n189 55.914
R1681 vbias2.t99 vbias2.n192 55.914
R1682 vbias2.t107 vbias2.n198 55.914
R1683 vbias2.t70 vbias2.n201 55.914
R1684 vbias2.t77 vbias2.n207 55.914
R1685 vbias2.t36 vbias2.n210 55.914
R1686 vbias2.t49 vbias2.n216 55.914
R1687 vbias2.t124 vbias2.n219 55.914
R1688 vbias2.t132 vbias2.n225 55.914
R1689 vbias2.t91 vbias2.n477 55.914
R1690 vbias2.t101 vbias2.n267 55.914
R1691 vbias2.t63 vbias2.n475 55.914
R1692 vbias2.t105 vbias2.n25 55.914
R1693 vbias2.t97 vbias2.n490 55.914
R1694 vbias2.t8 vbias2.n473 55.914
R1695 vbias2.t41 vbias2.n470 55.914
R1696 vbias2.t58 vbias2.n7 55.914
R1697 vbias2.t2 vbias2.n495 55.914
R1698 vbias2.t18 vbias2.n303 55.914
R1699 vbias2.t28 vbias2.n462 55.914
R1700 vbias2.t67 vbias2.n454 55.914
R1701 vbias2.t75 vbias2.n459 55.914
R1702 vbias2.t82 vbias2.n446 55.914
R1703 vbias2.t88 vbias2.n451 55.914
R1704 vbias2.t117 vbias2.n438 55.914
R1705 vbias2.t125 vbias2.n443 55.914
R1706 vbias2.t139 vbias2.n430 55.914
R1707 vbias2.t151 vbias2.n435 55.914
R1708 vbias2.t35 vbias2.n422 55.914
R1709 vbias2.t51 vbias2.n427 55.914
R1710 vbias2.t106 vbias2.n414 55.914
R1711 vbias2.t115 vbias2.n419 55.914
R1712 vbias2.t127 vbias2.n406 55.914
R1713 vbias2.t136 vbias2.n411 55.914
R1714 vbias2.t39 vbias2.n398 55.914
R1715 vbias2.t56 vbias2.n403 55.914
R1716 vbias2.t73 vbias2.n390 55.914
R1717 vbias2.t79 vbias2.n395 55.914
R1718 vbias2.t45 vbias2.n382 55.914
R1719 vbias2.t62 vbias2.n387 55.914
R1720 vbias2.t113 vbias2.n374 55.914
R1721 vbias2.t121 vbias2.n379 55.914
R1722 vbias2.t133 vbias2.n366 55.914
R1723 vbias2.t145 vbias2.n371 55.914
R1724 vbias2.t52 vbias2.n358 55.914
R1725 vbias2.t66 vbias2.n363 55.914
R1726 vbias2.t78 vbias2.n350 55.914
R1727 vbias2.t81 vbias2.n355 55.914
R1728 vbias2.t149 vbias2.n342 55.914
R1729 vbias2.t26 vbias2.n347 55.914
R1730 vbias2.t89 vbias2.n334 55.914
R1731 vbias2.t100 vbias2.n339 55.914
R1732 vbias2.t114 vbias2.n326 55.914
R1733 vbias2.t122 vbias2.n331 55.914
R1734 vbias2.t38 vbias2.n467 55.914
R1735 vbias2.t14 vbias2.n35 55.914
R1736 vbias2.t72 vbias2.n48 55.914
R1737 vbias2.t20 vbias2.n485 55.914
R1738 vbias2.t12 vbias2.n237 55.914
R1739 vbias2.t10 vbias2.n251 55.914
R1740 vbias2.t0 vbias2.n284 55.914
R1741 vbias2.t116 vbias2.n323 55.914
R1742 vbias2.t108 vbias2.n318 55.914
R1743 vbias2.n478 vbias2.t91 55.912
R1744 vbias2.n268 vbias2.t101 55.912
R1745 vbias2.n261 vbias2.t95 55.912
R1746 vbias2.t95 vbias2.n260 55.912
R1747 vbias2.n26 vbias2.t105 55.912
R1748 vbias2.n19 vbias2.t102 55.912
R1749 vbias2.n39 vbias2.t4 55.912
R1750 vbias2.n11 vbias2.t48 55.912
R1751 vbias2.n8 vbias2.t58 55.912
R1752 vbias2.n308 vbias2.t6 55.912
R1753 vbias2.n304 vbias2.t18 55.912
R1754 vbias2.n36 vbias2.t14 55.912
R1755 vbias2.n49 vbias2.t72 55.912
R1756 vbias2.n52 vbias2.t68 55.912
R1757 vbias2.n278 vbias2.t22 55.912
R1758 vbias2.n244 vbias2.t16 55.912
R1759 vbias2.n252 vbias2.t10 55.912
R1760 vbias2.n285 vbias2.t0 55.912
R1761 vbias2.n250 vbias2.n249 54.492
R1762 vbias2.n300 vbias2.n299 52.343
R1763 vbias2.n297 vbias2.n0 48.571
R1764 vbias2.n294 vbias2.n293 45.634
R1765 vbias2.n289 vbias2.n288 37.195
R1766 vbias2.n290 vbias2.n289 37.195
R1767 vbias2.n293 vbias2.n290 37.195
R1768 vbias2.n293 vbias2.n292 37.195
R1769 vbias2.n292 vbias2.n291 32.954
R1770 vbias2.n240 vbias2.n239 19.786
R1771 vbias2.n500 vbias2.n499 19.786
R1772 vbias2.n316 vbias2.n315 16.988
R1773 vbias2.n16 vbias2.n15 12.2
R1774 vbias2.n276 vbias2.n275 12.2
R1775 vbias2.n257 vbias2.n256 12.2
R1776 vbias2.n233 vbias2.n232 12.2
R1777 vbias2.n229 vbias2.t17 7.141
R1778 vbias2.n238 vbias2.t13 7.141
R1779 vbias2.n290 vbias2.t23 7.141
R1780 vbias2.n290 vbias2.t5 7.141
R1781 vbias2.n288 vbias2.t9 7.141
R1782 vbias2.n288 vbias2.t21 7.141
R1783 vbias2.n292 vbias2.t1 7.141
R1784 vbias2.n292 vbias2.t15 7.141
R1785 vbias2.n313 vbias2.t7 7.141
R1786 vbias2.n498 vbias2.t3 7.141
R1787 vbias2.n230 vbias2.t11 7.141
R1788 vbias2.n314 vbias2.t19 7.141
R1789 vbias2.n18 vbias2.n17 3.897
R1790 vbias2.n31 vbias2.n29 3.897
R1791 vbias2.n31 vbias2.n30 3.897
R1792 vbias2.n18 vbias2.n16 3.897
R1793 vbias2.n3 vbias2.n1 3.897
R1794 vbias2.n3 vbias2.n2 3.897
R1795 vbias2.n44 vbias2.n42 3.897
R1796 vbias2.n277 vbias2.n274 3.897
R1797 vbias2.n277 vbias2.n276 3.897
R1798 vbias2.n44 vbias2.n43 3.897
R1799 vbias2.n259 vbias2.n257 3.897
R1800 vbias2.n259 vbias2.n258 3.897
R1801 vbias2.n235 vbias2.n233 3.897
R1802 vbias2.n235 vbias2.n234 3.897
R1803 vbias2.n232 vbias2.n231 3.275
R1804 vbias2.n312 vbias2.n297 0.55
R1805 vbias2.n65 vbias2.n64 0.548
R1806 vbias2.n484 vbias2.n483 0.547
R1807 vbias2.n497 vbias2.n493 0.546
R1808 vbias2.n492 vbias2.n489 0.546
R1809 vbias2.n487 vbias2.n484 0.546
R1810 vbias2.n493 vbias2.n492 0.545
R1811 vbias2.n503 vbias2.n502 0.545
R1812 vbias2.n502 vbias2.n501 0.544
R1813 vbias2.n341 vbias2.n333 0.544
R1814 vbias2.n349 vbias2.n341 0.544
R1815 vbias2.n357 vbias2.n349 0.544
R1816 vbias2.n365 vbias2.n357 0.544
R1817 vbias2.n373 vbias2.n365 0.544
R1818 vbias2.n381 vbias2.n373 0.544
R1819 vbias2.n389 vbias2.n381 0.544
R1820 vbias2.n397 vbias2.n389 0.544
R1821 vbias2.n405 vbias2.n397 0.544
R1822 vbias2.n413 vbias2.n405 0.544
R1823 vbias2.n421 vbias2.n413 0.544
R1824 vbias2.n429 vbias2.n421 0.544
R1825 vbias2.n437 vbias2.n429 0.544
R1826 vbias2.n445 vbias2.n437 0.544
R1827 vbias2.n453 vbias2.n445 0.544
R1828 vbias2.n461 vbias2.n453 0.544
R1829 vbias2.n469 vbias2.n461 0.544
R1830 vbias2.n333 vbias2.n325 0.544
R1831 vbias2.n523 vbias2.n469 0.544
R1832 vbias2.n504 vbias2.n503 0.544
R1833 vbias2.n505 vbias2.n504 0.544
R1834 vbias2.n506 vbias2.n505 0.544
R1835 vbias2.n507 vbias2.n506 0.544
R1836 vbias2.n508 vbias2.n507 0.544
R1837 vbias2.n509 vbias2.n508 0.544
R1838 vbias2.n510 vbias2.n509 0.544
R1839 vbias2.n511 vbias2.n510 0.544
R1840 vbias2.n512 vbias2.n511 0.544
R1841 vbias2.n513 vbias2.n512 0.544
R1842 vbias2.n514 vbias2.n513 0.544
R1843 vbias2.n515 vbias2.n514 0.544
R1844 vbias2.n516 vbias2.n515 0.544
R1845 vbias2.n517 vbias2.n516 0.544
R1846 vbias2.n518 vbias2.n517 0.544
R1847 vbias2.n519 vbias2.n518 0.544
R1848 vbias2.n520 vbias2.n519 0.544
R1849 vbias2.n297 vbias2.n296 0.542
R1850 vbias2.n296 vbias2.n295 0.542
R1851 vbias2.n295 vbias2.n294 0.542
R1852 vbias2.n294 vbias2.n273 0.542
R1853 vbias2.n255 vbias2.n228 0.542
R1854 vbias2.n272 vbias2.n255 0.542
R1855 vbias2.n273 vbias2.n272 0.542
R1856 vbias2.n83 vbias2.n74 0.537
R1857 vbias2.n92 vbias2.n83 0.537
R1858 vbias2.n101 vbias2.n92 0.537
R1859 vbias2.n110 vbias2.n101 0.537
R1860 vbias2.n119 vbias2.n110 0.537
R1861 vbias2.n128 vbias2.n119 0.537
R1862 vbias2.n137 vbias2.n128 0.537
R1863 vbias2.n146 vbias2.n137 0.537
R1864 vbias2.n155 vbias2.n146 0.537
R1865 vbias2.n164 vbias2.n155 0.537
R1866 vbias2.n173 vbias2.n164 0.537
R1867 vbias2.n182 vbias2.n173 0.537
R1868 vbias2.n191 vbias2.n182 0.537
R1869 vbias2.n200 vbias2.n191 0.537
R1870 vbias2.n209 vbias2.n200 0.537
R1871 vbias2.n218 vbias2.n209 0.537
R1872 vbias2.n227 vbias2.n218 0.537
R1873 vbias2.n74 vbias2.n65 0.537
R1874 vbias2.n473 vbias2.n472 0.498
R1875 vbias2.n237 vbias2.n236 0.381
R1876 vbias2.n520 vbias2 0.335
R1877 vbias2.n325 vbias2.n316 0.311
R1878 vbias2.n501 vbias2.n500 0.277
R1879 vbias2.n489 vbias2.n488 0.274
R1880 vbias2.n488 vbias2.n487 0.273
R1881 vbias2.n242 vbias2.n240 0.268
R1882 vbias2.n500 vbias2.n497 0.268
R1883 vbias2.n316 vbias2.n312 0.228
R1884 vbias2.n310 vbias2.n306 0.176
R1885 vbias2.n51 vbias2.n44 0.175
R1886 vbias2.n280 vbias2.n277 0.175
R1887 vbias2.n10 vbias2.n3 0.175
R1888 vbias2.n38 vbias2.n31 0.175
R1889 vbias2.n21 vbias2.n18 0.175
R1890 vbias2.n263 vbias2.n259 0.175
R1891 vbias2.n246 vbias2.n235 0.175
R1892 vbias2.n61 vbias2.n60 0.033
R1893 vbias2.n224 vbias2.n223 0.027
R1894 vbias2.n206 vbias2.n205 0.027
R1895 vbias2.n188 vbias2.n187 0.027
R1896 vbias2.n170 vbias2.n169 0.027
R1897 vbias2.n152 vbias2.n151 0.027
R1898 vbias2.n134 vbias2.n133 0.027
R1899 vbias2.n116 vbias2.n115 0.027
R1900 vbias2.n98 vbias2.n97 0.027
R1901 vbias2.n80 vbias2.n79 0.027
R1902 vbias2.n71 vbias2.n70 0.027
R1903 vbias2.n89 vbias2.n88 0.027
R1904 vbias2.n107 vbias2.n106 0.027
R1905 vbias2.n125 vbias2.n124 0.027
R1906 vbias2.n143 vbias2.n142 0.027
R1907 vbias2.n161 vbias2.n160 0.027
R1908 vbias2.n179 vbias2.n178 0.027
R1909 vbias2.n197 vbias2.n196 0.027
R1910 vbias2.n215 vbias2.n214 0.027
R1911 vbias2.n283 vbias2.n282 0.027
R1912 vbias2.n47 vbias2.n46 0.027
R1913 vbias2.n266 vbias2.n265 0.027
R1914 vbias2.n24 vbias2.n23 0.027
R1915 vbias2.n6 vbias2.n5 0.027
R1916 vbias2.n302 vbias2.n301 0.027
R1917 vbias2.n34 vbias2.n33 0.027
R1918 vbias2.n250 vbias2.n248 0.027
R1919 vbias2.n467 vbias2.n466 0.024
R1920 vbias2.n311 vbias2.n305 0.021
R1921 vbias2.n38 vbias2.n37 0.021
R1922 vbias2.n21 vbias2.n20 0.021
R1923 vbias2.n10 vbias2.n9 0.021
R1924 vbias2.n310 vbias2.n309 0.021
R1925 vbias2.n280 vbias2.n279 0.021
R1926 vbias2.n51 vbias2.n50 0.021
R1927 vbias2.n263 vbias2.n262 0.021
R1928 vbias2.n246 vbias2.n245 0.021
R1929 vbias2.n28 vbias2.n27 0.02
R1930 vbias2.n41 vbias2.n40 0.02
R1931 vbias2.n13 vbias2.n12 0.02
R1932 vbias2.n54 vbias2.n53 0.02
R1933 vbias2.n287 vbias2.n286 0.02
R1934 vbias2.n270 vbias2.n269 0.02
R1935 vbias2.n254 vbias2.n253 0.02
R1936 vbias2.n458 vbias2.n457 0.018
R1937 vbias2.n442 vbias2.n441 0.018
R1938 vbias2.n426 vbias2.n425 0.018
R1939 vbias2.n410 vbias2.n409 0.018
R1940 vbias2.n394 vbias2.n393 0.018
R1941 vbias2.n378 vbias2.n377 0.018
R1942 vbias2.n362 vbias2.n361 0.018
R1943 vbias2.n346 vbias2.n345 0.018
R1944 vbias2.n330 vbias2.n329 0.018
R1945 vbias2.n338 vbias2.n337 0.018
R1946 vbias2.n354 vbias2.n353 0.018
R1947 vbias2.n370 vbias2.n369 0.018
R1948 vbias2.n386 vbias2.n385 0.018
R1949 vbias2.n402 vbias2.n401 0.018
R1950 vbias2.n418 vbias2.n417 0.018
R1951 vbias2.n434 vbias2.n433 0.018
R1952 vbias2.n450 vbias2.n449 0.018
R1953 vbias2.n322 vbias2.n321 0.018
R1954 vbias2.n296 vbias2.n14 0.014
R1955 vbias2.n272 vbias2.n271 0.014
R1956 vbias2.n227 vbias2.n226 0.014
R1957 vbias2.n218 vbias2.n217 0.014
R1958 vbias2.n209 vbias2.n208 0.014
R1959 vbias2.n200 vbias2.n199 0.014
R1960 vbias2.n191 vbias2.n190 0.014
R1961 vbias2.n182 vbias2.n181 0.014
R1962 vbias2.n173 vbias2.n172 0.014
R1963 vbias2.n164 vbias2.n163 0.014
R1964 vbias2.n155 vbias2.n154 0.014
R1965 vbias2.n146 vbias2.n145 0.014
R1966 vbias2.n137 vbias2.n136 0.014
R1967 vbias2.n128 vbias2.n127 0.014
R1968 vbias2.n119 vbias2.n118 0.014
R1969 vbias2.n110 vbias2.n109 0.014
R1970 vbias2.n101 vbias2.n100 0.014
R1971 vbias2.n92 vbias2.n91 0.014
R1972 vbias2.n83 vbias2.n82 0.014
R1973 vbias2.n74 vbias2.n73 0.014
R1974 vbias2.n65 vbias2.n62 0.014
R1975 vbias2.n303 vbias2.n302 0.006
R1976 vbias2.n7 vbias2.n6 0.006
R1977 vbias2.n25 vbias2.n24 0.006
R1978 vbias2.n35 vbias2.n34 0.006
R1979 vbias2.n251 vbias2.n250 0.006
R1980 vbias2.n267 vbias2.n266 0.006
R1981 vbias2.n48 vbias2.n47 0.006
R1982 vbias2.n284 vbias2.n283 0.006
R1983 vbias2.n312 vbias2.n311 0.006
R1984 vbias2.n331 vbias2.n330 0.006
R1985 vbias2.n339 vbias2.n338 0.006
R1986 vbias2.n347 vbias2.n346 0.006
R1987 vbias2.n355 vbias2.n354 0.006
R1988 vbias2.n363 vbias2.n362 0.006
R1989 vbias2.n371 vbias2.n370 0.006
R1990 vbias2.n379 vbias2.n378 0.006
R1991 vbias2.n387 vbias2.n386 0.006
R1992 vbias2.n395 vbias2.n394 0.006
R1993 vbias2.n403 vbias2.n402 0.006
R1994 vbias2.n411 vbias2.n410 0.006
R1995 vbias2.n419 vbias2.n418 0.006
R1996 vbias2.n427 vbias2.n426 0.006
R1997 vbias2.n435 vbias2.n434 0.006
R1998 vbias2.n443 vbias2.n442 0.006
R1999 vbias2.n451 vbias2.n450 0.006
R2000 vbias2.n459 vbias2.n458 0.006
R2001 vbias2.n323 vbias2.n322 0.006
R2002 vbias2.n72 vbias2.n71 0.006
R2003 vbias2.n81 vbias2.n80 0.006
R2004 vbias2.n90 vbias2.n89 0.006
R2005 vbias2.n99 vbias2.n98 0.006
R2006 vbias2.n108 vbias2.n107 0.006
R2007 vbias2.n117 vbias2.n116 0.006
R2008 vbias2.n126 vbias2.n125 0.006
R2009 vbias2.n135 vbias2.n134 0.006
R2010 vbias2.n144 vbias2.n143 0.006
R2011 vbias2.n153 vbias2.n152 0.006
R2012 vbias2.n162 vbias2.n161 0.006
R2013 vbias2.n171 vbias2.n170 0.006
R2014 vbias2.n180 vbias2.n179 0.006
R2015 vbias2.n189 vbias2.n188 0.006
R2016 vbias2.n198 vbias2.n197 0.006
R2017 vbias2.n207 vbias2.n206 0.006
R2018 vbias2.n216 vbias2.n215 0.006
R2019 vbias2.n225 vbias2.n224 0.006
R2020 vbias2.n27 vbias2.n26 0.002
R2021 vbias2.n309 vbias2.n308 0.002
R2022 vbias2.n40 vbias2.n39 0.002
R2023 vbias2.n37 vbias2.n36 0.002
R2024 vbias2.n20 vbias2.n19 0.002
R2025 vbias2.n12 vbias2.n11 0.002
R2026 vbias2.n9 vbias2.n8 0.002
R2027 vbias2.n305 vbias2.n304 0.002
R2028 vbias2.n53 vbias2.n52 0.002
R2029 vbias2.n479 vbias2.n478 0.002
R2030 vbias2.n286 vbias2.n285 0.002
R2031 vbias2.n279 vbias2.n278 0.002
R2032 vbias2.n50 vbias2.n49 0.002
R2033 vbias2.n269 vbias2.n268 0.002
R2034 vbias2.n262 vbias2.n261 0.002
R2035 vbias2.n253 vbias2.n252 0.002
R2036 vbias2.n245 vbias2.n244 0.002
R2037 vbias2.n480 vbias2.n479 0.001
R2038 vbias2.n294 vbias2.n287 0.001
R2039 vbias2.n297 vbias2.n13 0.001
R2040 vbias2.n295 vbias2.n41 0.001
R2041 vbias2.n296 vbias2.n28 0.001
R2042 vbias2.n272 vbias2.n270 0.001
R2043 vbias2.n255 vbias2.n254 0.001
R2044 vbias2.n273 vbias2.n54 0.001
R2045 vbias2.n318 vbias2.n317 0.001
R2046 vbias2.n333 vbias2.n332 0.001
R2047 vbias2.n341 vbias2.n340 0.001
R2048 vbias2.n349 vbias2.n348 0.001
R2049 vbias2.n357 vbias2.n356 0.001
R2050 vbias2.n365 vbias2.n364 0.001
R2051 vbias2.n373 vbias2.n372 0.001
R2052 vbias2.n381 vbias2.n380 0.001
R2053 vbias2.n389 vbias2.n388 0.001
R2054 vbias2.n397 vbias2.n396 0.001
R2055 vbias2.n405 vbias2.n404 0.001
R2056 vbias2.n413 vbias2.n412 0.001
R2057 vbias2.n421 vbias2.n420 0.001
R2058 vbias2.n429 vbias2.n428 0.001
R2059 vbias2.n437 vbias2.n436 0.001
R2060 vbias2.n445 vbias2.n444 0.001
R2061 vbias2.n453 vbias2.n452 0.001
R2062 vbias2.n461 vbias2.n460 0.001
R2063 vbias2.n469 vbias2.n468 0.001
R2064 vbias2.n523 vbias2.n522 0.001
R2065 vbias2.n325 vbias2.n324 0.001
R2066 vbias2.n521 vbias2.n520 0.001
R2067 vbias2.n57 vbias2.n56 0.001
R2068 vbias2.n68 vbias2.n67 0.001
R2069 vbias2.n77 vbias2.n76 0.001
R2070 vbias2.n86 vbias2.n85 0.001
R2071 vbias2.n95 vbias2.n94 0.001
R2072 vbias2.n104 vbias2.n103 0.001
R2073 vbias2.n113 vbias2.n112 0.001
R2074 vbias2.n122 vbias2.n121 0.001
R2075 vbias2.n131 vbias2.n130 0.001
R2076 vbias2.n140 vbias2.n139 0.001
R2077 vbias2.n149 vbias2.n148 0.001
R2078 vbias2.n158 vbias2.n157 0.001
R2079 vbias2.n167 vbias2.n166 0.001
R2080 vbias2.n176 vbias2.n175 0.001
R2081 vbias2.n185 vbias2.n184 0.001
R2082 vbias2.n194 vbias2.n193 0.001
R2083 vbias2.n203 vbias2.n202 0.001
R2084 vbias2.n212 vbias2.n211 0.001
R2085 vbias2.n221 vbias2.n220 0.001
R2086 vbias2 vbias2.n523 0.001
R2087 vbias2.n60 vbias2.n59 0.001
R2088 vbias2.n466 vbias2.n465 0.001
R2089 vbias2.n311 vbias2.n310 0.001
R2090 vbias2.n54 vbias2.n51 0.001
R2091 vbias2.n28 vbias2.n21 0.001
R2092 vbias2.n41 vbias2.n38 0.001
R2093 vbias2.n13 vbias2.n10 0.001
R2094 vbias2.n287 vbias2.n280 0.001
R2095 vbias2.n270 vbias2.n263 0.001
R2096 vbias2.n254 vbias2.n246 0.001
R2097 vbias2.n228 vbias2.n227 0.001
R2098 vbias2.n481 vbias2.n480 0.001
R2099 vbias2.n484 vbias2.n476 0.001
R2100 vbias2.n487 vbias2.n486 0.001
R2101 vbias2.n497 vbias2.n496 0.001
R2102 vbias2.n493 vbias2.n471 0.001
R2103 vbias2.n492 vbias2.n491 0.001
R2104 vbias2.n489 vbias2.n474 0.001
R2105 vbias2.n243 vbias2.n242 0.001
R2106 vbias2.n223 vbias2.n222 0.001
R2107 vbias2.n205 vbias2.n204 0.001
R2108 vbias2.n187 vbias2.n186 0.001
R2109 vbias2.n169 vbias2.n168 0.001
R2110 vbias2.n151 vbias2.n150 0.001
R2111 vbias2.n133 vbias2.n132 0.001
R2112 vbias2.n115 vbias2.n114 0.001
R2113 vbias2.n97 vbias2.n96 0.001
R2114 vbias2.n79 vbias2.n78 0.001
R2115 vbias2.n59 vbias2.n58 0.001
R2116 vbias2.n70 vbias2.n69 0.001
R2117 vbias2.n88 vbias2.n87 0.001
R2118 vbias2.n106 vbias2.n105 0.001
R2119 vbias2.n124 vbias2.n123 0.001
R2120 vbias2.n142 vbias2.n141 0.001
R2121 vbias2.n160 vbias2.n159 0.001
R2122 vbias2.n178 vbias2.n177 0.001
R2123 vbias2.n196 vbias2.n195 0.001
R2124 vbias2.n214 vbias2.n213 0.001
R2125 vbias2.n282 vbias2.n281 0.001
R2126 vbias2.n46 vbias2.n45 0.001
R2127 vbias2.n265 vbias2.n264 0.001
R2128 vbias2.n23 vbias2.n22 0.001
R2129 vbias2.n5 vbias2.n4 0.001
R2130 vbias2.n301 vbias2.n300 0.001
R2131 vbias2.n457 vbias2.n456 0.001
R2132 vbias2.n441 vbias2.n440 0.001
R2133 vbias2.n425 vbias2.n424 0.001
R2134 vbias2.n409 vbias2.n408 0.001
R2135 vbias2.n393 vbias2.n392 0.001
R2136 vbias2.n377 vbias2.n376 0.001
R2137 vbias2.n361 vbias2.n360 0.001
R2138 vbias2.n345 vbias2.n344 0.001
R2139 vbias2.n329 vbias2.n328 0.001
R2140 vbias2.n337 vbias2.n336 0.001
R2141 vbias2.n353 vbias2.n352 0.001
R2142 vbias2.n369 vbias2.n368 0.001
R2143 vbias2.n385 vbias2.n384 0.001
R2144 vbias2.n401 vbias2.n400 0.001
R2145 vbias2.n417 vbias2.n416 0.001
R2146 vbias2.n433 vbias2.n432 0.001
R2147 vbias2.n449 vbias2.n448 0.001
R2148 vbias2.n465 vbias2.n464 0.001
R2149 vbias2.n33 vbias2.n32 0.001
R2150 vbias2.n483 vbias2.n482 0.001
R2151 vbias2.n248 vbias2.n247 0.001
R2152 vbias2.n321 vbias2.n320 0.001
R2153 vbias2.n483 vbias2.n481 0.001
R2154 vdd.n210 vdd.n209 13465.4
R2155 vdd.n164 vdd.n159 380.99
R2156 vdd.n210 vdd.n205 344.236
R2157 vdd.n209 vdd.n115 344.236
R2158 vdd.n119 vdd.n115 344.236
R2159 vdd.n131 vdd.n127 344.236
R2160 vdd.n135 vdd.n131 344.236
R2161 vdd.n142 vdd.n135 344.236
R2162 vdd.n143 vdd.n142 344.236
R2163 vdd.n147 vdd.n143 344.236
R2164 vdd.n151 vdd.n147 344.236
R2165 vdd.n173 vdd.n169 344.236
R2166 vdd.n177 vdd.n173 344.236
R2167 vdd.n181 vdd.n177 344.236
R2168 vdd.n185 vdd.n181 344.236
R2169 vdd.n189 vdd.n185 344.236
R2170 vdd.n193 vdd.n189 344.236
R2171 vdd.n197 vdd.n193 344.236
R2172 vdd.n201 vdd.n197 344.236
R2173 vdd.n205 vdd.n201 344.236
R2174 vdd.n79 vdd.n78 344.236
R2175 vdd.n126 vdd.n119 341.409
R2176 vdd.n127 vdd.n126 340.106
R2177 vdd.n94 vdd.n93 340.106
R2178 vdd.n169 vdd.n168 327.477
R2179 vdd.n167 vdd.n151 326.862
R2180 vdd.n168 vdd.n167 308.856
R2181 vdd.n208 vdd.t230 7.146
R2182 vdd.n208 vdd.t283 7.146
R2183 vdd.n207 vdd.t225 7.146
R2184 vdd.n207 vdd.t278 7.146
R2185 vdd.n206 vdd.t262 7.146
R2186 vdd.n206 vdd.t279 7.146
R2187 vdd.n204 vdd.t238 7.146
R2188 vdd.n204 vdd.t199 7.146
R2189 vdd.n203 vdd.t234 7.146
R2190 vdd.n203 vdd.t285 7.146
R2191 vdd.n202 vdd.t223 7.146
R2192 vdd.n202 vdd.t152 7.146
R2193 vdd.n200 vdd.t254 7.146
R2194 vdd.n200 vdd.t266 7.146
R2195 vdd.n199 vdd.t248 7.146
R2196 vdd.n199 vdd.t263 7.146
R2197 vdd.n198 vdd.t184 7.146
R2198 vdd.n198 vdd.t209 7.146
R2199 vdd.n196 vdd.t161 7.146
R2200 vdd.n196 vdd.t271 7.146
R2201 vdd.n195 vdd.t157 7.146
R2202 vdd.n195 vdd.t268 7.146
R2203 vdd.n194 vdd.t146 7.146
R2204 vdd.n194 vdd.t188 7.146
R2205 vdd.n192 vdd.t168 7.146
R2206 vdd.n192 vdd.t160 7.146
R2207 vdd.n191 vdd.t164 7.146
R2208 vdd.n191 vdd.t154 7.146
R2209 vdd.n190 vdd.t270 7.146
R2210 vdd.n190 vdd.t193 7.146
R2211 vdd.n188 vdd.t175 7.146
R2212 vdd.n188 vdd.t227 7.146
R2213 vdd.n187 vdd.t169 7.146
R2214 vdd.n187 vdd.t220 7.146
R2215 vdd.n186 vdd.t214 7.146
R2216 vdd.n186 vdd.t149 7.146
R2217 vdd.n184 vdd.t185 7.146
R2218 vdd.n184 vdd.t237 7.146
R2219 vdd.n183 vdd.t178 7.146
R2220 vdd.n183 vdd.t229 7.146
R2221 vdd.n182 vdd.t253 7.146
R2222 vdd.n182 vdd.t274 7.146
R2223 vdd.n180 vdd.t275 7.146
R2224 vdd.n180 vdd.t286 7.146
R2225 vdd.n179 vdd.t273 7.146
R2226 vdd.n179 vdd.t281 7.146
R2227 vdd.n178 vdd.t159 7.146
R2228 vdd.n178 vdd.t201 7.146
R2229 vdd.n176 vdd.t249 7.146
R2230 vdd.n176 vdd.t231 7.146
R2231 vdd.n175 vdd.t189 7.146
R2232 vdd.n175 vdd.t224 7.146
R2233 vdd.n174 vdd.t216 7.146
R2234 vdd.n174 vdd.t210 7.146
R2235 vdd.n172 vdd.t145 7.146
R2236 vdd.n172 vdd.t239 7.146
R2237 vdd.n171 vdd.t144 7.146
R2238 vdd.n171 vdd.t233 7.146
R2239 vdd.n170 vdd.t247 7.146
R2240 vdd.n170 vdd.t191 7.146
R2241 vdd.n154 vdd.t272 7.146
R2242 vdd.n154 vdd.t243 7.146
R2243 vdd.n153 vdd.t269 7.146
R2244 vdd.n153 vdd.t244 7.146
R2245 vdd.n152 vdd.t203 7.146
R2246 vdd.n152 vdd.t195 7.146
R2247 vdd.n150 vdd.t217 7.146
R2248 vdd.n150 vdd.t176 7.146
R2249 vdd.n149 vdd.t211 7.146
R2250 vdd.n149 vdd.t171 7.146
R2251 vdd.n148 vdd.t236 7.146
R2252 vdd.n148 vdd.t182 7.146
R2253 vdd.n146 vdd.t228 7.146
R2254 vdd.n146 vdd.t186 7.146
R2255 vdd.n145 vdd.t219 7.146
R2256 vdd.n145 vdd.t179 7.146
R2257 vdd.n144 vdd.t265 7.146
R2258 vdd.n144 vdd.t207 7.146
R2259 vdd.n141 vdd.t204 7.146
R2260 vdd.n141 vdd.t187 7.146
R2261 vdd.n140 vdd.t200 7.146
R2262 vdd.n140 vdd.t181 7.146
R2263 vdd.n139 vdd.t165 7.146
R2264 vdd.n139 vdd.t208 7.146
R2265 vdd.n138 vdd.t287 7.146
R2266 vdd.n138 vdd.t250 7.146
R2267 vdd.n137 vdd.t280 7.146
R2268 vdd.n137 vdd.t190 7.146
R2269 vdd.n136 vdd.t151 7.146
R2270 vdd.n136 vdd.t183 7.146
R2271 vdd.n134 vdd.t232 7.146
R2272 vdd.n134 vdd.t256 7.146
R2273 vdd.n133 vdd.t226 7.146
R2274 vdd.n133 vdd.t251 7.146
R2275 vdd.n132 vdd.t174 7.146
R2276 vdd.n132 vdd.t196 7.146
R2277 vdd.n130 vdd.t205 7.146
R2278 vdd.n130 vdd.t261 7.146
R2279 vdd.n129 vdd.t202 7.146
R2280 vdd.n129 vdd.t257 7.146
R2281 vdd.n128 vdd.t235 7.146
R2282 vdd.n128 vdd.t158 7.146
R2283 vdd.n125 vdd.t155 7.146
R2284 vdd.n125 vdd.t267 7.146
R2285 vdd.n124 vdd.t150 7.146
R2286 vdd.n124 vdd.t264 7.146
R2287 vdd.n123 vdd.t192 7.146
R2288 vdd.n123 vdd.t282 7.146
R2289 vdd.n122 vdd.t221 7.146
R2290 vdd.n122 vdd.t180 7.146
R2291 vdd.n121 vdd.t213 7.146
R2292 vdd.n121 vdd.t172 7.146
R2293 vdd.n120 vdd.t148 7.146
R2294 vdd.n120 vdd.t252 7.146
R2295 vdd.n118 vdd.t167 7.146
R2296 vdd.n118 vdd.t218 7.146
R2297 vdd.n117 vdd.t163 7.146
R2298 vdd.n117 vdd.t212 7.146
R2299 vdd.n116 vdd.t166 7.146
R2300 vdd.n116 vdd.t255 7.146
R2301 vdd.n113 vdd.t177 7.146
R2302 vdd.n113 vdd.t198 7.146
R2303 vdd.n112 vdd.t170 7.146
R2304 vdd.n112 vdd.t284 7.146
R2305 vdd.n111 vdd.t197 7.146
R2306 vdd.n111 vdd.t153 7.146
R2307 vdd.n157 vdd.t240 7.146
R2308 vdd.n157 vdd.t162 7.146
R2309 vdd.n156 vdd.t241 7.146
R2310 vdd.n156 vdd.t156 7.146
R2311 vdd.n155 vdd.t242 7.146
R2312 vdd.n155 vdd.t259 7.146
R2313 vdd.n162 vdd.t260 7.146
R2314 vdd.n162 vdd.t245 7.146
R2315 vdd.n161 vdd.t258 7.146
R2316 vdd.n161 vdd.t246 7.146
R2317 vdd.n160 vdd.t206 7.146
R2318 vdd.n160 vdd.t194 7.146
R2319 vdd.n213 vdd.t222 7.146
R2320 vdd.n213 vdd.t277 7.146
R2321 vdd.n212 vdd.t215 7.146
R2322 vdd.n212 vdd.t276 7.146
R2323 vdd.n211 vdd.t147 7.146
R2324 vdd.n211 vdd.t173 7.146
R2325 vdd.n3 vdd.t13 7.146
R2326 vdd.n3 vdd.t126 7.146
R2327 vdd.n2 vdd.t21 7.146
R2328 vdd.n2 vdd.t133 7.146
R2329 vdd.n1 vdd.t27 7.146
R2330 vdd.n1 vdd.t138 7.146
R2331 vdd.n6 vdd.t89 7.146
R2332 vdd.n6 vdd.t76 7.146
R2333 vdd.n5 vdd.t93 7.146
R2334 vdd.n5 vdd.t80 7.146
R2335 vdd.n4 vdd.t97 7.146
R2336 vdd.n4 vdd.t82 7.146
R2337 vdd.n12 vdd.t34 7.146
R2338 vdd.n12 vdd.t4 7.146
R2339 vdd.n11 vdd.t40 7.146
R2340 vdd.n11 vdd.t12 7.146
R2341 vdd.n10 vdd.t44 7.146
R2342 vdd.n10 vdd.t16 7.146
R2343 vdd.n15 vdd.t113 7.146
R2344 vdd.n15 vdd.t46 7.146
R2345 vdd.n14 vdd.t120 7.146
R2346 vdd.n14 vdd.t52 7.146
R2347 vdd.n13 vdd.t130 7.146
R2348 vdd.n13 vdd.t57 7.146
R2349 vdd.n21 vdd.t20 7.146
R2350 vdd.n21 vdd.t108 7.146
R2351 vdd.n20 vdd.t26 7.146
R2352 vdd.n20 vdd.t117 7.146
R2353 vdd.n19 vdd.t31 7.146
R2354 vdd.n19 vdd.t125 7.146
R2355 vdd.n24 vdd.t85 7.146
R2356 vdd.n24 vdd.t102 7.146
R2357 vdd.n23 vdd.t88 7.146
R2358 vdd.n23 vdd.t110 7.146
R2359 vdd.n22 vdd.t91 7.146
R2360 vdd.n22 vdd.t119 7.146
R2361 vdd.n30 vdd.t39 7.146
R2362 vdd.n30 vdd.t10 7.146
R2363 vdd.n29 vdd.t43 7.146
R2364 vdd.n29 vdd.t18 7.146
R2365 vdd.n28 vdd.t48 7.146
R2366 vdd.n28 vdd.t23 7.146
R2367 vdd.n33 vdd.t98 7.146
R2368 vdd.n33 vdd.t83 7.146
R2369 vdd.n32 vdd.t105 7.146
R2370 vdd.n32 vdd.t84 7.146
R2371 vdd.n31 vdd.t112 7.146
R2372 vdd.n31 vdd.t86 7.146
R2373 vdd.n39 vdd.t141 7.146
R2374 vdd.n39 vdd.t64 7.146
R2375 vdd.n38 vdd.t1 7.146
R2376 vdd.n38 vdd.t70 7.146
R2377 vdd.n37 vdd.t6 7.146
R2378 vdd.n37 vdd.t75 7.146
R2379 vdd.n42 vdd.t38 7.146
R2380 vdd.n42 vdd.t45 7.146
R2381 vdd.n41 vdd.t42 7.146
R2382 vdd.n41 vdd.t51 7.146
R2383 vdd.n40 vdd.t47 7.146
R2384 vdd.n40 vdd.t55 7.146
R2385 vdd.n48 vdd.t19 7.146
R2386 vdd.n48 vdd.t106 7.146
R2387 vdd.n47 vdd.t25 7.146
R2388 vdd.n47 vdd.t116 7.146
R2389 vdd.n46 vdd.t29 7.146
R2390 vdd.n46 vdd.t123 7.146
R2391 vdd.n65 vdd.t63 7.146
R2392 vdd.n65 vdd.t50 7.146
R2393 vdd.n64 vdd.t69 7.146
R2394 vdd.n64 vdd.t53 7.146
R2395 vdd.n63 vdd.t73 7.146
R2396 vdd.n63 vdd.t60 7.146
R2397 vdd.n71 vdd.t24 7.146
R2398 vdd.n71 vdd.t115 7.146
R2399 vdd.n70 vdd.t30 7.146
R2400 vdd.n70 vdd.t121 7.146
R2401 vdd.n69 vdd.t35 7.146
R2402 vdd.n69 vdd.t129 7.146
R2403 vdd.n74 vdd.t87 7.146
R2404 vdd.n74 vdd.t56 7.146
R2405 vdd.n73 vdd.t90 7.146
R2406 vdd.n73 vdd.t61 7.146
R2407 vdd.n72 vdd.t94 7.146
R2408 vdd.n72 vdd.t65 7.146
R2409 vdd.n77 vdd.t135 7.146
R2410 vdd.n77 vdd.t49 7.146
R2411 vdd.n76 vdd.t139 7.146
R2412 vdd.n76 vdd.t54 7.146
R2413 vdd.n75 vdd.t0 7.146
R2414 vdd.n75 vdd.t59 7.146
R2415 vdd.n84 vdd.t5 7.146
R2416 vdd.n84 vdd.t114 7.146
R2417 vdd.n83 vdd.t9 7.146
R2418 vdd.n83 vdd.t122 7.146
R2419 vdd.n82 vdd.t15 7.146
R2420 vdd.n82 vdd.t128 7.146
R2421 vdd.n87 vdd.t124 7.146
R2422 vdd.n87 vdd.t68 7.146
R2423 vdd.n86 vdd.t131 7.146
R2424 vdd.n86 vdd.t72 7.146
R2425 vdd.n85 vdd.t137 7.146
R2426 vdd.n85 vdd.t78 7.146
R2427 vdd.n97 vdd.t28 7.146
R2428 vdd.n97 vdd.t142 7.146
R2429 vdd.n96 vdd.t32 7.146
R2430 vdd.n96 vdd.t2 7.146
R2431 vdd.n95 vdd.t37 7.146
R2432 vdd.n95 vdd.t8 7.146
R2433 vdd.n92 vdd.t103 7.146
R2434 vdd.n92 vdd.t74 7.146
R2435 vdd.n91 vdd.t109 7.146
R2436 vdd.n91 vdd.t79 7.146
R2437 vdd.n90 vdd.t118 7.146
R2438 vdd.n90 vdd.t81 7.146
R2439 vdd.n100 vdd.t11 7.146
R2440 vdd.n100 vdd.t99 7.146
R2441 vdd.n99 vdd.t17 7.146
R2442 vdd.n99 vdd.t104 7.146
R2443 vdd.n98 vdd.t22 7.146
R2444 vdd.n98 vdd.t111 7.146
R2445 vdd.n106 vdd.t132 7.146
R2446 vdd.n106 vdd.t95 7.146
R2447 vdd.n105 vdd.t136 7.146
R2448 vdd.n105 vdd.t100 7.146
R2449 vdd.n104 vdd.t143 7.146
R2450 vdd.n104 vdd.t107 7.146
R2451 vdd.n58 vdd.t127 7.146
R2452 vdd.n58 vdd.t92 7.146
R2453 vdd.n57 vdd.t134 7.146
R2454 vdd.n57 vdd.t96 7.146
R2455 vdd.n56 vdd.t140 7.146
R2456 vdd.n56 vdd.t101 7.146
R2457 vdd.n51 vdd.t58 7.146
R2458 vdd.n51 vdd.t33 7.146
R2459 vdd.n50 vdd.t62 7.146
R2460 vdd.n50 vdd.t36 7.146
R2461 vdd.n49 vdd.t67 7.146
R2462 vdd.n49 vdd.t41 7.146
R2463 vdd.n110 vdd.t66 7.146
R2464 vdd.n110 vdd.t3 7.146
R2465 vdd.n109 vdd.t71 7.146
R2466 vdd.n109 vdd.t7 7.146
R2467 vdd.n108 vdd.t77 7.146
R2468 vdd.n108 vdd.t14 7.146
R2469 vdd.n158 vdd.n157 0.916
R2470 vdd.n163 vdd.n162 0.916
R2471 vdd.n59 vdd.n58 0.916
R2472 vdd.n52 vdd.n51 0.916
R2473 vdd.n215 vdd.n208 0.898
R2474 vdd.n216 vdd.n204 0.898
R2475 vdd.n217 vdd.n200 0.898
R2476 vdd.n218 vdd.n196 0.898
R2477 vdd.n219 vdd.n192 0.898
R2478 vdd.n220 vdd.n188 0.898
R2479 vdd.n221 vdd.n184 0.898
R2480 vdd.n222 vdd.n180 0.898
R2481 vdd.n223 vdd.n176 0.898
R2482 vdd.n224 vdd.n172 0.898
R2483 vdd.n227 vdd.n154 0.898
R2484 vdd.n228 vdd.n150 0.898
R2485 vdd.n229 vdd.n146 0.898
R2486 vdd.n230 vdd.n138 0.898
R2487 vdd.n231 vdd.n134 0.898
R2488 vdd.n232 vdd.n130 0.898
R2489 vdd.n233 vdd.n122 0.898
R2490 vdd.n234 vdd.n118 0.898
R2491 vdd.n114 vdd.n113 0.898
R2492 vdd.n214 vdd.n213 0.898
R2493 vdd.n257 vdd.n3 0.898
R2494 vdd.n8 vdd.n6 0.898
R2495 vdd.n255 vdd.n12 0.898
R2496 vdd.n17 vdd.n15 0.898
R2497 vdd.n253 vdd.n21 0.898
R2498 vdd.n26 vdd.n24 0.898
R2499 vdd.n251 vdd.n30 0.898
R2500 vdd.n35 vdd.n33 0.898
R2501 vdd.n249 vdd.n39 0.898
R2502 vdd.n44 vdd.n42 0.898
R2503 vdd.n247 vdd.n48 0.898
R2504 vdd.n67 vdd.n65 0.898
R2505 vdd.n243 vdd.n71 0.898
R2506 vdd.n80 vdd.n74 0.898
R2507 vdd.n241 vdd.n84 0.898
R2508 vdd.n89 vdd.n87 0.898
R2509 vdd.n239 vdd.n97 0.898
R2510 vdd.n102 vdd.n100 0.898
R2511 vdd.n237 vdd.n106 0.898
R2512 vdd.n236 vdd.n110 0.898
R2513 vdd.n142 vdd.n141 0.884
R2514 vdd.n78 vdd.n77 0.884
R2515 vdd.n126 vdd.n125 0.882
R2516 vdd.n93 vdd.n92 0.882
R2517 vdd.n207 vdd.n206 0.865
R2518 vdd.n208 vdd.n207 0.865
R2519 vdd.n203 vdd.n202 0.865
R2520 vdd.n204 vdd.n203 0.865
R2521 vdd.n199 vdd.n198 0.865
R2522 vdd.n200 vdd.n199 0.865
R2523 vdd.n195 vdd.n194 0.865
R2524 vdd.n196 vdd.n195 0.865
R2525 vdd.n191 vdd.n190 0.865
R2526 vdd.n192 vdd.n191 0.865
R2527 vdd.n187 vdd.n186 0.865
R2528 vdd.n188 vdd.n187 0.865
R2529 vdd.n183 vdd.n182 0.865
R2530 vdd.n184 vdd.n183 0.865
R2531 vdd.n179 vdd.n178 0.865
R2532 vdd.n180 vdd.n179 0.865
R2533 vdd.n175 vdd.n174 0.865
R2534 vdd.n176 vdd.n175 0.865
R2535 vdd.n171 vdd.n170 0.865
R2536 vdd.n172 vdd.n171 0.865
R2537 vdd.n153 vdd.n152 0.865
R2538 vdd.n154 vdd.n153 0.865
R2539 vdd.n149 vdd.n148 0.865
R2540 vdd.n150 vdd.n149 0.865
R2541 vdd.n145 vdd.n144 0.865
R2542 vdd.n146 vdd.n145 0.865
R2543 vdd.n140 vdd.n139 0.865
R2544 vdd.n141 vdd.n140 0.865
R2545 vdd.n137 vdd.n136 0.865
R2546 vdd.n138 vdd.n137 0.865
R2547 vdd.n133 vdd.n132 0.865
R2548 vdd.n134 vdd.n133 0.865
R2549 vdd.n129 vdd.n128 0.865
R2550 vdd.n130 vdd.n129 0.865
R2551 vdd.n124 vdd.n123 0.865
R2552 vdd.n125 vdd.n124 0.865
R2553 vdd.n121 vdd.n120 0.865
R2554 vdd.n122 vdd.n121 0.865
R2555 vdd.n117 vdd.n116 0.865
R2556 vdd.n118 vdd.n117 0.865
R2557 vdd.n112 vdd.n111 0.865
R2558 vdd.n113 vdd.n112 0.865
R2559 vdd.n156 vdd.n155 0.865
R2560 vdd.n157 vdd.n156 0.865
R2561 vdd.n161 vdd.n160 0.865
R2562 vdd.n162 vdd.n161 0.865
R2563 vdd.n212 vdd.n211 0.865
R2564 vdd.n213 vdd.n212 0.865
R2565 vdd.n2 vdd.n1 0.865
R2566 vdd.n3 vdd.n2 0.865
R2567 vdd.n5 vdd.n4 0.865
R2568 vdd.n6 vdd.n5 0.865
R2569 vdd.n11 vdd.n10 0.865
R2570 vdd.n12 vdd.n11 0.865
R2571 vdd.n14 vdd.n13 0.865
R2572 vdd.n15 vdd.n14 0.865
R2573 vdd.n20 vdd.n19 0.865
R2574 vdd.n21 vdd.n20 0.865
R2575 vdd.n23 vdd.n22 0.865
R2576 vdd.n24 vdd.n23 0.865
R2577 vdd.n29 vdd.n28 0.865
R2578 vdd.n30 vdd.n29 0.865
R2579 vdd.n32 vdd.n31 0.865
R2580 vdd.n33 vdd.n32 0.865
R2581 vdd.n38 vdd.n37 0.865
R2582 vdd.n39 vdd.n38 0.865
R2583 vdd.n41 vdd.n40 0.865
R2584 vdd.n42 vdd.n41 0.865
R2585 vdd.n47 vdd.n46 0.865
R2586 vdd.n48 vdd.n47 0.865
R2587 vdd.n64 vdd.n63 0.865
R2588 vdd.n65 vdd.n64 0.865
R2589 vdd.n70 vdd.n69 0.865
R2590 vdd.n71 vdd.n70 0.865
R2591 vdd.n73 vdd.n72 0.865
R2592 vdd.n74 vdd.n73 0.865
R2593 vdd.n76 vdd.n75 0.865
R2594 vdd.n77 vdd.n76 0.865
R2595 vdd.n83 vdd.n82 0.865
R2596 vdd.n84 vdd.n83 0.865
R2597 vdd.n86 vdd.n85 0.865
R2598 vdd.n87 vdd.n86 0.865
R2599 vdd.n96 vdd.n95 0.865
R2600 vdd.n97 vdd.n96 0.865
R2601 vdd.n91 vdd.n90 0.865
R2602 vdd.n92 vdd.n91 0.865
R2603 vdd.n99 vdd.n98 0.865
R2604 vdd.n100 vdd.n99 0.865
R2605 vdd.n105 vdd.n104 0.865
R2606 vdd.n106 vdd.n105 0.865
R2607 vdd.n57 vdd.n56 0.865
R2608 vdd.n58 vdd.n57 0.865
R2609 vdd.n50 vdd.n49 0.865
R2610 vdd.n51 vdd.n50 0.865
R2611 vdd.n109 vdd.n108 0.865
R2612 vdd.n110 vdd.n109 0.865
R2613 vdd.n236 vdd 0.682
R2614 vdd.n166 vdd.n158 0.5
R2615 vdd.n165 vdd.n163 0.5
R2616 vdd vdd.n235 0.115
R2617 vdd.n233 vdd.n232 0.072
R2618 vdd.n230 vdd.n229 0.072
R2619 vdd.n239 vdd.n238 0.072
R2620 vdd.n242 vdd.n241 0.072
R2621 vdd.n214 vdd 0.059
R2622 vdd.n226 vdd.n159 0.05
R2623 vdd.n225 vdd.n164 0.05
R2624 vdd.n245 vdd.n62 0.05
R2625 vdd.n246 vdd.n55 0.05
R2626 vdd vdd.n257 0.05
R2627 vdd.n235 vdd.n234 0.036
R2628 vdd.n234 vdd.n233 0.036
R2629 vdd.n232 vdd.n231 0.036
R2630 vdd.n231 vdd.n230 0.036
R2631 vdd.n229 vdd.n228 0.036
R2632 vdd.n228 vdd.n227 0.036
R2633 vdd.n227 vdd.n226 0.036
R2634 vdd.n226 vdd.n225 0.036
R2635 vdd.n225 vdd.n224 0.036
R2636 vdd.n224 vdd.n223 0.036
R2637 vdd.n223 vdd.n222 0.036
R2638 vdd.n222 vdd.n221 0.036
R2639 vdd.n221 vdd.n220 0.036
R2640 vdd.n220 vdd.n219 0.036
R2641 vdd.n219 vdd.n218 0.036
R2642 vdd.n218 vdd.n217 0.036
R2643 vdd.n217 vdd.n216 0.036
R2644 vdd.n216 vdd.n215 0.036
R2645 vdd.n215 vdd.n214 0.036
R2646 vdd.n237 vdd.n236 0.036
R2647 vdd.n238 vdd.n237 0.036
R2648 vdd.n240 vdd.n239 0.036
R2649 vdd.n241 vdd.n240 0.036
R2650 vdd.n243 vdd.n242 0.036
R2651 vdd.n244 vdd.n243 0.036
R2652 vdd.n245 vdd.n244 0.036
R2653 vdd.n246 vdd.n245 0.036
R2654 vdd.n247 vdd.n246 0.036
R2655 vdd.n248 vdd.n247 0.036
R2656 vdd.n249 vdd.n248 0.036
R2657 vdd.n250 vdd.n249 0.036
R2658 vdd.n251 vdd.n250 0.036
R2659 vdd.n252 vdd.n251 0.036
R2660 vdd.n253 vdd.n252 0.036
R2661 vdd.n254 vdd.n253 0.036
R2662 vdd.n255 vdd.n254 0.036
R2663 vdd.n256 vdd.n255 0.036
R2664 vdd.n257 vdd.n256 0.036
R2665 vdd.n235 vdd.n114 0.002
R2666 vdd.n238 vdd.n102 0.002
R2667 vdd.n240 vdd.n89 0.002
R2668 vdd.n242 vdd.n80 0.002
R2669 vdd.n244 vdd.n67 0.002
R2670 vdd.n248 vdd.n44 0.002
R2671 vdd.n250 vdd.n35 0.002
R2672 vdd.n252 vdd.n26 0.002
R2673 vdd.n254 vdd.n17 0.002
R2674 vdd.n256 vdd.n8 0.002
R2675 vdd.n166 vdd.n159 0.001
R2676 vdd.n165 vdd.n164 0.001
R2677 vdd.n62 vdd.n61 0.001
R2678 vdd.n55 vdd.n54 0.001
R2679 vdd.n234 vdd.n115 0.001
R2680 vdd.n231 vdd.n131 0.001
R2681 vdd.n230 vdd.n135 0.001
R2682 vdd.n229 vdd.n143 0.001
R2683 vdd.n228 vdd.n147 0.001
R2684 vdd.n227 vdd.n151 0.001
R2685 vdd.n224 vdd.n169 0.001
R2686 vdd.n223 vdd.n173 0.001
R2687 vdd.n222 vdd.n177 0.001
R2688 vdd.n221 vdd.n181 0.001
R2689 vdd.n220 vdd.n185 0.001
R2690 vdd.n219 vdd.n189 0.001
R2691 vdd.n218 vdd.n193 0.001
R2692 vdd.n217 vdd.n197 0.001
R2693 vdd.n216 vdd.n201 0.001
R2694 vdd.n215 vdd.n205 0.001
R2695 vdd.n237 vdd.n103 0.001
R2696 vdd.n89 vdd.n88 0.001
R2697 vdd.n241 vdd.n81 0.001
R2698 vdd.n80 vdd.n79 0.001
R2699 vdd.n243 vdd.n68 0.001
R2700 vdd.n67 vdd.n66 0.001
R2701 vdd.n247 vdd.n45 0.001
R2702 vdd.n44 vdd.n43 0.001
R2703 vdd.n249 vdd.n36 0.001
R2704 vdd.n35 vdd.n34 0.001
R2705 vdd.n251 vdd.n27 0.001
R2706 vdd.n26 vdd.n25 0.001
R2707 vdd.n253 vdd.n18 0.001
R2708 vdd.n17 vdd.n16 0.001
R2709 vdd.n255 vdd.n9 0.001
R2710 vdd.n8 vdd.n7 0.001
R2711 vdd.n233 vdd.n119 0.001
R2712 vdd.n102 vdd.n101 0.001
R2713 vdd.n232 vdd.n127 0.001
R2714 vdd.n239 vdd.n94 0.001
R2715 vdd.n209 vdd.n114 0.001
R2716 vdd.n236 vdd.n107 0.001
R2717 vdd.n214 vdd.n210 0.001
R2718 vdd.n257 vdd.n0 0.001
R2719 vdd.n168 vdd.n165 0.001
R2720 vdd.n54 vdd.n53 0.001
R2721 vdd.n167 vdd.n166 0.001
R2722 vdd.n61 vdd.n60 0.001
R2723 vdd.n226 vdd.n158 0.001
R2724 vdd.n225 vdd.n163 0.001
R2725 vdd.n245 vdd.n59 0.001
R2726 vdd.n246 vdd.n52 0.001
R2727 vref.n25 vref.t18 348.723
R2728 vref.n25 vref.t21 348.588
R2729 vref.n14 vref.t3 348.416
R2730 vref.n27 vref.t1 348.416
R2731 vref.n15 vref.t15 348.416
R2732 vref.t23 vref.n21 348.416
R2733 vref.t13 vref.n20 348.416
R2734 vref.n24 vref.t11 348.416
R2735 vref.n23 vref.t20 348.416
R2736 vref.t10 vref.n30 348.416
R2737 vref.t2 vref.n29 348.416
R2738 vref.t8 vref.n28 348.416
R2739 vref.n7 vref.t4 347.346
R2740 vref.t20 vref.n22 347.336
R2741 vref.n7 vref.t14 347.211
R2742 vref.n22 vref.t23 347.202
R2743 vref.n9 vref.t0 347.04
R2744 vref.t3 vref.n13 347.039
R2745 vref.t1 vref.n15 347.039
R2746 vref.t15 vref.n14 347.039
R2747 vref.n21 vref.t13 347.039
R2748 vref.n20 vref.t21 347.039
R2749 vref.t18 vref.n24 347.039
R2750 vref.t11 vref.n23 347.039
R2751 vref.n31 vref.t10 347.039
R2752 vref.n30 vref.t2 347.039
R2753 vref.n29 vref.t8 347.039
R2754 vref.n2 vref.t22 347.039
R2755 vref.n38 vref.t6 347.039
R2756 vref.n42 vref.t16 347.039
R2757 vref.n0 vref.t7 347.039
R2758 vref.n8 vref.t12 347.039
R2759 vref.n1 vref.t19 347.039
R2760 vref.n37 vref.t5 347.039
R2761 vref.n39 vref.t17 347.039
R2762 vref.n3 vref.t9 347.039
R2763 vref.n29 vref.n15 24.584
R2764 vref.n30 vref.n14 24.584
R2765 vref.n28 vref.n27 24.584
R2766 vref vref.n34 8.877
R2767 vref.n35 vref 5.333
R2768 vref.n49 vref.n48 1.667
R2769 vref.n17 vref.n16 1.296
R2770 vref.n19 vref.n18 1.296
R2771 vref.n26 vref.n25 1.296
R2772 vref.n22 vref.n13 1.289
R2773 vref.n35 vref.n9 1.232
R2774 vref.n49 vref.n43 1.082
R2775 vref.n36 vref.n6 1.079
R2776 vref.n32 vref.n31 1.058
R2777 vref.n32 vref.n12 0.555
R2778 vref.n33 vref.n11 0.555
R2779 vref.n34 vref.n10 0.555
R2780 vref vref.n49 0.543
R2781 vref.n34 vref.n33 0.509
R2782 vref.n33 vref 0.367
R2783 vref.n24 vref.n17 0.307
R2784 vref.n23 vref.n19 0.307
R2785 vref.n4 vref.n3 0.307
R2786 vref.n40 vref.n39 0.307
R2787 vref.n5 vref.n4 0.246
R2788 vref.n47 vref.n46 0.241
R2789 vref.n41 vref.n40 0.24
R2790 vref.n8 vref.n7 0.236
R2791 vref.n27 vref.n26 0.175
R2792 vref.n18 vref.n14 0.175
R2793 vref.n29 vref.n11 0.175
R2794 vref.n16 vref.n15 0.175
R2795 vref.n30 vref.n12 0.175
R2796 vref.n28 vref.n10 0.175
R2797 vref.n5 vref.n1 0.175
R2798 vref.n6 vref.n0 0.175
R2799 vref.n47 vref.n45 0.175
R2800 vref.n48 vref.n44 0.175
R2801 vref.n20 vref.n17 0.172
R2802 vref.n21 vref.n19 0.172
R2803 vref.n4 vref.n2 0.172
R2804 vref.n40 vref.n38 0.172
R2805 vref.n41 vref.n37 0.166
R2806 vref.n43 vref.n42 0.166
R2807 vref vref.n32 0.141
R2808 vref.n16 vref.n11 0.138
R2809 vref.n18 vref.n12 0.138
R2810 vref.n26 vref.n10 0.138
R2811 vref.n48 vref.n47 0.138
R2812 vref.n6 vref.n5 0.136
R2813 vref.n43 vref.n41 0.136
R2814 vref.n36 vref.n35 0.134
R2815 vref.n9 vref.n8 0.087
R2816 vref.n31 vref.n13 0.086
R2817 vref vref.n36 0.041
R2818 a_23370_8306.n12 a_23370_8306.t21 8.207
R2819 a_23370_8306.n0 a_23370_8306.t12 8.207
R2820 a_23370_8306.n23 a_23370_8306.t20 7.146
R2821 a_23370_8306.n4 a_23370_8306.t25 7.146
R2822 a_23370_8306.n4 a_23370_8306.t35 7.146
R2823 a_23370_8306.n3 a_23370_8306.t24 7.146
R2824 a_23370_8306.n3 a_23370_8306.t34 7.146
R2825 a_23370_8306.n2 a_23370_8306.t32 7.146
R2826 a_23370_8306.n2 a_23370_8306.t27 7.146
R2827 a_23370_8306.n16 a_23370_8306.t33 7.146
R2828 a_23370_8306.n16 a_23370_8306.t30 7.146
R2829 a_23370_8306.n15 a_23370_8306.t31 7.146
R2830 a_23370_8306.n15 a_23370_8306.t29 7.146
R2831 a_23370_8306.n14 a_23370_8306.t26 7.146
R2832 a_23370_8306.n14 a_23370_8306.t28 7.146
R2833 a_23370_8306.n13 a_23370_8306.t14 7.146
R2834 a_23370_8306.n12 a_23370_8306.t17 7.146
R2835 a_23370_8306.n11 a_23370_8306.t10 7.146
R2836 a_23370_8306.n11 a_23370_8306.t16 7.146
R2837 a_23370_8306.n10 a_23370_8306.t6 7.146
R2838 a_23370_8306.n10 a_23370_8306.t22 7.146
R2839 a_23370_8306.n9 a_23370_8306.t2 7.146
R2840 a_23370_8306.n9 a_23370_8306.t23 7.146
R2841 a_23370_8306.n8 a_23370_8306.t5 7.146
R2842 a_23370_8306.n8 a_23370_8306.t4 7.146
R2843 a_23370_8306.n7 a_23370_8306.t1 7.146
R2844 a_23370_8306.n7 a_23370_8306.t0 7.146
R2845 a_23370_8306.n6 a_23370_8306.t9 7.146
R2846 a_23370_8306.n6 a_23370_8306.t8 7.146
R2847 a_23370_8306.n1 a_23370_8306.t15 7.146
R2848 a_23370_8306.n0 a_23370_8306.t19 7.146
R2849 a_23370_8306.n22 a_23370_8306.t18 7.146
R2850 a_23370_8306.n22 a_23370_8306.t7 7.146
R2851 a_23370_8306.n21 a_23370_8306.t13 7.146
R2852 a_23370_8306.n21 a_23370_8306.t3 7.146
R2853 a_23370_8306.t11 a_23370_8306.n23 7.146
R2854 a_23370_8306.n5 a_23370_8306.n4 1.938
R2855 a_23370_8306.n17 a_23370_8306.n16 1.938
R2856 a_23370_8306.n17 a_23370_8306.n13 1.493
R2857 a_23370_8306.n5 a_23370_8306.n1 1.493
R2858 a_23370_8306.n18 a_23370_8306.n11 1.386
R2859 a_23370_8306.n19 a_23370_8306.n8 1.386
R2860 a_23370_8306.n23 a_23370_8306.n20 1.386
R2861 a_23370_8306.n13 a_23370_8306.n12 1.061
R2862 a_23370_8306.n1 a_23370_8306.n0 1.061
R2863 a_23370_8306.n3 a_23370_8306.n2 0.865
R2864 a_23370_8306.n4 a_23370_8306.n3 0.865
R2865 a_23370_8306.n15 a_23370_8306.n14 0.865
R2866 a_23370_8306.n16 a_23370_8306.n15 0.865
R2867 a_23370_8306.n20 a_23370_8306.n5 0.831
R2868 a_23370_8306.n20 a_23370_8306.n19 0.831
R2869 a_23370_8306.n19 a_23370_8306.n18 0.831
R2870 a_23370_8306.n18 a_23370_8306.n17 0.831
R2871 a_23370_8306.n10 a_23370_8306.n9 0.827
R2872 a_23370_8306.n11 a_23370_8306.n10 0.827
R2873 a_23370_8306.n7 a_23370_8306.n6 0.827
R2874 a_23370_8306.n8 a_23370_8306.n7 0.827
R2875 a_23370_8306.n22 a_23370_8306.n21 0.827
R2876 a_23370_8306.n23 a_23370_8306.n22 0.827
R2877 vbias1.n446 vbias1.n441 160.035
R2878 vbias1.n296 vbias1.n295 160.035
R2879 vbias1.n452 vbias1.n448 160.035
R2880 vbias1.n446 vbias1.n445 160.035
R2881 vbias1.n304 vbias1.n303 160.035
R2882 vbias1.n296 vbias1.n294 160.035
R2883 vbias1.n77 vbias1.n76 62.435
R2884 vbias1.n72 vbias1.n53 62.435
R2885 vbias1.n337 vbias1.n336 62.435
R2886 vbias1.n329 vbias1.n326 62.435
R2887 vbias1.n401 vbias1.n400 62.435
R2888 vbias1.n393 vbias1.n378 62.435
R2889 vbias1.n348 vbias1.n342 62.435
R2890 vbias1.n340 vbias1.n324 62.435
R2891 vbias1.n69 vbias1.n54 62.435
R2892 vbias1.n61 vbias1.n55 62.435
R2893 vbias1.t128 vbias1.n74 55.951
R2894 vbias1.t127 vbias1.n362 55.945
R2895 vbias1.t59 vbias1.n458 55.942
R2896 vbias1.t117 vbias1.n470 55.942
R2897 vbias1.t154 vbias1.n482 55.942
R2898 vbias1.t143 vbias1.n494 55.942
R2899 vbias1.t65 vbias1.n506 55.942
R2900 vbias1.t107 vbias1.n518 55.942
R2901 vbias1.t55 vbias1.n530 55.942
R2902 vbias1.t97 vbias1.n542 55.942
R2903 vbias1.t82 vbias1.n554 55.942
R2904 vbias1.t90 vbias1.n566 55.942
R2905 vbias1.t139 vbias1.n578 55.942
R2906 vbias1.t83 vbias1.n590 55.942
R2907 vbias1.t134 vbias1.n602 55.942
R2908 vbias1.t122 vbias1.n614 55.942
R2909 vbias1.t27 vbias1.n626 55.942
R2910 vbias1.t66 vbias1.n638 55.942
R2911 vbias1.t151 vbias1.n650 55.942
R2912 vbias1.t31 vbias1.n327 55.94
R2913 vbias1.t22 vbias1.n300 55.94
R2914 vbias1.t25 vbias1.n84 55.94
R2915 vbias1.t123 vbias1.n94 55.94
R2916 vbias1.t88 vbias1.n106 55.94
R2917 vbias1.t120 vbias1.n116 55.94
R2918 vbias1.t70 vbias1.n128 55.94
R2919 vbias1.t150 vbias1.n138 55.94
R2920 vbias1.t114 vbias1.n150 55.94
R2921 vbias1.t80 vbias1.n160 55.94
R2922 vbias1.t63 vbias1.n172 55.94
R2923 vbias1.t24 vbias1.n182 55.94
R2924 vbias1.t96 vbias1.n194 55.94
R2925 vbias1.t105 vbias1.n204 55.94
R2926 vbias1.t73 vbias1.n216 55.94
R2927 vbias1.t36 vbias1.n226 55.94
R2928 vbias1.t87 vbias1.n238 55.94
R2929 vbias1.t35 vbias1.n248 55.94
R2930 vbias1.t133 vbias1.n260 55.94
R2931 vbias1.t104 vbias1.n270 55.94
R2932 vbias1.t0 vbias1.n20 55.935
R2933 vbias1.t14 vbias1.n423 55.935
R2934 vbias1.t18 vbias1.n3 55.934
R2935 vbias1.t64 vbias1.n283 55.92
R2936 vbias1.t8 vbias1.n381 55.92
R2937 vbias1.t58 vbias1.n663 55.92
R2938 vbias1.t43 vbias1.n686 55.915
R2939 vbias1.n679 vbias1.t144 55.915
R2940 vbias1.n664 vbias1.t58 55.915
R2941 vbias1.n651 vbias1.t146 55.915
R2942 vbias1.n639 vbias1.t66 55.915
R2943 vbias1.n627 vbias1.t153 55.915
R2944 vbias1.n615 vbias1.t122 55.915
R2945 vbias1.n603 vbias1.t131 55.915
R2946 vbias1.n591 vbias1.t83 55.915
R2947 vbias1.n579 vbias1.t136 55.915
R2948 vbias1.n567 vbias1.t90 55.915
R2949 vbias1.n555 vbias1.t76 55.915
R2950 vbias1.n543 vbias1.t97 55.915
R2951 vbias1.n531 vbias1.t48 55.915
R2952 vbias1.n519 vbias1.t107 55.915
R2953 vbias1.n507 vbias1.t57 55.915
R2954 vbias1.n495 vbias1.t143 55.915
R2955 vbias1.n483 vbias1.t149 55.915
R2956 vbias1.n471 vbias1.t117 55.915
R2957 vbias1.n459 vbias1.t52 55.915
R2958 vbias1.n687 vbias1.t43 55.915
R2959 vbias1.n291 vbias1.t39 55.915
R2960 vbias1.n280 vbias1.t98 55.915
R2961 vbias1.n268 vbias1.t47 55.915
R2962 vbias1.n258 vbias1.t108 55.915
R2963 vbias1.n246 vbias1.t28 55.915
R2964 vbias1.n236 vbias1.t109 55.915
R2965 vbias1.n224 vbias1.t148 55.915
R2966 vbias1.n214 vbias1.t118 55.915
R2967 vbias1.n202 vbias1.t54 55.915
R2968 vbias1.n192 vbias1.t124 55.915
R2969 vbias1.n180 vbias1.t30 55.915
R2970 vbias1.n170 vbias1.t129 55.915
R2971 vbias1.n158 vbias1.t72 55.915
R2972 vbias1.n148 vbias1.t135 55.915
R2973 vbias1.n136 vbias1.t41 55.915
R2974 vbias1.n126 vbias1.t102 55.915
R2975 vbias1.n114 vbias1.t85 55.915
R2976 vbias1.n104 vbias1.t46 55.915
R2977 vbias1.n92 vbias1.t92 55.915
R2978 vbias1.n83 vbias1.t26 55.915
R2979 vbias1.n674 vbias1.t95 55.915
R2980 vbias1.n661 vbias1.t130 55.915
R2981 vbias1.t146 vbias1.n649 55.915
R2982 vbias1.n637 vbias1.t51 55.915
R2983 vbias1.n625 vbias1.t74 55.915
R2984 vbias1.t116 vbias1.n613 55.915
R2985 vbias1.n601 vbias1.t37 55.915
R2986 vbias1.n589 vbias1.t68 55.915
R2987 vbias1.t136 vbias1.n577 55.915
R2988 vbias1.n565 vbias1.t138 55.915
R2989 vbias1.n553 vbias1.t115 55.915
R2990 vbias1.t91 vbias1.n541 55.915
R2991 vbias1.n529 vbias1.t71 55.915
R2992 vbias1.n517 vbias1.t121 55.915
R2993 vbias1.t57 vbias1.n505 55.915
R2994 vbias1.n493 vbias1.t81 55.915
R2995 vbias1.n481 vbias1.t29 55.915
R2996 vbias1.t111 vbias1.n469 55.915
R2997 vbias1.n457 vbias1.t38 55.915
R2998 vbias1.t39 vbias1.n286 55.915
R2999 vbias1.t93 vbias1.n275 55.915
R3000 vbias1.t47 vbias1.n263 55.915
R3001 vbias1.t101 vbias1.n253 55.915
R3002 vbias1.t28 vbias1.n241 55.915
R3003 vbias1.t103 vbias1.n231 55.915
R3004 vbias1.t148 vbias1.n219 55.915
R3005 vbias1.t112 vbias1.n209 55.915
R3006 vbias1.t54 vbias1.n197 55.915
R3007 vbias1.t119 vbias1.n187 55.915
R3008 vbias1.t30 vbias1.n175 55.915
R3009 vbias1.t125 vbias1.n165 55.915
R3010 vbias1.t72 vbias1.n153 55.915
R3011 vbias1.t132 vbias1.n143 55.915
R3012 vbias1.t41 vbias1.n131 55.915
R3013 vbias1.t94 vbias1.n121 55.915
R3014 vbias1.t85 vbias1.n109 55.915
R3015 vbias1.t40 vbias1.n99 55.915
R3016 vbias1.t92 vbias1.n87 55.915
R3017 vbias1.t152 vbias1.n82 55.915
R3018 vbias1.n82 vbias1.t75 55.915
R3019 vbias1.n83 vbias1.t152 55.915
R3020 vbias1.n87 vbias1.t25 55.915
R3021 vbias1.n92 vbias1.t99 55.915
R3022 vbias1.n99 vbias1.t123 55.915
R3023 vbias1.n104 vbias1.t40 55.915
R3024 vbias1.n109 vbias1.t88 55.915
R3025 vbias1.n114 vbias1.t89 55.915
R3026 vbias1.n121 vbias1.t120 55.915
R3027 vbias1.n126 vbias1.t94 55.915
R3028 vbias1.n131 vbias1.t70 55.915
R3029 vbias1.n136 vbias1.t49 55.915
R3030 vbias1.n143 vbias1.t150 55.915
R3031 vbias1.n148 vbias1.t132 55.915
R3032 vbias1.n153 vbias1.t114 55.915
R3033 vbias1.n158 vbias1.t77 55.915
R3034 vbias1.n165 vbias1.t80 55.915
R3035 vbias1.n170 vbias1.t125 55.915
R3036 vbias1.n175 vbias1.t63 55.915
R3037 vbias1.n180 vbias1.t33 55.915
R3038 vbias1.n187 vbias1.t24 55.915
R3039 vbias1.n192 vbias1.t119 55.915
R3040 vbias1.n197 vbias1.t96 55.915
R3041 vbias1.n202 vbias1.t60 55.915
R3042 vbias1.n209 vbias1.t105 55.915
R3043 vbias1.n214 vbias1.t112 55.915
R3044 vbias1.n219 vbias1.t73 55.915
R3045 vbias1.n224 vbias1.t155 55.915
R3046 vbias1.n231 vbias1.t36 55.915
R3047 vbias1.n236 vbias1.t103 55.915
R3048 vbias1.n241 vbias1.t87 55.915
R3049 vbias1.n246 vbias1.t32 55.915
R3050 vbias1.n253 vbias1.t35 55.915
R3051 vbias1.n258 vbias1.t101 55.915
R3052 vbias1.n263 vbias1.t133 55.915
R3053 vbias1.n268 vbias1.t56 55.915
R3054 vbias1.n275 vbias1.t104 55.915
R3055 vbias1.n280 vbias1.t93 55.915
R3056 vbias1.n286 vbias1.t64 55.915
R3057 vbias1.n291 vbias1.t45 55.915
R3058 vbias1.t144 vbias1.n674 55.915
R3059 vbias1.t53 vbias1.n661 55.915
R3060 vbias1.n664 vbias1.t53 55.915
R3061 vbias1.n649 vbias1.t147 55.915
R3062 vbias1.n651 vbias1.t151 55.915
R3063 vbias1.t62 vbias1.n637 55.915
R3064 vbias1.n639 vbias1.t62 55.915
R3065 vbias1.t153 vbias1.n625 55.915
R3066 vbias1.n627 vbias1.t27 55.915
R3067 vbias1.n613 vbias1.t106 55.915
R3068 vbias1.n615 vbias1.t116 55.915
R3069 vbias1.t131 vbias1.n601 55.915
R3070 vbias1.n603 vbias1.t134 55.915
R3071 vbias1.t79 vbias1.n589 55.915
R3072 vbias1.n591 vbias1.t79 55.915
R3073 vbias1.n577 vbias1.t110 55.915
R3074 vbias1.n579 vbias1.t139 55.915
R3075 vbias1.t86 vbias1.n565 55.915
R3076 vbias1.n567 vbias1.t86 55.915
R3077 vbias1.t76 vbias1.n553 55.915
R3078 vbias1.n555 vbias1.t82 55.915
R3079 vbias1.n541 vbias1.t42 55.915
R3080 vbias1.n543 vbias1.t91 55.915
R3081 vbias1.t48 vbias1.n529 55.915
R3082 vbias1.n531 vbias1.t55 55.915
R3083 vbias1.t100 vbias1.n517 55.915
R3084 vbias1.n519 vbias1.t100 55.915
R3085 vbias1.n505 vbias1.t142 55.915
R3086 vbias1.n507 vbias1.t65 55.915
R3087 vbias1.t141 vbias1.n493 55.915
R3088 vbias1.n495 vbias1.t141 55.915
R3089 vbias1.t149 vbias1.n481 55.915
R3090 vbias1.n483 vbias1.t154 55.915
R3091 vbias1.n469 vbias1.t44 55.915
R3092 vbias1.n471 vbias1.t111 55.915
R3093 vbias1.t52 vbias1.n457 55.915
R3094 vbias1.n459 vbias1.t59 55.915
R3095 vbias1.n687 vbias1.t50 55.915
R3096 vbias1.n679 vbias1.t145 55.915
R3097 vbias1.n686 vbias1.t69 55.914
R3098 vbias1.t99 vbias1.n91 55.914
R3099 vbias1.t46 vbias1.n103 55.914
R3100 vbias1.t89 vbias1.n113 55.914
R3101 vbias1.t102 vbias1.n125 55.914
R3102 vbias1.t49 vbias1.n135 55.914
R3103 vbias1.t135 vbias1.n147 55.914
R3104 vbias1.t77 vbias1.n157 55.914
R3105 vbias1.t129 vbias1.n169 55.914
R3106 vbias1.t33 vbias1.n179 55.914
R3107 vbias1.t124 vbias1.n191 55.914
R3108 vbias1.t60 vbias1.n201 55.914
R3109 vbias1.t118 vbias1.n213 55.914
R3110 vbias1.t155 vbias1.n223 55.914
R3111 vbias1.t109 vbias1.n235 55.914
R3112 vbias1.t32 vbias1.n245 55.914
R3113 vbias1.t108 vbias1.n257 55.914
R3114 vbias1.t56 vbias1.n267 55.914
R3115 vbias1.t98 vbias1.n279 55.914
R3116 vbias1.t45 vbias1.n290 55.914
R3117 vbias1.t140 vbias1.n346 55.914
R3118 vbias1.t20 vbias1.n411 55.914
R3119 vbias1.t34 vbias1.n59 55.914
R3120 vbias1.t95 vbias1.n669 55.914
R3121 vbias1.t130 vbias1.n656 55.914
R3122 vbias1.t147 vbias1.n644 55.914
R3123 vbias1.t51 vbias1.n632 55.914
R3124 vbias1.t74 vbias1.n620 55.914
R3125 vbias1.t106 vbias1.n608 55.914
R3126 vbias1.t37 vbias1.n596 55.914
R3127 vbias1.t68 vbias1.n584 55.914
R3128 vbias1.t110 vbias1.n572 55.914
R3129 vbias1.t138 vbias1.n560 55.914
R3130 vbias1.t115 vbias1.n548 55.914
R3131 vbias1.t42 vbias1.n536 55.914
R3132 vbias1.t71 vbias1.n524 55.914
R3133 vbias1.t121 vbias1.n512 55.914
R3134 vbias1.t142 vbias1.n500 55.914
R3135 vbias1.t81 vbias1.n488 55.914
R3136 vbias1.t29 vbias1.n476 55.914
R3137 vbias1.t44 vbias1.n464 55.914
R3138 vbias1.t38 vbias1.n447 55.914
R3139 vbias1.t145 vbias1.n678 55.914
R3140 vbias1.t84 vbias1.n358 55.914
R3141 vbias1.t10 vbias1.n318 55.914
R3142 vbias1.t4 vbias1.n398 55.914
R3143 vbias1.t67 vbias1.n31 55.914
R3144 vbias1.t113 vbias1.n38 55.914
R3145 vbias1.n328 vbias1.t31 55.912
R3146 vbias1.n347 vbias1.t140 55.912
R3147 vbias1.n339 vbias1.t137 55.912
R3148 vbias1.t137 vbias1.n338 55.912
R3149 vbias1.n363 vbias1.t127 55.912
R3150 vbias1.n412 vbias1.t20 55.912
R3151 vbias1.t16 vbias1.n418 55.912
R3152 vbias1.n419 vbias1.t16 55.912
R3153 vbias1.n424 vbias1.t14 55.912
R3154 vbias1.n60 vbias1.t34 55.912
R3155 vbias1.t126 vbias1.n70 55.912
R3156 vbias1.n71 vbias1.t126 55.912
R3157 vbias1.n75 vbias1.t128 55.912
R3158 vbias1.n4 vbias1.t18 55.912
R3159 vbias1.t2 vbias1.n14 55.912
R3160 vbias1.n15 vbias1.t2 55.912
R3161 vbias1.n21 vbias1.t0 55.912
R3162 vbias1.n359 vbias1.t84 55.912
R3163 vbias1.n372 vbias1.t78 55.912
R3164 vbias1.t78 vbias1.n371 55.912
R3165 vbias1.n382 vbias1.t8 55.912
R3166 vbias1.t6 vbias1.n391 55.912
R3167 vbias1.n392 vbias1.t6 55.912
R3168 vbias1.n301 vbias1.t22 55.912
R3169 vbias1.t12 vbias1.n310 55.912
R3170 vbias1.n311 vbias1.t12 55.912
R3171 vbias1.n319 vbias1.t10 55.912
R3172 vbias1.n399 vbias1.t4 55.912
R3173 vbias1.n32 vbias1.t67 55.912
R3174 vbias1.n48 vbias1.t61 55.912
R3175 vbias1.t61 vbias1.n47 55.912
R3176 vbias1.n39 vbias1.t113 55.912
R3177 vbias1.n299 vbias1.n298 52.349
R3178 vbias1.n440 vbias1.n26 47.684
R3179 vbias1.n438 vbias1.n81 47.684
R3180 vbias1.n406 vbias1.n405 47.684
R3181 vbias1.n353 vbias1.n352 47.684
R3182 vbias1.n9 vbias1.n8 47.509
R3183 vbias1.n65 vbias1.n64 47.509
R3184 vbias1.n387 vbias1.n386 47.509
R3185 vbias1.n334 vbias1.n333 47.509
R3186 vbias1.n432 vbias1.n429 45.929
R3187 vbias1.n432 vbias1.n428 45.929
R3188 vbias1.n437 vbias1.n436 44.747
R3189 vbias1.n432 vbias1.n431 37.195
R3190 vbias1.n433 vbias1.n432 37.195
R3191 vbias1.n436 vbias1.n433 37.195
R3192 vbias1.n436 vbias1.n435 37.195
R3193 vbias1.n455 vbias1.n452 36.608
R3194 vbias1.n431 vbias1.n430 32.954
R3195 vbias1.n435 vbias1.n434 32.954
R3196 vbias1.n322 vbias1.n296 29.722
R3197 vbias1.n305 vbias1.n304 29.547
R3198 vbias1.n461 vbias1.n446 23.454
R3199 vbias1.n317 vbias1.n314 16.084
R3200 vbias1.n8 vbias1.n6 9.329
R3201 vbias1.n333 vbias1.n331 9.329
R3202 vbias1.n64 vbias1.n62 9.329
R3203 vbias1.n26 vbias1.n24 9.329
R3204 vbias1.n444 vbias1.n443 9.329
R3205 vbias1.n444 vbias1.n442 9.329
R3206 vbias1.n26 vbias1.n25 9.329
R3207 vbias1.n81 vbias1.n80 9.329
R3208 vbias1.n81 vbias1.n79 9.329
R3209 vbias1.n405 vbias1.n403 9.329
R3210 vbias1.n386 vbias1.n384 9.329
R3211 vbias1.n386 vbias1.n385 9.329
R3212 vbias1.n333 vbias1.n332 9.329
R3213 vbias1.n405 vbias1.n404 9.329
R3214 vbias1.n352 vbias1.n351 9.329
R3215 vbias1.n352 vbias1.n350 9.329
R3216 vbias1.n451 vbias1.n450 9.329
R3217 vbias1.n451 vbias1.n449 9.329
R3218 vbias1.n8 vbias1.n7 9.329
R3219 vbias1.n64 vbias1.n63 9.329
R3220 vbias1.n294 vbias1.t13 7.141
R3221 vbias1.n303 vbias1.t23 7.141
R3222 vbias1.n433 vbias1.t17 7.141
R3223 vbias1.n431 vbias1.t21 7.141
R3224 vbias1.n431 vbias1.t9 7.141
R3225 vbias1.n433 vbias1.t7 7.141
R3226 vbias1.n435 vbias1.t5 7.141
R3227 vbias1.n435 vbias1.t15 7.141
R3228 vbias1.n445 vbias1.t3 7.141
R3229 vbias1.n448 vbias1.t19 7.141
R3230 vbias1.n295 vbias1.t11 7.141
R3231 vbias1.n441 vbias1.t1 7.141
R3232 vbias1.n446 vbias1.n444 3.275
R3233 vbias1.n452 vbias1.n451 3.275
R3234 vbias1.n93 vbias1.n83 0.399
R3235 vbias1.n463 vbias1.n440 0.394
R3236 vbias1.n322 vbias1.n293 0.386
R3237 vbias1.n353 vbias1.n322 0.386
R3238 vbias1.n376 vbias1.n353 0.386
R3239 vbias1.n406 vbias1.n376 0.386
R3240 vbias1.n437 vbias1.n406 0.386
R3241 vbias1.n438 vbias1.n437 0.386
R3242 vbias1.n439 vbias1.n438 0.386
R3243 vbias1.n440 vbias1.n439 0.386
R3244 vbias1.n475 vbias1.n463 0.386
R3245 vbias1.n487 vbias1.n475 0.386
R3246 vbias1.n499 vbias1.n487 0.386
R3247 vbias1.n511 vbias1.n499 0.386
R3248 vbias1.n523 vbias1.n511 0.386
R3249 vbias1.n535 vbias1.n523 0.386
R3250 vbias1.n547 vbias1.n535 0.386
R3251 vbias1.n559 vbias1.n547 0.386
R3252 vbias1.n571 vbias1.n559 0.386
R3253 vbias1.n583 vbias1.n571 0.386
R3254 vbias1.n595 vbias1.n583 0.386
R3255 vbias1.n607 vbias1.n595 0.386
R3256 vbias1.n619 vbias1.n607 0.386
R3257 vbias1.n631 vbias1.n619 0.386
R3258 vbias1.n643 vbias1.n631 0.386
R3259 vbias1.n655 vbias1.n643 0.386
R3260 vbias1.n668 vbias1.n655 0.386
R3261 vbias1.n683 vbias1.n668 0.386
R3262 vbias1.n690 vbias1.n683 0.386
R3263 vbias1.n105 vbias1.n93 0.384
R3264 vbias1.n115 vbias1.n105 0.384
R3265 vbias1.n127 vbias1.n115 0.384
R3266 vbias1.n137 vbias1.n127 0.384
R3267 vbias1.n149 vbias1.n137 0.384
R3268 vbias1.n159 vbias1.n149 0.384
R3269 vbias1.n171 vbias1.n159 0.384
R3270 vbias1.n181 vbias1.n171 0.384
R3271 vbias1.n193 vbias1.n181 0.384
R3272 vbias1.n203 vbias1.n193 0.384
R3273 vbias1.n215 vbias1.n203 0.384
R3274 vbias1.n225 vbias1.n215 0.384
R3275 vbias1.n237 vbias1.n225 0.384
R3276 vbias1.n247 vbias1.n237 0.384
R3277 vbias1.n259 vbias1.n247 0.384
R3278 vbias1.n269 vbias1.n259 0.384
R3279 vbias1.n281 vbias1.n269 0.384
R3280 vbias1.n293 vbias1.n281 0.384
R3281 vbias1.n684 vbias1 0.367
R3282 vbias1.n68 vbias1.n67 0.181
R3283 vbias1.n12 vbias1.n11 0.181
R3284 vbias1.n42 vbias1.n41 0.181
R3285 vbias1.n308 vbias1.n307 0.181
R3286 vbias1.n330 vbias1.n325 0.181
R3287 vbias1.n369 vbias1.n368 0.181
R3288 vbias1.n414 vbias1.n407 0.181
R3289 vbias1.n389 vbias1.n379 0.181
R3290 vbias1.n73 vbias1.n52 0.135
R3291 vbias1.n34 vbias1.n27 0.135
R3292 vbias1.n17 vbias1.n0 0.135
R3293 vbias1.n426 vbias1.n421 0.135
R3294 vbias1.n394 vbias1.n377 0.135
R3295 vbias1.n361 vbias1.n354 0.135
R3296 vbias1.n341 vbias1.n323 0.135
R3297 vbias1.n313 vbias1.n297 0.135
R3298 vbias1.n19 vbias1.n18 0.109
R3299 vbias1.n2 vbias1.n1 0.091
R3300 vbias1.n31 vbias1.n30 0.036
R3301 vbias1.n91 vbias1.n90 0.036
R3302 vbias1.n678 vbias1.n677 0.027
R3303 vbias1.n318 vbias1.n317 0.021
R3304 vbias1.n346 vbias1.n345 0.021
R3305 vbias1.n358 vbias1.n357 0.021
R3306 vbias1.n398 vbias1.n397 0.021
R3307 vbias1.n103 vbias1.n102 0.021
R3308 vbias1.n113 vbias1.n112 0.021
R3309 vbias1.n125 vbias1.n124 0.021
R3310 vbias1.n135 vbias1.n134 0.021
R3311 vbias1.n147 vbias1.n146 0.021
R3312 vbias1.n157 vbias1.n156 0.021
R3313 vbias1.n169 vbias1.n168 0.021
R3314 vbias1.n179 vbias1.n178 0.021
R3315 vbias1.n191 vbias1.n190 0.021
R3316 vbias1.n201 vbias1.n200 0.021
R3317 vbias1.n213 vbias1.n212 0.021
R3318 vbias1.n223 vbias1.n222 0.021
R3319 vbias1.n235 vbias1.n234 0.021
R3320 vbias1.n245 vbias1.n244 0.021
R3321 vbias1.n257 vbias1.n256 0.021
R3322 vbias1.n267 vbias1.n266 0.021
R3323 vbias1.n279 vbias1.n278 0.021
R3324 vbias1.n290 vbias1.n289 0.021
R3325 vbias1.n663 vbias1.n662 0.021
R3326 vbias1.n306 vbias1.n302 0.021
R3327 vbias1.n417 vbias1.n416 0.021
R3328 vbias1.n367 vbias1.n364 0.021
R3329 vbias1.n388 vbias1.n383 0.021
R3330 vbias1.n337 vbias1.n335 0.021
R3331 vbias1.n10 vbias1.n5 0.021
R3332 vbias1.n46 vbias1.n45 0.021
R3333 vbias1.n66 vbias1.n61 0.021
R3334 vbias1.n17 vbias1.n16 0.021
R3335 vbias1.n73 vbias1.n72 0.021
R3336 vbias1.n426 vbias1.n425 0.021
R3337 vbias1.n390 vbias1.n389 0.021
R3338 vbias1.n370 vbias1.n369 0.021
R3339 vbias1.n330 vbias1.n329 0.021
R3340 vbias1.n309 vbias1.n308 0.021
R3341 vbias1.n394 vbias1.n393 0.021
R3342 vbias1.n361 vbias1.n360 0.021
R3343 vbias1.n341 vbias1.n340 0.021
R3344 vbias1.n313 vbias1.n312 0.021
R3345 vbias1.n34 vbias1.n33 0.021
R3346 vbias1.n42 vbias1.n40 0.021
R3347 vbias1.n13 vbias1.n12 0.021
R3348 vbias1.n69 vbias1.n68 0.021
R3349 vbias1.n414 vbias1.n413 0.021
R3350 vbias1.n50 vbias1.n49 0.021
R3351 vbias1.n23 vbias1.n22 0.021
R3352 vbias1.n78 vbias1.n77 0.021
R3353 vbias1.n427 vbias1.n420 0.021
R3354 vbias1.n374 vbias1.n373 0.021
R3355 vbias1.n402 vbias1.n401 0.021
R3356 vbias1.n349 vbias1.n348 0.021
R3357 vbias1.n321 vbias1.n320 0.021
R3358 vbias1.n38 vbias1.n37 0.02
R3359 vbias1.n283 vbias1.n282 0.019
R3360 vbias1.n58 vbias1.n57 0.018
R3361 vbias1.n381 vbias1.n380 0.016
R3362 vbias1.n410 vbias1.n409 0.016
R3363 vbias1.n44 vbias1.n43 0.016
R3364 vbias1.n366 vbias1.n365 0.016
R3365 vbias1.n423 vbias1.n422 0.015
R3366 vbias1.n20 vbias1.n19 0.015
R3367 vbias1.n274 vbias1.n273 0.015
R3368 vbias1.n252 vbias1.n251 0.015
R3369 vbias1.n230 vbias1.n229 0.015
R3370 vbias1.n208 vbias1.n207 0.015
R3371 vbias1.n186 vbias1.n185 0.015
R3372 vbias1.n164 vbias1.n163 0.015
R3373 vbias1.n142 vbias1.n141 0.015
R3374 vbias1.n120 vbias1.n119 0.015
R3375 vbias1.n98 vbias1.n97 0.015
R3376 vbias1.n278 vbias1.n277 0.015
R3377 vbias1.n256 vbias1.n255 0.015
R3378 vbias1.n234 vbias1.n233 0.015
R3379 vbias1.n212 vbias1.n211 0.015
R3380 vbias1.n190 vbias1.n189 0.015
R3381 vbias1.n168 vbias1.n167 0.015
R3382 vbias1.n146 vbias1.n145 0.015
R3383 vbias1.n124 vbias1.n123 0.015
R3384 vbias1.n102 vbias1.n101 0.015
R3385 vbias1.n112 vbias1.n111 0.015
R3386 vbias1.n134 vbias1.n133 0.015
R3387 vbias1.n156 vbias1.n155 0.015
R3388 vbias1.n178 vbias1.n177 0.015
R3389 vbias1.n200 vbias1.n199 0.015
R3390 vbias1.n222 vbias1.n221 0.015
R3391 vbias1.n244 vbias1.n243 0.015
R3392 vbias1.n266 vbias1.n265 0.015
R3393 vbias1.n289 vbias1.n288 0.015
R3394 vbias1.n357 vbias1.n356 0.015
R3395 vbias1.n345 vbias1.n344 0.015
R3396 vbias1.n317 vbias1.n316 0.015
R3397 vbias1.n397 vbias1.n396 0.015
R3398 vbias1 vbias1.n691 0.014
R3399 vbias1.n281 vbias1.n280 0.014
R3400 vbias1.n269 vbias1.n268 0.014
R3401 vbias1.n259 vbias1.n258 0.014
R3402 vbias1.n247 vbias1.n246 0.014
R3403 vbias1.n237 vbias1.n236 0.014
R3404 vbias1.n225 vbias1.n224 0.014
R3405 vbias1.n215 vbias1.n214 0.014
R3406 vbias1.n203 vbias1.n202 0.014
R3407 vbias1.n193 vbias1.n192 0.014
R3408 vbias1.n181 vbias1.n180 0.014
R3409 vbias1.n171 vbias1.n170 0.014
R3410 vbias1.n159 vbias1.n158 0.014
R3411 vbias1.n149 vbias1.n148 0.014
R3412 vbias1.n137 vbias1.n136 0.014
R3413 vbias1.n127 vbias1.n126 0.014
R3414 vbias1.n115 vbias1.n114 0.014
R3415 vbias1.n105 vbias1.n104 0.014
R3416 vbias1.n93 vbias1.n92 0.014
R3417 vbias1.n439 vbias1.n51 0.012
R3418 vbias1.n376 vbias1.n375 0.012
R3419 vbias1.n86 vbias1.n85 0.012
R3420 vbias1.n108 vbias1.n107 0.012
R3421 vbias1.n130 vbias1.n129 0.012
R3422 vbias1.n152 vbias1.n151 0.012
R3423 vbias1.n174 vbias1.n173 0.012
R3424 vbias1.n196 vbias1.n195 0.012
R3425 vbias1.n218 vbias1.n217 0.012
R3426 vbias1.n240 vbias1.n239 0.012
R3427 vbias1.n262 vbias1.n261 0.012
R3428 vbias1.n285 vbias1.n284 0.012
R3429 vbias1.n681 vbias1.n680 0.011
R3430 vbias1.n666 vbias1.n665 0.011
R3431 vbias1.n653 vbias1.n652 0.011
R3432 vbias1.n641 vbias1.n640 0.011
R3433 vbias1.n629 vbias1.n628 0.011
R3434 vbias1.n617 vbias1.n616 0.011
R3435 vbias1.n605 vbias1.n604 0.011
R3436 vbias1.n593 vbias1.n592 0.011
R3437 vbias1.n581 vbias1.n580 0.011
R3438 vbias1.n569 vbias1.n568 0.011
R3439 vbias1.n557 vbias1.n556 0.011
R3440 vbias1.n545 vbias1.n544 0.011
R3441 vbias1.n533 vbias1.n532 0.011
R3442 vbias1.n521 vbias1.n520 0.011
R3443 vbias1.n509 vbias1.n508 0.011
R3444 vbias1.n497 vbias1.n496 0.011
R3445 vbias1.n485 vbias1.n484 0.011
R3446 vbias1.n473 vbias1.n472 0.011
R3447 vbias1.n461 vbias1.n460 0.011
R3448 vbias1.n689 vbias1.n688 0.011
R3449 vbias1.n293 vbias1.n292 0.01
R3450 vbias1.n672 vbias1.n671 0.01
R3451 vbias1.n635 vbias1.n634 0.01
R3452 vbias1.n599 vbias1.n598 0.01
R3453 vbias1.n563 vbias1.n562 0.01
R3454 vbias1.n527 vbias1.n526 0.01
R3455 vbias1.n491 vbias1.n490 0.01
R3456 vbias1.n455 vbias1.n454 0.01
R3457 vbias1.n467 vbias1.n466 0.01
R3458 vbias1.n503 vbias1.n502 0.01
R3459 vbias1.n539 vbias1.n538 0.01
R3460 vbias1.n575 vbias1.n574 0.01
R3461 vbias1.n611 vbias1.n610 0.01
R3462 vbias1.n647 vbias1.n646 0.01
R3463 vbias1.n479 vbias1.n478 0.01
R3464 vbias1.n515 vbias1.n514 0.01
R3465 vbias1.n551 vbias1.n550 0.01
R3466 vbias1.n587 vbias1.n586 0.01
R3467 vbias1.n623 vbias1.n622 0.01
R3468 vbias1.n659 vbias1.n658 0.01
R3469 vbias1.n685 vbias1.n684 0.009
R3470 vbias1.n683 vbias1.n681 0.008
R3471 vbias1.n668 vbias1.n666 0.008
R3472 vbias1.n655 vbias1.n653 0.008
R3473 vbias1.n643 vbias1.n641 0.008
R3474 vbias1.n631 vbias1.n629 0.008
R3475 vbias1.n619 vbias1.n617 0.008
R3476 vbias1.n607 vbias1.n605 0.008
R3477 vbias1.n595 vbias1.n593 0.008
R3478 vbias1.n583 vbias1.n581 0.008
R3479 vbias1.n571 vbias1.n569 0.008
R3480 vbias1.n559 vbias1.n557 0.008
R3481 vbias1.n547 vbias1.n545 0.008
R3482 vbias1.n535 vbias1.n533 0.008
R3483 vbias1.n523 vbias1.n521 0.008
R3484 vbias1.n511 vbias1.n509 0.008
R3485 vbias1.n499 vbias1.n497 0.008
R3486 vbias1.n487 vbias1.n485 0.008
R3487 vbias1.n475 vbias1.n473 0.008
R3488 vbias1.n463 vbias1.n461 0.008
R3489 vbias1.n690 vbias1.n689 0.008
R3490 vbias1.n411 vbias1.n410 0.007
R3491 vbias1.n59 vbias1.n58 0.007
R3492 vbias1.n87 vbias1.n86 0.004
R3493 vbias1.n109 vbias1.n108 0.004
R3494 vbias1.n131 vbias1.n130 0.004
R3495 vbias1.n153 vbias1.n152 0.004
R3496 vbias1.n175 vbias1.n174 0.004
R3497 vbias1.n197 vbias1.n196 0.004
R3498 vbias1.n219 vbias1.n218 0.004
R3499 vbias1.n241 vbias1.n240 0.004
R3500 vbias1.n263 vbias1.n262 0.004
R3501 vbias1.n286 vbias1.n285 0.004
R3502 vbias1.n37 vbias1.n36 0.004
R3503 vbias1.n292 vbias1.n291 0.004
R3504 vbias1.n686 vbias1.n685 0.004
R3505 vbias1.n45 vbias1.n44 0.003
R3506 vbias1.n306 vbias1.n305 0.003
R3507 vbias1.n335 vbias1.n334 0.003
R3508 vbias1.n416 vbias1.n415 0.003
R3509 vbias1.n367 vbias1.n366 0.003
R3510 vbias1.n388 vbias1.n387 0.003
R3511 vbias1.n10 vbias1.n9 0.003
R3512 vbias1.n66 vbias1.n65 0.003
R3513 vbias1.n3 vbias1.n2 0.003
R3514 vbias1.n456 vbias1.n455 0.003
R3515 vbias1.n468 vbias1.n467 0.003
R3516 vbias1.n492 vbias1.n491 0.003
R3517 vbias1.n504 vbias1.n503 0.003
R3518 vbias1.n528 vbias1.n527 0.003
R3519 vbias1.n540 vbias1.n539 0.003
R3520 vbias1.n564 vbias1.n563 0.003
R3521 vbias1.n576 vbias1.n575 0.003
R3522 vbias1.n600 vbias1.n599 0.003
R3523 vbias1.n612 vbias1.n611 0.003
R3524 vbias1.n636 vbias1.n635 0.003
R3525 vbias1.n648 vbias1.n647 0.003
R3526 vbias1.n673 vbias1.n672 0.003
R3527 vbias1.n480 vbias1.n479 0.003
R3528 vbias1.n516 vbias1.n515 0.003
R3529 vbias1.n552 vbias1.n551 0.003
R3530 vbias1.n588 vbias1.n587 0.003
R3531 vbias1.n624 vbias1.n623 0.003
R3532 vbias1.n660 vbias1.n659 0.003
R3533 vbias1.n418 vbias1.n417 0.002
R3534 vbias1.n22 vbias1.n21 0.002
R3535 vbias1.n16 vbias1.n15 0.002
R3536 vbias1.n77 vbias1.n75 0.002
R3537 vbias1.n72 vbias1.n71 0.002
R3538 vbias1.n425 vbias1.n424 0.002
R3539 vbias1.n420 vbias1.n419 0.002
R3540 vbias1.n373 vbias1.n372 0.002
R3541 vbias1.n364 vbias1.n363 0.002
R3542 vbias1.n391 vbias1.n390 0.002
R3543 vbias1.n383 vbias1.n382 0.002
R3544 vbias1.n371 vbias1.n370 0.002
R3545 vbias1.n338 vbias1.n337 0.002
R3546 vbias1.n329 vbias1.n328 0.002
R3547 vbias1.n310 vbias1.n309 0.002
R3548 vbias1.n302 vbias1.n301 0.002
R3549 vbias1.n401 vbias1.n399 0.002
R3550 vbias1.n393 vbias1.n392 0.002
R3551 vbias1.n360 vbias1.n359 0.002
R3552 vbias1.n348 vbias1.n347 0.002
R3553 vbias1.n340 vbias1.n339 0.002
R3554 vbias1.n320 vbias1.n319 0.002
R3555 vbias1.n312 vbias1.n311 0.002
R3556 vbias1.n49 vbias1.n48 0.002
R3557 vbias1.n33 vbias1.n32 0.002
R3558 vbias1.n40 vbias1.n39 0.002
R3559 vbias1.n14 vbias1.n13 0.002
R3560 vbias1.n5 vbias1.n4 0.002
R3561 vbias1.n47 vbias1.n46 0.002
R3562 vbias1.n70 vbias1.n69 0.002
R3563 vbias1.n61 vbias1.n60 0.002
R3564 vbias1.n413 vbias1.n412 0.002
R3565 vbias1.n438 vbias1.n78 0.001
R3566 vbias1.n439 vbias1.n50 0.001
R3567 vbias1.n440 vbias1.n23 0.001
R3568 vbias1.n437 vbias1.n427 0.001
R3569 vbias1.n406 vbias1.n402 0.001
R3570 vbias1.n376 vbias1.n374 0.001
R3571 vbias1.n353 vbias1.n349 0.001
R3572 vbias1.n322 vbias1.n321 0.001
R3573 vbias1.n680 vbias1.n679 0.001
R3574 vbias1.n665 vbias1.n664 0.001
R3575 vbias1.n652 vbias1.n651 0.001
R3576 vbias1.n640 vbias1.n639 0.001
R3577 vbias1.n628 vbias1.n627 0.001
R3578 vbias1.n616 vbias1.n615 0.001
R3579 vbias1.n604 vbias1.n603 0.001
R3580 vbias1.n592 vbias1.n591 0.001
R3581 vbias1.n580 vbias1.n579 0.001
R3582 vbias1.n568 vbias1.n567 0.001
R3583 vbias1.n556 vbias1.n555 0.001
R3584 vbias1.n544 vbias1.n543 0.001
R3585 vbias1.n532 vbias1.n531 0.001
R3586 vbias1.n520 vbias1.n519 0.001
R3587 vbias1.n508 vbias1.n507 0.001
R3588 vbias1.n496 vbias1.n495 0.001
R3589 vbias1.n484 vbias1.n483 0.001
R3590 vbias1.n472 vbias1.n471 0.001
R3591 vbias1.n460 vbias1.n459 0.001
R3592 vbias1.n688 vbias1.n687 0.001
R3593 vbias1.n674 vbias1.n673 0.001
R3594 vbias1.n637 vbias1.n636 0.001
R3595 vbias1.n601 vbias1.n600 0.001
R3596 vbias1.n565 vbias1.n564 0.001
R3597 vbias1.n529 vbias1.n528 0.001
R3598 vbias1.n493 vbias1.n492 0.001
R3599 vbias1.n457 vbias1.n456 0.001
R3600 vbias1.n469 vbias1.n468 0.001
R3601 vbias1.n481 vbias1.n480 0.001
R3602 vbias1.n505 vbias1.n504 0.001
R3603 vbias1.n517 vbias1.n516 0.001
R3604 vbias1.n541 vbias1.n540 0.001
R3605 vbias1.n553 vbias1.n552 0.001
R3606 vbias1.n577 vbias1.n576 0.001
R3607 vbias1.n589 vbias1.n588 0.001
R3608 vbias1.n613 vbias1.n612 0.001
R3609 vbias1.n625 vbias1.n624 0.001
R3610 vbias1.n649 vbias1.n648 0.001
R3611 vbias1.n661 vbias1.n660 0.001
R3612 vbias1.n99 vbias1.n98 0.001
R3613 vbias1.n121 vbias1.n120 0.001
R3614 vbias1.n143 vbias1.n142 0.001
R3615 vbias1.n165 vbias1.n164 0.001
R3616 vbias1.n187 vbias1.n186 0.001
R3617 vbias1.n209 vbias1.n208 0.001
R3618 vbias1.n231 vbias1.n230 0.001
R3619 vbias1.n253 vbias1.n252 0.001
R3620 vbias1.n275 vbias1.n274 0.001
R3621 vbias1.n668 vbias1.n667 0.001
R3622 vbias1.n643 vbias1.n642 0.001
R3623 vbias1.n619 vbias1.n618 0.001
R3624 vbias1.n595 vbias1.n594 0.001
R3625 vbias1.n571 vbias1.n570 0.001
R3626 vbias1.n547 vbias1.n546 0.001
R3627 vbias1.n523 vbias1.n522 0.001
R3628 vbias1.n499 vbias1.n498 0.001
R3629 vbias1.n475 vbias1.n474 0.001
R3630 vbias1.n683 vbias1.n682 0.001
R3631 vbias1.n655 vbias1.n654 0.001
R3632 vbias1.n631 vbias1.n630 0.001
R3633 vbias1.n607 vbias1.n606 0.001
R3634 vbias1.n583 vbias1.n582 0.001
R3635 vbias1.n559 vbias1.n558 0.001
R3636 vbias1.n535 vbias1.n534 0.001
R3637 vbias1.n511 vbias1.n510 0.001
R3638 vbias1.n487 vbias1.n486 0.001
R3639 vbias1.n463 vbias1.n462 0.001
R3640 vbias1.n90 vbias1.n89 0.001
R3641 vbias1.n30 vbias1.n29 0.001
R3642 vbias1.n677 vbias1.n676 0.001
R3643 vbias1.n273 vbias1.n272 0.001
R3644 vbias1.n251 vbias1.n250 0.001
R3645 vbias1.n229 vbias1.n228 0.001
R3646 vbias1.n207 vbias1.n206 0.001
R3647 vbias1.n185 vbias1.n184 0.001
R3648 vbias1.n163 vbias1.n162 0.001
R3649 vbias1.n141 vbias1.n140 0.001
R3650 vbias1.n119 vbias1.n118 0.001
R3651 vbias1.n97 vbias1.n96 0.001
R3652 vbias1.n300 vbias1.n299 0.001
R3653 vbias1.n68 vbias1.n66 0.001
R3654 vbias1.n12 vbias1.n10 0.001
R3655 vbias1.n369 vbias1.n367 0.001
R3656 vbias1.n416 vbias1.n414 0.001
R3657 vbias1.n389 vbias1.n388 0.001
R3658 vbias1.n335 vbias1.n330 0.001
R3659 vbias1.n308 vbias1.n306 0.001
R3660 vbias1.n45 vbias1.n42 0.001
R3661 vbias1.n23 vbias1.n17 0.001
R3662 vbias1.n78 vbias1.n73 0.001
R3663 vbias1.n427 vbias1.n426 0.001
R3664 vbias1.n374 vbias1.n361 0.001
R3665 vbias1.n402 vbias1.n394 0.001
R3666 vbias1.n349 vbias1.n341 0.001
R3667 vbias1.n321 vbias1.n313 0.001
R3668 vbias1.n50 vbias1.n34 0.001
R3669 vbias1.n691 vbias1.n690 0.001
R3670 vbias1.n272 vbias1.n271 0.001
R3671 vbias1.n250 vbias1.n249 0.001
R3672 vbias1.n228 vbias1.n227 0.001
R3673 vbias1.n206 vbias1.n205 0.001
R3674 vbias1.n184 vbias1.n183 0.001
R3675 vbias1.n162 vbias1.n161 0.001
R3676 vbias1.n140 vbias1.n139 0.001
R3677 vbias1.n118 vbias1.n117 0.001
R3678 vbias1.n96 vbias1.n95 0.001
R3679 vbias1.n466 vbias1.n465 0.001
R3680 vbias1.n502 vbias1.n501 0.001
R3681 vbias1.n538 vbias1.n537 0.001
R3682 vbias1.n574 vbias1.n573 0.001
R3683 vbias1.n610 vbias1.n609 0.001
R3684 vbias1.n646 vbias1.n645 0.001
R3685 vbias1.n57 vbias1.n56 0.001
R3686 vbias1.n29 vbias1.n28 0.001
R3687 vbias1.n277 vbias1.n276 0.001
R3688 vbias1.n255 vbias1.n254 0.001
R3689 vbias1.n233 vbias1.n232 0.001
R3690 vbias1.n211 vbias1.n210 0.001
R3691 vbias1.n189 vbias1.n188 0.001
R3692 vbias1.n167 vbias1.n166 0.001
R3693 vbias1.n145 vbias1.n144 0.001
R3694 vbias1.n123 vbias1.n122 0.001
R3695 vbias1.n101 vbias1.n100 0.001
R3696 vbias1.n89 vbias1.n88 0.001
R3697 vbias1.n111 vbias1.n110 0.001
R3698 vbias1.n133 vbias1.n132 0.001
R3699 vbias1.n155 vbias1.n154 0.001
R3700 vbias1.n177 vbias1.n176 0.001
R3701 vbias1.n199 vbias1.n198 0.001
R3702 vbias1.n221 vbias1.n220 0.001
R3703 vbias1.n243 vbias1.n242 0.001
R3704 vbias1.n265 vbias1.n264 0.001
R3705 vbias1.n288 vbias1.n287 0.001
R3706 vbias1.n396 vbias1.n395 0.001
R3707 vbias1.n356 vbias1.n355 0.001
R3708 vbias1.n344 vbias1.n343 0.001
R3709 vbias1.n316 vbias1.n315 0.001
R3710 vbias1.n676 vbias1.n675 0.001
R3711 vbias1.n36 vbias1.n35 0.001
R3712 vbias1.n409 vbias1.n408 0.001
R3713 vbias1.n454 vbias1.n453 0.001
R3714 vbias1.n478 vbias1.n477 0.001
R3715 vbias1.n490 vbias1.n489 0.001
R3716 vbias1.n514 vbias1.n513 0.001
R3717 vbias1.n526 vbias1.n525 0.001
R3718 vbias1.n550 vbias1.n549 0.001
R3719 vbias1.n562 vbias1.n561 0.001
R3720 vbias1.n586 vbias1.n585 0.001
R3721 vbias1.n598 vbias1.n597 0.001
R3722 vbias1.n622 vbias1.n621 0.001
R3723 vbias1.n634 vbias1.n633 0.001
R3724 vbias1.n658 vbias1.n657 0.001
R3725 vbias1.n671 vbias1.n670 0.001
R3726 a_23744_20184.n20 a_23744_20184.t18 278.182
R3727 a_23744_20184.n17 a_23744_20184.t12 278.182
R3728 a_23744_20184.n6 a_23744_20184.t20 278.182
R3729 a_23744_20184.n7 a_23744_20184.t23 278.182
R3730 a_23744_20184.n0 a_23744_20184.t14 276.116
R3731 a_23744_20184.n1 a_23744_20184.t16 276.116
R3732 a_23744_20184.n1 a_23744_20184.t22 276.116
R3733 a_23744_20184.n0 a_23744_20184.t21 276.116
R3734 a_23744_20184.n2 a_23744_20184.n0 127.197
R3735 a_23744_20184.n1 a_23744_20184.n3 127.197
R3736 a_23744_20184.n21 a_23744_20184.n20 127.197
R3737 a_23744_20184.n21 a_23744_20184.n9 121.282
R3738 a_23744_20184.n0 a_23744_20184.n1 22.632
R3739 a_23744_20184.n6 a_23744_20184.n5 22.181
R3740 a_23744_20184.n7 a_23744_20184.n6 22.181
R3741 a_23744_20184.n8 a_23744_20184.n7 22.181
R3742 a_23744_20184.n18 a_23744_20184.n17 22.181
R3743 a_23744_20184.n19 a_23744_20184.n18 22.181
R3744 a_23744_20184.n20 a_23744_20184.n19 22.181
R3745 a_23744_20184.n12 a_23744_20184.t1 7.146
R3746 a_23744_20184.n12 a_23744_20184.t9 7.146
R3747 a_23744_20184.n11 a_23744_20184.t11 7.146
R3748 a_23744_20184.n11 a_23744_20184.t8 7.146
R3749 a_23744_20184.n10 a_23744_20184.t5 7.146
R3750 a_23744_20184.n10 a_23744_20184.t0 7.146
R3751 a_23744_20184.n15 a_23744_20184.t4 7.146
R3752 a_23744_20184.n15 a_23744_20184.t10 7.146
R3753 a_23744_20184.n14 a_23744_20184.t7 7.146
R3754 a_23744_20184.n14 a_23744_20184.t6 7.146
R3755 a_23744_20184.n13 a_23744_20184.t3 7.146
R3756 a_23744_20184.n13 a_23744_20184.t2 7.146
R3757 a_23744_20184.n5 a_23744_20184.n4 5.915
R3758 a_23744_20184.n9 a_23744_20184.n8 5.915
R3759 a_23744_20184.n16 a_23744_20184.t13 5.801
R3760 a_23744_20184.n2 a_23744_20184.t15 5.801
R3761 a_23744_20184.n3 a_23744_20184.t17 5.801
R3762 a_23744_20184.t19 a_23744_20184.n21 5.801
R3763 a_23744_20184.n2 a_23744_20184.n12 3.315
R3764 a_23744_20184.n3 a_23744_20184.n15 3.278
R3765 a_23744_20184.n21 a_23744_20184.n2 1.365
R3766 a_23744_20184.n3 a_23744_20184.n16 1.313
R3767 a_23744_20184.n11 a_23744_20184.n10 0.827
R3768 a_23744_20184.n12 a_23744_20184.n11 0.827
R3769 a_23744_20184.n14 a_23744_20184.n13 0.827
R3770 a_23744_20184.n15 a_23744_20184.n14 0.827
R3771 a_23370_24650.n14 a_23370_24650.t8 8.207
R3772 a_23370_24650.n6 a_23370_24650.t3 8.207
R3773 a_23370_24650.n23 a_23370_24650.t25 7.146
R3774 a_23370_24650.n22 a_23370_24650.t30 7.146
R3775 a_23370_24650.n22 a_23370_24650.t4 7.146
R3776 a_23370_24650.n21 a_23370_24650.t24 7.146
R3777 a_23370_24650.n21 a_23370_24650.t9 7.146
R3778 a_23370_24650.n10 a_23370_24650.t18 7.146
R3779 a_23370_24650.n10 a_23370_24650.t14 7.146
R3780 a_23370_24650.n9 a_23370_24650.t19 7.146
R3781 a_23370_24650.n9 a_23370_24650.t16 7.146
R3782 a_23370_24650.n8 a_23370_24650.t20 7.146
R3783 a_23370_24650.n8 a_23370_24650.t17 7.146
R3784 a_23370_24650.n18 a_23370_24650.t12 7.146
R3785 a_23370_24650.n18 a_23370_24650.t21 7.146
R3786 a_23370_24650.n17 a_23370_24650.t13 7.146
R3787 a_23370_24650.n17 a_23370_24650.t22 7.146
R3788 a_23370_24650.n16 a_23370_24650.t23 7.146
R3789 a_23370_24650.n16 a_23370_24650.t15 7.146
R3790 a_23370_24650.n15 a_23370_24650.t7 7.146
R3791 a_23370_24650.n14 a_23370_24650.t10 7.146
R3792 a_23370_24650.n2 a_23370_24650.t34 7.146
R3793 a_23370_24650.n2 a_23370_24650.t32 7.146
R3794 a_23370_24650.n1 a_23370_24650.t27 7.146
R3795 a_23370_24650.n1 a_23370_24650.t26 7.146
R3796 a_23370_24650.n0 a_23370_24650.t35 7.146
R3797 a_23370_24650.n0 a_23370_24650.t33 7.146
R3798 a_23370_24650.n5 a_23370_24650.t0 7.146
R3799 a_23370_24650.n5 a_23370_24650.t28 7.146
R3800 a_23370_24650.n4 a_23370_24650.t5 7.146
R3801 a_23370_24650.n4 a_23370_24650.t31 7.146
R3802 a_23370_24650.n3 a_23370_24650.t1 7.146
R3803 a_23370_24650.n3 a_23370_24650.t29 7.146
R3804 a_23370_24650.n7 a_23370_24650.t2 7.146
R3805 a_23370_24650.n6 a_23370_24650.t6 7.146
R3806 a_23370_24650.t11 a_23370_24650.n23 7.146
R3807 a_23370_24650.n11 a_23370_24650.n10 1.938
R3808 a_23370_24650.n19 a_23370_24650.n18 1.938
R3809 a_23370_24650.n19 a_23370_24650.n15 1.493
R3810 a_23370_24650.n11 a_23370_24650.n7 1.493
R3811 a_23370_24650.n13 a_23370_24650.n2 1.386
R3812 a_23370_24650.n12 a_23370_24650.n5 1.386
R3813 a_23370_24650.n21 a_23370_24650.n20 1.386
R3814 a_23370_24650.n15 a_23370_24650.n14 1.061
R3815 a_23370_24650.n7 a_23370_24650.n6 1.061
R3816 a_23370_24650.n9 a_23370_24650.n8 0.865
R3817 a_23370_24650.n10 a_23370_24650.n9 0.865
R3818 a_23370_24650.n17 a_23370_24650.n16 0.865
R3819 a_23370_24650.n18 a_23370_24650.n17 0.865
R3820 a_23370_24650.n12 a_23370_24650.n11 0.831
R3821 a_23370_24650.n13 a_23370_24650.n12 0.831
R3822 a_23370_24650.n20 a_23370_24650.n13 0.831
R3823 a_23370_24650.n20 a_23370_24650.n19 0.831
R3824 a_23370_24650.n1 a_23370_24650.n0 0.827
R3825 a_23370_24650.n2 a_23370_24650.n1 0.827
R3826 a_23370_24650.n4 a_23370_24650.n3 0.827
R3827 a_23370_24650.n5 a_23370_24650.n4 0.827
R3828 a_23370_24650.n22 a_23370_24650.n21 0.827
R3829 a_23370_24650.n23 a_23370_24650.n22 0.827
R3830 a_23744_3840.n18 a_23744_3840.t14 278.182
R3831 a_23744_3840.n21 a_23744_3840.t18 278.182
R3832 a_23744_3840.n20 a_23744_3840.t23 278.182
R3833 a_23744_3840.n19 a_23744_3840.t22 278.182
R3834 a_23744_3840.n13 a_23744_3840.t12 276.116
R3835 a_23744_3840.n16 a_23744_3840.t16 276.116
R3836 a_23744_3840.n15 a_23744_3840.t21 276.116
R3837 a_23744_3840.n14 a_23744_3840.t20 276.116
R3838 a_23744_3840.n13 a_23744_3840.n0 127.197
R3839 a_23744_3840.n1 a_23744_3840.n16 127.197
R3840 a_23744_3840.n8 a_23744_3840.n7 127.197
R3841 a_23744_3840.n1 a_23744_3840.n22 121.282
R3842 a_23744_3840.n15 a_23744_3840.n14 22.181
R3843 a_23744_3840.n21 a_23744_3840.n20 22.181
R3844 a_23744_3840.n20 a_23744_3840.n19 22.181
R3845 a_23744_3840.n19 a_23744_3840.n18 22.181
R3846 a_23744_3840.n7 a_23744_3840.n6 22.181
R3847 a_23744_3840.n6 a_23744_3840.n5 22.181
R3848 a_23744_3840.n5 a_23744_3840.n4 22.181
R3849 a_23744_3840.n23 a_23744_3840.t10 7.146
R3850 a_23744_3840.n3 a_23744_3840.t2 7.146
R3851 a_23744_3840.n3 a_23744_3840.t3 7.146
R3852 a_23744_3840.n2 a_23744_3840.t6 7.146
R3853 a_23744_3840.n2 a_23744_3840.t7 7.146
R3854 a_23744_3840.n11 a_23744_3840.t5 7.146
R3855 a_23744_3840.n11 a_23744_3840.t8 7.146
R3856 a_23744_3840.n10 a_23744_3840.t9 7.146
R3857 a_23744_3840.n10 a_23744_3840.t0 7.146
R3858 a_23744_3840.n9 a_23744_3840.t4 7.146
R3859 a_23744_3840.n9 a_23744_3840.t1 7.146
R3860 a_23744_3840.t11 a_23744_3840.n23 7.146
R3861 a_23744_3840.n22 a_23744_3840.n21 5.915
R3862 a_23744_3840.n18 a_23744_3840.n17 5.915
R3863 a_23744_3840.n8 a_23744_3840.t19 5.801
R3864 a_23744_3840.n12 a_23744_3840.t15 5.801
R3865 a_23744_3840.n0 a_23744_3840.t13 5.801
R3866 a_23744_3840.n1 a_23744_3840.t17 5.801
R3867 a_23744_3840.n0 a_23744_3840.n11 3.315
R3868 a_23744_3840.n23 a_23744_3840.n1 3.278
R3869 a_23744_3840.n0 a_23744_3840.n12 1.365
R3870 a_23744_3840.n1 a_23744_3840.n8 1.313
R3871 a_23744_3840.n3 a_23744_3840.n2 0.827
R3872 a_23744_3840.n23 a_23744_3840.n3 0.827
R3873 a_23744_3840.n10 a_23744_3840.n9 0.827
R3874 a_23744_3840.n11 a_23744_3840.n10 0.827
R3875 a_23744_3840.n14 a_23744_3840.n13 0.226
R3876 a_23744_3840.n16 a_23744_3840.n15 0.226
C16 a_30793_4721# vss 9.53fF
C17 vbias1 vss 92.36fF
C18 a_30831_20339# vss 7.40fF
C19 vt vss 151.29fF
C20 vref vss 101.71fF
C21 OTA_0/vp vss 16.15fF
C22 vbias2 vss 89.96fF
C23 OTA_tri_0/vn vss 91.85fF
C24 vsquare vss 132.70fF
C25 vdd vss 1007.47fF
C26 a_23744_3840.n0 vss 1.56fF $ **FLOATING
C27 a_23744_3840.n1 vss 1.59fF $ **FLOATING
C28 a_23744_3840.n2 vss 2.69fF $ **FLOATING
C29 a_23744_3840.n3 vss 2.78fF $ **FLOATING
C30 a_23744_3840.n9 vss 2.69fF $ **FLOATING
C31 a_23744_3840.n10 vss 2.78fF $ **FLOATING
C32 a_23744_3840.n11 vss 3.35fF $ **FLOATING
C33 a_23744_3840.n23 vss 3.34fF $ **FLOATING
C34 a_23370_24650.n0 vss 2.20fF $ **FLOATING
C35 a_23370_24650.n1 vss 2.27fF $ **FLOATING
C36 a_23370_24650.n2 vss 2.32fF $ **FLOATING
C37 a_23370_24650.n3 vss 2.20fF $ **FLOATING
C38 a_23370_24650.n4 vss 2.27fF $ **FLOATING
C39 a_23370_24650.n5 vss 2.32fF $ **FLOATING
C40 a_23370_24650.n6 vss 2.65fF $ **FLOATING
C41 a_23370_24650.n7 vss 1.50fF $ **FLOATING
C42 a_23370_24650.n8 vss 2.14fF $ **FLOATING
C43 a_23370_24650.n9 vss 2.20fF $ **FLOATING
C44 a_23370_24650.n10 vss 2.33fF $ **FLOATING
C45 a_23370_24650.n14 vss 2.65fF $ **FLOATING
C46 a_23370_24650.n15 vss 1.50fF $ **FLOATING
C47 a_23370_24650.n16 vss 2.14fF $ **FLOATING
C48 a_23370_24650.n17 vss 2.20fF $ **FLOATING
C49 a_23370_24650.n18 vss 2.33fF $ **FLOATING
C50 a_23370_24650.n21 vss 2.32fF $ **FLOATING
C51 a_23370_24650.n22 vss 2.27fF $ **FLOATING
C52 a_23370_24650.n23 vss 2.20fF $ **FLOATING
C53 a_23744_20184.n0 vss 1.44fF $ **FLOATING
C54 a_23744_20184.n1 vss 1.44fF $ **FLOATING
C55 a_23744_20184.n2 vss 1.67fF $ **FLOATING
C56 a_23744_20184.n3 vss 1.70fF $ **FLOATING
C57 a_23744_20184.n10 vss 2.88fF $ **FLOATING
C58 a_23744_20184.n11 vss 2.97fF $ **FLOATING
C59 a_23744_20184.n12 vss 3.58fF $ **FLOATING
C60 a_23744_20184.n13 vss 2.88fF $ **FLOATING
C61 a_23744_20184.n14 vss 2.97fF $ **FLOATING
C62 a_23744_20184.n15 vss 3.57fF $ **FLOATING
C63 a_23744_20184.n16 vss 1.03fF $ **FLOATING
C64 vbias1.n84 vss 1.09fF $ **FLOATING
C65 a_23370_8306.n0 vss 2.67fF $ **FLOATING
C66 a_23370_8306.n1 vss 1.50fF $ **FLOATING
C67 a_23370_8306.n2 vss 2.15fF $ **FLOATING
C68 a_23370_8306.n3 vss 2.21fF $ **FLOATING
C69 a_23370_8306.n4 vss 2.34fF $ **FLOATING
C70 a_23370_8306.n6 vss 2.21fF $ **FLOATING
C71 a_23370_8306.n7 vss 2.28fF $ **FLOATING
C72 a_23370_8306.n8 vss 2.33fF $ **FLOATING
C73 a_23370_8306.n9 vss 2.21fF $ **FLOATING
C74 a_23370_8306.n10 vss 2.28fF $ **FLOATING
C75 a_23370_8306.n11 vss 2.33fF $ **FLOATING
C76 a_23370_8306.n12 vss 2.67fF $ **FLOATING
C77 a_23370_8306.n13 vss 1.50fF $ **FLOATING
C78 a_23370_8306.n14 vss 2.15fF $ **FLOATING
C79 a_23370_8306.n15 vss 2.21fF $ **FLOATING
C80 a_23370_8306.n16 vss 2.34fF $ **FLOATING
C81 a_23370_8306.n21 vss 2.21fF $ **FLOATING
C82 a_23370_8306.n22 vss 2.28fF $ **FLOATING
C83 a_23370_8306.n23 vss 2.33fF $ **FLOATING
C84 vref.n34 vss 10.93fF $ **FLOATING
C85 vref.n35 vss 14.94fF $ **FLOATING
C86 vdd.n0 vss 7.61fF $ **FLOATING
C87 vdd.n1 vss 1.61fF $ **FLOATING
C88 vdd.n2 vss 1.66fF $ **FLOATING
C89 vdd.n3 vss 1.59fF $ **FLOATING
C90 vdd.n4 vss 1.61fF $ **FLOATING
C91 vdd.n5 vss 1.66fF $ **FLOATING
C92 vdd.n6 vss 1.59fF $ **FLOATING
C93 vdd.n10 vss 1.61fF $ **FLOATING
C94 vdd.n11 vss 1.66fF $ **FLOATING
C95 vdd.n12 vss 1.59fF $ **FLOATING
C96 vdd.n13 vss 1.61fF $ **FLOATING
C97 vdd.n14 vss 1.66fF $ **FLOATING
C98 vdd.n15 vss 1.59fF $ **FLOATING
C99 vdd.n19 vss 1.61fF $ **FLOATING
C100 vdd.n20 vss 1.66fF $ **FLOATING
C101 vdd.n21 vss 1.59fF $ **FLOATING
C102 vdd.n22 vss 1.61fF $ **FLOATING
C103 vdd.n23 vss 1.66fF $ **FLOATING
C104 vdd.n24 vss 1.59fF $ **FLOATING
C105 vdd.n28 vss 1.61fF $ **FLOATING
C106 vdd.n29 vss 1.66fF $ **FLOATING
C107 vdd.n30 vss 1.59fF $ **FLOATING
C108 vdd.n31 vss 1.61fF $ **FLOATING
C109 vdd.n32 vss 1.66fF $ **FLOATING
C110 vdd.n33 vss 1.59fF $ **FLOATING
C111 vdd.n37 vss 1.61fF $ **FLOATING
C112 vdd.n38 vss 1.66fF $ **FLOATING
C113 vdd.n39 vss 1.59fF $ **FLOATING
C114 vdd.n40 vss 1.61fF $ **FLOATING
C115 vdd.n41 vss 1.66fF $ **FLOATING
C116 vdd.n42 vss 1.59fF $ **FLOATING
C117 vdd.n46 vss 1.61fF $ **FLOATING
C118 vdd.n47 vss 1.66fF $ **FLOATING
C119 vdd.n48 vss 1.59fF $ **FLOATING
C120 vdd.n49 vss 1.61fF $ **FLOATING
C121 vdd.n50 vss 1.66fF $ **FLOATING
C122 vdd.n51 vss 1.60fF $ **FLOATING
C123 vdd.n55 vss 3.65fF $ **FLOATING
C124 vdd.n56 vss 1.61fF $ **FLOATING
C125 vdd.n57 vss 1.66fF $ **FLOATING
C126 vdd.n58 vss 1.60fF $ **FLOATING
C127 vdd.n62 vss 3.65fF $ **FLOATING
C128 vdd.n63 vss 1.61fF $ **FLOATING
C129 vdd.n64 vss 1.66fF $ **FLOATING
C130 vdd.n65 vss 1.59fF $ **FLOATING
C131 vdd.n69 vss 1.61fF $ **FLOATING
C132 vdd.n70 vss 1.66fF $ **FLOATING
C133 vdd.n71 vss 1.59fF $ **FLOATING
C134 vdd.n72 vss 1.61fF $ **FLOATING
C135 vdd.n73 vss 1.66fF $ **FLOATING
C136 vdd.n74 vss 1.59fF $ **FLOATING
C137 vdd.n75 vss 1.61fF $ **FLOATING
C138 vdd.n76 vss 1.66fF $ **FLOATING
C139 vdd.n77 vss 1.59fF $ **FLOATING
C140 vdd.n82 vss 1.61fF $ **FLOATING
C141 vdd.n83 vss 1.66fF $ **FLOATING
C142 vdd.n84 vss 1.59fF $ **FLOATING
C143 vdd.n85 vss 1.61fF $ **FLOATING
C144 vdd.n86 vss 1.66fF $ **FLOATING
C145 vdd.n87 vss 1.59fF $ **FLOATING
C146 vdd.n90 vss 1.61fF $ **FLOATING
C147 vdd.n91 vss 1.66fF $ **FLOATING
C148 vdd.n92 vss 1.59fF $ **FLOATING
C149 vdd.n95 vss 1.61fF $ **FLOATING
C150 vdd.n96 vss 1.66fF $ **FLOATING
C151 vdd.n97 vss 1.59fF $ **FLOATING
C152 vdd.n98 vss 1.61fF $ **FLOATING
C153 vdd.n99 vss 1.66fF $ **FLOATING
C154 vdd.n100 vss 1.59fF $ **FLOATING
C155 vdd.n104 vss 1.61fF $ **FLOATING
C156 vdd.n105 vss 1.66fF $ **FLOATING
C157 vdd.n106 vss 1.59fF $ **FLOATING
C158 vdd.n107 vss 7.61fF $ **FLOATING
C159 vdd.n108 vss 1.61fF $ **FLOATING
C160 vdd.n109 vss 1.66fF $ **FLOATING
C161 vdd.n110 vss 1.59fF $ **FLOATING
C162 vdd.n111 vss 1.61fF $ **FLOATING
C163 vdd.n112 vss 1.66fF $ **FLOATING
C164 vdd.n113 vss 1.59fF $ **FLOATING
C165 vdd.n116 vss 1.61fF $ **FLOATING
C166 vdd.n117 vss 1.66fF $ **FLOATING
C167 vdd.n118 vss 1.59fF $ **FLOATING
C168 vdd.n120 vss 1.61fF $ **FLOATING
C169 vdd.n121 vss 1.66fF $ **FLOATING
C170 vdd.n122 vss 1.59fF $ **FLOATING
C171 vdd.n123 vss 1.61fF $ **FLOATING
C172 vdd.n124 vss 1.66fF $ **FLOATING
C173 vdd.n125 vss 1.59fF $ **FLOATING
C174 vdd.n128 vss 1.61fF $ **FLOATING
C175 vdd.n129 vss 1.66fF $ **FLOATING
C176 vdd.n130 vss 1.59fF $ **FLOATING
C177 vdd.n132 vss 1.61fF $ **FLOATING
C178 vdd.n133 vss 1.66fF $ **FLOATING
C179 vdd.n134 vss 1.59fF $ **FLOATING
C180 vdd.n136 vss 1.61fF $ **FLOATING
C181 vdd.n137 vss 1.66fF $ **FLOATING
C182 vdd.n138 vss 1.59fF $ **FLOATING
C183 vdd.n139 vss 1.61fF $ **FLOATING
C184 vdd.n140 vss 1.66fF $ **FLOATING
C185 vdd.n141 vss 1.59fF $ **FLOATING
C186 vdd.n144 vss 1.61fF $ **FLOATING
C187 vdd.n145 vss 1.66fF $ **FLOATING
C188 vdd.n146 vss 1.59fF $ **FLOATING
C189 vdd.n148 vss 1.61fF $ **FLOATING
C190 vdd.n149 vss 1.66fF $ **FLOATING
C191 vdd.n150 vss 1.59fF $ **FLOATING
C192 vdd.n152 vss 1.61fF $ **FLOATING
C193 vdd.n153 vss 1.66fF $ **FLOATING
C194 vdd.n154 vss 1.59fF $ **FLOATING
C195 vdd.n155 vss 1.61fF $ **FLOATING
C196 vdd.n156 vss 1.66fF $ **FLOATING
C197 vdd.n157 vss 1.60fF $ **FLOATING
C198 vdd.n159 vss 3.65fF $ **FLOATING
C199 vdd.n160 vss 1.61fF $ **FLOATING
C200 vdd.n161 vss 1.66fF $ **FLOATING
C201 vdd.n162 vss 1.60fF $ **FLOATING
C202 vdd.n164 vss 3.65fF $ **FLOATING
C203 vdd.n170 vss 1.61fF $ **FLOATING
C204 vdd.n171 vss 1.66fF $ **FLOATING
C205 vdd.n172 vss 1.59fF $ **FLOATING
C206 vdd.n174 vss 1.61fF $ **FLOATING
C207 vdd.n175 vss 1.66fF $ **FLOATING
C208 vdd.n176 vss 1.59fF $ **FLOATING
C209 vdd.n178 vss 1.61fF $ **FLOATING
C210 vdd.n179 vss 1.66fF $ **FLOATING
C211 vdd.n180 vss 1.59fF $ **FLOATING
C212 vdd.n182 vss 1.61fF $ **FLOATING
C213 vdd.n183 vss 1.66fF $ **FLOATING
C214 vdd.n184 vss 1.59fF $ **FLOATING
C215 vdd.n186 vss 1.61fF $ **FLOATING
C216 vdd.n187 vss 1.66fF $ **FLOATING
C217 vdd.n188 vss 1.59fF $ **FLOATING
C218 vdd.n190 vss 1.61fF $ **FLOATING
C219 vdd.n191 vss 1.66fF $ **FLOATING
C220 vdd.n192 vss 1.59fF $ **FLOATING
C221 vdd.n194 vss 1.61fF $ **FLOATING
C222 vdd.n195 vss 1.66fF $ **FLOATING
C223 vdd.n196 vss 1.59fF $ **FLOATING
C224 vdd.n198 vss 1.61fF $ **FLOATING
C225 vdd.n199 vss 1.66fF $ **FLOATING
C226 vdd.n200 vss 1.59fF $ **FLOATING
C227 vdd.n202 vss 1.61fF $ **FLOATING
C228 vdd.n203 vss 1.66fF $ **FLOATING
C229 vdd.n204 vss 1.59fF $ **FLOATING
C230 vdd.n206 vss 1.61fF $ **FLOATING
C231 vdd.n207 vss 1.66fF $ **FLOATING
C232 vdd.n208 vss 1.59fF $ **FLOATING
C233 vdd.n209 vss 7.61fF $ **FLOATING
C234 vdd.n210 vss 7.61fF $ **FLOATING
C235 vdd.n211 vss 1.61fF $ **FLOATING
C236 vdd.n212 vss 1.66fF $ **FLOATING
C237 vdd.n213 vss 1.59fF $ **FLOATING
C238 vdd.n214 vss 14.83fF $ **FLOATING
C239 vdd.n215 vss 11.39fF $ **FLOATING
C240 vdd.n216 vss 11.39fF $ **FLOATING
C241 vdd.n217 vss 11.39fF $ **FLOATING
C242 vdd.n218 vss 11.39fF $ **FLOATING
C243 vdd.n219 vss 11.39fF $ **FLOATING
C244 vdd.n220 vss 11.39fF $ **FLOATING
C245 vdd.n221 vss 11.39fF $ **FLOATING
C246 vdd.n222 vss 11.39fF $ **FLOATING
C247 vdd.n223 vss 11.39fF $ **FLOATING
C248 vdd.n224 vss 11.39fF $ **FLOATING
C249 vdd.n225 vss 10.96fF $ **FLOATING
C250 vdd.n226 vss 10.96fF $ **FLOATING
C251 vdd.n227 vss 11.39fF $ **FLOATING
C252 vdd.n228 vss 11.39fF $ **FLOATING
C253 vdd.n229 vss 16.69fF $ **FLOATING
C254 vdd.n230 vss 16.69fF $ **FLOATING
C255 vdd.n231 vss 11.39fF $ **FLOATING
C256 vdd.n232 vss 16.68fF $ **FLOATING
C257 vdd.n233 vss 16.68fF $ **FLOATING
C258 vdd.n234 vss 11.39fF $ **FLOATING
C259 vdd.n235 vss 22.60fF $ **FLOATING
C260 vdd.n236 vss 95.23fF $ **FLOATING
C261 vdd.n237 vss 11.39fF $ **FLOATING
C262 vdd.n238 vss 16.23fF $ **FLOATING
C263 vdd.n239 vss 16.68fF $ **FLOATING
C264 vdd.n240 vss 10.94fF $ **FLOATING
C265 vdd.n241 vss 16.69fF $ **FLOATING
C266 vdd.n242 vss 16.23fF $ **FLOATING
C267 vdd.n243 vss 11.39fF $ **FLOATING
C268 vdd.n244 vss 10.94fF $ **FLOATING
C269 vdd.n245 vss 10.96fF $ **FLOATING
C270 vdd.n246 vss 10.96fF $ **FLOATING
C271 vdd.n247 vss 11.39fF $ **FLOATING
C272 vdd.n248 vss 10.94fF $ **FLOATING
C273 vdd.n249 vss 11.39fF $ **FLOATING
C274 vdd.n250 vss 10.94fF $ **FLOATING
C275 vdd.n251 vss 11.39fF $ **FLOATING
C276 vdd.n252 vss 10.94fF $ **FLOATING
C277 vdd.n253 vss 11.39fF $ **FLOATING
C278 vdd.n254 vss 10.94fF $ **FLOATING
C279 vdd.n255 vss 11.39fF $ **FLOATING
C280 vdd.n256 vss 10.94fF $ **FLOATING
C281 vdd.n257 vss 13.54fF $ **FLOATING
C282 vsquare.n2 vss 1.04fF $ **FLOATING
C283 vsquare.n3 vss 1.18fF $ **FLOATING
C284 vsquare.n5 vss 3.59fF $ **FLOATING
C285 vsquare.n6 vss 2.40fF $ **FLOATING
C286 vsquare.n9 vss 1.04fF $ **FLOATING
C287 vsquare.n12 vss 1.04fF $ **FLOATING
C288 vsquare.n15 vss 1.04fF $ **FLOATING
C289 vsquare.n18 vss 1.04fF $ **FLOATING
C290 vsquare.n21 vss 1.04fF $ **FLOATING
C291 vsquare.n24 vss 1.04fF $ **FLOATING
C292 vsquare.n28 vss 1.04fF $ **FLOATING
C293 vsquare.n35 vss 1.04fF $ **FLOATING
C294 vsquare.n72 vss 1.04fF $ **FLOATING
C295 vsquare.n79 vss 1.04fF $ **FLOATING
C296 vsquare.n83 vss 1.04fF $ **FLOATING
C297 vsquare.n86 vss 1.04fF $ **FLOATING
C298 vsquare.n89 vss 1.04fF $ **FLOATING
C299 vsquare.n92 vss 1.04fF $ **FLOATING
C300 vsquare.n95 vss 1.04fF $ **FLOATING
C301 vsquare.n98 vss 1.04fF $ **FLOATING
C302 vsquare.n101 vss 1.04fF $ **FLOATING
C303 vsquare.n102 vss 1.18fF $ **FLOATING
C304 vsquare.n104 vss 8.83fF $ **FLOATING
C305 vsquare.n105 vss 3.71fF $ **FLOATING
C306 vsquare.n106 vss 3.71fF $ **FLOATING
C307 vsquare.n107 vss 3.71fF $ **FLOATING
C308 vsquare.n108 vss 3.71fF $ **FLOATING
C309 vsquare.n109 vss 3.71fF $ **FLOATING
C310 vsquare.n110 vss 3.71fF $ **FLOATING
C311 vsquare.n111 vss 3.56fF $ **FLOATING
C312 vsquare.n112 vss 1.90fF $ **FLOATING
C313 vsquare.n114 vss 1.41fF $ **FLOATING
C314 vsquare.n115 vss 1.30fF $ **FLOATING
C315 vsquare.n117 vss 1.08fF $ **FLOATING
C316 vsquare.n118 vss 1.55fF $ **FLOATING
C317 vsquare.n121 vss 1.52fF $ **FLOATING
C318 vsquare.n122 vss 1.55fF $ **FLOATING
C319 vsquare.n123 vss 1.55fF $ **FLOATING
C320 vsquare.n124 vss 1.55fF $ **FLOATING
C321 vsquare.n125 vss 1.55fF $ **FLOATING
C322 vsquare.n126 vss 1.55fF $ **FLOATING
C323 vsquare.n127 vss 1.55fF $ **FLOATING
C324 vsquare.n128 vss 1.55fF $ **FLOATING
C325 vsquare.n129 vss 1.52fF $ **FLOATING
C326 vsquare.n132 vss 1.55fF $ **FLOATING
C327 vsquare.n133 vss 1.08fF $ **FLOATING
C328 vsquare.n135 vss 1.30fF $ **FLOATING
C329 vsquare.n136 vss 1.40fF $ **FLOATING
C330 vsquare.n138 vss 1.90fF $ **FLOATING
C331 vsquare.n139 vss 3.55fF $ **FLOATING
C332 vsquare.n140 vss 3.71fF $ **FLOATING
C333 vsquare.n141 vss 3.71fF $ **FLOATING
C334 vsquare.n142 vss 41.58fF $ **FLOATING
C335 vsquare.n143 vss 14.99fF $ **FLOATING
C336 vsquare.n144 vss 3.19fF $ **FLOATING
C337 a_19926_29936.n0 vss 2.85fF $ **FLOATING
C338 a_19926_29936.n1 vss 1.99fF $ **FLOATING
C339 a_19926_29936.n2 vss 4.18fF $ **FLOATING
C340 a_19926_29936.n3 vss 1.99fF $ **FLOATING
C341 a_19926_29936.n4 vss 4.18fF $ **FLOATING
C342 a_19926_29936.n5 vss 5.60fF $ **FLOATING
C343 a_19926_29936.n6 vss 7.19fF $ **FLOATING
C344 a_19926_29936.n7 vss 5.60fF $ **FLOATING
C345 a_19926_29936.n8 vss 5.60fF $ **FLOATING
C346 a_19926_29936.n9 vss 4.03fF $ **FLOATING
C347 a_19926_29936.n10 vss 6.10fF $ **FLOATING
C348 a_19926_29936.n11 vss 7.82fF $ **FLOATING
C349 a_19926_29936.n12 vss 6.10fF $ **FLOATING
C350 a_19926_29936.n13 vss 6.10fF $ **FLOATING
C351 a_19926_29936.n14 vss 4.41fF $ **FLOATING
C352 a_19926_29936.n15 vss 46.82fF $ **FLOATING
C353 a_19926_29936.n16 vss 4.47fF $ **FLOATING
C354 a_19926_29936.n17 vss 17.93fF $ **FLOATING
C355 vt.n5 vss 1.45fF $ **FLOATING
C356 vt.n6 vss 1.58fF $ **FLOATING
C357 vt.n103 vss 12.15fF $ **FLOATING
C358 vt.n104 vss 452.58fF $ **FLOATING
C359 vt.n105 vss 2.45fF $ **FLOATING
C360 vt.n106 vss 2.45fF $ **FLOATING
C361 vt.n107 vss 2.45fF $ **FLOATING
C362 vt.n108 vss 2.45fF $ **FLOATING
C363 vt.n109 vss 2.45fF $ **FLOATING
C364 vt.n110 vss 2.35fF $ **FLOATING
C365 vt.n111 vss 1.26fF $ **FLOATING
C366 vt.n117 vss 1.03fF $ **FLOATING
C367 vt.n120 vss 1.01fF $ **FLOATING
C368 vt.n121 vss 1.03fF $ **FLOATING
C369 vt.n122 vss 1.03fF $ **FLOATING
C370 vt.n123 vss 1.03fF $ **FLOATING
C371 vt.n124 vss 1.03fF $ **FLOATING
C372 vt.n125 vss 1.03fF $ **FLOATING
C373 vt.n126 vss 1.03fF $ **FLOATING
C374 vt.n127 vss 1.03fF $ **FLOATING
C375 vt.n128 vss 1.00fF $ **FLOATING
C376 vt.n131 vss 1.03fF $ **FLOATING
C377 vt.n137 vss 1.26fF $ **FLOATING
C378 vt.n138 vss 2.35fF $ **FLOATING
C379 vt.n139 vss 2.45fF $ **FLOATING
C380 vt.n140 vss 2.45fF $ **FLOATING
C381 vt.n141 vss 33.12fF $ **FLOATING
C382 vt.n142 vss 11.43fF $ **FLOATING
C383 vt.n143 vss 2.15fF $ **FLOATING
C384 a_19926_13536.n0 vss 2.72fF $ **FLOATING
C385 a_19926_13536.n1 vss 1.91fF $ **FLOATING
C386 a_19926_13536.n2 vss 4.00fF $ **FLOATING
C387 a_19926_13536.n3 vss 1.91fF $ **FLOATING
C388 a_19926_13536.n4 vss 4.00fF $ **FLOATING
C389 a_19926_13536.n5 vss 5.36fF $ **FLOATING
C390 a_19926_13536.n6 vss 6.88fF $ **FLOATING
C391 a_19926_13536.n7 vss 5.36fF $ **FLOATING
C392 a_19926_13536.n8 vss 5.36fF $ **FLOATING
C393 a_19926_13536.n9 vss 3.86fF $ **FLOATING
C394 a_19926_13536.n10 vss 5.83fF $ **FLOATING
C395 a_19926_13536.n11 vss 7.48fF $ **FLOATING
C396 a_19926_13536.n12 vss 5.83fF $ **FLOATING
C397 a_19926_13536.n13 vss 5.83fF $ **FLOATING
C398 a_19926_13536.n14 vss 4.22fF $ **FLOATING
C399 a_19926_13536.n15 vss 44.47fF $ **FLOATING
C400 a_19926_13536.n16 vss 4.18fF $ **FLOATING
C401 a_19926_13536.n17 vss 24.71fF $ **FLOATING
.ends
