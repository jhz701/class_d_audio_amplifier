magic
tech sky130A
magscale 1 2
timestamp 1627227727
<< nwell >>
rect 11200 27492 11620 27570
rect 11788 27492 12208 27570
rect 12376 27492 12796 27570
rect 12964 27492 13384 27570
rect 13552 27492 13972 27570
rect 14140 27492 14560 27570
rect 14728 27492 15148 27570
rect 15316 27492 15736 27570
rect 15904 27492 16324 27570
rect 16492 27492 16912 27570
rect 17080 27492 17500 27570
rect 17668 27492 18088 27570
rect 18256 27492 18676 27570
rect 18844 27492 19264 27570
rect 19432 27492 19852 27570
rect 20020 27492 20440 27570
rect 20608 27492 21028 27570
rect 21196 27492 21616 27570
rect 22974 27490 23366 27564
rect 23562 27490 23954 27564
rect 24150 27490 24542 27564
rect 24738 27490 25130 27564
rect 25326 27490 25718 27564
rect 25914 27490 26306 27564
rect 26502 27490 26894 27564
rect 27090 27490 27482 27564
rect 27678 27490 28070 27564
rect 28266 27490 28658 27564
rect 28854 27490 29246 27564
rect 29442 27490 29834 27564
rect 30030 27490 30422 27564
rect 30618 27490 31010 27564
rect 31206 27490 31598 27564
rect 31794 27490 32186 27564
rect 32382 27490 32774 27564
rect 32970 27490 33362 27564
rect 33558 27490 33950 27564
rect 34146 27490 34538 27564
rect 34734 27490 35126 27564
rect 35322 27490 35714 27564
rect 35910 27490 36302 27564
rect 36498 27490 36890 27564
rect 37086 27490 37478 27564
rect 37674 27490 38066 27564
rect 38262 27490 38654 27564
rect 11214 26492 11606 26626
rect 11802 26492 12194 26626
rect 12390 26492 12782 26626
rect 12978 26492 13370 26626
rect 13566 26492 13958 26626
rect 14154 26492 14546 26626
rect 14742 26492 15134 26626
rect 15330 26492 15722 26626
rect 15918 26492 16310 26626
rect 16506 26492 16898 26626
rect 17094 26492 17486 26626
rect 17682 26492 18074 26626
rect 18270 26492 18662 26626
rect 18858 26492 19250 26626
rect 19446 26492 19838 26626
rect 20034 26492 20426 26626
rect 20622 26492 21014 26626
rect 21210 26492 21602 26626
rect 21798 26492 22190 26626
rect 22974 26498 23354 26626
rect 23562 26498 23942 26626
rect 24150 26498 24530 26626
rect 24738 26498 25118 26626
rect 25326 26498 25706 26626
rect 25914 26498 26294 26626
rect 26502 26498 26882 26626
rect 27090 26498 27470 26626
rect 27678 26498 28058 26626
rect 28266 26498 28646 26626
rect 28854 26498 29234 26626
rect 29442 26498 29822 26626
rect 30030 26498 30410 26626
rect 30618 26498 30998 26626
rect 31206 26498 31586 26626
rect 31794 26498 32174 26626
rect 32382 26498 32762 26626
rect 32970 26498 33350 26626
rect 33558 26498 33938 26626
rect 34146 26498 34526 26626
rect 34734 26498 35114 26626
rect 35322 26498 35702 26626
rect 35910 26498 36290 26626
rect 36498 26498 36878 26626
rect 37086 26498 37466 26626
rect 37674 26498 38054 26626
rect 38262 26498 38642 26626
rect 10638 25498 11006 25626
rect 11226 25498 11594 25626
rect 11814 25498 12182 25626
rect 12402 25498 12770 25626
rect 12990 25498 13358 25626
rect 13578 25498 13946 25626
rect 14166 25498 14534 25626
rect 14754 25498 15122 25626
rect 15342 25498 15710 25626
rect 15930 25498 16298 25626
rect 16518 25498 16886 25626
rect 17106 25498 17474 25626
rect 17694 25498 18062 25626
rect 18282 25498 18650 25626
rect 18870 25498 19238 25626
rect 19458 25498 19826 25626
rect 20046 25498 20414 25626
rect 20634 25498 21002 25626
rect 21222 25498 21590 25626
rect 21810 25498 22178 25626
rect 23574 25496 23942 25628
rect 24162 25496 24530 25628
rect 24750 25496 25118 25628
rect 25338 25496 25706 25628
rect 25926 25496 26294 25628
rect 26514 25496 26882 25628
rect 27102 25496 27470 25628
rect 27690 25496 28058 25628
rect 28278 25496 28646 25628
rect 28866 25496 29234 25628
rect 29454 25496 29822 25628
rect 30042 25496 30410 25628
rect 30630 25496 30998 25628
rect 31218 25496 31586 25628
rect 31806 25496 32174 25628
rect 32394 25496 32762 25628
rect 32982 25496 33350 25628
rect 33570 25496 33938 25628
rect 34158 25496 34526 25628
rect 34746 25496 35114 25628
rect 35334 25496 35702 25628
rect 35922 25496 36290 25628
rect 36510 25496 36878 25628
rect 37098 25496 37466 25628
rect 37686 25496 38054 25628
rect 38274 25496 38642 25628
rect 11210 24562 11594 24634
rect 11798 24562 12182 24634
rect 12386 24562 12770 24634
rect 12974 24562 13358 24634
rect 13562 24562 13946 24634
rect 14150 24562 14534 24634
rect 14738 24562 15122 24634
rect 15326 24562 15710 24634
rect 15914 24562 16298 24634
rect 16502 24562 16886 24634
rect 17090 24562 17474 24634
rect 17678 24562 18062 24634
rect 18266 24562 18650 24634
rect 18854 24562 19238 24634
rect 19442 24562 19826 24634
rect 20030 24562 20414 24634
rect 20618 24562 21002 24634
rect 21206 24562 21590 24634
rect 21794 24562 22178 24634
rect 22986 24556 23354 24644
rect 23574 24556 23942 24644
rect 24162 24556 24530 24644
rect 24750 24556 25118 24644
rect 25338 24556 25706 24644
rect 25926 24556 26294 24644
rect 26514 24556 26882 24644
rect 27102 24556 27470 24644
rect 27690 24556 28058 24644
rect 28278 24556 28646 24644
rect 28866 24556 29234 24644
rect 29454 24556 29822 24644
rect 30042 24556 30410 24644
rect 30630 24556 30998 24644
rect 31218 24556 31586 24644
rect 31806 24556 32174 24644
rect 32394 24556 32762 24644
rect 32982 24556 33350 24644
rect 33570 24556 33938 24644
rect 34158 24556 34526 24644
rect 34746 24556 35114 24644
rect 35334 24556 35702 24644
rect 35922 24556 36290 24644
rect 36510 24556 36878 24644
rect 37098 24556 37466 24644
rect 37686 24556 38054 24644
rect 38274 24556 38642 24644
rect 11226 11134 11594 11206
rect 11814 11134 12182 11206
rect 12402 11134 12770 11206
rect 12990 11134 13358 11206
rect 13578 11134 13946 11206
rect 14166 11134 14534 11206
rect 14754 11134 15122 11206
rect 15342 11134 15710 11206
rect 15930 11134 16298 11206
rect 16518 11134 16886 11206
rect 17106 11134 17474 11206
rect 17694 11134 18062 11206
rect 18282 11134 18650 11206
rect 18870 11134 19238 11206
rect 19458 11134 19826 11206
rect 20046 11134 20414 11206
rect 20634 11134 21002 11206
rect 21222 11134 21590 11206
rect 21810 11134 22178 11206
rect 26502 11116 26894 11238
rect 27090 11116 27482 11238
rect 27678 11116 28070 11238
rect 28266 11116 28658 11238
rect 28854 11116 29246 11238
rect 29442 11116 29834 11238
rect 30030 11116 30422 11238
rect 30618 11116 31010 11238
rect 31206 11116 31598 11238
rect 31794 11116 32186 11238
rect 32382 11116 32774 11238
rect 32970 11116 33362 11238
rect 33558 11116 33950 11238
rect 34146 11116 34538 11238
rect 34734 11116 35126 11238
rect 35322 11116 35714 11238
rect 35910 11116 36302 11238
rect 36498 11116 36890 11238
rect 37086 11116 37478 11238
rect 37674 11116 38066 11238
rect 38262 11116 38654 11238
rect 11214 10138 11606 10276
rect 11802 10138 12194 10276
rect 12390 10138 12782 10276
rect 12978 10138 13370 10276
rect 13566 10138 13958 10276
rect 14154 10138 14546 10276
rect 14742 10138 15134 10276
rect 15330 10138 15722 10276
rect 15918 10138 16310 10276
rect 16506 10138 16898 10276
rect 17094 10138 17486 10276
rect 17682 10138 18074 10276
rect 18270 10138 18662 10276
rect 18858 10138 19250 10276
rect 19446 10138 19838 10276
rect 20034 10138 20426 10276
rect 20622 10138 21014 10276
rect 21210 10138 21602 10276
rect 21798 10138 22190 10276
rect 22974 10136 23354 10276
rect 23562 10136 23942 10276
rect 24150 10136 24530 10276
rect 24738 10136 25118 10276
rect 25326 10136 25706 10276
rect 25914 10136 26294 10276
rect 26502 10136 26882 10276
rect 27090 10136 27470 10276
rect 27678 10136 28058 10276
rect 28266 10136 28646 10276
rect 28854 10136 29234 10276
rect 29442 10136 29822 10276
rect 30030 10136 30410 10276
rect 30618 10136 30998 10276
rect 31206 10136 31586 10276
rect 31794 10136 32174 10276
rect 32382 10136 32762 10276
rect 32970 10136 33350 10276
rect 33558 10136 33938 10276
rect 34146 10136 34526 10276
rect 34734 10136 35114 10276
rect 35322 10136 35702 10276
rect 35910 10136 36290 10276
rect 36498 10136 36878 10276
rect 37086 10136 37466 10276
rect 37674 10136 38054 10276
rect 38262 10136 38642 10276
rect 10638 9118 11006 9286
rect 11226 9118 11594 9286
rect 11814 9118 12182 9286
rect 12402 9118 12770 9286
rect 12990 9118 13358 9286
rect 13578 9118 13946 9286
rect 14166 9118 14534 9286
rect 14754 9118 15122 9286
rect 15342 9118 15710 9286
rect 15930 9118 16298 9286
rect 16518 9118 16886 9286
rect 17106 9118 17474 9286
rect 17694 9118 18062 9286
rect 18282 9118 18650 9286
rect 18870 9118 19238 9286
rect 19458 9118 19826 9286
rect 20046 9118 20414 9286
rect 20634 9118 21002 9286
rect 21222 9118 21590 9286
rect 21810 9118 22178 9286
rect 22986 9116 23354 9298
rect 23574 9116 23942 9298
rect 24162 9116 24530 9298
rect 24750 9116 25118 9298
rect 25338 9116 25706 9298
rect 25926 9116 26294 9298
rect 26514 9116 26882 9298
rect 27102 9116 27470 9298
rect 27690 9116 28058 9298
rect 28278 9116 28646 9298
rect 28866 9116 29234 9298
rect 29454 9116 29822 9298
rect 30042 9116 30410 9298
rect 30630 9116 30998 9298
rect 31218 9116 31586 9298
rect 31806 9116 32174 9298
rect 32394 9116 32762 9298
rect 32982 9116 33350 9298
rect 33570 9116 33938 9298
rect 34158 9116 34526 9298
rect 34746 9116 35114 9298
rect 35334 9116 35702 9298
rect 35922 9116 36290 9298
rect 36510 9116 36878 9298
rect 37098 9116 37466 9298
rect 37686 9116 38054 9298
rect 38274 9116 38642 9298
rect 11226 8198 11594 8286
rect 11814 8198 12182 8286
rect 12402 8198 12770 8286
rect 12990 8198 13358 8286
rect 13578 8198 13946 8286
rect 14166 8198 14534 8286
rect 14754 8198 15122 8286
rect 15342 8198 15710 8286
rect 15930 8198 16298 8286
rect 16518 8198 16886 8286
rect 17106 8198 17474 8286
rect 17694 8198 18062 8286
rect 18282 8198 18650 8286
rect 18870 8198 19238 8286
rect 19458 8198 19826 8286
rect 20046 8198 20414 8286
rect 20634 8198 21002 8286
rect 21222 8198 21590 8286
rect 21810 8198 22178 8286
rect 22986 8186 23354 8284
rect 23574 8186 23942 8284
rect 24162 8186 24530 8284
rect 24750 8186 25118 8284
rect 25338 8186 25706 8284
rect 25926 8186 26294 8284
rect 26514 8186 26882 8284
rect 27102 8186 27470 8284
rect 27690 8186 28058 8284
rect 28278 8186 28646 8284
rect 28866 8186 29234 8284
rect 29454 8186 29822 8284
rect 30042 8186 30410 8284
rect 30630 8186 30998 8284
rect 31218 8186 31586 8284
rect 31806 8186 32174 8284
rect 32394 8186 32762 8284
rect 32982 8186 33350 8284
rect 33570 8186 33938 8284
rect 34158 8186 34526 8284
rect 34746 8186 35114 8284
rect 35334 8186 35702 8284
rect 35922 8186 36290 8284
rect 36510 8186 36878 8284
rect 37098 8186 37466 8284
rect 37686 8186 38054 8284
rect 38274 8186 38642 8284
<< pwell >>
rect 6619 24731 7021 29327
rect 39623 23861 40025 26857
rect 39623 20849 40025 22845
<< psubdiff >>
rect 6655 29257 6751 29291
rect 6889 29257 6985 29291
rect 6655 29195 6689 29257
rect 6951 29195 6985 29257
rect 6655 24801 6689 24863
rect 39659 26787 39755 26821
rect 39893 26787 39989 26821
rect 39659 26725 39693 26787
rect 6951 24801 6985 24863
rect 6655 24767 6751 24801
rect 6889 24767 6985 24801
rect 39955 26725 39989 26787
rect 39659 23931 39693 23993
rect 39955 23931 39989 23993
rect 39659 23897 39755 23931
rect 39893 23897 39989 23931
rect 39659 22775 39755 22809
rect 39893 22775 39989 22809
rect 39659 22713 39693 22775
rect 39955 22713 39989 22775
rect 39659 20919 39693 20981
rect 39955 20919 39989 20981
rect 39659 20885 39755 20919
rect 39893 20885 39989 20919
<< psubdiffcont >>
rect 6751 29257 6889 29291
rect 6655 24863 6689 29195
rect 6951 24863 6985 29195
rect 39755 26787 39893 26821
rect 6751 24767 6889 24801
rect 39659 23993 39693 26725
rect 39955 23993 39989 26725
rect 39755 23897 39893 23931
rect 39755 22775 39893 22809
rect 39659 20981 39693 22713
rect 39955 20981 39989 22713
rect 39755 20885 39893 20919
<< poly >>
rect 11210 27531 11610 27547
rect 11210 27497 11226 27531
rect 11594 27497 11610 27531
rect 11210 27480 11610 27497
rect 11798 27531 12198 27547
rect 11798 27497 11814 27531
rect 12182 27497 12198 27531
rect 11798 27480 12198 27497
rect 12386 27531 12786 27547
rect 12386 27497 12402 27531
rect 12770 27497 12786 27531
rect 12386 27480 12786 27497
rect 12974 27531 13374 27547
rect 12974 27497 12990 27531
rect 13358 27497 13374 27531
rect 12974 27480 13374 27497
rect 13562 27531 13962 27547
rect 13562 27497 13578 27531
rect 13946 27497 13962 27531
rect 13562 27480 13962 27497
rect 14150 27531 14550 27547
rect 14150 27497 14166 27531
rect 14534 27497 14550 27531
rect 14150 27480 14550 27497
rect 14738 27531 15138 27547
rect 14738 27497 14754 27531
rect 15122 27497 15138 27531
rect 14738 27480 15138 27497
rect 15326 27531 15726 27547
rect 15326 27497 15342 27531
rect 15710 27497 15726 27531
rect 15326 27480 15726 27497
rect 15914 27531 16314 27547
rect 15914 27497 15930 27531
rect 16298 27497 16314 27531
rect 15914 27480 16314 27497
rect 16502 27531 16902 27547
rect 16502 27497 16518 27531
rect 16886 27497 16902 27531
rect 16502 27480 16902 27497
rect 17090 27531 17490 27547
rect 17090 27497 17106 27531
rect 17474 27497 17490 27531
rect 17090 27480 17490 27497
rect 17678 27531 18078 27547
rect 17678 27497 17694 27531
rect 18062 27497 18078 27531
rect 17678 27480 18078 27497
rect 18266 27531 18666 27547
rect 18266 27497 18282 27531
rect 18650 27497 18666 27531
rect 18266 27480 18666 27497
rect 18854 27531 19254 27547
rect 18854 27497 18870 27531
rect 19238 27497 19254 27531
rect 18854 27480 19254 27497
rect 19442 27531 19842 27547
rect 19442 27497 19458 27531
rect 19826 27497 19842 27531
rect 19442 27480 19842 27497
rect 20030 27531 20430 27547
rect 20030 27497 20046 27531
rect 20414 27497 20430 27531
rect 20030 27480 20430 27497
rect 20618 27531 21018 27547
rect 20618 27497 20634 27531
rect 21002 27497 21018 27531
rect 20618 27480 21018 27497
rect 21206 27531 21606 27547
rect 21206 27497 21222 27531
rect 21590 27497 21606 27531
rect 21206 27480 21606 27497
rect 22974 27531 23366 27547
rect 22974 27497 22986 27531
rect 23354 27497 23366 27531
rect 22974 27478 23366 27497
rect 23562 27531 23954 27547
rect 23562 27497 23574 27531
rect 23942 27497 23954 27531
rect 23562 27478 23954 27497
rect 24150 27531 24542 27547
rect 24150 27497 24162 27531
rect 24530 27497 24542 27531
rect 24150 27478 24542 27497
rect 24738 27531 25130 27547
rect 24738 27497 24750 27531
rect 25118 27497 25130 27531
rect 24738 27478 25130 27497
rect 25326 27531 25718 27547
rect 25326 27497 25338 27531
rect 25706 27497 25718 27531
rect 25326 27478 25718 27497
rect 25914 27531 26306 27547
rect 25914 27497 25926 27531
rect 26294 27497 26306 27531
rect 25914 27478 26306 27497
rect 26502 27531 26894 27547
rect 26502 27497 26514 27531
rect 26882 27497 26894 27531
rect 26502 27478 26894 27497
rect 27090 27531 27482 27547
rect 27090 27497 27102 27531
rect 27470 27497 27482 27531
rect 27090 27478 27482 27497
rect 27678 27531 28070 27547
rect 27678 27497 27690 27531
rect 28058 27497 28070 27531
rect 27678 27478 28070 27497
rect 28266 27531 28658 27547
rect 28266 27497 28278 27531
rect 28646 27497 28658 27531
rect 28266 27478 28658 27497
rect 28854 27531 29246 27547
rect 28854 27497 28866 27531
rect 29234 27497 29246 27531
rect 28854 27478 29246 27497
rect 29442 27531 29834 27547
rect 29442 27497 29454 27531
rect 29822 27497 29834 27531
rect 29442 27478 29834 27497
rect 30030 27531 30422 27547
rect 30030 27497 30042 27531
rect 30410 27497 30422 27531
rect 30030 27478 30422 27497
rect 30618 27531 31010 27547
rect 30618 27497 30630 27531
rect 30998 27497 31010 27531
rect 30618 27478 31010 27497
rect 31206 27531 31598 27547
rect 31206 27497 31218 27531
rect 31586 27497 31598 27531
rect 31206 27478 31598 27497
rect 31794 27531 32186 27547
rect 31794 27497 31806 27531
rect 32174 27497 32186 27531
rect 31794 27478 32186 27497
rect 32382 27531 32774 27547
rect 32382 27497 32394 27531
rect 32762 27497 32774 27531
rect 32382 27478 32774 27497
rect 32970 27531 33362 27547
rect 32970 27497 32982 27531
rect 33350 27497 33362 27531
rect 32970 27478 33362 27497
rect 33558 27531 33950 27547
rect 33558 27497 33570 27531
rect 33938 27497 33950 27531
rect 33558 27478 33950 27497
rect 34146 27531 34538 27547
rect 34146 27497 34158 27531
rect 34526 27497 34538 27531
rect 34146 27478 34538 27497
rect 34734 27531 35126 27547
rect 34734 27497 34746 27531
rect 35114 27497 35126 27531
rect 34734 27478 35126 27497
rect 35322 27531 35714 27547
rect 35322 27497 35334 27531
rect 35702 27497 35714 27531
rect 35322 27478 35714 27497
rect 35910 27531 36302 27547
rect 35910 27497 35922 27531
rect 36290 27497 36302 27531
rect 35910 27478 36302 27497
rect 36498 27531 36890 27547
rect 36498 27497 36510 27531
rect 36878 27497 36890 27531
rect 36498 27478 36890 27497
rect 37086 27531 37478 27547
rect 37086 27497 37098 27531
rect 37466 27497 37478 27531
rect 37086 27478 37478 27497
rect 37674 27531 38066 27547
rect 37674 27497 37686 27531
rect 38054 27497 38066 27531
rect 37674 27478 38066 27497
rect 38262 27531 38654 27547
rect 38262 27497 38274 27531
rect 38642 27497 38654 27531
rect 38262 27478 38654 27497
rect 11214 26603 11606 26614
rect 11214 26569 11226 26603
rect 11594 26569 11606 26603
rect 11214 26531 11606 26569
rect 11214 26497 11226 26531
rect 11594 26497 11606 26531
rect 11214 26480 11606 26497
rect 11802 26603 12194 26614
rect 11802 26569 11814 26603
rect 12182 26569 12194 26603
rect 11802 26531 12194 26569
rect 11802 26497 11814 26531
rect 12182 26497 12194 26531
rect 11802 26480 12194 26497
rect 12390 26603 12782 26614
rect 12390 26569 12402 26603
rect 12770 26569 12782 26603
rect 12390 26531 12782 26569
rect 12390 26497 12402 26531
rect 12770 26497 12782 26531
rect 12390 26480 12782 26497
rect 12978 26603 13370 26614
rect 12978 26569 12990 26603
rect 13358 26569 13370 26603
rect 12978 26531 13370 26569
rect 12978 26497 12990 26531
rect 13358 26497 13370 26531
rect 12978 26480 13370 26497
rect 13566 26603 13958 26614
rect 13566 26569 13578 26603
rect 13946 26569 13958 26603
rect 13566 26531 13958 26569
rect 13566 26497 13578 26531
rect 13946 26497 13958 26531
rect 13566 26480 13958 26497
rect 14154 26603 14546 26614
rect 14154 26569 14166 26603
rect 14534 26569 14546 26603
rect 14154 26531 14546 26569
rect 14154 26497 14166 26531
rect 14534 26497 14546 26531
rect 14154 26480 14546 26497
rect 14742 26603 15134 26614
rect 14742 26569 14754 26603
rect 15122 26569 15134 26603
rect 14742 26531 15134 26569
rect 14742 26497 14754 26531
rect 15122 26497 15134 26531
rect 14742 26480 15134 26497
rect 15330 26603 15722 26614
rect 15330 26569 15342 26603
rect 15710 26569 15722 26603
rect 15330 26531 15722 26569
rect 15330 26497 15342 26531
rect 15710 26497 15722 26531
rect 15330 26480 15722 26497
rect 15918 26603 16310 26614
rect 15918 26569 15930 26603
rect 16298 26569 16310 26603
rect 15918 26531 16310 26569
rect 15918 26497 15930 26531
rect 16298 26497 16310 26531
rect 15918 26480 16310 26497
rect 16506 26603 16898 26614
rect 16506 26569 16518 26603
rect 16886 26569 16898 26603
rect 16506 26531 16898 26569
rect 16506 26497 16518 26531
rect 16886 26497 16898 26531
rect 16506 26480 16898 26497
rect 17094 26603 17486 26614
rect 17094 26569 17106 26603
rect 17474 26569 17486 26603
rect 17094 26531 17486 26569
rect 17094 26497 17106 26531
rect 17474 26497 17486 26531
rect 17094 26480 17486 26497
rect 17682 26603 18074 26614
rect 17682 26569 17694 26603
rect 18062 26569 18074 26603
rect 17682 26531 18074 26569
rect 17682 26497 17694 26531
rect 18062 26497 18074 26531
rect 17682 26480 18074 26497
rect 18270 26603 18662 26614
rect 18270 26569 18282 26603
rect 18650 26569 18662 26603
rect 18270 26531 18662 26569
rect 18270 26497 18282 26531
rect 18650 26497 18662 26531
rect 18270 26480 18662 26497
rect 18858 26603 19250 26614
rect 18858 26569 18870 26603
rect 19238 26569 19250 26603
rect 18858 26531 19250 26569
rect 18858 26497 18870 26531
rect 19238 26497 19250 26531
rect 18858 26480 19250 26497
rect 19446 26603 19838 26614
rect 19446 26569 19458 26603
rect 19826 26569 19838 26603
rect 19446 26531 19838 26569
rect 19446 26497 19458 26531
rect 19826 26497 19838 26531
rect 19446 26480 19838 26497
rect 20034 26603 20426 26614
rect 20034 26569 20046 26603
rect 20414 26569 20426 26603
rect 20034 26531 20426 26569
rect 20034 26497 20046 26531
rect 20414 26497 20426 26531
rect 20034 26480 20426 26497
rect 20622 26603 21014 26614
rect 20622 26569 20634 26603
rect 21002 26569 21014 26603
rect 20622 26531 21014 26569
rect 20622 26497 20634 26531
rect 21002 26497 21014 26531
rect 20622 26480 21014 26497
rect 21210 26603 21602 26614
rect 21210 26569 21222 26603
rect 21590 26569 21602 26603
rect 21210 26531 21602 26569
rect 21210 26497 21222 26531
rect 21590 26497 21602 26531
rect 21210 26480 21602 26497
rect 21798 26603 22190 26614
rect 21798 26569 21810 26603
rect 22178 26569 22190 26603
rect 21798 26531 22190 26569
rect 21798 26497 21810 26531
rect 22178 26497 22190 26531
rect 21798 26480 22190 26497
rect 22974 26603 23354 26614
rect 22974 26569 22986 26603
rect 22974 26531 23354 26569
rect 22974 26497 22986 26531
rect 22974 26486 23354 26497
rect 23562 26603 23942 26614
rect 23562 26569 23574 26603
rect 23562 26531 23942 26569
rect 23562 26497 23574 26531
rect 23562 26486 23942 26497
rect 24150 26603 24530 26614
rect 24150 26569 24162 26603
rect 24150 26531 24530 26569
rect 24150 26497 24162 26531
rect 24150 26486 24530 26497
rect 24738 26603 25118 26614
rect 24738 26569 24750 26603
rect 24738 26531 25118 26569
rect 24738 26497 24750 26531
rect 24738 26486 25118 26497
rect 25326 26603 25706 26614
rect 25326 26569 25338 26603
rect 25326 26531 25706 26569
rect 25326 26497 25338 26531
rect 25326 26486 25706 26497
rect 25914 26603 26294 26614
rect 25914 26569 25926 26603
rect 25914 26531 26294 26569
rect 25914 26497 25926 26531
rect 25914 26486 26294 26497
rect 26502 26603 26882 26614
rect 26502 26569 26514 26603
rect 26502 26531 26882 26569
rect 26502 26497 26514 26531
rect 26502 26486 26882 26497
rect 27090 26603 27470 26614
rect 27090 26569 27102 26603
rect 27090 26531 27470 26569
rect 27090 26497 27102 26531
rect 27090 26486 27470 26497
rect 27678 26603 28058 26614
rect 27678 26569 27690 26603
rect 27678 26531 28058 26569
rect 27678 26497 27690 26531
rect 27678 26486 28058 26497
rect 28266 26603 28646 26614
rect 28266 26569 28278 26603
rect 28266 26531 28646 26569
rect 28266 26497 28278 26531
rect 28266 26486 28646 26497
rect 28854 26603 29234 26614
rect 28854 26569 28866 26603
rect 28854 26531 29234 26569
rect 28854 26497 28866 26531
rect 28854 26486 29234 26497
rect 29442 26603 29822 26614
rect 29442 26569 29454 26603
rect 29442 26531 29822 26569
rect 29442 26497 29454 26531
rect 29442 26486 29822 26497
rect 30030 26603 30410 26614
rect 30030 26569 30042 26603
rect 30030 26531 30410 26569
rect 30030 26497 30042 26531
rect 30030 26486 30410 26497
rect 30618 26603 30998 26614
rect 30618 26569 30630 26603
rect 30618 26531 30998 26569
rect 30618 26497 30630 26531
rect 30618 26486 30998 26497
rect 31206 26603 31586 26614
rect 31206 26569 31218 26603
rect 31206 26531 31586 26569
rect 31206 26497 31218 26531
rect 31206 26486 31586 26497
rect 31794 26603 32174 26614
rect 31794 26569 31806 26603
rect 31794 26531 32174 26569
rect 31794 26497 31806 26531
rect 31794 26486 32174 26497
rect 32382 26603 32762 26614
rect 32382 26569 32394 26603
rect 32382 26531 32762 26569
rect 32382 26497 32394 26531
rect 32382 26486 32762 26497
rect 32970 26603 33350 26614
rect 32970 26569 32982 26603
rect 32970 26531 33350 26569
rect 32970 26497 32982 26531
rect 32970 26486 33350 26497
rect 33558 26603 33938 26614
rect 33558 26569 33570 26603
rect 33558 26531 33938 26569
rect 33558 26497 33570 26531
rect 33558 26486 33938 26497
rect 34146 26603 34526 26614
rect 34146 26569 34158 26603
rect 34146 26531 34526 26569
rect 34146 26497 34158 26531
rect 34146 26486 34526 26497
rect 34734 26603 35114 26614
rect 34734 26569 34746 26603
rect 34734 26531 35114 26569
rect 34734 26497 34746 26531
rect 34734 26486 35114 26497
rect 35322 26603 35702 26614
rect 35322 26569 35334 26603
rect 35322 26531 35702 26569
rect 35322 26497 35334 26531
rect 35322 26486 35702 26497
rect 35910 26603 36290 26614
rect 35910 26569 35922 26603
rect 35910 26531 36290 26569
rect 35910 26497 35922 26531
rect 35910 26486 36290 26497
rect 36498 26603 36878 26614
rect 36498 26569 36510 26603
rect 36498 26531 36878 26569
rect 36498 26497 36510 26531
rect 36498 26486 36878 26497
rect 37086 26603 37466 26614
rect 37086 26569 37098 26603
rect 37086 26531 37466 26569
rect 37086 26497 37098 26531
rect 37086 26486 37466 26497
rect 37674 26603 38054 26614
rect 37674 26569 37686 26603
rect 37674 26531 38054 26569
rect 37674 26497 37686 26531
rect 37674 26486 38054 26497
rect 38262 26603 38642 26614
rect 38262 26569 38274 26603
rect 38262 26531 38642 26569
rect 38262 26497 38274 26531
rect 38262 26486 38642 26497
rect 10638 25603 11006 25614
rect 10638 25531 11006 25569
rect 10638 25486 11006 25497
rect 11226 25603 11594 25614
rect 11226 25531 11594 25569
rect 11226 25486 11594 25497
rect 11814 25603 12182 25614
rect 11814 25531 12182 25569
rect 11814 25486 12182 25497
rect 12402 25603 12770 25614
rect 12402 25531 12770 25569
rect 12402 25486 12770 25497
rect 12990 25603 13358 25614
rect 12990 25531 13358 25569
rect 12990 25486 13358 25497
rect 13578 25603 13946 25614
rect 13578 25531 13946 25569
rect 13578 25486 13946 25497
rect 14166 25603 14534 25614
rect 14166 25531 14534 25569
rect 14166 25486 14534 25497
rect 14754 25603 15122 25614
rect 14754 25531 15122 25569
rect 14754 25486 15122 25497
rect 15342 25603 15710 25614
rect 15342 25531 15710 25569
rect 15342 25486 15710 25497
rect 15930 25603 16298 25614
rect 15930 25531 16298 25569
rect 15930 25486 16298 25497
rect 16518 25603 16886 25614
rect 16518 25531 16886 25569
rect 16518 25486 16886 25497
rect 17106 25603 17474 25614
rect 17106 25531 17474 25569
rect 17106 25486 17474 25497
rect 17694 25603 18062 25614
rect 17694 25531 18062 25569
rect 17694 25486 18062 25497
rect 18282 25603 18650 25614
rect 18282 25531 18650 25569
rect 18282 25486 18650 25497
rect 18870 25603 19238 25614
rect 18870 25531 19238 25569
rect 18870 25486 19238 25497
rect 19458 25603 19826 25614
rect 19458 25531 19826 25569
rect 19458 25486 19826 25497
rect 20046 25603 20414 25614
rect 20046 25531 20414 25569
rect 20046 25486 20414 25497
rect 20634 25603 21002 25614
rect 20634 25531 21002 25569
rect 20634 25486 21002 25497
rect 21222 25603 21590 25614
rect 21222 25531 21590 25569
rect 21222 25486 21590 25497
rect 21810 25603 22178 25614
rect 21810 25531 22178 25569
rect 21810 25486 22178 25497
rect 23574 25603 23942 25616
rect 23574 25531 23942 25569
rect 23574 25484 23942 25497
rect 24162 25603 24530 25616
rect 24162 25531 24530 25569
rect 24162 25484 24530 25497
rect 24750 25603 25118 25616
rect 24750 25531 25118 25569
rect 24750 25484 25118 25497
rect 25338 25603 25706 25616
rect 25338 25531 25706 25569
rect 25338 25484 25706 25497
rect 25926 25603 26294 25616
rect 25926 25531 26294 25569
rect 25926 25484 26294 25497
rect 26514 25603 26882 25616
rect 26514 25531 26882 25569
rect 26514 25484 26882 25497
rect 27102 25603 27470 25616
rect 27102 25531 27470 25569
rect 27102 25484 27470 25497
rect 27690 25603 28058 25616
rect 27690 25531 28058 25569
rect 27690 25484 28058 25497
rect 28278 25603 28646 25616
rect 28278 25531 28646 25569
rect 28278 25484 28646 25497
rect 28866 25603 29234 25616
rect 28866 25531 29234 25569
rect 28866 25484 29234 25497
rect 29454 25603 29822 25616
rect 29454 25531 29822 25569
rect 29454 25484 29822 25497
rect 30042 25603 30410 25616
rect 30042 25531 30410 25569
rect 30042 25484 30410 25497
rect 30630 25603 30998 25616
rect 30630 25531 30998 25569
rect 30630 25484 30998 25497
rect 31218 25603 31586 25616
rect 31218 25531 31586 25569
rect 31218 25484 31586 25497
rect 31806 25603 32174 25616
rect 31806 25531 32174 25569
rect 31806 25484 32174 25497
rect 32394 25603 32762 25616
rect 32394 25531 32762 25569
rect 32394 25484 32762 25497
rect 32982 25603 33350 25616
rect 32982 25531 33350 25569
rect 32982 25484 33350 25497
rect 33570 25603 33938 25616
rect 33570 25531 33938 25569
rect 33570 25484 33938 25497
rect 34158 25603 34526 25616
rect 34158 25531 34526 25569
rect 34158 25484 34526 25497
rect 34746 25603 35114 25616
rect 34746 25531 35114 25569
rect 34746 25484 35114 25497
rect 35334 25603 35702 25616
rect 35334 25531 35702 25569
rect 35334 25484 35702 25497
rect 35922 25603 36290 25616
rect 35922 25531 36290 25569
rect 35922 25484 36290 25497
rect 36510 25603 36878 25616
rect 36510 25531 36878 25569
rect 36510 25484 36878 25497
rect 37098 25603 37466 25616
rect 37098 25531 37466 25569
rect 37098 25484 37466 25497
rect 37686 25603 38054 25616
rect 37686 25531 38054 25569
rect 37686 25484 38054 25497
rect 38274 25603 38642 25616
rect 38274 25531 38642 25569
rect 38274 25484 38642 25497
rect 11210 24603 11594 24622
rect 11210 24569 11226 24603
rect 11210 24553 11594 24569
rect 11798 24603 12182 24622
rect 11798 24569 11814 24603
rect 11798 24553 12182 24569
rect 12386 24603 12770 24622
rect 12386 24569 12402 24603
rect 12386 24553 12770 24569
rect 12974 24603 13358 24622
rect 12974 24569 12990 24603
rect 12974 24553 13358 24569
rect 13562 24603 13946 24622
rect 13562 24569 13578 24603
rect 13562 24553 13946 24569
rect 14150 24603 14534 24622
rect 14150 24569 14166 24603
rect 14150 24553 14534 24569
rect 14738 24603 15122 24622
rect 14738 24569 14754 24603
rect 14738 24553 15122 24569
rect 15326 24603 15710 24622
rect 15326 24569 15342 24603
rect 15326 24553 15710 24569
rect 15914 24603 16298 24622
rect 15914 24569 15930 24603
rect 15914 24553 16298 24569
rect 16502 24603 16886 24622
rect 16502 24569 16518 24603
rect 16502 24553 16886 24569
rect 17090 24603 17474 24622
rect 17090 24569 17106 24603
rect 17090 24553 17474 24569
rect 17678 24603 18062 24622
rect 17678 24569 17694 24603
rect 17678 24553 18062 24569
rect 18266 24603 18650 24622
rect 18266 24569 18282 24603
rect 18266 24553 18650 24569
rect 18854 24603 19238 24622
rect 18854 24569 18870 24603
rect 18854 24553 19238 24569
rect 19442 24603 19826 24622
rect 19442 24569 19458 24603
rect 19442 24553 19826 24569
rect 20030 24603 20414 24622
rect 20030 24569 20046 24603
rect 20030 24553 20414 24569
rect 20618 24603 21002 24622
rect 20618 24569 20634 24603
rect 20618 24553 21002 24569
rect 21206 24603 21590 24622
rect 21206 24569 21222 24603
rect 21206 24553 21590 24569
rect 21794 24603 22178 24622
rect 21794 24569 21810 24603
rect 21794 24553 22178 24569
rect 22986 24603 23354 24632
rect 22986 24553 23354 24569
rect 23574 24603 23942 24632
rect 23574 24553 23942 24569
rect 24162 24603 24530 24632
rect 24162 24553 24530 24569
rect 24750 24603 25118 24632
rect 24750 24553 25118 24569
rect 25338 24603 25706 24632
rect 25338 24553 25706 24569
rect 25926 24603 26294 24632
rect 25926 24553 26294 24569
rect 26514 24603 26882 24632
rect 26514 24553 26882 24569
rect 27102 24603 27470 24632
rect 27102 24553 27470 24569
rect 27690 24603 28058 24632
rect 27690 24553 28058 24569
rect 28278 24603 28646 24632
rect 28278 24553 28646 24569
rect 28866 24603 29234 24632
rect 28866 24553 29234 24569
rect 29454 24603 29822 24632
rect 29454 24553 29822 24569
rect 30042 24603 30410 24632
rect 30042 24553 30410 24569
rect 30630 24603 30998 24632
rect 30630 24553 30998 24569
rect 31218 24603 31586 24632
rect 31218 24553 31586 24569
rect 31806 24603 32174 24632
rect 31806 24553 32174 24569
rect 32394 24603 32762 24632
rect 32394 24553 32762 24569
rect 32982 24603 33350 24632
rect 32982 24553 33350 24569
rect 33570 24603 33938 24632
rect 33570 24553 33938 24569
rect 34158 24603 34526 24632
rect 34158 24553 34526 24569
rect 34746 24603 35114 24632
rect 34746 24553 35114 24569
rect 35334 24603 35702 24632
rect 35334 24553 35702 24569
rect 35922 24603 36290 24632
rect 35922 24553 36290 24569
rect 36510 24603 36878 24632
rect 36510 24553 36878 24569
rect 37098 24603 37466 24632
rect 37098 24553 37466 24569
rect 37686 24603 38054 24632
rect 37686 24553 38054 24569
rect 38274 24603 38642 24632
rect 38274 24553 38642 24569
rect 11226 11187 11594 11203
rect 11226 11134 11594 11153
rect 11814 11187 12182 11203
rect 11814 11134 12182 11153
rect 12402 11187 12770 11203
rect 12402 11134 12770 11153
rect 12990 11187 13358 11203
rect 12990 11134 13358 11153
rect 13578 11187 13946 11203
rect 13578 11134 13946 11153
rect 14166 11187 14534 11203
rect 14166 11134 14534 11153
rect 14754 11187 15122 11203
rect 14754 11134 15122 11153
rect 15342 11187 15710 11203
rect 15342 11134 15710 11153
rect 15930 11187 16298 11203
rect 15930 11134 16298 11153
rect 16518 11187 16886 11203
rect 16518 11134 16886 11153
rect 17106 11187 17474 11203
rect 17106 11134 17474 11153
rect 17694 11187 18062 11203
rect 17694 11134 18062 11153
rect 18282 11187 18650 11203
rect 18282 11134 18650 11153
rect 18870 11187 19238 11203
rect 18870 11134 19238 11153
rect 19458 11187 19826 11203
rect 19458 11134 19826 11153
rect 20046 11187 20414 11203
rect 20046 11134 20414 11153
rect 20634 11187 21002 11203
rect 20634 11134 21002 11153
rect 21222 11187 21590 11203
rect 21222 11134 21590 11153
rect 21810 11187 22178 11203
rect 21810 11134 22178 11153
rect 26502 11187 26894 11203
rect 26502 11153 26514 11187
rect 26882 11153 26894 11187
rect 26502 11116 26894 11153
rect 27090 11187 27482 11203
rect 27090 11153 27102 11187
rect 27470 11153 27482 11187
rect 27090 11116 27482 11153
rect 27678 11187 28070 11203
rect 27678 11153 27690 11187
rect 28058 11153 28070 11187
rect 27678 11116 28070 11153
rect 28266 11187 28658 11203
rect 28266 11153 28278 11187
rect 28646 11153 28658 11187
rect 28266 11116 28658 11153
rect 28854 11187 29246 11203
rect 28854 11153 28866 11187
rect 29234 11153 29246 11187
rect 28854 11116 29246 11153
rect 29442 11187 29834 11203
rect 29442 11153 29454 11187
rect 29822 11153 29834 11187
rect 29442 11116 29834 11153
rect 30030 11187 30422 11203
rect 30030 11153 30042 11187
rect 30410 11153 30422 11187
rect 30030 11116 30422 11153
rect 30618 11187 31010 11203
rect 30618 11153 30630 11187
rect 30998 11153 31010 11187
rect 30618 11116 31010 11153
rect 31206 11187 31598 11203
rect 31206 11153 31218 11187
rect 31586 11153 31598 11187
rect 31206 11116 31598 11153
rect 31794 11187 32186 11203
rect 31794 11153 31806 11187
rect 32174 11153 32186 11187
rect 31794 11116 32186 11153
rect 32382 11187 32774 11203
rect 32382 11153 32394 11187
rect 32762 11153 32774 11187
rect 32382 11116 32774 11153
rect 32970 11187 33362 11203
rect 32970 11153 32982 11187
rect 33350 11153 33362 11187
rect 32970 11116 33362 11153
rect 33558 11187 33950 11203
rect 33558 11153 33570 11187
rect 33938 11153 33950 11187
rect 33558 11116 33950 11153
rect 34146 11187 34538 11203
rect 34146 11153 34158 11187
rect 34526 11153 34538 11187
rect 34146 11116 34538 11153
rect 34734 11187 35126 11203
rect 34734 11153 34746 11187
rect 35114 11153 35126 11187
rect 34734 11116 35126 11153
rect 35322 11187 35714 11203
rect 35322 11153 35334 11187
rect 35702 11153 35714 11187
rect 35322 11116 35714 11153
rect 35910 11187 36302 11203
rect 35910 11153 35922 11187
rect 36290 11153 36302 11187
rect 35910 11116 36302 11153
rect 36498 11187 36890 11203
rect 36498 11153 36510 11187
rect 36878 11153 36890 11187
rect 36498 11116 36890 11153
rect 37086 11187 37478 11203
rect 37086 11153 37098 11187
rect 37466 11153 37478 11187
rect 37086 11116 37478 11153
rect 37674 11187 38066 11203
rect 37674 11153 37686 11187
rect 38054 11153 38066 11187
rect 37674 11116 38066 11153
rect 38262 11187 38654 11203
rect 38262 11153 38274 11187
rect 38642 11153 38654 11187
rect 38262 11116 38654 11153
rect 11214 10259 11606 10276
rect 11214 10225 11226 10259
rect 11594 10225 11606 10259
rect 11214 10187 11606 10225
rect 11214 10153 11226 10187
rect 11594 10153 11606 10187
rect 11214 10138 11606 10153
rect 11802 10259 12194 10276
rect 11802 10225 11814 10259
rect 12182 10225 12194 10259
rect 11802 10187 12194 10225
rect 11802 10153 11814 10187
rect 12182 10153 12194 10187
rect 11802 10138 12194 10153
rect 12390 10259 12782 10276
rect 12390 10225 12402 10259
rect 12770 10225 12782 10259
rect 12390 10187 12782 10225
rect 12390 10153 12402 10187
rect 12770 10153 12782 10187
rect 12390 10138 12782 10153
rect 12978 10259 13370 10276
rect 12978 10225 12990 10259
rect 13358 10225 13370 10259
rect 12978 10187 13370 10225
rect 12978 10153 12990 10187
rect 13358 10153 13370 10187
rect 12978 10138 13370 10153
rect 13566 10259 13958 10276
rect 13566 10225 13578 10259
rect 13946 10225 13958 10259
rect 13566 10187 13958 10225
rect 13566 10153 13578 10187
rect 13946 10153 13958 10187
rect 13566 10138 13958 10153
rect 14154 10259 14546 10276
rect 14154 10225 14166 10259
rect 14534 10225 14546 10259
rect 14154 10187 14546 10225
rect 14154 10153 14166 10187
rect 14534 10153 14546 10187
rect 14154 10138 14546 10153
rect 14742 10259 15134 10276
rect 14742 10225 14754 10259
rect 15122 10225 15134 10259
rect 14742 10187 15134 10225
rect 14742 10153 14754 10187
rect 15122 10153 15134 10187
rect 14742 10138 15134 10153
rect 15330 10259 15722 10276
rect 15330 10225 15342 10259
rect 15710 10225 15722 10259
rect 15330 10187 15722 10225
rect 15330 10153 15342 10187
rect 15710 10153 15722 10187
rect 15330 10138 15722 10153
rect 15918 10259 16310 10276
rect 15918 10225 15930 10259
rect 16298 10225 16310 10259
rect 15918 10187 16310 10225
rect 15918 10153 15930 10187
rect 16298 10153 16310 10187
rect 15918 10138 16310 10153
rect 16506 10259 16898 10276
rect 16506 10225 16518 10259
rect 16886 10225 16898 10259
rect 16506 10187 16898 10225
rect 16506 10153 16518 10187
rect 16886 10153 16898 10187
rect 16506 10138 16898 10153
rect 17094 10259 17486 10276
rect 17094 10225 17106 10259
rect 17474 10225 17486 10259
rect 17094 10187 17486 10225
rect 17094 10153 17106 10187
rect 17474 10153 17486 10187
rect 17094 10138 17486 10153
rect 17682 10259 18074 10276
rect 17682 10225 17694 10259
rect 18062 10225 18074 10259
rect 17682 10187 18074 10225
rect 17682 10153 17694 10187
rect 18062 10153 18074 10187
rect 17682 10138 18074 10153
rect 18270 10259 18662 10276
rect 18270 10225 18282 10259
rect 18650 10225 18662 10259
rect 18270 10187 18662 10225
rect 18270 10153 18282 10187
rect 18650 10153 18662 10187
rect 18270 10138 18662 10153
rect 18858 10259 19250 10276
rect 18858 10225 18870 10259
rect 19238 10225 19250 10259
rect 18858 10187 19250 10225
rect 18858 10153 18870 10187
rect 19238 10153 19250 10187
rect 18858 10138 19250 10153
rect 19446 10259 19838 10276
rect 19446 10225 19458 10259
rect 19826 10225 19838 10259
rect 19446 10187 19838 10225
rect 19446 10153 19458 10187
rect 19826 10153 19838 10187
rect 19446 10138 19838 10153
rect 20034 10259 20426 10276
rect 20034 10225 20046 10259
rect 20414 10225 20426 10259
rect 20034 10187 20426 10225
rect 20034 10153 20046 10187
rect 20414 10153 20426 10187
rect 20034 10138 20426 10153
rect 20622 10259 21014 10276
rect 20622 10225 20634 10259
rect 21002 10225 21014 10259
rect 20622 10187 21014 10225
rect 20622 10153 20634 10187
rect 21002 10153 21014 10187
rect 20622 10138 21014 10153
rect 21210 10259 21602 10276
rect 21210 10225 21222 10259
rect 21590 10225 21602 10259
rect 21210 10187 21602 10225
rect 21210 10153 21222 10187
rect 21590 10153 21602 10187
rect 21210 10138 21602 10153
rect 21798 10259 22190 10276
rect 21798 10225 21810 10259
rect 22178 10225 22190 10259
rect 21798 10187 22190 10225
rect 21798 10153 21810 10187
rect 22178 10153 22190 10187
rect 21798 10138 22190 10153
rect 22974 10259 23354 10276
rect 22974 10225 22986 10259
rect 22974 10187 23354 10225
rect 22974 10153 22986 10187
rect 22974 10136 23354 10153
rect 23562 10259 23942 10276
rect 23562 10225 23574 10259
rect 23562 10187 23942 10225
rect 23562 10153 23574 10187
rect 23562 10136 23942 10153
rect 24150 10259 24530 10276
rect 24150 10225 24162 10259
rect 24150 10187 24530 10225
rect 24150 10153 24162 10187
rect 24150 10136 24530 10153
rect 24738 10259 25118 10276
rect 24738 10225 24750 10259
rect 24738 10187 25118 10225
rect 24738 10153 24750 10187
rect 24738 10136 25118 10153
rect 25326 10259 25706 10276
rect 25326 10225 25338 10259
rect 25326 10187 25706 10225
rect 25326 10153 25338 10187
rect 25326 10136 25706 10153
rect 25914 10259 26294 10276
rect 25914 10225 25926 10259
rect 25914 10187 26294 10225
rect 25914 10153 25926 10187
rect 25914 10136 26294 10153
rect 26502 10259 26882 10276
rect 26502 10225 26514 10259
rect 26502 10187 26882 10225
rect 26502 10153 26514 10187
rect 26502 10136 26882 10153
rect 27090 10259 27470 10276
rect 27090 10225 27102 10259
rect 27090 10187 27470 10225
rect 27090 10153 27102 10187
rect 27090 10136 27470 10153
rect 27678 10259 28058 10276
rect 27678 10225 27690 10259
rect 27678 10187 28058 10225
rect 27678 10153 27690 10187
rect 27678 10136 28058 10153
rect 28266 10259 28646 10276
rect 28266 10225 28278 10259
rect 28266 10187 28646 10225
rect 28266 10153 28278 10187
rect 28266 10136 28646 10153
rect 28854 10259 29234 10276
rect 28854 10225 28866 10259
rect 28854 10187 29234 10225
rect 28854 10153 28866 10187
rect 28854 10136 29234 10153
rect 29442 10259 29822 10276
rect 29442 10225 29454 10259
rect 29442 10187 29822 10225
rect 29442 10153 29454 10187
rect 29442 10136 29822 10153
rect 30030 10259 30410 10276
rect 30030 10225 30042 10259
rect 30030 10187 30410 10225
rect 30030 10153 30042 10187
rect 30030 10136 30410 10153
rect 30618 10259 30998 10276
rect 30618 10225 30630 10259
rect 30618 10187 30998 10225
rect 30618 10153 30630 10187
rect 30618 10136 30998 10153
rect 31206 10259 31586 10276
rect 31206 10225 31218 10259
rect 31206 10187 31586 10225
rect 31206 10153 31218 10187
rect 31206 10136 31586 10153
rect 31794 10259 32174 10276
rect 31794 10225 31806 10259
rect 31794 10187 32174 10225
rect 31794 10153 31806 10187
rect 31794 10136 32174 10153
rect 32382 10259 32762 10276
rect 32382 10225 32394 10259
rect 32382 10187 32762 10225
rect 32382 10153 32394 10187
rect 32382 10136 32762 10153
rect 32970 10259 33350 10276
rect 32970 10225 32982 10259
rect 32970 10187 33350 10225
rect 32970 10153 32982 10187
rect 32970 10136 33350 10153
rect 33558 10259 33938 10276
rect 33558 10225 33570 10259
rect 33558 10187 33938 10225
rect 33558 10153 33570 10187
rect 33558 10136 33938 10153
rect 34146 10259 34526 10276
rect 34146 10225 34158 10259
rect 34146 10187 34526 10225
rect 34146 10153 34158 10187
rect 34146 10136 34526 10153
rect 34734 10259 35114 10276
rect 34734 10225 34746 10259
rect 34734 10187 35114 10225
rect 34734 10153 34746 10187
rect 34734 10136 35114 10153
rect 35322 10259 35702 10276
rect 35322 10225 35334 10259
rect 35322 10187 35702 10225
rect 35322 10153 35334 10187
rect 35322 10136 35702 10153
rect 35910 10259 36290 10276
rect 35910 10225 35922 10259
rect 35910 10187 36290 10225
rect 35910 10153 35922 10187
rect 35910 10136 36290 10153
rect 36498 10259 36878 10276
rect 36498 10225 36510 10259
rect 36498 10187 36878 10225
rect 36498 10153 36510 10187
rect 36498 10136 36878 10153
rect 37086 10259 37466 10276
rect 37086 10225 37098 10259
rect 37086 10187 37466 10225
rect 37086 10153 37098 10187
rect 37086 10136 37466 10153
rect 37674 10259 38054 10276
rect 37674 10225 37686 10259
rect 37674 10187 38054 10225
rect 37674 10153 37686 10187
rect 37674 10136 38054 10153
rect 38262 10259 38642 10276
rect 38262 10225 38274 10259
rect 38262 10187 38642 10225
rect 38262 10153 38274 10187
rect 38262 10136 38642 10153
rect 10638 9259 11006 9286
rect 10638 9187 11006 9225
rect 10638 9118 11006 9153
rect 11226 9259 11594 9286
rect 11226 9187 11594 9225
rect 11226 9118 11594 9153
rect 11814 9259 12182 9286
rect 11814 9187 12182 9225
rect 11814 9118 12182 9153
rect 12402 9259 12770 9286
rect 12402 9187 12770 9225
rect 12402 9118 12770 9153
rect 12990 9259 13358 9286
rect 12990 9187 13358 9225
rect 12990 9118 13358 9153
rect 13578 9259 13946 9286
rect 13578 9187 13946 9225
rect 13578 9118 13946 9153
rect 14166 9259 14534 9286
rect 14166 9187 14534 9225
rect 14166 9118 14534 9153
rect 14754 9259 15122 9286
rect 14754 9187 15122 9225
rect 14754 9118 15122 9153
rect 15342 9259 15710 9286
rect 15342 9187 15710 9225
rect 15342 9118 15710 9153
rect 15930 9259 16298 9286
rect 15930 9187 16298 9225
rect 15930 9118 16298 9153
rect 16518 9259 16886 9286
rect 16518 9187 16886 9225
rect 16518 9118 16886 9153
rect 17106 9259 17474 9286
rect 17106 9187 17474 9225
rect 17106 9118 17474 9153
rect 17694 9259 18062 9286
rect 17694 9187 18062 9225
rect 17694 9118 18062 9153
rect 18282 9259 18650 9286
rect 18282 9187 18650 9225
rect 18282 9118 18650 9153
rect 18870 9259 19238 9286
rect 18870 9187 19238 9225
rect 18870 9118 19238 9153
rect 19458 9259 19826 9286
rect 19458 9187 19826 9225
rect 19458 9118 19826 9153
rect 20046 9259 20414 9286
rect 20046 9187 20414 9225
rect 20046 9118 20414 9153
rect 20634 9259 21002 9286
rect 20634 9187 21002 9225
rect 20634 9118 21002 9153
rect 21222 9259 21590 9286
rect 21222 9187 21590 9225
rect 21222 9118 21590 9153
rect 21810 9259 22178 9286
rect 21810 9187 22178 9225
rect 21810 9118 22178 9153
rect 22986 9259 23354 9298
rect 22986 9187 23354 9225
rect 22986 9116 23354 9153
rect 23574 9259 23942 9298
rect 23574 9187 23942 9225
rect 23574 9116 23942 9153
rect 24162 9259 24530 9298
rect 24162 9187 24530 9225
rect 24162 9116 24530 9153
rect 24750 9259 25118 9298
rect 24750 9187 25118 9225
rect 24750 9116 25118 9153
rect 25338 9259 25706 9298
rect 25338 9187 25706 9225
rect 25338 9116 25706 9153
rect 25926 9259 26294 9298
rect 25926 9187 26294 9225
rect 25926 9116 26294 9153
rect 26514 9259 26882 9298
rect 26514 9187 26882 9225
rect 26514 9116 26882 9153
rect 27102 9259 27470 9298
rect 27102 9187 27470 9225
rect 27102 9116 27470 9153
rect 27690 9259 28058 9298
rect 27690 9187 28058 9225
rect 27690 9116 28058 9153
rect 28278 9259 28646 9298
rect 28278 9187 28646 9225
rect 28278 9116 28646 9153
rect 28866 9259 29234 9298
rect 28866 9187 29234 9225
rect 28866 9116 29234 9153
rect 29454 9259 29822 9298
rect 29454 9187 29822 9225
rect 29454 9116 29822 9153
rect 30042 9259 30410 9298
rect 30042 9187 30410 9225
rect 30042 9116 30410 9153
rect 30630 9259 30998 9298
rect 30630 9187 30998 9225
rect 30630 9116 30998 9153
rect 31218 9259 31586 9298
rect 31218 9187 31586 9225
rect 31218 9116 31586 9153
rect 31806 9259 32174 9298
rect 31806 9187 32174 9225
rect 31806 9116 32174 9153
rect 32394 9259 32762 9298
rect 32394 9187 32762 9225
rect 32394 9116 32762 9153
rect 32982 9259 33350 9298
rect 32982 9187 33350 9225
rect 32982 9116 33350 9153
rect 33570 9259 33938 9298
rect 33570 9187 33938 9225
rect 33570 9116 33938 9153
rect 34158 9259 34526 9298
rect 34158 9187 34526 9225
rect 34158 9116 34526 9153
rect 34746 9259 35114 9298
rect 34746 9187 35114 9225
rect 34746 9116 35114 9153
rect 35334 9259 35702 9298
rect 35334 9187 35702 9225
rect 35334 9116 35702 9153
rect 35922 9259 36290 9298
rect 35922 9187 36290 9225
rect 35922 9116 36290 9153
rect 36510 9259 36878 9298
rect 36510 9187 36878 9225
rect 36510 9116 36878 9153
rect 37098 9259 37466 9298
rect 37098 9187 37466 9225
rect 37098 9116 37466 9153
rect 37686 9259 38054 9298
rect 37686 9187 38054 9225
rect 37686 9116 38054 9153
rect 38274 9259 38642 9298
rect 38274 9187 38642 9225
rect 38274 9116 38642 9153
rect 11226 8259 11594 8286
rect 11226 8209 11594 8225
rect 11814 8259 12182 8286
rect 11814 8209 12182 8225
rect 12402 8259 12770 8286
rect 12402 8209 12770 8225
rect 12990 8259 13358 8286
rect 12990 8209 13358 8225
rect 13578 8259 13946 8286
rect 13578 8209 13946 8225
rect 14166 8259 14534 8286
rect 14166 8209 14534 8225
rect 14754 8259 15122 8286
rect 14754 8209 15122 8225
rect 15342 8259 15710 8286
rect 15342 8209 15710 8225
rect 15930 8259 16298 8286
rect 15930 8209 16298 8225
rect 16518 8259 16886 8286
rect 16518 8209 16886 8225
rect 17106 8259 17474 8286
rect 17106 8209 17474 8225
rect 17694 8259 18062 8286
rect 17694 8209 18062 8225
rect 18282 8259 18650 8286
rect 18282 8209 18650 8225
rect 18870 8259 19238 8286
rect 18870 8209 19238 8225
rect 19458 8259 19826 8286
rect 19458 8209 19826 8225
rect 20046 8259 20414 8286
rect 20046 8209 20414 8225
rect 20634 8259 21002 8286
rect 20634 8209 21002 8225
rect 21222 8259 21590 8286
rect 21222 8209 21590 8225
rect 21810 8259 22178 8286
rect 21810 8209 22178 8225
rect 22986 8259 23354 8284
rect 22986 8209 23354 8225
rect 23574 8259 23942 8284
rect 23574 8209 23942 8225
rect 24162 8259 24530 8284
rect 24162 8209 24530 8225
rect 24750 8259 25118 8284
rect 24750 8209 25118 8225
rect 25338 8259 25706 8284
rect 25338 8209 25706 8225
rect 25926 8259 26294 8284
rect 25926 8209 26294 8225
rect 26514 8259 26882 8284
rect 26514 8209 26882 8225
rect 27102 8259 27470 8284
rect 27102 8209 27470 8225
rect 27690 8259 28058 8284
rect 27690 8209 28058 8225
rect 28278 8259 28646 8284
rect 28278 8209 28646 8225
rect 28866 8259 29234 8284
rect 28866 8209 29234 8225
rect 29454 8259 29822 8284
rect 29454 8209 29822 8225
rect 30042 8259 30410 8284
rect 30042 8209 30410 8225
rect 30630 8259 30998 8284
rect 30630 8209 30998 8225
rect 31218 8259 31586 8284
rect 31218 8209 31586 8225
rect 31806 8259 32174 8284
rect 31806 8209 32174 8225
rect 32394 8259 32762 8284
rect 32394 8209 32762 8225
rect 32982 8259 33350 8284
rect 32982 8209 33350 8225
rect 33570 8259 33938 8284
rect 33570 8209 33938 8225
rect 34158 8259 34526 8284
rect 34158 8209 34526 8225
rect 34746 8259 35114 8284
rect 34746 8209 35114 8225
rect 35334 8259 35702 8284
rect 35334 8209 35702 8225
rect 35922 8259 36290 8284
rect 35922 8209 36290 8225
rect 36510 8259 36878 8284
rect 36510 8209 36878 8225
rect 37098 8259 37466 8284
rect 37098 8209 37466 8225
rect 37686 8259 38054 8284
rect 37686 8209 38054 8225
rect 38274 8259 38642 8284
rect 38274 8209 38642 8225
<< polycont >>
rect 11226 27497 11594 27531
rect 11814 27497 12182 27531
rect 12402 27497 12770 27531
rect 12990 27497 13358 27531
rect 13578 27497 13946 27531
rect 14166 27497 14534 27531
rect 14754 27497 15122 27531
rect 15342 27497 15710 27531
rect 15930 27497 16298 27531
rect 16518 27497 16886 27531
rect 17106 27497 17474 27531
rect 17694 27497 18062 27531
rect 18282 27497 18650 27531
rect 18870 27497 19238 27531
rect 19458 27497 19826 27531
rect 20046 27497 20414 27531
rect 20634 27497 21002 27531
rect 21222 27497 21590 27531
rect 22986 27497 23354 27531
rect 23574 27497 23942 27531
rect 24162 27497 24530 27531
rect 24750 27497 25118 27531
rect 25338 27497 25706 27531
rect 25926 27497 26294 27531
rect 26514 27497 26882 27531
rect 27102 27497 27470 27531
rect 27690 27497 28058 27531
rect 28278 27497 28646 27531
rect 28866 27497 29234 27531
rect 29454 27497 29822 27531
rect 30042 27497 30410 27531
rect 30630 27497 30998 27531
rect 31218 27497 31586 27531
rect 31806 27497 32174 27531
rect 32394 27497 32762 27531
rect 32982 27497 33350 27531
rect 33570 27497 33938 27531
rect 34158 27497 34526 27531
rect 34746 27497 35114 27531
rect 35334 27497 35702 27531
rect 35922 27497 36290 27531
rect 36510 27497 36878 27531
rect 37098 27497 37466 27531
rect 37686 27497 38054 27531
rect 38274 27497 38642 27531
rect 11226 26569 11594 26603
rect 11226 26497 11594 26531
rect 11814 26569 12182 26603
rect 11814 26497 12182 26531
rect 12402 26569 12770 26603
rect 12402 26497 12770 26531
rect 12990 26569 13358 26603
rect 12990 26497 13358 26531
rect 13578 26569 13946 26603
rect 13578 26497 13946 26531
rect 14166 26569 14534 26603
rect 14166 26497 14534 26531
rect 14754 26569 15122 26603
rect 14754 26497 15122 26531
rect 15342 26569 15710 26603
rect 15342 26497 15710 26531
rect 15930 26569 16298 26603
rect 15930 26497 16298 26531
rect 16518 26569 16886 26603
rect 16518 26497 16886 26531
rect 17106 26569 17474 26603
rect 17106 26497 17474 26531
rect 17694 26569 18062 26603
rect 17694 26497 18062 26531
rect 18282 26569 18650 26603
rect 18282 26497 18650 26531
rect 18870 26569 19238 26603
rect 18870 26497 19238 26531
rect 19458 26569 19826 26603
rect 19458 26497 19826 26531
rect 20046 26569 20414 26603
rect 20046 26497 20414 26531
rect 20634 26569 21002 26603
rect 20634 26497 21002 26531
rect 21222 26569 21590 26603
rect 21222 26497 21590 26531
rect 21810 26569 22178 26603
rect 21810 26497 22178 26531
rect 22986 26569 23354 26603
rect 22986 26497 23354 26531
rect 23574 26569 23942 26603
rect 23574 26497 23942 26531
rect 24162 26569 24530 26603
rect 24162 26497 24530 26531
rect 24750 26569 25118 26603
rect 24750 26497 25118 26531
rect 25338 26569 25706 26603
rect 25338 26497 25706 26531
rect 25926 26569 26294 26603
rect 25926 26497 26294 26531
rect 26514 26569 26882 26603
rect 26514 26497 26882 26531
rect 27102 26569 27470 26603
rect 27102 26497 27470 26531
rect 27690 26569 28058 26603
rect 27690 26497 28058 26531
rect 28278 26569 28646 26603
rect 28278 26497 28646 26531
rect 28866 26569 29234 26603
rect 28866 26497 29234 26531
rect 29454 26569 29822 26603
rect 29454 26497 29822 26531
rect 30042 26569 30410 26603
rect 30042 26497 30410 26531
rect 30630 26569 30998 26603
rect 30630 26497 30998 26531
rect 31218 26569 31586 26603
rect 31218 26497 31586 26531
rect 31806 26569 32174 26603
rect 31806 26497 32174 26531
rect 32394 26569 32762 26603
rect 32394 26497 32762 26531
rect 32982 26569 33350 26603
rect 32982 26497 33350 26531
rect 33570 26569 33938 26603
rect 33570 26497 33938 26531
rect 34158 26569 34526 26603
rect 34158 26497 34526 26531
rect 34746 26569 35114 26603
rect 34746 26497 35114 26531
rect 35334 26569 35702 26603
rect 35334 26497 35702 26531
rect 35922 26569 36290 26603
rect 35922 26497 36290 26531
rect 36510 26569 36878 26603
rect 36510 26497 36878 26531
rect 37098 26569 37466 26603
rect 37098 26497 37466 26531
rect 37686 26569 38054 26603
rect 37686 26497 38054 26531
rect 38274 26569 38642 26603
rect 38274 26497 38642 26531
rect 10638 25569 11006 25603
rect 10638 25497 11006 25531
rect 11226 25569 11594 25603
rect 11226 25497 11594 25531
rect 11814 25569 12182 25603
rect 11814 25497 12182 25531
rect 12402 25569 12770 25603
rect 12402 25497 12770 25531
rect 12990 25569 13358 25603
rect 12990 25497 13358 25531
rect 13578 25569 13946 25603
rect 13578 25497 13946 25531
rect 14166 25569 14534 25603
rect 14166 25497 14534 25531
rect 14754 25569 15122 25603
rect 14754 25497 15122 25531
rect 15342 25569 15710 25603
rect 15342 25497 15710 25531
rect 15930 25569 16298 25603
rect 15930 25497 16298 25531
rect 16518 25569 16886 25603
rect 16518 25497 16886 25531
rect 17106 25569 17474 25603
rect 17106 25497 17474 25531
rect 17694 25569 18062 25603
rect 17694 25497 18062 25531
rect 18282 25569 18650 25603
rect 18282 25497 18650 25531
rect 18870 25569 19238 25603
rect 18870 25497 19238 25531
rect 19458 25569 19826 25603
rect 19458 25497 19826 25531
rect 20046 25569 20414 25603
rect 20046 25497 20414 25531
rect 20634 25569 21002 25603
rect 20634 25497 21002 25531
rect 21222 25569 21590 25603
rect 21222 25497 21590 25531
rect 21810 25569 22178 25603
rect 21810 25497 22178 25531
rect 23574 25569 23942 25603
rect 23574 25497 23942 25531
rect 24162 25569 24530 25603
rect 24162 25497 24530 25531
rect 24750 25569 25118 25603
rect 24750 25497 25118 25531
rect 25338 25569 25706 25603
rect 25338 25497 25706 25531
rect 25926 25569 26294 25603
rect 25926 25497 26294 25531
rect 26514 25569 26882 25603
rect 26514 25497 26882 25531
rect 27102 25569 27470 25603
rect 27102 25497 27470 25531
rect 27690 25569 28058 25603
rect 27690 25497 28058 25531
rect 28278 25569 28646 25603
rect 28278 25497 28646 25531
rect 28866 25569 29234 25603
rect 28866 25497 29234 25531
rect 29454 25569 29822 25603
rect 29454 25497 29822 25531
rect 30042 25569 30410 25603
rect 30042 25497 30410 25531
rect 30630 25569 30998 25603
rect 30630 25497 30998 25531
rect 31218 25569 31586 25603
rect 31218 25497 31586 25531
rect 31806 25569 32174 25603
rect 31806 25497 32174 25531
rect 32394 25569 32762 25603
rect 32394 25497 32762 25531
rect 32982 25569 33350 25603
rect 32982 25497 33350 25531
rect 33570 25569 33938 25603
rect 33570 25497 33938 25531
rect 34158 25569 34526 25603
rect 34158 25497 34526 25531
rect 34746 25569 35114 25603
rect 34746 25497 35114 25531
rect 35334 25569 35702 25603
rect 35334 25497 35702 25531
rect 35922 25569 36290 25603
rect 35922 25497 36290 25531
rect 36510 25569 36878 25603
rect 36510 25497 36878 25531
rect 37098 25569 37466 25603
rect 37098 25497 37466 25531
rect 37686 25569 38054 25603
rect 37686 25497 38054 25531
rect 38274 25569 38642 25603
rect 38274 25497 38642 25531
rect 11226 24569 11594 24603
rect 11814 24569 12182 24603
rect 12402 24569 12770 24603
rect 12990 24569 13358 24603
rect 13578 24569 13946 24603
rect 14166 24569 14534 24603
rect 14754 24569 15122 24603
rect 15342 24569 15710 24603
rect 15930 24569 16298 24603
rect 16518 24569 16886 24603
rect 17106 24569 17474 24603
rect 17694 24569 18062 24603
rect 18282 24569 18650 24603
rect 18870 24569 19238 24603
rect 19458 24569 19826 24603
rect 20046 24569 20414 24603
rect 20634 24569 21002 24603
rect 21222 24569 21590 24603
rect 21810 24569 22178 24603
rect 22986 24569 23354 24603
rect 23574 24569 23942 24603
rect 24162 24569 24530 24603
rect 24750 24569 25118 24603
rect 25338 24569 25706 24603
rect 25926 24569 26294 24603
rect 26514 24569 26882 24603
rect 27102 24569 27470 24603
rect 27690 24569 28058 24603
rect 28278 24569 28646 24603
rect 28866 24569 29234 24603
rect 29454 24569 29822 24603
rect 30042 24569 30410 24603
rect 30630 24569 30998 24603
rect 31218 24569 31586 24603
rect 31806 24569 32174 24603
rect 32394 24569 32762 24603
rect 32982 24569 33350 24603
rect 33570 24569 33938 24603
rect 34158 24569 34526 24603
rect 34746 24569 35114 24603
rect 35334 24569 35702 24603
rect 35922 24569 36290 24603
rect 36510 24569 36878 24603
rect 37098 24569 37466 24603
rect 37686 24569 38054 24603
rect 38274 24569 38642 24603
rect 11226 11153 11594 11187
rect 11814 11153 12182 11187
rect 12402 11153 12770 11187
rect 12990 11153 13358 11187
rect 13578 11153 13946 11187
rect 14166 11153 14534 11187
rect 14754 11153 15122 11187
rect 15342 11153 15710 11187
rect 15930 11153 16298 11187
rect 16518 11153 16886 11187
rect 17106 11153 17474 11187
rect 17694 11153 18062 11187
rect 18282 11153 18650 11187
rect 18870 11153 19238 11187
rect 19458 11153 19826 11187
rect 20046 11153 20414 11187
rect 20634 11153 21002 11187
rect 21222 11153 21590 11187
rect 21810 11153 22178 11187
rect 26514 11153 26882 11187
rect 27102 11153 27470 11187
rect 27690 11153 28058 11187
rect 28278 11153 28646 11187
rect 28866 11153 29234 11187
rect 29454 11153 29822 11187
rect 30042 11153 30410 11187
rect 30630 11153 30998 11187
rect 31218 11153 31586 11187
rect 31806 11153 32174 11187
rect 32394 11153 32762 11187
rect 32982 11153 33350 11187
rect 33570 11153 33938 11187
rect 34158 11153 34526 11187
rect 34746 11153 35114 11187
rect 35334 11153 35702 11187
rect 35922 11153 36290 11187
rect 36510 11153 36878 11187
rect 37098 11153 37466 11187
rect 37686 11153 38054 11187
rect 38274 11153 38642 11187
rect 11226 10225 11594 10259
rect 11226 10153 11594 10187
rect 11814 10225 12182 10259
rect 11814 10153 12182 10187
rect 12402 10225 12770 10259
rect 12402 10153 12770 10187
rect 12990 10225 13358 10259
rect 12990 10153 13358 10187
rect 13578 10225 13946 10259
rect 13578 10153 13946 10187
rect 14166 10225 14534 10259
rect 14166 10153 14534 10187
rect 14754 10225 15122 10259
rect 14754 10153 15122 10187
rect 15342 10225 15710 10259
rect 15342 10153 15710 10187
rect 15930 10225 16298 10259
rect 15930 10153 16298 10187
rect 16518 10225 16886 10259
rect 16518 10153 16886 10187
rect 17106 10225 17474 10259
rect 17106 10153 17474 10187
rect 17694 10225 18062 10259
rect 17694 10153 18062 10187
rect 18282 10225 18650 10259
rect 18282 10153 18650 10187
rect 18870 10225 19238 10259
rect 18870 10153 19238 10187
rect 19458 10225 19826 10259
rect 19458 10153 19826 10187
rect 20046 10225 20414 10259
rect 20046 10153 20414 10187
rect 20634 10225 21002 10259
rect 20634 10153 21002 10187
rect 21222 10225 21590 10259
rect 21222 10153 21590 10187
rect 21810 10225 22178 10259
rect 21810 10153 22178 10187
rect 22986 10225 23354 10259
rect 22986 10153 23354 10187
rect 23574 10225 23942 10259
rect 23574 10153 23942 10187
rect 24162 10225 24530 10259
rect 24162 10153 24530 10187
rect 24750 10225 25118 10259
rect 24750 10153 25118 10187
rect 25338 10225 25706 10259
rect 25338 10153 25706 10187
rect 25926 10225 26294 10259
rect 25926 10153 26294 10187
rect 26514 10225 26882 10259
rect 26514 10153 26882 10187
rect 27102 10225 27470 10259
rect 27102 10153 27470 10187
rect 27690 10225 28058 10259
rect 27690 10153 28058 10187
rect 28278 10225 28646 10259
rect 28278 10153 28646 10187
rect 28866 10225 29234 10259
rect 28866 10153 29234 10187
rect 29454 10225 29822 10259
rect 29454 10153 29822 10187
rect 30042 10225 30410 10259
rect 30042 10153 30410 10187
rect 30630 10225 30998 10259
rect 30630 10153 30998 10187
rect 31218 10225 31586 10259
rect 31218 10153 31586 10187
rect 31806 10225 32174 10259
rect 31806 10153 32174 10187
rect 32394 10225 32762 10259
rect 32394 10153 32762 10187
rect 32982 10225 33350 10259
rect 32982 10153 33350 10187
rect 33570 10225 33938 10259
rect 33570 10153 33938 10187
rect 34158 10225 34526 10259
rect 34158 10153 34526 10187
rect 34746 10225 35114 10259
rect 34746 10153 35114 10187
rect 35334 10225 35702 10259
rect 35334 10153 35702 10187
rect 35922 10225 36290 10259
rect 35922 10153 36290 10187
rect 36510 10225 36878 10259
rect 36510 10153 36878 10187
rect 37098 10225 37466 10259
rect 37098 10153 37466 10187
rect 37686 10225 38054 10259
rect 37686 10153 38054 10187
rect 38274 10225 38642 10259
rect 38274 10153 38642 10187
rect 10638 9225 11006 9259
rect 10638 9153 11006 9187
rect 11226 9225 11594 9259
rect 11226 9153 11594 9187
rect 11814 9225 12182 9259
rect 11814 9153 12182 9187
rect 12402 9225 12770 9259
rect 12402 9153 12770 9187
rect 12990 9225 13358 9259
rect 12990 9153 13358 9187
rect 13578 9225 13946 9259
rect 13578 9153 13946 9187
rect 14166 9225 14534 9259
rect 14166 9153 14534 9187
rect 14754 9225 15122 9259
rect 14754 9153 15122 9187
rect 15342 9225 15710 9259
rect 15342 9153 15710 9187
rect 15930 9225 16298 9259
rect 15930 9153 16298 9187
rect 16518 9225 16886 9259
rect 16518 9153 16886 9187
rect 17106 9225 17474 9259
rect 17106 9153 17474 9187
rect 17694 9225 18062 9259
rect 17694 9153 18062 9187
rect 18282 9225 18650 9259
rect 18282 9153 18650 9187
rect 18870 9225 19238 9259
rect 18870 9153 19238 9187
rect 19458 9225 19826 9259
rect 19458 9153 19826 9187
rect 20046 9225 20414 9259
rect 20046 9153 20414 9187
rect 20634 9225 21002 9259
rect 20634 9153 21002 9187
rect 21222 9225 21590 9259
rect 21222 9153 21590 9187
rect 21810 9225 22178 9259
rect 21810 9153 22178 9187
rect 22986 9225 23354 9259
rect 22986 9153 23354 9187
rect 23574 9225 23942 9259
rect 23574 9153 23942 9187
rect 24162 9225 24530 9259
rect 24162 9153 24530 9187
rect 24750 9225 25118 9259
rect 24750 9153 25118 9187
rect 25338 9225 25706 9259
rect 25338 9153 25706 9187
rect 25926 9225 26294 9259
rect 25926 9153 26294 9187
rect 26514 9225 26882 9259
rect 26514 9153 26882 9187
rect 27102 9225 27470 9259
rect 27102 9153 27470 9187
rect 27690 9225 28058 9259
rect 27690 9153 28058 9187
rect 28278 9225 28646 9259
rect 28278 9153 28646 9187
rect 28866 9225 29234 9259
rect 28866 9153 29234 9187
rect 29454 9225 29822 9259
rect 29454 9153 29822 9187
rect 30042 9225 30410 9259
rect 30042 9153 30410 9187
rect 30630 9225 30998 9259
rect 30630 9153 30998 9187
rect 31218 9225 31586 9259
rect 31218 9153 31586 9187
rect 31806 9225 32174 9259
rect 31806 9153 32174 9187
rect 32394 9225 32762 9259
rect 32394 9153 32762 9187
rect 32982 9225 33350 9259
rect 32982 9153 33350 9187
rect 33570 9225 33938 9259
rect 33570 9153 33938 9187
rect 34158 9225 34526 9259
rect 34158 9153 34526 9187
rect 34746 9225 35114 9259
rect 34746 9153 35114 9187
rect 35334 9225 35702 9259
rect 35334 9153 35702 9187
rect 35922 9225 36290 9259
rect 35922 9153 36290 9187
rect 36510 9225 36878 9259
rect 36510 9153 36878 9187
rect 37098 9225 37466 9259
rect 37098 9153 37466 9187
rect 37686 9225 38054 9259
rect 37686 9153 38054 9187
rect 38274 9225 38642 9259
rect 38274 9153 38642 9187
rect 11226 8225 11594 8259
rect 11814 8225 12182 8259
rect 12402 8225 12770 8259
rect 12990 8225 13358 8259
rect 13578 8225 13946 8259
rect 14166 8225 14534 8259
rect 14754 8225 15122 8259
rect 15342 8225 15710 8259
rect 15930 8225 16298 8259
rect 16518 8225 16886 8259
rect 17106 8225 17474 8259
rect 17694 8225 18062 8259
rect 18282 8225 18650 8259
rect 18870 8225 19238 8259
rect 19458 8225 19826 8259
rect 20046 8225 20414 8259
rect 20634 8225 21002 8259
rect 21222 8225 21590 8259
rect 21810 8225 22178 8259
rect 22986 8225 23354 8259
rect 23574 8225 23942 8259
rect 24162 8225 24530 8259
rect 24750 8225 25118 8259
rect 25338 8225 25706 8259
rect 25926 8225 26294 8259
rect 26514 8225 26882 8259
rect 27102 8225 27470 8259
rect 27690 8225 28058 8259
rect 28278 8225 28646 8259
rect 28866 8225 29234 8259
rect 29454 8225 29822 8259
rect 30042 8225 30410 8259
rect 30630 8225 30998 8259
rect 31218 8225 31586 8259
rect 31806 8225 32174 8259
rect 32394 8225 32762 8259
rect 32982 8225 33350 8259
rect 33570 8225 33938 8259
rect 34158 8225 34526 8259
rect 34746 8225 35114 8259
rect 35334 8225 35702 8259
rect 35922 8225 36290 8259
rect 36510 8225 36878 8259
rect 37098 8225 37466 8259
rect 37686 8225 38054 8259
rect 38274 8225 38642 8259
<< xpolycontact >>
rect 6785 28729 6855 29161
rect 6785 24897 6855 25329
rect 39789 26259 39859 26691
rect 39789 24027 39859 24459
rect 39789 22247 39859 22679
rect 39789 21015 39859 21447
<< xpolyres >>
rect 6785 25329 6855 28729
rect 39789 24459 39859 26259
rect 39789 21447 39859 22247
<< locali >>
rect 6655 29257 6751 29291
rect 6889 29257 6985 29291
rect 6655 29195 6689 29257
rect 6951 29195 6985 29257
rect 6655 24801 6689 24863
rect 11210 27531 11620 27532
rect 11210 27497 11226 27531
rect 11594 27497 11620 27531
rect 11210 27496 11620 27497
rect 11798 27531 12208 27532
rect 11798 27497 11814 27531
rect 12182 27497 12208 27531
rect 11798 27496 12208 27497
rect 12386 27531 12796 27532
rect 12386 27497 12402 27531
rect 12770 27497 12796 27531
rect 12386 27496 12796 27497
rect 12974 27531 13384 27532
rect 12974 27497 12990 27531
rect 13358 27497 13384 27531
rect 12974 27496 13384 27497
rect 13562 27531 13972 27532
rect 13562 27497 13578 27531
rect 13946 27497 13972 27531
rect 13562 27496 13972 27497
rect 14150 27531 14560 27532
rect 14150 27497 14166 27531
rect 14534 27497 14560 27531
rect 14150 27496 14560 27497
rect 14738 27531 15148 27532
rect 14738 27497 14754 27531
rect 15122 27497 15148 27531
rect 14738 27496 15148 27497
rect 15326 27531 15736 27532
rect 15326 27497 15342 27531
rect 15710 27497 15736 27531
rect 15326 27496 15736 27497
rect 15914 27531 16324 27532
rect 15914 27497 15930 27531
rect 16298 27497 16324 27531
rect 15914 27496 16324 27497
rect 16502 27531 16912 27532
rect 16502 27497 16518 27531
rect 16886 27497 16912 27531
rect 16502 27496 16912 27497
rect 17090 27531 17500 27532
rect 17090 27497 17106 27531
rect 17474 27497 17500 27531
rect 17090 27496 17500 27497
rect 17678 27531 18088 27532
rect 17678 27497 17694 27531
rect 18062 27497 18088 27531
rect 17678 27496 18088 27497
rect 18266 27531 18676 27532
rect 18266 27497 18282 27531
rect 18650 27497 18676 27531
rect 18266 27496 18676 27497
rect 18854 27531 19264 27532
rect 18854 27497 18870 27531
rect 19238 27497 19264 27531
rect 18854 27496 19264 27497
rect 19442 27531 19852 27532
rect 19442 27497 19458 27531
rect 19826 27497 19852 27531
rect 19442 27496 19852 27497
rect 20030 27531 20440 27532
rect 20030 27497 20046 27531
rect 20414 27497 20440 27531
rect 20030 27496 20440 27497
rect 20618 27531 21028 27532
rect 20618 27497 20634 27531
rect 21002 27497 21028 27531
rect 20618 27496 21028 27497
rect 21206 27531 21616 27532
rect 21206 27497 21222 27531
rect 21590 27497 21616 27531
rect 22974 27497 22986 27531
rect 23354 27497 23366 27531
rect 23562 27497 23574 27531
rect 23942 27497 23954 27531
rect 24150 27497 24162 27531
rect 24530 27497 24542 27531
rect 24738 27497 24750 27531
rect 25118 27497 25130 27531
rect 25326 27497 25338 27531
rect 25706 27497 25718 27531
rect 25914 27497 25926 27531
rect 26294 27497 26306 27531
rect 26502 27497 26514 27531
rect 26882 27497 26894 27531
rect 27090 27497 27102 27531
rect 27470 27497 27482 27531
rect 27678 27497 27690 27531
rect 28058 27497 28070 27531
rect 28266 27497 28278 27531
rect 28646 27497 28658 27531
rect 28854 27497 28866 27531
rect 29234 27497 29246 27531
rect 29442 27497 29454 27531
rect 29822 27497 29834 27531
rect 30030 27497 30042 27531
rect 30410 27497 30422 27531
rect 30618 27497 30630 27531
rect 30998 27497 31010 27531
rect 31206 27497 31218 27531
rect 31586 27497 31598 27531
rect 31794 27497 31806 27531
rect 32174 27497 32186 27531
rect 32382 27497 32394 27531
rect 32762 27497 32774 27531
rect 32970 27497 32982 27531
rect 33350 27497 33362 27531
rect 33558 27497 33570 27531
rect 33938 27497 33950 27531
rect 34146 27497 34158 27531
rect 34526 27497 34538 27531
rect 34734 27497 34746 27531
rect 35114 27497 35126 27531
rect 35322 27497 35334 27531
rect 35702 27497 35714 27531
rect 35910 27497 35922 27531
rect 36290 27497 36302 27531
rect 36498 27497 36510 27531
rect 36878 27497 36890 27531
rect 37086 27497 37098 27531
rect 37466 27497 37478 27531
rect 37674 27497 37686 27531
rect 38054 27497 38066 27531
rect 38262 27497 38274 27531
rect 38642 27497 38654 27531
rect 21206 27496 21616 27497
rect 39659 26787 39755 26821
rect 39893 26787 39989 26821
rect 39659 26725 39693 26787
rect 11214 26603 11606 26604
rect 11214 26569 11226 26603
rect 11594 26569 11606 26603
rect 11214 26531 11606 26569
rect 11214 26497 11226 26531
rect 11594 26497 11606 26531
rect 11214 26496 11606 26497
rect 11802 26603 12194 26604
rect 11802 26569 11814 26603
rect 12182 26569 12194 26603
rect 11802 26531 12194 26569
rect 11802 26497 11814 26531
rect 12182 26497 12194 26531
rect 11802 26496 12194 26497
rect 12390 26603 12782 26604
rect 12390 26569 12402 26603
rect 12770 26569 12782 26603
rect 12390 26531 12782 26569
rect 12390 26497 12402 26531
rect 12770 26497 12782 26531
rect 12390 26496 12782 26497
rect 12978 26603 13370 26604
rect 12978 26569 12990 26603
rect 13358 26569 13370 26603
rect 12978 26531 13370 26569
rect 12978 26497 12990 26531
rect 13358 26497 13370 26531
rect 12978 26496 13370 26497
rect 13566 26603 13958 26604
rect 13566 26569 13578 26603
rect 13946 26569 13958 26603
rect 13566 26531 13958 26569
rect 13566 26497 13578 26531
rect 13946 26497 13958 26531
rect 13566 26496 13958 26497
rect 14154 26603 14546 26604
rect 14154 26569 14166 26603
rect 14534 26569 14546 26603
rect 14154 26531 14546 26569
rect 14154 26497 14166 26531
rect 14534 26497 14546 26531
rect 14154 26496 14546 26497
rect 14742 26603 15134 26604
rect 14742 26569 14754 26603
rect 15122 26569 15134 26603
rect 14742 26531 15134 26569
rect 14742 26497 14754 26531
rect 15122 26497 15134 26531
rect 14742 26496 15134 26497
rect 15330 26603 15722 26604
rect 15330 26569 15342 26603
rect 15710 26569 15722 26603
rect 15330 26531 15722 26569
rect 15330 26497 15342 26531
rect 15710 26497 15722 26531
rect 15330 26496 15722 26497
rect 15918 26603 16310 26604
rect 15918 26569 15930 26603
rect 16298 26569 16310 26603
rect 15918 26531 16310 26569
rect 15918 26497 15930 26531
rect 16298 26497 16310 26531
rect 15918 26496 16310 26497
rect 16506 26603 16898 26604
rect 16506 26569 16518 26603
rect 16886 26569 16898 26603
rect 16506 26531 16898 26569
rect 16506 26497 16518 26531
rect 16886 26497 16898 26531
rect 16506 26496 16898 26497
rect 17094 26603 17486 26604
rect 17094 26569 17106 26603
rect 17474 26569 17486 26603
rect 17094 26531 17486 26569
rect 17094 26497 17106 26531
rect 17474 26497 17486 26531
rect 17094 26496 17486 26497
rect 17682 26603 18074 26604
rect 17682 26569 17694 26603
rect 18062 26569 18074 26603
rect 17682 26531 18074 26569
rect 17682 26497 17694 26531
rect 18062 26497 18074 26531
rect 17682 26496 18074 26497
rect 18270 26603 18662 26604
rect 18270 26569 18282 26603
rect 18650 26569 18662 26603
rect 18270 26531 18662 26569
rect 18270 26497 18282 26531
rect 18650 26497 18662 26531
rect 18270 26496 18662 26497
rect 18858 26603 19250 26604
rect 18858 26569 18870 26603
rect 19238 26569 19250 26603
rect 18858 26531 19250 26569
rect 18858 26497 18870 26531
rect 19238 26497 19250 26531
rect 18858 26496 19250 26497
rect 19446 26603 19838 26604
rect 19446 26569 19458 26603
rect 19826 26569 19838 26603
rect 19446 26531 19838 26569
rect 19446 26497 19458 26531
rect 19826 26497 19838 26531
rect 19446 26496 19838 26497
rect 20034 26603 20426 26604
rect 20034 26569 20046 26603
rect 20414 26569 20426 26603
rect 20034 26531 20426 26569
rect 20034 26497 20046 26531
rect 20414 26497 20426 26531
rect 20034 26496 20426 26497
rect 20622 26603 21014 26604
rect 20622 26569 20634 26603
rect 21002 26569 21014 26603
rect 20622 26531 21014 26569
rect 20622 26497 20634 26531
rect 21002 26497 21014 26531
rect 20622 26496 21014 26497
rect 21210 26603 21602 26604
rect 21210 26569 21222 26603
rect 21590 26569 21602 26603
rect 21210 26531 21602 26569
rect 21210 26497 21222 26531
rect 21590 26497 21602 26531
rect 21210 26496 21602 26497
rect 21798 26603 22190 26604
rect 21798 26569 21810 26603
rect 22178 26569 22190 26603
rect 22974 26569 22986 26603
rect 23562 26569 23574 26603
rect 24150 26569 24162 26603
rect 24738 26569 24750 26603
rect 25326 26569 25338 26603
rect 25914 26569 25926 26603
rect 26502 26569 26514 26603
rect 27090 26569 27102 26603
rect 27678 26569 27690 26603
rect 28266 26569 28278 26603
rect 28854 26569 28866 26603
rect 29442 26569 29454 26603
rect 30030 26569 30042 26603
rect 30618 26569 30630 26603
rect 31206 26569 31218 26603
rect 31794 26569 31806 26603
rect 32382 26569 32394 26603
rect 32970 26569 32982 26603
rect 33558 26569 33570 26603
rect 34146 26569 34158 26603
rect 34734 26569 34746 26603
rect 35322 26569 35334 26603
rect 35910 26569 35922 26603
rect 36498 26569 36510 26603
rect 37086 26569 37098 26603
rect 37674 26569 37686 26603
rect 38262 26569 38274 26603
rect 21798 26531 22190 26569
rect 21798 26497 21810 26531
rect 22178 26497 22190 26531
rect 22974 26497 22986 26531
rect 23562 26497 23574 26531
rect 24150 26497 24162 26531
rect 24738 26497 24750 26531
rect 25326 26497 25338 26531
rect 25914 26497 25926 26531
rect 26502 26497 26514 26531
rect 27090 26497 27102 26531
rect 27678 26497 27690 26531
rect 28266 26497 28278 26531
rect 28854 26497 28866 26531
rect 29442 26497 29454 26531
rect 30030 26497 30042 26531
rect 30618 26497 30630 26531
rect 31206 26497 31218 26531
rect 31794 26497 31806 26531
rect 32382 26497 32394 26531
rect 32970 26497 32982 26531
rect 33558 26497 33570 26531
rect 34146 26497 34158 26531
rect 34734 26497 34746 26531
rect 35322 26497 35334 26531
rect 35910 26497 35922 26531
rect 36498 26497 36510 26531
rect 37086 26497 37098 26531
rect 37674 26497 37686 26531
rect 38262 26497 38274 26531
rect 21798 26496 22190 26497
rect 10638 25603 11006 25604
rect 10638 25531 11006 25569
rect 10638 25496 11006 25497
rect 11226 25603 11594 25604
rect 11226 25531 11594 25569
rect 11226 25496 11594 25497
rect 11814 25603 12182 25604
rect 11814 25531 12182 25569
rect 11814 25496 12182 25497
rect 12402 25603 12770 25604
rect 12402 25531 12770 25569
rect 12402 25496 12770 25497
rect 12990 25603 13358 25604
rect 12990 25531 13358 25569
rect 12990 25496 13358 25497
rect 13578 25603 13946 25604
rect 13578 25531 13946 25569
rect 13578 25496 13946 25497
rect 14166 25603 14534 25604
rect 14166 25531 14534 25569
rect 14166 25496 14534 25497
rect 14754 25603 15122 25604
rect 14754 25531 15122 25569
rect 14754 25496 15122 25497
rect 15342 25603 15710 25604
rect 15342 25531 15710 25569
rect 15342 25496 15710 25497
rect 15930 25603 16298 25604
rect 15930 25531 16298 25569
rect 15930 25496 16298 25497
rect 16518 25603 16886 25604
rect 16518 25531 16886 25569
rect 16518 25496 16886 25497
rect 17106 25603 17474 25604
rect 17106 25531 17474 25569
rect 17106 25496 17474 25497
rect 17694 25603 18062 25604
rect 17694 25531 18062 25569
rect 17694 25496 18062 25497
rect 18282 25603 18650 25604
rect 18282 25531 18650 25569
rect 18282 25496 18650 25497
rect 18870 25603 19238 25604
rect 18870 25531 19238 25569
rect 18870 25496 19238 25497
rect 19458 25603 19826 25604
rect 19458 25531 19826 25569
rect 19458 25496 19826 25497
rect 20046 25603 20414 25604
rect 20046 25531 20414 25569
rect 20046 25496 20414 25497
rect 20634 25603 21002 25604
rect 20634 25531 21002 25569
rect 20634 25496 21002 25497
rect 21222 25603 21590 25604
rect 21222 25531 21590 25569
rect 21222 25496 21590 25497
rect 21810 25603 22178 25604
rect 21810 25531 22178 25569
rect 21810 25496 22178 25497
rect 6951 24801 6985 24863
rect 6655 24767 6751 24801
rect 6889 24767 6985 24801
rect 11210 24603 11594 24604
rect 11210 24569 11226 24603
rect 11210 24568 11594 24569
rect 11798 24603 12182 24604
rect 11798 24569 11814 24603
rect 11798 24568 12182 24569
rect 12386 24603 12770 24604
rect 12386 24569 12402 24603
rect 12386 24568 12770 24569
rect 12974 24603 13358 24604
rect 12974 24569 12990 24603
rect 12974 24568 13358 24569
rect 13562 24603 13946 24604
rect 13562 24569 13578 24603
rect 13562 24568 13946 24569
rect 14150 24603 14534 24604
rect 14150 24569 14166 24603
rect 14150 24568 14534 24569
rect 14738 24603 15122 24604
rect 14738 24569 14754 24603
rect 14738 24568 15122 24569
rect 15326 24603 15710 24604
rect 15326 24569 15342 24603
rect 15326 24568 15710 24569
rect 15914 24603 16298 24604
rect 15914 24569 15930 24603
rect 15914 24568 16298 24569
rect 16502 24603 16886 24604
rect 16502 24569 16518 24603
rect 16502 24568 16886 24569
rect 17090 24603 17474 24604
rect 17090 24569 17106 24603
rect 17090 24568 17474 24569
rect 17678 24603 18062 24604
rect 17678 24569 17694 24603
rect 17678 24568 18062 24569
rect 18266 24603 18650 24604
rect 18266 24569 18282 24603
rect 18266 24568 18650 24569
rect 18854 24603 19238 24604
rect 18854 24569 18870 24603
rect 18854 24568 19238 24569
rect 19442 24603 19826 24604
rect 19442 24569 19458 24603
rect 19442 24568 19826 24569
rect 20030 24603 20414 24604
rect 20030 24569 20046 24603
rect 20030 24568 20414 24569
rect 20618 24603 21002 24604
rect 20618 24569 20634 24603
rect 20618 24568 21002 24569
rect 21206 24603 21590 24604
rect 21206 24569 21222 24603
rect 21206 24568 21590 24569
rect 21794 24603 22178 24604
rect 21794 24569 21810 24603
rect 21794 24568 22178 24569
rect 39955 26725 39989 26787
rect 39659 23986 39693 23993
rect 38978 23931 39693 23986
rect 39955 23931 39989 23993
rect 38978 23900 39755 23931
rect 39659 23897 39755 23900
rect 39893 23897 39989 23931
rect 39659 22775 39755 22809
rect 39893 22775 39989 22809
rect 39659 22713 39693 22775
rect 38980 21368 39659 21606
rect 39955 22713 39989 22775
rect 39659 20919 39693 20981
rect 39955 20919 39989 20981
rect 39659 20885 39755 20919
rect 39893 20885 39989 20919
rect 11226 11187 11594 11188
rect 11226 11152 11594 11153
rect 11814 11187 12182 11188
rect 11814 11152 12182 11153
rect 12402 11187 12770 11188
rect 12402 11152 12770 11153
rect 12990 11187 13358 11188
rect 12990 11152 13358 11153
rect 13578 11187 13946 11188
rect 13578 11152 13946 11153
rect 14166 11187 14534 11188
rect 14166 11152 14534 11153
rect 14754 11187 15122 11188
rect 14754 11152 15122 11153
rect 15342 11187 15710 11188
rect 15342 11152 15710 11153
rect 15930 11187 16298 11188
rect 15930 11152 16298 11153
rect 16518 11187 16886 11188
rect 16518 11152 16886 11153
rect 17106 11187 17474 11188
rect 17106 11152 17474 11153
rect 17694 11187 18062 11188
rect 17694 11152 18062 11153
rect 18282 11187 18650 11188
rect 18282 11152 18650 11153
rect 18870 11187 19238 11188
rect 18870 11152 19238 11153
rect 19458 11187 19826 11188
rect 19458 11152 19826 11153
rect 20046 11187 20414 11188
rect 20046 11152 20414 11153
rect 20634 11187 21002 11188
rect 20634 11152 21002 11153
rect 21222 11187 21590 11188
rect 21222 11152 21590 11153
rect 21810 11187 22178 11188
rect 26502 11153 26514 11187
rect 26882 11153 26894 11187
rect 27090 11153 27102 11187
rect 27470 11153 27482 11187
rect 27678 11153 27690 11187
rect 28058 11153 28070 11187
rect 28266 11153 28278 11187
rect 28646 11153 28658 11187
rect 28854 11153 28866 11187
rect 29234 11153 29246 11187
rect 29442 11153 29454 11187
rect 29822 11153 29834 11187
rect 30030 11153 30042 11187
rect 30410 11153 30422 11187
rect 30618 11153 30630 11187
rect 30998 11153 31010 11187
rect 31206 11153 31218 11187
rect 31586 11153 31598 11187
rect 31794 11153 31806 11187
rect 32174 11153 32186 11187
rect 32382 11153 32394 11187
rect 32762 11153 32774 11187
rect 32970 11153 32982 11187
rect 33350 11153 33362 11187
rect 33558 11153 33570 11187
rect 33938 11153 33950 11187
rect 34146 11153 34158 11187
rect 34526 11153 34538 11187
rect 34734 11153 34746 11187
rect 35114 11153 35126 11187
rect 35322 11153 35334 11187
rect 35702 11153 35714 11187
rect 35910 11153 35922 11187
rect 36290 11153 36302 11187
rect 36498 11153 36510 11187
rect 36878 11153 36890 11187
rect 37086 11153 37098 11187
rect 37466 11153 37478 11187
rect 37674 11153 37686 11187
rect 38054 11153 38066 11187
rect 38262 11153 38274 11187
rect 38642 11153 38654 11187
rect 21810 11152 22178 11153
rect 11214 10259 11606 10260
rect 11214 10225 11226 10259
rect 11594 10225 11606 10259
rect 11214 10187 11606 10225
rect 11214 10153 11226 10187
rect 11594 10153 11606 10187
rect 11214 10152 11606 10153
rect 11802 10259 12194 10260
rect 11802 10225 11814 10259
rect 12182 10225 12194 10259
rect 11802 10187 12194 10225
rect 11802 10153 11814 10187
rect 12182 10153 12194 10187
rect 11802 10152 12194 10153
rect 12390 10259 12782 10260
rect 12390 10225 12402 10259
rect 12770 10225 12782 10259
rect 12390 10187 12782 10225
rect 12390 10153 12402 10187
rect 12770 10153 12782 10187
rect 12390 10152 12782 10153
rect 12978 10259 13370 10260
rect 12978 10225 12990 10259
rect 13358 10225 13370 10259
rect 12978 10187 13370 10225
rect 12978 10153 12990 10187
rect 13358 10153 13370 10187
rect 12978 10152 13370 10153
rect 13566 10259 13958 10260
rect 13566 10225 13578 10259
rect 13946 10225 13958 10259
rect 13566 10187 13958 10225
rect 13566 10153 13578 10187
rect 13946 10153 13958 10187
rect 13566 10152 13958 10153
rect 14154 10259 14546 10260
rect 14154 10225 14166 10259
rect 14534 10225 14546 10259
rect 14154 10187 14546 10225
rect 14154 10153 14166 10187
rect 14534 10153 14546 10187
rect 14154 10152 14546 10153
rect 14742 10259 15134 10260
rect 14742 10225 14754 10259
rect 15122 10225 15134 10259
rect 14742 10187 15134 10225
rect 14742 10153 14754 10187
rect 15122 10153 15134 10187
rect 14742 10152 15134 10153
rect 15330 10259 15722 10260
rect 15330 10225 15342 10259
rect 15710 10225 15722 10259
rect 15330 10187 15722 10225
rect 15330 10153 15342 10187
rect 15710 10153 15722 10187
rect 15330 10152 15722 10153
rect 15918 10259 16310 10260
rect 15918 10225 15930 10259
rect 16298 10225 16310 10259
rect 15918 10187 16310 10225
rect 15918 10153 15930 10187
rect 16298 10153 16310 10187
rect 15918 10152 16310 10153
rect 16506 10259 16898 10260
rect 16506 10225 16518 10259
rect 16886 10225 16898 10259
rect 16506 10187 16898 10225
rect 16506 10153 16518 10187
rect 16886 10153 16898 10187
rect 16506 10152 16898 10153
rect 17094 10259 17486 10260
rect 17094 10225 17106 10259
rect 17474 10225 17486 10259
rect 17094 10187 17486 10225
rect 17094 10153 17106 10187
rect 17474 10153 17486 10187
rect 17094 10152 17486 10153
rect 17682 10259 18074 10260
rect 17682 10225 17694 10259
rect 18062 10225 18074 10259
rect 17682 10187 18074 10225
rect 17682 10153 17694 10187
rect 18062 10153 18074 10187
rect 17682 10152 18074 10153
rect 18270 10259 18662 10260
rect 18270 10225 18282 10259
rect 18650 10225 18662 10259
rect 18270 10187 18662 10225
rect 18270 10153 18282 10187
rect 18650 10153 18662 10187
rect 18270 10152 18662 10153
rect 18858 10259 19250 10260
rect 18858 10225 18870 10259
rect 19238 10225 19250 10259
rect 18858 10187 19250 10225
rect 18858 10153 18870 10187
rect 19238 10153 19250 10187
rect 18858 10152 19250 10153
rect 19446 10259 19838 10260
rect 19446 10225 19458 10259
rect 19826 10225 19838 10259
rect 19446 10187 19838 10225
rect 19446 10153 19458 10187
rect 19826 10153 19838 10187
rect 19446 10152 19838 10153
rect 20034 10259 20426 10260
rect 20034 10225 20046 10259
rect 20414 10225 20426 10259
rect 20034 10187 20426 10225
rect 20034 10153 20046 10187
rect 20414 10153 20426 10187
rect 20034 10152 20426 10153
rect 20622 10259 21014 10260
rect 20622 10225 20634 10259
rect 21002 10225 21014 10259
rect 20622 10187 21014 10225
rect 20622 10153 20634 10187
rect 21002 10153 21014 10187
rect 20622 10152 21014 10153
rect 21210 10259 21602 10260
rect 21210 10225 21222 10259
rect 21590 10225 21602 10259
rect 21210 10187 21602 10225
rect 21210 10153 21222 10187
rect 21590 10153 21602 10187
rect 21210 10152 21602 10153
rect 21798 10259 22190 10260
rect 21798 10225 21810 10259
rect 22178 10225 22190 10259
rect 22974 10225 22986 10259
rect 23562 10225 23574 10259
rect 24150 10225 24162 10259
rect 24738 10225 24750 10259
rect 25326 10225 25338 10259
rect 25914 10225 25926 10259
rect 26502 10225 26514 10259
rect 27090 10225 27102 10259
rect 27678 10225 27690 10259
rect 28266 10225 28278 10259
rect 28854 10225 28866 10259
rect 29442 10225 29454 10259
rect 30030 10225 30042 10259
rect 30618 10225 30630 10259
rect 31206 10225 31218 10259
rect 31794 10225 31806 10259
rect 32382 10225 32394 10259
rect 32970 10225 32982 10259
rect 33558 10225 33570 10259
rect 34146 10225 34158 10259
rect 34734 10225 34746 10259
rect 35322 10225 35334 10259
rect 35910 10225 35922 10259
rect 36498 10225 36510 10259
rect 37086 10225 37098 10259
rect 37674 10225 37686 10259
rect 38262 10225 38274 10259
rect 21798 10187 22190 10225
rect 21798 10153 21810 10187
rect 22178 10153 22190 10187
rect 22974 10153 22986 10187
rect 23562 10153 23574 10187
rect 24150 10153 24162 10187
rect 24738 10153 24750 10187
rect 25326 10153 25338 10187
rect 25914 10153 25926 10187
rect 26502 10153 26514 10187
rect 27090 10153 27102 10187
rect 27678 10153 27690 10187
rect 28266 10153 28278 10187
rect 28854 10153 28866 10187
rect 29442 10153 29454 10187
rect 30030 10153 30042 10187
rect 30618 10153 30630 10187
rect 31206 10153 31218 10187
rect 31794 10153 31806 10187
rect 32382 10153 32394 10187
rect 32970 10153 32982 10187
rect 33558 10153 33570 10187
rect 34146 10153 34158 10187
rect 34734 10153 34746 10187
rect 35322 10153 35334 10187
rect 35910 10153 35922 10187
rect 36498 10153 36510 10187
rect 37086 10153 37098 10187
rect 37674 10153 37686 10187
rect 38262 10153 38274 10187
rect 21798 10152 22190 10153
rect 10638 9259 11006 9260
rect 10638 9187 11006 9225
rect 10638 9152 11006 9153
rect 11226 9259 11594 9260
rect 11226 9187 11594 9225
rect 11226 9152 11594 9153
rect 11814 9259 12182 9260
rect 11814 9187 12182 9225
rect 11814 9152 12182 9153
rect 12402 9259 12770 9260
rect 12402 9187 12770 9225
rect 12402 9152 12770 9153
rect 12990 9259 13358 9260
rect 12990 9187 13358 9225
rect 12990 9152 13358 9153
rect 13578 9259 13946 9260
rect 13578 9187 13946 9225
rect 13578 9152 13946 9153
rect 14166 9259 14534 9260
rect 14166 9187 14534 9225
rect 14166 9152 14534 9153
rect 14754 9259 15122 9260
rect 14754 9187 15122 9225
rect 14754 9152 15122 9153
rect 15342 9259 15710 9260
rect 15342 9187 15710 9225
rect 15342 9152 15710 9153
rect 15930 9259 16298 9260
rect 15930 9187 16298 9225
rect 15930 9152 16298 9153
rect 16518 9259 16886 9260
rect 16518 9187 16886 9225
rect 16518 9152 16886 9153
rect 17106 9259 17474 9260
rect 17106 9187 17474 9225
rect 17106 9152 17474 9153
rect 17694 9259 18062 9260
rect 17694 9187 18062 9225
rect 17694 9152 18062 9153
rect 18282 9259 18650 9260
rect 18282 9187 18650 9225
rect 18282 9152 18650 9153
rect 18870 9259 19238 9260
rect 18870 9187 19238 9225
rect 18870 9152 19238 9153
rect 19458 9259 19826 9260
rect 19458 9187 19826 9225
rect 19458 9152 19826 9153
rect 20046 9259 20414 9260
rect 20046 9187 20414 9225
rect 20046 9152 20414 9153
rect 20634 9259 21002 9260
rect 20634 9187 21002 9225
rect 20634 9152 21002 9153
rect 21222 9259 21590 9260
rect 21222 9187 21590 9225
rect 21222 9152 21590 9153
rect 21810 9259 22178 9260
rect 21810 9187 22178 9225
rect 21810 9152 22178 9153
rect 11226 8259 11594 8260
rect 11226 8224 11594 8225
rect 11814 8259 12182 8260
rect 11814 8224 12182 8225
rect 12402 8259 12770 8260
rect 12402 8224 12770 8225
rect 12990 8259 13358 8260
rect 12990 8224 13358 8225
rect 13578 8259 13946 8260
rect 13578 8224 13946 8225
rect 14166 8259 14534 8260
rect 14166 8224 14534 8225
rect 14754 8259 15122 8260
rect 14754 8224 15122 8225
rect 15342 8259 15710 8260
rect 15342 8224 15710 8225
rect 15930 8259 16298 8260
rect 15930 8224 16298 8225
rect 16518 8259 16886 8260
rect 16518 8224 16886 8225
rect 17106 8259 17474 8260
rect 17106 8224 17474 8225
rect 17694 8259 18062 8260
rect 17694 8224 18062 8225
rect 18282 8259 18650 8260
rect 18282 8224 18650 8225
rect 18870 8259 19238 8260
rect 18870 8224 19238 8225
rect 19458 8259 19826 8260
rect 19458 8224 19826 8225
rect 20046 8259 20414 8260
rect 20046 8224 20414 8225
rect 20634 8259 21002 8260
rect 20634 8224 21002 8225
rect 21222 8259 21590 8260
rect 21222 8224 21590 8225
rect 21810 8259 22178 8260
rect 21810 8224 22178 8225
<< viali >>
rect 6801 28746 6839 29143
rect 6801 24915 6839 25312
rect 11226 27497 11594 27531
rect 11814 27497 12182 27531
rect 12402 27497 12770 27531
rect 12990 27497 13358 27531
rect 13578 27497 13946 27531
rect 14166 27497 14534 27531
rect 14754 27497 15122 27531
rect 15342 27497 15710 27531
rect 15930 27497 16298 27531
rect 16518 27497 16886 27531
rect 17106 27497 17474 27531
rect 17694 27497 18062 27531
rect 18282 27497 18650 27531
rect 18870 27497 19238 27531
rect 19458 27497 19826 27531
rect 20046 27497 20414 27531
rect 20634 27497 21002 27531
rect 21222 27497 21590 27531
rect 22986 27497 23354 27531
rect 23574 27497 23942 27531
rect 24162 27497 24530 27531
rect 24750 27497 25118 27531
rect 25338 27497 25706 27531
rect 25926 27497 26294 27531
rect 26514 27497 26882 27531
rect 27102 27497 27470 27531
rect 27690 27497 28058 27531
rect 28278 27497 28646 27531
rect 28866 27497 29234 27531
rect 29454 27497 29822 27531
rect 30042 27497 30410 27531
rect 30630 27497 30998 27531
rect 31218 27497 31586 27531
rect 31806 27497 32174 27531
rect 32394 27497 32762 27531
rect 32982 27497 33350 27531
rect 33570 27497 33938 27531
rect 34158 27497 34526 27531
rect 34746 27497 35114 27531
rect 35334 27497 35702 27531
rect 35922 27497 36290 27531
rect 36510 27497 36878 27531
rect 37098 27497 37466 27531
rect 37686 27497 38054 27531
rect 38274 27497 38642 27531
rect 11226 26569 11594 26603
rect 11226 26497 11594 26531
rect 11814 26569 12182 26603
rect 11814 26497 12182 26531
rect 12402 26569 12770 26603
rect 12402 26497 12770 26531
rect 12990 26569 13358 26603
rect 12990 26497 13358 26531
rect 13578 26569 13946 26603
rect 13578 26497 13946 26531
rect 14166 26569 14534 26603
rect 14166 26497 14534 26531
rect 14754 26569 15122 26603
rect 14754 26497 15122 26531
rect 15342 26569 15710 26603
rect 15342 26497 15710 26531
rect 15930 26569 16298 26603
rect 15930 26497 16298 26531
rect 16518 26569 16886 26603
rect 16518 26497 16886 26531
rect 17106 26569 17474 26603
rect 17106 26497 17474 26531
rect 17694 26569 18062 26603
rect 17694 26497 18062 26531
rect 18282 26569 18650 26603
rect 18282 26497 18650 26531
rect 18870 26569 19238 26603
rect 18870 26497 19238 26531
rect 19458 26569 19826 26603
rect 19458 26497 19826 26531
rect 20046 26569 20414 26603
rect 20046 26497 20414 26531
rect 20634 26569 21002 26603
rect 20634 26497 21002 26531
rect 21222 26569 21590 26603
rect 21222 26497 21590 26531
rect 21810 26569 22178 26603
rect 22986 26569 23354 26603
rect 23574 26569 23942 26603
rect 24162 26569 24530 26603
rect 24750 26569 25118 26603
rect 25338 26569 25706 26603
rect 25926 26569 26294 26603
rect 26514 26569 26882 26603
rect 27102 26569 27470 26603
rect 27690 26569 28058 26603
rect 28278 26569 28646 26603
rect 28866 26569 29234 26603
rect 29454 26569 29822 26603
rect 30042 26569 30410 26603
rect 30630 26569 30998 26603
rect 31218 26569 31586 26603
rect 31806 26569 32174 26603
rect 32394 26569 32762 26603
rect 32982 26569 33350 26603
rect 33570 26569 33938 26603
rect 34158 26569 34526 26603
rect 34746 26569 35114 26603
rect 35334 26569 35702 26603
rect 35922 26569 36290 26603
rect 36510 26569 36878 26603
rect 37098 26569 37466 26603
rect 37686 26569 38054 26603
rect 38274 26569 38642 26603
rect 21810 26497 22178 26531
rect 22986 26497 23354 26531
rect 23574 26497 23942 26531
rect 24162 26497 24530 26531
rect 24750 26497 25118 26531
rect 25338 26497 25706 26531
rect 25926 26497 26294 26531
rect 26514 26497 26882 26531
rect 27102 26497 27470 26531
rect 27690 26497 28058 26531
rect 28278 26497 28646 26531
rect 28866 26497 29234 26531
rect 29454 26497 29822 26531
rect 30042 26497 30410 26531
rect 30630 26497 30998 26531
rect 31218 26497 31586 26531
rect 31806 26497 32174 26531
rect 32394 26497 32762 26531
rect 32982 26497 33350 26531
rect 33570 26497 33938 26531
rect 34158 26497 34526 26531
rect 34746 26497 35114 26531
rect 35334 26497 35702 26531
rect 35922 26497 36290 26531
rect 36510 26497 36878 26531
rect 37098 26497 37466 26531
rect 37686 26497 38054 26531
rect 38274 26497 38642 26531
rect 10638 25569 11006 25603
rect 10638 25497 11006 25531
rect 11226 25569 11594 25603
rect 11226 25497 11594 25531
rect 11814 25569 12182 25603
rect 11814 25497 12182 25531
rect 12402 25569 12770 25603
rect 12402 25497 12770 25531
rect 12990 25569 13358 25603
rect 12990 25497 13358 25531
rect 13578 25569 13946 25603
rect 13578 25497 13946 25531
rect 14166 25569 14534 25603
rect 14166 25497 14534 25531
rect 14754 25569 15122 25603
rect 14754 25497 15122 25531
rect 15342 25569 15710 25603
rect 15342 25497 15710 25531
rect 15930 25569 16298 25603
rect 15930 25497 16298 25531
rect 16518 25569 16886 25603
rect 16518 25497 16886 25531
rect 17106 25569 17474 25603
rect 17106 25497 17474 25531
rect 17694 25569 18062 25603
rect 17694 25497 18062 25531
rect 18282 25569 18650 25603
rect 18282 25497 18650 25531
rect 18870 25569 19238 25603
rect 18870 25497 19238 25531
rect 19458 25569 19826 25603
rect 19458 25497 19826 25531
rect 20046 25569 20414 25603
rect 20046 25497 20414 25531
rect 20634 25569 21002 25603
rect 20634 25497 21002 25531
rect 21222 25569 21590 25603
rect 21222 25497 21590 25531
rect 21810 25569 22178 25603
rect 23574 25569 23942 25603
rect 24162 25569 24530 25603
rect 24750 25569 25118 25603
rect 25338 25569 25706 25603
rect 25926 25569 26294 25603
rect 26514 25569 26882 25603
rect 27102 25569 27470 25603
rect 27690 25569 28058 25603
rect 28278 25569 28646 25603
rect 28866 25569 29234 25603
rect 29454 25569 29822 25603
rect 30042 25569 30410 25603
rect 30630 25569 30998 25603
rect 31218 25569 31586 25603
rect 31806 25569 32174 25603
rect 32394 25569 32762 25603
rect 32982 25569 33350 25603
rect 33570 25569 33938 25603
rect 34158 25569 34526 25603
rect 34746 25569 35114 25603
rect 35334 25569 35702 25603
rect 35922 25569 36290 25603
rect 36510 25569 36878 25603
rect 37098 25569 37466 25603
rect 37686 25569 38054 25603
rect 38274 25569 38642 25603
rect 21810 25497 22178 25531
rect 23574 25497 23942 25531
rect 24162 25497 24530 25531
rect 24750 25497 25118 25531
rect 25338 25497 25706 25531
rect 25926 25497 26294 25531
rect 26514 25497 26882 25531
rect 27102 25497 27470 25531
rect 27690 25497 28058 25531
rect 28278 25497 28646 25531
rect 28866 25497 29234 25531
rect 29454 25497 29822 25531
rect 30042 25497 30410 25531
rect 30630 25497 30998 25531
rect 31218 25497 31586 25531
rect 31806 25497 32174 25531
rect 32394 25497 32762 25531
rect 32982 25497 33350 25531
rect 33570 25497 33938 25531
rect 34158 25497 34526 25531
rect 34746 25497 35114 25531
rect 35334 25497 35702 25531
rect 35922 25497 36290 25531
rect 36510 25497 36878 25531
rect 37098 25497 37466 25531
rect 37686 25497 38054 25531
rect 38274 25497 38642 25531
rect 11226 24569 11594 24603
rect 11814 24569 12182 24603
rect 12402 24569 12770 24603
rect 12990 24569 13358 24603
rect 13578 24569 13946 24603
rect 14166 24569 14534 24603
rect 14754 24569 15122 24603
rect 15342 24569 15710 24603
rect 15930 24569 16298 24603
rect 16518 24569 16886 24603
rect 17106 24569 17474 24603
rect 17694 24569 18062 24603
rect 18282 24569 18650 24603
rect 18870 24569 19238 24603
rect 19458 24569 19826 24603
rect 20046 24569 20414 24603
rect 20634 24569 21002 24603
rect 21222 24569 21590 24603
rect 21810 24569 22178 24603
rect 22986 24569 23354 24603
rect 23574 24569 23942 24603
rect 24162 24569 24530 24603
rect 24750 24569 25118 24603
rect 25338 24569 25706 24603
rect 25926 24569 26294 24603
rect 26514 24569 26882 24603
rect 27102 24569 27470 24603
rect 27690 24569 28058 24603
rect 28278 24569 28646 24603
rect 28866 24569 29234 24603
rect 29454 24569 29822 24603
rect 30042 24569 30410 24603
rect 30630 24569 30998 24603
rect 31218 24569 31586 24603
rect 31806 24569 32174 24603
rect 32394 24569 32762 24603
rect 32982 24569 33350 24603
rect 33570 24569 33938 24603
rect 34158 24569 34526 24603
rect 34746 24569 35114 24603
rect 35334 24569 35702 24603
rect 35922 24569 36290 24603
rect 36510 24569 36878 24603
rect 37098 24569 37466 24603
rect 37686 24569 38054 24603
rect 38274 24569 38642 24603
rect 38666 23772 38978 24038
rect 39805 26276 39843 26673
rect 39805 24045 39843 24442
rect 37832 20906 38980 22370
rect 39805 22264 39843 22661
rect 39805 21033 39843 21430
rect 11226 11153 11594 11187
rect 11814 11153 12182 11187
rect 12402 11153 12770 11187
rect 12990 11153 13358 11187
rect 13578 11153 13946 11187
rect 14166 11153 14534 11187
rect 14754 11153 15122 11187
rect 15342 11153 15710 11187
rect 15930 11153 16298 11187
rect 16518 11153 16886 11187
rect 17106 11153 17474 11187
rect 17694 11153 18062 11187
rect 18282 11153 18650 11187
rect 18870 11153 19238 11187
rect 19458 11153 19826 11187
rect 20046 11153 20414 11187
rect 20634 11153 21002 11187
rect 21222 11153 21590 11187
rect 21810 11153 22178 11187
rect 26514 11153 26882 11187
rect 27102 11153 27470 11187
rect 27690 11153 28058 11187
rect 28278 11153 28646 11187
rect 28866 11153 29234 11187
rect 29454 11153 29822 11187
rect 30042 11153 30410 11187
rect 30630 11153 30998 11187
rect 31218 11153 31586 11187
rect 31806 11153 32174 11187
rect 32394 11153 32762 11187
rect 32982 11153 33350 11187
rect 33570 11153 33938 11187
rect 34158 11153 34526 11187
rect 34746 11153 35114 11187
rect 35334 11153 35702 11187
rect 35922 11153 36290 11187
rect 36510 11153 36878 11187
rect 37098 11153 37466 11187
rect 37686 11153 38054 11187
rect 38274 11153 38642 11187
rect 11226 10225 11594 10259
rect 11226 10153 11594 10187
rect 11814 10225 12182 10259
rect 11814 10153 12182 10187
rect 12402 10225 12770 10259
rect 12402 10153 12770 10187
rect 12990 10225 13358 10259
rect 12990 10153 13358 10187
rect 13578 10225 13946 10259
rect 13578 10153 13946 10187
rect 14166 10225 14534 10259
rect 14166 10153 14534 10187
rect 14754 10225 15122 10259
rect 14754 10153 15122 10187
rect 15342 10225 15710 10259
rect 15342 10153 15710 10187
rect 15930 10225 16298 10259
rect 15930 10153 16298 10187
rect 16518 10225 16886 10259
rect 16518 10153 16886 10187
rect 17106 10225 17474 10259
rect 17106 10153 17474 10187
rect 17694 10225 18062 10259
rect 17694 10153 18062 10187
rect 18282 10225 18650 10259
rect 18282 10153 18650 10187
rect 18870 10225 19238 10259
rect 18870 10153 19238 10187
rect 19458 10225 19826 10259
rect 19458 10153 19826 10187
rect 20046 10225 20414 10259
rect 20046 10153 20414 10187
rect 20634 10225 21002 10259
rect 20634 10153 21002 10187
rect 21222 10225 21590 10259
rect 21222 10153 21590 10187
rect 21810 10225 22178 10259
rect 22986 10225 23354 10259
rect 23574 10225 23942 10259
rect 24162 10225 24530 10259
rect 24750 10225 25118 10259
rect 25338 10225 25706 10259
rect 25926 10225 26294 10259
rect 26514 10225 26882 10259
rect 27102 10225 27470 10259
rect 27690 10225 28058 10259
rect 28278 10225 28646 10259
rect 28866 10225 29234 10259
rect 29454 10225 29822 10259
rect 30042 10225 30410 10259
rect 30630 10225 30998 10259
rect 31218 10225 31586 10259
rect 31806 10225 32174 10259
rect 32394 10225 32762 10259
rect 32982 10225 33350 10259
rect 33570 10225 33938 10259
rect 34158 10225 34526 10259
rect 34746 10225 35114 10259
rect 35334 10225 35702 10259
rect 35922 10225 36290 10259
rect 36510 10225 36878 10259
rect 37098 10225 37466 10259
rect 37686 10225 38054 10259
rect 38274 10225 38642 10259
rect 21810 10153 22178 10187
rect 22986 10153 23354 10187
rect 23574 10153 23942 10187
rect 24162 10153 24530 10187
rect 24750 10153 25118 10187
rect 25338 10153 25706 10187
rect 25926 10153 26294 10187
rect 26514 10153 26882 10187
rect 27102 10153 27470 10187
rect 27690 10153 28058 10187
rect 28278 10153 28646 10187
rect 28866 10153 29234 10187
rect 29454 10153 29822 10187
rect 30042 10153 30410 10187
rect 30630 10153 30998 10187
rect 31218 10153 31586 10187
rect 31806 10153 32174 10187
rect 32394 10153 32762 10187
rect 32982 10153 33350 10187
rect 33570 10153 33938 10187
rect 34158 10153 34526 10187
rect 34746 10153 35114 10187
rect 35334 10153 35702 10187
rect 35922 10153 36290 10187
rect 36510 10153 36878 10187
rect 37098 10153 37466 10187
rect 37686 10153 38054 10187
rect 38274 10153 38642 10187
rect 10638 9225 11006 9259
rect 10638 9153 11006 9187
rect 11226 9225 11594 9259
rect 11226 9153 11594 9187
rect 11814 9225 12182 9259
rect 11814 9153 12182 9187
rect 12402 9225 12770 9259
rect 12402 9153 12770 9187
rect 12990 9225 13358 9259
rect 12990 9153 13358 9187
rect 13578 9225 13946 9259
rect 13578 9153 13946 9187
rect 14166 9225 14534 9259
rect 14166 9153 14534 9187
rect 14754 9225 15122 9259
rect 14754 9153 15122 9187
rect 15342 9225 15710 9259
rect 15342 9153 15710 9187
rect 15930 9225 16298 9259
rect 15930 9153 16298 9187
rect 16518 9225 16886 9259
rect 16518 9153 16886 9187
rect 17106 9225 17474 9259
rect 17106 9153 17474 9187
rect 17694 9225 18062 9259
rect 17694 9153 18062 9187
rect 18282 9225 18650 9259
rect 18282 9153 18650 9187
rect 18870 9225 19238 9259
rect 18870 9153 19238 9187
rect 19458 9225 19826 9259
rect 19458 9153 19826 9187
rect 20046 9225 20414 9259
rect 20046 9153 20414 9187
rect 20634 9225 21002 9259
rect 20634 9153 21002 9187
rect 21222 9225 21590 9259
rect 21222 9153 21590 9187
rect 21810 9225 22178 9259
rect 22986 9225 23354 9259
rect 23574 9225 23942 9259
rect 24162 9225 24530 9259
rect 24750 9225 25118 9259
rect 25338 9225 25706 9259
rect 25926 9225 26294 9259
rect 26514 9225 26882 9259
rect 27102 9225 27470 9259
rect 27690 9225 28058 9259
rect 28278 9225 28646 9259
rect 28866 9225 29234 9259
rect 29454 9225 29822 9259
rect 30042 9225 30410 9259
rect 30630 9225 30998 9259
rect 31218 9225 31586 9259
rect 31806 9225 32174 9259
rect 32394 9225 32762 9259
rect 32982 9225 33350 9259
rect 33570 9225 33938 9259
rect 34158 9225 34526 9259
rect 34746 9225 35114 9259
rect 35334 9225 35702 9259
rect 35922 9225 36290 9259
rect 36510 9225 36878 9259
rect 37098 9225 37466 9259
rect 37686 9225 38054 9259
rect 38274 9225 38642 9259
rect 21810 9153 22178 9187
rect 22986 9153 23354 9187
rect 23574 9153 23942 9187
rect 24162 9153 24530 9187
rect 24750 9153 25118 9187
rect 25338 9153 25706 9187
rect 25926 9153 26294 9187
rect 26514 9153 26882 9187
rect 27102 9153 27470 9187
rect 27690 9153 28058 9187
rect 28278 9153 28646 9187
rect 28866 9153 29234 9187
rect 29454 9153 29822 9187
rect 30042 9153 30410 9187
rect 30630 9153 30998 9187
rect 31218 9153 31586 9187
rect 31806 9153 32174 9187
rect 32394 9153 32762 9187
rect 32982 9153 33350 9187
rect 33570 9153 33938 9187
rect 34158 9153 34526 9187
rect 34746 9153 35114 9187
rect 35334 9153 35702 9187
rect 35922 9153 36290 9187
rect 36510 9153 36878 9187
rect 37098 9153 37466 9187
rect 37686 9153 38054 9187
rect 38274 9153 38642 9187
rect 11226 8225 11594 8259
rect 11814 8225 12182 8259
rect 12402 8225 12770 8259
rect 12990 8225 13358 8259
rect 13578 8225 13946 8259
rect 14166 8225 14534 8259
rect 14754 8225 15122 8259
rect 15342 8225 15710 8259
rect 15930 8225 16298 8259
rect 16518 8225 16886 8259
rect 17106 8225 17474 8259
rect 17694 8225 18062 8259
rect 18282 8225 18650 8259
rect 18870 8225 19238 8259
rect 19458 8225 19826 8259
rect 20046 8225 20414 8259
rect 20634 8225 21002 8259
rect 21222 8225 21590 8259
rect 21810 8225 22178 8259
rect 22986 8225 23354 8259
rect 23574 8225 23942 8259
rect 24162 8225 24530 8259
rect 24750 8225 25118 8259
rect 25338 8225 25706 8259
rect 25926 8225 26294 8259
rect 26514 8225 26882 8259
rect 27102 8225 27470 8259
rect 27690 8225 28058 8259
rect 28278 8225 28646 8259
rect 28866 8225 29234 8259
rect 29454 8225 29822 8259
rect 30042 8225 30410 8259
rect 30630 8225 30998 8259
rect 31218 8225 31586 8259
rect 31806 8225 32174 8259
rect 32394 8225 32762 8259
rect 32982 8225 33350 8259
rect 33570 8225 33938 8259
rect 34158 8225 34526 8259
rect 34746 8225 35114 8259
rect 35334 8225 35702 8259
rect 35922 8225 36290 8259
rect 36510 8225 36878 8259
rect 37098 8225 37466 8259
rect 37686 8225 38054 8259
rect 38274 8225 38642 8259
<< metal1 >>
rect 6784 29143 10486 29250
rect 6784 28746 6801 29143
rect 6839 28746 10486 29143
rect 6784 28728 10486 28746
rect 36888 28402 37756 29084
rect 38416 28388 39860 28662
rect 10612 27490 10622 27548
rect 11022 27490 11032 27548
rect 11200 27490 11210 27548
rect 11610 27490 11620 27548
rect 11788 27490 11798 27548
rect 12198 27490 12208 27548
rect 12376 27490 12386 27548
rect 12786 27490 12796 27548
rect 12964 27490 12974 27548
rect 13374 27490 13384 27548
rect 13552 27490 13562 27548
rect 13962 27490 13972 27548
rect 14140 27490 14150 27548
rect 14550 27490 14560 27548
rect 14728 27490 14738 27548
rect 15138 27490 15148 27548
rect 15316 27490 15326 27548
rect 15726 27490 15736 27548
rect 15904 27490 15914 27548
rect 16314 27490 16324 27548
rect 16492 27490 16502 27548
rect 16902 27490 16912 27548
rect 17080 27490 17090 27548
rect 17490 27490 17500 27548
rect 17668 27490 17678 27548
rect 18078 27490 18088 27548
rect 18256 27490 18266 27548
rect 18666 27490 18676 27548
rect 18844 27490 18854 27548
rect 19254 27490 19264 27548
rect 19432 27490 19442 27548
rect 19842 27490 19852 27548
rect 20020 27490 20030 27548
rect 20430 27490 20440 27548
rect 20608 27490 20618 27548
rect 21018 27490 21028 27548
rect 21196 27490 21206 27548
rect 21606 27490 21616 27548
rect 21792 27486 21802 27542
rect 22178 27486 22188 27542
rect 22388 27488 22398 27542
rect 22766 27488 22776 27542
rect 22976 27537 22986 27542
rect 22974 27491 22986 27537
rect 23354 27537 23364 27542
rect 23564 27537 23574 27542
rect 22976 27488 22986 27491
rect 23354 27491 23366 27537
rect 23562 27491 23574 27537
rect 23942 27537 23952 27542
rect 24152 27537 24162 27542
rect 23354 27488 23364 27491
rect 23564 27488 23574 27491
rect 23942 27491 23954 27537
rect 24150 27491 24162 27537
rect 24530 27537 24540 27542
rect 24740 27537 24750 27542
rect 23942 27488 23952 27491
rect 24152 27488 24162 27491
rect 24530 27491 24542 27537
rect 24738 27491 24750 27537
rect 25118 27537 25128 27542
rect 25328 27537 25338 27542
rect 24530 27488 24540 27491
rect 24740 27488 24750 27491
rect 25118 27491 25130 27537
rect 25326 27491 25338 27537
rect 25706 27537 25716 27542
rect 25916 27537 25926 27542
rect 25118 27488 25128 27491
rect 25328 27488 25338 27491
rect 25706 27491 25718 27537
rect 25914 27491 25926 27537
rect 26294 27537 26304 27542
rect 26504 27537 26514 27542
rect 25706 27488 25716 27491
rect 25916 27488 25926 27491
rect 26294 27491 26306 27537
rect 26502 27491 26514 27537
rect 26882 27537 26892 27542
rect 27092 27537 27102 27542
rect 26294 27488 26304 27491
rect 26504 27488 26514 27491
rect 26882 27491 26894 27537
rect 27090 27491 27102 27537
rect 27470 27537 27480 27542
rect 27680 27537 27690 27542
rect 26882 27488 26892 27491
rect 27092 27488 27102 27491
rect 27470 27491 27482 27537
rect 27678 27491 27690 27537
rect 28058 27537 28068 27542
rect 28268 27537 28278 27542
rect 27470 27488 27480 27491
rect 27680 27488 27690 27491
rect 28058 27491 28070 27537
rect 28266 27491 28278 27537
rect 28646 27537 28656 27542
rect 28856 27537 28866 27542
rect 28058 27488 28068 27491
rect 28268 27488 28278 27491
rect 28646 27491 28658 27537
rect 28854 27491 28866 27537
rect 29234 27537 29244 27542
rect 29444 27537 29454 27542
rect 28646 27488 28656 27491
rect 28856 27488 28866 27491
rect 29234 27491 29246 27537
rect 29442 27491 29454 27537
rect 29822 27537 29832 27542
rect 30032 27537 30042 27542
rect 29234 27488 29244 27491
rect 29444 27488 29454 27491
rect 29822 27491 29834 27537
rect 30030 27491 30042 27537
rect 30410 27537 30420 27542
rect 30620 27537 30630 27542
rect 29822 27488 29832 27491
rect 30032 27488 30042 27491
rect 30410 27491 30422 27537
rect 30618 27491 30630 27537
rect 30998 27537 31008 27542
rect 31208 27537 31218 27542
rect 30410 27488 30420 27491
rect 30620 27488 30630 27491
rect 30998 27491 31010 27537
rect 31206 27491 31218 27537
rect 31586 27537 31596 27542
rect 31796 27537 31806 27542
rect 30998 27488 31008 27491
rect 31208 27488 31218 27491
rect 31586 27491 31598 27537
rect 31794 27491 31806 27537
rect 32174 27537 32184 27542
rect 32384 27537 32394 27542
rect 31586 27488 31596 27491
rect 31796 27488 31806 27491
rect 32174 27491 32186 27537
rect 32382 27491 32394 27537
rect 32762 27537 32772 27542
rect 32972 27537 32982 27542
rect 32174 27488 32184 27491
rect 32384 27488 32394 27491
rect 32762 27491 32774 27537
rect 32970 27491 32982 27537
rect 33350 27537 33360 27542
rect 33560 27537 33570 27542
rect 32762 27488 32772 27491
rect 32972 27488 32982 27491
rect 33350 27491 33362 27537
rect 33558 27491 33570 27537
rect 33938 27537 33948 27542
rect 34148 27537 34158 27542
rect 33350 27488 33360 27491
rect 33560 27488 33570 27491
rect 33938 27491 33950 27537
rect 34146 27491 34158 27537
rect 34526 27537 34536 27542
rect 34736 27537 34746 27542
rect 33938 27488 33948 27491
rect 34148 27488 34158 27491
rect 34526 27491 34538 27537
rect 34734 27491 34746 27537
rect 35114 27537 35124 27542
rect 35324 27537 35334 27542
rect 34526 27488 34536 27491
rect 34736 27488 34746 27491
rect 35114 27491 35126 27537
rect 35322 27491 35334 27537
rect 35702 27537 35712 27542
rect 35912 27537 35922 27542
rect 35114 27488 35124 27491
rect 35324 27488 35334 27491
rect 35702 27491 35714 27537
rect 35910 27491 35922 27537
rect 36290 27537 36300 27542
rect 36500 27537 36510 27542
rect 35702 27488 35712 27491
rect 35912 27488 35922 27491
rect 36290 27491 36302 27537
rect 36498 27491 36510 27537
rect 36878 27537 36888 27542
rect 37088 27537 37098 27542
rect 36290 27488 36300 27491
rect 36500 27488 36510 27491
rect 36878 27491 36890 27537
rect 37086 27491 37098 27537
rect 37466 27537 37476 27542
rect 37676 27537 37686 27542
rect 36878 27488 36888 27491
rect 37088 27488 37098 27491
rect 37466 27491 37478 27537
rect 37674 27491 37686 27537
rect 38054 27537 38064 27542
rect 38264 27537 38274 27542
rect 37466 27488 37476 27491
rect 37676 27488 37686 27491
rect 38054 27491 38066 27537
rect 38262 27491 38274 27537
rect 38642 27537 38652 27542
rect 38054 27488 38064 27491
rect 38264 27488 38274 27491
rect 38642 27491 38654 27537
rect 38642 27488 38652 27491
rect 39788 26673 39860 28388
rect 39788 26662 39805 26673
rect 11214 26604 11606 26609
rect 10628 26490 10638 26604
rect 11006 26490 11016 26604
rect 11214 26491 11226 26604
rect 11216 26490 11226 26491
rect 11594 26491 11606 26604
rect 11802 26604 12194 26609
rect 11802 26491 11814 26604
rect 11594 26490 11604 26491
rect 11804 26490 11814 26491
rect 12182 26491 12194 26604
rect 12390 26604 12782 26609
rect 12390 26491 12402 26604
rect 12182 26490 12192 26491
rect 12392 26490 12402 26491
rect 12770 26491 12782 26604
rect 12978 26604 13370 26609
rect 12978 26491 12990 26604
rect 12770 26490 12780 26491
rect 12980 26490 12990 26491
rect 13358 26491 13370 26604
rect 13566 26604 13958 26609
rect 13566 26491 13578 26604
rect 13358 26490 13368 26491
rect 13568 26490 13578 26491
rect 13946 26491 13958 26604
rect 14154 26604 14546 26609
rect 14154 26491 14166 26604
rect 13946 26490 13956 26491
rect 14156 26490 14166 26491
rect 14534 26491 14546 26604
rect 14742 26604 15134 26609
rect 14742 26491 14754 26604
rect 14534 26490 14544 26491
rect 14744 26490 14754 26491
rect 15122 26491 15134 26604
rect 15330 26604 15722 26609
rect 15330 26491 15342 26604
rect 15122 26490 15132 26491
rect 15332 26490 15342 26491
rect 15710 26491 15722 26604
rect 15918 26604 16310 26609
rect 15918 26491 15930 26604
rect 15710 26490 15720 26491
rect 15920 26490 15930 26491
rect 16298 26491 16310 26604
rect 16506 26604 16898 26609
rect 16506 26491 16518 26604
rect 16298 26490 16308 26491
rect 16508 26490 16518 26491
rect 16886 26491 16898 26604
rect 17094 26604 17486 26609
rect 17094 26491 17106 26604
rect 16886 26490 16896 26491
rect 17096 26490 17106 26491
rect 17474 26491 17486 26604
rect 17682 26604 18074 26609
rect 17682 26491 17694 26604
rect 17474 26490 17484 26491
rect 17684 26490 17694 26491
rect 18062 26491 18074 26604
rect 18270 26604 18662 26609
rect 18270 26491 18282 26604
rect 18062 26490 18072 26491
rect 18272 26490 18282 26491
rect 18650 26491 18662 26604
rect 18858 26604 19250 26609
rect 18858 26491 18870 26604
rect 18650 26490 18660 26491
rect 18860 26490 18870 26491
rect 19238 26491 19250 26604
rect 19446 26604 19838 26609
rect 19446 26491 19458 26604
rect 19238 26490 19248 26491
rect 19448 26490 19458 26491
rect 19826 26491 19838 26604
rect 20034 26604 20426 26609
rect 20034 26491 20046 26604
rect 19826 26490 19836 26491
rect 20036 26490 20046 26491
rect 20414 26491 20426 26604
rect 20622 26604 21014 26609
rect 20622 26491 20634 26604
rect 20414 26490 20424 26491
rect 20624 26490 20634 26491
rect 21002 26491 21014 26604
rect 21210 26604 21602 26609
rect 21210 26491 21222 26604
rect 21002 26490 21012 26491
rect 21212 26490 21222 26491
rect 21590 26491 21602 26604
rect 21798 26604 22190 26609
rect 22974 26604 23354 26609
rect 21798 26491 21810 26604
rect 21590 26490 21600 26491
rect 21800 26490 21810 26491
rect 22178 26491 22190 26604
rect 22388 26496 22398 26604
rect 22766 26496 22776 26604
rect 22974 26496 22986 26604
rect 22974 26491 23354 26496
rect 23562 26604 23942 26609
rect 23562 26496 23574 26604
rect 23562 26491 23942 26496
rect 24150 26604 24530 26609
rect 24150 26496 24162 26604
rect 24150 26491 24530 26496
rect 24738 26604 25118 26609
rect 24738 26496 24750 26604
rect 24738 26491 25118 26496
rect 25326 26604 25706 26609
rect 25326 26496 25338 26604
rect 25326 26491 25706 26496
rect 25914 26604 26294 26609
rect 25914 26496 25926 26604
rect 25914 26491 26294 26496
rect 26502 26604 26882 26609
rect 26502 26496 26514 26604
rect 26502 26491 26882 26496
rect 27090 26604 27470 26609
rect 27090 26496 27102 26604
rect 27090 26491 27470 26496
rect 27678 26604 28058 26609
rect 27678 26496 27690 26604
rect 27678 26491 28058 26496
rect 28266 26604 28646 26609
rect 28266 26496 28278 26604
rect 28266 26491 28646 26496
rect 28854 26604 29234 26609
rect 28854 26496 28866 26604
rect 28854 26491 29234 26496
rect 29442 26604 29822 26609
rect 29442 26496 29454 26604
rect 29442 26491 29822 26496
rect 30030 26604 30410 26609
rect 30030 26496 30042 26604
rect 30030 26491 30410 26496
rect 30618 26604 30998 26609
rect 30618 26496 30630 26604
rect 30618 26491 30998 26496
rect 31206 26604 31586 26609
rect 31206 26496 31218 26604
rect 31206 26491 31586 26496
rect 31794 26604 32174 26609
rect 31794 26496 31806 26604
rect 31794 26491 32174 26496
rect 32382 26604 32762 26609
rect 32382 26496 32394 26604
rect 32382 26491 32762 26496
rect 32970 26604 33350 26609
rect 32970 26496 32982 26604
rect 32970 26491 33350 26496
rect 33558 26604 33938 26609
rect 33558 26496 33570 26604
rect 33558 26491 33938 26496
rect 34146 26604 34526 26609
rect 34146 26496 34158 26604
rect 34146 26491 34526 26496
rect 34734 26604 35114 26609
rect 34734 26496 34746 26604
rect 34734 26491 35114 26496
rect 35322 26604 35702 26609
rect 35322 26496 35334 26604
rect 35322 26491 35702 26496
rect 35910 26604 36290 26609
rect 35910 26496 35922 26604
rect 35910 26491 36290 26496
rect 36498 26604 36878 26609
rect 36498 26496 36510 26604
rect 36498 26491 36878 26496
rect 37086 26604 37466 26609
rect 37086 26496 37098 26604
rect 37086 26491 37466 26496
rect 37674 26604 38054 26609
rect 37674 26496 37686 26604
rect 37674 26491 38054 26496
rect 38262 26604 38642 26609
rect 38262 26496 38274 26604
rect 38262 26491 38642 26496
rect 22178 26490 22188 26491
rect 39799 26276 39805 26662
rect 39843 26662 39860 26673
rect 39843 26276 39849 26662
rect 39799 26264 39849 26276
rect 10638 25604 11006 25609
rect 11226 25604 11594 25609
rect 11814 25604 12182 25609
rect 11216 25496 11226 25604
rect 11594 25496 11604 25604
rect 10638 25491 11006 25496
rect 11226 25491 11594 25496
rect 11814 25491 12182 25496
rect 12402 25604 12770 25609
rect 12402 25491 12770 25496
rect 12990 25604 13358 25609
rect 12990 25491 13358 25496
rect 13578 25604 13946 25609
rect 13578 25491 13946 25496
rect 14166 25604 14534 25609
rect 14166 25491 14534 25496
rect 14754 25604 15122 25609
rect 14754 25491 15122 25496
rect 15342 25604 15710 25609
rect 15342 25491 15710 25496
rect 15930 25604 16298 25609
rect 15930 25491 16298 25496
rect 16518 25604 16886 25609
rect 16518 25491 16886 25496
rect 17106 25604 17474 25609
rect 17106 25491 17474 25496
rect 17694 25604 18062 25609
rect 17694 25491 18062 25496
rect 18282 25604 18650 25609
rect 18282 25491 18650 25496
rect 18870 25604 19238 25609
rect 18870 25491 19238 25496
rect 19458 25604 19826 25609
rect 19458 25491 19826 25496
rect 20046 25604 20414 25609
rect 20046 25491 20414 25496
rect 20634 25604 21002 25609
rect 20634 25491 21002 25496
rect 21222 25604 21590 25609
rect 21222 25491 21590 25496
rect 21810 25604 22178 25609
rect 23574 25606 23942 25609
rect 22410 25496 22420 25604
rect 22732 25496 22742 25604
rect 21810 25491 22178 25496
rect 23010 25494 23020 25606
rect 23318 25494 23328 25606
rect 23574 25603 23608 25606
rect 23906 25603 23942 25606
rect 23574 25531 23608 25569
rect 23906 25531 23942 25569
rect 23574 25494 23608 25497
rect 23906 25494 23942 25497
rect 23574 25491 23942 25494
rect 24162 25606 24530 25609
rect 24162 25603 24196 25606
rect 24494 25603 24530 25606
rect 24162 25531 24196 25569
rect 24494 25531 24530 25569
rect 24162 25494 24196 25497
rect 24494 25494 24530 25497
rect 24162 25491 24530 25494
rect 24750 25606 25118 25609
rect 24750 25603 24784 25606
rect 25082 25603 25118 25606
rect 24750 25531 24784 25569
rect 25082 25531 25118 25569
rect 24750 25494 24784 25497
rect 25082 25494 25118 25497
rect 24750 25491 25118 25494
rect 25338 25606 25706 25609
rect 25338 25603 25372 25606
rect 25670 25603 25706 25606
rect 25338 25531 25372 25569
rect 25670 25531 25706 25569
rect 25338 25494 25372 25497
rect 25670 25494 25706 25497
rect 25338 25491 25706 25494
rect 25926 25606 26294 25609
rect 25926 25603 25960 25606
rect 26258 25603 26294 25606
rect 25926 25531 25960 25569
rect 26258 25531 26294 25569
rect 25926 25494 25960 25497
rect 26258 25494 26294 25497
rect 25926 25491 26294 25494
rect 26514 25606 26882 25609
rect 26514 25603 26548 25606
rect 26846 25603 26882 25606
rect 26514 25531 26548 25569
rect 26846 25531 26882 25569
rect 26514 25494 26548 25497
rect 26846 25494 26882 25497
rect 26514 25491 26882 25494
rect 27102 25606 27470 25609
rect 27102 25603 27136 25606
rect 27434 25603 27470 25606
rect 27102 25531 27136 25569
rect 27434 25531 27470 25569
rect 27102 25494 27136 25497
rect 27434 25494 27470 25497
rect 27102 25491 27470 25494
rect 27690 25606 28058 25609
rect 27690 25603 27724 25606
rect 28022 25603 28058 25606
rect 27690 25531 27724 25569
rect 28022 25531 28058 25569
rect 27690 25494 27724 25497
rect 28022 25494 28058 25497
rect 27690 25491 28058 25494
rect 28278 25606 28646 25609
rect 28278 25603 28312 25606
rect 28610 25603 28646 25606
rect 28278 25531 28312 25569
rect 28610 25531 28646 25569
rect 28278 25494 28312 25497
rect 28610 25494 28646 25497
rect 28278 25491 28646 25494
rect 28866 25606 29234 25609
rect 28866 25603 28900 25606
rect 29198 25603 29234 25606
rect 28866 25531 28900 25569
rect 29198 25531 29234 25569
rect 28866 25494 28900 25497
rect 29198 25494 29234 25497
rect 28866 25491 29234 25494
rect 29454 25606 29822 25609
rect 29454 25603 29488 25606
rect 29786 25603 29822 25606
rect 29454 25531 29488 25569
rect 29786 25531 29822 25569
rect 29454 25494 29488 25497
rect 29786 25494 29822 25497
rect 29454 25491 29822 25494
rect 30042 25606 30410 25609
rect 30042 25603 30076 25606
rect 30374 25603 30410 25606
rect 30042 25531 30076 25569
rect 30374 25531 30410 25569
rect 30042 25494 30076 25497
rect 30374 25494 30410 25497
rect 30042 25491 30410 25494
rect 30630 25606 30998 25609
rect 30630 25603 30664 25606
rect 30962 25603 30998 25606
rect 30630 25531 30664 25569
rect 30962 25531 30998 25569
rect 30630 25494 30664 25497
rect 30962 25494 30998 25497
rect 30630 25491 30998 25494
rect 31218 25606 31586 25609
rect 31218 25603 31252 25606
rect 31550 25603 31586 25606
rect 31218 25531 31252 25569
rect 31550 25531 31586 25569
rect 31218 25494 31252 25497
rect 31550 25494 31586 25497
rect 31218 25491 31586 25494
rect 31806 25606 32174 25609
rect 31806 25603 31840 25606
rect 32138 25603 32174 25606
rect 31806 25531 31840 25569
rect 32138 25531 32174 25569
rect 31806 25494 31840 25497
rect 32138 25494 32174 25497
rect 31806 25491 32174 25494
rect 32394 25606 32762 25609
rect 32394 25603 32428 25606
rect 32726 25603 32762 25606
rect 32394 25531 32428 25569
rect 32726 25531 32762 25569
rect 32394 25494 32428 25497
rect 32726 25494 32762 25497
rect 32394 25491 32762 25494
rect 32982 25606 33350 25609
rect 32982 25603 33016 25606
rect 33314 25603 33350 25606
rect 32982 25531 33016 25569
rect 33314 25531 33350 25569
rect 32982 25494 33016 25497
rect 33314 25494 33350 25497
rect 32982 25491 33350 25494
rect 33570 25606 33938 25609
rect 33570 25603 33604 25606
rect 33902 25603 33938 25606
rect 33570 25531 33604 25569
rect 33902 25531 33938 25569
rect 33570 25494 33604 25497
rect 33902 25494 33938 25497
rect 33570 25491 33938 25494
rect 34158 25606 34526 25609
rect 34158 25603 34192 25606
rect 34490 25603 34526 25606
rect 34158 25531 34192 25569
rect 34490 25531 34526 25569
rect 34158 25494 34192 25497
rect 34490 25494 34526 25497
rect 34158 25491 34526 25494
rect 34746 25606 35114 25609
rect 34746 25603 34780 25606
rect 35078 25603 35114 25606
rect 34746 25531 34780 25569
rect 35078 25531 35114 25569
rect 34746 25494 34780 25497
rect 35078 25494 35114 25497
rect 34746 25491 35114 25494
rect 35334 25606 35702 25609
rect 35334 25603 35368 25606
rect 35666 25603 35702 25606
rect 35334 25531 35368 25569
rect 35666 25531 35702 25569
rect 35334 25494 35368 25497
rect 35666 25494 35702 25497
rect 35334 25491 35702 25494
rect 35922 25606 36290 25609
rect 35922 25603 35956 25606
rect 36254 25603 36290 25606
rect 35922 25531 35956 25569
rect 36254 25531 36290 25569
rect 35922 25494 35956 25497
rect 36254 25494 36290 25497
rect 35922 25491 36290 25494
rect 36510 25606 36878 25609
rect 36510 25603 36544 25606
rect 36842 25603 36878 25606
rect 36510 25531 36544 25569
rect 36842 25531 36878 25569
rect 36510 25494 36544 25497
rect 36842 25494 36878 25497
rect 36510 25491 36878 25494
rect 37098 25606 37466 25609
rect 37098 25603 37132 25606
rect 37430 25603 37466 25606
rect 37098 25531 37132 25569
rect 37430 25531 37466 25569
rect 37098 25494 37132 25497
rect 37430 25494 37466 25497
rect 37098 25491 37466 25494
rect 37686 25606 38054 25609
rect 37686 25603 37720 25606
rect 38018 25603 38054 25606
rect 37686 25531 37720 25569
rect 38018 25531 38054 25569
rect 37686 25494 37720 25497
rect 38018 25494 38054 25497
rect 37686 25491 38054 25494
rect 38274 25606 38642 25609
rect 38274 25603 38308 25606
rect 38606 25603 38642 25606
rect 38274 25531 38308 25569
rect 38606 25531 38642 25569
rect 38274 25494 38308 25497
rect 38606 25494 38642 25497
rect 38274 25491 38642 25494
rect 6795 25312 6845 25324
rect 6795 24932 6801 25312
rect 6784 24915 6801 24932
rect 6839 24932 6845 25312
rect 6839 24915 6856 24932
rect 3536 11952 3546 13186
rect 5048 11952 5058 13186
rect 6784 4988 6856 24915
rect 10648 24560 10658 24612
rect 10988 24560 10998 24612
rect 11236 24609 11246 24612
rect 11214 24603 11246 24609
rect 11576 24609 11586 24612
rect 11824 24609 11834 24612
rect 11576 24603 11594 24609
rect 11214 24569 11226 24603
rect 11214 24563 11246 24569
rect 11236 24560 11246 24563
rect 11576 24563 11594 24569
rect 11802 24603 11834 24609
rect 12164 24609 12174 24612
rect 12412 24609 12422 24612
rect 12164 24603 12182 24609
rect 11802 24569 11814 24603
rect 11802 24563 11834 24569
rect 11576 24560 11586 24563
rect 11824 24560 11834 24563
rect 12164 24563 12182 24569
rect 12390 24603 12422 24609
rect 12752 24609 12762 24612
rect 13000 24609 13010 24612
rect 12752 24603 12770 24609
rect 12390 24569 12402 24603
rect 12390 24563 12422 24569
rect 12164 24560 12174 24563
rect 12412 24560 12422 24563
rect 12752 24563 12770 24569
rect 12978 24603 13010 24609
rect 13340 24609 13350 24612
rect 13588 24609 13598 24612
rect 13340 24603 13358 24609
rect 12978 24569 12990 24603
rect 12978 24563 13010 24569
rect 12752 24560 12762 24563
rect 13000 24560 13010 24563
rect 13340 24563 13358 24569
rect 13566 24603 13598 24609
rect 13928 24609 13938 24612
rect 14176 24609 14186 24612
rect 13928 24603 13946 24609
rect 13566 24569 13578 24603
rect 13566 24563 13598 24569
rect 13340 24560 13350 24563
rect 13588 24560 13598 24563
rect 13928 24563 13946 24569
rect 14154 24603 14186 24609
rect 14516 24609 14526 24612
rect 14764 24609 14774 24612
rect 14516 24603 14534 24609
rect 14154 24569 14166 24603
rect 14154 24563 14186 24569
rect 13928 24560 13938 24563
rect 14176 24560 14186 24563
rect 14516 24563 14534 24569
rect 14742 24603 14774 24609
rect 15104 24609 15114 24612
rect 15352 24609 15362 24612
rect 15104 24603 15122 24609
rect 14742 24569 14754 24603
rect 14742 24563 14774 24569
rect 14516 24560 14526 24563
rect 14764 24560 14774 24563
rect 15104 24563 15122 24569
rect 15330 24603 15362 24609
rect 15692 24609 15702 24612
rect 15940 24609 15950 24612
rect 15692 24603 15710 24609
rect 15330 24569 15342 24603
rect 15330 24563 15362 24569
rect 15104 24560 15114 24563
rect 15352 24560 15362 24563
rect 15692 24563 15710 24569
rect 15918 24603 15950 24609
rect 16280 24609 16290 24612
rect 16528 24609 16538 24612
rect 16280 24603 16298 24609
rect 15918 24569 15930 24603
rect 15918 24563 15950 24569
rect 15692 24560 15702 24563
rect 15940 24560 15950 24563
rect 16280 24563 16298 24569
rect 16506 24603 16538 24609
rect 16868 24609 16878 24612
rect 17116 24609 17126 24612
rect 16868 24603 16886 24609
rect 16506 24569 16518 24603
rect 16506 24563 16538 24569
rect 16280 24560 16290 24563
rect 16528 24560 16538 24563
rect 16868 24563 16886 24569
rect 17094 24603 17126 24609
rect 17456 24609 17466 24612
rect 17704 24609 17714 24612
rect 17456 24603 17474 24609
rect 17094 24569 17106 24603
rect 17094 24563 17126 24569
rect 16868 24560 16878 24563
rect 17116 24560 17126 24563
rect 17456 24563 17474 24569
rect 17682 24603 17714 24609
rect 18044 24609 18054 24612
rect 18292 24609 18302 24612
rect 18044 24603 18062 24609
rect 17682 24569 17694 24603
rect 17682 24563 17714 24569
rect 17456 24560 17466 24563
rect 17704 24560 17714 24563
rect 18044 24563 18062 24569
rect 18270 24603 18302 24609
rect 18632 24609 18642 24612
rect 18880 24609 18890 24612
rect 18632 24603 18650 24609
rect 18270 24569 18282 24603
rect 18270 24563 18302 24569
rect 18044 24560 18054 24563
rect 18292 24560 18302 24563
rect 18632 24563 18650 24569
rect 18858 24603 18890 24609
rect 19220 24609 19230 24612
rect 19468 24609 19478 24612
rect 19220 24603 19238 24609
rect 18858 24569 18870 24603
rect 18858 24563 18890 24569
rect 18632 24560 18642 24563
rect 18880 24560 18890 24563
rect 19220 24563 19238 24569
rect 19446 24603 19478 24609
rect 19808 24609 19818 24612
rect 20056 24609 20066 24612
rect 19808 24603 19826 24609
rect 19446 24569 19458 24603
rect 19446 24563 19478 24569
rect 19220 24560 19230 24563
rect 19468 24560 19478 24563
rect 19808 24563 19826 24569
rect 20034 24603 20066 24609
rect 20396 24609 20406 24612
rect 20644 24609 20654 24612
rect 20396 24603 20414 24609
rect 20034 24569 20046 24603
rect 20034 24563 20066 24569
rect 19808 24560 19818 24563
rect 20056 24560 20066 24563
rect 20396 24563 20414 24569
rect 20622 24603 20654 24609
rect 20984 24609 20994 24612
rect 21232 24609 21242 24612
rect 20984 24603 21002 24609
rect 20622 24569 20634 24603
rect 20622 24563 20654 24569
rect 20396 24560 20406 24563
rect 20644 24560 20654 24563
rect 20984 24563 21002 24569
rect 21210 24603 21242 24609
rect 21572 24609 21582 24612
rect 21820 24609 21830 24612
rect 21572 24603 21590 24609
rect 21210 24569 21222 24603
rect 21210 24563 21242 24569
rect 20984 24560 20994 24563
rect 21232 24560 21242 24563
rect 21572 24563 21590 24569
rect 21798 24603 21830 24609
rect 22160 24609 22170 24612
rect 22160 24603 22178 24609
rect 21798 24569 21810 24603
rect 21798 24563 21830 24569
rect 21572 24560 21582 24563
rect 21820 24560 21830 24563
rect 22160 24563 22178 24569
rect 22160 24560 22170 24563
rect 22406 24554 22416 24622
rect 22736 24554 22746 24622
rect 22994 24609 23004 24622
rect 22986 24603 23004 24609
rect 23324 24609 23334 24622
rect 23582 24609 23592 24622
rect 23324 24603 23354 24609
rect 22986 24563 23004 24569
rect 22994 24554 23004 24563
rect 23324 24563 23354 24569
rect 23574 24603 23592 24609
rect 23912 24609 23922 24622
rect 24170 24609 24180 24622
rect 23912 24603 23942 24609
rect 23574 24563 23592 24569
rect 23324 24554 23334 24563
rect 23582 24554 23592 24563
rect 23912 24563 23942 24569
rect 24162 24603 24180 24609
rect 24500 24609 24510 24622
rect 24758 24609 24768 24622
rect 24500 24603 24530 24609
rect 24162 24563 24180 24569
rect 23912 24554 23922 24563
rect 24170 24554 24180 24563
rect 24500 24563 24530 24569
rect 24750 24603 24768 24609
rect 25088 24609 25098 24622
rect 25346 24609 25356 24622
rect 25088 24603 25118 24609
rect 24750 24563 24768 24569
rect 24500 24554 24510 24563
rect 24758 24554 24768 24563
rect 25088 24563 25118 24569
rect 25338 24603 25356 24609
rect 25676 24609 25686 24622
rect 25934 24609 25944 24622
rect 25676 24603 25706 24609
rect 25338 24563 25356 24569
rect 25088 24554 25098 24563
rect 25346 24554 25356 24563
rect 25676 24563 25706 24569
rect 25926 24603 25944 24609
rect 26264 24609 26274 24622
rect 26522 24609 26532 24622
rect 26264 24603 26294 24609
rect 25926 24563 25944 24569
rect 25676 24554 25686 24563
rect 25934 24554 25944 24563
rect 26264 24563 26294 24569
rect 26514 24603 26532 24609
rect 26852 24609 26862 24622
rect 27110 24609 27120 24622
rect 26852 24603 26882 24609
rect 26514 24563 26532 24569
rect 26264 24554 26274 24563
rect 26522 24554 26532 24563
rect 26852 24563 26882 24569
rect 27102 24603 27120 24609
rect 27440 24609 27450 24622
rect 27698 24609 27708 24622
rect 27440 24603 27470 24609
rect 27102 24563 27120 24569
rect 26852 24554 26862 24563
rect 27110 24554 27120 24563
rect 27440 24563 27470 24569
rect 27690 24603 27708 24609
rect 28028 24609 28038 24622
rect 28286 24609 28296 24622
rect 28028 24603 28058 24609
rect 27690 24563 27708 24569
rect 27440 24554 27450 24563
rect 27698 24554 27708 24563
rect 28028 24563 28058 24569
rect 28278 24603 28296 24609
rect 28616 24609 28626 24622
rect 28874 24609 28884 24622
rect 28616 24603 28646 24609
rect 28278 24563 28296 24569
rect 28028 24554 28038 24563
rect 28286 24554 28296 24563
rect 28616 24563 28646 24569
rect 28866 24603 28884 24609
rect 29204 24609 29214 24622
rect 29462 24609 29472 24622
rect 29204 24603 29234 24609
rect 28866 24563 28884 24569
rect 28616 24554 28626 24563
rect 28874 24554 28884 24563
rect 29204 24563 29234 24569
rect 29454 24603 29472 24609
rect 29792 24609 29802 24622
rect 30050 24609 30060 24622
rect 29792 24603 29822 24609
rect 29454 24563 29472 24569
rect 29204 24554 29214 24563
rect 29462 24554 29472 24563
rect 29792 24563 29822 24569
rect 30042 24603 30060 24609
rect 30380 24609 30390 24622
rect 30638 24609 30648 24622
rect 30380 24603 30410 24609
rect 30042 24563 30060 24569
rect 29792 24554 29802 24563
rect 30050 24554 30060 24563
rect 30380 24563 30410 24569
rect 30630 24603 30648 24609
rect 30968 24609 30978 24622
rect 31226 24609 31236 24622
rect 30968 24603 30998 24609
rect 30630 24563 30648 24569
rect 30380 24554 30390 24563
rect 30638 24554 30648 24563
rect 30968 24563 30998 24569
rect 31218 24603 31236 24609
rect 31556 24609 31566 24622
rect 31814 24609 31824 24622
rect 31556 24603 31586 24609
rect 31218 24563 31236 24569
rect 30968 24554 30978 24563
rect 31226 24554 31236 24563
rect 31556 24563 31586 24569
rect 31806 24603 31824 24609
rect 32144 24609 32154 24622
rect 32402 24609 32412 24622
rect 32144 24603 32174 24609
rect 31806 24563 31824 24569
rect 31556 24554 31566 24563
rect 31814 24554 31824 24563
rect 32144 24563 32174 24569
rect 32394 24603 32412 24609
rect 32732 24609 32742 24622
rect 32990 24609 33000 24622
rect 32732 24603 32762 24609
rect 32394 24563 32412 24569
rect 32144 24554 32154 24563
rect 32402 24554 32412 24563
rect 32732 24563 32762 24569
rect 32982 24603 33000 24609
rect 33320 24609 33330 24622
rect 33578 24609 33588 24622
rect 33320 24603 33350 24609
rect 32982 24563 33000 24569
rect 32732 24554 32742 24563
rect 32990 24554 33000 24563
rect 33320 24563 33350 24569
rect 33570 24603 33588 24609
rect 33908 24609 33918 24622
rect 34166 24609 34176 24622
rect 33908 24603 33938 24609
rect 33570 24563 33588 24569
rect 33320 24554 33330 24563
rect 33578 24554 33588 24563
rect 33908 24563 33938 24569
rect 34158 24603 34176 24609
rect 34496 24609 34506 24622
rect 34754 24609 34764 24622
rect 34496 24603 34526 24609
rect 34158 24563 34176 24569
rect 33908 24554 33918 24563
rect 34166 24554 34176 24563
rect 34496 24563 34526 24569
rect 34746 24603 34764 24609
rect 35084 24609 35094 24622
rect 35342 24609 35352 24622
rect 35084 24603 35114 24609
rect 34746 24563 34764 24569
rect 34496 24554 34506 24563
rect 34754 24554 34764 24563
rect 35084 24563 35114 24569
rect 35334 24603 35352 24609
rect 35672 24609 35682 24622
rect 35930 24609 35940 24622
rect 35672 24603 35702 24609
rect 35334 24563 35352 24569
rect 35084 24554 35094 24563
rect 35342 24554 35352 24563
rect 35672 24563 35702 24569
rect 35922 24603 35940 24609
rect 36260 24609 36270 24622
rect 36518 24609 36528 24622
rect 36260 24603 36290 24609
rect 35922 24563 35940 24569
rect 35672 24554 35682 24563
rect 35930 24554 35940 24563
rect 36260 24563 36290 24569
rect 36510 24603 36528 24609
rect 36848 24609 36858 24622
rect 37106 24609 37116 24622
rect 36848 24603 36878 24609
rect 36510 24563 36528 24569
rect 36260 24554 36270 24563
rect 36518 24554 36528 24563
rect 36848 24563 36878 24569
rect 37098 24603 37116 24609
rect 37436 24609 37446 24622
rect 37694 24609 37704 24622
rect 37436 24603 37466 24609
rect 37098 24563 37116 24569
rect 36848 24554 36858 24563
rect 37106 24554 37116 24563
rect 37436 24563 37466 24569
rect 37686 24603 37704 24609
rect 38024 24609 38034 24622
rect 38282 24609 38292 24622
rect 38024 24603 38054 24609
rect 37686 24563 37704 24569
rect 37436 24554 37446 24563
rect 37694 24554 37704 24563
rect 38024 24563 38054 24569
rect 38274 24603 38292 24609
rect 38612 24609 38622 24622
rect 38612 24603 38642 24609
rect 38274 24563 38292 24569
rect 38024 24554 38034 24563
rect 38282 24554 38292 24563
rect 38612 24563 38642 24569
rect 38612 24554 38622 24563
rect 39799 24442 39849 24454
rect 39799 24074 39805 24442
rect 39788 24045 39805 24074
rect 39843 24074 39849 24442
rect 39843 24045 39860 24074
rect 38654 24038 38990 24044
rect 38654 23772 38666 24038
rect 38978 23772 38990 24038
rect 38654 23766 38990 23772
rect 38666 22382 38854 23766
rect 39788 23424 39860 24045
rect 39572 22924 39582 23424
rect 39860 22924 39870 23424
rect 39788 22661 39860 22924
rect 39788 22656 39805 22661
rect 37826 22370 38986 22382
rect 37822 20906 37832 22370
rect 38980 20906 38990 22370
rect 39799 22264 39805 22656
rect 39843 22656 39860 22661
rect 39843 22264 39849 22656
rect 39799 22252 39849 22264
rect 39799 21430 39849 21442
rect 39799 21033 39805 21430
rect 39843 21033 39849 21430
rect 39799 21032 39849 21033
rect 37826 20894 38986 20906
rect 10472 12046 10482 12856
rect 11158 12850 11168 12856
rect 39788 12850 39860 21032
rect 44302 18676 44312 19484
rect 45378 18676 45388 19484
rect 12288 12046 12298 12850
rect 38794 12252 39860 12850
rect 10640 11144 10650 11196
rect 10994 11144 11004 11196
rect 11228 11193 11238 11196
rect 11226 11187 11238 11193
rect 11582 11193 11592 11196
rect 11816 11193 11826 11196
rect 11582 11187 11594 11193
rect 11226 11147 11238 11153
rect 11228 11144 11238 11147
rect 11582 11147 11594 11153
rect 11814 11187 11826 11193
rect 12170 11193 12180 11196
rect 12404 11193 12414 11196
rect 12170 11187 12182 11193
rect 11814 11147 11826 11153
rect 11582 11144 11592 11147
rect 11816 11144 11826 11147
rect 12170 11147 12182 11153
rect 12402 11187 12414 11193
rect 12758 11193 12768 11196
rect 12992 11193 13002 11196
rect 12758 11187 12770 11193
rect 12402 11147 12414 11153
rect 12170 11144 12180 11147
rect 12404 11144 12414 11147
rect 12758 11147 12770 11153
rect 12990 11187 13002 11193
rect 13346 11193 13356 11196
rect 13580 11193 13590 11196
rect 13346 11187 13358 11193
rect 12990 11147 13002 11153
rect 12758 11144 12768 11147
rect 12992 11144 13002 11147
rect 13346 11147 13358 11153
rect 13578 11187 13590 11193
rect 13934 11193 13944 11196
rect 14168 11193 14178 11196
rect 13934 11187 13946 11193
rect 13578 11147 13590 11153
rect 13346 11144 13356 11147
rect 13580 11144 13590 11147
rect 13934 11147 13946 11153
rect 14166 11187 14178 11193
rect 14522 11193 14532 11196
rect 14756 11193 14766 11196
rect 14522 11187 14534 11193
rect 14166 11147 14178 11153
rect 13934 11144 13944 11147
rect 14168 11144 14178 11147
rect 14522 11147 14534 11153
rect 14754 11187 14766 11193
rect 15110 11193 15120 11196
rect 15344 11193 15354 11196
rect 15110 11187 15122 11193
rect 14754 11147 14766 11153
rect 14522 11144 14532 11147
rect 14756 11144 14766 11147
rect 15110 11147 15122 11153
rect 15342 11187 15354 11193
rect 15698 11193 15708 11196
rect 15932 11193 15942 11196
rect 15698 11187 15710 11193
rect 15342 11147 15354 11153
rect 15110 11144 15120 11147
rect 15344 11144 15354 11147
rect 15698 11147 15710 11153
rect 15930 11187 15942 11193
rect 16286 11193 16296 11196
rect 16520 11193 16530 11196
rect 16286 11187 16298 11193
rect 15930 11147 15942 11153
rect 15698 11144 15708 11147
rect 15932 11144 15942 11147
rect 16286 11147 16298 11153
rect 16518 11187 16530 11193
rect 16874 11193 16884 11196
rect 17108 11193 17118 11196
rect 16874 11187 16886 11193
rect 16518 11147 16530 11153
rect 16286 11144 16296 11147
rect 16520 11144 16530 11147
rect 16874 11147 16886 11153
rect 17106 11187 17118 11193
rect 17462 11193 17472 11196
rect 17696 11193 17706 11196
rect 17462 11187 17474 11193
rect 17106 11147 17118 11153
rect 16874 11144 16884 11147
rect 17108 11144 17118 11147
rect 17462 11147 17474 11153
rect 17694 11187 17706 11193
rect 18050 11193 18060 11196
rect 18284 11193 18294 11196
rect 18050 11187 18062 11193
rect 17694 11147 17706 11153
rect 17462 11144 17472 11147
rect 17696 11144 17706 11147
rect 18050 11147 18062 11153
rect 18282 11187 18294 11193
rect 18638 11193 18648 11196
rect 18872 11193 18882 11196
rect 18638 11187 18650 11193
rect 18282 11147 18294 11153
rect 18050 11144 18060 11147
rect 18284 11144 18294 11147
rect 18638 11147 18650 11153
rect 18870 11187 18882 11193
rect 19226 11193 19236 11196
rect 19460 11193 19470 11196
rect 19226 11187 19238 11193
rect 18870 11147 18882 11153
rect 18638 11144 18648 11147
rect 18872 11144 18882 11147
rect 19226 11147 19238 11153
rect 19458 11187 19470 11193
rect 19814 11193 19824 11196
rect 20048 11193 20058 11196
rect 19814 11187 19826 11193
rect 19458 11147 19470 11153
rect 19226 11144 19236 11147
rect 19460 11144 19470 11147
rect 19814 11147 19826 11153
rect 20046 11187 20058 11193
rect 20402 11193 20412 11196
rect 20636 11193 20646 11196
rect 20402 11187 20414 11193
rect 20046 11147 20058 11153
rect 19814 11144 19824 11147
rect 20048 11144 20058 11147
rect 20402 11147 20414 11153
rect 20634 11187 20646 11193
rect 20990 11193 21000 11196
rect 21224 11193 21234 11196
rect 20990 11187 21002 11193
rect 20634 11147 20646 11153
rect 20402 11144 20412 11147
rect 20636 11144 20646 11147
rect 20990 11147 21002 11153
rect 21222 11187 21234 11193
rect 21578 11193 21588 11196
rect 21812 11193 21822 11196
rect 21578 11187 21590 11193
rect 21222 11147 21234 11153
rect 20990 11144 21000 11147
rect 21224 11144 21234 11147
rect 21578 11147 21590 11153
rect 21810 11187 21822 11193
rect 22166 11193 22176 11196
rect 22166 11187 22178 11193
rect 21810 11147 21822 11153
rect 21578 11144 21588 11147
rect 21812 11144 21822 11147
rect 22166 11147 22178 11153
rect 22166 11144 22176 11147
rect 22436 11138 22446 11196
rect 22716 11138 22726 11196
rect 23010 11140 23020 11200
rect 23318 11140 23328 11200
rect 23590 11136 23600 11200
rect 23920 11136 23930 11200
rect 24168 11130 24178 11202
rect 24512 11130 24522 11202
rect 24766 11130 24776 11212
rect 25094 11130 25104 11212
rect 25350 11128 25360 11230
rect 25698 11128 25708 11230
rect 25934 11126 25944 11228
rect 26282 11126 26292 11228
rect 26522 11193 26532 11228
rect 26502 11187 26532 11193
rect 26870 11193 26880 11228
rect 27110 11193 27120 11228
rect 26870 11187 26894 11193
rect 26502 11153 26514 11187
rect 26882 11153 26894 11187
rect 26502 11147 26532 11153
rect 26522 11126 26532 11147
rect 26870 11147 26894 11153
rect 27090 11187 27120 11193
rect 27458 11193 27468 11228
rect 27698 11193 27708 11228
rect 27458 11187 27482 11193
rect 27090 11153 27102 11187
rect 27470 11153 27482 11187
rect 27090 11147 27120 11153
rect 26870 11126 26880 11147
rect 27110 11126 27120 11147
rect 27458 11147 27482 11153
rect 27678 11187 27708 11193
rect 28046 11193 28056 11228
rect 28286 11193 28296 11228
rect 28046 11187 28070 11193
rect 27678 11153 27690 11187
rect 28058 11153 28070 11187
rect 27678 11147 27708 11153
rect 27458 11126 27468 11147
rect 27698 11126 27708 11147
rect 28046 11147 28070 11153
rect 28266 11187 28296 11193
rect 28634 11193 28644 11228
rect 28874 11193 28884 11228
rect 28634 11187 28658 11193
rect 28266 11153 28278 11187
rect 28646 11153 28658 11187
rect 28266 11147 28296 11153
rect 28046 11126 28056 11147
rect 28286 11126 28296 11147
rect 28634 11147 28658 11153
rect 28854 11187 28884 11193
rect 29222 11193 29232 11228
rect 29462 11193 29472 11228
rect 29222 11187 29246 11193
rect 28854 11153 28866 11187
rect 29234 11153 29246 11187
rect 28854 11147 28884 11153
rect 28634 11126 28644 11147
rect 28874 11126 28884 11147
rect 29222 11147 29246 11153
rect 29442 11187 29472 11193
rect 29810 11193 29820 11228
rect 30050 11193 30060 11228
rect 29810 11187 29834 11193
rect 29442 11153 29454 11187
rect 29822 11153 29834 11187
rect 29442 11147 29472 11153
rect 29222 11126 29232 11147
rect 29462 11126 29472 11147
rect 29810 11147 29834 11153
rect 30030 11187 30060 11193
rect 30398 11193 30408 11228
rect 30638 11193 30648 11228
rect 30398 11187 30422 11193
rect 30030 11153 30042 11187
rect 30410 11153 30422 11187
rect 30030 11147 30060 11153
rect 29810 11126 29820 11147
rect 30050 11126 30060 11147
rect 30398 11147 30422 11153
rect 30618 11187 30648 11193
rect 30986 11193 30996 11228
rect 31226 11193 31236 11228
rect 30986 11187 31010 11193
rect 30618 11153 30630 11187
rect 30998 11153 31010 11187
rect 30618 11147 30648 11153
rect 30398 11126 30408 11147
rect 30638 11126 30648 11147
rect 30986 11147 31010 11153
rect 31206 11187 31236 11193
rect 31574 11193 31584 11228
rect 31814 11193 31824 11228
rect 31574 11187 31598 11193
rect 31206 11153 31218 11187
rect 31586 11153 31598 11187
rect 31206 11147 31236 11153
rect 30986 11126 30996 11147
rect 31226 11126 31236 11147
rect 31574 11147 31598 11153
rect 31794 11187 31824 11193
rect 32162 11193 32172 11228
rect 32402 11193 32412 11228
rect 32162 11187 32186 11193
rect 31794 11153 31806 11187
rect 32174 11153 32186 11187
rect 31794 11147 31824 11153
rect 31574 11126 31584 11147
rect 31814 11126 31824 11147
rect 32162 11147 32186 11153
rect 32382 11187 32412 11193
rect 32750 11193 32760 11228
rect 32990 11193 33000 11228
rect 32750 11187 32774 11193
rect 32382 11153 32394 11187
rect 32762 11153 32774 11187
rect 32382 11147 32412 11153
rect 32162 11126 32172 11147
rect 32402 11126 32412 11147
rect 32750 11147 32774 11153
rect 32970 11187 33000 11193
rect 33338 11193 33348 11228
rect 33578 11193 33588 11228
rect 33338 11187 33362 11193
rect 32970 11153 32982 11187
rect 33350 11153 33362 11187
rect 32970 11147 33000 11153
rect 32750 11126 32760 11147
rect 32990 11126 33000 11147
rect 33338 11147 33362 11153
rect 33558 11187 33588 11193
rect 33926 11193 33936 11228
rect 34166 11193 34176 11228
rect 33926 11187 33950 11193
rect 33558 11153 33570 11187
rect 33938 11153 33950 11187
rect 33558 11147 33588 11153
rect 33338 11126 33348 11147
rect 33578 11126 33588 11147
rect 33926 11147 33950 11153
rect 34146 11187 34176 11193
rect 34514 11193 34524 11228
rect 34754 11193 34764 11228
rect 34514 11187 34538 11193
rect 34146 11153 34158 11187
rect 34526 11153 34538 11187
rect 34146 11147 34176 11153
rect 33926 11126 33936 11147
rect 34166 11126 34176 11147
rect 34514 11147 34538 11153
rect 34734 11187 34764 11193
rect 35102 11193 35112 11228
rect 35342 11193 35352 11228
rect 35102 11187 35126 11193
rect 34734 11153 34746 11187
rect 35114 11153 35126 11187
rect 34734 11147 34764 11153
rect 34514 11126 34524 11147
rect 34754 11126 34764 11147
rect 35102 11147 35126 11153
rect 35322 11187 35352 11193
rect 35690 11193 35700 11228
rect 35930 11193 35940 11228
rect 35690 11187 35714 11193
rect 35322 11153 35334 11187
rect 35702 11153 35714 11187
rect 35322 11147 35352 11153
rect 35102 11126 35112 11147
rect 35342 11126 35352 11147
rect 35690 11147 35714 11153
rect 35910 11187 35940 11193
rect 36278 11193 36288 11228
rect 36518 11193 36528 11228
rect 36278 11187 36302 11193
rect 35910 11153 35922 11187
rect 36290 11153 36302 11187
rect 35910 11147 35940 11153
rect 35690 11126 35700 11147
rect 35930 11126 35940 11147
rect 36278 11147 36302 11153
rect 36498 11187 36528 11193
rect 36866 11193 36876 11228
rect 37106 11193 37116 11228
rect 36866 11187 36890 11193
rect 36498 11153 36510 11187
rect 36878 11153 36890 11187
rect 36498 11147 36528 11153
rect 36278 11126 36288 11147
rect 36518 11126 36528 11147
rect 36866 11147 36890 11153
rect 37086 11187 37116 11193
rect 37454 11193 37464 11228
rect 37694 11193 37704 11228
rect 37454 11187 37478 11193
rect 37086 11153 37098 11187
rect 37466 11153 37478 11187
rect 37086 11147 37116 11153
rect 36866 11126 36876 11147
rect 37106 11126 37116 11147
rect 37454 11147 37478 11153
rect 37674 11187 37704 11193
rect 38042 11193 38052 11228
rect 38282 11193 38292 11228
rect 38042 11187 38066 11193
rect 37674 11153 37686 11187
rect 38054 11153 38066 11187
rect 37674 11147 37704 11153
rect 37454 11126 37464 11147
rect 37694 11126 37704 11147
rect 38042 11147 38066 11153
rect 38262 11187 38292 11193
rect 38630 11193 38640 11228
rect 38630 11187 38654 11193
rect 38262 11153 38274 11187
rect 38642 11153 38654 11187
rect 38262 11147 38292 11153
rect 38042 11126 38052 11147
rect 38282 11126 38292 11147
rect 38630 11147 38654 11153
rect 38630 11126 38640 11147
rect 10650 10148 10660 10266
rect 10982 10148 10992 10266
rect 11238 10265 11248 10266
rect 11214 10259 11248 10265
rect 11570 10265 11580 10266
rect 11826 10265 11836 10266
rect 11570 10259 11606 10265
rect 11214 10225 11226 10259
rect 11594 10225 11606 10259
rect 11214 10187 11248 10225
rect 11570 10187 11606 10225
rect 11214 10153 11226 10187
rect 11594 10153 11606 10187
rect 11214 10148 11248 10153
rect 11570 10148 11606 10153
rect 11214 10147 11606 10148
rect 11802 10259 11836 10265
rect 12158 10265 12168 10266
rect 12414 10265 12424 10266
rect 12158 10259 12194 10265
rect 11802 10225 11814 10259
rect 12182 10225 12194 10259
rect 11802 10187 11836 10225
rect 12158 10187 12194 10225
rect 11802 10153 11814 10187
rect 12182 10153 12194 10187
rect 11802 10148 11836 10153
rect 12158 10148 12194 10153
rect 11802 10147 12194 10148
rect 12390 10259 12424 10265
rect 12746 10265 12756 10266
rect 13002 10265 13012 10266
rect 12746 10259 12782 10265
rect 12390 10225 12402 10259
rect 12770 10225 12782 10259
rect 12390 10187 12424 10225
rect 12746 10187 12782 10225
rect 12390 10153 12402 10187
rect 12770 10153 12782 10187
rect 12390 10148 12424 10153
rect 12746 10148 12782 10153
rect 12390 10147 12782 10148
rect 12978 10259 13012 10265
rect 13334 10265 13344 10266
rect 13590 10265 13600 10266
rect 13334 10259 13370 10265
rect 12978 10225 12990 10259
rect 13358 10225 13370 10259
rect 12978 10187 13012 10225
rect 13334 10187 13370 10225
rect 12978 10153 12990 10187
rect 13358 10153 13370 10187
rect 12978 10148 13012 10153
rect 13334 10148 13370 10153
rect 12978 10147 13370 10148
rect 13566 10259 13600 10265
rect 13922 10265 13932 10266
rect 14178 10265 14188 10266
rect 13922 10259 13958 10265
rect 13566 10225 13578 10259
rect 13946 10225 13958 10259
rect 13566 10187 13600 10225
rect 13922 10187 13958 10225
rect 13566 10153 13578 10187
rect 13946 10153 13958 10187
rect 13566 10148 13600 10153
rect 13922 10148 13958 10153
rect 13566 10147 13958 10148
rect 14154 10259 14188 10265
rect 14510 10265 14520 10266
rect 14766 10265 14776 10266
rect 14510 10259 14546 10265
rect 14154 10225 14166 10259
rect 14534 10225 14546 10259
rect 14154 10187 14188 10225
rect 14510 10187 14546 10225
rect 14154 10153 14166 10187
rect 14534 10153 14546 10187
rect 14154 10148 14188 10153
rect 14510 10148 14546 10153
rect 14154 10147 14546 10148
rect 14742 10259 14776 10265
rect 15098 10265 15108 10266
rect 15354 10265 15364 10266
rect 15098 10259 15134 10265
rect 14742 10225 14754 10259
rect 15122 10225 15134 10259
rect 14742 10187 14776 10225
rect 15098 10187 15134 10225
rect 14742 10153 14754 10187
rect 15122 10153 15134 10187
rect 14742 10148 14776 10153
rect 15098 10148 15134 10153
rect 14742 10147 15134 10148
rect 15330 10259 15364 10265
rect 15686 10265 15696 10266
rect 15942 10265 15952 10266
rect 15686 10259 15722 10265
rect 15330 10225 15342 10259
rect 15710 10225 15722 10259
rect 15330 10187 15364 10225
rect 15686 10187 15722 10225
rect 15330 10153 15342 10187
rect 15710 10153 15722 10187
rect 15330 10148 15364 10153
rect 15686 10148 15722 10153
rect 15330 10147 15722 10148
rect 15918 10259 15952 10265
rect 16274 10265 16284 10266
rect 16530 10265 16540 10266
rect 16274 10259 16310 10265
rect 15918 10225 15930 10259
rect 16298 10225 16310 10259
rect 15918 10187 15952 10225
rect 16274 10187 16310 10225
rect 15918 10153 15930 10187
rect 16298 10153 16310 10187
rect 15918 10148 15952 10153
rect 16274 10148 16310 10153
rect 15918 10147 16310 10148
rect 16506 10259 16540 10265
rect 16862 10265 16872 10266
rect 17118 10265 17128 10266
rect 16862 10259 16898 10265
rect 16506 10225 16518 10259
rect 16886 10225 16898 10259
rect 16506 10187 16540 10225
rect 16862 10187 16898 10225
rect 16506 10153 16518 10187
rect 16886 10153 16898 10187
rect 16506 10148 16540 10153
rect 16862 10148 16898 10153
rect 16506 10147 16898 10148
rect 17094 10259 17128 10265
rect 17450 10265 17460 10266
rect 17706 10265 17716 10266
rect 17450 10259 17486 10265
rect 17094 10225 17106 10259
rect 17474 10225 17486 10259
rect 17094 10187 17128 10225
rect 17450 10187 17486 10225
rect 17094 10153 17106 10187
rect 17474 10153 17486 10187
rect 17094 10148 17128 10153
rect 17450 10148 17486 10153
rect 17094 10147 17486 10148
rect 17682 10259 17716 10265
rect 18038 10265 18048 10266
rect 18294 10265 18304 10266
rect 18038 10259 18074 10265
rect 17682 10225 17694 10259
rect 18062 10225 18074 10259
rect 17682 10187 17716 10225
rect 18038 10187 18074 10225
rect 17682 10153 17694 10187
rect 18062 10153 18074 10187
rect 17682 10148 17716 10153
rect 18038 10148 18074 10153
rect 17682 10147 18074 10148
rect 18270 10259 18304 10265
rect 18626 10265 18636 10266
rect 18882 10265 18892 10266
rect 18626 10259 18662 10265
rect 18270 10225 18282 10259
rect 18650 10225 18662 10259
rect 18270 10187 18304 10225
rect 18626 10187 18662 10225
rect 18270 10153 18282 10187
rect 18650 10153 18662 10187
rect 18270 10148 18304 10153
rect 18626 10148 18662 10153
rect 18270 10147 18662 10148
rect 18858 10259 18892 10265
rect 19214 10265 19224 10266
rect 19470 10265 19480 10266
rect 19214 10259 19250 10265
rect 18858 10225 18870 10259
rect 19238 10225 19250 10259
rect 18858 10187 18892 10225
rect 19214 10187 19250 10225
rect 18858 10153 18870 10187
rect 19238 10153 19250 10187
rect 18858 10148 18892 10153
rect 19214 10148 19250 10153
rect 18858 10147 19250 10148
rect 19446 10259 19480 10265
rect 19802 10265 19812 10266
rect 20058 10265 20068 10266
rect 19802 10259 19838 10265
rect 19446 10225 19458 10259
rect 19826 10225 19838 10259
rect 19446 10187 19480 10225
rect 19802 10187 19838 10225
rect 19446 10153 19458 10187
rect 19826 10153 19838 10187
rect 19446 10148 19480 10153
rect 19802 10148 19838 10153
rect 19446 10147 19838 10148
rect 20034 10259 20068 10265
rect 20390 10265 20400 10266
rect 20646 10265 20656 10266
rect 20390 10259 20426 10265
rect 20034 10225 20046 10259
rect 20414 10225 20426 10259
rect 20034 10187 20068 10225
rect 20390 10187 20426 10225
rect 20034 10153 20046 10187
rect 20414 10153 20426 10187
rect 20034 10148 20068 10153
rect 20390 10148 20426 10153
rect 20034 10147 20426 10148
rect 20622 10259 20656 10265
rect 20978 10265 20988 10266
rect 21234 10265 21244 10266
rect 20978 10259 21014 10265
rect 20622 10225 20634 10259
rect 21002 10225 21014 10259
rect 20622 10187 20656 10225
rect 20978 10187 21014 10225
rect 20622 10153 20634 10187
rect 21002 10153 21014 10187
rect 20622 10148 20656 10153
rect 20978 10148 21014 10153
rect 20622 10147 21014 10148
rect 21210 10259 21244 10265
rect 21566 10265 21576 10266
rect 21822 10265 21832 10266
rect 21566 10259 21602 10265
rect 21210 10225 21222 10259
rect 21590 10225 21602 10259
rect 21210 10187 21244 10225
rect 21566 10187 21602 10225
rect 21210 10153 21222 10187
rect 21590 10153 21602 10187
rect 21210 10148 21244 10153
rect 21566 10148 21602 10153
rect 21210 10147 21602 10148
rect 21798 10259 21832 10265
rect 22154 10265 22164 10266
rect 22154 10259 22190 10265
rect 21798 10225 21810 10259
rect 22178 10225 22190 10259
rect 21798 10187 21832 10225
rect 22154 10187 22190 10225
rect 21798 10153 21810 10187
rect 22178 10153 22190 10187
rect 21798 10148 21832 10153
rect 22154 10148 22190 10153
rect 21798 10147 22190 10148
rect 22408 10146 22418 10266
rect 22752 10146 22762 10266
rect 22996 10265 23006 10266
rect 22974 10259 23006 10265
rect 23340 10265 23350 10266
rect 23584 10265 23594 10266
rect 23340 10259 23354 10265
rect 22974 10225 22986 10259
rect 22974 10187 23006 10225
rect 23340 10187 23354 10225
rect 22974 10153 22986 10187
rect 22974 10147 23006 10153
rect 22996 10146 23006 10147
rect 23340 10147 23354 10153
rect 23562 10259 23594 10265
rect 23928 10265 23938 10266
rect 24172 10265 24182 10266
rect 23928 10259 23942 10265
rect 23562 10225 23574 10259
rect 23562 10187 23594 10225
rect 23928 10187 23942 10225
rect 23562 10153 23574 10187
rect 23562 10147 23594 10153
rect 23340 10146 23350 10147
rect 23584 10146 23594 10147
rect 23928 10147 23942 10153
rect 24150 10259 24182 10265
rect 24516 10265 24526 10266
rect 24760 10265 24770 10266
rect 24516 10259 24530 10265
rect 24150 10225 24162 10259
rect 24150 10187 24182 10225
rect 24516 10187 24530 10225
rect 24150 10153 24162 10187
rect 24150 10147 24182 10153
rect 23928 10146 23938 10147
rect 24172 10146 24182 10147
rect 24516 10147 24530 10153
rect 24738 10259 24770 10265
rect 25104 10265 25114 10266
rect 25348 10265 25358 10266
rect 25104 10259 25118 10265
rect 24738 10225 24750 10259
rect 24738 10187 24770 10225
rect 25104 10187 25118 10225
rect 24738 10153 24750 10187
rect 24738 10147 24770 10153
rect 24516 10146 24526 10147
rect 24760 10146 24770 10147
rect 25104 10147 25118 10153
rect 25326 10259 25358 10265
rect 25692 10265 25702 10266
rect 25936 10265 25946 10266
rect 25692 10259 25706 10265
rect 25326 10225 25338 10259
rect 25326 10187 25358 10225
rect 25692 10187 25706 10225
rect 25326 10153 25338 10187
rect 25326 10147 25358 10153
rect 25104 10146 25114 10147
rect 25348 10146 25358 10147
rect 25692 10147 25706 10153
rect 25914 10259 25946 10265
rect 26280 10265 26290 10266
rect 26524 10265 26534 10266
rect 26280 10259 26294 10265
rect 25914 10225 25926 10259
rect 25914 10187 25946 10225
rect 26280 10187 26294 10225
rect 25914 10153 25926 10187
rect 25914 10147 25946 10153
rect 25692 10146 25702 10147
rect 25936 10146 25946 10147
rect 26280 10147 26294 10153
rect 26502 10259 26534 10265
rect 26868 10265 26878 10266
rect 27112 10265 27122 10266
rect 26868 10259 26882 10265
rect 26502 10225 26514 10259
rect 26502 10187 26534 10225
rect 26868 10187 26882 10225
rect 26502 10153 26514 10187
rect 26502 10147 26534 10153
rect 26280 10146 26290 10147
rect 26524 10146 26534 10147
rect 26868 10147 26882 10153
rect 27090 10259 27122 10265
rect 27456 10265 27466 10266
rect 27700 10265 27710 10266
rect 27456 10259 27470 10265
rect 27090 10225 27102 10259
rect 27090 10187 27122 10225
rect 27456 10187 27470 10225
rect 27090 10153 27102 10187
rect 27090 10147 27122 10153
rect 26868 10146 26878 10147
rect 27112 10146 27122 10147
rect 27456 10147 27470 10153
rect 27678 10259 27710 10265
rect 28044 10265 28054 10266
rect 28288 10265 28298 10266
rect 28044 10259 28058 10265
rect 27678 10225 27690 10259
rect 27678 10187 27710 10225
rect 28044 10187 28058 10225
rect 27678 10153 27690 10187
rect 27678 10147 27710 10153
rect 27456 10146 27466 10147
rect 27700 10146 27710 10147
rect 28044 10147 28058 10153
rect 28266 10259 28298 10265
rect 28632 10265 28642 10266
rect 28876 10265 28886 10266
rect 28632 10259 28646 10265
rect 28266 10225 28278 10259
rect 28266 10187 28298 10225
rect 28632 10187 28646 10225
rect 28266 10153 28278 10187
rect 28266 10147 28298 10153
rect 28044 10146 28054 10147
rect 28288 10146 28298 10147
rect 28632 10147 28646 10153
rect 28854 10259 28886 10265
rect 29220 10265 29230 10266
rect 29464 10265 29474 10266
rect 29220 10259 29234 10265
rect 28854 10225 28866 10259
rect 28854 10187 28886 10225
rect 29220 10187 29234 10225
rect 28854 10153 28866 10187
rect 28854 10147 28886 10153
rect 28632 10146 28642 10147
rect 28876 10146 28886 10147
rect 29220 10147 29234 10153
rect 29442 10259 29474 10265
rect 29808 10265 29818 10266
rect 30052 10265 30062 10266
rect 29808 10259 29822 10265
rect 29442 10225 29454 10259
rect 29442 10187 29474 10225
rect 29808 10187 29822 10225
rect 29442 10153 29454 10187
rect 29442 10147 29474 10153
rect 29220 10146 29230 10147
rect 29464 10146 29474 10147
rect 29808 10147 29822 10153
rect 30030 10259 30062 10265
rect 30396 10265 30406 10266
rect 30640 10265 30650 10266
rect 30396 10259 30410 10265
rect 30030 10225 30042 10259
rect 30030 10187 30062 10225
rect 30396 10187 30410 10225
rect 30030 10153 30042 10187
rect 30030 10147 30062 10153
rect 29808 10146 29818 10147
rect 30052 10146 30062 10147
rect 30396 10147 30410 10153
rect 30618 10259 30650 10265
rect 30984 10265 30994 10266
rect 31228 10265 31238 10266
rect 30984 10259 30998 10265
rect 30618 10225 30630 10259
rect 30618 10187 30650 10225
rect 30984 10187 30998 10225
rect 30618 10153 30630 10187
rect 30618 10147 30650 10153
rect 30396 10146 30406 10147
rect 30640 10146 30650 10147
rect 30984 10147 30998 10153
rect 31206 10259 31238 10265
rect 31572 10265 31582 10266
rect 31816 10265 31826 10266
rect 31572 10259 31586 10265
rect 31206 10225 31218 10259
rect 31206 10187 31238 10225
rect 31572 10187 31586 10225
rect 31206 10153 31218 10187
rect 31206 10147 31238 10153
rect 30984 10146 30994 10147
rect 31228 10146 31238 10147
rect 31572 10147 31586 10153
rect 31794 10259 31826 10265
rect 32160 10265 32170 10266
rect 32404 10265 32414 10266
rect 32160 10259 32174 10265
rect 31794 10225 31806 10259
rect 31794 10187 31826 10225
rect 32160 10187 32174 10225
rect 31794 10153 31806 10187
rect 31794 10147 31826 10153
rect 31572 10146 31582 10147
rect 31816 10146 31826 10147
rect 32160 10147 32174 10153
rect 32382 10259 32414 10265
rect 32748 10265 32758 10266
rect 32992 10265 33002 10266
rect 32748 10259 32762 10265
rect 32382 10225 32394 10259
rect 32382 10187 32414 10225
rect 32748 10187 32762 10225
rect 32382 10153 32394 10187
rect 32382 10147 32414 10153
rect 32160 10146 32170 10147
rect 32404 10146 32414 10147
rect 32748 10147 32762 10153
rect 32970 10259 33002 10265
rect 33336 10265 33346 10266
rect 33580 10265 33590 10266
rect 33336 10259 33350 10265
rect 32970 10225 32982 10259
rect 32970 10187 33002 10225
rect 33336 10187 33350 10225
rect 32970 10153 32982 10187
rect 32970 10147 33002 10153
rect 32748 10146 32758 10147
rect 32992 10146 33002 10147
rect 33336 10147 33350 10153
rect 33558 10259 33590 10265
rect 33924 10265 33934 10266
rect 34168 10265 34178 10266
rect 33924 10259 33938 10265
rect 33558 10225 33570 10259
rect 33558 10187 33590 10225
rect 33924 10187 33938 10225
rect 33558 10153 33570 10187
rect 33558 10147 33590 10153
rect 33336 10146 33346 10147
rect 33580 10146 33590 10147
rect 33924 10147 33938 10153
rect 34146 10259 34178 10265
rect 34512 10265 34522 10266
rect 34756 10265 34766 10266
rect 34512 10259 34526 10265
rect 34146 10225 34158 10259
rect 34146 10187 34178 10225
rect 34512 10187 34526 10225
rect 34146 10153 34158 10187
rect 34146 10147 34178 10153
rect 33924 10146 33934 10147
rect 34168 10146 34178 10147
rect 34512 10147 34526 10153
rect 34734 10259 34766 10265
rect 35100 10265 35110 10266
rect 35344 10265 35354 10266
rect 35100 10259 35114 10265
rect 34734 10225 34746 10259
rect 34734 10187 34766 10225
rect 35100 10187 35114 10225
rect 34734 10153 34746 10187
rect 34734 10147 34766 10153
rect 34512 10146 34522 10147
rect 34756 10146 34766 10147
rect 35100 10147 35114 10153
rect 35322 10259 35354 10265
rect 35688 10265 35698 10266
rect 35932 10265 35942 10266
rect 35688 10259 35702 10265
rect 35322 10225 35334 10259
rect 35322 10187 35354 10225
rect 35688 10187 35702 10225
rect 35322 10153 35334 10187
rect 35322 10147 35354 10153
rect 35100 10146 35110 10147
rect 35344 10146 35354 10147
rect 35688 10147 35702 10153
rect 35910 10259 35942 10265
rect 36276 10265 36286 10266
rect 36520 10265 36530 10266
rect 36276 10259 36290 10265
rect 35910 10225 35922 10259
rect 35910 10187 35942 10225
rect 36276 10187 36290 10225
rect 35910 10153 35922 10187
rect 35910 10147 35942 10153
rect 35688 10146 35698 10147
rect 35932 10146 35942 10147
rect 36276 10147 36290 10153
rect 36498 10259 36530 10265
rect 36864 10265 36874 10266
rect 37108 10265 37118 10266
rect 36864 10259 36878 10265
rect 36498 10225 36510 10259
rect 36498 10187 36530 10225
rect 36864 10187 36878 10225
rect 36498 10153 36510 10187
rect 36498 10147 36530 10153
rect 36276 10146 36286 10147
rect 36520 10146 36530 10147
rect 36864 10147 36878 10153
rect 37086 10259 37118 10265
rect 37452 10265 37462 10266
rect 37696 10265 37706 10266
rect 37452 10259 37466 10265
rect 37086 10225 37098 10259
rect 37086 10187 37118 10225
rect 37452 10187 37466 10225
rect 37086 10153 37098 10187
rect 37086 10147 37118 10153
rect 36864 10146 36874 10147
rect 37108 10146 37118 10147
rect 37452 10147 37466 10153
rect 37674 10259 37706 10265
rect 38040 10265 38050 10266
rect 38284 10265 38294 10266
rect 38040 10259 38054 10265
rect 37674 10225 37686 10259
rect 37674 10187 37706 10225
rect 38040 10187 38054 10225
rect 37674 10153 37686 10187
rect 37674 10147 37706 10153
rect 37452 10146 37462 10147
rect 37696 10146 37706 10147
rect 38040 10147 38054 10153
rect 38262 10259 38294 10265
rect 38628 10265 38638 10266
rect 38628 10259 38642 10265
rect 38262 10225 38274 10259
rect 38262 10187 38294 10225
rect 38628 10187 38642 10225
rect 38262 10153 38274 10187
rect 38262 10147 38294 10153
rect 38040 10146 38050 10147
rect 38284 10146 38294 10147
rect 38628 10147 38642 10153
rect 38628 10146 38638 10147
rect 10670 9265 10680 9276
rect 10638 9259 10680 9265
rect 10946 9265 10956 9276
rect 11258 9265 11268 9276
rect 10946 9259 11006 9265
rect 10638 9187 10680 9225
rect 10946 9187 11006 9225
rect 10638 9147 10680 9153
rect 10670 9128 10680 9147
rect 10946 9147 11006 9153
rect 11226 9259 11268 9265
rect 11534 9265 11544 9276
rect 11846 9265 11856 9276
rect 11534 9259 11594 9265
rect 11226 9187 11268 9225
rect 11534 9187 11594 9225
rect 11226 9147 11268 9153
rect 10946 9128 10956 9147
rect 11258 9128 11268 9147
rect 11534 9147 11594 9153
rect 11814 9259 11856 9265
rect 12122 9265 12132 9276
rect 12434 9265 12444 9276
rect 12122 9259 12182 9265
rect 11814 9187 11856 9225
rect 12122 9187 12182 9225
rect 11814 9147 11856 9153
rect 11534 9128 11544 9147
rect 11846 9128 11856 9147
rect 12122 9147 12182 9153
rect 12402 9259 12444 9265
rect 12710 9265 12720 9276
rect 13022 9265 13032 9276
rect 12710 9259 12770 9265
rect 12402 9187 12444 9225
rect 12710 9187 12770 9225
rect 12402 9147 12444 9153
rect 12122 9128 12132 9147
rect 12434 9128 12444 9147
rect 12710 9147 12770 9153
rect 12990 9259 13032 9265
rect 13298 9265 13308 9276
rect 13610 9265 13620 9276
rect 13298 9259 13358 9265
rect 12990 9187 13032 9225
rect 13298 9187 13358 9225
rect 12990 9147 13032 9153
rect 12710 9128 12720 9147
rect 13022 9128 13032 9147
rect 13298 9147 13358 9153
rect 13578 9259 13620 9265
rect 13886 9265 13896 9276
rect 14198 9265 14208 9276
rect 13886 9259 13946 9265
rect 13578 9187 13620 9225
rect 13886 9187 13946 9225
rect 13578 9147 13620 9153
rect 13298 9128 13308 9147
rect 13610 9128 13620 9147
rect 13886 9147 13946 9153
rect 14166 9259 14208 9265
rect 14474 9265 14484 9276
rect 14786 9265 14796 9276
rect 14474 9259 14534 9265
rect 14166 9187 14208 9225
rect 14474 9187 14534 9225
rect 14166 9147 14208 9153
rect 13886 9128 13896 9147
rect 14198 9128 14208 9147
rect 14474 9147 14534 9153
rect 14754 9259 14796 9265
rect 15062 9265 15072 9276
rect 15374 9265 15384 9276
rect 15062 9259 15122 9265
rect 14754 9187 14796 9225
rect 15062 9187 15122 9225
rect 14754 9147 14796 9153
rect 14474 9128 14484 9147
rect 14786 9128 14796 9147
rect 15062 9147 15122 9153
rect 15342 9259 15384 9265
rect 15650 9265 15660 9276
rect 15962 9265 15972 9276
rect 15650 9259 15710 9265
rect 15342 9187 15384 9225
rect 15650 9187 15710 9225
rect 15342 9147 15384 9153
rect 15062 9128 15072 9147
rect 15374 9128 15384 9147
rect 15650 9147 15710 9153
rect 15930 9259 15972 9265
rect 16238 9265 16248 9276
rect 16550 9265 16560 9276
rect 16238 9259 16298 9265
rect 15930 9187 15972 9225
rect 16238 9187 16298 9225
rect 15930 9147 15972 9153
rect 15650 9128 15660 9147
rect 15962 9128 15972 9147
rect 16238 9147 16298 9153
rect 16518 9259 16560 9265
rect 16826 9265 16836 9276
rect 17138 9265 17148 9276
rect 16826 9259 16886 9265
rect 16518 9187 16560 9225
rect 16826 9187 16886 9225
rect 16518 9147 16560 9153
rect 16238 9128 16248 9147
rect 16550 9128 16560 9147
rect 16826 9147 16886 9153
rect 17106 9259 17148 9265
rect 17414 9265 17424 9276
rect 17726 9265 17736 9276
rect 17414 9259 17474 9265
rect 17106 9187 17148 9225
rect 17414 9187 17474 9225
rect 17106 9147 17148 9153
rect 16826 9128 16836 9147
rect 17138 9128 17148 9147
rect 17414 9147 17474 9153
rect 17694 9259 17736 9265
rect 18002 9265 18012 9276
rect 18314 9265 18324 9276
rect 18002 9259 18062 9265
rect 17694 9187 17736 9225
rect 18002 9187 18062 9225
rect 17694 9147 17736 9153
rect 17414 9128 17424 9147
rect 17726 9128 17736 9147
rect 18002 9147 18062 9153
rect 18282 9259 18324 9265
rect 18590 9265 18600 9276
rect 18902 9265 18912 9276
rect 18590 9259 18650 9265
rect 18282 9187 18324 9225
rect 18590 9187 18650 9225
rect 18282 9147 18324 9153
rect 18002 9128 18012 9147
rect 18314 9128 18324 9147
rect 18590 9147 18650 9153
rect 18870 9259 18912 9265
rect 19178 9265 19188 9276
rect 19490 9265 19500 9276
rect 19178 9259 19238 9265
rect 18870 9187 18912 9225
rect 19178 9187 19238 9225
rect 18870 9147 18912 9153
rect 18590 9128 18600 9147
rect 18902 9128 18912 9147
rect 19178 9147 19238 9153
rect 19458 9259 19500 9265
rect 19766 9265 19776 9276
rect 20078 9265 20088 9276
rect 19766 9259 19826 9265
rect 19458 9187 19500 9225
rect 19766 9187 19826 9225
rect 19458 9147 19500 9153
rect 19178 9128 19188 9147
rect 19490 9128 19500 9147
rect 19766 9147 19826 9153
rect 20046 9259 20088 9265
rect 20354 9265 20364 9276
rect 20666 9265 20676 9276
rect 20354 9259 20414 9265
rect 20046 9187 20088 9225
rect 20354 9187 20414 9225
rect 20046 9147 20088 9153
rect 19766 9128 19776 9147
rect 20078 9128 20088 9147
rect 20354 9147 20414 9153
rect 20634 9259 20676 9265
rect 20942 9265 20952 9276
rect 21254 9265 21264 9276
rect 20942 9259 21002 9265
rect 20634 9187 20676 9225
rect 20942 9187 21002 9225
rect 20634 9147 20676 9153
rect 20354 9128 20364 9147
rect 20666 9128 20676 9147
rect 20942 9147 21002 9153
rect 21222 9259 21264 9265
rect 21530 9265 21540 9276
rect 21842 9265 21852 9276
rect 21530 9259 21590 9265
rect 21222 9187 21264 9225
rect 21530 9187 21590 9225
rect 21222 9147 21264 9153
rect 20942 9128 20952 9147
rect 21254 9128 21264 9147
rect 21530 9147 21590 9153
rect 21810 9259 21852 9265
rect 22118 9265 22128 9276
rect 22118 9259 22178 9265
rect 21810 9187 21852 9225
rect 22118 9187 22178 9225
rect 21810 9147 21852 9153
rect 21530 9128 21540 9147
rect 21842 9128 21852 9147
rect 22118 9147 22178 9153
rect 22118 9128 22128 9147
rect 22408 9126 22418 9286
rect 22750 9126 22760 9286
rect 22996 9265 23006 9286
rect 22986 9259 23006 9265
rect 23338 9265 23348 9286
rect 23584 9265 23594 9286
rect 23338 9259 23354 9265
rect 22986 9187 23006 9225
rect 23338 9187 23354 9225
rect 22986 9147 23006 9153
rect 22996 9126 23006 9147
rect 23338 9147 23354 9153
rect 23574 9259 23594 9265
rect 23926 9265 23936 9286
rect 24172 9265 24182 9286
rect 23926 9259 23942 9265
rect 23574 9187 23594 9225
rect 23926 9187 23942 9225
rect 23574 9147 23594 9153
rect 23338 9126 23348 9147
rect 23584 9126 23594 9147
rect 23926 9147 23942 9153
rect 24162 9259 24182 9265
rect 24514 9265 24524 9286
rect 24760 9265 24770 9286
rect 24514 9259 24530 9265
rect 24162 9187 24182 9225
rect 24514 9187 24530 9225
rect 24162 9147 24182 9153
rect 23926 9126 23936 9147
rect 24172 9126 24182 9147
rect 24514 9147 24530 9153
rect 24750 9259 24770 9265
rect 25102 9265 25112 9286
rect 25348 9265 25358 9286
rect 25102 9259 25118 9265
rect 24750 9187 24770 9225
rect 25102 9187 25118 9225
rect 24750 9147 24770 9153
rect 24514 9126 24524 9147
rect 24760 9126 24770 9147
rect 25102 9147 25118 9153
rect 25338 9259 25358 9265
rect 25690 9265 25700 9286
rect 25936 9265 25946 9286
rect 25690 9259 25706 9265
rect 25338 9187 25358 9225
rect 25690 9187 25706 9225
rect 25338 9147 25358 9153
rect 25102 9126 25112 9147
rect 25348 9126 25358 9147
rect 25690 9147 25706 9153
rect 25926 9259 25946 9265
rect 26278 9265 26288 9286
rect 26524 9265 26534 9286
rect 26278 9259 26294 9265
rect 25926 9187 25946 9225
rect 26278 9187 26294 9225
rect 25926 9147 25946 9153
rect 25690 9126 25700 9147
rect 25936 9126 25946 9147
rect 26278 9147 26294 9153
rect 26514 9259 26534 9265
rect 26866 9265 26876 9286
rect 27112 9265 27122 9286
rect 26866 9259 26882 9265
rect 26514 9187 26534 9225
rect 26866 9187 26882 9225
rect 26514 9147 26534 9153
rect 26278 9126 26288 9147
rect 26524 9126 26534 9147
rect 26866 9147 26882 9153
rect 27102 9259 27122 9265
rect 27454 9265 27464 9286
rect 27700 9265 27710 9286
rect 27454 9259 27470 9265
rect 27102 9187 27122 9225
rect 27454 9187 27470 9225
rect 27102 9147 27122 9153
rect 26866 9126 26876 9147
rect 27112 9126 27122 9147
rect 27454 9147 27470 9153
rect 27690 9259 27710 9265
rect 28042 9265 28052 9286
rect 28288 9265 28298 9286
rect 28042 9259 28058 9265
rect 27690 9187 27710 9225
rect 28042 9187 28058 9225
rect 27690 9147 27710 9153
rect 27454 9126 27464 9147
rect 27700 9126 27710 9147
rect 28042 9147 28058 9153
rect 28278 9259 28298 9265
rect 28630 9265 28640 9286
rect 28876 9265 28886 9286
rect 28630 9259 28646 9265
rect 28278 9187 28298 9225
rect 28630 9187 28646 9225
rect 28278 9147 28298 9153
rect 28042 9126 28052 9147
rect 28288 9126 28298 9147
rect 28630 9147 28646 9153
rect 28866 9259 28886 9265
rect 29218 9265 29228 9286
rect 29464 9265 29474 9286
rect 29218 9259 29234 9265
rect 28866 9187 28886 9225
rect 29218 9187 29234 9225
rect 28866 9147 28886 9153
rect 28630 9126 28640 9147
rect 28876 9126 28886 9147
rect 29218 9147 29234 9153
rect 29454 9259 29474 9265
rect 29806 9265 29816 9286
rect 30052 9265 30062 9286
rect 29806 9259 29822 9265
rect 29454 9187 29474 9225
rect 29806 9187 29822 9225
rect 29454 9147 29474 9153
rect 29218 9126 29228 9147
rect 29464 9126 29474 9147
rect 29806 9147 29822 9153
rect 30042 9259 30062 9265
rect 30394 9265 30404 9286
rect 30640 9265 30650 9286
rect 30394 9259 30410 9265
rect 30042 9187 30062 9225
rect 30394 9187 30410 9225
rect 30042 9147 30062 9153
rect 29806 9126 29816 9147
rect 30052 9126 30062 9147
rect 30394 9147 30410 9153
rect 30630 9259 30650 9265
rect 30982 9265 30992 9286
rect 31228 9265 31238 9286
rect 30982 9259 30998 9265
rect 30630 9187 30650 9225
rect 30982 9187 30998 9225
rect 30630 9147 30650 9153
rect 30394 9126 30404 9147
rect 30640 9126 30650 9147
rect 30982 9147 30998 9153
rect 31218 9259 31238 9265
rect 31570 9265 31580 9286
rect 31816 9265 31826 9286
rect 31570 9259 31586 9265
rect 31218 9187 31238 9225
rect 31570 9187 31586 9225
rect 31218 9147 31238 9153
rect 30982 9126 30992 9147
rect 31228 9126 31238 9147
rect 31570 9147 31586 9153
rect 31806 9259 31826 9265
rect 32158 9265 32168 9286
rect 32404 9265 32414 9286
rect 32158 9259 32174 9265
rect 31806 9187 31826 9225
rect 32158 9187 32174 9225
rect 31806 9147 31826 9153
rect 31570 9126 31580 9147
rect 31816 9126 31826 9147
rect 32158 9147 32174 9153
rect 32394 9259 32414 9265
rect 32746 9265 32756 9286
rect 32992 9265 33002 9286
rect 32746 9259 32762 9265
rect 32394 9187 32414 9225
rect 32746 9187 32762 9225
rect 32394 9147 32414 9153
rect 32158 9126 32168 9147
rect 32404 9126 32414 9147
rect 32746 9147 32762 9153
rect 32982 9259 33002 9265
rect 33334 9265 33344 9286
rect 33580 9265 33590 9286
rect 33334 9259 33350 9265
rect 32982 9187 33002 9225
rect 33334 9187 33350 9225
rect 32982 9147 33002 9153
rect 32746 9126 32756 9147
rect 32992 9126 33002 9147
rect 33334 9147 33350 9153
rect 33570 9259 33590 9265
rect 33922 9265 33932 9286
rect 34168 9265 34178 9286
rect 33922 9259 33938 9265
rect 33570 9187 33590 9225
rect 33922 9187 33938 9225
rect 33570 9147 33590 9153
rect 33334 9126 33344 9147
rect 33580 9126 33590 9147
rect 33922 9147 33938 9153
rect 34158 9259 34178 9265
rect 34510 9265 34520 9286
rect 34756 9265 34766 9286
rect 34510 9259 34526 9265
rect 34158 9187 34178 9225
rect 34510 9187 34526 9225
rect 34158 9147 34178 9153
rect 33922 9126 33932 9147
rect 34168 9126 34178 9147
rect 34510 9147 34526 9153
rect 34746 9259 34766 9265
rect 35098 9265 35108 9286
rect 35344 9265 35354 9286
rect 35098 9259 35114 9265
rect 34746 9187 34766 9225
rect 35098 9187 35114 9225
rect 34746 9147 34766 9153
rect 34510 9126 34520 9147
rect 34756 9126 34766 9147
rect 35098 9147 35114 9153
rect 35334 9259 35354 9265
rect 35686 9265 35696 9286
rect 35932 9265 35942 9286
rect 35686 9259 35702 9265
rect 35334 9187 35354 9225
rect 35686 9187 35702 9225
rect 35334 9147 35354 9153
rect 35098 9126 35108 9147
rect 35344 9126 35354 9147
rect 35686 9147 35702 9153
rect 35922 9259 35942 9265
rect 36274 9265 36284 9286
rect 36520 9265 36530 9286
rect 36274 9259 36290 9265
rect 35922 9187 35942 9225
rect 36274 9187 36290 9225
rect 35922 9147 35942 9153
rect 35686 9126 35696 9147
rect 35932 9126 35942 9147
rect 36274 9147 36290 9153
rect 36510 9259 36530 9265
rect 36862 9265 36872 9286
rect 37108 9265 37118 9286
rect 36862 9259 36878 9265
rect 36510 9187 36530 9225
rect 36862 9187 36878 9225
rect 36510 9147 36530 9153
rect 36274 9126 36284 9147
rect 36520 9126 36530 9147
rect 36862 9147 36878 9153
rect 37098 9259 37118 9265
rect 37450 9265 37460 9286
rect 37696 9265 37706 9286
rect 37450 9259 37466 9265
rect 37098 9187 37118 9225
rect 37450 9187 37466 9225
rect 37098 9147 37118 9153
rect 36862 9126 36872 9147
rect 37108 9126 37118 9147
rect 37450 9147 37466 9153
rect 37686 9259 37706 9265
rect 38038 9265 38048 9286
rect 38284 9265 38294 9286
rect 38038 9259 38054 9265
rect 37686 9187 37706 9225
rect 38038 9187 38054 9225
rect 37686 9147 37706 9153
rect 37450 9126 37460 9147
rect 37696 9126 37706 9147
rect 38038 9147 38054 9153
rect 38274 9259 38294 9265
rect 38626 9265 38636 9286
rect 38626 9259 38642 9265
rect 38274 9187 38294 9225
rect 38626 9187 38642 9225
rect 38274 9147 38294 9153
rect 38038 9126 38048 9147
rect 38284 9126 38294 9147
rect 38626 9147 38642 9153
rect 38626 9126 38636 9147
rect 10656 8208 10666 8276
rect 10984 8208 10994 8276
rect 11244 8265 11254 8276
rect 11226 8259 11254 8265
rect 11572 8265 11582 8276
rect 11832 8265 11842 8276
rect 11572 8259 11594 8265
rect 11226 8219 11254 8225
rect 11244 8208 11254 8219
rect 11572 8219 11594 8225
rect 11814 8259 11842 8265
rect 12160 8265 12170 8276
rect 12420 8265 12430 8276
rect 12160 8259 12182 8265
rect 11814 8219 11842 8225
rect 11572 8208 11582 8219
rect 11832 8208 11842 8219
rect 12160 8219 12182 8225
rect 12402 8259 12430 8265
rect 12748 8265 12758 8276
rect 13008 8265 13018 8276
rect 12748 8259 12770 8265
rect 12402 8219 12430 8225
rect 12160 8208 12170 8219
rect 12420 8208 12430 8219
rect 12748 8219 12770 8225
rect 12990 8259 13018 8265
rect 13336 8265 13346 8276
rect 13596 8265 13606 8276
rect 13336 8259 13358 8265
rect 12990 8219 13018 8225
rect 12748 8208 12758 8219
rect 13008 8208 13018 8219
rect 13336 8219 13358 8225
rect 13578 8259 13606 8265
rect 13924 8265 13934 8276
rect 14184 8265 14194 8276
rect 13924 8259 13946 8265
rect 13578 8219 13606 8225
rect 13336 8208 13346 8219
rect 13596 8208 13606 8219
rect 13924 8219 13946 8225
rect 14166 8259 14194 8265
rect 14512 8265 14522 8276
rect 14772 8265 14782 8276
rect 14512 8259 14534 8265
rect 14166 8219 14194 8225
rect 13924 8208 13934 8219
rect 14184 8208 14194 8219
rect 14512 8219 14534 8225
rect 14754 8259 14782 8265
rect 15100 8265 15110 8276
rect 15360 8265 15370 8276
rect 15100 8259 15122 8265
rect 14754 8219 14782 8225
rect 14512 8208 14522 8219
rect 14772 8208 14782 8219
rect 15100 8219 15122 8225
rect 15342 8259 15370 8265
rect 15688 8265 15698 8276
rect 15948 8265 15958 8276
rect 15688 8259 15710 8265
rect 15342 8219 15370 8225
rect 15100 8208 15110 8219
rect 15360 8208 15370 8219
rect 15688 8219 15710 8225
rect 15930 8259 15958 8265
rect 16276 8265 16286 8276
rect 16536 8265 16546 8276
rect 16276 8259 16298 8265
rect 15930 8219 15958 8225
rect 15688 8208 15698 8219
rect 15948 8208 15958 8219
rect 16276 8219 16298 8225
rect 16518 8259 16546 8265
rect 16864 8265 16874 8276
rect 17124 8265 17134 8276
rect 16864 8259 16886 8265
rect 16518 8219 16546 8225
rect 16276 8208 16286 8219
rect 16536 8208 16546 8219
rect 16864 8219 16886 8225
rect 17106 8259 17134 8265
rect 17452 8265 17462 8276
rect 17712 8265 17722 8276
rect 17452 8259 17474 8265
rect 17106 8219 17134 8225
rect 16864 8208 16874 8219
rect 17124 8208 17134 8219
rect 17452 8219 17474 8225
rect 17694 8259 17722 8265
rect 18040 8265 18050 8276
rect 18300 8265 18310 8276
rect 18040 8259 18062 8265
rect 17694 8219 17722 8225
rect 17452 8208 17462 8219
rect 17712 8208 17722 8219
rect 18040 8219 18062 8225
rect 18282 8259 18310 8265
rect 18628 8265 18638 8276
rect 18888 8265 18898 8276
rect 18628 8259 18650 8265
rect 18282 8219 18310 8225
rect 18040 8208 18050 8219
rect 18300 8208 18310 8219
rect 18628 8219 18650 8225
rect 18870 8259 18898 8265
rect 19216 8265 19226 8276
rect 19476 8265 19486 8276
rect 19216 8259 19238 8265
rect 18870 8219 18898 8225
rect 18628 8208 18638 8219
rect 18888 8208 18898 8219
rect 19216 8219 19238 8225
rect 19458 8259 19486 8265
rect 19804 8265 19814 8276
rect 20064 8265 20074 8276
rect 19804 8259 19826 8265
rect 19458 8219 19486 8225
rect 19216 8208 19226 8219
rect 19476 8208 19486 8219
rect 19804 8219 19826 8225
rect 20046 8259 20074 8265
rect 20392 8265 20402 8276
rect 20652 8265 20662 8276
rect 20392 8259 20414 8265
rect 20046 8219 20074 8225
rect 19804 8208 19814 8219
rect 20064 8208 20074 8219
rect 20392 8219 20414 8225
rect 20634 8259 20662 8265
rect 20980 8265 20990 8276
rect 21240 8265 21250 8276
rect 20980 8259 21002 8265
rect 20634 8219 20662 8225
rect 20392 8208 20402 8219
rect 20652 8208 20662 8219
rect 20980 8219 21002 8225
rect 21222 8259 21250 8265
rect 21568 8265 21578 8276
rect 21828 8265 21838 8276
rect 21568 8259 21590 8265
rect 21222 8219 21250 8225
rect 20980 8208 20990 8219
rect 21240 8208 21250 8219
rect 21568 8219 21590 8225
rect 21810 8259 21838 8265
rect 22156 8265 22166 8276
rect 22156 8259 22178 8265
rect 21810 8219 21838 8225
rect 21568 8208 21578 8219
rect 21828 8208 21838 8219
rect 22156 8219 22178 8225
rect 22156 8208 22166 8219
rect 22424 8196 22434 8274
rect 22712 8196 22722 8274
rect 23012 8265 23022 8274
rect 22986 8259 23022 8265
rect 23300 8265 23310 8274
rect 23600 8265 23610 8274
rect 23300 8259 23354 8265
rect 22986 8219 23022 8225
rect 23012 8196 23022 8219
rect 23300 8219 23354 8225
rect 23574 8259 23610 8265
rect 23888 8265 23898 8274
rect 24188 8265 24198 8274
rect 23888 8259 23942 8265
rect 23574 8219 23610 8225
rect 23300 8196 23310 8219
rect 23600 8196 23610 8219
rect 23888 8219 23942 8225
rect 24162 8259 24198 8265
rect 24476 8265 24486 8274
rect 24776 8265 24786 8274
rect 24476 8259 24530 8265
rect 24162 8219 24198 8225
rect 23888 8196 23898 8219
rect 24188 8196 24198 8219
rect 24476 8219 24530 8225
rect 24750 8259 24786 8265
rect 25064 8265 25074 8274
rect 25364 8265 25374 8274
rect 25064 8259 25118 8265
rect 24750 8219 24786 8225
rect 24476 8196 24486 8219
rect 24776 8196 24786 8219
rect 25064 8219 25118 8225
rect 25338 8259 25374 8265
rect 25652 8265 25662 8274
rect 25952 8265 25962 8274
rect 25652 8259 25706 8265
rect 25338 8219 25374 8225
rect 25064 8196 25074 8219
rect 25364 8196 25374 8219
rect 25652 8219 25706 8225
rect 25926 8259 25962 8265
rect 26240 8265 26250 8274
rect 26540 8265 26550 8274
rect 26240 8259 26294 8265
rect 25926 8219 25962 8225
rect 25652 8196 25662 8219
rect 25952 8196 25962 8219
rect 26240 8219 26294 8225
rect 26514 8259 26550 8265
rect 26828 8265 26838 8274
rect 27128 8265 27138 8274
rect 26828 8259 26882 8265
rect 26514 8219 26550 8225
rect 26240 8196 26250 8219
rect 26540 8196 26550 8219
rect 26828 8219 26882 8225
rect 27102 8259 27138 8265
rect 27416 8265 27426 8274
rect 27716 8265 27726 8274
rect 27416 8259 27470 8265
rect 27102 8219 27138 8225
rect 26828 8196 26838 8219
rect 27128 8196 27138 8219
rect 27416 8219 27470 8225
rect 27690 8259 27726 8265
rect 28004 8265 28014 8274
rect 28304 8265 28314 8274
rect 28004 8259 28058 8265
rect 27690 8219 27726 8225
rect 27416 8196 27426 8219
rect 27716 8196 27726 8219
rect 28004 8219 28058 8225
rect 28278 8259 28314 8265
rect 28592 8265 28602 8274
rect 28892 8265 28902 8274
rect 28592 8259 28646 8265
rect 28278 8219 28314 8225
rect 28004 8196 28014 8219
rect 28304 8196 28314 8219
rect 28592 8219 28646 8225
rect 28866 8259 28902 8265
rect 29180 8265 29190 8274
rect 29480 8265 29490 8274
rect 29180 8259 29234 8265
rect 28866 8219 28902 8225
rect 28592 8196 28602 8219
rect 28892 8196 28902 8219
rect 29180 8219 29234 8225
rect 29454 8259 29490 8265
rect 29768 8265 29778 8274
rect 30068 8265 30078 8274
rect 29768 8259 29822 8265
rect 29454 8219 29490 8225
rect 29180 8196 29190 8219
rect 29480 8196 29490 8219
rect 29768 8219 29822 8225
rect 30042 8259 30078 8265
rect 30356 8265 30366 8274
rect 30656 8265 30666 8274
rect 30356 8259 30410 8265
rect 30042 8219 30078 8225
rect 29768 8196 29778 8219
rect 30068 8196 30078 8219
rect 30356 8219 30410 8225
rect 30630 8259 30666 8265
rect 30944 8265 30954 8274
rect 31244 8265 31254 8274
rect 30944 8259 30998 8265
rect 30630 8219 30666 8225
rect 30356 8196 30366 8219
rect 30656 8196 30666 8219
rect 30944 8219 30998 8225
rect 31218 8259 31254 8265
rect 31532 8265 31542 8274
rect 31832 8265 31842 8274
rect 31532 8259 31586 8265
rect 31218 8219 31254 8225
rect 30944 8196 30954 8219
rect 31244 8196 31254 8219
rect 31532 8219 31586 8225
rect 31806 8259 31842 8265
rect 32120 8265 32130 8274
rect 32420 8265 32430 8274
rect 32120 8259 32174 8265
rect 31806 8219 31842 8225
rect 31532 8196 31542 8219
rect 31832 8196 31842 8219
rect 32120 8219 32174 8225
rect 32394 8259 32430 8265
rect 32708 8265 32718 8274
rect 33008 8265 33018 8274
rect 32708 8259 32762 8265
rect 32394 8219 32430 8225
rect 32120 8196 32130 8219
rect 32420 8196 32430 8219
rect 32708 8219 32762 8225
rect 32982 8259 33018 8265
rect 33296 8265 33306 8274
rect 33596 8265 33606 8274
rect 33296 8259 33350 8265
rect 32982 8219 33018 8225
rect 32708 8196 32718 8219
rect 33008 8196 33018 8219
rect 33296 8219 33350 8225
rect 33570 8259 33606 8265
rect 33884 8265 33894 8274
rect 34184 8265 34194 8274
rect 33884 8259 33938 8265
rect 33570 8219 33606 8225
rect 33296 8196 33306 8219
rect 33596 8196 33606 8219
rect 33884 8219 33938 8225
rect 34158 8259 34194 8265
rect 34472 8265 34482 8274
rect 34772 8265 34782 8274
rect 34472 8259 34526 8265
rect 34158 8219 34194 8225
rect 33884 8196 33894 8219
rect 34184 8196 34194 8219
rect 34472 8219 34526 8225
rect 34746 8259 34782 8265
rect 35060 8265 35070 8274
rect 35360 8265 35370 8274
rect 35060 8259 35114 8265
rect 34746 8219 34782 8225
rect 34472 8196 34482 8219
rect 34772 8196 34782 8219
rect 35060 8219 35114 8225
rect 35334 8259 35370 8265
rect 35648 8265 35658 8274
rect 35948 8265 35958 8274
rect 35648 8259 35702 8265
rect 35334 8219 35370 8225
rect 35060 8196 35070 8219
rect 35360 8196 35370 8219
rect 35648 8219 35702 8225
rect 35922 8259 35958 8265
rect 36236 8265 36246 8274
rect 36536 8265 36546 8274
rect 36236 8259 36290 8265
rect 35922 8219 35958 8225
rect 35648 8196 35658 8219
rect 35948 8196 35958 8219
rect 36236 8219 36290 8225
rect 36510 8259 36546 8265
rect 36824 8265 36834 8274
rect 37124 8265 37134 8274
rect 36824 8259 36878 8265
rect 36510 8219 36546 8225
rect 36236 8196 36246 8219
rect 36536 8196 36546 8219
rect 36824 8219 36878 8225
rect 37098 8259 37134 8265
rect 37412 8265 37422 8274
rect 37712 8265 37722 8274
rect 37412 8259 37466 8265
rect 37098 8219 37134 8225
rect 36824 8196 36834 8219
rect 37124 8196 37134 8219
rect 37412 8219 37466 8225
rect 37686 8259 37722 8265
rect 38000 8265 38010 8274
rect 38300 8265 38310 8274
rect 38000 8259 38054 8265
rect 37686 8219 37722 8225
rect 37412 8196 37422 8219
rect 37712 8196 37722 8219
rect 38000 8219 38054 8225
rect 38274 8259 38310 8265
rect 38588 8265 38598 8274
rect 38588 8259 38642 8265
rect 38274 8219 38310 8225
rect 38000 8196 38010 8219
rect 38300 8196 38310 8219
rect 38588 8219 38642 8225
rect 38588 8196 38598 8219
rect 44370 6952 45388 18676
rect 44370 6144 44380 6952
rect 45446 6144 45456 6952
rect 6268 3996 6278 4988
rect 7030 3996 7040 4988
<< via1 >>
rect 10622 27490 11022 27548
rect 11210 27531 11610 27548
rect 11210 27497 11226 27531
rect 11226 27497 11594 27531
rect 11594 27497 11610 27531
rect 11210 27490 11610 27497
rect 11798 27531 12198 27548
rect 11798 27497 11814 27531
rect 11814 27497 12182 27531
rect 12182 27497 12198 27531
rect 11798 27490 12198 27497
rect 12386 27531 12786 27548
rect 12386 27497 12402 27531
rect 12402 27497 12770 27531
rect 12770 27497 12786 27531
rect 12386 27490 12786 27497
rect 12974 27531 13374 27548
rect 12974 27497 12990 27531
rect 12990 27497 13358 27531
rect 13358 27497 13374 27531
rect 12974 27490 13374 27497
rect 13562 27531 13962 27548
rect 13562 27497 13578 27531
rect 13578 27497 13946 27531
rect 13946 27497 13962 27531
rect 13562 27490 13962 27497
rect 14150 27531 14550 27548
rect 14150 27497 14166 27531
rect 14166 27497 14534 27531
rect 14534 27497 14550 27531
rect 14150 27490 14550 27497
rect 14738 27531 15138 27548
rect 14738 27497 14754 27531
rect 14754 27497 15122 27531
rect 15122 27497 15138 27531
rect 14738 27490 15138 27497
rect 15326 27531 15726 27548
rect 15326 27497 15342 27531
rect 15342 27497 15710 27531
rect 15710 27497 15726 27531
rect 15326 27490 15726 27497
rect 15914 27531 16314 27548
rect 15914 27497 15930 27531
rect 15930 27497 16298 27531
rect 16298 27497 16314 27531
rect 15914 27490 16314 27497
rect 16502 27531 16902 27548
rect 16502 27497 16518 27531
rect 16518 27497 16886 27531
rect 16886 27497 16902 27531
rect 16502 27490 16902 27497
rect 17090 27531 17490 27548
rect 17090 27497 17106 27531
rect 17106 27497 17474 27531
rect 17474 27497 17490 27531
rect 17090 27490 17490 27497
rect 17678 27531 18078 27548
rect 17678 27497 17694 27531
rect 17694 27497 18062 27531
rect 18062 27497 18078 27531
rect 17678 27490 18078 27497
rect 18266 27531 18666 27548
rect 18266 27497 18282 27531
rect 18282 27497 18650 27531
rect 18650 27497 18666 27531
rect 18266 27490 18666 27497
rect 18854 27531 19254 27548
rect 18854 27497 18870 27531
rect 18870 27497 19238 27531
rect 19238 27497 19254 27531
rect 18854 27490 19254 27497
rect 19442 27531 19842 27548
rect 19442 27497 19458 27531
rect 19458 27497 19826 27531
rect 19826 27497 19842 27531
rect 19442 27490 19842 27497
rect 20030 27531 20430 27548
rect 20030 27497 20046 27531
rect 20046 27497 20414 27531
rect 20414 27497 20430 27531
rect 20030 27490 20430 27497
rect 20618 27531 21018 27548
rect 20618 27497 20634 27531
rect 20634 27497 21002 27531
rect 21002 27497 21018 27531
rect 20618 27490 21018 27497
rect 21206 27531 21606 27548
rect 21206 27497 21222 27531
rect 21222 27497 21590 27531
rect 21590 27497 21606 27531
rect 21206 27490 21606 27497
rect 21802 27486 22178 27542
rect 22398 27488 22766 27542
rect 22986 27531 23354 27542
rect 22986 27497 23354 27531
rect 22986 27488 23354 27497
rect 23574 27531 23942 27542
rect 23574 27497 23942 27531
rect 23574 27488 23942 27497
rect 24162 27531 24530 27542
rect 24162 27497 24530 27531
rect 24162 27488 24530 27497
rect 24750 27531 25118 27542
rect 24750 27497 25118 27531
rect 24750 27488 25118 27497
rect 25338 27531 25706 27542
rect 25338 27497 25706 27531
rect 25338 27488 25706 27497
rect 25926 27531 26294 27542
rect 25926 27497 26294 27531
rect 25926 27488 26294 27497
rect 26514 27531 26882 27542
rect 26514 27497 26882 27531
rect 26514 27488 26882 27497
rect 27102 27531 27470 27542
rect 27102 27497 27470 27531
rect 27102 27488 27470 27497
rect 27690 27531 28058 27542
rect 27690 27497 28058 27531
rect 27690 27488 28058 27497
rect 28278 27531 28646 27542
rect 28278 27497 28646 27531
rect 28278 27488 28646 27497
rect 28866 27531 29234 27542
rect 28866 27497 29234 27531
rect 28866 27488 29234 27497
rect 29454 27531 29822 27542
rect 29454 27497 29822 27531
rect 29454 27488 29822 27497
rect 30042 27531 30410 27542
rect 30042 27497 30410 27531
rect 30042 27488 30410 27497
rect 30630 27531 30998 27542
rect 30630 27497 30998 27531
rect 30630 27488 30998 27497
rect 31218 27531 31586 27542
rect 31218 27497 31586 27531
rect 31218 27488 31586 27497
rect 31806 27531 32174 27542
rect 31806 27497 32174 27531
rect 31806 27488 32174 27497
rect 32394 27531 32762 27542
rect 32394 27497 32762 27531
rect 32394 27488 32762 27497
rect 32982 27531 33350 27542
rect 32982 27497 33350 27531
rect 32982 27488 33350 27497
rect 33570 27531 33938 27542
rect 33570 27497 33938 27531
rect 33570 27488 33938 27497
rect 34158 27531 34526 27542
rect 34158 27497 34526 27531
rect 34158 27488 34526 27497
rect 34746 27531 35114 27542
rect 34746 27497 35114 27531
rect 34746 27488 35114 27497
rect 35334 27531 35702 27542
rect 35334 27497 35702 27531
rect 35334 27488 35702 27497
rect 35922 27531 36290 27542
rect 35922 27497 36290 27531
rect 35922 27488 36290 27497
rect 36510 27531 36878 27542
rect 36510 27497 36878 27531
rect 36510 27488 36878 27497
rect 37098 27531 37466 27542
rect 37098 27497 37466 27531
rect 37098 27488 37466 27497
rect 37686 27531 38054 27542
rect 37686 27497 38054 27531
rect 37686 27488 38054 27497
rect 38274 27531 38642 27542
rect 38274 27497 38642 27531
rect 38274 27488 38642 27497
rect 10638 26490 11006 26604
rect 11226 26603 11594 26604
rect 11226 26569 11594 26603
rect 11226 26531 11594 26569
rect 11226 26497 11594 26531
rect 11226 26490 11594 26497
rect 11814 26603 12182 26604
rect 11814 26569 12182 26603
rect 11814 26531 12182 26569
rect 11814 26497 12182 26531
rect 11814 26490 12182 26497
rect 12402 26603 12770 26604
rect 12402 26569 12770 26603
rect 12402 26531 12770 26569
rect 12402 26497 12770 26531
rect 12402 26490 12770 26497
rect 12990 26603 13358 26604
rect 12990 26569 13358 26603
rect 12990 26531 13358 26569
rect 12990 26497 13358 26531
rect 12990 26490 13358 26497
rect 13578 26603 13946 26604
rect 13578 26569 13946 26603
rect 13578 26531 13946 26569
rect 13578 26497 13946 26531
rect 13578 26490 13946 26497
rect 14166 26603 14534 26604
rect 14166 26569 14534 26603
rect 14166 26531 14534 26569
rect 14166 26497 14534 26531
rect 14166 26490 14534 26497
rect 14754 26603 15122 26604
rect 14754 26569 15122 26603
rect 14754 26531 15122 26569
rect 14754 26497 15122 26531
rect 14754 26490 15122 26497
rect 15342 26603 15710 26604
rect 15342 26569 15710 26603
rect 15342 26531 15710 26569
rect 15342 26497 15710 26531
rect 15342 26490 15710 26497
rect 15930 26603 16298 26604
rect 15930 26569 16298 26603
rect 15930 26531 16298 26569
rect 15930 26497 16298 26531
rect 15930 26490 16298 26497
rect 16518 26603 16886 26604
rect 16518 26569 16886 26603
rect 16518 26531 16886 26569
rect 16518 26497 16886 26531
rect 16518 26490 16886 26497
rect 17106 26603 17474 26604
rect 17106 26569 17474 26603
rect 17106 26531 17474 26569
rect 17106 26497 17474 26531
rect 17106 26490 17474 26497
rect 17694 26603 18062 26604
rect 17694 26569 18062 26603
rect 17694 26531 18062 26569
rect 17694 26497 18062 26531
rect 17694 26490 18062 26497
rect 18282 26603 18650 26604
rect 18282 26569 18650 26603
rect 18282 26531 18650 26569
rect 18282 26497 18650 26531
rect 18282 26490 18650 26497
rect 18870 26603 19238 26604
rect 18870 26569 19238 26603
rect 18870 26531 19238 26569
rect 18870 26497 19238 26531
rect 18870 26490 19238 26497
rect 19458 26603 19826 26604
rect 19458 26569 19826 26603
rect 19458 26531 19826 26569
rect 19458 26497 19826 26531
rect 19458 26490 19826 26497
rect 20046 26603 20414 26604
rect 20046 26569 20414 26603
rect 20046 26531 20414 26569
rect 20046 26497 20414 26531
rect 20046 26490 20414 26497
rect 20634 26603 21002 26604
rect 20634 26569 21002 26603
rect 20634 26531 21002 26569
rect 20634 26497 21002 26531
rect 20634 26490 21002 26497
rect 21222 26603 21590 26604
rect 21222 26569 21590 26603
rect 21222 26531 21590 26569
rect 21222 26497 21590 26531
rect 21222 26490 21590 26497
rect 21810 26603 22178 26604
rect 21810 26569 22178 26603
rect 21810 26531 22178 26569
rect 21810 26497 22178 26531
rect 21810 26490 22178 26497
rect 22398 26496 22766 26604
rect 22986 26603 23354 26604
rect 22986 26569 23354 26603
rect 22986 26531 23354 26569
rect 22986 26497 23354 26531
rect 22986 26496 23354 26497
rect 23574 26603 23942 26604
rect 23574 26569 23942 26603
rect 23574 26531 23942 26569
rect 23574 26497 23942 26531
rect 23574 26496 23942 26497
rect 24162 26603 24530 26604
rect 24162 26569 24530 26603
rect 24162 26531 24530 26569
rect 24162 26497 24530 26531
rect 24162 26496 24530 26497
rect 24750 26603 25118 26604
rect 24750 26569 25118 26603
rect 24750 26531 25118 26569
rect 24750 26497 25118 26531
rect 24750 26496 25118 26497
rect 25338 26603 25706 26604
rect 25338 26569 25706 26603
rect 25338 26531 25706 26569
rect 25338 26497 25706 26531
rect 25338 26496 25706 26497
rect 25926 26603 26294 26604
rect 25926 26569 26294 26603
rect 25926 26531 26294 26569
rect 25926 26497 26294 26531
rect 25926 26496 26294 26497
rect 26514 26603 26882 26604
rect 26514 26569 26882 26603
rect 26514 26531 26882 26569
rect 26514 26497 26882 26531
rect 26514 26496 26882 26497
rect 27102 26603 27470 26604
rect 27102 26569 27470 26603
rect 27102 26531 27470 26569
rect 27102 26497 27470 26531
rect 27102 26496 27470 26497
rect 27690 26603 28058 26604
rect 27690 26569 28058 26603
rect 27690 26531 28058 26569
rect 27690 26497 28058 26531
rect 27690 26496 28058 26497
rect 28278 26603 28646 26604
rect 28278 26569 28646 26603
rect 28278 26531 28646 26569
rect 28278 26497 28646 26531
rect 28278 26496 28646 26497
rect 28866 26603 29234 26604
rect 28866 26569 29234 26603
rect 28866 26531 29234 26569
rect 28866 26497 29234 26531
rect 28866 26496 29234 26497
rect 29454 26603 29822 26604
rect 29454 26569 29822 26603
rect 29454 26531 29822 26569
rect 29454 26497 29822 26531
rect 29454 26496 29822 26497
rect 30042 26603 30410 26604
rect 30042 26569 30410 26603
rect 30042 26531 30410 26569
rect 30042 26497 30410 26531
rect 30042 26496 30410 26497
rect 30630 26603 30998 26604
rect 30630 26569 30998 26603
rect 30630 26531 30998 26569
rect 30630 26497 30998 26531
rect 30630 26496 30998 26497
rect 31218 26603 31586 26604
rect 31218 26569 31586 26603
rect 31218 26531 31586 26569
rect 31218 26497 31586 26531
rect 31218 26496 31586 26497
rect 31806 26603 32174 26604
rect 31806 26569 32174 26603
rect 31806 26531 32174 26569
rect 31806 26497 32174 26531
rect 31806 26496 32174 26497
rect 32394 26603 32762 26604
rect 32394 26569 32762 26603
rect 32394 26531 32762 26569
rect 32394 26497 32762 26531
rect 32394 26496 32762 26497
rect 32982 26603 33350 26604
rect 32982 26569 33350 26603
rect 32982 26531 33350 26569
rect 32982 26497 33350 26531
rect 32982 26496 33350 26497
rect 33570 26603 33938 26604
rect 33570 26569 33938 26603
rect 33570 26531 33938 26569
rect 33570 26497 33938 26531
rect 33570 26496 33938 26497
rect 34158 26603 34526 26604
rect 34158 26569 34526 26603
rect 34158 26531 34526 26569
rect 34158 26497 34526 26531
rect 34158 26496 34526 26497
rect 34746 26603 35114 26604
rect 34746 26569 35114 26603
rect 34746 26531 35114 26569
rect 34746 26497 35114 26531
rect 34746 26496 35114 26497
rect 35334 26603 35702 26604
rect 35334 26569 35702 26603
rect 35334 26531 35702 26569
rect 35334 26497 35702 26531
rect 35334 26496 35702 26497
rect 35922 26603 36290 26604
rect 35922 26569 36290 26603
rect 35922 26531 36290 26569
rect 35922 26497 36290 26531
rect 35922 26496 36290 26497
rect 36510 26603 36878 26604
rect 36510 26569 36878 26603
rect 36510 26531 36878 26569
rect 36510 26497 36878 26531
rect 36510 26496 36878 26497
rect 37098 26603 37466 26604
rect 37098 26569 37466 26603
rect 37098 26531 37466 26569
rect 37098 26497 37466 26531
rect 37098 26496 37466 26497
rect 37686 26603 38054 26604
rect 37686 26569 38054 26603
rect 37686 26531 38054 26569
rect 37686 26497 38054 26531
rect 37686 26496 38054 26497
rect 38274 26603 38642 26604
rect 38274 26569 38642 26603
rect 38274 26531 38642 26569
rect 38274 26497 38642 26531
rect 38274 26496 38642 26497
rect 10638 25603 11006 25604
rect 10638 25569 11006 25603
rect 10638 25531 11006 25569
rect 10638 25497 11006 25531
rect 10638 25496 11006 25497
rect 11226 25603 11594 25604
rect 11226 25569 11594 25603
rect 11226 25531 11594 25569
rect 11226 25497 11594 25531
rect 11226 25496 11594 25497
rect 11814 25603 12182 25604
rect 11814 25569 12182 25603
rect 11814 25531 12182 25569
rect 11814 25497 12182 25531
rect 11814 25496 12182 25497
rect 12402 25603 12770 25604
rect 12402 25569 12770 25603
rect 12402 25531 12770 25569
rect 12402 25497 12770 25531
rect 12402 25496 12770 25497
rect 12990 25603 13358 25604
rect 12990 25569 13358 25603
rect 12990 25531 13358 25569
rect 12990 25497 13358 25531
rect 12990 25496 13358 25497
rect 13578 25603 13946 25604
rect 13578 25569 13946 25603
rect 13578 25531 13946 25569
rect 13578 25497 13946 25531
rect 13578 25496 13946 25497
rect 14166 25603 14534 25604
rect 14166 25569 14534 25603
rect 14166 25531 14534 25569
rect 14166 25497 14534 25531
rect 14166 25496 14534 25497
rect 14754 25603 15122 25604
rect 14754 25569 15122 25603
rect 14754 25531 15122 25569
rect 14754 25497 15122 25531
rect 14754 25496 15122 25497
rect 15342 25603 15710 25604
rect 15342 25569 15710 25603
rect 15342 25531 15710 25569
rect 15342 25497 15710 25531
rect 15342 25496 15710 25497
rect 15930 25603 16298 25604
rect 15930 25569 16298 25603
rect 15930 25531 16298 25569
rect 15930 25497 16298 25531
rect 15930 25496 16298 25497
rect 16518 25603 16886 25604
rect 16518 25569 16886 25603
rect 16518 25531 16886 25569
rect 16518 25497 16886 25531
rect 16518 25496 16886 25497
rect 17106 25603 17474 25604
rect 17106 25569 17474 25603
rect 17106 25531 17474 25569
rect 17106 25497 17474 25531
rect 17106 25496 17474 25497
rect 17694 25603 18062 25604
rect 17694 25569 18062 25603
rect 17694 25531 18062 25569
rect 17694 25497 18062 25531
rect 17694 25496 18062 25497
rect 18282 25603 18650 25604
rect 18282 25569 18650 25603
rect 18282 25531 18650 25569
rect 18282 25497 18650 25531
rect 18282 25496 18650 25497
rect 18870 25603 19238 25604
rect 18870 25569 19238 25603
rect 18870 25531 19238 25569
rect 18870 25497 19238 25531
rect 18870 25496 19238 25497
rect 19458 25603 19826 25604
rect 19458 25569 19826 25603
rect 19458 25531 19826 25569
rect 19458 25497 19826 25531
rect 19458 25496 19826 25497
rect 20046 25603 20414 25604
rect 20046 25569 20414 25603
rect 20046 25531 20414 25569
rect 20046 25497 20414 25531
rect 20046 25496 20414 25497
rect 20634 25603 21002 25604
rect 20634 25569 21002 25603
rect 20634 25531 21002 25569
rect 20634 25497 21002 25531
rect 20634 25496 21002 25497
rect 21222 25603 21590 25604
rect 21222 25569 21590 25603
rect 21222 25531 21590 25569
rect 21222 25497 21590 25531
rect 21222 25496 21590 25497
rect 21810 25603 22178 25604
rect 21810 25569 22178 25603
rect 21810 25531 22178 25569
rect 21810 25497 22178 25531
rect 21810 25496 22178 25497
rect 22420 25496 22732 25604
rect 23020 25494 23318 25606
rect 23608 25603 23906 25606
rect 23608 25569 23906 25603
rect 23608 25531 23906 25569
rect 23608 25497 23906 25531
rect 23608 25494 23906 25497
rect 24196 25603 24494 25606
rect 24196 25569 24494 25603
rect 24196 25531 24494 25569
rect 24196 25497 24494 25531
rect 24196 25494 24494 25497
rect 24784 25603 25082 25606
rect 24784 25569 25082 25603
rect 24784 25531 25082 25569
rect 24784 25497 25082 25531
rect 24784 25494 25082 25497
rect 25372 25603 25670 25606
rect 25372 25569 25670 25603
rect 25372 25531 25670 25569
rect 25372 25497 25670 25531
rect 25372 25494 25670 25497
rect 25960 25603 26258 25606
rect 25960 25569 26258 25603
rect 25960 25531 26258 25569
rect 25960 25497 26258 25531
rect 25960 25494 26258 25497
rect 26548 25603 26846 25606
rect 26548 25569 26846 25603
rect 26548 25531 26846 25569
rect 26548 25497 26846 25531
rect 26548 25494 26846 25497
rect 27136 25603 27434 25606
rect 27136 25569 27434 25603
rect 27136 25531 27434 25569
rect 27136 25497 27434 25531
rect 27136 25494 27434 25497
rect 27724 25603 28022 25606
rect 27724 25569 28022 25603
rect 27724 25531 28022 25569
rect 27724 25497 28022 25531
rect 27724 25494 28022 25497
rect 28312 25603 28610 25606
rect 28312 25569 28610 25603
rect 28312 25531 28610 25569
rect 28312 25497 28610 25531
rect 28312 25494 28610 25497
rect 28900 25603 29198 25606
rect 28900 25569 29198 25603
rect 28900 25531 29198 25569
rect 28900 25497 29198 25531
rect 28900 25494 29198 25497
rect 29488 25603 29786 25606
rect 29488 25569 29786 25603
rect 29488 25531 29786 25569
rect 29488 25497 29786 25531
rect 29488 25494 29786 25497
rect 30076 25603 30374 25606
rect 30076 25569 30374 25603
rect 30076 25531 30374 25569
rect 30076 25497 30374 25531
rect 30076 25494 30374 25497
rect 30664 25603 30962 25606
rect 30664 25569 30962 25603
rect 30664 25531 30962 25569
rect 30664 25497 30962 25531
rect 30664 25494 30962 25497
rect 31252 25603 31550 25606
rect 31252 25569 31550 25603
rect 31252 25531 31550 25569
rect 31252 25497 31550 25531
rect 31252 25494 31550 25497
rect 31840 25603 32138 25606
rect 31840 25569 32138 25603
rect 31840 25531 32138 25569
rect 31840 25497 32138 25531
rect 31840 25494 32138 25497
rect 32428 25603 32726 25606
rect 32428 25569 32726 25603
rect 32428 25531 32726 25569
rect 32428 25497 32726 25531
rect 32428 25494 32726 25497
rect 33016 25603 33314 25606
rect 33016 25569 33314 25603
rect 33016 25531 33314 25569
rect 33016 25497 33314 25531
rect 33016 25494 33314 25497
rect 33604 25603 33902 25606
rect 33604 25569 33902 25603
rect 33604 25531 33902 25569
rect 33604 25497 33902 25531
rect 33604 25494 33902 25497
rect 34192 25603 34490 25606
rect 34192 25569 34490 25603
rect 34192 25531 34490 25569
rect 34192 25497 34490 25531
rect 34192 25494 34490 25497
rect 34780 25603 35078 25606
rect 34780 25569 35078 25603
rect 34780 25531 35078 25569
rect 34780 25497 35078 25531
rect 34780 25494 35078 25497
rect 35368 25603 35666 25606
rect 35368 25569 35666 25603
rect 35368 25531 35666 25569
rect 35368 25497 35666 25531
rect 35368 25494 35666 25497
rect 35956 25603 36254 25606
rect 35956 25569 36254 25603
rect 35956 25531 36254 25569
rect 35956 25497 36254 25531
rect 35956 25494 36254 25497
rect 36544 25603 36842 25606
rect 36544 25569 36842 25603
rect 36544 25531 36842 25569
rect 36544 25497 36842 25531
rect 36544 25494 36842 25497
rect 37132 25603 37430 25606
rect 37132 25569 37430 25603
rect 37132 25531 37430 25569
rect 37132 25497 37430 25531
rect 37132 25494 37430 25497
rect 37720 25603 38018 25606
rect 37720 25569 38018 25603
rect 37720 25531 38018 25569
rect 37720 25497 38018 25531
rect 37720 25494 38018 25497
rect 38308 25603 38606 25606
rect 38308 25569 38606 25603
rect 38308 25531 38606 25569
rect 38308 25497 38606 25531
rect 38308 25494 38606 25497
rect 3546 11952 5048 13186
rect 10658 24560 10988 24612
rect 11246 24603 11576 24612
rect 11246 24569 11576 24603
rect 11246 24560 11576 24569
rect 11834 24603 12164 24612
rect 11834 24569 12164 24603
rect 11834 24560 12164 24569
rect 12422 24603 12752 24612
rect 12422 24569 12752 24603
rect 12422 24560 12752 24569
rect 13010 24603 13340 24612
rect 13010 24569 13340 24603
rect 13010 24560 13340 24569
rect 13598 24603 13928 24612
rect 13598 24569 13928 24603
rect 13598 24560 13928 24569
rect 14186 24603 14516 24612
rect 14186 24569 14516 24603
rect 14186 24560 14516 24569
rect 14774 24603 15104 24612
rect 14774 24569 15104 24603
rect 14774 24560 15104 24569
rect 15362 24603 15692 24612
rect 15362 24569 15692 24603
rect 15362 24560 15692 24569
rect 15950 24603 16280 24612
rect 15950 24569 16280 24603
rect 15950 24560 16280 24569
rect 16538 24603 16868 24612
rect 16538 24569 16868 24603
rect 16538 24560 16868 24569
rect 17126 24603 17456 24612
rect 17126 24569 17456 24603
rect 17126 24560 17456 24569
rect 17714 24603 18044 24612
rect 17714 24569 18044 24603
rect 17714 24560 18044 24569
rect 18302 24603 18632 24612
rect 18302 24569 18632 24603
rect 18302 24560 18632 24569
rect 18890 24603 19220 24612
rect 18890 24569 19220 24603
rect 18890 24560 19220 24569
rect 19478 24603 19808 24612
rect 19478 24569 19808 24603
rect 19478 24560 19808 24569
rect 20066 24603 20396 24612
rect 20066 24569 20396 24603
rect 20066 24560 20396 24569
rect 20654 24603 20984 24612
rect 20654 24569 20984 24603
rect 20654 24560 20984 24569
rect 21242 24603 21572 24612
rect 21242 24569 21572 24603
rect 21242 24560 21572 24569
rect 21830 24603 22160 24612
rect 21830 24569 22160 24603
rect 21830 24560 22160 24569
rect 22416 24554 22736 24622
rect 23004 24603 23324 24622
rect 23004 24569 23324 24603
rect 23004 24554 23324 24569
rect 23592 24603 23912 24622
rect 23592 24569 23912 24603
rect 23592 24554 23912 24569
rect 24180 24603 24500 24622
rect 24180 24569 24500 24603
rect 24180 24554 24500 24569
rect 24768 24603 25088 24622
rect 24768 24569 25088 24603
rect 24768 24554 25088 24569
rect 25356 24603 25676 24622
rect 25356 24569 25676 24603
rect 25356 24554 25676 24569
rect 25944 24603 26264 24622
rect 25944 24569 26264 24603
rect 25944 24554 26264 24569
rect 26532 24603 26852 24622
rect 26532 24569 26852 24603
rect 26532 24554 26852 24569
rect 27120 24603 27440 24622
rect 27120 24569 27440 24603
rect 27120 24554 27440 24569
rect 27708 24603 28028 24622
rect 27708 24569 28028 24603
rect 27708 24554 28028 24569
rect 28296 24603 28616 24622
rect 28296 24569 28616 24603
rect 28296 24554 28616 24569
rect 28884 24603 29204 24622
rect 28884 24569 29204 24603
rect 28884 24554 29204 24569
rect 29472 24603 29792 24622
rect 29472 24569 29792 24603
rect 29472 24554 29792 24569
rect 30060 24603 30380 24622
rect 30060 24569 30380 24603
rect 30060 24554 30380 24569
rect 30648 24603 30968 24622
rect 30648 24569 30968 24603
rect 30648 24554 30968 24569
rect 31236 24603 31556 24622
rect 31236 24569 31556 24603
rect 31236 24554 31556 24569
rect 31824 24603 32144 24622
rect 31824 24569 32144 24603
rect 31824 24554 32144 24569
rect 32412 24603 32732 24622
rect 32412 24569 32732 24603
rect 32412 24554 32732 24569
rect 33000 24603 33320 24622
rect 33000 24569 33320 24603
rect 33000 24554 33320 24569
rect 33588 24603 33908 24622
rect 33588 24569 33908 24603
rect 33588 24554 33908 24569
rect 34176 24603 34496 24622
rect 34176 24569 34496 24603
rect 34176 24554 34496 24569
rect 34764 24603 35084 24622
rect 34764 24569 35084 24603
rect 34764 24554 35084 24569
rect 35352 24603 35672 24622
rect 35352 24569 35672 24603
rect 35352 24554 35672 24569
rect 35940 24603 36260 24622
rect 35940 24569 36260 24603
rect 35940 24554 36260 24569
rect 36528 24603 36848 24622
rect 36528 24569 36848 24603
rect 36528 24554 36848 24569
rect 37116 24603 37436 24622
rect 37116 24569 37436 24603
rect 37116 24554 37436 24569
rect 37704 24603 38024 24622
rect 37704 24569 38024 24603
rect 37704 24554 38024 24569
rect 38292 24603 38612 24622
rect 38292 24569 38612 24603
rect 38292 24554 38612 24569
rect 39582 22924 39860 23424
rect 37832 20906 38980 22370
rect 10482 12850 11158 12856
rect 44312 18676 45378 19484
rect 10482 12046 12288 12850
rect 10650 11144 10994 11196
rect 11238 11187 11582 11196
rect 11238 11153 11582 11187
rect 11238 11144 11582 11153
rect 11826 11187 12170 11196
rect 11826 11153 12170 11187
rect 11826 11144 12170 11153
rect 12414 11187 12758 11196
rect 12414 11153 12758 11187
rect 12414 11144 12758 11153
rect 13002 11187 13346 11196
rect 13002 11153 13346 11187
rect 13002 11144 13346 11153
rect 13590 11187 13934 11196
rect 13590 11153 13934 11187
rect 13590 11144 13934 11153
rect 14178 11187 14522 11196
rect 14178 11153 14522 11187
rect 14178 11144 14522 11153
rect 14766 11187 15110 11196
rect 14766 11153 15110 11187
rect 14766 11144 15110 11153
rect 15354 11187 15698 11196
rect 15354 11153 15698 11187
rect 15354 11144 15698 11153
rect 15942 11187 16286 11196
rect 15942 11153 16286 11187
rect 15942 11144 16286 11153
rect 16530 11187 16874 11196
rect 16530 11153 16874 11187
rect 16530 11144 16874 11153
rect 17118 11187 17462 11196
rect 17118 11153 17462 11187
rect 17118 11144 17462 11153
rect 17706 11187 18050 11196
rect 17706 11153 18050 11187
rect 17706 11144 18050 11153
rect 18294 11187 18638 11196
rect 18294 11153 18638 11187
rect 18294 11144 18638 11153
rect 18882 11187 19226 11196
rect 18882 11153 19226 11187
rect 18882 11144 19226 11153
rect 19470 11187 19814 11196
rect 19470 11153 19814 11187
rect 19470 11144 19814 11153
rect 20058 11187 20402 11196
rect 20058 11153 20402 11187
rect 20058 11144 20402 11153
rect 20646 11187 20990 11196
rect 20646 11153 20990 11187
rect 20646 11144 20990 11153
rect 21234 11187 21578 11196
rect 21234 11153 21578 11187
rect 21234 11144 21578 11153
rect 21822 11187 22166 11196
rect 21822 11153 22166 11187
rect 21822 11144 22166 11153
rect 22446 11138 22716 11196
rect 23020 11140 23318 11200
rect 23600 11136 23920 11200
rect 24178 11130 24512 11202
rect 24776 11130 25094 11212
rect 25360 11128 25698 11230
rect 25944 11126 26282 11228
rect 26532 11187 26870 11228
rect 26532 11153 26870 11187
rect 26532 11126 26870 11153
rect 27120 11187 27458 11228
rect 27120 11153 27458 11187
rect 27120 11126 27458 11153
rect 27708 11187 28046 11228
rect 27708 11153 28046 11187
rect 27708 11126 28046 11153
rect 28296 11187 28634 11228
rect 28296 11153 28634 11187
rect 28296 11126 28634 11153
rect 28884 11187 29222 11228
rect 28884 11153 29222 11187
rect 28884 11126 29222 11153
rect 29472 11187 29810 11228
rect 29472 11153 29810 11187
rect 29472 11126 29810 11153
rect 30060 11187 30398 11228
rect 30060 11153 30398 11187
rect 30060 11126 30398 11153
rect 30648 11187 30986 11228
rect 30648 11153 30986 11187
rect 30648 11126 30986 11153
rect 31236 11187 31574 11228
rect 31236 11153 31574 11187
rect 31236 11126 31574 11153
rect 31824 11187 32162 11228
rect 31824 11153 32162 11187
rect 31824 11126 32162 11153
rect 32412 11187 32750 11228
rect 32412 11153 32750 11187
rect 32412 11126 32750 11153
rect 33000 11187 33338 11228
rect 33000 11153 33338 11187
rect 33000 11126 33338 11153
rect 33588 11187 33926 11228
rect 33588 11153 33926 11187
rect 33588 11126 33926 11153
rect 34176 11187 34514 11228
rect 34176 11153 34514 11187
rect 34176 11126 34514 11153
rect 34764 11187 35102 11228
rect 34764 11153 35102 11187
rect 34764 11126 35102 11153
rect 35352 11187 35690 11228
rect 35352 11153 35690 11187
rect 35352 11126 35690 11153
rect 35940 11187 36278 11228
rect 35940 11153 36278 11187
rect 35940 11126 36278 11153
rect 36528 11187 36866 11228
rect 36528 11153 36866 11187
rect 36528 11126 36866 11153
rect 37116 11187 37454 11228
rect 37116 11153 37454 11187
rect 37116 11126 37454 11153
rect 37704 11187 38042 11228
rect 37704 11153 38042 11187
rect 37704 11126 38042 11153
rect 38292 11187 38630 11228
rect 38292 11153 38630 11187
rect 38292 11126 38630 11153
rect 10660 10148 10982 10266
rect 11248 10259 11570 10266
rect 11248 10225 11570 10259
rect 11248 10187 11570 10225
rect 11248 10153 11570 10187
rect 11248 10148 11570 10153
rect 11836 10259 12158 10266
rect 11836 10225 12158 10259
rect 11836 10187 12158 10225
rect 11836 10153 12158 10187
rect 11836 10148 12158 10153
rect 12424 10259 12746 10266
rect 12424 10225 12746 10259
rect 12424 10187 12746 10225
rect 12424 10153 12746 10187
rect 12424 10148 12746 10153
rect 13012 10259 13334 10266
rect 13012 10225 13334 10259
rect 13012 10187 13334 10225
rect 13012 10153 13334 10187
rect 13012 10148 13334 10153
rect 13600 10259 13922 10266
rect 13600 10225 13922 10259
rect 13600 10187 13922 10225
rect 13600 10153 13922 10187
rect 13600 10148 13922 10153
rect 14188 10259 14510 10266
rect 14188 10225 14510 10259
rect 14188 10187 14510 10225
rect 14188 10153 14510 10187
rect 14188 10148 14510 10153
rect 14776 10259 15098 10266
rect 14776 10225 15098 10259
rect 14776 10187 15098 10225
rect 14776 10153 15098 10187
rect 14776 10148 15098 10153
rect 15364 10259 15686 10266
rect 15364 10225 15686 10259
rect 15364 10187 15686 10225
rect 15364 10153 15686 10187
rect 15364 10148 15686 10153
rect 15952 10259 16274 10266
rect 15952 10225 16274 10259
rect 15952 10187 16274 10225
rect 15952 10153 16274 10187
rect 15952 10148 16274 10153
rect 16540 10259 16862 10266
rect 16540 10225 16862 10259
rect 16540 10187 16862 10225
rect 16540 10153 16862 10187
rect 16540 10148 16862 10153
rect 17128 10259 17450 10266
rect 17128 10225 17450 10259
rect 17128 10187 17450 10225
rect 17128 10153 17450 10187
rect 17128 10148 17450 10153
rect 17716 10259 18038 10266
rect 17716 10225 18038 10259
rect 17716 10187 18038 10225
rect 17716 10153 18038 10187
rect 17716 10148 18038 10153
rect 18304 10259 18626 10266
rect 18304 10225 18626 10259
rect 18304 10187 18626 10225
rect 18304 10153 18626 10187
rect 18304 10148 18626 10153
rect 18892 10259 19214 10266
rect 18892 10225 19214 10259
rect 18892 10187 19214 10225
rect 18892 10153 19214 10187
rect 18892 10148 19214 10153
rect 19480 10259 19802 10266
rect 19480 10225 19802 10259
rect 19480 10187 19802 10225
rect 19480 10153 19802 10187
rect 19480 10148 19802 10153
rect 20068 10259 20390 10266
rect 20068 10225 20390 10259
rect 20068 10187 20390 10225
rect 20068 10153 20390 10187
rect 20068 10148 20390 10153
rect 20656 10259 20978 10266
rect 20656 10225 20978 10259
rect 20656 10187 20978 10225
rect 20656 10153 20978 10187
rect 20656 10148 20978 10153
rect 21244 10259 21566 10266
rect 21244 10225 21566 10259
rect 21244 10187 21566 10225
rect 21244 10153 21566 10187
rect 21244 10148 21566 10153
rect 21832 10259 22154 10266
rect 21832 10225 22154 10259
rect 21832 10187 22154 10225
rect 21832 10153 22154 10187
rect 21832 10148 22154 10153
rect 22418 10146 22752 10266
rect 23006 10259 23340 10266
rect 23006 10225 23340 10259
rect 23006 10187 23340 10225
rect 23006 10153 23340 10187
rect 23006 10146 23340 10153
rect 23594 10259 23928 10266
rect 23594 10225 23928 10259
rect 23594 10187 23928 10225
rect 23594 10153 23928 10187
rect 23594 10146 23928 10153
rect 24182 10259 24516 10266
rect 24182 10225 24516 10259
rect 24182 10187 24516 10225
rect 24182 10153 24516 10187
rect 24182 10146 24516 10153
rect 24770 10259 25104 10266
rect 24770 10225 25104 10259
rect 24770 10187 25104 10225
rect 24770 10153 25104 10187
rect 24770 10146 25104 10153
rect 25358 10259 25692 10266
rect 25358 10225 25692 10259
rect 25358 10187 25692 10225
rect 25358 10153 25692 10187
rect 25358 10146 25692 10153
rect 25946 10259 26280 10266
rect 25946 10225 26280 10259
rect 25946 10187 26280 10225
rect 25946 10153 26280 10187
rect 25946 10146 26280 10153
rect 26534 10259 26868 10266
rect 26534 10225 26868 10259
rect 26534 10187 26868 10225
rect 26534 10153 26868 10187
rect 26534 10146 26868 10153
rect 27122 10259 27456 10266
rect 27122 10225 27456 10259
rect 27122 10187 27456 10225
rect 27122 10153 27456 10187
rect 27122 10146 27456 10153
rect 27710 10259 28044 10266
rect 27710 10225 28044 10259
rect 27710 10187 28044 10225
rect 27710 10153 28044 10187
rect 27710 10146 28044 10153
rect 28298 10259 28632 10266
rect 28298 10225 28632 10259
rect 28298 10187 28632 10225
rect 28298 10153 28632 10187
rect 28298 10146 28632 10153
rect 28886 10259 29220 10266
rect 28886 10225 29220 10259
rect 28886 10187 29220 10225
rect 28886 10153 29220 10187
rect 28886 10146 29220 10153
rect 29474 10259 29808 10266
rect 29474 10225 29808 10259
rect 29474 10187 29808 10225
rect 29474 10153 29808 10187
rect 29474 10146 29808 10153
rect 30062 10259 30396 10266
rect 30062 10225 30396 10259
rect 30062 10187 30396 10225
rect 30062 10153 30396 10187
rect 30062 10146 30396 10153
rect 30650 10259 30984 10266
rect 30650 10225 30984 10259
rect 30650 10187 30984 10225
rect 30650 10153 30984 10187
rect 30650 10146 30984 10153
rect 31238 10259 31572 10266
rect 31238 10225 31572 10259
rect 31238 10187 31572 10225
rect 31238 10153 31572 10187
rect 31238 10146 31572 10153
rect 31826 10259 32160 10266
rect 31826 10225 32160 10259
rect 31826 10187 32160 10225
rect 31826 10153 32160 10187
rect 31826 10146 32160 10153
rect 32414 10259 32748 10266
rect 32414 10225 32748 10259
rect 32414 10187 32748 10225
rect 32414 10153 32748 10187
rect 32414 10146 32748 10153
rect 33002 10259 33336 10266
rect 33002 10225 33336 10259
rect 33002 10187 33336 10225
rect 33002 10153 33336 10187
rect 33002 10146 33336 10153
rect 33590 10259 33924 10266
rect 33590 10225 33924 10259
rect 33590 10187 33924 10225
rect 33590 10153 33924 10187
rect 33590 10146 33924 10153
rect 34178 10259 34512 10266
rect 34178 10225 34512 10259
rect 34178 10187 34512 10225
rect 34178 10153 34512 10187
rect 34178 10146 34512 10153
rect 34766 10259 35100 10266
rect 34766 10225 35100 10259
rect 34766 10187 35100 10225
rect 34766 10153 35100 10187
rect 34766 10146 35100 10153
rect 35354 10259 35688 10266
rect 35354 10225 35688 10259
rect 35354 10187 35688 10225
rect 35354 10153 35688 10187
rect 35354 10146 35688 10153
rect 35942 10259 36276 10266
rect 35942 10225 36276 10259
rect 35942 10187 36276 10225
rect 35942 10153 36276 10187
rect 35942 10146 36276 10153
rect 36530 10259 36864 10266
rect 36530 10225 36864 10259
rect 36530 10187 36864 10225
rect 36530 10153 36864 10187
rect 36530 10146 36864 10153
rect 37118 10259 37452 10266
rect 37118 10225 37452 10259
rect 37118 10187 37452 10225
rect 37118 10153 37452 10187
rect 37118 10146 37452 10153
rect 37706 10259 38040 10266
rect 37706 10225 38040 10259
rect 37706 10187 38040 10225
rect 37706 10153 38040 10187
rect 37706 10146 38040 10153
rect 38294 10259 38628 10266
rect 38294 10225 38628 10259
rect 38294 10187 38628 10225
rect 38294 10153 38628 10187
rect 38294 10146 38628 10153
rect 10680 9259 10946 9276
rect 10680 9225 10946 9259
rect 10680 9187 10946 9225
rect 10680 9153 10946 9187
rect 10680 9128 10946 9153
rect 11268 9259 11534 9276
rect 11268 9225 11534 9259
rect 11268 9187 11534 9225
rect 11268 9153 11534 9187
rect 11268 9128 11534 9153
rect 11856 9259 12122 9276
rect 11856 9225 12122 9259
rect 11856 9187 12122 9225
rect 11856 9153 12122 9187
rect 11856 9128 12122 9153
rect 12444 9259 12710 9276
rect 12444 9225 12710 9259
rect 12444 9187 12710 9225
rect 12444 9153 12710 9187
rect 12444 9128 12710 9153
rect 13032 9259 13298 9276
rect 13032 9225 13298 9259
rect 13032 9187 13298 9225
rect 13032 9153 13298 9187
rect 13032 9128 13298 9153
rect 13620 9259 13886 9276
rect 13620 9225 13886 9259
rect 13620 9187 13886 9225
rect 13620 9153 13886 9187
rect 13620 9128 13886 9153
rect 14208 9259 14474 9276
rect 14208 9225 14474 9259
rect 14208 9187 14474 9225
rect 14208 9153 14474 9187
rect 14208 9128 14474 9153
rect 14796 9259 15062 9276
rect 14796 9225 15062 9259
rect 14796 9187 15062 9225
rect 14796 9153 15062 9187
rect 14796 9128 15062 9153
rect 15384 9259 15650 9276
rect 15384 9225 15650 9259
rect 15384 9187 15650 9225
rect 15384 9153 15650 9187
rect 15384 9128 15650 9153
rect 15972 9259 16238 9276
rect 15972 9225 16238 9259
rect 15972 9187 16238 9225
rect 15972 9153 16238 9187
rect 15972 9128 16238 9153
rect 16560 9259 16826 9276
rect 16560 9225 16826 9259
rect 16560 9187 16826 9225
rect 16560 9153 16826 9187
rect 16560 9128 16826 9153
rect 17148 9259 17414 9276
rect 17148 9225 17414 9259
rect 17148 9187 17414 9225
rect 17148 9153 17414 9187
rect 17148 9128 17414 9153
rect 17736 9259 18002 9276
rect 17736 9225 18002 9259
rect 17736 9187 18002 9225
rect 17736 9153 18002 9187
rect 17736 9128 18002 9153
rect 18324 9259 18590 9276
rect 18324 9225 18590 9259
rect 18324 9187 18590 9225
rect 18324 9153 18590 9187
rect 18324 9128 18590 9153
rect 18912 9259 19178 9276
rect 18912 9225 19178 9259
rect 18912 9187 19178 9225
rect 18912 9153 19178 9187
rect 18912 9128 19178 9153
rect 19500 9259 19766 9276
rect 19500 9225 19766 9259
rect 19500 9187 19766 9225
rect 19500 9153 19766 9187
rect 19500 9128 19766 9153
rect 20088 9259 20354 9276
rect 20088 9225 20354 9259
rect 20088 9187 20354 9225
rect 20088 9153 20354 9187
rect 20088 9128 20354 9153
rect 20676 9259 20942 9276
rect 20676 9225 20942 9259
rect 20676 9187 20942 9225
rect 20676 9153 20942 9187
rect 20676 9128 20942 9153
rect 21264 9259 21530 9276
rect 21264 9225 21530 9259
rect 21264 9187 21530 9225
rect 21264 9153 21530 9187
rect 21264 9128 21530 9153
rect 21852 9259 22118 9276
rect 21852 9225 22118 9259
rect 21852 9187 22118 9225
rect 21852 9153 22118 9187
rect 21852 9128 22118 9153
rect 22418 9126 22750 9286
rect 23006 9259 23338 9286
rect 23006 9225 23338 9259
rect 23006 9187 23338 9225
rect 23006 9153 23338 9187
rect 23006 9126 23338 9153
rect 23594 9259 23926 9286
rect 23594 9225 23926 9259
rect 23594 9187 23926 9225
rect 23594 9153 23926 9187
rect 23594 9126 23926 9153
rect 24182 9259 24514 9286
rect 24182 9225 24514 9259
rect 24182 9187 24514 9225
rect 24182 9153 24514 9187
rect 24182 9126 24514 9153
rect 24770 9259 25102 9286
rect 24770 9225 25102 9259
rect 24770 9187 25102 9225
rect 24770 9153 25102 9187
rect 24770 9126 25102 9153
rect 25358 9259 25690 9286
rect 25358 9225 25690 9259
rect 25358 9187 25690 9225
rect 25358 9153 25690 9187
rect 25358 9126 25690 9153
rect 25946 9259 26278 9286
rect 25946 9225 26278 9259
rect 25946 9187 26278 9225
rect 25946 9153 26278 9187
rect 25946 9126 26278 9153
rect 26534 9259 26866 9286
rect 26534 9225 26866 9259
rect 26534 9187 26866 9225
rect 26534 9153 26866 9187
rect 26534 9126 26866 9153
rect 27122 9259 27454 9286
rect 27122 9225 27454 9259
rect 27122 9187 27454 9225
rect 27122 9153 27454 9187
rect 27122 9126 27454 9153
rect 27710 9259 28042 9286
rect 27710 9225 28042 9259
rect 27710 9187 28042 9225
rect 27710 9153 28042 9187
rect 27710 9126 28042 9153
rect 28298 9259 28630 9286
rect 28298 9225 28630 9259
rect 28298 9187 28630 9225
rect 28298 9153 28630 9187
rect 28298 9126 28630 9153
rect 28886 9259 29218 9286
rect 28886 9225 29218 9259
rect 28886 9187 29218 9225
rect 28886 9153 29218 9187
rect 28886 9126 29218 9153
rect 29474 9259 29806 9286
rect 29474 9225 29806 9259
rect 29474 9187 29806 9225
rect 29474 9153 29806 9187
rect 29474 9126 29806 9153
rect 30062 9259 30394 9286
rect 30062 9225 30394 9259
rect 30062 9187 30394 9225
rect 30062 9153 30394 9187
rect 30062 9126 30394 9153
rect 30650 9259 30982 9286
rect 30650 9225 30982 9259
rect 30650 9187 30982 9225
rect 30650 9153 30982 9187
rect 30650 9126 30982 9153
rect 31238 9259 31570 9286
rect 31238 9225 31570 9259
rect 31238 9187 31570 9225
rect 31238 9153 31570 9187
rect 31238 9126 31570 9153
rect 31826 9259 32158 9286
rect 31826 9225 32158 9259
rect 31826 9187 32158 9225
rect 31826 9153 32158 9187
rect 31826 9126 32158 9153
rect 32414 9259 32746 9286
rect 32414 9225 32746 9259
rect 32414 9187 32746 9225
rect 32414 9153 32746 9187
rect 32414 9126 32746 9153
rect 33002 9259 33334 9286
rect 33002 9225 33334 9259
rect 33002 9187 33334 9225
rect 33002 9153 33334 9187
rect 33002 9126 33334 9153
rect 33590 9259 33922 9286
rect 33590 9225 33922 9259
rect 33590 9187 33922 9225
rect 33590 9153 33922 9187
rect 33590 9126 33922 9153
rect 34178 9259 34510 9286
rect 34178 9225 34510 9259
rect 34178 9187 34510 9225
rect 34178 9153 34510 9187
rect 34178 9126 34510 9153
rect 34766 9259 35098 9286
rect 34766 9225 35098 9259
rect 34766 9187 35098 9225
rect 34766 9153 35098 9187
rect 34766 9126 35098 9153
rect 35354 9259 35686 9286
rect 35354 9225 35686 9259
rect 35354 9187 35686 9225
rect 35354 9153 35686 9187
rect 35354 9126 35686 9153
rect 35942 9259 36274 9286
rect 35942 9225 36274 9259
rect 35942 9187 36274 9225
rect 35942 9153 36274 9187
rect 35942 9126 36274 9153
rect 36530 9259 36862 9286
rect 36530 9225 36862 9259
rect 36530 9187 36862 9225
rect 36530 9153 36862 9187
rect 36530 9126 36862 9153
rect 37118 9259 37450 9286
rect 37118 9225 37450 9259
rect 37118 9187 37450 9225
rect 37118 9153 37450 9187
rect 37118 9126 37450 9153
rect 37706 9259 38038 9286
rect 37706 9225 38038 9259
rect 37706 9187 38038 9225
rect 37706 9153 38038 9187
rect 37706 9126 38038 9153
rect 38294 9259 38626 9286
rect 38294 9225 38626 9259
rect 38294 9187 38626 9225
rect 38294 9153 38626 9187
rect 38294 9126 38626 9153
rect 10666 8208 10984 8276
rect 11254 8259 11572 8276
rect 11254 8225 11572 8259
rect 11254 8208 11572 8225
rect 11842 8259 12160 8276
rect 11842 8225 12160 8259
rect 11842 8208 12160 8225
rect 12430 8259 12748 8276
rect 12430 8225 12748 8259
rect 12430 8208 12748 8225
rect 13018 8259 13336 8276
rect 13018 8225 13336 8259
rect 13018 8208 13336 8225
rect 13606 8259 13924 8276
rect 13606 8225 13924 8259
rect 13606 8208 13924 8225
rect 14194 8259 14512 8276
rect 14194 8225 14512 8259
rect 14194 8208 14512 8225
rect 14782 8259 15100 8276
rect 14782 8225 15100 8259
rect 14782 8208 15100 8225
rect 15370 8259 15688 8276
rect 15370 8225 15688 8259
rect 15370 8208 15688 8225
rect 15958 8259 16276 8276
rect 15958 8225 16276 8259
rect 15958 8208 16276 8225
rect 16546 8259 16864 8276
rect 16546 8225 16864 8259
rect 16546 8208 16864 8225
rect 17134 8259 17452 8276
rect 17134 8225 17452 8259
rect 17134 8208 17452 8225
rect 17722 8259 18040 8276
rect 17722 8225 18040 8259
rect 17722 8208 18040 8225
rect 18310 8259 18628 8276
rect 18310 8225 18628 8259
rect 18310 8208 18628 8225
rect 18898 8259 19216 8276
rect 18898 8225 19216 8259
rect 18898 8208 19216 8225
rect 19486 8259 19804 8276
rect 19486 8225 19804 8259
rect 19486 8208 19804 8225
rect 20074 8259 20392 8276
rect 20074 8225 20392 8259
rect 20074 8208 20392 8225
rect 20662 8259 20980 8276
rect 20662 8225 20980 8259
rect 20662 8208 20980 8225
rect 21250 8259 21568 8276
rect 21250 8225 21568 8259
rect 21250 8208 21568 8225
rect 21838 8259 22156 8276
rect 21838 8225 22156 8259
rect 21838 8208 22156 8225
rect 22434 8196 22712 8274
rect 23022 8259 23300 8274
rect 23022 8225 23300 8259
rect 23022 8196 23300 8225
rect 23610 8259 23888 8274
rect 23610 8225 23888 8259
rect 23610 8196 23888 8225
rect 24198 8259 24476 8274
rect 24198 8225 24476 8259
rect 24198 8196 24476 8225
rect 24786 8259 25064 8274
rect 24786 8225 25064 8259
rect 24786 8196 25064 8225
rect 25374 8259 25652 8274
rect 25374 8225 25652 8259
rect 25374 8196 25652 8225
rect 25962 8259 26240 8274
rect 25962 8225 26240 8259
rect 25962 8196 26240 8225
rect 26550 8259 26828 8274
rect 26550 8225 26828 8259
rect 26550 8196 26828 8225
rect 27138 8259 27416 8274
rect 27138 8225 27416 8259
rect 27138 8196 27416 8225
rect 27726 8259 28004 8274
rect 27726 8225 28004 8259
rect 27726 8196 28004 8225
rect 28314 8259 28592 8274
rect 28314 8225 28592 8259
rect 28314 8196 28592 8225
rect 28902 8259 29180 8274
rect 28902 8225 29180 8259
rect 28902 8196 29180 8225
rect 29490 8259 29768 8274
rect 29490 8225 29768 8259
rect 29490 8196 29768 8225
rect 30078 8259 30356 8274
rect 30078 8225 30356 8259
rect 30078 8196 30356 8225
rect 30666 8259 30944 8274
rect 30666 8225 30944 8259
rect 30666 8196 30944 8225
rect 31254 8259 31532 8274
rect 31254 8225 31532 8259
rect 31254 8196 31532 8225
rect 31842 8259 32120 8274
rect 31842 8225 32120 8259
rect 31842 8196 32120 8225
rect 32430 8259 32708 8274
rect 32430 8225 32708 8259
rect 32430 8196 32708 8225
rect 33018 8259 33296 8274
rect 33018 8225 33296 8259
rect 33018 8196 33296 8225
rect 33606 8259 33884 8274
rect 33606 8225 33884 8259
rect 33606 8196 33884 8225
rect 34194 8259 34472 8274
rect 34194 8225 34472 8259
rect 34194 8196 34472 8225
rect 34782 8259 35060 8274
rect 34782 8225 35060 8259
rect 34782 8196 35060 8225
rect 35370 8259 35648 8274
rect 35370 8225 35648 8259
rect 35370 8196 35648 8225
rect 35958 8259 36236 8274
rect 35958 8225 36236 8259
rect 35958 8196 36236 8225
rect 36546 8259 36824 8274
rect 36546 8225 36824 8259
rect 36546 8196 36824 8225
rect 37134 8259 37412 8274
rect 37134 8225 37412 8259
rect 37134 8196 37412 8225
rect 37722 8259 38000 8274
rect 37722 8225 38000 8259
rect 37722 8196 38000 8225
rect 38310 8259 38588 8274
rect 38310 8225 38588 8259
rect 38310 8196 38588 8225
rect 44380 6144 45446 6952
rect 6278 3996 7030 4988
<< metal2 >>
rect 10622 27552 11022 27558
rect 11210 27552 11610 27558
rect 11798 27552 12198 27558
rect 12386 27552 12786 27558
rect 12974 27552 13374 27558
rect 13562 27552 13962 27558
rect 14150 27552 14550 27558
rect 14738 27552 15138 27558
rect 15326 27552 15726 27558
rect 15914 27552 16314 27558
rect 16502 27552 16902 27558
rect 17090 27552 17490 27558
rect 17678 27552 18078 27558
rect 18266 27552 18666 27558
rect 18854 27552 19254 27558
rect 19442 27552 19842 27558
rect 20030 27552 20430 27558
rect 20618 27552 21018 27558
rect 21206 27552 21606 27558
rect 10612 27548 38650 27552
rect 10612 27490 10622 27548
rect 11022 27490 11210 27548
rect 11610 27490 11798 27548
rect 12198 27490 12386 27548
rect 12786 27490 12974 27548
rect 13374 27490 13562 27548
rect 13962 27490 14150 27548
rect 14550 27490 14738 27548
rect 15138 27490 15326 27548
rect 15726 27490 15914 27548
rect 16314 27490 16502 27548
rect 16902 27490 17090 27548
rect 17490 27490 17678 27548
rect 18078 27490 18266 27548
rect 18666 27490 18854 27548
rect 19254 27490 19442 27548
rect 19842 27490 20030 27548
rect 20430 27490 20618 27548
rect 21018 27490 21206 27548
rect 21606 27542 38650 27548
rect 21606 27490 21802 27542
rect 10612 27486 21802 27490
rect 22178 27488 22398 27542
rect 22766 27488 22986 27542
rect 23354 27488 23574 27542
rect 23942 27488 24162 27542
rect 24530 27488 24750 27542
rect 25118 27488 25338 27542
rect 25706 27488 25926 27542
rect 26294 27488 26514 27542
rect 26882 27488 27102 27542
rect 27470 27488 27690 27542
rect 28058 27488 28278 27542
rect 28646 27488 28866 27542
rect 29234 27488 29454 27542
rect 29822 27488 30042 27542
rect 30410 27488 30630 27542
rect 30998 27488 31218 27542
rect 31586 27488 31806 27542
rect 32174 27488 32394 27542
rect 32762 27488 32982 27542
rect 33350 27488 33570 27542
rect 33938 27488 34158 27542
rect 34526 27488 34746 27542
rect 35114 27488 35334 27542
rect 35702 27488 35922 27542
rect 36290 27488 36510 27542
rect 36878 27488 37098 27542
rect 37466 27488 37686 27542
rect 38054 27488 38274 27542
rect 38642 27488 38650 27542
rect 22178 27486 38650 27488
rect 10612 27480 38650 27486
rect 21802 27476 22178 27480
rect 22398 27478 22766 27480
rect 22986 27478 23354 27480
rect 23574 27478 23942 27480
rect 24162 27478 24530 27480
rect 24750 27478 25118 27480
rect 25338 27478 25706 27480
rect 25926 27478 26294 27480
rect 26514 27478 26882 27480
rect 27102 27478 27470 27480
rect 27690 27478 28058 27480
rect 28278 27478 28646 27480
rect 28866 27478 29234 27480
rect 29454 27478 29822 27480
rect 30042 27478 30410 27480
rect 30630 27478 30998 27480
rect 31218 27478 31586 27480
rect 31806 27478 32174 27480
rect 32394 27478 32762 27480
rect 32982 27478 33350 27480
rect 33570 27478 33938 27480
rect 34158 27478 34526 27480
rect 34746 27478 35114 27480
rect 35334 27478 35702 27480
rect 35922 27478 36290 27480
rect 36510 27478 36878 27480
rect 37098 27478 37466 27480
rect 37686 27478 38054 27480
rect 38274 27478 38650 27480
rect 10436 26604 38650 26614
rect 10436 26490 10638 26604
rect 11006 26490 11226 26604
rect 11594 26490 11814 26604
rect 12182 26490 12402 26604
rect 12770 26490 12990 26604
rect 13358 26490 13578 26604
rect 13946 26490 14166 26604
rect 14534 26490 14754 26604
rect 15122 26490 15342 26604
rect 15710 26490 15930 26604
rect 16298 26490 16518 26604
rect 16886 26490 17106 26604
rect 17474 26490 17694 26604
rect 18062 26490 18282 26604
rect 18650 26490 18870 26604
rect 19238 26490 19458 26604
rect 19826 26490 20046 26604
rect 20414 26490 20634 26604
rect 21002 26490 21222 26604
rect 21590 26490 21810 26604
rect 22178 26496 22398 26604
rect 22766 26496 22986 26604
rect 23354 26496 23574 26604
rect 23942 26496 24162 26604
rect 24530 26496 24750 26604
rect 25118 26496 25338 26604
rect 25706 26496 25926 26604
rect 26294 26496 26514 26604
rect 26882 26496 27102 26604
rect 27470 26496 27690 26604
rect 28058 26496 28278 26604
rect 28646 26496 28866 26604
rect 29234 26496 29454 26604
rect 29822 26496 30042 26604
rect 30410 26496 30630 26604
rect 30998 26496 31218 26604
rect 31586 26496 31806 26604
rect 32174 26496 32394 26604
rect 32762 26496 32982 26604
rect 33350 26496 33570 26604
rect 33938 26496 34158 26604
rect 34526 26496 34746 26604
rect 35114 26496 35334 26604
rect 35702 26496 35922 26604
rect 36290 26496 36510 26604
rect 36878 26496 37098 26604
rect 37466 26496 37686 26604
rect 38054 26496 38274 26604
rect 38642 26496 38650 26604
rect 22178 26490 38650 26496
rect 10436 26480 38650 26490
rect 10638 25606 38650 25620
rect 10638 25604 23020 25606
rect 11006 25496 11226 25604
rect 11594 25496 11814 25604
rect 12182 25496 12402 25604
rect 12770 25496 12990 25604
rect 13358 25496 13578 25604
rect 13946 25496 14166 25604
rect 14534 25496 14754 25604
rect 15122 25496 15342 25604
rect 15710 25496 15930 25604
rect 16298 25496 16518 25604
rect 16886 25496 17106 25604
rect 17474 25496 17694 25604
rect 18062 25496 18282 25604
rect 18650 25496 18870 25604
rect 19238 25496 19458 25604
rect 19826 25496 20046 25604
rect 20414 25496 20634 25604
rect 21002 25496 21222 25604
rect 21590 25496 21810 25604
rect 22178 25496 22420 25604
rect 22732 25496 23020 25604
rect 10638 25494 23020 25496
rect 23318 25494 23608 25606
rect 23906 25494 24196 25606
rect 24494 25494 24784 25606
rect 25082 25494 25372 25606
rect 25670 25494 25960 25606
rect 26258 25494 26548 25606
rect 26846 25494 27136 25606
rect 27434 25494 27724 25606
rect 28022 25494 28312 25606
rect 28610 25494 28900 25606
rect 29198 25494 29488 25606
rect 29786 25494 30076 25606
rect 30374 25494 30664 25606
rect 30962 25494 31252 25606
rect 31550 25494 31840 25606
rect 32138 25494 32428 25606
rect 32726 25494 33016 25606
rect 33314 25494 33604 25606
rect 33902 25494 34192 25606
rect 34490 25494 34780 25606
rect 35078 25494 35368 25606
rect 35666 25494 35956 25606
rect 36254 25494 36544 25606
rect 36842 25494 37132 25606
rect 37430 25494 37720 25606
rect 38018 25494 38308 25606
rect 38606 25494 38650 25606
rect 10638 25486 38650 25494
rect 23020 25484 23318 25486
rect 23608 25484 23906 25486
rect 24196 25484 24494 25486
rect 24784 25484 25082 25486
rect 25372 25484 25670 25486
rect 25960 25484 26258 25486
rect 26548 25484 26846 25486
rect 27136 25484 27434 25486
rect 27724 25484 28022 25486
rect 28312 25484 28610 25486
rect 28900 25484 29198 25486
rect 29488 25484 29786 25486
rect 30076 25484 30374 25486
rect 30664 25484 30962 25486
rect 31252 25484 31550 25486
rect 31840 25484 32138 25486
rect 32428 25484 32726 25486
rect 33016 25484 33314 25486
rect 33604 25484 33902 25486
rect 34192 25484 34490 25486
rect 34780 25484 35078 25486
rect 35368 25484 35666 25486
rect 35956 25484 36254 25486
rect 36544 25484 36842 25486
rect 37132 25484 37430 25486
rect 37720 25484 38018 25486
rect 38308 25484 38606 25486
rect 10638 24622 38650 24638
rect 10638 24612 22416 24622
rect 10638 24560 10658 24612
rect 10988 24560 11246 24612
rect 11576 24560 11834 24612
rect 12164 24560 12422 24612
rect 12752 24560 13010 24612
rect 13340 24560 13598 24612
rect 13928 24560 14186 24612
rect 14516 24560 14774 24612
rect 15104 24560 15362 24612
rect 15692 24560 15950 24612
rect 16280 24560 16538 24612
rect 16868 24560 17126 24612
rect 17456 24560 17714 24612
rect 18044 24560 18302 24612
rect 18632 24560 18890 24612
rect 19220 24560 19478 24612
rect 19808 24560 20066 24612
rect 20396 24560 20654 24612
rect 20984 24560 21242 24612
rect 21572 24560 21830 24612
rect 22160 24560 22416 24612
rect 10638 24554 22416 24560
rect 22736 24554 23004 24622
rect 23324 24554 23592 24622
rect 23912 24554 24180 24622
rect 24500 24554 24768 24622
rect 25088 24554 25356 24622
rect 25676 24554 25944 24622
rect 26264 24554 26532 24622
rect 26852 24554 27120 24622
rect 27440 24554 27708 24622
rect 28028 24554 28296 24622
rect 28616 24554 28884 24622
rect 29204 24554 29472 24622
rect 29792 24554 30060 24622
rect 30380 24554 30648 24622
rect 30968 24554 31236 24622
rect 31556 24554 31824 24622
rect 32144 24554 32412 24622
rect 32732 24554 33000 24622
rect 33320 24554 33588 24622
rect 33908 24554 34176 24622
rect 34496 24554 34764 24622
rect 35084 24554 35352 24622
rect 35672 24554 35940 24622
rect 36260 24554 36528 24622
rect 36848 24554 37116 24622
rect 37436 24554 37704 24622
rect 38024 24554 38292 24622
rect 38612 24554 38650 24622
rect 10638 24548 38650 24554
rect 22416 24544 22736 24548
rect 23004 24544 23324 24548
rect 23592 24544 23912 24548
rect 24180 24544 24500 24548
rect 24768 24544 25088 24548
rect 25356 24544 25676 24548
rect 25944 24544 26264 24548
rect 26532 24544 26852 24548
rect 27120 24544 27440 24548
rect 27708 24544 28028 24548
rect 28296 24544 28616 24548
rect 28884 24544 29204 24548
rect 29472 24544 29792 24548
rect 30060 24544 30380 24548
rect 30648 24544 30968 24548
rect 31236 24544 31556 24548
rect 31824 24544 32144 24548
rect 32412 24544 32732 24548
rect 33000 24544 33320 24548
rect 33588 24544 33908 24548
rect 34176 24544 34496 24548
rect 34764 24544 35084 24548
rect 35352 24544 35672 24548
rect 35940 24544 36260 24548
rect 36528 24544 36848 24548
rect 37116 24544 37436 24548
rect 37704 24544 38024 24548
rect 38292 24544 38612 24548
rect 39582 23424 39860 23434
rect 26390 22924 39582 23424
rect 39582 22914 39860 22924
rect 37832 22370 38980 22380
rect 37832 20896 38980 20906
rect 22888 19020 23128 19866
rect 44312 19484 45378 19494
rect 30754 19020 30924 19324
rect 22888 18676 44312 19020
rect 22888 18672 45378 18676
rect 44312 18666 45378 18672
rect 3546 13186 5048 13196
rect 5048 12860 11210 12882
rect 5048 12856 12288 12860
rect 5048 12046 10482 12856
rect 11158 12850 12288 12856
rect 5048 12036 12288 12046
rect 5048 12014 11210 12036
rect 3546 11942 5048 11952
rect 10624 11230 38642 11240
rect 10624 11212 25360 11230
rect 10624 11202 24776 11212
rect 10624 11200 24178 11202
rect 10624 11196 23020 11200
rect 10624 11144 10650 11196
rect 10994 11144 11238 11196
rect 11582 11144 11826 11196
rect 12170 11144 12414 11196
rect 12758 11144 13002 11196
rect 13346 11144 13590 11196
rect 13934 11144 14178 11196
rect 14522 11144 14766 11196
rect 15110 11144 15354 11196
rect 15698 11144 15942 11196
rect 16286 11144 16530 11196
rect 16874 11144 17118 11196
rect 17462 11144 17706 11196
rect 18050 11144 18294 11196
rect 18638 11144 18882 11196
rect 19226 11144 19470 11196
rect 19814 11144 20058 11196
rect 20402 11144 20646 11196
rect 20990 11144 21234 11196
rect 21578 11144 21822 11196
rect 22166 11144 22446 11196
rect 10624 11138 22446 11144
rect 22716 11140 23020 11196
rect 23318 11140 23600 11200
rect 22716 11138 23600 11140
rect 10624 11136 23600 11138
rect 23920 11136 24178 11200
rect 10624 11134 24178 11136
rect 22446 11128 22716 11134
rect 23020 11130 23318 11134
rect 23600 11126 23920 11134
rect 24512 11134 24776 11202
rect 24178 11120 24512 11130
rect 25094 11134 25360 11212
rect 24776 11120 25094 11130
rect 25698 11228 38642 11230
rect 25698 11134 25944 11228
rect 25360 11118 25698 11128
rect 26282 11134 26532 11228
rect 25944 11116 26282 11126
rect 26870 11134 27120 11228
rect 26532 11116 26870 11126
rect 27458 11134 27708 11228
rect 27120 11116 27458 11126
rect 28046 11134 28296 11228
rect 27708 11116 28046 11126
rect 28634 11134 28884 11228
rect 28296 11116 28634 11126
rect 29222 11134 29472 11228
rect 28884 11116 29222 11126
rect 29810 11134 30060 11228
rect 29472 11116 29810 11126
rect 30398 11134 30648 11228
rect 30060 11116 30398 11126
rect 30986 11134 31236 11228
rect 30648 11116 30986 11126
rect 31574 11134 31824 11228
rect 31236 11116 31574 11126
rect 32162 11134 32412 11228
rect 31824 11116 32162 11126
rect 32750 11134 33000 11228
rect 32412 11116 32750 11126
rect 33338 11134 33588 11228
rect 33000 11116 33338 11126
rect 33926 11134 34176 11228
rect 33588 11116 33926 11126
rect 34514 11134 34764 11228
rect 34176 11116 34514 11126
rect 35102 11134 35352 11228
rect 34764 11116 35102 11126
rect 35690 11134 35940 11228
rect 35352 11116 35690 11126
rect 36278 11134 36528 11228
rect 35940 11116 36278 11126
rect 36866 11134 37116 11228
rect 36528 11116 36866 11126
rect 37454 11134 37704 11228
rect 37116 11116 37454 11126
rect 38042 11134 38292 11228
rect 37704 11116 38042 11126
rect 38630 11134 38642 11228
rect 38292 11116 38630 11126
rect 10342 10266 38642 10284
rect 10342 10148 10660 10266
rect 10982 10148 11248 10266
rect 11570 10148 11836 10266
rect 12158 10148 12424 10266
rect 12746 10148 13012 10266
rect 13334 10148 13600 10266
rect 13922 10148 14188 10266
rect 14510 10148 14776 10266
rect 15098 10148 15364 10266
rect 15686 10148 15952 10266
rect 16274 10148 16540 10266
rect 16862 10148 17128 10266
rect 17450 10148 17716 10266
rect 18038 10148 18304 10266
rect 18626 10148 18892 10266
rect 19214 10148 19480 10266
rect 19802 10148 20068 10266
rect 20390 10148 20656 10266
rect 20978 10148 21244 10266
rect 21566 10148 21832 10266
rect 22154 10148 22418 10266
rect 10342 10146 22418 10148
rect 22752 10146 23006 10266
rect 23340 10146 23594 10266
rect 23928 10146 24182 10266
rect 24516 10146 24770 10266
rect 25104 10146 25358 10266
rect 25692 10146 25946 10266
rect 26280 10146 26534 10266
rect 26868 10146 27122 10266
rect 27456 10146 27710 10266
rect 28044 10146 28298 10266
rect 28632 10146 28886 10266
rect 29220 10146 29474 10266
rect 29808 10146 30062 10266
rect 30396 10146 30650 10266
rect 30984 10146 31238 10266
rect 31572 10146 31826 10266
rect 32160 10146 32414 10266
rect 32748 10146 33002 10266
rect 33336 10146 33590 10266
rect 33924 10146 34178 10266
rect 34512 10146 34766 10266
rect 35100 10146 35354 10266
rect 35688 10146 35942 10266
rect 36276 10146 36530 10266
rect 36864 10146 37118 10266
rect 37452 10146 37706 10266
rect 38040 10146 38294 10266
rect 38628 10146 38642 10266
rect 10342 10136 38642 10146
rect 10668 9286 38642 9300
rect 10668 9276 22418 9286
rect 10668 9128 10680 9276
rect 10946 9128 11268 9276
rect 11534 9128 11856 9276
rect 12122 9128 12444 9276
rect 12710 9128 13032 9276
rect 13298 9128 13620 9276
rect 13886 9128 14208 9276
rect 14474 9128 14796 9276
rect 15062 9128 15384 9276
rect 15650 9128 15972 9276
rect 16238 9128 16560 9276
rect 16826 9128 17148 9276
rect 17414 9128 17736 9276
rect 18002 9128 18324 9276
rect 18590 9128 18912 9276
rect 19178 9128 19500 9276
rect 19766 9128 20088 9276
rect 20354 9128 20676 9276
rect 20942 9128 21264 9276
rect 21530 9128 21852 9276
rect 22118 9128 22418 9276
rect 10668 9126 22418 9128
rect 22750 9126 23006 9286
rect 23338 9126 23594 9286
rect 23926 9126 24182 9286
rect 24514 9126 24770 9286
rect 25102 9126 25358 9286
rect 25690 9126 25946 9286
rect 26278 9126 26534 9286
rect 26866 9126 27122 9286
rect 27454 9126 27710 9286
rect 28042 9126 28298 9286
rect 28630 9126 28886 9286
rect 29218 9126 29474 9286
rect 29806 9126 30062 9286
rect 30394 9126 30650 9286
rect 30982 9126 31238 9286
rect 31570 9126 31826 9286
rect 32158 9126 32414 9286
rect 32746 9126 33002 9286
rect 33334 9126 33590 9286
rect 33922 9126 34178 9286
rect 34510 9126 34766 9286
rect 35098 9126 35354 9286
rect 35686 9126 35942 9286
rect 36274 9126 36530 9286
rect 36862 9126 37118 9286
rect 37450 9126 37706 9286
rect 38038 9126 38294 9286
rect 38626 9126 38642 9286
rect 10668 9110 38642 9126
rect 10658 8276 38642 8286
rect 10658 8208 10666 8276
rect 10984 8208 11254 8276
rect 11572 8208 11842 8276
rect 12160 8208 12430 8276
rect 12748 8208 13018 8276
rect 13336 8208 13606 8276
rect 13924 8208 14194 8276
rect 14512 8208 14782 8276
rect 15100 8208 15370 8276
rect 15688 8208 15958 8276
rect 16276 8208 16546 8276
rect 16864 8208 17134 8276
rect 17452 8208 17722 8276
rect 18040 8208 18310 8276
rect 18628 8208 18898 8276
rect 19216 8208 19486 8276
rect 19804 8208 20074 8276
rect 20392 8208 20662 8276
rect 20980 8208 21250 8276
rect 21568 8208 21838 8276
rect 22156 8274 38642 8276
rect 22156 8208 22434 8274
rect 10658 8196 22434 8208
rect 22712 8196 23022 8274
rect 23300 8196 23610 8274
rect 23888 8196 24198 8274
rect 24476 8196 24786 8274
rect 25064 8196 25374 8274
rect 25652 8196 25962 8274
rect 26240 8196 26550 8274
rect 26828 8196 27138 8274
rect 27416 8196 27726 8274
rect 28004 8196 28314 8274
rect 28592 8196 28902 8274
rect 29180 8196 29490 8274
rect 29768 8196 30078 8274
rect 30356 8196 30666 8274
rect 30944 8196 31254 8274
rect 31532 8196 31842 8274
rect 32120 8196 32430 8274
rect 32708 8196 33018 8274
rect 33296 8196 33606 8274
rect 33884 8196 34194 8274
rect 34472 8196 34782 8274
rect 35060 8196 35370 8274
rect 35648 8196 35958 8274
rect 36236 8196 36546 8274
rect 36824 8196 37134 8274
rect 37412 8196 37722 8274
rect 38000 8196 38310 8274
rect 38588 8196 38642 8274
rect 22434 8186 22712 8196
rect 23022 8186 23300 8196
rect 23610 8186 23888 8196
rect 24198 8186 24476 8196
rect 24786 8186 25064 8196
rect 25374 8186 25652 8196
rect 25962 8186 26240 8196
rect 26550 8186 26828 8196
rect 27138 8186 27416 8196
rect 27726 8186 28004 8196
rect 28314 8186 28592 8196
rect 28902 8186 29180 8196
rect 29490 8186 29768 8196
rect 30078 8186 30356 8196
rect 30666 8186 30944 8196
rect 31254 8186 31532 8196
rect 31842 8186 32120 8196
rect 32430 8186 32708 8196
rect 33018 8186 33296 8196
rect 33606 8186 33884 8196
rect 34194 8186 34472 8196
rect 34782 8186 35060 8196
rect 35370 8186 35648 8196
rect 35958 8186 36236 8196
rect 36546 8186 36824 8196
rect 37134 8186 37412 8196
rect 37722 8186 38000 8196
rect 38310 8186 38588 8196
rect 44380 6952 45446 6962
rect 26232 6240 44380 6750
rect 44380 6134 45446 6144
rect 5800 5160 7070 5170
rect 5288 3996 5800 4988
rect 22920 4392 22938 4436
rect 7070 3996 22938 4392
rect 5800 3788 7070 3798
<< via2 >>
rect 37832 20906 38980 22370
rect 3546 11952 5048 13186
rect 5800 4988 7070 5160
rect 5800 3996 6278 4988
rect 6278 3996 7030 4988
rect 7030 3996 7070 4988
rect 5800 3798 7070 3996
<< metal3 >>
rect 37822 22370 38990 22375
rect 37822 20906 37832 22370
rect 38980 20906 38990 22370
rect 37822 20901 38990 20906
rect 37896 17768 38708 20901
rect 37330 16240 37340 17768
rect 39154 16240 39164 17768
rect -10524 4988 2588 15568
rect 3536 13186 5058 13191
rect 3536 11952 3546 13186
rect 5048 11952 5058 13186
rect 3536 11947 5058 11952
rect 5790 5160 7080 5165
rect 5790 4988 5800 5160
rect -10524 3996 5800 4988
rect -10524 2468 2588 3996
rect 5790 3798 5800 3996
rect 7070 3798 7080 5160
rect 5790 3793 7080 3798
<< via3 >>
rect 37340 16240 39154 17768
rect 3546 11952 5048 13186
<< mimcap >>
rect -10423 15428 -7423 15468
rect -10423 12508 -10383 15428
rect -7463 12508 -7423 15428
rect -10423 12468 -7423 12508
rect -7104 15428 -4104 15468
rect -7104 12508 -7064 15428
rect -4144 12508 -4104 15428
rect -7104 12468 -4104 12508
rect -3785 15428 -785 15468
rect -3785 12508 -3745 15428
rect -825 12508 -785 15428
rect -3785 12468 -785 12508
rect -466 15428 2534 15468
rect -466 12508 -426 15428
rect 2494 12508 2534 15428
rect -466 12468 2534 12508
rect -10423 12128 -7423 12168
rect -10423 9208 -10383 12128
rect -7463 9208 -7423 12128
rect -10423 9168 -7423 9208
rect -7104 12128 -4104 12168
rect -7104 9208 -7064 12128
rect -4144 9208 -4104 12128
rect -7104 9168 -4104 9208
rect -3785 12128 -785 12168
rect -3785 9208 -3745 12128
rect -825 9208 -785 12128
rect -3785 9168 -785 9208
rect -466 12128 2534 12168
rect -466 9208 -426 12128
rect 2494 9208 2534 12128
rect -466 9168 2534 9208
rect -10423 8828 -7423 8868
rect -10423 5908 -10383 8828
rect -7463 5908 -7423 8828
rect -10423 5868 -7423 5908
rect -7104 8828 -4104 8868
rect -7104 5908 -7064 8828
rect -4144 5908 -4104 8828
rect -7104 5868 -4104 5908
rect -3785 8828 -785 8868
rect -3785 5908 -3745 8828
rect -825 5908 -785 8828
rect -3785 5868 -785 5908
rect -466 8828 2534 8868
rect -466 5908 -426 8828
rect 2494 5908 2534 8828
rect -466 5868 2534 5908
rect -10423 5528 -7423 5568
rect -10423 2608 -10383 5528
rect -7463 2608 -7423 5528
rect -10423 2568 -7423 2608
rect -7104 5528 -4104 5568
rect -7104 2608 -7064 5528
rect -4144 2608 -4104 5528
rect -7104 2568 -4104 2608
rect -3785 5528 -785 5568
rect -3785 2608 -3745 5528
rect -825 2608 -785 5528
rect -3785 2568 -785 2608
rect -466 5528 2534 5568
rect -466 2608 -426 5528
rect 2494 2608 2534 5528
rect -466 2568 2534 2608
<< mimcapcontact >>
rect -10383 12508 -7463 15428
rect -7064 12508 -4144 15428
rect -3745 12508 -825 15428
rect -426 12508 2494 15428
rect -10383 9208 -7463 12128
rect -7064 9208 -4144 12128
rect -3745 9208 -825 12128
rect -426 9208 2494 12128
rect -10383 5908 -7463 8828
rect -7064 5908 -4144 8828
rect -3745 5908 -825 8828
rect -426 5908 2494 8828
rect -10383 2608 -7463 5528
rect -7064 2608 -4144 5528
rect -3745 2608 -825 5528
rect -426 2608 2494 5528
<< metal4 >>
rect 11210 24550 11594 24622
rect 11798 24550 12182 24622
rect 12386 24550 12770 24622
rect 12974 24550 13358 24622
rect 13562 24550 13946 24622
rect 14150 24550 14534 24622
rect 14738 24550 15122 24622
rect 15326 24550 15710 24622
rect 15914 24550 16298 24622
rect 16502 24550 16886 24622
rect 17090 24550 17474 24622
rect 17678 24550 18062 24622
rect 18266 24550 18650 24622
rect 18854 24550 19238 24622
rect 19442 24550 19826 24622
rect 20030 24550 20414 24622
rect 20618 24550 21002 24622
rect 21206 24550 21590 24622
rect 21794 24550 22178 24622
rect 22986 24544 23354 24632
rect 23574 24544 23942 24632
rect 24162 24544 24530 24632
rect 24750 24544 25118 24632
rect 25338 24544 25706 24632
rect 25926 24544 26294 24632
rect 26514 24544 26882 24632
rect 27102 24544 27470 24632
rect 27690 24544 28058 24632
rect 28278 24544 28646 24632
rect 28866 24544 29234 24632
rect 29454 24544 29822 24632
rect 30042 24544 30410 24632
rect 30630 24544 30998 24632
rect 31218 24544 31586 24632
rect 31806 24544 32174 24632
rect 32394 24544 32762 24632
rect 32982 24544 33350 24632
rect 33570 24544 33938 24632
rect 34158 24544 34526 24632
rect 34746 24544 35114 24632
rect 35334 24544 35702 24632
rect 35922 24544 36290 24632
rect 36510 24544 36878 24632
rect 37098 24544 37466 24632
rect 37686 24544 38054 24632
rect 38274 24544 38642 24632
rect 39290 23634 43290 25164
rect 37339 17768 39155 17769
rect -8975 15568 -8871 15618
rect -5656 15568 -5552 15618
rect -2337 15568 -2233 15618
rect 982 15568 1086 15618
rect -10524 15428 2588 15568
rect -10524 12508 -10383 15428
rect -7463 12508 -7064 15428
rect -4144 12508 -3745 15428
rect -825 12508 -426 15428
rect 2494 13040 2588 15428
rect 8002 15326 9108 16946
rect 37339 16240 37340 17768
rect 39154 16240 39155 17768
rect 37339 16239 39155 16240
rect 3545 13186 5049 13187
rect 3545 13040 3546 13186
rect 2494 12508 3546 13040
rect -10524 12128 3546 12508
rect -10524 9208 -10383 12128
rect -7463 9208 -7064 12128
rect -4144 9208 -3745 12128
rect -825 9208 -426 12128
rect 2494 11990 3546 12128
rect 2494 9208 2588 11990
rect 3545 11952 3546 11990
rect 5048 11952 5049 13186
rect 3545 11951 5049 11952
rect -10524 8828 2588 9208
rect -10524 5908 -10383 8828
rect -7463 5908 -7064 8828
rect -4144 5908 -3745 8828
rect -825 5908 -426 8828
rect 2494 5908 2588 8828
rect 41964 8818 43290 23634
rect 11226 8198 11594 8286
rect 11814 8198 12182 8286
rect 12402 8198 12770 8286
rect 12990 8198 13358 8286
rect 13578 8198 13946 8286
rect 14166 8198 14534 8286
rect 14754 8198 15122 8286
rect 15342 8198 15710 8286
rect 15930 8198 16298 8286
rect 16518 8198 16886 8286
rect 17106 8198 17474 8286
rect 17694 8198 18062 8286
rect 18282 8198 18650 8286
rect 18870 8198 19238 8286
rect 19458 8198 19826 8286
rect 20046 8198 20414 8286
rect 20634 8198 21002 8286
rect 21222 8198 21590 8286
rect 21810 8198 22178 8286
rect 22986 8186 23354 8284
rect 23574 8186 23942 8284
rect 24162 8186 24530 8284
rect 24750 8186 25118 8284
rect 25338 8186 25706 8284
rect 25926 8186 26294 8284
rect 26514 8186 26882 8284
rect 27102 8186 27470 8284
rect 27690 8186 28058 8284
rect 28278 8186 28646 8284
rect 28866 8186 29234 8284
rect 29454 8186 29822 8284
rect 30042 8186 30410 8284
rect 30630 8186 30998 8284
rect 31218 8186 31586 8284
rect 31806 8186 32174 8284
rect 32394 8186 32762 8284
rect 32982 8186 33350 8284
rect 33570 8186 33938 8284
rect 34158 8186 34526 8284
rect 34746 8186 35114 8284
rect 35334 8186 35702 8284
rect 35922 8186 36290 8284
rect 36510 8186 36878 8284
rect 37098 8186 37466 8284
rect 37686 8186 38054 8284
rect 38274 8186 38642 8284
rect 39448 7288 43290 8818
rect -10524 5528 2588 5908
rect -10524 2608 -10383 5528
rect -7463 2608 -7064 5528
rect -4144 2608 -3745 5528
rect -825 2608 -426 5528
rect 2494 2608 2588 5528
rect -10524 2468 2588 2608
rect -8975 2418 -8871 2468
rect -5656 2418 -5552 2468
rect -2337 2418 -2233 2468
rect 982 2418 1086 2468
<< comment >>
rect 30580 19352 31202 19420
rect 30580 18898 30674 19352
rect 31138 18898 31202 19352
rect 30580 18796 31202 18898
use OTA_tri  OTA_tri_0 ~/magic/class_d_audio_amplifier/OTA
timestamp 1627023135
transform 1 0 12 0 1 -6
box 7082 6 39470 16350
use OTA  OTA_0 ~/magic/class_d_audio_amplifier/OTA
timestamp 1627028181
transform 1 0 26464 0 1 35750
box -19208 -19408 12858 -3006
<< labels >>
flabel metal4 8616 16242 8616 16242 0 FreeSans 3200 0 0 0 vss
flabel metal4 41924 8146 41924 8146 0 FreeSans 3200 0 0 0 vdd
flabel metal1 38930 12424 38930 12424 0 FreeSans 3200 0 0 0 vt
flabel metal1 44814 13146 44814 13146 0 FreeSans 3200 0 0 0 vref
flabel metal2 10462 26556 10462 26556 0 FreeSans 3200 0 0 0 vbias2
flabel metal2 10386 10184 10386 10184 0 FreeSans 3200 0 0 0 vbias1
flabel metal1 37232 28710 37232 28710 0 FreeSans 3200 0 0 0 vsquare
<< end >>
