magic
tech sky130A
magscale 1 2
timestamp 1627028181
<< nwell >>
rect -16334 -11632 12686 -7768
rect -3322 -16172 -326 -12142
<< pwell >>
rect -7030 -6248 3384 -3612
rect 4201 -16109 4603 -14813
rect -2710 -18950 -936 -16334
<< pmoslvt >>
rect -15842 -9100 -15442 -8300
rect -15254 -9100 -14854 -8300
rect -14666 -9100 -14266 -8300
rect -14078 -9100 -13678 -8300
rect -13490 -9100 -13090 -8300
rect -12902 -9100 -12502 -8300
rect -12314 -9100 -11914 -8300
rect -11726 -9100 -11326 -8300
rect -11138 -9100 -10738 -8300
rect -10550 -9100 -10150 -8300
rect -9962 -9100 -9562 -8300
rect -9374 -9100 -8974 -8300
rect -8786 -9100 -8386 -8300
rect -8198 -9100 -7798 -8300
rect -7610 -9100 -7210 -8300
rect -7022 -9100 -6622 -8300
rect -6434 -9100 -6034 -8300
rect -5846 -9100 -5446 -8300
rect -5258 -9100 -4858 -8300
rect -4670 -9100 -4270 -8300
rect -4082 -9100 -3682 -8300
rect -3494 -9100 -3094 -8300
rect -2906 -9100 -2506 -8300
rect -2318 -9100 -1918 -8300
rect -1730 -9100 -1330 -8300
rect -1142 -9100 -742 -8300
rect -554 -9100 -154 -8300
rect 34 -9100 434 -8300
rect 622 -9100 1022 -8300
rect 1210 -9100 1610 -8300
rect 1798 -9100 2198 -8300
rect 2386 -9100 2786 -8300
rect 2974 -9100 3374 -8300
rect 3562 -9100 3962 -8300
rect 4150 -9100 4550 -8300
rect 4738 -9100 5138 -8300
rect 5326 -9100 5726 -8300
rect 5914 -9100 6314 -8300
rect 6502 -9100 6902 -8300
rect 7090 -9100 7490 -8300
rect 7678 -9100 8078 -8300
rect 8266 -9100 8666 -8300
rect 8854 -9100 9254 -8300
rect 9442 -9100 9842 -8300
rect 10030 -9100 10430 -8300
rect 10618 -9100 11018 -8300
rect 11206 -9100 11606 -8300
rect 11794 -9100 12194 -8300
rect -15842 -10100 -15442 -9300
rect -15254 -10100 -14854 -9300
rect -14666 -10100 -14266 -9300
rect -14078 -10100 -13678 -9300
rect -13490 -10100 -13090 -9300
rect -12902 -10100 -12502 -9300
rect -12314 -10100 -11914 -9300
rect -11726 -10100 -11326 -9300
rect -11138 -10100 -10738 -9300
rect -10550 -10100 -10150 -9300
rect -9962 -10100 -9562 -9300
rect -9374 -10100 -8974 -9300
rect -8786 -10100 -8386 -9300
rect -8198 -10100 -7798 -9300
rect -7610 -10100 -7210 -9300
rect -7022 -10100 -6622 -9300
rect -6434 -10100 -6034 -9300
rect -5846 -10100 -5446 -9300
rect -5258 -10100 -4858 -9300
rect -4670 -10100 -4270 -9300
rect -4082 -10100 -3682 -9300
rect -3494 -10100 -3094 -9300
rect -2906 -10100 -2506 -9300
rect -2318 -10100 -1918 -9300
rect -1730 -10100 -1330 -9300
rect -1142 -10100 -742 -9300
rect -554 -10100 -154 -9300
rect 34 -10100 434 -9300
rect 622 -10100 1022 -9300
rect 1210 -10100 1610 -9300
rect 1798 -10100 2198 -9300
rect 2386 -10100 2786 -9300
rect 2974 -10100 3374 -9300
rect 3562 -10100 3962 -9300
rect 4150 -10100 4550 -9300
rect 4738 -10100 5138 -9300
rect 5326 -10100 5726 -9300
rect 5914 -10100 6314 -9300
rect 6502 -10100 6902 -9300
rect 7090 -10100 7490 -9300
rect 7678 -10100 8078 -9300
rect 8266 -10100 8666 -9300
rect 8854 -10100 9254 -9300
rect 9442 -10100 9842 -9300
rect 10030 -10100 10430 -9300
rect 10618 -10100 11018 -9300
rect 11206 -10100 11606 -9300
rect 11794 -10100 12194 -9300
rect -15842 -11100 -15442 -10300
rect -15254 -11100 -14854 -10300
rect -14666 -11100 -14266 -10300
rect -14078 -11100 -13678 -10300
rect -13490 -11100 -13090 -10300
rect -12902 -11100 -12502 -10300
rect -12314 -11100 -11914 -10300
rect -11726 -11100 -11326 -10300
rect -11138 -11100 -10738 -10300
rect -10550 -11100 -10150 -10300
rect -9962 -11100 -9562 -10300
rect -9374 -11100 -8974 -10300
rect -8786 -11100 -8386 -10300
rect -8198 -11100 -7798 -10300
rect -7610 -11100 -7210 -10300
rect -7022 -11100 -6622 -10300
rect -6434 -11100 -6034 -10300
rect -5846 -11100 -5446 -10300
rect -5258 -11100 -4858 -10300
rect -4670 -11100 -4270 -10300
rect -4082 -11100 -3682 -10300
rect -3494 -11100 -3094 -10300
rect -2906 -11100 -2506 -10300
rect -2318 -11100 -1918 -10300
rect -1730 -11100 -1330 -10300
rect -1142 -11100 -742 -10300
rect -554 -11100 -154 -10300
rect 34 -11100 434 -10300
rect 622 -11100 1022 -10300
rect 1210 -11100 1610 -10300
rect 1798 -11100 2198 -10300
rect 2386 -11100 2786 -10300
rect 2974 -11100 3374 -10300
rect 3562 -11100 3962 -10300
rect 4150 -11100 4550 -10300
rect 4738 -11100 5138 -10300
rect 5326 -11100 5726 -10300
rect 5914 -11100 6314 -10300
rect 6502 -11100 6902 -10300
rect 7090 -11100 7490 -10300
rect 7678 -11100 8078 -10300
rect 8266 -11100 8666 -10300
rect 8854 -11100 9254 -10300
rect 9442 -11100 9842 -10300
rect 10030 -11100 10430 -10300
rect 10618 -11100 11018 -10300
rect 11206 -11100 11606 -10300
rect 11794 -11100 12194 -10300
rect -2790 -13546 -2720 -12746
rect -2524 -13546 -2454 -12746
rect -2258 -13546 -2188 -12746
rect -1992 -13546 -1922 -12746
rect -1726 -13546 -1656 -12746
rect -1460 -13546 -1390 -12746
rect -1194 -13546 -1124 -12746
rect -928 -13546 -858 -12746
rect -2790 -14556 -2720 -13756
rect -2524 -14556 -2454 -13756
rect -2258 -14556 -2188 -13756
rect -1992 -14556 -1922 -13756
rect -1726 -14556 -1656 -13756
rect -1460 -14556 -1390 -13756
rect -1194 -14556 -1124 -13756
rect -928 -14556 -858 -13756
rect -2790 -15566 -2720 -14766
rect -2524 -15566 -2454 -14766
rect -2258 -15566 -2188 -14766
rect -1992 -15566 -1922 -14766
rect -1726 -15566 -1656 -14766
rect -1460 -15566 -1390 -14766
rect -1194 -15566 -1124 -14766
rect -928 -15566 -858 -14766
<< nmoslvt >>
rect -6538 -4826 -6468 -4226
rect -6298 -4826 -6228 -4226
rect -6058 -4826 -5988 -4226
rect -5818 -4826 -5748 -4226
rect -5578 -4826 -5508 -4226
rect -5338 -4826 -5268 -4226
rect -5098 -4826 -5028 -4226
rect -4858 -4826 -4788 -4226
rect -4618 -4826 -4548 -4226
rect -4378 -4826 -4308 -4226
rect -4138 -4826 -4068 -4226
rect -3898 -4826 -3828 -4226
rect -3658 -4826 -3588 -4226
rect -3418 -4826 -3348 -4226
rect -3178 -4826 -3108 -4226
rect -2938 -4826 -2868 -4226
rect -2698 -4826 -2628 -4226
rect -2458 -4826 -2388 -4226
rect -2218 -4826 -2148 -4226
rect -1978 -4826 -1908 -4226
rect -1738 -4826 -1668 -4226
rect -1498 -4826 -1428 -4226
rect -1258 -4826 -1188 -4226
rect -1018 -4826 -948 -4226
rect -778 -4826 -708 -4226
rect -538 -4826 -468 -4226
rect -298 -4826 -228 -4226
rect -58 -4826 12 -4226
rect 182 -4826 252 -4226
rect 422 -4826 492 -4226
rect 662 -4826 732 -4226
rect 902 -4826 972 -4226
rect 1142 -4826 1212 -4226
rect 1382 -4826 1452 -4226
rect 1622 -4826 1692 -4226
rect 1862 -4826 1932 -4226
rect 2102 -4826 2172 -4226
rect 2342 -4826 2412 -4226
rect 2582 -4826 2652 -4226
rect 2822 -4826 2892 -4226
rect -6538 -5634 -6468 -5034
rect -6298 -5634 -6228 -5034
rect -6058 -5634 -5988 -5034
rect -5818 -5634 -5748 -5034
rect -5578 -5634 -5508 -5034
rect -5338 -5634 -5268 -5034
rect -5098 -5634 -5028 -5034
rect -4858 -5634 -4788 -5034
rect -4618 -5634 -4548 -5034
rect -4378 -5634 -4308 -5034
rect -4138 -5634 -4068 -5034
rect -3898 -5634 -3828 -5034
rect -3658 -5634 -3588 -5034
rect -3418 -5634 -3348 -5034
rect -3178 -5634 -3108 -5034
rect -2938 -5634 -2868 -5034
rect -2698 -5634 -2628 -5034
rect -2458 -5634 -2388 -5034
rect -2218 -5634 -2148 -5034
rect -1978 -5634 -1908 -5034
rect -1738 -5634 -1668 -5034
rect -1498 -5634 -1428 -5034
rect -1258 -5634 -1188 -5034
rect -1018 -5634 -948 -5034
rect -778 -5634 -708 -5034
rect -538 -5634 -468 -5034
rect -298 -5634 -228 -5034
rect -58 -5634 12 -5034
rect 182 -5634 252 -5034
rect 422 -5634 492 -5034
rect 662 -5634 732 -5034
rect 902 -5634 972 -5034
rect 1142 -5634 1212 -5034
rect 1382 -5634 1452 -5034
rect 1622 -5634 1692 -5034
rect 1862 -5634 1932 -5034
rect 2102 -5634 2172 -5034
rect 2342 -5634 2412 -5034
rect 2582 -5634 2652 -5034
rect 2822 -5634 2892 -5034
rect -2218 -17538 -2148 -16938
rect -1978 -17538 -1908 -16938
rect -1738 -17538 -1668 -16938
rect -1498 -17538 -1428 -16938
rect -2218 -18346 -2148 -17746
rect -1978 -18346 -1908 -17746
rect -1738 -18346 -1668 -17746
rect -1498 -18346 -1428 -17746
<< ndiff >>
rect -6596 -4238 -6538 -4226
rect -6596 -4814 -6584 -4238
rect -6550 -4814 -6538 -4238
rect -6596 -4826 -6538 -4814
rect -6468 -4238 -6410 -4226
rect -6468 -4814 -6456 -4238
rect -6422 -4814 -6410 -4238
rect -6468 -4826 -6410 -4814
rect -6356 -4238 -6298 -4226
rect -6356 -4814 -6344 -4238
rect -6310 -4814 -6298 -4238
rect -6356 -4826 -6298 -4814
rect -6228 -4238 -6170 -4226
rect -6228 -4814 -6216 -4238
rect -6182 -4814 -6170 -4238
rect -6228 -4826 -6170 -4814
rect -6116 -4238 -6058 -4226
rect -6116 -4814 -6104 -4238
rect -6070 -4814 -6058 -4238
rect -6116 -4826 -6058 -4814
rect -5988 -4238 -5930 -4226
rect -5988 -4814 -5976 -4238
rect -5942 -4814 -5930 -4238
rect -5988 -4826 -5930 -4814
rect -5876 -4238 -5818 -4226
rect -5876 -4814 -5864 -4238
rect -5830 -4814 -5818 -4238
rect -5876 -4826 -5818 -4814
rect -5748 -4238 -5690 -4226
rect -5748 -4814 -5736 -4238
rect -5702 -4814 -5690 -4238
rect -5748 -4826 -5690 -4814
rect -5636 -4238 -5578 -4226
rect -5636 -4814 -5624 -4238
rect -5590 -4814 -5578 -4238
rect -5636 -4826 -5578 -4814
rect -5508 -4238 -5450 -4226
rect -5508 -4814 -5496 -4238
rect -5462 -4814 -5450 -4238
rect -5508 -4826 -5450 -4814
rect -5396 -4238 -5338 -4226
rect -5396 -4814 -5384 -4238
rect -5350 -4814 -5338 -4238
rect -5396 -4826 -5338 -4814
rect -5268 -4238 -5210 -4226
rect -5268 -4814 -5256 -4238
rect -5222 -4814 -5210 -4238
rect -5268 -4826 -5210 -4814
rect -5156 -4238 -5098 -4226
rect -5156 -4814 -5144 -4238
rect -5110 -4814 -5098 -4238
rect -5156 -4826 -5098 -4814
rect -5028 -4238 -4970 -4226
rect -5028 -4814 -5016 -4238
rect -4982 -4814 -4970 -4238
rect -5028 -4826 -4970 -4814
rect -4916 -4238 -4858 -4226
rect -4916 -4814 -4904 -4238
rect -4870 -4814 -4858 -4238
rect -4916 -4826 -4858 -4814
rect -4788 -4238 -4730 -4226
rect -4788 -4814 -4776 -4238
rect -4742 -4814 -4730 -4238
rect -4788 -4826 -4730 -4814
rect -4676 -4238 -4618 -4226
rect -4676 -4814 -4664 -4238
rect -4630 -4814 -4618 -4238
rect -4676 -4826 -4618 -4814
rect -4548 -4238 -4490 -4226
rect -4548 -4814 -4536 -4238
rect -4502 -4814 -4490 -4238
rect -4548 -4826 -4490 -4814
rect -4436 -4238 -4378 -4226
rect -4436 -4814 -4424 -4238
rect -4390 -4814 -4378 -4238
rect -4436 -4826 -4378 -4814
rect -4308 -4238 -4250 -4226
rect -4308 -4814 -4296 -4238
rect -4262 -4814 -4250 -4238
rect -4308 -4826 -4250 -4814
rect -4196 -4238 -4138 -4226
rect -4196 -4814 -4184 -4238
rect -4150 -4814 -4138 -4238
rect -4196 -4826 -4138 -4814
rect -4068 -4238 -4010 -4226
rect -4068 -4814 -4056 -4238
rect -4022 -4814 -4010 -4238
rect -4068 -4826 -4010 -4814
rect -3956 -4238 -3898 -4226
rect -3956 -4814 -3944 -4238
rect -3910 -4814 -3898 -4238
rect -3956 -4826 -3898 -4814
rect -3828 -4238 -3770 -4226
rect -3828 -4814 -3816 -4238
rect -3782 -4814 -3770 -4238
rect -3828 -4826 -3770 -4814
rect -3716 -4238 -3658 -4226
rect -3716 -4814 -3704 -4238
rect -3670 -4814 -3658 -4238
rect -3716 -4826 -3658 -4814
rect -3588 -4238 -3530 -4226
rect -3588 -4814 -3576 -4238
rect -3542 -4814 -3530 -4238
rect -3588 -4826 -3530 -4814
rect -3476 -4238 -3418 -4226
rect -3476 -4814 -3464 -4238
rect -3430 -4814 -3418 -4238
rect -3476 -4826 -3418 -4814
rect -3348 -4238 -3290 -4226
rect -3348 -4814 -3336 -4238
rect -3302 -4814 -3290 -4238
rect -3348 -4826 -3290 -4814
rect -3236 -4238 -3178 -4226
rect -3236 -4814 -3224 -4238
rect -3190 -4814 -3178 -4238
rect -3236 -4826 -3178 -4814
rect -3108 -4238 -3050 -4226
rect -3108 -4814 -3096 -4238
rect -3062 -4814 -3050 -4238
rect -3108 -4826 -3050 -4814
rect -2996 -4238 -2938 -4226
rect -2996 -4814 -2984 -4238
rect -2950 -4814 -2938 -4238
rect -2996 -4826 -2938 -4814
rect -2868 -4238 -2810 -4226
rect -2868 -4814 -2856 -4238
rect -2822 -4814 -2810 -4238
rect -2868 -4826 -2810 -4814
rect -2756 -4238 -2698 -4226
rect -2756 -4814 -2744 -4238
rect -2710 -4814 -2698 -4238
rect -2756 -4826 -2698 -4814
rect -2628 -4238 -2570 -4226
rect -2628 -4814 -2616 -4238
rect -2582 -4814 -2570 -4238
rect -2628 -4826 -2570 -4814
rect -2516 -4238 -2458 -4226
rect -2516 -4814 -2504 -4238
rect -2470 -4814 -2458 -4238
rect -2516 -4826 -2458 -4814
rect -2388 -4238 -2330 -4226
rect -2388 -4814 -2376 -4238
rect -2342 -4814 -2330 -4238
rect -2388 -4826 -2330 -4814
rect -2276 -4238 -2218 -4226
rect -2276 -4814 -2264 -4238
rect -2230 -4814 -2218 -4238
rect -2276 -4826 -2218 -4814
rect -2148 -4238 -2090 -4226
rect -2148 -4814 -2136 -4238
rect -2102 -4814 -2090 -4238
rect -2148 -4826 -2090 -4814
rect -2036 -4238 -1978 -4226
rect -2036 -4814 -2024 -4238
rect -1990 -4814 -1978 -4238
rect -2036 -4826 -1978 -4814
rect -1908 -4238 -1850 -4226
rect -1908 -4814 -1896 -4238
rect -1862 -4814 -1850 -4238
rect -1908 -4826 -1850 -4814
rect -1796 -4238 -1738 -4226
rect -1796 -4814 -1784 -4238
rect -1750 -4814 -1738 -4238
rect -1796 -4826 -1738 -4814
rect -1668 -4238 -1610 -4226
rect -1668 -4814 -1656 -4238
rect -1622 -4814 -1610 -4238
rect -1668 -4826 -1610 -4814
rect -1556 -4238 -1498 -4226
rect -1556 -4814 -1544 -4238
rect -1510 -4814 -1498 -4238
rect -1556 -4826 -1498 -4814
rect -1428 -4238 -1370 -4226
rect -1428 -4814 -1416 -4238
rect -1382 -4814 -1370 -4238
rect -1428 -4826 -1370 -4814
rect -1316 -4238 -1258 -4226
rect -1316 -4814 -1304 -4238
rect -1270 -4814 -1258 -4238
rect -1316 -4826 -1258 -4814
rect -1188 -4238 -1130 -4226
rect -1188 -4814 -1176 -4238
rect -1142 -4814 -1130 -4238
rect -1188 -4826 -1130 -4814
rect -1076 -4238 -1018 -4226
rect -1076 -4814 -1064 -4238
rect -1030 -4814 -1018 -4238
rect -1076 -4826 -1018 -4814
rect -948 -4238 -890 -4226
rect -948 -4814 -936 -4238
rect -902 -4814 -890 -4238
rect -948 -4826 -890 -4814
rect -836 -4238 -778 -4226
rect -836 -4814 -824 -4238
rect -790 -4814 -778 -4238
rect -836 -4826 -778 -4814
rect -708 -4238 -650 -4226
rect -708 -4814 -696 -4238
rect -662 -4814 -650 -4238
rect -708 -4826 -650 -4814
rect -596 -4238 -538 -4226
rect -596 -4814 -584 -4238
rect -550 -4814 -538 -4238
rect -596 -4826 -538 -4814
rect -468 -4238 -410 -4226
rect -468 -4814 -456 -4238
rect -422 -4814 -410 -4238
rect -468 -4826 -410 -4814
rect -356 -4238 -298 -4226
rect -356 -4814 -344 -4238
rect -310 -4814 -298 -4238
rect -356 -4826 -298 -4814
rect -228 -4238 -170 -4226
rect -228 -4814 -216 -4238
rect -182 -4814 -170 -4238
rect -228 -4826 -170 -4814
rect -116 -4238 -58 -4226
rect -116 -4814 -104 -4238
rect -70 -4814 -58 -4238
rect -116 -4826 -58 -4814
rect 12 -4238 70 -4226
rect 12 -4814 24 -4238
rect 58 -4814 70 -4238
rect 12 -4826 70 -4814
rect 124 -4238 182 -4226
rect 124 -4814 136 -4238
rect 170 -4814 182 -4238
rect 124 -4826 182 -4814
rect 252 -4238 310 -4226
rect 252 -4814 264 -4238
rect 298 -4814 310 -4238
rect 252 -4826 310 -4814
rect 364 -4238 422 -4226
rect 364 -4814 376 -4238
rect 410 -4814 422 -4238
rect 364 -4826 422 -4814
rect 492 -4238 550 -4226
rect 492 -4814 504 -4238
rect 538 -4814 550 -4238
rect 492 -4826 550 -4814
rect 604 -4238 662 -4226
rect 604 -4814 616 -4238
rect 650 -4814 662 -4238
rect 604 -4826 662 -4814
rect 732 -4238 790 -4226
rect 732 -4814 744 -4238
rect 778 -4814 790 -4238
rect 732 -4826 790 -4814
rect 844 -4238 902 -4226
rect 844 -4814 856 -4238
rect 890 -4814 902 -4238
rect 844 -4826 902 -4814
rect 972 -4238 1030 -4226
rect 972 -4814 984 -4238
rect 1018 -4814 1030 -4238
rect 972 -4826 1030 -4814
rect 1084 -4238 1142 -4226
rect 1084 -4814 1096 -4238
rect 1130 -4814 1142 -4238
rect 1084 -4826 1142 -4814
rect 1212 -4238 1270 -4226
rect 1212 -4814 1224 -4238
rect 1258 -4814 1270 -4238
rect 1212 -4826 1270 -4814
rect 1324 -4238 1382 -4226
rect 1324 -4814 1336 -4238
rect 1370 -4814 1382 -4238
rect 1324 -4826 1382 -4814
rect 1452 -4238 1510 -4226
rect 1452 -4814 1464 -4238
rect 1498 -4814 1510 -4238
rect 1452 -4826 1510 -4814
rect 1564 -4238 1622 -4226
rect 1564 -4814 1576 -4238
rect 1610 -4814 1622 -4238
rect 1564 -4826 1622 -4814
rect 1692 -4238 1750 -4226
rect 1692 -4814 1704 -4238
rect 1738 -4814 1750 -4238
rect 1692 -4826 1750 -4814
rect 1804 -4238 1862 -4226
rect 1804 -4814 1816 -4238
rect 1850 -4814 1862 -4238
rect 1804 -4826 1862 -4814
rect 1932 -4238 1990 -4226
rect 1932 -4814 1944 -4238
rect 1978 -4814 1990 -4238
rect 1932 -4826 1990 -4814
rect 2044 -4238 2102 -4226
rect 2044 -4814 2056 -4238
rect 2090 -4814 2102 -4238
rect 2044 -4826 2102 -4814
rect 2172 -4238 2230 -4226
rect 2172 -4814 2184 -4238
rect 2218 -4814 2230 -4238
rect 2172 -4826 2230 -4814
rect 2284 -4238 2342 -4226
rect 2284 -4814 2296 -4238
rect 2330 -4814 2342 -4238
rect 2284 -4826 2342 -4814
rect 2412 -4238 2470 -4226
rect 2412 -4814 2424 -4238
rect 2458 -4814 2470 -4238
rect 2412 -4826 2470 -4814
rect 2524 -4238 2582 -4226
rect 2524 -4814 2536 -4238
rect 2570 -4814 2582 -4238
rect 2524 -4826 2582 -4814
rect 2652 -4238 2710 -4226
rect 2652 -4814 2664 -4238
rect 2698 -4814 2710 -4238
rect 2652 -4826 2710 -4814
rect 2764 -4238 2822 -4226
rect 2764 -4814 2776 -4238
rect 2810 -4814 2822 -4238
rect 2764 -4826 2822 -4814
rect 2892 -4238 2950 -4226
rect 2892 -4814 2904 -4238
rect 2938 -4814 2950 -4238
rect 2892 -4826 2950 -4814
rect -6596 -5046 -6538 -5034
rect -6596 -5622 -6584 -5046
rect -6550 -5622 -6538 -5046
rect -6596 -5634 -6538 -5622
rect -6468 -5046 -6410 -5034
rect -6468 -5622 -6456 -5046
rect -6422 -5622 -6410 -5046
rect -6468 -5634 -6410 -5622
rect -6356 -5046 -6298 -5034
rect -6356 -5622 -6344 -5046
rect -6310 -5622 -6298 -5046
rect -6356 -5634 -6298 -5622
rect -6228 -5046 -6170 -5034
rect -6228 -5622 -6216 -5046
rect -6182 -5622 -6170 -5046
rect -6228 -5634 -6170 -5622
rect -6116 -5046 -6058 -5034
rect -6116 -5622 -6104 -5046
rect -6070 -5622 -6058 -5046
rect -6116 -5634 -6058 -5622
rect -5988 -5046 -5930 -5034
rect -5988 -5622 -5976 -5046
rect -5942 -5622 -5930 -5046
rect -5988 -5634 -5930 -5622
rect -5876 -5046 -5818 -5034
rect -5876 -5622 -5864 -5046
rect -5830 -5622 -5818 -5046
rect -5876 -5634 -5818 -5622
rect -5748 -5046 -5690 -5034
rect -5748 -5622 -5736 -5046
rect -5702 -5622 -5690 -5046
rect -5748 -5634 -5690 -5622
rect -5636 -5046 -5578 -5034
rect -5636 -5622 -5624 -5046
rect -5590 -5622 -5578 -5046
rect -5636 -5634 -5578 -5622
rect -5508 -5046 -5450 -5034
rect -5508 -5622 -5496 -5046
rect -5462 -5622 -5450 -5046
rect -5508 -5634 -5450 -5622
rect -5396 -5046 -5338 -5034
rect -5396 -5622 -5384 -5046
rect -5350 -5622 -5338 -5046
rect -5396 -5634 -5338 -5622
rect -5268 -5046 -5210 -5034
rect -5268 -5622 -5256 -5046
rect -5222 -5622 -5210 -5046
rect -5268 -5634 -5210 -5622
rect -5156 -5046 -5098 -5034
rect -5156 -5622 -5144 -5046
rect -5110 -5622 -5098 -5046
rect -5156 -5634 -5098 -5622
rect -5028 -5046 -4970 -5034
rect -5028 -5622 -5016 -5046
rect -4982 -5622 -4970 -5046
rect -5028 -5634 -4970 -5622
rect -4916 -5046 -4858 -5034
rect -4916 -5622 -4904 -5046
rect -4870 -5622 -4858 -5046
rect -4916 -5634 -4858 -5622
rect -4788 -5046 -4730 -5034
rect -4788 -5622 -4776 -5046
rect -4742 -5622 -4730 -5046
rect -4788 -5634 -4730 -5622
rect -4676 -5046 -4618 -5034
rect -4676 -5622 -4664 -5046
rect -4630 -5622 -4618 -5046
rect -4676 -5634 -4618 -5622
rect -4548 -5046 -4490 -5034
rect -4548 -5622 -4536 -5046
rect -4502 -5622 -4490 -5046
rect -4548 -5634 -4490 -5622
rect -4436 -5046 -4378 -5034
rect -4436 -5622 -4424 -5046
rect -4390 -5622 -4378 -5046
rect -4436 -5634 -4378 -5622
rect -4308 -5046 -4250 -5034
rect -4308 -5622 -4296 -5046
rect -4262 -5622 -4250 -5046
rect -4308 -5634 -4250 -5622
rect -4196 -5046 -4138 -5034
rect -4196 -5622 -4184 -5046
rect -4150 -5622 -4138 -5046
rect -4196 -5634 -4138 -5622
rect -4068 -5046 -4010 -5034
rect -4068 -5622 -4056 -5046
rect -4022 -5622 -4010 -5046
rect -4068 -5634 -4010 -5622
rect -3956 -5046 -3898 -5034
rect -3956 -5622 -3944 -5046
rect -3910 -5622 -3898 -5046
rect -3956 -5634 -3898 -5622
rect -3828 -5046 -3770 -5034
rect -3828 -5622 -3816 -5046
rect -3782 -5622 -3770 -5046
rect -3828 -5634 -3770 -5622
rect -3716 -5046 -3658 -5034
rect -3716 -5622 -3704 -5046
rect -3670 -5622 -3658 -5046
rect -3716 -5634 -3658 -5622
rect -3588 -5046 -3530 -5034
rect -3588 -5622 -3576 -5046
rect -3542 -5622 -3530 -5046
rect -3588 -5634 -3530 -5622
rect -3476 -5046 -3418 -5034
rect -3476 -5622 -3464 -5046
rect -3430 -5622 -3418 -5046
rect -3476 -5634 -3418 -5622
rect -3348 -5046 -3290 -5034
rect -3348 -5622 -3336 -5046
rect -3302 -5622 -3290 -5046
rect -3348 -5634 -3290 -5622
rect -3236 -5046 -3178 -5034
rect -3236 -5622 -3224 -5046
rect -3190 -5622 -3178 -5046
rect -3236 -5634 -3178 -5622
rect -3108 -5046 -3050 -5034
rect -3108 -5622 -3096 -5046
rect -3062 -5622 -3050 -5046
rect -3108 -5634 -3050 -5622
rect -2996 -5046 -2938 -5034
rect -2996 -5622 -2984 -5046
rect -2950 -5622 -2938 -5046
rect -2996 -5634 -2938 -5622
rect -2868 -5046 -2810 -5034
rect -2868 -5622 -2856 -5046
rect -2822 -5622 -2810 -5046
rect -2868 -5634 -2810 -5622
rect -2756 -5046 -2698 -5034
rect -2756 -5622 -2744 -5046
rect -2710 -5622 -2698 -5046
rect -2756 -5634 -2698 -5622
rect -2628 -5046 -2570 -5034
rect -2628 -5622 -2616 -5046
rect -2582 -5622 -2570 -5046
rect -2628 -5634 -2570 -5622
rect -2516 -5046 -2458 -5034
rect -2516 -5622 -2504 -5046
rect -2470 -5622 -2458 -5046
rect -2516 -5634 -2458 -5622
rect -2388 -5046 -2330 -5034
rect -2388 -5622 -2376 -5046
rect -2342 -5622 -2330 -5046
rect -2388 -5634 -2330 -5622
rect -2276 -5046 -2218 -5034
rect -2276 -5622 -2264 -5046
rect -2230 -5622 -2218 -5046
rect -2276 -5634 -2218 -5622
rect -2148 -5046 -2090 -5034
rect -2148 -5622 -2136 -5046
rect -2102 -5622 -2090 -5046
rect -2148 -5634 -2090 -5622
rect -2036 -5046 -1978 -5034
rect -2036 -5622 -2024 -5046
rect -1990 -5622 -1978 -5046
rect -2036 -5634 -1978 -5622
rect -1908 -5046 -1850 -5034
rect -1908 -5622 -1896 -5046
rect -1862 -5622 -1850 -5046
rect -1908 -5634 -1850 -5622
rect -1796 -5046 -1738 -5034
rect -1796 -5622 -1784 -5046
rect -1750 -5622 -1738 -5046
rect -1796 -5634 -1738 -5622
rect -1668 -5046 -1610 -5034
rect -1668 -5622 -1656 -5046
rect -1622 -5622 -1610 -5046
rect -1668 -5634 -1610 -5622
rect -1556 -5046 -1498 -5034
rect -1556 -5622 -1544 -5046
rect -1510 -5622 -1498 -5046
rect -1556 -5634 -1498 -5622
rect -1428 -5046 -1370 -5034
rect -1428 -5622 -1416 -5046
rect -1382 -5622 -1370 -5046
rect -1428 -5634 -1370 -5622
rect -1316 -5046 -1258 -5034
rect -1316 -5622 -1304 -5046
rect -1270 -5622 -1258 -5046
rect -1316 -5634 -1258 -5622
rect -1188 -5046 -1130 -5034
rect -1188 -5622 -1176 -5046
rect -1142 -5622 -1130 -5046
rect -1188 -5634 -1130 -5622
rect -1076 -5046 -1018 -5034
rect -1076 -5622 -1064 -5046
rect -1030 -5622 -1018 -5046
rect -1076 -5634 -1018 -5622
rect -948 -5046 -890 -5034
rect -948 -5622 -936 -5046
rect -902 -5622 -890 -5046
rect -948 -5634 -890 -5622
rect -836 -5046 -778 -5034
rect -836 -5622 -824 -5046
rect -790 -5622 -778 -5046
rect -836 -5634 -778 -5622
rect -708 -5046 -650 -5034
rect -708 -5622 -696 -5046
rect -662 -5622 -650 -5046
rect -708 -5634 -650 -5622
rect -596 -5046 -538 -5034
rect -596 -5622 -584 -5046
rect -550 -5622 -538 -5046
rect -596 -5634 -538 -5622
rect -468 -5046 -410 -5034
rect -468 -5622 -456 -5046
rect -422 -5622 -410 -5046
rect -468 -5634 -410 -5622
rect -356 -5046 -298 -5034
rect -356 -5622 -344 -5046
rect -310 -5622 -298 -5046
rect -356 -5634 -298 -5622
rect -228 -5046 -170 -5034
rect -228 -5622 -216 -5046
rect -182 -5622 -170 -5046
rect -228 -5634 -170 -5622
rect -116 -5046 -58 -5034
rect -116 -5622 -104 -5046
rect -70 -5622 -58 -5046
rect -116 -5634 -58 -5622
rect 12 -5046 70 -5034
rect 12 -5622 24 -5046
rect 58 -5622 70 -5046
rect 12 -5634 70 -5622
rect 124 -5046 182 -5034
rect 124 -5622 136 -5046
rect 170 -5622 182 -5046
rect 124 -5634 182 -5622
rect 252 -5046 310 -5034
rect 252 -5622 264 -5046
rect 298 -5622 310 -5046
rect 252 -5634 310 -5622
rect 364 -5046 422 -5034
rect 364 -5622 376 -5046
rect 410 -5622 422 -5046
rect 364 -5634 422 -5622
rect 492 -5046 550 -5034
rect 492 -5622 504 -5046
rect 538 -5622 550 -5046
rect 492 -5634 550 -5622
rect 604 -5046 662 -5034
rect 604 -5622 616 -5046
rect 650 -5622 662 -5046
rect 604 -5634 662 -5622
rect 732 -5046 790 -5034
rect 732 -5622 744 -5046
rect 778 -5622 790 -5046
rect 732 -5634 790 -5622
rect 844 -5046 902 -5034
rect 844 -5622 856 -5046
rect 890 -5622 902 -5046
rect 844 -5634 902 -5622
rect 972 -5046 1030 -5034
rect 972 -5622 984 -5046
rect 1018 -5622 1030 -5046
rect 972 -5634 1030 -5622
rect 1084 -5046 1142 -5034
rect 1084 -5622 1096 -5046
rect 1130 -5622 1142 -5046
rect 1084 -5634 1142 -5622
rect 1212 -5046 1270 -5034
rect 1212 -5622 1224 -5046
rect 1258 -5622 1270 -5046
rect 1212 -5634 1270 -5622
rect 1324 -5046 1382 -5034
rect 1324 -5622 1336 -5046
rect 1370 -5622 1382 -5046
rect 1324 -5634 1382 -5622
rect 1452 -5046 1510 -5034
rect 1452 -5622 1464 -5046
rect 1498 -5622 1510 -5046
rect 1452 -5634 1510 -5622
rect 1564 -5046 1622 -5034
rect 1564 -5622 1576 -5046
rect 1610 -5622 1622 -5046
rect 1564 -5634 1622 -5622
rect 1692 -5046 1750 -5034
rect 1692 -5622 1704 -5046
rect 1738 -5622 1750 -5046
rect 1692 -5634 1750 -5622
rect 1804 -5046 1862 -5034
rect 1804 -5622 1816 -5046
rect 1850 -5622 1862 -5046
rect 1804 -5634 1862 -5622
rect 1932 -5046 1990 -5034
rect 1932 -5622 1944 -5046
rect 1978 -5622 1990 -5046
rect 1932 -5634 1990 -5622
rect 2044 -5046 2102 -5034
rect 2044 -5622 2056 -5046
rect 2090 -5622 2102 -5046
rect 2044 -5634 2102 -5622
rect 2172 -5046 2230 -5034
rect 2172 -5622 2184 -5046
rect 2218 -5622 2230 -5046
rect 2172 -5634 2230 -5622
rect 2284 -5046 2342 -5034
rect 2284 -5622 2296 -5046
rect 2330 -5622 2342 -5046
rect 2284 -5634 2342 -5622
rect 2412 -5046 2470 -5034
rect 2412 -5622 2424 -5046
rect 2458 -5622 2470 -5046
rect 2412 -5634 2470 -5622
rect 2524 -5046 2582 -5034
rect 2524 -5622 2536 -5046
rect 2570 -5622 2582 -5046
rect 2524 -5634 2582 -5622
rect 2652 -5046 2710 -5034
rect 2652 -5622 2664 -5046
rect 2698 -5622 2710 -5046
rect 2652 -5634 2710 -5622
rect 2764 -5046 2822 -5034
rect 2764 -5622 2776 -5046
rect 2810 -5622 2822 -5046
rect 2764 -5634 2822 -5622
rect 2892 -5046 2950 -5034
rect 2892 -5622 2904 -5046
rect 2938 -5622 2950 -5046
rect 2892 -5634 2950 -5622
rect -2276 -16950 -2218 -16938
rect -2276 -17526 -2264 -16950
rect -2230 -17526 -2218 -16950
rect -2276 -17538 -2218 -17526
rect -2148 -16950 -2090 -16938
rect -2148 -17526 -2136 -16950
rect -2102 -17526 -2090 -16950
rect -2148 -17538 -2090 -17526
rect -2036 -16950 -1978 -16938
rect -2036 -17526 -2024 -16950
rect -1990 -17526 -1978 -16950
rect -2036 -17538 -1978 -17526
rect -1908 -16950 -1850 -16938
rect -1908 -17526 -1896 -16950
rect -1862 -17526 -1850 -16950
rect -1908 -17538 -1850 -17526
rect -1796 -16950 -1738 -16938
rect -1796 -17526 -1784 -16950
rect -1750 -17526 -1738 -16950
rect -1796 -17538 -1738 -17526
rect -1668 -16950 -1610 -16938
rect -1668 -17526 -1656 -16950
rect -1622 -17526 -1610 -16950
rect -1668 -17538 -1610 -17526
rect -1556 -16950 -1498 -16938
rect -1556 -17526 -1544 -16950
rect -1510 -17526 -1498 -16950
rect -1556 -17538 -1498 -17526
rect -1428 -16950 -1370 -16938
rect -1428 -17526 -1416 -16950
rect -1382 -17526 -1370 -16950
rect -1428 -17538 -1370 -17526
rect -2276 -17758 -2218 -17746
rect -2276 -18334 -2264 -17758
rect -2230 -18334 -2218 -17758
rect -2276 -18346 -2218 -18334
rect -2148 -17758 -2090 -17746
rect -2148 -18334 -2136 -17758
rect -2102 -18334 -2090 -17758
rect -2148 -18346 -2090 -18334
rect -2036 -17758 -1978 -17746
rect -2036 -18334 -2024 -17758
rect -1990 -18334 -1978 -17758
rect -2036 -18346 -1978 -18334
rect -1908 -17758 -1850 -17746
rect -1908 -18334 -1896 -17758
rect -1862 -18334 -1850 -17758
rect -1908 -18346 -1850 -18334
rect -1796 -17758 -1738 -17746
rect -1796 -18334 -1784 -17758
rect -1750 -18334 -1738 -17758
rect -1796 -18346 -1738 -18334
rect -1668 -17758 -1610 -17746
rect -1668 -18334 -1656 -17758
rect -1622 -18334 -1610 -17758
rect -1668 -18346 -1610 -18334
rect -1556 -17758 -1498 -17746
rect -1556 -18334 -1544 -17758
rect -1510 -18334 -1498 -17758
rect -1556 -18346 -1498 -18334
rect -1428 -17758 -1370 -17746
rect -1428 -18334 -1416 -17758
rect -1382 -18334 -1370 -17758
rect -1428 -18346 -1370 -18334
<< pdiff >>
rect -15900 -8312 -15842 -8300
rect -15900 -9088 -15888 -8312
rect -15854 -9088 -15842 -8312
rect -15900 -9100 -15842 -9088
rect -15442 -8312 -15384 -8300
rect -15442 -9088 -15430 -8312
rect -15396 -9088 -15384 -8312
rect -15442 -9100 -15384 -9088
rect -15312 -8312 -15254 -8300
rect -15312 -9088 -15300 -8312
rect -15266 -9088 -15254 -8312
rect -15312 -9100 -15254 -9088
rect -14854 -8312 -14796 -8300
rect -14854 -9088 -14842 -8312
rect -14808 -9088 -14796 -8312
rect -14854 -9100 -14796 -9088
rect -14724 -8312 -14666 -8300
rect -14724 -9088 -14712 -8312
rect -14678 -9088 -14666 -8312
rect -14724 -9100 -14666 -9088
rect -14266 -8312 -14208 -8300
rect -14266 -9088 -14254 -8312
rect -14220 -9088 -14208 -8312
rect -14266 -9100 -14208 -9088
rect -14136 -8312 -14078 -8300
rect -14136 -9088 -14124 -8312
rect -14090 -9088 -14078 -8312
rect -14136 -9100 -14078 -9088
rect -13678 -8312 -13620 -8300
rect -13678 -9088 -13666 -8312
rect -13632 -9088 -13620 -8312
rect -13678 -9100 -13620 -9088
rect -13548 -8312 -13490 -8300
rect -13548 -9088 -13536 -8312
rect -13502 -9088 -13490 -8312
rect -13548 -9100 -13490 -9088
rect -13090 -8312 -13032 -8300
rect -13090 -9088 -13078 -8312
rect -13044 -9088 -13032 -8312
rect -13090 -9100 -13032 -9088
rect -12960 -8312 -12902 -8300
rect -12960 -9088 -12948 -8312
rect -12914 -9088 -12902 -8312
rect -12960 -9100 -12902 -9088
rect -12502 -8312 -12444 -8300
rect -12502 -9088 -12490 -8312
rect -12456 -9088 -12444 -8312
rect -12502 -9100 -12444 -9088
rect -12372 -8312 -12314 -8300
rect -12372 -9088 -12360 -8312
rect -12326 -9088 -12314 -8312
rect -12372 -9100 -12314 -9088
rect -11914 -8312 -11856 -8300
rect -11914 -9088 -11902 -8312
rect -11868 -9088 -11856 -8312
rect -11914 -9100 -11856 -9088
rect -11784 -8312 -11726 -8300
rect -11784 -9088 -11772 -8312
rect -11738 -9088 -11726 -8312
rect -11784 -9100 -11726 -9088
rect -11326 -8312 -11268 -8300
rect -11326 -9088 -11314 -8312
rect -11280 -9088 -11268 -8312
rect -11326 -9100 -11268 -9088
rect -11196 -8312 -11138 -8300
rect -11196 -9088 -11184 -8312
rect -11150 -9088 -11138 -8312
rect -11196 -9100 -11138 -9088
rect -10738 -8312 -10680 -8300
rect -10738 -9088 -10726 -8312
rect -10692 -9088 -10680 -8312
rect -10738 -9100 -10680 -9088
rect -10608 -8312 -10550 -8300
rect -10608 -9088 -10596 -8312
rect -10562 -9088 -10550 -8312
rect -10608 -9100 -10550 -9088
rect -10150 -8312 -10092 -8300
rect -10150 -9088 -10138 -8312
rect -10104 -9088 -10092 -8312
rect -10150 -9100 -10092 -9088
rect -10020 -8312 -9962 -8300
rect -10020 -9088 -10008 -8312
rect -9974 -9088 -9962 -8312
rect -10020 -9100 -9962 -9088
rect -9562 -8312 -9504 -8300
rect -9562 -9088 -9550 -8312
rect -9516 -9088 -9504 -8312
rect -9562 -9100 -9504 -9088
rect -9432 -8312 -9374 -8300
rect -9432 -9088 -9420 -8312
rect -9386 -9088 -9374 -8312
rect -9432 -9100 -9374 -9088
rect -8974 -8312 -8916 -8300
rect -8974 -9088 -8962 -8312
rect -8928 -9088 -8916 -8312
rect -8974 -9100 -8916 -9088
rect -8844 -8312 -8786 -8300
rect -8844 -9088 -8832 -8312
rect -8798 -9088 -8786 -8312
rect -8844 -9100 -8786 -9088
rect -8386 -8312 -8328 -8300
rect -8386 -9088 -8374 -8312
rect -8340 -9088 -8328 -8312
rect -8386 -9100 -8328 -9088
rect -8256 -8312 -8198 -8300
rect -8256 -9088 -8244 -8312
rect -8210 -9088 -8198 -8312
rect -8256 -9100 -8198 -9088
rect -7798 -8312 -7740 -8300
rect -7798 -9088 -7786 -8312
rect -7752 -9088 -7740 -8312
rect -7798 -9100 -7740 -9088
rect -7668 -8312 -7610 -8300
rect -7668 -9088 -7656 -8312
rect -7622 -9088 -7610 -8312
rect -7668 -9100 -7610 -9088
rect -7210 -8312 -7152 -8300
rect -7210 -9088 -7198 -8312
rect -7164 -9088 -7152 -8312
rect -7210 -9100 -7152 -9088
rect -7080 -8312 -7022 -8300
rect -7080 -9088 -7068 -8312
rect -7034 -9088 -7022 -8312
rect -7080 -9100 -7022 -9088
rect -6622 -8312 -6564 -8300
rect -6622 -9088 -6610 -8312
rect -6576 -9088 -6564 -8312
rect -6622 -9100 -6564 -9088
rect -6492 -8312 -6434 -8300
rect -6492 -9088 -6480 -8312
rect -6446 -9088 -6434 -8312
rect -6492 -9100 -6434 -9088
rect -6034 -8312 -5976 -8300
rect -6034 -9088 -6022 -8312
rect -5988 -9088 -5976 -8312
rect -6034 -9100 -5976 -9088
rect -5904 -8312 -5846 -8300
rect -5904 -9088 -5892 -8312
rect -5858 -9088 -5846 -8312
rect -5904 -9100 -5846 -9088
rect -5446 -8312 -5388 -8300
rect -5446 -9088 -5434 -8312
rect -5400 -9088 -5388 -8312
rect -5446 -9100 -5388 -9088
rect -5316 -8312 -5258 -8300
rect -5316 -9088 -5304 -8312
rect -5270 -9088 -5258 -8312
rect -5316 -9100 -5258 -9088
rect -4858 -8312 -4800 -8300
rect -4858 -9088 -4846 -8312
rect -4812 -9088 -4800 -8312
rect -4858 -9100 -4800 -9088
rect -4728 -8312 -4670 -8300
rect -4728 -9088 -4716 -8312
rect -4682 -9088 -4670 -8312
rect -4728 -9100 -4670 -9088
rect -4270 -8312 -4212 -8300
rect -4270 -9088 -4258 -8312
rect -4224 -9088 -4212 -8312
rect -4270 -9100 -4212 -9088
rect -4140 -8312 -4082 -8300
rect -4140 -9088 -4128 -8312
rect -4094 -9088 -4082 -8312
rect -4140 -9100 -4082 -9088
rect -3682 -8312 -3624 -8300
rect -3682 -9088 -3670 -8312
rect -3636 -9088 -3624 -8312
rect -3682 -9100 -3624 -9088
rect -3552 -8312 -3494 -8300
rect -3552 -9088 -3540 -8312
rect -3506 -9088 -3494 -8312
rect -3552 -9100 -3494 -9088
rect -3094 -8312 -3036 -8300
rect -3094 -9088 -3082 -8312
rect -3048 -9088 -3036 -8312
rect -3094 -9100 -3036 -9088
rect -2964 -8312 -2906 -8300
rect -2964 -9088 -2952 -8312
rect -2918 -9088 -2906 -8312
rect -2964 -9100 -2906 -9088
rect -2506 -8312 -2448 -8300
rect -2506 -9088 -2494 -8312
rect -2460 -9088 -2448 -8312
rect -2506 -9100 -2448 -9088
rect -2376 -8312 -2318 -8300
rect -2376 -9088 -2364 -8312
rect -2330 -9088 -2318 -8312
rect -2376 -9100 -2318 -9088
rect -1918 -8312 -1860 -8300
rect -1918 -9088 -1906 -8312
rect -1872 -9088 -1860 -8312
rect -1918 -9100 -1860 -9088
rect -1788 -8312 -1730 -8300
rect -1788 -9088 -1776 -8312
rect -1742 -9088 -1730 -8312
rect -1788 -9100 -1730 -9088
rect -1330 -8312 -1272 -8300
rect -1330 -9088 -1318 -8312
rect -1284 -9088 -1272 -8312
rect -1330 -9100 -1272 -9088
rect -1200 -8312 -1142 -8300
rect -1200 -9088 -1188 -8312
rect -1154 -9088 -1142 -8312
rect -1200 -9100 -1142 -9088
rect -742 -8312 -684 -8300
rect -742 -9088 -730 -8312
rect -696 -9088 -684 -8312
rect -742 -9100 -684 -9088
rect -612 -8312 -554 -8300
rect -612 -9088 -600 -8312
rect -566 -9088 -554 -8312
rect -612 -9100 -554 -9088
rect -154 -8312 -96 -8300
rect -154 -9088 -142 -8312
rect -108 -9088 -96 -8312
rect -154 -9100 -96 -9088
rect -24 -8312 34 -8300
rect -24 -9088 -12 -8312
rect 22 -9088 34 -8312
rect -24 -9100 34 -9088
rect 434 -8312 492 -8300
rect 434 -9088 446 -8312
rect 480 -9088 492 -8312
rect 434 -9100 492 -9088
rect 564 -8312 622 -8300
rect 564 -9088 576 -8312
rect 610 -9088 622 -8312
rect 564 -9100 622 -9088
rect 1022 -8312 1080 -8300
rect 1022 -9088 1034 -8312
rect 1068 -9088 1080 -8312
rect 1022 -9100 1080 -9088
rect 1152 -8312 1210 -8300
rect 1152 -9088 1164 -8312
rect 1198 -9088 1210 -8312
rect 1152 -9100 1210 -9088
rect 1610 -8312 1668 -8300
rect 1610 -9088 1622 -8312
rect 1656 -9088 1668 -8312
rect 1610 -9100 1668 -9088
rect 1740 -8312 1798 -8300
rect 1740 -9088 1752 -8312
rect 1786 -9088 1798 -8312
rect 1740 -9100 1798 -9088
rect 2198 -8312 2256 -8300
rect 2198 -9088 2210 -8312
rect 2244 -9088 2256 -8312
rect 2198 -9100 2256 -9088
rect 2328 -8312 2386 -8300
rect 2328 -9088 2340 -8312
rect 2374 -9088 2386 -8312
rect 2328 -9100 2386 -9088
rect 2786 -8312 2844 -8300
rect 2786 -9088 2798 -8312
rect 2832 -9088 2844 -8312
rect 2786 -9100 2844 -9088
rect 2916 -8312 2974 -8300
rect 2916 -9088 2928 -8312
rect 2962 -9088 2974 -8312
rect 2916 -9100 2974 -9088
rect 3374 -8312 3432 -8300
rect 3374 -9088 3386 -8312
rect 3420 -9088 3432 -8312
rect 3374 -9100 3432 -9088
rect 3504 -8312 3562 -8300
rect 3504 -9088 3516 -8312
rect 3550 -9088 3562 -8312
rect 3504 -9100 3562 -9088
rect 3962 -8312 4020 -8300
rect 3962 -9088 3974 -8312
rect 4008 -9088 4020 -8312
rect 3962 -9100 4020 -9088
rect 4092 -8312 4150 -8300
rect 4092 -9088 4104 -8312
rect 4138 -9088 4150 -8312
rect 4092 -9100 4150 -9088
rect 4550 -8312 4608 -8300
rect 4550 -9088 4562 -8312
rect 4596 -9088 4608 -8312
rect 4550 -9100 4608 -9088
rect 4680 -8312 4738 -8300
rect 4680 -9088 4692 -8312
rect 4726 -9088 4738 -8312
rect 4680 -9100 4738 -9088
rect 5138 -8312 5196 -8300
rect 5138 -9088 5150 -8312
rect 5184 -9088 5196 -8312
rect 5138 -9100 5196 -9088
rect 5268 -8312 5326 -8300
rect 5268 -9088 5280 -8312
rect 5314 -9088 5326 -8312
rect 5268 -9100 5326 -9088
rect 5726 -8312 5784 -8300
rect 5726 -9088 5738 -8312
rect 5772 -9088 5784 -8312
rect 5726 -9100 5784 -9088
rect 5856 -8312 5914 -8300
rect 5856 -9088 5868 -8312
rect 5902 -9088 5914 -8312
rect 5856 -9100 5914 -9088
rect 6314 -8312 6372 -8300
rect 6314 -9088 6326 -8312
rect 6360 -9088 6372 -8312
rect 6314 -9100 6372 -9088
rect 6444 -8312 6502 -8300
rect 6444 -9088 6456 -8312
rect 6490 -9088 6502 -8312
rect 6444 -9100 6502 -9088
rect 6902 -8312 6960 -8300
rect 6902 -9088 6914 -8312
rect 6948 -9088 6960 -8312
rect 6902 -9100 6960 -9088
rect 7032 -8312 7090 -8300
rect 7032 -9088 7044 -8312
rect 7078 -9088 7090 -8312
rect 7032 -9100 7090 -9088
rect 7490 -8312 7548 -8300
rect 7490 -9088 7502 -8312
rect 7536 -9088 7548 -8312
rect 7490 -9100 7548 -9088
rect 7620 -8312 7678 -8300
rect 7620 -9088 7632 -8312
rect 7666 -9088 7678 -8312
rect 7620 -9100 7678 -9088
rect 8078 -8312 8136 -8300
rect 8078 -9088 8090 -8312
rect 8124 -9088 8136 -8312
rect 8078 -9100 8136 -9088
rect 8208 -8312 8266 -8300
rect 8208 -9088 8220 -8312
rect 8254 -9088 8266 -8312
rect 8208 -9100 8266 -9088
rect 8666 -8312 8724 -8300
rect 8666 -9088 8678 -8312
rect 8712 -9088 8724 -8312
rect 8666 -9100 8724 -9088
rect 8796 -8312 8854 -8300
rect 8796 -9088 8808 -8312
rect 8842 -9088 8854 -8312
rect 8796 -9100 8854 -9088
rect 9254 -8312 9312 -8300
rect 9254 -9088 9266 -8312
rect 9300 -9088 9312 -8312
rect 9254 -9100 9312 -9088
rect 9384 -8312 9442 -8300
rect 9384 -9088 9396 -8312
rect 9430 -9088 9442 -8312
rect 9384 -9100 9442 -9088
rect 9842 -8312 9900 -8300
rect 9842 -9088 9854 -8312
rect 9888 -9088 9900 -8312
rect 9842 -9100 9900 -9088
rect 9972 -8312 10030 -8300
rect 9972 -9088 9984 -8312
rect 10018 -9088 10030 -8312
rect 9972 -9100 10030 -9088
rect 10430 -8312 10488 -8300
rect 10430 -9088 10442 -8312
rect 10476 -9088 10488 -8312
rect 10430 -9100 10488 -9088
rect 10560 -8312 10618 -8300
rect 10560 -9088 10572 -8312
rect 10606 -9088 10618 -8312
rect 10560 -9100 10618 -9088
rect 11018 -8312 11076 -8300
rect 11018 -9088 11030 -8312
rect 11064 -9088 11076 -8312
rect 11018 -9100 11076 -9088
rect 11148 -8312 11206 -8300
rect 11148 -9088 11160 -8312
rect 11194 -9088 11206 -8312
rect 11148 -9100 11206 -9088
rect 11606 -8312 11664 -8300
rect 11606 -9088 11618 -8312
rect 11652 -9088 11664 -8312
rect 11606 -9100 11664 -9088
rect 11736 -8312 11794 -8300
rect 11736 -9088 11748 -8312
rect 11782 -9088 11794 -8312
rect 11736 -9100 11794 -9088
rect 12194 -8312 12252 -8300
rect 12194 -9088 12206 -8312
rect 12240 -9088 12252 -8312
rect 12194 -9100 12252 -9088
rect -15900 -9312 -15842 -9300
rect -15900 -10088 -15888 -9312
rect -15854 -10088 -15842 -9312
rect -15900 -10100 -15842 -10088
rect -15442 -9312 -15384 -9300
rect -15442 -10088 -15430 -9312
rect -15396 -10088 -15384 -9312
rect -15442 -10100 -15384 -10088
rect -15312 -9312 -15254 -9300
rect -15312 -10088 -15300 -9312
rect -15266 -10088 -15254 -9312
rect -15312 -10100 -15254 -10088
rect -14854 -9312 -14796 -9300
rect -14854 -10088 -14842 -9312
rect -14808 -10088 -14796 -9312
rect -14854 -10100 -14796 -10088
rect -14724 -9312 -14666 -9300
rect -14724 -10088 -14712 -9312
rect -14678 -10088 -14666 -9312
rect -14724 -10100 -14666 -10088
rect -14266 -9312 -14208 -9300
rect -14266 -10088 -14254 -9312
rect -14220 -10088 -14208 -9312
rect -14266 -10100 -14208 -10088
rect -14136 -9312 -14078 -9300
rect -14136 -10088 -14124 -9312
rect -14090 -10088 -14078 -9312
rect -14136 -10100 -14078 -10088
rect -13678 -9312 -13620 -9300
rect -13678 -10088 -13666 -9312
rect -13632 -10088 -13620 -9312
rect -13678 -10100 -13620 -10088
rect -13548 -9312 -13490 -9300
rect -13548 -10088 -13536 -9312
rect -13502 -10088 -13490 -9312
rect -13548 -10100 -13490 -10088
rect -13090 -9312 -13032 -9300
rect -13090 -10088 -13078 -9312
rect -13044 -10088 -13032 -9312
rect -13090 -10100 -13032 -10088
rect -12960 -9312 -12902 -9300
rect -12960 -10088 -12948 -9312
rect -12914 -10088 -12902 -9312
rect -12960 -10100 -12902 -10088
rect -12502 -9312 -12444 -9300
rect -12502 -10088 -12490 -9312
rect -12456 -10088 -12444 -9312
rect -12502 -10100 -12444 -10088
rect -12372 -9312 -12314 -9300
rect -12372 -10088 -12360 -9312
rect -12326 -10088 -12314 -9312
rect -12372 -10100 -12314 -10088
rect -11914 -9312 -11856 -9300
rect -11914 -10088 -11902 -9312
rect -11868 -10088 -11856 -9312
rect -11914 -10100 -11856 -10088
rect -11784 -9312 -11726 -9300
rect -11784 -10088 -11772 -9312
rect -11738 -10088 -11726 -9312
rect -11784 -10100 -11726 -10088
rect -11326 -9312 -11268 -9300
rect -11326 -10088 -11314 -9312
rect -11280 -10088 -11268 -9312
rect -11326 -10100 -11268 -10088
rect -11196 -9312 -11138 -9300
rect -11196 -10088 -11184 -9312
rect -11150 -10088 -11138 -9312
rect -11196 -10100 -11138 -10088
rect -10738 -9312 -10680 -9300
rect -10738 -10088 -10726 -9312
rect -10692 -10088 -10680 -9312
rect -10738 -10100 -10680 -10088
rect -10608 -9312 -10550 -9300
rect -10608 -10088 -10596 -9312
rect -10562 -10088 -10550 -9312
rect -10608 -10100 -10550 -10088
rect -10150 -9312 -10092 -9300
rect -10150 -10088 -10138 -9312
rect -10104 -10088 -10092 -9312
rect -10150 -10100 -10092 -10088
rect -10020 -9312 -9962 -9300
rect -10020 -10088 -10008 -9312
rect -9974 -10088 -9962 -9312
rect -10020 -10100 -9962 -10088
rect -9562 -9312 -9504 -9300
rect -9562 -10088 -9550 -9312
rect -9516 -10088 -9504 -9312
rect -9562 -10100 -9504 -10088
rect -9432 -9312 -9374 -9300
rect -9432 -10088 -9420 -9312
rect -9386 -10088 -9374 -9312
rect -9432 -10100 -9374 -10088
rect -8974 -9312 -8916 -9300
rect -8974 -10088 -8962 -9312
rect -8928 -10088 -8916 -9312
rect -8974 -10100 -8916 -10088
rect -8844 -9312 -8786 -9300
rect -8844 -10088 -8832 -9312
rect -8798 -10088 -8786 -9312
rect -8844 -10100 -8786 -10088
rect -8386 -9312 -8328 -9300
rect -8386 -10088 -8374 -9312
rect -8340 -10088 -8328 -9312
rect -8386 -10100 -8328 -10088
rect -8256 -9312 -8198 -9300
rect -8256 -10088 -8244 -9312
rect -8210 -10088 -8198 -9312
rect -8256 -10100 -8198 -10088
rect -7798 -9312 -7740 -9300
rect -7798 -10088 -7786 -9312
rect -7752 -10088 -7740 -9312
rect -7798 -10100 -7740 -10088
rect -7668 -9312 -7610 -9300
rect -7668 -10088 -7656 -9312
rect -7622 -10088 -7610 -9312
rect -7668 -10100 -7610 -10088
rect -7210 -9312 -7152 -9300
rect -7210 -10088 -7198 -9312
rect -7164 -10088 -7152 -9312
rect -7210 -10100 -7152 -10088
rect -7080 -9312 -7022 -9300
rect -7080 -10088 -7068 -9312
rect -7034 -10088 -7022 -9312
rect -7080 -10100 -7022 -10088
rect -6622 -9312 -6564 -9300
rect -6622 -10088 -6610 -9312
rect -6576 -10088 -6564 -9312
rect -6622 -10100 -6564 -10088
rect -6492 -9312 -6434 -9300
rect -6492 -10088 -6480 -9312
rect -6446 -10088 -6434 -9312
rect -6492 -10100 -6434 -10088
rect -6034 -9312 -5976 -9300
rect -6034 -10088 -6022 -9312
rect -5988 -10088 -5976 -9312
rect -6034 -10100 -5976 -10088
rect -5904 -9312 -5846 -9300
rect -5904 -10088 -5892 -9312
rect -5858 -10088 -5846 -9312
rect -5904 -10100 -5846 -10088
rect -5446 -9312 -5388 -9300
rect -5446 -10088 -5434 -9312
rect -5400 -10088 -5388 -9312
rect -5446 -10100 -5388 -10088
rect -5316 -9312 -5258 -9300
rect -5316 -10088 -5304 -9312
rect -5270 -10088 -5258 -9312
rect -5316 -10100 -5258 -10088
rect -4858 -9312 -4800 -9300
rect -4858 -10088 -4846 -9312
rect -4812 -10088 -4800 -9312
rect -4858 -10100 -4800 -10088
rect -4728 -9312 -4670 -9300
rect -4728 -10088 -4716 -9312
rect -4682 -10088 -4670 -9312
rect -4728 -10100 -4670 -10088
rect -4270 -9312 -4212 -9300
rect -4270 -10088 -4258 -9312
rect -4224 -10088 -4212 -9312
rect -4270 -10100 -4212 -10088
rect -4140 -9312 -4082 -9300
rect -4140 -10088 -4128 -9312
rect -4094 -10088 -4082 -9312
rect -4140 -10100 -4082 -10088
rect -3682 -9312 -3624 -9300
rect -3682 -10088 -3670 -9312
rect -3636 -10088 -3624 -9312
rect -3682 -10100 -3624 -10088
rect -3552 -9312 -3494 -9300
rect -3552 -10088 -3540 -9312
rect -3506 -10088 -3494 -9312
rect -3552 -10100 -3494 -10088
rect -3094 -9312 -3036 -9300
rect -3094 -10088 -3082 -9312
rect -3048 -10088 -3036 -9312
rect -3094 -10100 -3036 -10088
rect -2964 -9312 -2906 -9300
rect -2964 -10088 -2952 -9312
rect -2918 -10088 -2906 -9312
rect -2964 -10100 -2906 -10088
rect -2506 -9312 -2448 -9300
rect -2506 -10088 -2494 -9312
rect -2460 -10088 -2448 -9312
rect -2506 -10100 -2448 -10088
rect -2376 -9312 -2318 -9300
rect -2376 -10088 -2364 -9312
rect -2330 -10088 -2318 -9312
rect -2376 -10100 -2318 -10088
rect -1918 -9312 -1860 -9300
rect -1918 -10088 -1906 -9312
rect -1872 -10088 -1860 -9312
rect -1918 -10100 -1860 -10088
rect -1788 -9312 -1730 -9300
rect -1788 -10088 -1776 -9312
rect -1742 -10088 -1730 -9312
rect -1788 -10100 -1730 -10088
rect -1330 -9312 -1272 -9300
rect -1330 -10088 -1318 -9312
rect -1284 -10088 -1272 -9312
rect -1330 -10100 -1272 -10088
rect -1200 -9312 -1142 -9300
rect -1200 -10088 -1188 -9312
rect -1154 -10088 -1142 -9312
rect -1200 -10100 -1142 -10088
rect -742 -9312 -684 -9300
rect -742 -10088 -730 -9312
rect -696 -10088 -684 -9312
rect -742 -10100 -684 -10088
rect -612 -9312 -554 -9300
rect -612 -10088 -600 -9312
rect -566 -10088 -554 -9312
rect -612 -10100 -554 -10088
rect -154 -9312 -96 -9300
rect -154 -10088 -142 -9312
rect -108 -10088 -96 -9312
rect -154 -10100 -96 -10088
rect -24 -9312 34 -9300
rect -24 -10088 -12 -9312
rect 22 -10088 34 -9312
rect -24 -10100 34 -10088
rect 434 -9312 492 -9300
rect 434 -10088 446 -9312
rect 480 -10088 492 -9312
rect 434 -10100 492 -10088
rect 564 -9312 622 -9300
rect 564 -10088 576 -9312
rect 610 -10088 622 -9312
rect 564 -10100 622 -10088
rect 1022 -9312 1080 -9300
rect 1022 -10088 1034 -9312
rect 1068 -10088 1080 -9312
rect 1022 -10100 1080 -10088
rect 1152 -9312 1210 -9300
rect 1152 -10088 1164 -9312
rect 1198 -10088 1210 -9312
rect 1152 -10100 1210 -10088
rect 1610 -9312 1668 -9300
rect 1610 -10088 1622 -9312
rect 1656 -10088 1668 -9312
rect 1610 -10100 1668 -10088
rect 1740 -9312 1798 -9300
rect 1740 -10088 1752 -9312
rect 1786 -10088 1798 -9312
rect 1740 -10100 1798 -10088
rect 2198 -9312 2256 -9300
rect 2198 -10088 2210 -9312
rect 2244 -10088 2256 -9312
rect 2198 -10100 2256 -10088
rect 2328 -9312 2386 -9300
rect 2328 -10088 2340 -9312
rect 2374 -10088 2386 -9312
rect 2328 -10100 2386 -10088
rect 2786 -9312 2844 -9300
rect 2786 -10088 2798 -9312
rect 2832 -10088 2844 -9312
rect 2786 -10100 2844 -10088
rect 2916 -9312 2974 -9300
rect 2916 -10088 2928 -9312
rect 2962 -10088 2974 -9312
rect 2916 -10100 2974 -10088
rect 3374 -9312 3432 -9300
rect 3374 -10088 3386 -9312
rect 3420 -10088 3432 -9312
rect 3374 -10100 3432 -10088
rect 3504 -9312 3562 -9300
rect 3504 -10088 3516 -9312
rect 3550 -10088 3562 -9312
rect 3504 -10100 3562 -10088
rect 3962 -9312 4020 -9300
rect 3962 -10088 3974 -9312
rect 4008 -10088 4020 -9312
rect 3962 -10100 4020 -10088
rect 4092 -9312 4150 -9300
rect 4092 -10088 4104 -9312
rect 4138 -10088 4150 -9312
rect 4092 -10100 4150 -10088
rect 4550 -9312 4608 -9300
rect 4550 -10088 4562 -9312
rect 4596 -10088 4608 -9312
rect 4550 -10100 4608 -10088
rect 4680 -9312 4738 -9300
rect 4680 -10088 4692 -9312
rect 4726 -10088 4738 -9312
rect 4680 -10100 4738 -10088
rect 5138 -9312 5196 -9300
rect 5138 -10088 5150 -9312
rect 5184 -10088 5196 -9312
rect 5138 -10100 5196 -10088
rect 5268 -9312 5326 -9300
rect 5268 -10088 5280 -9312
rect 5314 -10088 5326 -9312
rect 5268 -10100 5326 -10088
rect 5726 -9312 5784 -9300
rect 5726 -10088 5738 -9312
rect 5772 -10088 5784 -9312
rect 5726 -10100 5784 -10088
rect 5856 -9312 5914 -9300
rect 5856 -10088 5868 -9312
rect 5902 -10088 5914 -9312
rect 5856 -10100 5914 -10088
rect 6314 -9312 6372 -9300
rect 6314 -10088 6326 -9312
rect 6360 -10088 6372 -9312
rect 6314 -10100 6372 -10088
rect 6444 -9312 6502 -9300
rect 6444 -10088 6456 -9312
rect 6490 -10088 6502 -9312
rect 6444 -10100 6502 -10088
rect 6902 -9312 6960 -9300
rect 6902 -10088 6914 -9312
rect 6948 -10088 6960 -9312
rect 6902 -10100 6960 -10088
rect 7032 -9312 7090 -9300
rect 7032 -10088 7044 -9312
rect 7078 -10088 7090 -9312
rect 7032 -10100 7090 -10088
rect 7490 -9312 7548 -9300
rect 7490 -10088 7502 -9312
rect 7536 -10088 7548 -9312
rect 7490 -10100 7548 -10088
rect 7620 -9312 7678 -9300
rect 7620 -10088 7632 -9312
rect 7666 -10088 7678 -9312
rect 7620 -10100 7678 -10088
rect 8078 -9312 8136 -9300
rect 8078 -10088 8090 -9312
rect 8124 -10088 8136 -9312
rect 8078 -10100 8136 -10088
rect 8208 -9312 8266 -9300
rect 8208 -10088 8220 -9312
rect 8254 -10088 8266 -9312
rect 8208 -10100 8266 -10088
rect 8666 -9312 8724 -9300
rect 8666 -10088 8678 -9312
rect 8712 -10088 8724 -9312
rect 8666 -10100 8724 -10088
rect 8796 -9312 8854 -9300
rect 8796 -10088 8808 -9312
rect 8842 -10088 8854 -9312
rect 8796 -10100 8854 -10088
rect 9254 -9312 9312 -9300
rect 9254 -10088 9266 -9312
rect 9300 -10088 9312 -9312
rect 9254 -10100 9312 -10088
rect 9384 -9312 9442 -9300
rect 9384 -10088 9396 -9312
rect 9430 -10088 9442 -9312
rect 9384 -10100 9442 -10088
rect 9842 -9312 9900 -9300
rect 9842 -10088 9854 -9312
rect 9888 -10088 9900 -9312
rect 9842 -10100 9900 -10088
rect 9972 -9312 10030 -9300
rect 9972 -10088 9984 -9312
rect 10018 -10088 10030 -9312
rect 9972 -10100 10030 -10088
rect 10430 -9312 10488 -9300
rect 10430 -10088 10442 -9312
rect 10476 -10088 10488 -9312
rect 10430 -10100 10488 -10088
rect 10560 -9312 10618 -9300
rect 10560 -10088 10572 -9312
rect 10606 -10088 10618 -9312
rect 10560 -10100 10618 -10088
rect 11018 -9312 11076 -9300
rect 11018 -10088 11030 -9312
rect 11064 -10088 11076 -9312
rect 11018 -10100 11076 -10088
rect 11148 -9312 11206 -9300
rect 11148 -10088 11160 -9312
rect 11194 -10088 11206 -9312
rect 11148 -10100 11206 -10088
rect 11606 -9312 11664 -9300
rect 11606 -10088 11618 -9312
rect 11652 -10088 11664 -9312
rect 11606 -10100 11664 -10088
rect 11736 -9312 11794 -9300
rect 11736 -10088 11748 -9312
rect 11782 -10088 11794 -9312
rect 11736 -10100 11794 -10088
rect 12194 -9312 12252 -9300
rect 12194 -10088 12206 -9312
rect 12240 -10088 12252 -9312
rect 12194 -10100 12252 -10088
rect -15900 -10312 -15842 -10300
rect -15900 -11088 -15888 -10312
rect -15854 -11088 -15842 -10312
rect -15900 -11100 -15842 -11088
rect -15442 -10312 -15384 -10300
rect -15442 -11088 -15430 -10312
rect -15396 -11088 -15384 -10312
rect -15442 -11100 -15384 -11088
rect -15312 -10312 -15254 -10300
rect -15312 -11088 -15300 -10312
rect -15266 -11088 -15254 -10312
rect -15312 -11100 -15254 -11088
rect -14854 -10312 -14796 -10300
rect -14854 -11088 -14842 -10312
rect -14808 -11088 -14796 -10312
rect -14854 -11100 -14796 -11088
rect -14724 -10312 -14666 -10300
rect -14724 -11088 -14712 -10312
rect -14678 -11088 -14666 -10312
rect -14724 -11100 -14666 -11088
rect -14266 -10312 -14208 -10300
rect -14266 -11088 -14254 -10312
rect -14220 -11088 -14208 -10312
rect -14266 -11100 -14208 -11088
rect -14136 -10312 -14078 -10300
rect -14136 -11088 -14124 -10312
rect -14090 -11088 -14078 -10312
rect -14136 -11100 -14078 -11088
rect -13678 -10312 -13620 -10300
rect -13678 -11088 -13666 -10312
rect -13632 -11088 -13620 -10312
rect -13678 -11100 -13620 -11088
rect -13548 -10312 -13490 -10300
rect -13548 -11088 -13536 -10312
rect -13502 -11088 -13490 -10312
rect -13548 -11100 -13490 -11088
rect -13090 -10312 -13032 -10300
rect -13090 -11088 -13078 -10312
rect -13044 -11088 -13032 -10312
rect -13090 -11100 -13032 -11088
rect -12960 -10312 -12902 -10300
rect -12960 -11088 -12948 -10312
rect -12914 -11088 -12902 -10312
rect -12960 -11100 -12902 -11088
rect -12502 -10312 -12444 -10300
rect -12502 -11088 -12490 -10312
rect -12456 -11088 -12444 -10312
rect -12502 -11100 -12444 -11088
rect -12372 -10312 -12314 -10300
rect -12372 -11088 -12360 -10312
rect -12326 -11088 -12314 -10312
rect -12372 -11100 -12314 -11088
rect -11914 -10312 -11856 -10300
rect -11914 -11088 -11902 -10312
rect -11868 -11088 -11856 -10312
rect -11914 -11100 -11856 -11088
rect -11784 -10312 -11726 -10300
rect -11784 -11088 -11772 -10312
rect -11738 -11088 -11726 -10312
rect -11784 -11100 -11726 -11088
rect -11326 -10312 -11268 -10300
rect -11326 -11088 -11314 -10312
rect -11280 -11088 -11268 -10312
rect -11326 -11100 -11268 -11088
rect -11196 -10312 -11138 -10300
rect -11196 -11088 -11184 -10312
rect -11150 -11088 -11138 -10312
rect -11196 -11100 -11138 -11088
rect -10738 -10312 -10680 -10300
rect -10738 -11088 -10726 -10312
rect -10692 -11088 -10680 -10312
rect -10738 -11100 -10680 -11088
rect -10608 -10312 -10550 -10300
rect -10608 -11088 -10596 -10312
rect -10562 -11088 -10550 -10312
rect -10608 -11100 -10550 -11088
rect -10150 -10312 -10092 -10300
rect -10150 -11088 -10138 -10312
rect -10104 -11088 -10092 -10312
rect -10150 -11100 -10092 -11088
rect -10020 -10312 -9962 -10300
rect -10020 -11088 -10008 -10312
rect -9974 -11088 -9962 -10312
rect -10020 -11100 -9962 -11088
rect -9562 -10312 -9504 -10300
rect -9562 -11088 -9550 -10312
rect -9516 -11088 -9504 -10312
rect -9562 -11100 -9504 -11088
rect -9432 -10312 -9374 -10300
rect -9432 -11088 -9420 -10312
rect -9386 -11088 -9374 -10312
rect -9432 -11100 -9374 -11088
rect -8974 -10312 -8916 -10300
rect -8974 -11088 -8962 -10312
rect -8928 -11088 -8916 -10312
rect -8974 -11100 -8916 -11088
rect -8844 -10312 -8786 -10300
rect -8844 -11088 -8832 -10312
rect -8798 -11088 -8786 -10312
rect -8844 -11100 -8786 -11088
rect -8386 -10312 -8328 -10300
rect -8386 -11088 -8374 -10312
rect -8340 -11088 -8328 -10312
rect -8386 -11100 -8328 -11088
rect -8256 -10312 -8198 -10300
rect -8256 -11088 -8244 -10312
rect -8210 -11088 -8198 -10312
rect -8256 -11100 -8198 -11088
rect -7798 -10312 -7740 -10300
rect -7798 -11088 -7786 -10312
rect -7752 -11088 -7740 -10312
rect -7798 -11100 -7740 -11088
rect -7668 -10312 -7610 -10300
rect -7668 -11088 -7656 -10312
rect -7622 -11088 -7610 -10312
rect -7668 -11100 -7610 -11088
rect -7210 -10312 -7152 -10300
rect -7210 -11088 -7198 -10312
rect -7164 -11088 -7152 -10312
rect -7210 -11100 -7152 -11088
rect -7080 -10312 -7022 -10300
rect -7080 -11088 -7068 -10312
rect -7034 -11088 -7022 -10312
rect -7080 -11100 -7022 -11088
rect -6622 -10312 -6564 -10300
rect -6622 -11088 -6610 -10312
rect -6576 -11088 -6564 -10312
rect -6622 -11100 -6564 -11088
rect -6492 -10312 -6434 -10300
rect -6492 -11088 -6480 -10312
rect -6446 -11088 -6434 -10312
rect -6492 -11100 -6434 -11088
rect -6034 -10312 -5976 -10300
rect -6034 -11088 -6022 -10312
rect -5988 -11088 -5976 -10312
rect -6034 -11100 -5976 -11088
rect -5904 -10312 -5846 -10300
rect -5904 -11088 -5892 -10312
rect -5858 -11088 -5846 -10312
rect -5904 -11100 -5846 -11088
rect -5446 -10312 -5388 -10300
rect -5446 -11088 -5434 -10312
rect -5400 -11088 -5388 -10312
rect -5446 -11100 -5388 -11088
rect -5316 -10312 -5258 -10300
rect -5316 -11088 -5304 -10312
rect -5270 -11088 -5258 -10312
rect -5316 -11100 -5258 -11088
rect -4858 -10312 -4800 -10300
rect -4858 -11088 -4846 -10312
rect -4812 -11088 -4800 -10312
rect -4858 -11100 -4800 -11088
rect -4728 -10312 -4670 -10300
rect -4728 -11088 -4716 -10312
rect -4682 -11088 -4670 -10312
rect -4728 -11100 -4670 -11088
rect -4270 -10312 -4212 -10300
rect -4270 -11088 -4258 -10312
rect -4224 -11088 -4212 -10312
rect -4270 -11100 -4212 -11088
rect -4140 -10312 -4082 -10300
rect -4140 -11088 -4128 -10312
rect -4094 -11088 -4082 -10312
rect -4140 -11100 -4082 -11088
rect -3682 -10312 -3624 -10300
rect -3682 -11088 -3670 -10312
rect -3636 -11088 -3624 -10312
rect -3682 -11100 -3624 -11088
rect -3552 -10312 -3494 -10300
rect -3552 -11088 -3540 -10312
rect -3506 -11088 -3494 -10312
rect -3552 -11100 -3494 -11088
rect -3094 -10312 -3036 -10300
rect -3094 -11088 -3082 -10312
rect -3048 -11088 -3036 -10312
rect -3094 -11100 -3036 -11088
rect -2964 -10312 -2906 -10300
rect -2964 -11088 -2952 -10312
rect -2918 -11088 -2906 -10312
rect -2964 -11100 -2906 -11088
rect -2506 -10312 -2448 -10300
rect -2506 -11088 -2494 -10312
rect -2460 -11088 -2448 -10312
rect -2506 -11100 -2448 -11088
rect -2376 -10312 -2318 -10300
rect -2376 -11088 -2364 -10312
rect -2330 -11088 -2318 -10312
rect -2376 -11100 -2318 -11088
rect -1918 -10312 -1860 -10300
rect -1918 -11088 -1906 -10312
rect -1872 -11088 -1860 -10312
rect -1918 -11100 -1860 -11088
rect -1788 -10312 -1730 -10300
rect -1788 -11088 -1776 -10312
rect -1742 -11088 -1730 -10312
rect -1788 -11100 -1730 -11088
rect -1330 -10312 -1272 -10300
rect -1330 -11088 -1318 -10312
rect -1284 -11088 -1272 -10312
rect -1330 -11100 -1272 -11088
rect -1200 -10312 -1142 -10300
rect -1200 -11088 -1188 -10312
rect -1154 -11088 -1142 -10312
rect -1200 -11100 -1142 -11088
rect -742 -10312 -684 -10300
rect -742 -11088 -730 -10312
rect -696 -11088 -684 -10312
rect -742 -11100 -684 -11088
rect -612 -10312 -554 -10300
rect -612 -11088 -600 -10312
rect -566 -11088 -554 -10312
rect -612 -11100 -554 -11088
rect -154 -10312 -96 -10300
rect -154 -11088 -142 -10312
rect -108 -11088 -96 -10312
rect -154 -11100 -96 -11088
rect -24 -10312 34 -10300
rect -24 -11088 -12 -10312
rect 22 -11088 34 -10312
rect -24 -11100 34 -11088
rect 434 -10312 492 -10300
rect 434 -11088 446 -10312
rect 480 -11088 492 -10312
rect 434 -11100 492 -11088
rect 564 -10312 622 -10300
rect 564 -11088 576 -10312
rect 610 -11088 622 -10312
rect 564 -11100 622 -11088
rect 1022 -10312 1080 -10300
rect 1022 -11088 1034 -10312
rect 1068 -11088 1080 -10312
rect 1022 -11100 1080 -11088
rect 1152 -10312 1210 -10300
rect 1152 -11088 1164 -10312
rect 1198 -11088 1210 -10312
rect 1152 -11100 1210 -11088
rect 1610 -10312 1668 -10300
rect 1610 -11088 1622 -10312
rect 1656 -11088 1668 -10312
rect 1610 -11100 1668 -11088
rect 1740 -10312 1798 -10300
rect 1740 -11088 1752 -10312
rect 1786 -11088 1798 -10312
rect 1740 -11100 1798 -11088
rect 2198 -10312 2256 -10300
rect 2198 -11088 2210 -10312
rect 2244 -11088 2256 -10312
rect 2198 -11100 2256 -11088
rect 2328 -10312 2386 -10300
rect 2328 -11088 2340 -10312
rect 2374 -11088 2386 -10312
rect 2328 -11100 2386 -11088
rect 2786 -10312 2844 -10300
rect 2786 -11088 2798 -10312
rect 2832 -11088 2844 -10312
rect 2786 -11100 2844 -11088
rect 2916 -10312 2974 -10300
rect 2916 -11088 2928 -10312
rect 2962 -11088 2974 -10312
rect 2916 -11100 2974 -11088
rect 3374 -10312 3432 -10300
rect 3374 -11088 3386 -10312
rect 3420 -11088 3432 -10312
rect 3374 -11100 3432 -11088
rect 3504 -10312 3562 -10300
rect 3504 -11088 3516 -10312
rect 3550 -11088 3562 -10312
rect 3504 -11100 3562 -11088
rect 3962 -10312 4020 -10300
rect 3962 -11088 3974 -10312
rect 4008 -11088 4020 -10312
rect 3962 -11100 4020 -11088
rect 4092 -10312 4150 -10300
rect 4092 -11088 4104 -10312
rect 4138 -11088 4150 -10312
rect 4092 -11100 4150 -11088
rect 4550 -10312 4608 -10300
rect 4550 -11088 4562 -10312
rect 4596 -11088 4608 -10312
rect 4550 -11100 4608 -11088
rect 4680 -10312 4738 -10300
rect 4680 -11088 4692 -10312
rect 4726 -11088 4738 -10312
rect 4680 -11100 4738 -11088
rect 5138 -10312 5196 -10300
rect 5138 -11088 5150 -10312
rect 5184 -11088 5196 -10312
rect 5138 -11100 5196 -11088
rect 5268 -10312 5326 -10300
rect 5268 -11088 5280 -10312
rect 5314 -11088 5326 -10312
rect 5268 -11100 5326 -11088
rect 5726 -10312 5784 -10300
rect 5726 -11088 5738 -10312
rect 5772 -11088 5784 -10312
rect 5726 -11100 5784 -11088
rect 5856 -10312 5914 -10300
rect 5856 -11088 5868 -10312
rect 5902 -11088 5914 -10312
rect 5856 -11100 5914 -11088
rect 6314 -10312 6372 -10300
rect 6314 -11088 6326 -10312
rect 6360 -11088 6372 -10312
rect 6314 -11100 6372 -11088
rect 6444 -10312 6502 -10300
rect 6444 -11088 6456 -10312
rect 6490 -11088 6502 -10312
rect 6444 -11100 6502 -11088
rect 6902 -10312 6960 -10300
rect 6902 -11088 6914 -10312
rect 6948 -11088 6960 -10312
rect 6902 -11100 6960 -11088
rect 7032 -10312 7090 -10300
rect 7032 -11088 7044 -10312
rect 7078 -11088 7090 -10312
rect 7032 -11100 7090 -11088
rect 7490 -10312 7548 -10300
rect 7490 -11088 7502 -10312
rect 7536 -11088 7548 -10312
rect 7490 -11100 7548 -11088
rect 7620 -10312 7678 -10300
rect 7620 -11088 7632 -10312
rect 7666 -11088 7678 -10312
rect 7620 -11100 7678 -11088
rect 8078 -10312 8136 -10300
rect 8078 -11088 8090 -10312
rect 8124 -11088 8136 -10312
rect 8078 -11100 8136 -11088
rect 8208 -10312 8266 -10300
rect 8208 -11088 8220 -10312
rect 8254 -11088 8266 -10312
rect 8208 -11100 8266 -11088
rect 8666 -10312 8724 -10300
rect 8666 -11088 8678 -10312
rect 8712 -11088 8724 -10312
rect 8666 -11100 8724 -11088
rect 8796 -10312 8854 -10300
rect 8796 -11088 8808 -10312
rect 8842 -11088 8854 -10312
rect 8796 -11100 8854 -11088
rect 9254 -10312 9312 -10300
rect 9254 -11088 9266 -10312
rect 9300 -11088 9312 -10312
rect 9254 -11100 9312 -11088
rect 9384 -10312 9442 -10300
rect 9384 -11088 9396 -10312
rect 9430 -11088 9442 -10312
rect 9384 -11100 9442 -11088
rect 9842 -10312 9900 -10300
rect 9842 -11088 9854 -10312
rect 9888 -11088 9900 -10312
rect 9842 -11100 9900 -11088
rect 9972 -10312 10030 -10300
rect 9972 -11088 9984 -10312
rect 10018 -11088 10030 -10312
rect 9972 -11100 10030 -11088
rect 10430 -10312 10488 -10300
rect 10430 -11088 10442 -10312
rect 10476 -11088 10488 -10312
rect 10430 -11100 10488 -11088
rect 10560 -10312 10618 -10300
rect 10560 -11088 10572 -10312
rect 10606 -11088 10618 -10312
rect 10560 -11100 10618 -11088
rect 11018 -10312 11076 -10300
rect 11018 -11088 11030 -10312
rect 11064 -11088 11076 -10312
rect 11018 -11100 11076 -11088
rect 11148 -10312 11206 -10300
rect 11148 -11088 11160 -10312
rect 11194 -11088 11206 -10312
rect 11148 -11100 11206 -11088
rect 11606 -10312 11664 -10300
rect 11606 -11088 11618 -10312
rect 11652 -11088 11664 -10312
rect 11606 -11100 11664 -11088
rect 11736 -10312 11794 -10300
rect 11736 -11088 11748 -10312
rect 11782 -11088 11794 -10312
rect 11736 -11100 11794 -11088
rect 12194 -10312 12252 -10300
rect 12194 -11088 12206 -10312
rect 12240 -11088 12252 -10312
rect 12194 -11100 12252 -11088
rect -2848 -12758 -2790 -12746
rect -2848 -13534 -2836 -12758
rect -2802 -13534 -2790 -12758
rect -2848 -13546 -2790 -13534
rect -2720 -12758 -2662 -12746
rect -2720 -13534 -2708 -12758
rect -2674 -13534 -2662 -12758
rect -2720 -13546 -2662 -13534
rect -2582 -12758 -2524 -12746
rect -2582 -13534 -2570 -12758
rect -2536 -13534 -2524 -12758
rect -2582 -13546 -2524 -13534
rect -2454 -12758 -2396 -12746
rect -2454 -13534 -2442 -12758
rect -2408 -13534 -2396 -12758
rect -2454 -13546 -2396 -13534
rect -2316 -12758 -2258 -12746
rect -2316 -13534 -2304 -12758
rect -2270 -13534 -2258 -12758
rect -2316 -13546 -2258 -13534
rect -2188 -12758 -2130 -12746
rect -2188 -13534 -2176 -12758
rect -2142 -13534 -2130 -12758
rect -2188 -13546 -2130 -13534
rect -2050 -12758 -1992 -12746
rect -2050 -13534 -2038 -12758
rect -2004 -13534 -1992 -12758
rect -2050 -13546 -1992 -13534
rect -1922 -12758 -1864 -12746
rect -1922 -13534 -1910 -12758
rect -1876 -13534 -1864 -12758
rect -1922 -13546 -1864 -13534
rect -1784 -12758 -1726 -12746
rect -1784 -13534 -1772 -12758
rect -1738 -13534 -1726 -12758
rect -1784 -13546 -1726 -13534
rect -1656 -12758 -1598 -12746
rect -1656 -13534 -1644 -12758
rect -1610 -13534 -1598 -12758
rect -1656 -13546 -1598 -13534
rect -1518 -12758 -1460 -12746
rect -1518 -13534 -1506 -12758
rect -1472 -13534 -1460 -12758
rect -1518 -13546 -1460 -13534
rect -1390 -12758 -1332 -12746
rect -1390 -13534 -1378 -12758
rect -1344 -13534 -1332 -12758
rect -1390 -13546 -1332 -13534
rect -1252 -12758 -1194 -12746
rect -1252 -13534 -1240 -12758
rect -1206 -13534 -1194 -12758
rect -1252 -13546 -1194 -13534
rect -1124 -12758 -1066 -12746
rect -1124 -13534 -1112 -12758
rect -1078 -13534 -1066 -12758
rect -1124 -13546 -1066 -13534
rect -986 -12758 -928 -12746
rect -986 -13534 -974 -12758
rect -940 -13534 -928 -12758
rect -986 -13546 -928 -13534
rect -858 -12758 -800 -12746
rect -858 -13534 -846 -12758
rect -812 -13534 -800 -12758
rect -858 -13546 -800 -13534
rect -2848 -13768 -2790 -13756
rect -2848 -14544 -2836 -13768
rect -2802 -14544 -2790 -13768
rect -2848 -14556 -2790 -14544
rect -2720 -13768 -2662 -13756
rect -2720 -14544 -2708 -13768
rect -2674 -14544 -2662 -13768
rect -2720 -14556 -2662 -14544
rect -2582 -13768 -2524 -13756
rect -2582 -14544 -2570 -13768
rect -2536 -14544 -2524 -13768
rect -2582 -14556 -2524 -14544
rect -2454 -13768 -2396 -13756
rect -2454 -14544 -2442 -13768
rect -2408 -14544 -2396 -13768
rect -2454 -14556 -2396 -14544
rect -2316 -13768 -2258 -13756
rect -2316 -14544 -2304 -13768
rect -2270 -14544 -2258 -13768
rect -2316 -14556 -2258 -14544
rect -2188 -13768 -2130 -13756
rect -2188 -14544 -2176 -13768
rect -2142 -14544 -2130 -13768
rect -2188 -14556 -2130 -14544
rect -2050 -13768 -1992 -13756
rect -2050 -14544 -2038 -13768
rect -2004 -14544 -1992 -13768
rect -2050 -14556 -1992 -14544
rect -1922 -13768 -1864 -13756
rect -1922 -14544 -1910 -13768
rect -1876 -14544 -1864 -13768
rect -1922 -14556 -1864 -14544
rect -1784 -13768 -1726 -13756
rect -1784 -14544 -1772 -13768
rect -1738 -14544 -1726 -13768
rect -1784 -14556 -1726 -14544
rect -1656 -13768 -1598 -13756
rect -1656 -14544 -1644 -13768
rect -1610 -14544 -1598 -13768
rect -1656 -14556 -1598 -14544
rect -1518 -13768 -1460 -13756
rect -1518 -14544 -1506 -13768
rect -1472 -14544 -1460 -13768
rect -1518 -14556 -1460 -14544
rect -1390 -13768 -1332 -13756
rect -1390 -14544 -1378 -13768
rect -1344 -14544 -1332 -13768
rect -1390 -14556 -1332 -14544
rect -1252 -13768 -1194 -13756
rect -1252 -14544 -1240 -13768
rect -1206 -14544 -1194 -13768
rect -1252 -14556 -1194 -14544
rect -1124 -13768 -1066 -13756
rect -1124 -14544 -1112 -13768
rect -1078 -14544 -1066 -13768
rect -1124 -14556 -1066 -14544
rect -986 -13768 -928 -13756
rect -986 -14544 -974 -13768
rect -940 -14544 -928 -13768
rect -986 -14556 -928 -14544
rect -858 -13768 -800 -13756
rect -858 -14544 -846 -13768
rect -812 -14544 -800 -13768
rect -858 -14556 -800 -14544
rect -2848 -14778 -2790 -14766
rect -2848 -15554 -2836 -14778
rect -2802 -15554 -2790 -14778
rect -2848 -15566 -2790 -15554
rect -2720 -14778 -2662 -14766
rect -2720 -15554 -2708 -14778
rect -2674 -15554 -2662 -14778
rect -2720 -15566 -2662 -15554
rect -2582 -14778 -2524 -14766
rect -2582 -15554 -2570 -14778
rect -2536 -15554 -2524 -14778
rect -2582 -15566 -2524 -15554
rect -2454 -14778 -2396 -14766
rect -2454 -15554 -2442 -14778
rect -2408 -15554 -2396 -14778
rect -2454 -15566 -2396 -15554
rect -2316 -14778 -2258 -14766
rect -2316 -15554 -2304 -14778
rect -2270 -15554 -2258 -14778
rect -2316 -15566 -2258 -15554
rect -2188 -14778 -2130 -14766
rect -2188 -15554 -2176 -14778
rect -2142 -15554 -2130 -14778
rect -2188 -15566 -2130 -15554
rect -2050 -14778 -1992 -14766
rect -2050 -15554 -2038 -14778
rect -2004 -15554 -1992 -14778
rect -2050 -15566 -1992 -15554
rect -1922 -14778 -1864 -14766
rect -1922 -15554 -1910 -14778
rect -1876 -15554 -1864 -14778
rect -1922 -15566 -1864 -15554
rect -1784 -14778 -1726 -14766
rect -1784 -15554 -1772 -14778
rect -1738 -15554 -1726 -14778
rect -1784 -15566 -1726 -15554
rect -1656 -14778 -1598 -14766
rect -1656 -15554 -1644 -14778
rect -1610 -15554 -1598 -14778
rect -1656 -15566 -1598 -15554
rect -1518 -14778 -1460 -14766
rect -1518 -15554 -1506 -14778
rect -1472 -15554 -1460 -14778
rect -1518 -15566 -1460 -15554
rect -1390 -14778 -1332 -14766
rect -1390 -15554 -1378 -14778
rect -1344 -15554 -1332 -14778
rect -1390 -15566 -1332 -15554
rect -1252 -14778 -1194 -14766
rect -1252 -15554 -1240 -14778
rect -1206 -15554 -1194 -14778
rect -1252 -15566 -1194 -15554
rect -1124 -14778 -1066 -14766
rect -1124 -15554 -1112 -14778
rect -1078 -15554 -1066 -14778
rect -1124 -15566 -1066 -15554
rect -986 -14778 -928 -14766
rect -986 -15554 -974 -14778
rect -940 -15554 -928 -14778
rect -986 -15566 -928 -15554
rect -858 -14778 -800 -14766
rect -858 -15554 -846 -14778
rect -812 -15554 -800 -14778
rect -858 -15566 -800 -15554
<< ndiffc >>
rect -6584 -4814 -6550 -4238
rect -6456 -4814 -6422 -4238
rect -6344 -4814 -6310 -4238
rect -6216 -4814 -6182 -4238
rect -6104 -4814 -6070 -4238
rect -5976 -4814 -5942 -4238
rect -5864 -4814 -5830 -4238
rect -5736 -4814 -5702 -4238
rect -5624 -4814 -5590 -4238
rect -5496 -4814 -5462 -4238
rect -5384 -4814 -5350 -4238
rect -5256 -4814 -5222 -4238
rect -5144 -4814 -5110 -4238
rect -5016 -4814 -4982 -4238
rect -4904 -4814 -4870 -4238
rect -4776 -4814 -4742 -4238
rect -4664 -4814 -4630 -4238
rect -4536 -4814 -4502 -4238
rect -4424 -4814 -4390 -4238
rect -4296 -4814 -4262 -4238
rect -4184 -4814 -4150 -4238
rect -4056 -4814 -4022 -4238
rect -3944 -4814 -3910 -4238
rect -3816 -4814 -3782 -4238
rect -3704 -4814 -3670 -4238
rect -3576 -4814 -3542 -4238
rect -3464 -4814 -3430 -4238
rect -3336 -4814 -3302 -4238
rect -3224 -4814 -3190 -4238
rect -3096 -4814 -3062 -4238
rect -2984 -4814 -2950 -4238
rect -2856 -4814 -2822 -4238
rect -2744 -4814 -2710 -4238
rect -2616 -4814 -2582 -4238
rect -2504 -4814 -2470 -4238
rect -2376 -4814 -2342 -4238
rect -2264 -4814 -2230 -4238
rect -2136 -4814 -2102 -4238
rect -2024 -4814 -1990 -4238
rect -1896 -4814 -1862 -4238
rect -1784 -4814 -1750 -4238
rect -1656 -4814 -1622 -4238
rect -1544 -4814 -1510 -4238
rect -1416 -4814 -1382 -4238
rect -1304 -4814 -1270 -4238
rect -1176 -4814 -1142 -4238
rect -1064 -4814 -1030 -4238
rect -936 -4814 -902 -4238
rect -824 -4814 -790 -4238
rect -696 -4814 -662 -4238
rect -584 -4814 -550 -4238
rect -456 -4814 -422 -4238
rect -344 -4814 -310 -4238
rect -216 -4814 -182 -4238
rect -104 -4814 -70 -4238
rect 24 -4814 58 -4238
rect 136 -4814 170 -4238
rect 264 -4814 298 -4238
rect 376 -4814 410 -4238
rect 504 -4814 538 -4238
rect 616 -4814 650 -4238
rect 744 -4814 778 -4238
rect 856 -4814 890 -4238
rect 984 -4814 1018 -4238
rect 1096 -4814 1130 -4238
rect 1224 -4814 1258 -4238
rect 1336 -4814 1370 -4238
rect 1464 -4814 1498 -4238
rect 1576 -4814 1610 -4238
rect 1704 -4814 1738 -4238
rect 1816 -4814 1850 -4238
rect 1944 -4814 1978 -4238
rect 2056 -4814 2090 -4238
rect 2184 -4814 2218 -4238
rect 2296 -4814 2330 -4238
rect 2424 -4814 2458 -4238
rect 2536 -4814 2570 -4238
rect 2664 -4814 2698 -4238
rect 2776 -4814 2810 -4238
rect 2904 -4814 2938 -4238
rect -6584 -5622 -6550 -5046
rect -6456 -5622 -6422 -5046
rect -6344 -5622 -6310 -5046
rect -6216 -5622 -6182 -5046
rect -6104 -5622 -6070 -5046
rect -5976 -5622 -5942 -5046
rect -5864 -5622 -5830 -5046
rect -5736 -5622 -5702 -5046
rect -5624 -5622 -5590 -5046
rect -5496 -5622 -5462 -5046
rect -5384 -5622 -5350 -5046
rect -5256 -5622 -5222 -5046
rect -5144 -5622 -5110 -5046
rect -5016 -5622 -4982 -5046
rect -4904 -5622 -4870 -5046
rect -4776 -5622 -4742 -5046
rect -4664 -5622 -4630 -5046
rect -4536 -5622 -4502 -5046
rect -4424 -5622 -4390 -5046
rect -4296 -5622 -4262 -5046
rect -4184 -5622 -4150 -5046
rect -4056 -5622 -4022 -5046
rect -3944 -5622 -3910 -5046
rect -3816 -5622 -3782 -5046
rect -3704 -5622 -3670 -5046
rect -3576 -5622 -3542 -5046
rect -3464 -5622 -3430 -5046
rect -3336 -5622 -3302 -5046
rect -3224 -5622 -3190 -5046
rect -3096 -5622 -3062 -5046
rect -2984 -5622 -2950 -5046
rect -2856 -5622 -2822 -5046
rect -2744 -5622 -2710 -5046
rect -2616 -5622 -2582 -5046
rect -2504 -5622 -2470 -5046
rect -2376 -5622 -2342 -5046
rect -2264 -5622 -2230 -5046
rect -2136 -5622 -2102 -5046
rect -2024 -5622 -1990 -5046
rect -1896 -5622 -1862 -5046
rect -1784 -5622 -1750 -5046
rect -1656 -5622 -1622 -5046
rect -1544 -5622 -1510 -5046
rect -1416 -5622 -1382 -5046
rect -1304 -5622 -1270 -5046
rect -1176 -5622 -1142 -5046
rect -1064 -5622 -1030 -5046
rect -936 -5622 -902 -5046
rect -824 -5622 -790 -5046
rect -696 -5622 -662 -5046
rect -584 -5622 -550 -5046
rect -456 -5622 -422 -5046
rect -344 -5622 -310 -5046
rect -216 -5622 -182 -5046
rect -104 -5622 -70 -5046
rect 24 -5622 58 -5046
rect 136 -5622 170 -5046
rect 264 -5622 298 -5046
rect 376 -5622 410 -5046
rect 504 -5622 538 -5046
rect 616 -5622 650 -5046
rect 744 -5622 778 -5046
rect 856 -5622 890 -5046
rect 984 -5622 1018 -5046
rect 1096 -5622 1130 -5046
rect 1224 -5622 1258 -5046
rect 1336 -5622 1370 -5046
rect 1464 -5622 1498 -5046
rect 1576 -5622 1610 -5046
rect 1704 -5622 1738 -5046
rect 1816 -5622 1850 -5046
rect 1944 -5622 1978 -5046
rect 2056 -5622 2090 -5046
rect 2184 -5622 2218 -5046
rect 2296 -5622 2330 -5046
rect 2424 -5622 2458 -5046
rect 2536 -5622 2570 -5046
rect 2664 -5622 2698 -5046
rect 2776 -5622 2810 -5046
rect 2904 -5622 2938 -5046
rect -2264 -17526 -2230 -16950
rect -2136 -17526 -2102 -16950
rect -2024 -17526 -1990 -16950
rect -1896 -17526 -1862 -16950
rect -1784 -17526 -1750 -16950
rect -1656 -17526 -1622 -16950
rect -1544 -17526 -1510 -16950
rect -1416 -17526 -1382 -16950
rect -2264 -18334 -2230 -17758
rect -2136 -18334 -2102 -17758
rect -2024 -18334 -1990 -17758
rect -1896 -18334 -1862 -17758
rect -1784 -18334 -1750 -17758
rect -1656 -18334 -1622 -17758
rect -1544 -18334 -1510 -17758
rect -1416 -18334 -1382 -17758
<< pdiffc >>
rect -15888 -9088 -15854 -8312
rect -15430 -9088 -15396 -8312
rect -15300 -9088 -15266 -8312
rect -14842 -9088 -14808 -8312
rect -14712 -9088 -14678 -8312
rect -14254 -9088 -14220 -8312
rect -14124 -9088 -14090 -8312
rect -13666 -9088 -13632 -8312
rect -13536 -9088 -13502 -8312
rect -13078 -9088 -13044 -8312
rect -12948 -9088 -12914 -8312
rect -12490 -9088 -12456 -8312
rect -12360 -9088 -12326 -8312
rect -11902 -9088 -11868 -8312
rect -11772 -9088 -11738 -8312
rect -11314 -9088 -11280 -8312
rect -11184 -9088 -11150 -8312
rect -10726 -9088 -10692 -8312
rect -10596 -9088 -10562 -8312
rect -10138 -9088 -10104 -8312
rect -10008 -9088 -9974 -8312
rect -9550 -9088 -9516 -8312
rect -9420 -9088 -9386 -8312
rect -8962 -9088 -8928 -8312
rect -8832 -9088 -8798 -8312
rect -8374 -9088 -8340 -8312
rect -8244 -9088 -8210 -8312
rect -7786 -9088 -7752 -8312
rect -7656 -9088 -7622 -8312
rect -7198 -9088 -7164 -8312
rect -7068 -9088 -7034 -8312
rect -6610 -9088 -6576 -8312
rect -6480 -9088 -6446 -8312
rect -6022 -9088 -5988 -8312
rect -5892 -9088 -5858 -8312
rect -5434 -9088 -5400 -8312
rect -5304 -9088 -5270 -8312
rect -4846 -9088 -4812 -8312
rect -4716 -9088 -4682 -8312
rect -4258 -9088 -4224 -8312
rect -4128 -9088 -4094 -8312
rect -3670 -9088 -3636 -8312
rect -3540 -9088 -3506 -8312
rect -3082 -9088 -3048 -8312
rect -2952 -9088 -2918 -8312
rect -2494 -9088 -2460 -8312
rect -2364 -9088 -2330 -8312
rect -1906 -9088 -1872 -8312
rect -1776 -9088 -1742 -8312
rect -1318 -9088 -1284 -8312
rect -1188 -9088 -1154 -8312
rect -730 -9088 -696 -8312
rect -600 -9088 -566 -8312
rect -142 -9088 -108 -8312
rect -12 -9088 22 -8312
rect 446 -9088 480 -8312
rect 576 -9088 610 -8312
rect 1034 -9088 1068 -8312
rect 1164 -9088 1198 -8312
rect 1622 -9088 1656 -8312
rect 1752 -9088 1786 -8312
rect 2210 -9088 2244 -8312
rect 2340 -9088 2374 -8312
rect 2798 -9088 2832 -8312
rect 2928 -9088 2962 -8312
rect 3386 -9088 3420 -8312
rect 3516 -9088 3550 -8312
rect 3974 -9088 4008 -8312
rect 4104 -9088 4138 -8312
rect 4562 -9088 4596 -8312
rect 4692 -9088 4726 -8312
rect 5150 -9088 5184 -8312
rect 5280 -9088 5314 -8312
rect 5738 -9088 5772 -8312
rect 5868 -9088 5902 -8312
rect 6326 -9088 6360 -8312
rect 6456 -9088 6490 -8312
rect 6914 -9088 6948 -8312
rect 7044 -9088 7078 -8312
rect 7502 -9088 7536 -8312
rect 7632 -9088 7666 -8312
rect 8090 -9088 8124 -8312
rect 8220 -9088 8254 -8312
rect 8678 -9088 8712 -8312
rect 8808 -9088 8842 -8312
rect 9266 -9088 9300 -8312
rect 9396 -9088 9430 -8312
rect 9854 -9088 9888 -8312
rect 9984 -9088 10018 -8312
rect 10442 -9088 10476 -8312
rect 10572 -9088 10606 -8312
rect 11030 -9088 11064 -8312
rect 11160 -9088 11194 -8312
rect 11618 -9088 11652 -8312
rect 11748 -9088 11782 -8312
rect 12206 -9088 12240 -8312
rect -15888 -10088 -15854 -9312
rect -15430 -10088 -15396 -9312
rect -15300 -10088 -15266 -9312
rect -14842 -10088 -14808 -9312
rect -14712 -10088 -14678 -9312
rect -14254 -10088 -14220 -9312
rect -14124 -10088 -14090 -9312
rect -13666 -10088 -13632 -9312
rect -13536 -10088 -13502 -9312
rect -13078 -10088 -13044 -9312
rect -12948 -10088 -12914 -9312
rect -12490 -10088 -12456 -9312
rect -12360 -10088 -12326 -9312
rect -11902 -10088 -11868 -9312
rect -11772 -10088 -11738 -9312
rect -11314 -10088 -11280 -9312
rect -11184 -10088 -11150 -9312
rect -10726 -10088 -10692 -9312
rect -10596 -10088 -10562 -9312
rect -10138 -10088 -10104 -9312
rect -10008 -10088 -9974 -9312
rect -9550 -10088 -9516 -9312
rect -9420 -10088 -9386 -9312
rect -8962 -10088 -8928 -9312
rect -8832 -10088 -8798 -9312
rect -8374 -10088 -8340 -9312
rect -8244 -10088 -8210 -9312
rect -7786 -10088 -7752 -9312
rect -7656 -10088 -7622 -9312
rect -7198 -10088 -7164 -9312
rect -7068 -10088 -7034 -9312
rect -6610 -10088 -6576 -9312
rect -6480 -10088 -6446 -9312
rect -6022 -10088 -5988 -9312
rect -5892 -10088 -5858 -9312
rect -5434 -10088 -5400 -9312
rect -5304 -10088 -5270 -9312
rect -4846 -10088 -4812 -9312
rect -4716 -10088 -4682 -9312
rect -4258 -10088 -4224 -9312
rect -4128 -10088 -4094 -9312
rect -3670 -10088 -3636 -9312
rect -3540 -10088 -3506 -9312
rect -3082 -10088 -3048 -9312
rect -2952 -10088 -2918 -9312
rect -2494 -10088 -2460 -9312
rect -2364 -10088 -2330 -9312
rect -1906 -10088 -1872 -9312
rect -1776 -10088 -1742 -9312
rect -1318 -10088 -1284 -9312
rect -1188 -10088 -1154 -9312
rect -730 -10088 -696 -9312
rect -600 -10088 -566 -9312
rect -142 -10088 -108 -9312
rect -12 -10088 22 -9312
rect 446 -10088 480 -9312
rect 576 -10088 610 -9312
rect 1034 -10088 1068 -9312
rect 1164 -10088 1198 -9312
rect 1622 -10088 1656 -9312
rect 1752 -10088 1786 -9312
rect 2210 -10088 2244 -9312
rect 2340 -10088 2374 -9312
rect 2798 -10088 2832 -9312
rect 2928 -10088 2962 -9312
rect 3386 -10088 3420 -9312
rect 3516 -10088 3550 -9312
rect 3974 -10088 4008 -9312
rect 4104 -10088 4138 -9312
rect 4562 -10088 4596 -9312
rect 4692 -10088 4726 -9312
rect 5150 -10088 5184 -9312
rect 5280 -10088 5314 -9312
rect 5738 -10088 5772 -9312
rect 5868 -10088 5902 -9312
rect 6326 -10088 6360 -9312
rect 6456 -10088 6490 -9312
rect 6914 -10088 6948 -9312
rect 7044 -10088 7078 -9312
rect 7502 -10088 7536 -9312
rect 7632 -10088 7666 -9312
rect 8090 -10088 8124 -9312
rect 8220 -10088 8254 -9312
rect 8678 -10088 8712 -9312
rect 8808 -10088 8842 -9312
rect 9266 -10088 9300 -9312
rect 9396 -10088 9430 -9312
rect 9854 -10088 9888 -9312
rect 9984 -10088 10018 -9312
rect 10442 -10088 10476 -9312
rect 10572 -10088 10606 -9312
rect 11030 -10088 11064 -9312
rect 11160 -10088 11194 -9312
rect 11618 -10088 11652 -9312
rect 11748 -10088 11782 -9312
rect 12206 -10088 12240 -9312
rect -15888 -11088 -15854 -10312
rect -15430 -11088 -15396 -10312
rect -15300 -11088 -15266 -10312
rect -14842 -11088 -14808 -10312
rect -14712 -11088 -14678 -10312
rect -14254 -11088 -14220 -10312
rect -14124 -11088 -14090 -10312
rect -13666 -11088 -13632 -10312
rect -13536 -11088 -13502 -10312
rect -13078 -11088 -13044 -10312
rect -12948 -11088 -12914 -10312
rect -12490 -11088 -12456 -10312
rect -12360 -11088 -12326 -10312
rect -11902 -11088 -11868 -10312
rect -11772 -11088 -11738 -10312
rect -11314 -11088 -11280 -10312
rect -11184 -11088 -11150 -10312
rect -10726 -11088 -10692 -10312
rect -10596 -11088 -10562 -10312
rect -10138 -11088 -10104 -10312
rect -10008 -11088 -9974 -10312
rect -9550 -11088 -9516 -10312
rect -9420 -11088 -9386 -10312
rect -8962 -11088 -8928 -10312
rect -8832 -11088 -8798 -10312
rect -8374 -11088 -8340 -10312
rect -8244 -11088 -8210 -10312
rect -7786 -11088 -7752 -10312
rect -7656 -11088 -7622 -10312
rect -7198 -11088 -7164 -10312
rect -7068 -11088 -7034 -10312
rect -6610 -11088 -6576 -10312
rect -6480 -11088 -6446 -10312
rect -6022 -11088 -5988 -10312
rect -5892 -11088 -5858 -10312
rect -5434 -11088 -5400 -10312
rect -5304 -11088 -5270 -10312
rect -4846 -11088 -4812 -10312
rect -4716 -11088 -4682 -10312
rect -4258 -11088 -4224 -10312
rect -4128 -11088 -4094 -10312
rect -3670 -11088 -3636 -10312
rect -3540 -11088 -3506 -10312
rect -3082 -11088 -3048 -10312
rect -2952 -11088 -2918 -10312
rect -2494 -11088 -2460 -10312
rect -2364 -11088 -2330 -10312
rect -1906 -11088 -1872 -10312
rect -1776 -11088 -1742 -10312
rect -1318 -11088 -1284 -10312
rect -1188 -11088 -1154 -10312
rect -730 -11088 -696 -10312
rect -600 -11088 -566 -10312
rect -142 -11088 -108 -10312
rect -12 -11088 22 -10312
rect 446 -11088 480 -10312
rect 576 -11088 610 -10312
rect 1034 -11088 1068 -10312
rect 1164 -11088 1198 -10312
rect 1622 -11088 1656 -10312
rect 1752 -11088 1786 -10312
rect 2210 -11088 2244 -10312
rect 2340 -11088 2374 -10312
rect 2798 -11088 2832 -10312
rect 2928 -11088 2962 -10312
rect 3386 -11088 3420 -10312
rect 3516 -11088 3550 -10312
rect 3974 -11088 4008 -10312
rect 4104 -11088 4138 -10312
rect 4562 -11088 4596 -10312
rect 4692 -11088 4726 -10312
rect 5150 -11088 5184 -10312
rect 5280 -11088 5314 -10312
rect 5738 -11088 5772 -10312
rect 5868 -11088 5902 -10312
rect 6326 -11088 6360 -10312
rect 6456 -11088 6490 -10312
rect 6914 -11088 6948 -10312
rect 7044 -11088 7078 -10312
rect 7502 -11088 7536 -10312
rect 7632 -11088 7666 -10312
rect 8090 -11088 8124 -10312
rect 8220 -11088 8254 -10312
rect 8678 -11088 8712 -10312
rect 8808 -11088 8842 -10312
rect 9266 -11088 9300 -10312
rect 9396 -11088 9430 -10312
rect 9854 -11088 9888 -10312
rect 9984 -11088 10018 -10312
rect 10442 -11088 10476 -10312
rect 10572 -11088 10606 -10312
rect 11030 -11088 11064 -10312
rect 11160 -11088 11194 -10312
rect 11618 -11088 11652 -10312
rect 11748 -11088 11782 -10312
rect 12206 -11088 12240 -10312
rect -2836 -13534 -2802 -12758
rect -2708 -13534 -2674 -12758
rect -2570 -13534 -2536 -12758
rect -2442 -13534 -2408 -12758
rect -2304 -13534 -2270 -12758
rect -2176 -13534 -2142 -12758
rect -2038 -13534 -2004 -12758
rect -1910 -13534 -1876 -12758
rect -1772 -13534 -1738 -12758
rect -1644 -13534 -1610 -12758
rect -1506 -13534 -1472 -12758
rect -1378 -13534 -1344 -12758
rect -1240 -13534 -1206 -12758
rect -1112 -13534 -1078 -12758
rect -974 -13534 -940 -12758
rect -846 -13534 -812 -12758
rect -2836 -14544 -2802 -13768
rect -2708 -14544 -2674 -13768
rect -2570 -14544 -2536 -13768
rect -2442 -14544 -2408 -13768
rect -2304 -14544 -2270 -13768
rect -2176 -14544 -2142 -13768
rect -2038 -14544 -2004 -13768
rect -1910 -14544 -1876 -13768
rect -1772 -14544 -1738 -13768
rect -1644 -14544 -1610 -13768
rect -1506 -14544 -1472 -13768
rect -1378 -14544 -1344 -13768
rect -1240 -14544 -1206 -13768
rect -1112 -14544 -1078 -13768
rect -974 -14544 -940 -13768
rect -846 -14544 -812 -13768
rect -2836 -15554 -2802 -14778
rect -2708 -15554 -2674 -14778
rect -2570 -15554 -2536 -14778
rect -2442 -15554 -2408 -14778
rect -2304 -15554 -2270 -14778
rect -2176 -15554 -2142 -14778
rect -2038 -15554 -2004 -14778
rect -1910 -15554 -1876 -14778
rect -1772 -15554 -1738 -14778
rect -1644 -15554 -1610 -14778
rect -1506 -15554 -1472 -14778
rect -1378 -15554 -1344 -14778
rect -1240 -15554 -1206 -14778
rect -1112 -15554 -1078 -14778
rect -974 -15554 -940 -14778
rect -846 -15554 -812 -14778
<< psubdiff >>
rect 4237 -14883 4333 -14849
rect 4471 -14883 4567 -14849
rect 4237 -14945 4271 -14883
rect 4533 -14945 4567 -14883
rect 4237 -16039 4271 -15977
rect 4533 -16039 4567 -15977
rect 4237 -16073 4333 -16039
rect 4471 -16073 4567 -16039
<< nsubdiff >>
rect -3222 -12276 -3188 -12242
rect -460 -12276 -426 -12242
rect -3222 -16072 -3188 -16038
rect -460 -16072 -426 -16038
<< psubdiffcont >>
rect -6842 -3746 3196 -3712
rect -6930 -6060 -6896 -3780
rect 3250 -6060 3284 -3778
rect -6896 -6148 3250 -6114
rect 4333 -14883 4471 -14849
rect 4237 -15977 4271 -14945
rect 4533 -15977 4567 -14945
rect 4333 -16073 4471 -16039
rect -2464 -16468 -1254 -16434
rect -2610 -18816 -2576 -16468
rect -1070 -18816 -1036 -16468
rect -2452 -18850 -1242 -18816
<< nsubdiffcont >>
rect -16074 -7902 12448 -7868
rect -16234 -11478 -16200 -7930
rect 12552 -11444 12586 -7896
rect -16116 -11532 12498 -11498
rect -3188 -12276 -460 -12242
rect -3222 -16038 -3188 -12276
rect -460 -16038 -426 -12276
rect -3188 -16072 -460 -16038
<< poly >>
rect -6538 -4056 -6468 -4046
rect -6538 -4188 -6522 -4056
rect -6484 -4188 -6468 -4056
rect -6538 -4226 -6468 -4188
rect -6298 -4056 -6228 -4046
rect -6298 -4188 -6282 -4056
rect -6244 -4188 -6228 -4056
rect -6298 -4226 -6228 -4188
rect -6058 -4056 -5988 -4046
rect -6058 -4188 -6042 -4056
rect -6004 -4188 -5988 -4056
rect -6058 -4226 -5988 -4188
rect -5818 -4056 -5748 -4046
rect -5818 -4188 -5802 -4056
rect -5764 -4188 -5748 -4056
rect -5818 -4226 -5748 -4188
rect -5578 -4056 -5508 -4046
rect -5578 -4188 -5562 -4056
rect -5524 -4188 -5508 -4056
rect -5578 -4226 -5508 -4188
rect -5338 -4056 -5268 -4046
rect -5338 -4188 -5322 -4056
rect -5284 -4188 -5268 -4056
rect -5338 -4226 -5268 -4188
rect -5098 -4056 -5028 -4046
rect -5098 -4188 -5082 -4056
rect -5044 -4188 -5028 -4056
rect -5098 -4226 -5028 -4188
rect -4858 -4056 -4788 -4046
rect -4858 -4188 -4842 -4056
rect -4804 -4188 -4788 -4056
rect -4858 -4226 -4788 -4188
rect -4618 -4056 -4548 -4046
rect -4618 -4188 -4602 -4056
rect -4564 -4188 -4548 -4056
rect -4618 -4226 -4548 -4188
rect -4378 -4056 -4308 -4046
rect -4378 -4188 -4362 -4056
rect -4324 -4188 -4308 -4056
rect -4378 -4226 -4308 -4188
rect -4138 -4056 -4068 -4046
rect -4138 -4188 -4122 -4056
rect -4084 -4188 -4068 -4056
rect -4138 -4226 -4068 -4188
rect -3898 -4056 -3828 -4046
rect -3898 -4188 -3882 -4056
rect -3844 -4188 -3828 -4056
rect -3898 -4226 -3828 -4188
rect -3658 -4056 -3588 -4046
rect -3658 -4188 -3642 -4056
rect -3604 -4188 -3588 -4056
rect -3658 -4226 -3588 -4188
rect -3418 -4056 -3348 -4046
rect -3418 -4188 -3402 -4056
rect -3364 -4188 -3348 -4056
rect -3418 -4226 -3348 -4188
rect -3178 -4056 -3108 -4046
rect -3178 -4188 -3162 -4056
rect -3124 -4188 -3108 -4056
rect -3178 -4226 -3108 -4188
rect -2938 -4056 -2868 -4046
rect -2938 -4188 -2922 -4056
rect -2884 -4188 -2868 -4056
rect -2938 -4226 -2868 -4188
rect -2698 -4056 -2628 -4046
rect -2698 -4188 -2682 -4056
rect -2644 -4188 -2628 -4056
rect -2698 -4226 -2628 -4188
rect -2458 -4056 -2388 -4046
rect -2458 -4188 -2442 -4056
rect -2404 -4188 -2388 -4056
rect -2458 -4226 -2388 -4188
rect -2218 -4056 -2148 -4046
rect -2218 -4188 -2202 -4056
rect -2164 -4188 -2148 -4056
rect -2218 -4226 -2148 -4188
rect -1978 -4056 -1908 -4046
rect -1978 -4188 -1962 -4056
rect -1924 -4188 -1908 -4056
rect -1978 -4226 -1908 -4188
rect -1738 -4056 -1668 -4046
rect -1738 -4188 -1722 -4056
rect -1684 -4188 -1668 -4056
rect -1738 -4226 -1668 -4188
rect -1498 -4056 -1428 -4046
rect -1498 -4188 -1482 -4056
rect -1444 -4188 -1428 -4056
rect -1498 -4226 -1428 -4188
rect -1258 -4056 -1188 -4046
rect -1258 -4188 -1242 -4056
rect -1204 -4188 -1188 -4056
rect -1258 -4226 -1188 -4188
rect -1018 -4056 -948 -4046
rect -1018 -4188 -1002 -4056
rect -964 -4188 -948 -4056
rect -1018 -4226 -948 -4188
rect -778 -4056 -708 -4046
rect -778 -4188 -762 -4056
rect -724 -4188 -708 -4056
rect -778 -4226 -708 -4188
rect -538 -4056 -468 -4046
rect -538 -4188 -522 -4056
rect -484 -4188 -468 -4056
rect -538 -4226 -468 -4188
rect -298 -4056 -228 -4046
rect -298 -4188 -282 -4056
rect -244 -4188 -228 -4056
rect -298 -4226 -228 -4188
rect -58 -4056 12 -4046
rect -58 -4188 -42 -4056
rect -4 -4188 12 -4056
rect -58 -4226 12 -4188
rect 182 -4056 252 -4046
rect 182 -4188 198 -4056
rect 236 -4188 252 -4056
rect 182 -4226 252 -4188
rect 422 -4056 492 -4046
rect 422 -4188 438 -4056
rect 476 -4188 492 -4056
rect 422 -4226 492 -4188
rect 662 -4056 732 -4046
rect 662 -4188 678 -4056
rect 716 -4188 732 -4056
rect 662 -4226 732 -4188
rect 902 -4056 972 -4046
rect 902 -4188 918 -4056
rect 956 -4188 972 -4056
rect 902 -4226 972 -4188
rect 1142 -4056 1212 -4046
rect 1142 -4188 1158 -4056
rect 1196 -4188 1212 -4056
rect 1142 -4226 1212 -4188
rect 1382 -4056 1452 -4046
rect 1382 -4188 1398 -4056
rect 1436 -4188 1452 -4056
rect 1382 -4226 1452 -4188
rect 1622 -4056 1692 -4046
rect 1622 -4188 1638 -4056
rect 1676 -4188 1692 -4056
rect 1622 -4226 1692 -4188
rect 1862 -4056 1932 -4046
rect 1862 -4188 1878 -4056
rect 1916 -4188 1932 -4056
rect 1862 -4226 1932 -4188
rect 2102 -4056 2172 -4046
rect 2102 -4188 2118 -4056
rect 2156 -4188 2172 -4056
rect 2102 -4226 2172 -4188
rect 2342 -4056 2412 -4046
rect 2342 -4188 2358 -4056
rect 2396 -4188 2412 -4056
rect 2342 -4226 2412 -4188
rect 2582 -4056 2652 -4046
rect 2582 -4188 2598 -4056
rect 2636 -4188 2652 -4056
rect 2582 -4226 2652 -4188
rect 2822 -4056 2892 -4046
rect 2822 -4188 2838 -4056
rect 2876 -4188 2892 -4056
rect 2822 -4226 2892 -4188
rect -6538 -4864 -6468 -4826
rect -6538 -4996 -6522 -4864
rect -6484 -4996 -6468 -4864
rect -6538 -5034 -6468 -4996
rect -6298 -4864 -6228 -4826
rect -6298 -4996 -6282 -4864
rect -6244 -4996 -6228 -4864
rect -6298 -5034 -6228 -4996
rect -6058 -4864 -5988 -4826
rect -6058 -4996 -6042 -4864
rect -6004 -4996 -5988 -4864
rect -6058 -5034 -5988 -4996
rect -5818 -4864 -5748 -4826
rect -5818 -4996 -5802 -4864
rect -5764 -4996 -5748 -4864
rect -5818 -5034 -5748 -4996
rect -5578 -4864 -5508 -4826
rect -5578 -4996 -5562 -4864
rect -5524 -4996 -5508 -4864
rect -5578 -5034 -5508 -4996
rect -5338 -4864 -5268 -4826
rect -5338 -4996 -5322 -4864
rect -5284 -4996 -5268 -4864
rect -5338 -5034 -5268 -4996
rect -5098 -4864 -5028 -4826
rect -5098 -4996 -5082 -4864
rect -5044 -4996 -5028 -4864
rect -5098 -5034 -5028 -4996
rect -4858 -4864 -4788 -4826
rect -4858 -4996 -4842 -4864
rect -4804 -4996 -4788 -4864
rect -4858 -5034 -4788 -4996
rect -4618 -4864 -4548 -4826
rect -4618 -4996 -4602 -4864
rect -4564 -4996 -4548 -4864
rect -4618 -5034 -4548 -4996
rect -4378 -4864 -4308 -4826
rect -4378 -4996 -4362 -4864
rect -4324 -4996 -4308 -4864
rect -4378 -5034 -4308 -4996
rect -4138 -4864 -4068 -4826
rect -4138 -4996 -4122 -4864
rect -4084 -4996 -4068 -4864
rect -4138 -5034 -4068 -4996
rect -3898 -4864 -3828 -4826
rect -3898 -4996 -3882 -4864
rect -3844 -4996 -3828 -4864
rect -3898 -5034 -3828 -4996
rect -3658 -4864 -3588 -4826
rect -3658 -4996 -3642 -4864
rect -3604 -4996 -3588 -4864
rect -3658 -5034 -3588 -4996
rect -3418 -4864 -3348 -4826
rect -3418 -4996 -3402 -4864
rect -3364 -4996 -3348 -4864
rect -3418 -5034 -3348 -4996
rect -3178 -4864 -3108 -4826
rect -3178 -4996 -3162 -4864
rect -3124 -4996 -3108 -4864
rect -3178 -5034 -3108 -4996
rect -2938 -4864 -2868 -4826
rect -2938 -4996 -2922 -4864
rect -2884 -4996 -2868 -4864
rect -2938 -5034 -2868 -4996
rect -2698 -4864 -2628 -4826
rect -2698 -4996 -2682 -4864
rect -2644 -4996 -2628 -4864
rect -2698 -5034 -2628 -4996
rect -2458 -4864 -2388 -4826
rect -2458 -4996 -2442 -4864
rect -2404 -4996 -2388 -4864
rect -2458 -5034 -2388 -4996
rect -2218 -4864 -2148 -4826
rect -2218 -4996 -2202 -4864
rect -2164 -4996 -2148 -4864
rect -2218 -5034 -2148 -4996
rect -1978 -4864 -1908 -4826
rect -1978 -4996 -1962 -4864
rect -1924 -4996 -1908 -4864
rect -1978 -5034 -1908 -4996
rect -1738 -4864 -1668 -4826
rect -1738 -4996 -1722 -4864
rect -1684 -4996 -1668 -4864
rect -1738 -5034 -1668 -4996
rect -1498 -4864 -1428 -4826
rect -1498 -4996 -1482 -4864
rect -1444 -4996 -1428 -4864
rect -1498 -5034 -1428 -4996
rect -1258 -4864 -1188 -4826
rect -1258 -4996 -1242 -4864
rect -1204 -4996 -1188 -4864
rect -1258 -5034 -1188 -4996
rect -1018 -4864 -948 -4826
rect -1018 -4996 -1002 -4864
rect -964 -4996 -948 -4864
rect -1018 -5034 -948 -4996
rect -778 -4864 -708 -4826
rect -778 -4996 -762 -4864
rect -724 -4996 -708 -4864
rect -778 -5034 -708 -4996
rect -538 -4864 -468 -4826
rect -538 -4996 -522 -4864
rect -484 -4996 -468 -4864
rect -538 -5034 -468 -4996
rect -298 -4864 -228 -4826
rect -298 -4996 -282 -4864
rect -244 -4996 -228 -4864
rect -298 -5034 -228 -4996
rect -58 -4864 12 -4826
rect -58 -4996 -42 -4864
rect -4 -4996 12 -4864
rect -58 -5034 12 -4996
rect 182 -4864 252 -4826
rect 182 -4996 198 -4864
rect 236 -4996 252 -4864
rect 182 -5034 252 -4996
rect 422 -4864 492 -4826
rect 422 -4996 438 -4864
rect 476 -4996 492 -4864
rect 422 -5034 492 -4996
rect 662 -4864 732 -4826
rect 662 -4996 678 -4864
rect 716 -4996 732 -4864
rect 662 -5034 732 -4996
rect 902 -4864 972 -4826
rect 902 -4996 918 -4864
rect 956 -4996 972 -4864
rect 902 -5034 972 -4996
rect 1142 -4864 1212 -4826
rect 1142 -4996 1158 -4864
rect 1196 -4996 1212 -4864
rect 1142 -5034 1212 -4996
rect 1382 -4864 1452 -4826
rect 1382 -4996 1398 -4864
rect 1436 -4996 1452 -4864
rect 1382 -5034 1452 -4996
rect 1622 -4864 1692 -4826
rect 1622 -4996 1638 -4864
rect 1676 -4996 1692 -4864
rect 1622 -5034 1692 -4996
rect 1862 -4864 1932 -4826
rect 1862 -4996 1878 -4864
rect 1916 -4996 1932 -4864
rect 1862 -5034 1932 -4996
rect 2102 -4864 2172 -4826
rect 2102 -4996 2118 -4864
rect 2156 -4996 2172 -4864
rect 2102 -5034 2172 -4996
rect 2342 -4864 2412 -4826
rect 2342 -4996 2358 -4864
rect 2396 -4996 2412 -4864
rect 2342 -5034 2412 -4996
rect 2582 -4864 2652 -4826
rect 2582 -4996 2598 -4864
rect 2636 -4996 2652 -4864
rect 2582 -5034 2652 -4996
rect 2822 -4864 2892 -4826
rect 2822 -4996 2838 -4864
rect 2876 -4996 2892 -4864
rect 2822 -5034 2892 -4996
rect -6538 -5672 -6468 -5634
rect -6538 -5804 -6522 -5672
rect -6484 -5804 -6468 -5672
rect -6538 -5814 -6468 -5804
rect -6298 -5672 -6228 -5634
rect -6298 -5804 -6282 -5672
rect -6244 -5804 -6228 -5672
rect -6298 -5814 -6228 -5804
rect -6058 -5672 -5988 -5634
rect -6058 -5804 -6042 -5672
rect -6004 -5804 -5988 -5672
rect -6058 -5814 -5988 -5804
rect -5818 -5672 -5748 -5634
rect -5818 -5804 -5802 -5672
rect -5764 -5804 -5748 -5672
rect -5818 -5814 -5748 -5804
rect -5578 -5672 -5508 -5634
rect -5578 -5804 -5562 -5672
rect -5524 -5804 -5508 -5672
rect -5578 -5814 -5508 -5804
rect -5338 -5672 -5268 -5634
rect -5338 -5804 -5322 -5672
rect -5284 -5804 -5268 -5672
rect -5338 -5814 -5268 -5804
rect -5098 -5672 -5028 -5634
rect -5098 -5804 -5082 -5672
rect -5044 -5804 -5028 -5672
rect -5098 -5814 -5028 -5804
rect -4858 -5672 -4788 -5634
rect -4858 -5804 -4842 -5672
rect -4804 -5804 -4788 -5672
rect -4858 -5814 -4788 -5804
rect -4618 -5672 -4548 -5634
rect -4618 -5804 -4602 -5672
rect -4564 -5804 -4548 -5672
rect -4618 -5814 -4548 -5804
rect -4378 -5672 -4308 -5634
rect -4378 -5804 -4362 -5672
rect -4324 -5804 -4308 -5672
rect -4378 -5814 -4308 -5804
rect -4138 -5672 -4068 -5634
rect -4138 -5804 -4122 -5672
rect -4084 -5804 -4068 -5672
rect -4138 -5814 -4068 -5804
rect -3898 -5672 -3828 -5634
rect -3898 -5804 -3882 -5672
rect -3844 -5804 -3828 -5672
rect -3898 -5814 -3828 -5804
rect -3658 -5672 -3588 -5634
rect -3658 -5804 -3642 -5672
rect -3604 -5804 -3588 -5672
rect -3658 -5814 -3588 -5804
rect -3418 -5672 -3348 -5634
rect -3418 -5804 -3402 -5672
rect -3364 -5804 -3348 -5672
rect -3418 -5814 -3348 -5804
rect -3178 -5672 -3108 -5634
rect -3178 -5804 -3162 -5672
rect -3124 -5804 -3108 -5672
rect -3178 -5814 -3108 -5804
rect -2938 -5672 -2868 -5634
rect -2938 -5804 -2922 -5672
rect -2884 -5804 -2868 -5672
rect -2938 -5814 -2868 -5804
rect -2698 -5672 -2628 -5634
rect -2698 -5804 -2682 -5672
rect -2644 -5804 -2628 -5672
rect -2698 -5814 -2628 -5804
rect -2458 -5672 -2388 -5634
rect -2458 -5804 -2442 -5672
rect -2404 -5804 -2388 -5672
rect -2458 -5814 -2388 -5804
rect -2218 -5672 -2148 -5634
rect -2218 -5804 -2202 -5672
rect -2164 -5804 -2148 -5672
rect -2218 -5814 -2148 -5804
rect -1978 -5672 -1908 -5634
rect -1978 -5804 -1962 -5672
rect -1924 -5804 -1908 -5672
rect -1978 -5814 -1908 -5804
rect -1738 -5672 -1668 -5634
rect -1738 -5804 -1722 -5672
rect -1684 -5804 -1668 -5672
rect -1738 -5814 -1668 -5804
rect -1498 -5672 -1428 -5634
rect -1498 -5804 -1482 -5672
rect -1444 -5804 -1428 -5672
rect -1498 -5814 -1428 -5804
rect -1258 -5672 -1188 -5634
rect -1258 -5804 -1242 -5672
rect -1204 -5804 -1188 -5672
rect -1258 -5814 -1188 -5804
rect -1018 -5672 -948 -5634
rect -1018 -5804 -1002 -5672
rect -964 -5804 -948 -5672
rect -1018 -5814 -948 -5804
rect -778 -5672 -708 -5634
rect -778 -5804 -762 -5672
rect -724 -5804 -708 -5672
rect -778 -5814 -708 -5804
rect -538 -5672 -468 -5634
rect -538 -5804 -522 -5672
rect -484 -5804 -468 -5672
rect -538 -5814 -468 -5804
rect -298 -5672 -228 -5634
rect -298 -5804 -282 -5672
rect -244 -5804 -228 -5672
rect -298 -5814 -228 -5804
rect -58 -5672 12 -5634
rect -58 -5804 -42 -5672
rect -4 -5804 12 -5672
rect -58 -5814 12 -5804
rect 182 -5672 252 -5634
rect 182 -5804 198 -5672
rect 236 -5804 252 -5672
rect 182 -5814 252 -5804
rect 422 -5672 492 -5634
rect 422 -5804 438 -5672
rect 476 -5804 492 -5672
rect 422 -5814 492 -5804
rect 662 -5672 732 -5634
rect 662 -5804 678 -5672
rect 716 -5804 732 -5672
rect 662 -5814 732 -5804
rect 902 -5672 972 -5634
rect 902 -5804 918 -5672
rect 956 -5804 972 -5672
rect 902 -5814 972 -5804
rect 1142 -5672 1212 -5634
rect 1142 -5804 1158 -5672
rect 1196 -5804 1212 -5672
rect 1142 -5814 1212 -5804
rect 1382 -5672 1452 -5634
rect 1382 -5804 1398 -5672
rect 1436 -5804 1452 -5672
rect 1382 -5814 1452 -5804
rect 1622 -5672 1692 -5634
rect 1622 -5804 1638 -5672
rect 1676 -5804 1692 -5672
rect 1622 -5814 1692 -5804
rect 1862 -5672 1932 -5634
rect 1862 -5804 1878 -5672
rect 1916 -5804 1932 -5672
rect 1862 -5814 1932 -5804
rect 2102 -5672 2172 -5634
rect 2102 -5804 2118 -5672
rect 2156 -5804 2172 -5672
rect 2102 -5814 2172 -5804
rect 2342 -5672 2412 -5634
rect 2342 -5804 2358 -5672
rect 2396 -5804 2412 -5672
rect 2342 -5814 2412 -5804
rect 2582 -5672 2652 -5634
rect 2582 -5804 2598 -5672
rect 2636 -5804 2652 -5672
rect 2582 -5814 2652 -5804
rect 2822 -5672 2892 -5634
rect 2822 -5804 2838 -5672
rect 2876 -5804 2892 -5672
rect 2822 -5814 2892 -5804
rect -15842 -8219 -15442 -8203
rect -15842 -8253 -15826 -8219
rect -15458 -8253 -15442 -8219
rect -15842 -8300 -15442 -8253
rect -15254 -8219 -14854 -8203
rect -15254 -8253 -15238 -8219
rect -14870 -8253 -14854 -8219
rect -15254 -8300 -14854 -8253
rect -14666 -8219 -14266 -8203
rect -14666 -8253 -14650 -8219
rect -14282 -8253 -14266 -8219
rect -14666 -8300 -14266 -8253
rect -14078 -8219 -13678 -8203
rect -14078 -8253 -14062 -8219
rect -13694 -8253 -13678 -8219
rect -14078 -8300 -13678 -8253
rect -13490 -8219 -13090 -8203
rect -13490 -8253 -13474 -8219
rect -13106 -8253 -13090 -8219
rect -13490 -8300 -13090 -8253
rect -12902 -8219 -12502 -8203
rect -12902 -8253 -12886 -8219
rect -12518 -8253 -12502 -8219
rect -12902 -8300 -12502 -8253
rect -12314 -8219 -11914 -8203
rect -12314 -8253 -12298 -8219
rect -11930 -8253 -11914 -8219
rect -12314 -8300 -11914 -8253
rect -11726 -8219 -11326 -8203
rect -11726 -8253 -11710 -8219
rect -11342 -8253 -11326 -8219
rect -11726 -8300 -11326 -8253
rect -11138 -8219 -10738 -8203
rect -11138 -8253 -11122 -8219
rect -10754 -8253 -10738 -8219
rect -11138 -8300 -10738 -8253
rect -10550 -8219 -10150 -8203
rect -10550 -8253 -10534 -8219
rect -10166 -8253 -10150 -8219
rect -10550 -8300 -10150 -8253
rect -9962 -8219 -9562 -8203
rect -9962 -8253 -9946 -8219
rect -9578 -8253 -9562 -8219
rect -9962 -8300 -9562 -8253
rect -9374 -8219 -8974 -8203
rect -9374 -8253 -9358 -8219
rect -8990 -8253 -8974 -8219
rect -9374 -8300 -8974 -8253
rect -8786 -8219 -8386 -8203
rect -8786 -8253 -8770 -8219
rect -8402 -8253 -8386 -8219
rect -8786 -8300 -8386 -8253
rect -8198 -8219 -7798 -8203
rect -8198 -8253 -8182 -8219
rect -7814 -8253 -7798 -8219
rect -8198 -8300 -7798 -8253
rect -7610 -8219 -7210 -8203
rect -7610 -8253 -7594 -8219
rect -7226 -8253 -7210 -8219
rect -7610 -8300 -7210 -8253
rect -7022 -8219 -6622 -8203
rect -7022 -8253 -7006 -8219
rect -6638 -8253 -6622 -8219
rect -7022 -8300 -6622 -8253
rect -6434 -8219 -6034 -8203
rect -6434 -8253 -6418 -8219
rect -6050 -8253 -6034 -8219
rect -6434 -8300 -6034 -8253
rect -5846 -8219 -5446 -8203
rect -5846 -8253 -5830 -8219
rect -5462 -8253 -5446 -8219
rect -5846 -8300 -5446 -8253
rect -5258 -8219 -4858 -8203
rect -5258 -8253 -5242 -8219
rect -4874 -8253 -4858 -8219
rect -5258 -8300 -4858 -8253
rect -4670 -8219 -4270 -8203
rect -4670 -8253 -4654 -8219
rect -4286 -8253 -4270 -8219
rect -4670 -8300 -4270 -8253
rect -4082 -8219 -3682 -8203
rect -4082 -8253 -4066 -8219
rect -3698 -8253 -3682 -8219
rect -4082 -8300 -3682 -8253
rect -3494 -8219 -3094 -8203
rect -3494 -8253 -3478 -8219
rect -3110 -8253 -3094 -8219
rect -3494 -8300 -3094 -8253
rect -2906 -8219 -2506 -8203
rect -2906 -8253 -2890 -8219
rect -2522 -8253 -2506 -8219
rect -2906 -8300 -2506 -8253
rect -2318 -8219 -1918 -8203
rect -2318 -8253 -2302 -8219
rect -1934 -8253 -1918 -8219
rect -2318 -8300 -1918 -8253
rect -1730 -8219 -1330 -8203
rect -1730 -8253 -1714 -8219
rect -1346 -8253 -1330 -8219
rect -1730 -8300 -1330 -8253
rect -1142 -8219 -742 -8203
rect -1142 -8253 -1126 -8219
rect -758 -8253 -742 -8219
rect -1142 -8300 -742 -8253
rect -554 -8219 -154 -8203
rect -554 -8253 -538 -8219
rect -170 -8253 -154 -8219
rect -554 -8300 -154 -8253
rect 34 -8219 434 -8203
rect 34 -8253 50 -8219
rect 418 -8253 434 -8219
rect 34 -8300 434 -8253
rect 622 -8219 1022 -8203
rect 622 -8253 638 -8219
rect 1006 -8253 1022 -8219
rect 622 -8300 1022 -8253
rect 1210 -8219 1610 -8203
rect 1210 -8253 1226 -8219
rect 1594 -8253 1610 -8219
rect 1210 -8300 1610 -8253
rect 1798 -8219 2198 -8203
rect 1798 -8253 1814 -8219
rect 2182 -8253 2198 -8219
rect 1798 -8300 2198 -8253
rect 2386 -8219 2786 -8203
rect 2386 -8253 2402 -8219
rect 2770 -8253 2786 -8219
rect 2386 -8300 2786 -8253
rect 2974 -8219 3374 -8203
rect 2974 -8253 2990 -8219
rect 3358 -8253 3374 -8219
rect 2974 -8300 3374 -8253
rect 3562 -8219 3962 -8203
rect 3562 -8253 3578 -8219
rect 3946 -8253 3962 -8219
rect 3562 -8300 3962 -8253
rect 4150 -8219 4550 -8203
rect 4150 -8253 4166 -8219
rect 4534 -8253 4550 -8219
rect 4150 -8300 4550 -8253
rect 4738 -8219 5138 -8203
rect 4738 -8253 4754 -8219
rect 5122 -8253 5138 -8219
rect 4738 -8300 5138 -8253
rect 5326 -8219 5726 -8203
rect 5326 -8253 5342 -8219
rect 5710 -8253 5726 -8219
rect 5326 -8300 5726 -8253
rect 5914 -8219 6314 -8203
rect 5914 -8253 5930 -8219
rect 6298 -8253 6314 -8219
rect 5914 -8300 6314 -8253
rect 6502 -8219 6902 -8203
rect 6502 -8253 6518 -8219
rect 6886 -8253 6902 -8219
rect 6502 -8300 6902 -8253
rect 7090 -8219 7490 -8203
rect 7090 -8253 7106 -8219
rect 7474 -8253 7490 -8219
rect 7090 -8300 7490 -8253
rect 7678 -8219 8078 -8203
rect 7678 -8253 7694 -8219
rect 8062 -8253 8078 -8219
rect 7678 -8300 8078 -8253
rect 8266 -8219 8666 -8203
rect 8266 -8253 8282 -8219
rect 8650 -8253 8666 -8219
rect 8266 -8300 8666 -8253
rect 8854 -8219 9254 -8203
rect 8854 -8253 8870 -8219
rect 9238 -8253 9254 -8219
rect 8854 -8300 9254 -8253
rect 9442 -8219 9842 -8203
rect 9442 -8253 9458 -8219
rect 9826 -8253 9842 -8219
rect 9442 -8300 9842 -8253
rect 10030 -8219 10430 -8203
rect 10030 -8253 10046 -8219
rect 10414 -8253 10430 -8219
rect 10030 -8300 10430 -8253
rect 10618 -8219 11018 -8203
rect 10618 -8253 10634 -8219
rect 11002 -8253 11018 -8219
rect 10618 -8300 11018 -8253
rect 11206 -8219 11606 -8203
rect 11206 -8253 11222 -8219
rect 11590 -8253 11606 -8219
rect 11206 -8300 11606 -8253
rect 11794 -8219 12194 -8203
rect 11794 -8253 11810 -8219
rect 12178 -8253 12194 -8219
rect 11794 -8300 12194 -8253
rect -15842 -9147 -15442 -9100
rect -15842 -9181 -15826 -9147
rect -15458 -9181 -15442 -9147
rect -15842 -9219 -15442 -9181
rect -15842 -9253 -15826 -9219
rect -15458 -9253 -15442 -9219
rect -15842 -9300 -15442 -9253
rect -15254 -9147 -14854 -9100
rect -15254 -9181 -15238 -9147
rect -14870 -9181 -14854 -9147
rect -15254 -9219 -14854 -9181
rect -15254 -9253 -15238 -9219
rect -14870 -9253 -14854 -9219
rect -15254 -9300 -14854 -9253
rect -14666 -9147 -14266 -9100
rect -14666 -9181 -14650 -9147
rect -14282 -9181 -14266 -9147
rect -14666 -9219 -14266 -9181
rect -14666 -9253 -14650 -9219
rect -14282 -9253 -14266 -9219
rect -14666 -9300 -14266 -9253
rect -14078 -9147 -13678 -9100
rect -14078 -9181 -14062 -9147
rect -13694 -9181 -13678 -9147
rect -14078 -9219 -13678 -9181
rect -14078 -9253 -14062 -9219
rect -13694 -9253 -13678 -9219
rect -14078 -9300 -13678 -9253
rect -13490 -9147 -13090 -9100
rect -13490 -9181 -13474 -9147
rect -13106 -9181 -13090 -9147
rect -13490 -9219 -13090 -9181
rect -13490 -9253 -13474 -9219
rect -13106 -9253 -13090 -9219
rect -13490 -9300 -13090 -9253
rect -12902 -9147 -12502 -9100
rect -12902 -9181 -12886 -9147
rect -12518 -9181 -12502 -9147
rect -12902 -9219 -12502 -9181
rect -12902 -9253 -12886 -9219
rect -12518 -9253 -12502 -9219
rect -12902 -9300 -12502 -9253
rect -12314 -9147 -11914 -9100
rect -12314 -9181 -12298 -9147
rect -11930 -9181 -11914 -9147
rect -12314 -9219 -11914 -9181
rect -12314 -9253 -12298 -9219
rect -11930 -9253 -11914 -9219
rect -12314 -9300 -11914 -9253
rect -11726 -9147 -11326 -9100
rect -11726 -9181 -11710 -9147
rect -11342 -9181 -11326 -9147
rect -11726 -9219 -11326 -9181
rect -11726 -9253 -11710 -9219
rect -11342 -9253 -11326 -9219
rect -11726 -9300 -11326 -9253
rect -11138 -9147 -10738 -9100
rect -11138 -9181 -11122 -9147
rect -10754 -9181 -10738 -9147
rect -11138 -9219 -10738 -9181
rect -11138 -9253 -11122 -9219
rect -10754 -9253 -10738 -9219
rect -11138 -9300 -10738 -9253
rect -10550 -9147 -10150 -9100
rect -10550 -9181 -10534 -9147
rect -10166 -9181 -10150 -9147
rect -10550 -9219 -10150 -9181
rect -10550 -9253 -10534 -9219
rect -10166 -9253 -10150 -9219
rect -10550 -9300 -10150 -9253
rect -9962 -9147 -9562 -9100
rect -9962 -9181 -9946 -9147
rect -9578 -9181 -9562 -9147
rect -9962 -9219 -9562 -9181
rect -9962 -9253 -9946 -9219
rect -9578 -9253 -9562 -9219
rect -9962 -9300 -9562 -9253
rect -9374 -9147 -8974 -9100
rect -9374 -9181 -9358 -9147
rect -8990 -9181 -8974 -9147
rect -9374 -9219 -8974 -9181
rect -9374 -9253 -9358 -9219
rect -8990 -9253 -8974 -9219
rect -9374 -9300 -8974 -9253
rect -8786 -9147 -8386 -9100
rect -8786 -9181 -8770 -9147
rect -8402 -9181 -8386 -9147
rect -8786 -9219 -8386 -9181
rect -8786 -9253 -8770 -9219
rect -8402 -9253 -8386 -9219
rect -8786 -9300 -8386 -9253
rect -8198 -9147 -7798 -9100
rect -8198 -9181 -8182 -9147
rect -7814 -9181 -7798 -9147
rect -8198 -9219 -7798 -9181
rect -8198 -9253 -8182 -9219
rect -7814 -9253 -7798 -9219
rect -8198 -9300 -7798 -9253
rect -7610 -9147 -7210 -9100
rect -7610 -9181 -7594 -9147
rect -7226 -9181 -7210 -9147
rect -7610 -9219 -7210 -9181
rect -7610 -9253 -7594 -9219
rect -7226 -9253 -7210 -9219
rect -7610 -9300 -7210 -9253
rect -7022 -9147 -6622 -9100
rect -7022 -9181 -7006 -9147
rect -6638 -9181 -6622 -9147
rect -7022 -9219 -6622 -9181
rect -7022 -9253 -7006 -9219
rect -6638 -9253 -6622 -9219
rect -7022 -9300 -6622 -9253
rect -6434 -9147 -6034 -9100
rect -6434 -9181 -6418 -9147
rect -6050 -9181 -6034 -9147
rect -6434 -9219 -6034 -9181
rect -6434 -9253 -6418 -9219
rect -6050 -9253 -6034 -9219
rect -6434 -9300 -6034 -9253
rect -5846 -9147 -5446 -9100
rect -5846 -9181 -5830 -9147
rect -5462 -9181 -5446 -9147
rect -5846 -9219 -5446 -9181
rect -5846 -9253 -5830 -9219
rect -5462 -9253 -5446 -9219
rect -5846 -9300 -5446 -9253
rect -5258 -9147 -4858 -9100
rect -5258 -9181 -5242 -9147
rect -4874 -9181 -4858 -9147
rect -5258 -9219 -4858 -9181
rect -5258 -9253 -5242 -9219
rect -4874 -9253 -4858 -9219
rect -5258 -9300 -4858 -9253
rect -4670 -9147 -4270 -9100
rect -4670 -9181 -4654 -9147
rect -4286 -9181 -4270 -9147
rect -4670 -9219 -4270 -9181
rect -4670 -9253 -4654 -9219
rect -4286 -9253 -4270 -9219
rect -4670 -9300 -4270 -9253
rect -4082 -9147 -3682 -9100
rect -4082 -9181 -4066 -9147
rect -3698 -9181 -3682 -9147
rect -4082 -9219 -3682 -9181
rect -4082 -9253 -4066 -9219
rect -3698 -9253 -3682 -9219
rect -4082 -9300 -3682 -9253
rect -3494 -9147 -3094 -9100
rect -3494 -9181 -3478 -9147
rect -3110 -9181 -3094 -9147
rect -3494 -9219 -3094 -9181
rect -3494 -9253 -3478 -9219
rect -3110 -9253 -3094 -9219
rect -3494 -9300 -3094 -9253
rect -2906 -9147 -2506 -9100
rect -2906 -9181 -2890 -9147
rect -2522 -9181 -2506 -9147
rect -2906 -9219 -2506 -9181
rect -2906 -9253 -2890 -9219
rect -2522 -9253 -2506 -9219
rect -2906 -9300 -2506 -9253
rect -2318 -9147 -1918 -9100
rect -2318 -9181 -2302 -9147
rect -1934 -9181 -1918 -9147
rect -2318 -9219 -1918 -9181
rect -2318 -9253 -2302 -9219
rect -1934 -9253 -1918 -9219
rect -2318 -9300 -1918 -9253
rect -1730 -9147 -1330 -9100
rect -1730 -9181 -1714 -9147
rect -1346 -9181 -1330 -9147
rect -1730 -9219 -1330 -9181
rect -1730 -9253 -1714 -9219
rect -1346 -9253 -1330 -9219
rect -1730 -9300 -1330 -9253
rect -1142 -9147 -742 -9100
rect -1142 -9181 -1126 -9147
rect -758 -9181 -742 -9147
rect -1142 -9219 -742 -9181
rect -1142 -9253 -1126 -9219
rect -758 -9253 -742 -9219
rect -1142 -9300 -742 -9253
rect -554 -9147 -154 -9100
rect -554 -9181 -538 -9147
rect -170 -9181 -154 -9147
rect -554 -9219 -154 -9181
rect -554 -9253 -538 -9219
rect -170 -9253 -154 -9219
rect -554 -9300 -154 -9253
rect 34 -9147 434 -9100
rect 34 -9181 50 -9147
rect 418 -9181 434 -9147
rect 34 -9219 434 -9181
rect 34 -9253 50 -9219
rect 418 -9253 434 -9219
rect 34 -9300 434 -9253
rect 622 -9147 1022 -9100
rect 622 -9181 638 -9147
rect 1006 -9181 1022 -9147
rect 622 -9219 1022 -9181
rect 622 -9253 638 -9219
rect 1006 -9253 1022 -9219
rect 622 -9300 1022 -9253
rect 1210 -9147 1610 -9100
rect 1210 -9181 1226 -9147
rect 1594 -9181 1610 -9147
rect 1210 -9219 1610 -9181
rect 1210 -9253 1226 -9219
rect 1594 -9253 1610 -9219
rect 1210 -9300 1610 -9253
rect 1798 -9147 2198 -9100
rect 1798 -9181 1814 -9147
rect 2182 -9181 2198 -9147
rect 1798 -9219 2198 -9181
rect 1798 -9253 1814 -9219
rect 2182 -9253 2198 -9219
rect 1798 -9300 2198 -9253
rect 2386 -9147 2786 -9100
rect 2386 -9181 2402 -9147
rect 2770 -9181 2786 -9147
rect 2386 -9219 2786 -9181
rect 2386 -9253 2402 -9219
rect 2770 -9253 2786 -9219
rect 2386 -9300 2786 -9253
rect 2974 -9147 3374 -9100
rect 2974 -9181 2990 -9147
rect 3358 -9181 3374 -9147
rect 2974 -9219 3374 -9181
rect 2974 -9253 2990 -9219
rect 3358 -9253 3374 -9219
rect 2974 -9300 3374 -9253
rect 3562 -9147 3962 -9100
rect 3562 -9181 3578 -9147
rect 3946 -9181 3962 -9147
rect 3562 -9219 3962 -9181
rect 3562 -9253 3578 -9219
rect 3946 -9253 3962 -9219
rect 3562 -9300 3962 -9253
rect 4150 -9147 4550 -9100
rect 4150 -9181 4166 -9147
rect 4534 -9181 4550 -9147
rect 4150 -9219 4550 -9181
rect 4150 -9253 4166 -9219
rect 4534 -9253 4550 -9219
rect 4150 -9300 4550 -9253
rect 4738 -9147 5138 -9100
rect 4738 -9181 4754 -9147
rect 5122 -9181 5138 -9147
rect 4738 -9219 5138 -9181
rect 4738 -9253 4754 -9219
rect 5122 -9253 5138 -9219
rect 4738 -9300 5138 -9253
rect 5326 -9147 5726 -9100
rect 5326 -9181 5342 -9147
rect 5710 -9181 5726 -9147
rect 5326 -9219 5726 -9181
rect 5326 -9253 5342 -9219
rect 5710 -9253 5726 -9219
rect 5326 -9300 5726 -9253
rect 5914 -9147 6314 -9100
rect 5914 -9181 5930 -9147
rect 6298 -9181 6314 -9147
rect 5914 -9219 6314 -9181
rect 5914 -9253 5930 -9219
rect 6298 -9253 6314 -9219
rect 5914 -9300 6314 -9253
rect 6502 -9147 6902 -9100
rect 6502 -9181 6518 -9147
rect 6886 -9181 6902 -9147
rect 6502 -9219 6902 -9181
rect 6502 -9253 6518 -9219
rect 6886 -9253 6902 -9219
rect 6502 -9300 6902 -9253
rect 7090 -9147 7490 -9100
rect 7090 -9181 7106 -9147
rect 7474 -9181 7490 -9147
rect 7090 -9219 7490 -9181
rect 7090 -9253 7106 -9219
rect 7474 -9253 7490 -9219
rect 7090 -9300 7490 -9253
rect 7678 -9147 8078 -9100
rect 7678 -9181 7694 -9147
rect 8062 -9181 8078 -9147
rect 7678 -9219 8078 -9181
rect 7678 -9253 7694 -9219
rect 8062 -9253 8078 -9219
rect 7678 -9300 8078 -9253
rect 8266 -9147 8666 -9100
rect 8266 -9181 8282 -9147
rect 8650 -9181 8666 -9147
rect 8266 -9219 8666 -9181
rect 8266 -9253 8282 -9219
rect 8650 -9253 8666 -9219
rect 8266 -9300 8666 -9253
rect 8854 -9147 9254 -9100
rect 8854 -9181 8870 -9147
rect 9238 -9181 9254 -9147
rect 8854 -9219 9254 -9181
rect 8854 -9253 8870 -9219
rect 9238 -9253 9254 -9219
rect 8854 -9300 9254 -9253
rect 9442 -9147 9842 -9100
rect 9442 -9181 9458 -9147
rect 9826 -9181 9842 -9147
rect 9442 -9219 9842 -9181
rect 9442 -9253 9458 -9219
rect 9826 -9253 9842 -9219
rect 9442 -9300 9842 -9253
rect 10030 -9147 10430 -9100
rect 10030 -9181 10046 -9147
rect 10414 -9181 10430 -9147
rect 10030 -9219 10430 -9181
rect 10030 -9253 10046 -9219
rect 10414 -9253 10430 -9219
rect 10030 -9300 10430 -9253
rect 10618 -9147 11018 -9100
rect 10618 -9181 10634 -9147
rect 11002 -9181 11018 -9147
rect 10618 -9219 11018 -9181
rect 10618 -9253 10634 -9219
rect 11002 -9253 11018 -9219
rect 10618 -9300 11018 -9253
rect 11206 -9147 11606 -9100
rect 11206 -9181 11222 -9147
rect 11590 -9181 11606 -9147
rect 11206 -9219 11606 -9181
rect 11206 -9253 11222 -9219
rect 11590 -9253 11606 -9219
rect 11206 -9300 11606 -9253
rect 11794 -9147 12194 -9100
rect 11794 -9181 11810 -9147
rect 12178 -9181 12194 -9147
rect 11794 -9219 12194 -9181
rect 11794 -9253 11810 -9219
rect 12178 -9253 12194 -9219
rect 11794 -9300 12194 -9253
rect -15842 -10147 -15442 -10100
rect -15842 -10181 -15826 -10147
rect -15458 -10181 -15442 -10147
rect -15842 -10219 -15442 -10181
rect -15842 -10253 -15826 -10219
rect -15458 -10253 -15442 -10219
rect -15842 -10300 -15442 -10253
rect -15254 -10147 -14854 -10100
rect -15254 -10181 -15238 -10147
rect -14870 -10181 -14854 -10147
rect -15254 -10219 -14854 -10181
rect -15254 -10253 -15238 -10219
rect -14870 -10253 -14854 -10219
rect -15254 -10300 -14854 -10253
rect -14666 -10147 -14266 -10100
rect -14666 -10181 -14650 -10147
rect -14282 -10181 -14266 -10147
rect -14666 -10219 -14266 -10181
rect -14666 -10253 -14650 -10219
rect -14282 -10253 -14266 -10219
rect -14666 -10300 -14266 -10253
rect -14078 -10147 -13678 -10100
rect -14078 -10181 -14062 -10147
rect -13694 -10181 -13678 -10147
rect -14078 -10219 -13678 -10181
rect -14078 -10253 -14062 -10219
rect -13694 -10253 -13678 -10219
rect -14078 -10300 -13678 -10253
rect -13490 -10147 -13090 -10100
rect -13490 -10181 -13474 -10147
rect -13106 -10181 -13090 -10147
rect -13490 -10219 -13090 -10181
rect -13490 -10253 -13474 -10219
rect -13106 -10253 -13090 -10219
rect -13490 -10300 -13090 -10253
rect -12902 -10147 -12502 -10100
rect -12902 -10181 -12886 -10147
rect -12518 -10181 -12502 -10147
rect -12902 -10219 -12502 -10181
rect -12902 -10253 -12886 -10219
rect -12518 -10253 -12502 -10219
rect -12902 -10300 -12502 -10253
rect -12314 -10147 -11914 -10100
rect -12314 -10181 -12298 -10147
rect -11930 -10181 -11914 -10147
rect -12314 -10219 -11914 -10181
rect -12314 -10253 -12298 -10219
rect -11930 -10253 -11914 -10219
rect -12314 -10300 -11914 -10253
rect -11726 -10147 -11326 -10100
rect -11726 -10181 -11710 -10147
rect -11342 -10181 -11326 -10147
rect -11726 -10219 -11326 -10181
rect -11726 -10253 -11710 -10219
rect -11342 -10253 -11326 -10219
rect -11726 -10300 -11326 -10253
rect -11138 -10147 -10738 -10100
rect -11138 -10181 -11122 -10147
rect -10754 -10181 -10738 -10147
rect -11138 -10219 -10738 -10181
rect -11138 -10253 -11122 -10219
rect -10754 -10253 -10738 -10219
rect -11138 -10300 -10738 -10253
rect -10550 -10147 -10150 -10100
rect -10550 -10181 -10534 -10147
rect -10166 -10181 -10150 -10147
rect -10550 -10219 -10150 -10181
rect -10550 -10253 -10534 -10219
rect -10166 -10253 -10150 -10219
rect -10550 -10300 -10150 -10253
rect -9962 -10147 -9562 -10100
rect -9962 -10181 -9946 -10147
rect -9578 -10181 -9562 -10147
rect -9962 -10219 -9562 -10181
rect -9962 -10253 -9946 -10219
rect -9578 -10253 -9562 -10219
rect -9962 -10300 -9562 -10253
rect -9374 -10147 -8974 -10100
rect -9374 -10181 -9358 -10147
rect -8990 -10181 -8974 -10147
rect -9374 -10219 -8974 -10181
rect -9374 -10253 -9358 -10219
rect -8990 -10253 -8974 -10219
rect -9374 -10300 -8974 -10253
rect -8786 -10147 -8386 -10100
rect -8786 -10181 -8770 -10147
rect -8402 -10181 -8386 -10147
rect -8786 -10219 -8386 -10181
rect -8786 -10253 -8770 -10219
rect -8402 -10253 -8386 -10219
rect -8786 -10300 -8386 -10253
rect -8198 -10147 -7798 -10100
rect -8198 -10181 -8182 -10147
rect -7814 -10181 -7798 -10147
rect -8198 -10219 -7798 -10181
rect -8198 -10253 -8182 -10219
rect -7814 -10253 -7798 -10219
rect -8198 -10300 -7798 -10253
rect -7610 -10147 -7210 -10100
rect -7610 -10181 -7594 -10147
rect -7226 -10181 -7210 -10147
rect -7610 -10219 -7210 -10181
rect -7610 -10253 -7594 -10219
rect -7226 -10253 -7210 -10219
rect -7610 -10300 -7210 -10253
rect -7022 -10147 -6622 -10100
rect -7022 -10181 -7006 -10147
rect -6638 -10181 -6622 -10147
rect -7022 -10219 -6622 -10181
rect -7022 -10253 -7006 -10219
rect -6638 -10253 -6622 -10219
rect -7022 -10300 -6622 -10253
rect -6434 -10147 -6034 -10100
rect -6434 -10181 -6418 -10147
rect -6050 -10181 -6034 -10147
rect -6434 -10219 -6034 -10181
rect -6434 -10253 -6418 -10219
rect -6050 -10253 -6034 -10219
rect -6434 -10300 -6034 -10253
rect -5846 -10147 -5446 -10100
rect -5846 -10181 -5830 -10147
rect -5462 -10181 -5446 -10147
rect -5846 -10219 -5446 -10181
rect -5846 -10253 -5830 -10219
rect -5462 -10253 -5446 -10219
rect -5846 -10300 -5446 -10253
rect -5258 -10147 -4858 -10100
rect -5258 -10181 -5242 -10147
rect -4874 -10181 -4858 -10147
rect -5258 -10219 -4858 -10181
rect -5258 -10253 -5242 -10219
rect -4874 -10253 -4858 -10219
rect -5258 -10300 -4858 -10253
rect -4670 -10147 -4270 -10100
rect -4670 -10181 -4654 -10147
rect -4286 -10181 -4270 -10147
rect -4670 -10219 -4270 -10181
rect -4670 -10253 -4654 -10219
rect -4286 -10253 -4270 -10219
rect -4670 -10300 -4270 -10253
rect -4082 -10147 -3682 -10100
rect -4082 -10181 -4066 -10147
rect -3698 -10181 -3682 -10147
rect -4082 -10219 -3682 -10181
rect -4082 -10253 -4066 -10219
rect -3698 -10253 -3682 -10219
rect -4082 -10300 -3682 -10253
rect -3494 -10147 -3094 -10100
rect -3494 -10181 -3478 -10147
rect -3110 -10181 -3094 -10147
rect -3494 -10219 -3094 -10181
rect -3494 -10253 -3478 -10219
rect -3110 -10253 -3094 -10219
rect -3494 -10300 -3094 -10253
rect -2906 -10147 -2506 -10100
rect -2906 -10181 -2890 -10147
rect -2522 -10181 -2506 -10147
rect -2906 -10219 -2506 -10181
rect -2906 -10253 -2890 -10219
rect -2522 -10253 -2506 -10219
rect -2906 -10300 -2506 -10253
rect -2318 -10147 -1918 -10100
rect -2318 -10181 -2302 -10147
rect -1934 -10181 -1918 -10147
rect -2318 -10219 -1918 -10181
rect -2318 -10253 -2302 -10219
rect -1934 -10253 -1918 -10219
rect -2318 -10300 -1918 -10253
rect -1730 -10147 -1330 -10100
rect -1730 -10181 -1714 -10147
rect -1346 -10181 -1330 -10147
rect -1730 -10219 -1330 -10181
rect -1730 -10253 -1714 -10219
rect -1346 -10253 -1330 -10219
rect -1730 -10300 -1330 -10253
rect -1142 -10147 -742 -10100
rect -1142 -10181 -1126 -10147
rect -758 -10181 -742 -10147
rect -1142 -10219 -742 -10181
rect -1142 -10253 -1126 -10219
rect -758 -10253 -742 -10219
rect -1142 -10300 -742 -10253
rect -554 -10147 -154 -10100
rect -554 -10181 -538 -10147
rect -170 -10181 -154 -10147
rect -554 -10219 -154 -10181
rect -554 -10253 -538 -10219
rect -170 -10253 -154 -10219
rect -554 -10300 -154 -10253
rect 34 -10147 434 -10100
rect 34 -10181 50 -10147
rect 418 -10181 434 -10147
rect 34 -10219 434 -10181
rect 34 -10253 50 -10219
rect 418 -10253 434 -10219
rect 34 -10300 434 -10253
rect 622 -10147 1022 -10100
rect 622 -10181 638 -10147
rect 1006 -10181 1022 -10147
rect 622 -10219 1022 -10181
rect 622 -10253 638 -10219
rect 1006 -10253 1022 -10219
rect 622 -10300 1022 -10253
rect 1210 -10147 1610 -10100
rect 1210 -10181 1226 -10147
rect 1594 -10181 1610 -10147
rect 1210 -10219 1610 -10181
rect 1210 -10253 1226 -10219
rect 1594 -10253 1610 -10219
rect 1210 -10300 1610 -10253
rect 1798 -10147 2198 -10100
rect 1798 -10181 1814 -10147
rect 2182 -10181 2198 -10147
rect 1798 -10219 2198 -10181
rect 1798 -10253 1814 -10219
rect 2182 -10253 2198 -10219
rect 1798 -10300 2198 -10253
rect 2386 -10147 2786 -10100
rect 2386 -10181 2402 -10147
rect 2770 -10181 2786 -10147
rect 2386 -10219 2786 -10181
rect 2386 -10253 2402 -10219
rect 2770 -10253 2786 -10219
rect 2386 -10300 2786 -10253
rect 2974 -10147 3374 -10100
rect 2974 -10181 2990 -10147
rect 3358 -10181 3374 -10147
rect 2974 -10219 3374 -10181
rect 2974 -10253 2990 -10219
rect 3358 -10253 3374 -10219
rect 2974 -10300 3374 -10253
rect 3562 -10147 3962 -10100
rect 3562 -10181 3578 -10147
rect 3946 -10181 3962 -10147
rect 3562 -10219 3962 -10181
rect 3562 -10253 3578 -10219
rect 3946 -10253 3962 -10219
rect 3562 -10300 3962 -10253
rect 4150 -10147 4550 -10100
rect 4150 -10181 4166 -10147
rect 4534 -10181 4550 -10147
rect 4150 -10219 4550 -10181
rect 4150 -10253 4166 -10219
rect 4534 -10253 4550 -10219
rect 4150 -10300 4550 -10253
rect 4738 -10147 5138 -10100
rect 4738 -10181 4754 -10147
rect 5122 -10181 5138 -10147
rect 4738 -10219 5138 -10181
rect 4738 -10253 4754 -10219
rect 5122 -10253 5138 -10219
rect 4738 -10300 5138 -10253
rect 5326 -10147 5726 -10100
rect 5326 -10181 5342 -10147
rect 5710 -10181 5726 -10147
rect 5326 -10219 5726 -10181
rect 5326 -10253 5342 -10219
rect 5710 -10253 5726 -10219
rect 5326 -10300 5726 -10253
rect 5914 -10147 6314 -10100
rect 5914 -10181 5930 -10147
rect 6298 -10181 6314 -10147
rect 5914 -10219 6314 -10181
rect 5914 -10253 5930 -10219
rect 6298 -10253 6314 -10219
rect 5914 -10300 6314 -10253
rect 6502 -10147 6902 -10100
rect 6502 -10181 6518 -10147
rect 6886 -10181 6902 -10147
rect 6502 -10219 6902 -10181
rect 6502 -10253 6518 -10219
rect 6886 -10253 6902 -10219
rect 6502 -10300 6902 -10253
rect 7090 -10147 7490 -10100
rect 7090 -10181 7106 -10147
rect 7474 -10181 7490 -10147
rect 7090 -10219 7490 -10181
rect 7090 -10253 7106 -10219
rect 7474 -10253 7490 -10219
rect 7090 -10300 7490 -10253
rect 7678 -10147 8078 -10100
rect 7678 -10181 7694 -10147
rect 8062 -10181 8078 -10147
rect 7678 -10219 8078 -10181
rect 7678 -10253 7694 -10219
rect 8062 -10253 8078 -10219
rect 7678 -10300 8078 -10253
rect 8266 -10147 8666 -10100
rect 8266 -10181 8282 -10147
rect 8650 -10181 8666 -10147
rect 8266 -10219 8666 -10181
rect 8266 -10253 8282 -10219
rect 8650 -10253 8666 -10219
rect 8266 -10300 8666 -10253
rect 8854 -10147 9254 -10100
rect 8854 -10181 8870 -10147
rect 9238 -10181 9254 -10147
rect 8854 -10219 9254 -10181
rect 8854 -10253 8870 -10219
rect 9238 -10253 9254 -10219
rect 8854 -10300 9254 -10253
rect 9442 -10147 9842 -10100
rect 9442 -10181 9458 -10147
rect 9826 -10181 9842 -10147
rect 9442 -10219 9842 -10181
rect 9442 -10253 9458 -10219
rect 9826 -10253 9842 -10219
rect 9442 -10300 9842 -10253
rect 10030 -10147 10430 -10100
rect 10030 -10181 10046 -10147
rect 10414 -10181 10430 -10147
rect 10030 -10219 10430 -10181
rect 10030 -10253 10046 -10219
rect 10414 -10253 10430 -10219
rect 10030 -10300 10430 -10253
rect 10618 -10147 11018 -10100
rect 10618 -10181 10634 -10147
rect 11002 -10181 11018 -10147
rect 10618 -10219 11018 -10181
rect 10618 -10253 10634 -10219
rect 11002 -10253 11018 -10219
rect 10618 -10300 11018 -10253
rect 11206 -10147 11606 -10100
rect 11206 -10181 11222 -10147
rect 11590 -10181 11606 -10147
rect 11206 -10219 11606 -10181
rect 11206 -10253 11222 -10219
rect 11590 -10253 11606 -10219
rect 11206 -10300 11606 -10253
rect 11794 -10147 12194 -10100
rect 11794 -10181 11810 -10147
rect 12178 -10181 12194 -10147
rect 11794 -10219 12194 -10181
rect 11794 -10253 11810 -10219
rect 12178 -10253 12194 -10219
rect 11794 -10300 12194 -10253
rect -15842 -11147 -15442 -11100
rect -15842 -11181 -15826 -11147
rect -15458 -11181 -15442 -11147
rect -15842 -11197 -15442 -11181
rect -15254 -11147 -14854 -11100
rect -15254 -11181 -15238 -11147
rect -14870 -11181 -14854 -11147
rect -15254 -11197 -14854 -11181
rect -14666 -11147 -14266 -11100
rect -14666 -11181 -14650 -11147
rect -14282 -11181 -14266 -11147
rect -14666 -11197 -14266 -11181
rect -14078 -11147 -13678 -11100
rect -14078 -11181 -14062 -11147
rect -13694 -11181 -13678 -11147
rect -14078 -11197 -13678 -11181
rect -13490 -11147 -13090 -11100
rect -13490 -11181 -13474 -11147
rect -13106 -11181 -13090 -11147
rect -13490 -11197 -13090 -11181
rect -12902 -11147 -12502 -11100
rect -12902 -11181 -12886 -11147
rect -12518 -11181 -12502 -11147
rect -12902 -11197 -12502 -11181
rect -12314 -11147 -11914 -11100
rect -12314 -11181 -12298 -11147
rect -11930 -11181 -11914 -11147
rect -12314 -11197 -11914 -11181
rect -11726 -11147 -11326 -11100
rect -11726 -11181 -11710 -11147
rect -11342 -11181 -11326 -11147
rect -11726 -11197 -11326 -11181
rect -11138 -11147 -10738 -11100
rect -11138 -11181 -11122 -11147
rect -10754 -11181 -10738 -11147
rect -11138 -11197 -10738 -11181
rect -10550 -11147 -10150 -11100
rect -10550 -11181 -10534 -11147
rect -10166 -11181 -10150 -11147
rect -10550 -11197 -10150 -11181
rect -9962 -11147 -9562 -11100
rect -9962 -11181 -9946 -11147
rect -9578 -11181 -9562 -11147
rect -9962 -11197 -9562 -11181
rect -9374 -11147 -8974 -11100
rect -9374 -11181 -9358 -11147
rect -8990 -11181 -8974 -11147
rect -9374 -11197 -8974 -11181
rect -8786 -11147 -8386 -11100
rect -8786 -11181 -8770 -11147
rect -8402 -11181 -8386 -11147
rect -8786 -11197 -8386 -11181
rect -8198 -11147 -7798 -11100
rect -8198 -11181 -8182 -11147
rect -7814 -11181 -7798 -11147
rect -8198 -11197 -7798 -11181
rect -7610 -11147 -7210 -11100
rect -7610 -11181 -7594 -11147
rect -7226 -11181 -7210 -11147
rect -7610 -11197 -7210 -11181
rect -7022 -11147 -6622 -11100
rect -7022 -11181 -7006 -11147
rect -6638 -11181 -6622 -11147
rect -7022 -11197 -6622 -11181
rect -6434 -11147 -6034 -11100
rect -6434 -11181 -6418 -11147
rect -6050 -11181 -6034 -11147
rect -6434 -11197 -6034 -11181
rect -5846 -11147 -5446 -11100
rect -5846 -11181 -5830 -11147
rect -5462 -11181 -5446 -11147
rect -5846 -11197 -5446 -11181
rect -5258 -11147 -4858 -11100
rect -5258 -11181 -5242 -11147
rect -4874 -11181 -4858 -11147
rect -5258 -11197 -4858 -11181
rect -4670 -11147 -4270 -11100
rect -4670 -11181 -4654 -11147
rect -4286 -11181 -4270 -11147
rect -4670 -11197 -4270 -11181
rect -4082 -11147 -3682 -11100
rect -4082 -11181 -4066 -11147
rect -3698 -11181 -3682 -11147
rect -4082 -11197 -3682 -11181
rect -3494 -11147 -3094 -11100
rect -3494 -11181 -3478 -11147
rect -3110 -11181 -3094 -11147
rect -3494 -11197 -3094 -11181
rect -2906 -11147 -2506 -11100
rect -2906 -11181 -2890 -11147
rect -2522 -11181 -2506 -11147
rect -2906 -11197 -2506 -11181
rect -2318 -11147 -1918 -11100
rect -2318 -11181 -2302 -11147
rect -1934 -11181 -1918 -11147
rect -2318 -11197 -1918 -11181
rect -1730 -11147 -1330 -11100
rect -1730 -11181 -1714 -11147
rect -1346 -11181 -1330 -11147
rect -1730 -11197 -1330 -11181
rect -1142 -11147 -742 -11100
rect -1142 -11181 -1126 -11147
rect -758 -11181 -742 -11147
rect -1142 -11197 -742 -11181
rect -554 -11147 -154 -11100
rect -554 -11181 -538 -11147
rect -170 -11181 -154 -11147
rect -554 -11197 -154 -11181
rect 34 -11147 434 -11100
rect 34 -11181 50 -11147
rect 418 -11181 434 -11147
rect 34 -11197 434 -11181
rect 622 -11147 1022 -11100
rect 622 -11181 638 -11147
rect 1006 -11181 1022 -11147
rect 622 -11197 1022 -11181
rect 1210 -11147 1610 -11100
rect 1210 -11181 1226 -11147
rect 1594 -11181 1610 -11147
rect 1210 -11197 1610 -11181
rect 1798 -11147 2198 -11100
rect 1798 -11181 1814 -11147
rect 2182 -11181 2198 -11147
rect 1798 -11197 2198 -11181
rect 2386 -11147 2786 -11100
rect 2386 -11181 2402 -11147
rect 2770 -11181 2786 -11147
rect 2386 -11197 2786 -11181
rect 2974 -11147 3374 -11100
rect 2974 -11181 2990 -11147
rect 3358 -11181 3374 -11147
rect 2974 -11197 3374 -11181
rect 3562 -11147 3962 -11100
rect 3562 -11181 3578 -11147
rect 3946 -11181 3962 -11147
rect 3562 -11197 3962 -11181
rect 4150 -11147 4550 -11100
rect 4150 -11181 4166 -11147
rect 4534 -11181 4550 -11147
rect 4150 -11197 4550 -11181
rect 4738 -11147 5138 -11100
rect 4738 -11181 4754 -11147
rect 5122 -11181 5138 -11147
rect 4738 -11197 5138 -11181
rect 5326 -11147 5726 -11100
rect 5326 -11181 5342 -11147
rect 5710 -11181 5726 -11147
rect 5326 -11197 5726 -11181
rect 5914 -11147 6314 -11100
rect 5914 -11181 5930 -11147
rect 6298 -11181 6314 -11147
rect 5914 -11197 6314 -11181
rect 6502 -11147 6902 -11100
rect 6502 -11181 6518 -11147
rect 6886 -11181 6902 -11147
rect 6502 -11197 6902 -11181
rect 7090 -11147 7490 -11100
rect 7090 -11181 7106 -11147
rect 7474 -11181 7490 -11147
rect 7090 -11197 7490 -11181
rect 7678 -11147 8078 -11100
rect 7678 -11181 7694 -11147
rect 8062 -11181 8078 -11147
rect 7678 -11197 8078 -11181
rect 8266 -11147 8666 -11100
rect 8266 -11181 8282 -11147
rect 8650 -11181 8666 -11147
rect 8266 -11197 8666 -11181
rect 8854 -11147 9254 -11100
rect 8854 -11181 8870 -11147
rect 9238 -11181 9254 -11147
rect 8854 -11197 9254 -11181
rect 9442 -11147 9842 -11100
rect 9442 -11181 9458 -11147
rect 9826 -11181 9842 -11147
rect 9442 -11197 9842 -11181
rect 10030 -11147 10430 -11100
rect 10030 -11181 10046 -11147
rect 10414 -11181 10430 -11147
rect 10030 -11197 10430 -11181
rect 10618 -11147 11018 -11100
rect 10618 -11181 10634 -11147
rect 11002 -11181 11018 -11147
rect 10618 -11197 11018 -11181
rect 11206 -11147 11606 -11100
rect 11206 -11181 11222 -11147
rect 11590 -11181 11606 -11147
rect 11206 -11197 11606 -11181
rect 11794 -11147 12194 -11100
rect 11794 -11181 11810 -11147
rect 12178 -11181 12194 -11147
rect 11794 -11197 12194 -11181
rect -2790 -12576 -2720 -12570
rect -2790 -12708 -2774 -12576
rect -2736 -12708 -2720 -12576
rect -2790 -12746 -2720 -12708
rect -2524 -12576 -2454 -12570
rect -2524 -12708 -2508 -12576
rect -2470 -12708 -2454 -12576
rect -2524 -12746 -2454 -12708
rect -2258 -12576 -2188 -12570
rect -2258 -12708 -2242 -12576
rect -2204 -12708 -2188 -12576
rect -2258 -12746 -2188 -12708
rect -1992 -12576 -1922 -12570
rect -1992 -12708 -1976 -12576
rect -1938 -12708 -1922 -12576
rect -1992 -12746 -1922 -12708
rect -1726 -12576 -1656 -12570
rect -1726 -12708 -1710 -12576
rect -1672 -12708 -1656 -12576
rect -1726 -12746 -1656 -12708
rect -1460 -12576 -1390 -12570
rect -1460 -12708 -1444 -12576
rect -1406 -12708 -1390 -12576
rect -1460 -12746 -1390 -12708
rect -1194 -12576 -1124 -12570
rect -1194 -12708 -1178 -12576
rect -1140 -12708 -1124 -12576
rect -1194 -12746 -1124 -12708
rect -928 -12576 -858 -12570
rect -928 -12708 -912 -12576
rect -874 -12708 -858 -12576
rect -928 -12746 -858 -12708
rect -2790 -13586 -2720 -13546
rect -2790 -13718 -2774 -13586
rect -2736 -13718 -2720 -13586
rect -2790 -13756 -2720 -13718
rect -2524 -13586 -2454 -13546
rect -2524 -13718 -2508 -13586
rect -2470 -13718 -2454 -13586
rect -2524 -13756 -2454 -13718
rect -2258 -13586 -2188 -13546
rect -2258 -13718 -2242 -13586
rect -2204 -13718 -2188 -13586
rect -2258 -13756 -2188 -13718
rect -1992 -13586 -1922 -13546
rect -1992 -13718 -1976 -13586
rect -1938 -13718 -1922 -13586
rect -1992 -13756 -1922 -13718
rect -1726 -13586 -1656 -13546
rect -1726 -13718 -1710 -13586
rect -1672 -13718 -1656 -13586
rect -1726 -13756 -1656 -13718
rect -1460 -13586 -1390 -13546
rect -1460 -13718 -1444 -13586
rect -1406 -13718 -1390 -13586
rect -1460 -13756 -1390 -13718
rect -1194 -13586 -1124 -13546
rect -1194 -13718 -1178 -13586
rect -1140 -13718 -1124 -13586
rect -1194 -13756 -1124 -13718
rect -928 -13586 -858 -13546
rect -928 -13718 -912 -13586
rect -874 -13718 -858 -13586
rect -928 -13756 -858 -13718
rect -2790 -14596 -2720 -14556
rect -2790 -14728 -2774 -14596
rect -2736 -14728 -2720 -14596
rect -2790 -14766 -2720 -14728
rect -2524 -14596 -2454 -14556
rect -2524 -14728 -2508 -14596
rect -2470 -14728 -2454 -14596
rect -2524 -14766 -2454 -14728
rect -2258 -14596 -2188 -14556
rect -2258 -14728 -2242 -14596
rect -2204 -14728 -2188 -14596
rect -2258 -14766 -2188 -14728
rect -1992 -14596 -1922 -14556
rect -1992 -14728 -1976 -14596
rect -1938 -14728 -1922 -14596
rect -1992 -14766 -1922 -14728
rect -1726 -14596 -1656 -14556
rect -1726 -14728 -1710 -14596
rect -1672 -14728 -1656 -14596
rect -1726 -14766 -1656 -14728
rect -1460 -14596 -1390 -14556
rect -1460 -14728 -1444 -14596
rect -1406 -14728 -1390 -14596
rect -1460 -14766 -1390 -14728
rect -1194 -14596 -1124 -14556
rect -1194 -14728 -1178 -14596
rect -1140 -14728 -1124 -14596
rect -1194 -14766 -1124 -14728
rect -928 -14596 -858 -14556
rect -928 -14728 -912 -14596
rect -874 -14728 -858 -14596
rect -928 -14766 -858 -14728
rect -2790 -15606 -2720 -15566
rect -2790 -15738 -2774 -15606
rect -2736 -15738 -2720 -15606
rect -2790 -15748 -2720 -15738
rect -2524 -15606 -2454 -15566
rect -2524 -15738 -2508 -15606
rect -2470 -15738 -2454 -15606
rect -2524 -15748 -2454 -15738
rect -2258 -15606 -2188 -15566
rect -2258 -15738 -2242 -15606
rect -2204 -15738 -2188 -15606
rect -2258 -15748 -2188 -15738
rect -1992 -15606 -1922 -15566
rect -1992 -15738 -1976 -15606
rect -1938 -15738 -1922 -15606
rect -1992 -15748 -1922 -15738
rect -1726 -15606 -1656 -15566
rect -1726 -15738 -1710 -15606
rect -1672 -15738 -1656 -15606
rect -1726 -15748 -1656 -15738
rect -1460 -15606 -1390 -15566
rect -1460 -15738 -1444 -15606
rect -1406 -15738 -1390 -15606
rect -1460 -15748 -1390 -15738
rect -1194 -15606 -1124 -15566
rect -1194 -15738 -1178 -15606
rect -1140 -15738 -1124 -15606
rect -1194 -15748 -1124 -15738
rect -928 -15606 -858 -15566
rect -928 -15738 -912 -15606
rect -874 -15738 -858 -15606
rect -928 -15748 -858 -15738
rect -2218 -16774 -2148 -16768
rect -2218 -16900 -2202 -16774
rect -2164 -16900 -2148 -16774
rect -2218 -16938 -2148 -16900
rect -1978 -16774 -1908 -16768
rect -1978 -16900 -1962 -16774
rect -1924 -16900 -1908 -16774
rect -1978 -16938 -1908 -16900
rect -1738 -16774 -1668 -16768
rect -1738 -16900 -1722 -16774
rect -1684 -16900 -1668 -16774
rect -1738 -16938 -1668 -16900
rect -1498 -16774 -1428 -16768
rect -1498 -16900 -1482 -16774
rect -1444 -16900 -1428 -16774
rect -1498 -16938 -1428 -16900
rect -2218 -17576 -2148 -17538
rect -2218 -17708 -2202 -17576
rect -2164 -17708 -2148 -17576
rect -2218 -17746 -2148 -17708
rect -1978 -17576 -1908 -17538
rect -1978 -17708 -1962 -17576
rect -1924 -17708 -1908 -17576
rect -1978 -17746 -1908 -17708
rect -1738 -17576 -1668 -17538
rect -1738 -17708 -1722 -17576
rect -1684 -17708 -1668 -17576
rect -1738 -17746 -1668 -17708
rect -1498 -17576 -1428 -17538
rect -1498 -17708 -1482 -17576
rect -1444 -17708 -1428 -17576
rect -1498 -17746 -1428 -17708
rect -2218 -18384 -2148 -18346
rect -2218 -18516 -2202 -18384
rect -2164 -18516 -2148 -18384
rect -1978 -18384 -1908 -18346
rect -1978 -18516 -1962 -18384
rect -1924 -18516 -1908 -18384
rect -1738 -18384 -1668 -18346
rect -1738 -18516 -1722 -18384
rect -1684 -18516 -1668 -18384
rect -1498 -18384 -1428 -18346
rect -1498 -18516 -1482 -18384
rect -1444 -18516 -1428 -18384
<< polycont >>
rect -6522 -4188 -6484 -4056
rect -6282 -4188 -6244 -4056
rect -6042 -4188 -6004 -4056
rect -5802 -4188 -5764 -4056
rect -5562 -4188 -5524 -4056
rect -5322 -4188 -5284 -4056
rect -5082 -4188 -5044 -4056
rect -4842 -4188 -4804 -4056
rect -4602 -4188 -4564 -4056
rect -4362 -4188 -4324 -4056
rect -4122 -4188 -4084 -4056
rect -3882 -4188 -3844 -4056
rect -3642 -4188 -3604 -4056
rect -3402 -4188 -3364 -4056
rect -3162 -4188 -3124 -4056
rect -2922 -4188 -2884 -4056
rect -2682 -4188 -2644 -4056
rect -2442 -4188 -2404 -4056
rect -2202 -4188 -2164 -4056
rect -1962 -4188 -1924 -4056
rect -1722 -4188 -1684 -4056
rect -1482 -4188 -1444 -4056
rect -1242 -4188 -1204 -4056
rect -1002 -4188 -964 -4056
rect -762 -4188 -724 -4056
rect -522 -4188 -484 -4056
rect -282 -4188 -244 -4056
rect -42 -4188 -4 -4056
rect 198 -4188 236 -4056
rect 438 -4188 476 -4056
rect 678 -4188 716 -4056
rect 918 -4188 956 -4056
rect 1158 -4188 1196 -4056
rect 1398 -4188 1436 -4056
rect 1638 -4188 1676 -4056
rect 1878 -4188 1916 -4056
rect 2118 -4188 2156 -4056
rect 2358 -4188 2396 -4056
rect 2598 -4188 2636 -4056
rect 2838 -4188 2876 -4056
rect -6522 -4996 -6484 -4864
rect -6282 -4996 -6244 -4864
rect -6042 -4996 -6004 -4864
rect -5802 -4996 -5764 -4864
rect -5562 -4996 -5524 -4864
rect -5322 -4996 -5284 -4864
rect -5082 -4996 -5044 -4864
rect -4842 -4996 -4804 -4864
rect -4602 -4996 -4564 -4864
rect -4362 -4996 -4324 -4864
rect -4122 -4996 -4084 -4864
rect -3882 -4996 -3844 -4864
rect -3642 -4996 -3604 -4864
rect -3402 -4996 -3364 -4864
rect -3162 -4996 -3124 -4864
rect -2922 -4996 -2884 -4864
rect -2682 -4996 -2644 -4864
rect -2442 -4996 -2404 -4864
rect -2202 -4996 -2164 -4864
rect -1962 -4996 -1924 -4864
rect -1722 -4996 -1684 -4864
rect -1482 -4996 -1444 -4864
rect -1242 -4996 -1204 -4864
rect -1002 -4996 -964 -4864
rect -762 -4996 -724 -4864
rect -522 -4996 -484 -4864
rect -282 -4996 -244 -4864
rect -42 -4996 -4 -4864
rect 198 -4996 236 -4864
rect 438 -4996 476 -4864
rect 678 -4996 716 -4864
rect 918 -4996 956 -4864
rect 1158 -4996 1196 -4864
rect 1398 -4996 1436 -4864
rect 1638 -4996 1676 -4864
rect 1878 -4996 1916 -4864
rect 2118 -4996 2156 -4864
rect 2358 -4996 2396 -4864
rect 2598 -4996 2636 -4864
rect 2838 -4996 2876 -4864
rect -6522 -5804 -6484 -5672
rect -6282 -5804 -6244 -5672
rect -6042 -5804 -6004 -5672
rect -5802 -5804 -5764 -5672
rect -5562 -5804 -5524 -5672
rect -5322 -5804 -5284 -5672
rect -5082 -5804 -5044 -5672
rect -4842 -5804 -4804 -5672
rect -4602 -5804 -4564 -5672
rect -4362 -5804 -4324 -5672
rect -4122 -5804 -4084 -5672
rect -3882 -5804 -3844 -5672
rect -3642 -5804 -3604 -5672
rect -3402 -5804 -3364 -5672
rect -3162 -5804 -3124 -5672
rect -2922 -5804 -2884 -5672
rect -2682 -5804 -2644 -5672
rect -2442 -5804 -2404 -5672
rect -2202 -5804 -2164 -5672
rect -1962 -5804 -1924 -5672
rect -1722 -5804 -1684 -5672
rect -1482 -5804 -1444 -5672
rect -1242 -5804 -1204 -5672
rect -1002 -5804 -964 -5672
rect -762 -5804 -724 -5672
rect -522 -5804 -484 -5672
rect -282 -5804 -244 -5672
rect -42 -5804 -4 -5672
rect 198 -5804 236 -5672
rect 438 -5804 476 -5672
rect 678 -5804 716 -5672
rect 918 -5804 956 -5672
rect 1158 -5804 1196 -5672
rect 1398 -5804 1436 -5672
rect 1638 -5804 1676 -5672
rect 1878 -5804 1916 -5672
rect 2118 -5804 2156 -5672
rect 2358 -5804 2396 -5672
rect 2598 -5804 2636 -5672
rect 2838 -5804 2876 -5672
rect -15826 -8253 -15458 -8219
rect -15238 -8253 -14870 -8219
rect -14650 -8253 -14282 -8219
rect -14062 -8253 -13694 -8219
rect -13474 -8253 -13106 -8219
rect -12886 -8253 -12518 -8219
rect -12298 -8253 -11930 -8219
rect -11710 -8253 -11342 -8219
rect -11122 -8253 -10754 -8219
rect -10534 -8253 -10166 -8219
rect -9946 -8253 -9578 -8219
rect -9358 -8253 -8990 -8219
rect -8770 -8253 -8402 -8219
rect -8182 -8253 -7814 -8219
rect -7594 -8253 -7226 -8219
rect -7006 -8253 -6638 -8219
rect -6418 -8253 -6050 -8219
rect -5830 -8253 -5462 -8219
rect -5242 -8253 -4874 -8219
rect -4654 -8253 -4286 -8219
rect -4066 -8253 -3698 -8219
rect -3478 -8253 -3110 -8219
rect -2890 -8253 -2522 -8219
rect -2302 -8253 -1934 -8219
rect -1714 -8253 -1346 -8219
rect -1126 -8253 -758 -8219
rect -538 -8253 -170 -8219
rect 50 -8253 418 -8219
rect 638 -8253 1006 -8219
rect 1226 -8253 1594 -8219
rect 1814 -8253 2182 -8219
rect 2402 -8253 2770 -8219
rect 2990 -8253 3358 -8219
rect 3578 -8253 3946 -8219
rect 4166 -8253 4534 -8219
rect 4754 -8253 5122 -8219
rect 5342 -8253 5710 -8219
rect 5930 -8253 6298 -8219
rect 6518 -8253 6886 -8219
rect 7106 -8253 7474 -8219
rect 7694 -8253 8062 -8219
rect 8282 -8253 8650 -8219
rect 8870 -8253 9238 -8219
rect 9458 -8253 9826 -8219
rect 10046 -8253 10414 -8219
rect 10634 -8253 11002 -8219
rect 11222 -8253 11590 -8219
rect 11810 -8253 12178 -8219
rect -15826 -9181 -15458 -9147
rect -15826 -9253 -15458 -9219
rect -15238 -9181 -14870 -9147
rect -15238 -9253 -14870 -9219
rect -14650 -9181 -14282 -9147
rect -14650 -9253 -14282 -9219
rect -14062 -9181 -13694 -9147
rect -14062 -9253 -13694 -9219
rect -13474 -9181 -13106 -9147
rect -13474 -9253 -13106 -9219
rect -12886 -9181 -12518 -9147
rect -12886 -9253 -12518 -9219
rect -12298 -9181 -11930 -9147
rect -12298 -9253 -11930 -9219
rect -11710 -9181 -11342 -9147
rect -11710 -9253 -11342 -9219
rect -11122 -9181 -10754 -9147
rect -11122 -9253 -10754 -9219
rect -10534 -9181 -10166 -9147
rect -10534 -9253 -10166 -9219
rect -9946 -9181 -9578 -9147
rect -9946 -9253 -9578 -9219
rect -9358 -9181 -8990 -9147
rect -9358 -9253 -8990 -9219
rect -8770 -9181 -8402 -9147
rect -8770 -9253 -8402 -9219
rect -8182 -9181 -7814 -9147
rect -8182 -9253 -7814 -9219
rect -7594 -9181 -7226 -9147
rect -7594 -9253 -7226 -9219
rect -7006 -9181 -6638 -9147
rect -7006 -9253 -6638 -9219
rect -6418 -9181 -6050 -9147
rect -6418 -9253 -6050 -9219
rect -5830 -9181 -5462 -9147
rect -5830 -9253 -5462 -9219
rect -5242 -9181 -4874 -9147
rect -5242 -9253 -4874 -9219
rect -4654 -9181 -4286 -9147
rect -4654 -9253 -4286 -9219
rect -4066 -9181 -3698 -9147
rect -4066 -9253 -3698 -9219
rect -3478 -9181 -3110 -9147
rect -3478 -9253 -3110 -9219
rect -2890 -9181 -2522 -9147
rect -2890 -9253 -2522 -9219
rect -2302 -9181 -1934 -9147
rect -2302 -9253 -1934 -9219
rect -1714 -9181 -1346 -9147
rect -1714 -9253 -1346 -9219
rect -1126 -9181 -758 -9147
rect -1126 -9253 -758 -9219
rect -538 -9181 -170 -9147
rect -538 -9253 -170 -9219
rect 50 -9181 418 -9147
rect 50 -9253 418 -9219
rect 638 -9181 1006 -9147
rect 638 -9253 1006 -9219
rect 1226 -9181 1594 -9147
rect 1226 -9253 1594 -9219
rect 1814 -9181 2182 -9147
rect 1814 -9253 2182 -9219
rect 2402 -9181 2770 -9147
rect 2402 -9253 2770 -9219
rect 2990 -9181 3358 -9147
rect 2990 -9253 3358 -9219
rect 3578 -9181 3946 -9147
rect 3578 -9253 3946 -9219
rect 4166 -9181 4534 -9147
rect 4166 -9253 4534 -9219
rect 4754 -9181 5122 -9147
rect 4754 -9253 5122 -9219
rect 5342 -9181 5710 -9147
rect 5342 -9253 5710 -9219
rect 5930 -9181 6298 -9147
rect 5930 -9253 6298 -9219
rect 6518 -9181 6886 -9147
rect 6518 -9253 6886 -9219
rect 7106 -9181 7474 -9147
rect 7106 -9253 7474 -9219
rect 7694 -9181 8062 -9147
rect 7694 -9253 8062 -9219
rect 8282 -9181 8650 -9147
rect 8282 -9253 8650 -9219
rect 8870 -9181 9238 -9147
rect 8870 -9253 9238 -9219
rect 9458 -9181 9826 -9147
rect 9458 -9253 9826 -9219
rect 10046 -9181 10414 -9147
rect 10046 -9253 10414 -9219
rect 10634 -9181 11002 -9147
rect 10634 -9253 11002 -9219
rect 11222 -9181 11590 -9147
rect 11222 -9253 11590 -9219
rect 11810 -9181 12178 -9147
rect 11810 -9253 12178 -9219
rect -15826 -10181 -15458 -10147
rect -15826 -10253 -15458 -10219
rect -15238 -10181 -14870 -10147
rect -15238 -10253 -14870 -10219
rect -14650 -10181 -14282 -10147
rect -14650 -10253 -14282 -10219
rect -14062 -10181 -13694 -10147
rect -14062 -10253 -13694 -10219
rect -13474 -10181 -13106 -10147
rect -13474 -10253 -13106 -10219
rect -12886 -10181 -12518 -10147
rect -12886 -10253 -12518 -10219
rect -12298 -10181 -11930 -10147
rect -12298 -10253 -11930 -10219
rect -11710 -10181 -11342 -10147
rect -11710 -10253 -11342 -10219
rect -11122 -10181 -10754 -10147
rect -11122 -10253 -10754 -10219
rect -10534 -10181 -10166 -10147
rect -10534 -10253 -10166 -10219
rect -9946 -10181 -9578 -10147
rect -9946 -10253 -9578 -10219
rect -9358 -10181 -8990 -10147
rect -9358 -10253 -8990 -10219
rect -8770 -10181 -8402 -10147
rect -8770 -10253 -8402 -10219
rect -8182 -10181 -7814 -10147
rect -8182 -10253 -7814 -10219
rect -7594 -10181 -7226 -10147
rect -7594 -10253 -7226 -10219
rect -7006 -10181 -6638 -10147
rect -7006 -10253 -6638 -10219
rect -6418 -10181 -6050 -10147
rect -6418 -10253 -6050 -10219
rect -5830 -10181 -5462 -10147
rect -5830 -10253 -5462 -10219
rect -5242 -10181 -4874 -10147
rect -5242 -10253 -4874 -10219
rect -4654 -10181 -4286 -10147
rect -4654 -10253 -4286 -10219
rect -4066 -10181 -3698 -10147
rect -4066 -10253 -3698 -10219
rect -3478 -10181 -3110 -10147
rect -3478 -10253 -3110 -10219
rect -2890 -10181 -2522 -10147
rect -2890 -10253 -2522 -10219
rect -2302 -10181 -1934 -10147
rect -2302 -10253 -1934 -10219
rect -1714 -10181 -1346 -10147
rect -1714 -10253 -1346 -10219
rect -1126 -10181 -758 -10147
rect -1126 -10253 -758 -10219
rect -538 -10181 -170 -10147
rect -538 -10253 -170 -10219
rect 50 -10181 418 -10147
rect 50 -10253 418 -10219
rect 638 -10181 1006 -10147
rect 638 -10253 1006 -10219
rect 1226 -10181 1594 -10147
rect 1226 -10253 1594 -10219
rect 1814 -10181 2182 -10147
rect 1814 -10253 2182 -10219
rect 2402 -10181 2770 -10147
rect 2402 -10253 2770 -10219
rect 2990 -10181 3358 -10147
rect 2990 -10253 3358 -10219
rect 3578 -10181 3946 -10147
rect 3578 -10253 3946 -10219
rect 4166 -10181 4534 -10147
rect 4166 -10253 4534 -10219
rect 4754 -10181 5122 -10147
rect 4754 -10253 5122 -10219
rect 5342 -10181 5710 -10147
rect 5342 -10253 5710 -10219
rect 5930 -10181 6298 -10147
rect 5930 -10253 6298 -10219
rect 6518 -10181 6886 -10147
rect 6518 -10253 6886 -10219
rect 7106 -10181 7474 -10147
rect 7106 -10253 7474 -10219
rect 7694 -10181 8062 -10147
rect 7694 -10253 8062 -10219
rect 8282 -10181 8650 -10147
rect 8282 -10253 8650 -10219
rect 8870 -10181 9238 -10147
rect 8870 -10253 9238 -10219
rect 9458 -10181 9826 -10147
rect 9458 -10253 9826 -10219
rect 10046 -10181 10414 -10147
rect 10046 -10253 10414 -10219
rect 10634 -10181 11002 -10147
rect 10634 -10253 11002 -10219
rect 11222 -10181 11590 -10147
rect 11222 -10253 11590 -10219
rect 11810 -10181 12178 -10147
rect 11810 -10253 12178 -10219
rect -15826 -11181 -15458 -11147
rect -15238 -11181 -14870 -11147
rect -14650 -11181 -14282 -11147
rect -14062 -11181 -13694 -11147
rect -13474 -11181 -13106 -11147
rect -12886 -11181 -12518 -11147
rect -12298 -11181 -11930 -11147
rect -11710 -11181 -11342 -11147
rect -11122 -11181 -10754 -11147
rect -10534 -11181 -10166 -11147
rect -9946 -11181 -9578 -11147
rect -9358 -11181 -8990 -11147
rect -8770 -11181 -8402 -11147
rect -8182 -11181 -7814 -11147
rect -7594 -11181 -7226 -11147
rect -7006 -11181 -6638 -11147
rect -6418 -11181 -6050 -11147
rect -5830 -11181 -5462 -11147
rect -5242 -11181 -4874 -11147
rect -4654 -11181 -4286 -11147
rect -4066 -11181 -3698 -11147
rect -3478 -11181 -3110 -11147
rect -2890 -11181 -2522 -11147
rect -2302 -11181 -1934 -11147
rect -1714 -11181 -1346 -11147
rect -1126 -11181 -758 -11147
rect -538 -11181 -170 -11147
rect 50 -11181 418 -11147
rect 638 -11181 1006 -11147
rect 1226 -11181 1594 -11147
rect 1814 -11181 2182 -11147
rect 2402 -11181 2770 -11147
rect 2990 -11181 3358 -11147
rect 3578 -11181 3946 -11147
rect 4166 -11181 4534 -11147
rect 4754 -11181 5122 -11147
rect 5342 -11181 5710 -11147
rect 5930 -11181 6298 -11147
rect 6518 -11181 6886 -11147
rect 7106 -11181 7474 -11147
rect 7694 -11181 8062 -11147
rect 8282 -11181 8650 -11147
rect 8870 -11181 9238 -11147
rect 9458 -11181 9826 -11147
rect 10046 -11181 10414 -11147
rect 10634 -11181 11002 -11147
rect 11222 -11181 11590 -11147
rect 11810 -11181 12178 -11147
rect -2774 -12708 -2736 -12576
rect -2508 -12708 -2470 -12576
rect -2242 -12708 -2204 -12576
rect -1976 -12708 -1938 -12576
rect -1710 -12708 -1672 -12576
rect -1444 -12708 -1406 -12576
rect -1178 -12708 -1140 -12576
rect -912 -12708 -874 -12576
rect -2774 -13718 -2736 -13586
rect -2508 -13718 -2470 -13586
rect -2242 -13718 -2204 -13586
rect -1976 -13718 -1938 -13586
rect -1710 -13718 -1672 -13586
rect -1444 -13718 -1406 -13586
rect -1178 -13718 -1140 -13586
rect -912 -13718 -874 -13586
rect -2774 -14728 -2736 -14596
rect -2508 -14728 -2470 -14596
rect -2242 -14728 -2204 -14596
rect -1976 -14728 -1938 -14596
rect -1710 -14728 -1672 -14596
rect -1444 -14728 -1406 -14596
rect -1178 -14728 -1140 -14596
rect -912 -14728 -874 -14596
rect -2774 -15738 -2736 -15606
rect -2508 -15738 -2470 -15606
rect -2242 -15738 -2204 -15606
rect -1976 -15738 -1938 -15606
rect -1710 -15738 -1672 -15606
rect -1444 -15738 -1406 -15606
rect -1178 -15738 -1140 -15606
rect -912 -15738 -874 -15606
rect -2202 -16900 -2164 -16774
rect -1962 -16900 -1924 -16774
rect -1722 -16900 -1684 -16774
rect -1482 -16900 -1444 -16774
rect -2202 -17708 -2164 -17576
rect -1962 -17708 -1924 -17576
rect -1722 -17708 -1684 -17576
rect -1482 -17708 -1444 -17576
rect -2202 -18516 -2164 -18384
rect -1962 -18516 -1924 -18384
rect -1722 -18516 -1684 -18384
rect -1482 -18516 -1444 -18384
<< xpolycontact >>
rect 4367 -15411 4437 -14979
rect 4367 -15943 4437 -15511
<< xpolyres >>
rect 4367 -15511 4437 -15411
<< locali >>
rect -6930 -3746 -6842 -3712
rect 3196 -3746 3284 -3712
rect -6930 -3780 -6896 -3746
rect 3250 -3778 3284 -3746
rect -6538 -4188 -6522 -4056
rect -6484 -4188 -6282 -4056
rect -6244 -4188 -6042 -4056
rect -6004 -4188 -5802 -4056
rect -5764 -4188 -5562 -4056
rect -5524 -4188 -5322 -4056
rect -5284 -4188 -5082 -4056
rect -5044 -4188 -4842 -4056
rect -4804 -4188 -4602 -4056
rect -4564 -4188 -4362 -4056
rect -4324 -4188 -4122 -4056
rect -4084 -4188 -3882 -4056
rect -3844 -4188 -3642 -4056
rect -3604 -4188 -3402 -4056
rect -3364 -4188 -3162 -4056
rect -3124 -4188 -2922 -4056
rect -2884 -4188 -2682 -4056
rect -2644 -4188 -2442 -4056
rect -2404 -4188 -2202 -4056
rect -2164 -4188 -1962 -4056
rect -1924 -4188 -1722 -4056
rect -1684 -4188 -1482 -4056
rect -1444 -4188 -1242 -4056
rect -1204 -4188 -1002 -4056
rect -964 -4188 -762 -4056
rect -724 -4188 -522 -4056
rect -484 -4188 -282 -4056
rect -244 -4188 -42 -4056
rect -4 -4188 198 -4056
rect 236 -4188 438 -4056
rect 476 -4188 678 -4056
rect 716 -4188 918 -4056
rect 956 -4188 1158 -4056
rect 1196 -4188 1398 -4056
rect 1436 -4188 1638 -4056
rect 1676 -4188 1878 -4056
rect 1916 -4188 2118 -4056
rect 2156 -4188 2358 -4056
rect 2396 -4188 2598 -4056
rect 2636 -4188 2838 -4056
rect 2876 -4188 2902 -4056
rect -6584 -4238 -6550 -4222
rect -6584 -4830 -6550 -4814
rect -6456 -4238 -6422 -4222
rect -6456 -4830 -6422 -4814
rect -6344 -4238 -6310 -4222
rect -6344 -4830 -6310 -4814
rect -6216 -4238 -6182 -4222
rect -6216 -4830 -6182 -4814
rect -6104 -4238 -6070 -4222
rect -6104 -4830 -6070 -4814
rect -5976 -4238 -5942 -4222
rect -5976 -4830 -5942 -4814
rect -5864 -4238 -5830 -4222
rect -5864 -4830 -5830 -4814
rect -5736 -4238 -5702 -4222
rect -5736 -4830 -5702 -4814
rect -5624 -4238 -5590 -4222
rect -5624 -4830 -5590 -4814
rect -5496 -4238 -5462 -4222
rect -5496 -4830 -5462 -4814
rect -5384 -4238 -5350 -4222
rect -5384 -4830 -5350 -4814
rect -5256 -4238 -5222 -4222
rect -5256 -4830 -5222 -4814
rect -5144 -4238 -5110 -4222
rect -5144 -4830 -5110 -4814
rect -5016 -4238 -4982 -4222
rect -5016 -4830 -4982 -4814
rect -4904 -4238 -4870 -4222
rect -4904 -4830 -4870 -4814
rect -4776 -4238 -4742 -4222
rect -4776 -4830 -4742 -4814
rect -4664 -4238 -4630 -4222
rect -4664 -4830 -4630 -4814
rect -4536 -4238 -4502 -4222
rect -4536 -4830 -4502 -4814
rect -4424 -4238 -4390 -4222
rect -4424 -4830 -4390 -4814
rect -4296 -4238 -4262 -4222
rect -4296 -4830 -4262 -4814
rect -4184 -4238 -4150 -4222
rect -4184 -4830 -4150 -4814
rect -4056 -4238 -4022 -4222
rect -4056 -4830 -4022 -4814
rect -3944 -4238 -3910 -4222
rect -3944 -4830 -3910 -4814
rect -3816 -4238 -3782 -4222
rect -3816 -4830 -3782 -4814
rect -3704 -4238 -3670 -4222
rect -3704 -4830 -3670 -4814
rect -3576 -4238 -3542 -4222
rect -3576 -4830 -3542 -4814
rect -3464 -4238 -3430 -4222
rect -3464 -4830 -3430 -4814
rect -3336 -4238 -3302 -4222
rect -3336 -4830 -3302 -4814
rect -3224 -4238 -3190 -4222
rect -3224 -4830 -3190 -4814
rect -3096 -4238 -3062 -4222
rect -3096 -4830 -3062 -4814
rect -2984 -4238 -2950 -4222
rect -2984 -4830 -2950 -4814
rect -2856 -4238 -2822 -4222
rect -2856 -4830 -2822 -4814
rect -2744 -4238 -2710 -4222
rect -2744 -4830 -2710 -4814
rect -2616 -4238 -2582 -4222
rect -2616 -4830 -2582 -4814
rect -2504 -4238 -2470 -4222
rect -2504 -4830 -2470 -4814
rect -2376 -4238 -2342 -4222
rect -2376 -4830 -2342 -4814
rect -2264 -4238 -2230 -4222
rect -2264 -4830 -2230 -4814
rect -2136 -4238 -2102 -4222
rect -2136 -4830 -2102 -4814
rect -2024 -4238 -1990 -4222
rect -2024 -4830 -1990 -4814
rect -1896 -4238 -1862 -4222
rect -1896 -4830 -1862 -4814
rect -1784 -4238 -1750 -4222
rect -1784 -4830 -1750 -4814
rect -1656 -4238 -1622 -4222
rect -1656 -4830 -1622 -4814
rect -1544 -4238 -1510 -4222
rect -1544 -4830 -1510 -4814
rect -1416 -4238 -1382 -4222
rect -1416 -4830 -1382 -4814
rect -1304 -4238 -1270 -4222
rect -1304 -4830 -1270 -4814
rect -1176 -4238 -1142 -4222
rect -1176 -4830 -1142 -4814
rect -1064 -4238 -1030 -4222
rect -1064 -4830 -1030 -4814
rect -936 -4238 -902 -4222
rect -936 -4830 -902 -4814
rect -824 -4238 -790 -4222
rect -824 -4830 -790 -4814
rect -696 -4238 -662 -4222
rect -696 -4830 -662 -4814
rect -584 -4238 -550 -4222
rect -584 -4830 -550 -4814
rect -456 -4238 -422 -4222
rect -456 -4830 -422 -4814
rect -344 -4238 -310 -4222
rect -344 -4830 -310 -4814
rect -216 -4238 -182 -4222
rect -216 -4830 -182 -4814
rect -104 -4238 -70 -4222
rect -104 -4830 -70 -4814
rect 24 -4238 58 -4222
rect 24 -4830 58 -4814
rect 136 -4238 170 -4222
rect 136 -4830 170 -4814
rect 264 -4238 298 -4222
rect 264 -4830 298 -4814
rect 376 -4238 410 -4222
rect 376 -4830 410 -4814
rect 504 -4238 538 -4222
rect 504 -4830 538 -4814
rect 616 -4238 650 -4222
rect 616 -4830 650 -4814
rect 744 -4238 778 -4222
rect 744 -4830 778 -4814
rect 856 -4238 890 -4222
rect 856 -4830 890 -4814
rect 984 -4238 1018 -4222
rect 984 -4830 1018 -4814
rect 1096 -4238 1130 -4222
rect 1096 -4830 1130 -4814
rect 1224 -4238 1258 -4222
rect 1224 -4830 1258 -4814
rect 1336 -4238 1370 -4222
rect 1336 -4830 1370 -4814
rect 1464 -4238 1498 -4222
rect 1464 -4830 1498 -4814
rect 1576 -4238 1610 -4222
rect 1576 -4830 1610 -4814
rect 1704 -4238 1738 -4222
rect 1704 -4830 1738 -4814
rect 1816 -4238 1850 -4222
rect 1816 -4830 1850 -4814
rect 1944 -4238 1978 -4222
rect 1944 -4830 1978 -4814
rect 2056 -4238 2090 -4222
rect 2056 -4830 2090 -4814
rect 2184 -4238 2218 -4222
rect 2184 -4830 2218 -4814
rect 2296 -4238 2330 -4222
rect 2296 -4830 2330 -4814
rect 2424 -4238 2458 -4222
rect 2424 -4830 2458 -4814
rect 2536 -4238 2570 -4222
rect 2536 -4830 2570 -4814
rect 2664 -4238 2698 -4222
rect 2664 -4830 2698 -4814
rect 2776 -4238 2810 -4222
rect 2776 -4830 2810 -4814
rect 2904 -4238 2938 -4222
rect 2904 -4830 2938 -4814
rect -6538 -4996 -6522 -4864
rect -6484 -4996 -6282 -4864
rect -6244 -4996 -6042 -4864
rect -6004 -4996 -5802 -4864
rect -5764 -4996 -5562 -4864
rect -5524 -4996 -5322 -4864
rect -5284 -4996 -5082 -4864
rect -5044 -4996 -4842 -4864
rect -4804 -4996 -4602 -4864
rect -4564 -4996 -4362 -4864
rect -4324 -4996 -4122 -4864
rect -4084 -4996 -3882 -4864
rect -3844 -4996 -3642 -4864
rect -3604 -4996 -3402 -4864
rect -3364 -4996 -3162 -4864
rect -3124 -4996 -2922 -4864
rect -2884 -4996 -2682 -4864
rect -2644 -4996 -2442 -4864
rect -2404 -4996 -2202 -4864
rect -2164 -4996 -1962 -4864
rect -1924 -4996 -1722 -4864
rect -1684 -4996 -1482 -4864
rect -1444 -4996 -1242 -4864
rect -1204 -4996 -1002 -4864
rect -964 -4996 -762 -4864
rect -724 -4996 -522 -4864
rect -484 -4996 -282 -4864
rect -244 -4996 -42 -4864
rect -4 -4996 198 -4864
rect 236 -4996 438 -4864
rect 476 -4996 678 -4864
rect 716 -4996 918 -4864
rect 956 -4996 1158 -4864
rect 1196 -4996 1398 -4864
rect 1436 -4996 1638 -4864
rect 1676 -4996 1878 -4864
rect 1916 -4996 2118 -4864
rect 2156 -4996 2358 -4864
rect 2396 -4996 2598 -4864
rect 2636 -4996 2838 -4864
rect 2876 -4996 2902 -4864
rect -6584 -5046 -6550 -5030
rect -6584 -5638 -6550 -5622
rect -6456 -5046 -6422 -5030
rect -6456 -5638 -6422 -5622
rect -6344 -5046 -6310 -5030
rect -6344 -5638 -6310 -5622
rect -6216 -5046 -6182 -5030
rect -6216 -5638 -6182 -5622
rect -6104 -5046 -6070 -5030
rect -6104 -5638 -6070 -5622
rect -5976 -5046 -5942 -5030
rect -5976 -5638 -5942 -5622
rect -5864 -5046 -5830 -5030
rect -5864 -5638 -5830 -5622
rect -5736 -5046 -5702 -5030
rect -5736 -5638 -5702 -5622
rect -5624 -5046 -5590 -5030
rect -5624 -5638 -5590 -5622
rect -5496 -5046 -5462 -5030
rect -5496 -5638 -5462 -5622
rect -5384 -5046 -5350 -5030
rect -5384 -5638 -5350 -5622
rect -5256 -5046 -5222 -5030
rect -5256 -5638 -5222 -5622
rect -5144 -5046 -5110 -5030
rect -5144 -5638 -5110 -5622
rect -5016 -5046 -4982 -5030
rect -5016 -5638 -4982 -5622
rect -4904 -5046 -4870 -5030
rect -4904 -5638 -4870 -5622
rect -4776 -5046 -4742 -5030
rect -4776 -5638 -4742 -5622
rect -4664 -5046 -4630 -5030
rect -4664 -5638 -4630 -5622
rect -4536 -5046 -4502 -5030
rect -4536 -5638 -4502 -5622
rect -4424 -5046 -4390 -5030
rect -4424 -5638 -4390 -5622
rect -4296 -5046 -4262 -5030
rect -4296 -5638 -4262 -5622
rect -4184 -5046 -4150 -5030
rect -4184 -5638 -4150 -5622
rect -4056 -5046 -4022 -5030
rect -4056 -5638 -4022 -5622
rect -3944 -5046 -3910 -5030
rect -3944 -5638 -3910 -5622
rect -3816 -5046 -3782 -5030
rect -3816 -5638 -3782 -5622
rect -3704 -5046 -3670 -5030
rect -3704 -5638 -3670 -5622
rect -3576 -5046 -3542 -5030
rect -3576 -5638 -3542 -5622
rect -3464 -5046 -3430 -5030
rect -3464 -5638 -3430 -5622
rect -3336 -5046 -3302 -5030
rect -3336 -5638 -3302 -5622
rect -3224 -5046 -3190 -5030
rect -3224 -5638 -3190 -5622
rect -3096 -5046 -3062 -5030
rect -3096 -5638 -3062 -5622
rect -2984 -5046 -2950 -5030
rect -2984 -5638 -2950 -5622
rect -2856 -5046 -2822 -5030
rect -2856 -5638 -2822 -5622
rect -2744 -5046 -2710 -5030
rect -2744 -5638 -2710 -5622
rect -2616 -5046 -2582 -5030
rect -2616 -5638 -2582 -5622
rect -2504 -5046 -2470 -5030
rect -2504 -5638 -2470 -5622
rect -2376 -5046 -2342 -5030
rect -2376 -5638 -2342 -5622
rect -2264 -5046 -2230 -5030
rect -2264 -5638 -2230 -5622
rect -2136 -5046 -2102 -5030
rect -2136 -5638 -2102 -5622
rect -2024 -5046 -1990 -5030
rect -2024 -5638 -1990 -5622
rect -1896 -5046 -1862 -5030
rect -1896 -5638 -1862 -5622
rect -1784 -5046 -1750 -5030
rect -1784 -5638 -1750 -5622
rect -1656 -5046 -1622 -5030
rect -1656 -5638 -1622 -5622
rect -1544 -5046 -1510 -5030
rect -1544 -5638 -1510 -5622
rect -1416 -5046 -1382 -5030
rect -1416 -5638 -1382 -5622
rect -1304 -5046 -1270 -5030
rect -1304 -5638 -1270 -5622
rect -1176 -5046 -1142 -5030
rect -1176 -5638 -1142 -5622
rect -1064 -5046 -1030 -5030
rect -1064 -5638 -1030 -5622
rect -936 -5046 -902 -5030
rect -936 -5638 -902 -5622
rect -824 -5046 -790 -5030
rect -824 -5638 -790 -5622
rect -696 -5046 -662 -5030
rect -696 -5638 -662 -5622
rect -584 -5046 -550 -5030
rect -584 -5638 -550 -5622
rect -456 -5046 -422 -5030
rect -456 -5638 -422 -5622
rect -344 -5046 -310 -5030
rect -344 -5638 -310 -5622
rect -216 -5046 -182 -5030
rect -216 -5638 -182 -5622
rect -104 -5046 -70 -5030
rect -104 -5638 -70 -5622
rect 24 -5046 58 -5030
rect 24 -5638 58 -5622
rect 136 -5046 170 -5030
rect 136 -5638 170 -5622
rect 264 -5046 298 -5030
rect 264 -5638 298 -5622
rect 376 -5046 410 -5030
rect 376 -5638 410 -5622
rect 504 -5046 538 -5030
rect 504 -5638 538 -5622
rect 616 -5046 650 -5030
rect 616 -5638 650 -5622
rect 744 -5046 778 -5030
rect 744 -5638 778 -5622
rect 856 -5046 890 -5030
rect 856 -5638 890 -5622
rect 984 -5046 1018 -5030
rect 984 -5638 1018 -5622
rect 1096 -5046 1130 -5030
rect 1096 -5638 1130 -5622
rect 1224 -5046 1258 -5030
rect 1224 -5638 1258 -5622
rect 1336 -5046 1370 -5030
rect 1336 -5638 1370 -5622
rect 1464 -5046 1498 -5030
rect 1464 -5638 1498 -5622
rect 1576 -5046 1610 -5030
rect 1576 -5638 1610 -5622
rect 1704 -5046 1738 -5030
rect 1704 -5638 1738 -5622
rect 1816 -5046 1850 -5030
rect 1816 -5638 1850 -5622
rect 1944 -5046 1978 -5030
rect 1944 -5638 1978 -5622
rect 2056 -5046 2090 -5030
rect 2056 -5638 2090 -5622
rect 2184 -5046 2218 -5030
rect 2184 -5638 2218 -5622
rect 2296 -5046 2330 -5030
rect 2296 -5638 2330 -5622
rect 2424 -5046 2458 -5030
rect 2424 -5638 2458 -5622
rect 2536 -5046 2570 -5030
rect 2536 -5638 2570 -5622
rect 2664 -5046 2698 -5030
rect 2664 -5638 2698 -5622
rect 2776 -5046 2810 -5030
rect 2776 -5638 2810 -5622
rect 2904 -5046 2938 -5030
rect 2904 -5638 2938 -5622
rect -6538 -5804 -6522 -5672
rect -6484 -5804 -6282 -5672
rect -6244 -5804 -6042 -5672
rect -6004 -5804 -5802 -5672
rect -5764 -5804 -5562 -5672
rect -5524 -5804 -5322 -5672
rect -5284 -5804 -5082 -5672
rect -5044 -5804 -4842 -5672
rect -4804 -5804 -4602 -5672
rect -4564 -5804 -4362 -5672
rect -4324 -5804 -4122 -5672
rect -4084 -5804 -3882 -5672
rect -3844 -5804 -3642 -5672
rect -3604 -5804 -3402 -5672
rect -3364 -5804 -3162 -5672
rect -3124 -5804 -2922 -5672
rect -2884 -5804 -2682 -5672
rect -2644 -5804 -2442 -5672
rect -2404 -5804 -2202 -5672
rect -2164 -5804 -1962 -5672
rect -1924 -5804 -1722 -5672
rect -1684 -5804 -1482 -5672
rect -1444 -5804 -1242 -5672
rect -1204 -5804 -1002 -5672
rect -964 -5804 -762 -5672
rect -724 -5804 -522 -5672
rect -484 -5804 -282 -5672
rect -244 -5804 -42 -5672
rect -4 -5804 198 -5672
rect 236 -5804 438 -5672
rect 476 -5804 678 -5672
rect 716 -5804 918 -5672
rect 956 -5804 1158 -5672
rect 1196 -5804 1398 -5672
rect 1436 -5804 1638 -5672
rect 1676 -5804 1878 -5672
rect 1916 -5804 2118 -5672
rect 2156 -5804 2358 -5672
rect 2396 -5804 2598 -5672
rect 2636 -5804 2838 -5672
rect 2876 -5804 2902 -5672
rect -6930 -6148 -6896 -6060
rect 3250 -6148 3284 -6060
rect -16234 -7902 -16074 -7868
rect 12448 -7896 12586 -7868
rect 12448 -7902 12552 -7896
rect -16234 -7930 -16200 -7902
rect -15842 -8219 -4082 -8218
rect -3682 -8219 -3494 -8218
rect -3094 -8219 -2906 -8218
rect -2506 -8219 -2318 -8218
rect -1918 -8219 -1730 -8218
rect -1330 -8219 -1142 -8218
rect -742 -8219 -554 -8218
rect -154 -8219 34 -8218
rect 434 -8219 12194 -8218
rect -15842 -8253 -15826 -8219
rect -15458 -8253 -15238 -8219
rect -14870 -8253 -14650 -8219
rect -14282 -8253 -14062 -8219
rect -13694 -8253 -13474 -8219
rect -13106 -8253 -12886 -8219
rect -12518 -8253 -12298 -8219
rect -11930 -8253 -11710 -8219
rect -11342 -8253 -11122 -8219
rect -10754 -8253 -10534 -8219
rect -10166 -8253 -9946 -8219
rect -9578 -8253 -9358 -8219
rect -8990 -8253 -8770 -8219
rect -8402 -8253 -8182 -8219
rect -7814 -8253 -7594 -8219
rect -7226 -8253 -7006 -8219
rect -6638 -8253 -6418 -8219
rect -6050 -8253 -5830 -8219
rect -5462 -8253 -5242 -8219
rect -4874 -8253 -4654 -8219
rect -4286 -8253 -4066 -8219
rect -3698 -8253 -3478 -8219
rect -3110 -8253 -2890 -8219
rect -2522 -8253 -2302 -8219
rect -1934 -8253 -1714 -8219
rect -1346 -8253 -1126 -8219
rect -758 -8253 -538 -8219
rect -170 -8253 50 -8219
rect 418 -8253 638 -8219
rect 1006 -8253 1226 -8219
rect 1594 -8253 1814 -8219
rect 2182 -8253 2402 -8219
rect 2770 -8253 2990 -8219
rect 3358 -8253 3578 -8219
rect 3946 -8253 4166 -8219
rect 4534 -8253 4754 -8219
rect 5122 -8253 5342 -8219
rect 5710 -8253 5930 -8219
rect 6298 -8253 6518 -8219
rect 6886 -8253 7106 -8219
rect 7474 -8253 7694 -8219
rect 8062 -8253 8282 -8219
rect 8650 -8253 8870 -8219
rect 9238 -8253 9458 -8219
rect 9826 -8253 10046 -8219
rect 10414 -8253 10634 -8219
rect 11002 -8253 11222 -8219
rect 11590 -8253 11810 -8219
rect 12178 -8253 12194 -8219
rect -15842 -8254 -4082 -8253
rect -3682 -8254 -3494 -8253
rect -3094 -8254 -2906 -8253
rect -2506 -8254 -2318 -8253
rect -4128 -8296 -4082 -8254
rect -1918 -8296 -1730 -8253
rect -1330 -8254 -1142 -8253
rect -742 -8254 -554 -8253
rect -154 -8254 34 -8253
rect 434 -8254 12194 -8253
rect 434 -8296 480 -8254
rect -15888 -8312 -15854 -8296
rect -15888 -9104 -15854 -9088
rect -15430 -8312 -15396 -8296
rect -15430 -9104 -15396 -9088
rect -15300 -8312 -15266 -8296
rect -15300 -9104 -15266 -9088
rect -14842 -8312 -14808 -8296
rect -14842 -9104 -14808 -9088
rect -14712 -8312 -14678 -8296
rect -14712 -9104 -14678 -9088
rect -14254 -8312 -14220 -8296
rect -14254 -9104 -14220 -9088
rect -14124 -8312 -14090 -8296
rect -14124 -9104 -14090 -9088
rect -13666 -8312 -13632 -8296
rect -13666 -9104 -13632 -9088
rect -13536 -8312 -13502 -8296
rect -13536 -9104 -13502 -9088
rect -13078 -8312 -13044 -8296
rect -13078 -9104 -13044 -9088
rect -12948 -8312 -12914 -8296
rect -12948 -9104 -12914 -9088
rect -12490 -8312 -12456 -8296
rect -12490 -9104 -12456 -9088
rect -12360 -8312 -12326 -8296
rect -12360 -9104 -12326 -9088
rect -11902 -8312 -11868 -8296
rect -11902 -9104 -11868 -9088
rect -11772 -8312 -11738 -8296
rect -11772 -9104 -11738 -9088
rect -11314 -8312 -11280 -8296
rect -11314 -9104 -11280 -9088
rect -11184 -8312 -11150 -8296
rect -11184 -9104 -11150 -9088
rect -10726 -8312 -10692 -8296
rect -10726 -9104 -10692 -9088
rect -10596 -8312 -10562 -8296
rect -10596 -9104 -10562 -9088
rect -10138 -8312 -10104 -8296
rect -10138 -9104 -10104 -9088
rect -10008 -8312 -9974 -8296
rect -10008 -9104 -9974 -9088
rect -9550 -8312 -9516 -8296
rect -9550 -9104 -9516 -9088
rect -9420 -8312 -9386 -8296
rect -9420 -9104 -9386 -9088
rect -8962 -8312 -8928 -8296
rect -8962 -9104 -8928 -9088
rect -8832 -8312 -8798 -8296
rect -8832 -9104 -8798 -9088
rect -8374 -8312 -8340 -8296
rect -8374 -9104 -8340 -9088
rect -8244 -8312 -8210 -8296
rect -8244 -9104 -8210 -9088
rect -7786 -8312 -7752 -8296
rect -7786 -9104 -7752 -9088
rect -7656 -8312 -7622 -8296
rect -7656 -9104 -7622 -9088
rect -7198 -8312 -7164 -8296
rect -7198 -9104 -7164 -9088
rect -7068 -8312 -7034 -8296
rect -7068 -9104 -7034 -9088
rect -6610 -8312 -6576 -8296
rect -6610 -9104 -6576 -9088
rect -6480 -8312 -6446 -8296
rect -6480 -9104 -6446 -9088
rect -6022 -8312 -5988 -8296
rect -6022 -9104 -5988 -9088
rect -5892 -8312 -5858 -8296
rect -5892 -9104 -5858 -9088
rect -5434 -8312 -5400 -8296
rect -5434 -9104 -5400 -9088
rect -5304 -8312 -5270 -8296
rect -5304 -9104 -5270 -9088
rect -4846 -8312 -4812 -8296
rect -4846 -9104 -4812 -9088
rect -4716 -8312 -4682 -8296
rect -4716 -9104 -4682 -9088
rect -4258 -8312 -4224 -8296
rect -4258 -9104 -4224 -9088
rect -4128 -8312 -4094 -8296
rect -4128 -9146 -4094 -9088
rect -3670 -8312 -3636 -8296
rect -3670 -9104 -3636 -9088
rect -3540 -8312 -3506 -8296
rect -3540 -9104 -3506 -9088
rect -3082 -8312 -3048 -8296
rect -3082 -9104 -3048 -9088
rect -2952 -8312 -2918 -8296
rect -2952 -9104 -2918 -9088
rect -2494 -8312 -2460 -8296
rect -2494 -9104 -2460 -9088
rect -2364 -8312 -2330 -8296
rect -2364 -9104 -2330 -9088
rect -1906 -8312 -1742 -8296
rect -1872 -9088 -1776 -8312
rect -1906 -9146 -1742 -9088
rect -1318 -8312 -1284 -8296
rect -1318 -9104 -1284 -9088
rect -1188 -8312 -1154 -8296
rect -1188 -9104 -1154 -9088
rect -730 -8312 -696 -8296
rect -730 -9104 -696 -9088
rect -600 -8312 -566 -8296
rect -600 -9104 -566 -9088
rect -142 -8312 -108 -8296
rect -142 -9104 -108 -9088
rect -12 -8312 22 -8296
rect -12 -9104 22 -9088
rect 446 -8312 480 -8296
rect 446 -9146 480 -9088
rect 576 -8312 610 -8296
rect 576 -9104 610 -9088
rect 1034 -8312 1068 -8296
rect 1034 -9104 1068 -9088
rect 1164 -8312 1198 -8296
rect 1164 -9104 1198 -9088
rect 1622 -8312 1656 -8296
rect 1622 -9104 1656 -9088
rect 1752 -8312 1786 -8296
rect 1752 -9104 1786 -9088
rect 2210 -8312 2244 -8296
rect 2210 -9104 2244 -9088
rect 2340 -8312 2374 -8296
rect 2340 -9104 2374 -9088
rect 2798 -8312 2832 -8296
rect 2798 -9104 2832 -9088
rect 2928 -8312 2962 -8296
rect 2928 -9104 2962 -9088
rect 3386 -8312 3420 -8296
rect 3386 -9104 3420 -9088
rect 3516 -8312 3550 -8296
rect 3516 -9104 3550 -9088
rect 3974 -8312 4008 -8296
rect 3974 -9104 4008 -9088
rect 4104 -8312 4138 -8296
rect 4104 -9104 4138 -9088
rect 4562 -8312 4596 -8296
rect 4562 -9104 4596 -9088
rect 4692 -8312 4726 -8296
rect 4692 -9104 4726 -9088
rect 5150 -8312 5184 -8296
rect 5150 -9104 5184 -9088
rect 5280 -8312 5314 -8296
rect 5280 -9104 5314 -9088
rect 5738 -8312 5772 -8296
rect 5738 -9104 5772 -9088
rect 5868 -8312 5902 -8296
rect 5868 -9104 5902 -9088
rect 6326 -8312 6360 -8296
rect 6326 -9104 6360 -9088
rect 6456 -8312 6490 -8296
rect 6456 -9104 6490 -9088
rect 6914 -8312 6948 -8296
rect 6914 -9104 6948 -9088
rect 7044 -8312 7078 -8296
rect 7044 -9104 7078 -9088
rect 7502 -8312 7536 -8296
rect 7502 -9104 7536 -9088
rect 7632 -8312 7666 -8296
rect 7632 -9104 7666 -9088
rect 8090 -8312 8124 -8296
rect 8090 -9104 8124 -9088
rect 8220 -8312 8254 -8296
rect 8220 -9104 8254 -9088
rect 8678 -8312 8712 -8296
rect 8678 -9104 8712 -9088
rect 8808 -8312 8842 -8296
rect 8808 -9104 8842 -9088
rect 9266 -8312 9300 -8296
rect 9266 -9104 9300 -9088
rect 9396 -8312 9430 -8296
rect 9396 -9104 9430 -9088
rect 9854 -8312 9888 -8296
rect 9854 -9104 9888 -9088
rect 9984 -8312 10018 -8296
rect 9984 -9104 10018 -9088
rect 10442 -8312 10476 -8296
rect 10442 -9104 10476 -9088
rect 10572 -8312 10606 -8296
rect 10572 -9104 10606 -9088
rect 11030 -8312 11064 -8296
rect 11030 -9104 11064 -9088
rect 11160 -8312 11194 -8296
rect 11160 -9104 11194 -9088
rect 11618 -8312 11652 -8296
rect 11618 -9104 11652 -9088
rect 11748 -8312 11782 -8296
rect 11748 -9104 11782 -9088
rect 12206 -8312 12240 -8296
rect 12206 -9104 12240 -9088
rect -15842 -9147 -4082 -9146
rect -3682 -9147 -3494 -9146
rect -3094 -9147 -2906 -9146
rect -2506 -9147 -2318 -9146
rect -1918 -9147 -1730 -9146
rect -1330 -9147 -1142 -9146
rect -742 -9147 -554 -9146
rect -154 -9147 34 -9146
rect 434 -9147 12194 -9146
rect -15842 -9181 -15826 -9147
rect -15458 -9181 -15238 -9147
rect -14870 -9181 -14650 -9147
rect -14282 -9181 -14062 -9147
rect -13694 -9181 -13474 -9147
rect -13106 -9181 -12886 -9147
rect -12518 -9181 -12298 -9147
rect -11930 -9181 -11710 -9147
rect -11342 -9181 -11122 -9147
rect -10754 -9181 -10534 -9147
rect -10166 -9181 -9946 -9147
rect -9578 -9181 -9358 -9147
rect -8990 -9181 -8770 -9147
rect -8402 -9181 -8182 -9147
rect -7814 -9181 -7594 -9147
rect -7226 -9181 -7006 -9147
rect -6638 -9181 -6418 -9147
rect -6050 -9181 -5830 -9147
rect -5462 -9181 -5242 -9147
rect -4874 -9181 -4654 -9147
rect -4286 -9181 -4066 -9147
rect -3698 -9181 -3478 -9147
rect -3110 -9181 -2890 -9147
rect -2522 -9181 -2302 -9147
rect -1934 -9181 -1714 -9147
rect -1346 -9181 -1126 -9147
rect -758 -9181 -538 -9147
rect -170 -9181 50 -9147
rect 418 -9181 638 -9147
rect 1006 -9181 1226 -9147
rect 1594 -9181 1814 -9147
rect 2182 -9181 2402 -9147
rect 2770 -9181 2990 -9147
rect 3358 -9181 3578 -9147
rect 3946 -9181 4166 -9147
rect 4534 -9181 4754 -9147
rect 5122 -9181 5342 -9147
rect 5710 -9181 5930 -9147
rect 6298 -9181 6518 -9147
rect 6886 -9181 7106 -9147
rect 7474 -9181 7694 -9147
rect 8062 -9181 8282 -9147
rect 8650 -9181 8870 -9147
rect 9238 -9181 9458 -9147
rect 9826 -9181 10046 -9147
rect 10414 -9181 10634 -9147
rect 11002 -9181 11222 -9147
rect 11590 -9181 11810 -9147
rect 12178 -9181 12194 -9147
rect -15842 -9219 -4082 -9181
rect -3682 -9219 -3494 -9181
rect -3094 -9182 -2906 -9181
rect -3094 -9219 -2906 -9218
rect -2506 -9219 -2318 -9181
rect -1918 -9219 -1730 -9181
rect -1330 -9219 -1142 -9181
rect -742 -9182 -554 -9181
rect -742 -9219 -554 -9218
rect -154 -9219 34 -9181
rect 434 -9219 12194 -9181
rect -15842 -9253 -15826 -9219
rect -15458 -9253 -15238 -9219
rect -14870 -9253 -14650 -9219
rect -14282 -9253 -14062 -9219
rect -13694 -9253 -13474 -9219
rect -13106 -9253 -12886 -9219
rect -12518 -9253 -12298 -9219
rect -11930 -9253 -11710 -9219
rect -11342 -9253 -11122 -9219
rect -10754 -9253 -10534 -9219
rect -10166 -9253 -9946 -9219
rect -9578 -9253 -9358 -9219
rect -8990 -9253 -8770 -9219
rect -8402 -9253 -8182 -9219
rect -7814 -9253 -7594 -9219
rect -7226 -9253 -7006 -9219
rect -6638 -9253 -6418 -9219
rect -6050 -9253 -5830 -9219
rect -5462 -9253 -5242 -9219
rect -4874 -9253 -4654 -9219
rect -4286 -9253 -4066 -9219
rect -3698 -9253 -3478 -9219
rect -3110 -9253 -2890 -9219
rect -2522 -9253 -2302 -9219
rect -1934 -9253 -1714 -9219
rect -1346 -9253 -1126 -9219
rect -758 -9253 -538 -9219
rect -170 -9253 50 -9219
rect 418 -9253 638 -9219
rect 1006 -9253 1226 -9219
rect 1594 -9253 1814 -9219
rect 2182 -9253 2402 -9219
rect 2770 -9253 2990 -9219
rect 3358 -9253 3578 -9219
rect 3946 -9253 4166 -9219
rect 4534 -9253 4754 -9219
rect 5122 -9253 5342 -9219
rect 5710 -9253 5930 -9219
rect 6298 -9253 6518 -9219
rect 6886 -9253 7106 -9219
rect 7474 -9253 7694 -9219
rect 8062 -9253 8282 -9219
rect 8650 -9253 8870 -9219
rect 9238 -9253 9458 -9219
rect 9826 -9253 10046 -9219
rect 10414 -9253 10634 -9219
rect 11002 -9253 11222 -9219
rect 11590 -9253 11810 -9219
rect 12178 -9253 12194 -9219
rect -15842 -9254 -4082 -9253
rect -3682 -9254 -3494 -9253
rect -3094 -9254 -2906 -9253
rect -2506 -9254 -2318 -9253
rect -1918 -9254 -1730 -9253
rect -1330 -9254 -1142 -9253
rect -742 -9254 -554 -9253
rect -154 -9254 34 -9253
rect 434 -9254 12194 -9253
rect -15888 -9312 -15854 -9296
rect -15888 -10104 -15854 -10088
rect -15430 -9312 -15396 -9296
rect -15430 -10104 -15396 -10088
rect -15300 -9312 -15266 -9296
rect -15300 -10104 -15266 -10088
rect -14842 -9312 -14808 -9296
rect -14842 -10104 -14808 -10088
rect -14712 -9312 -14678 -9296
rect -14712 -10104 -14678 -10088
rect -14254 -9312 -14220 -9296
rect -14254 -10104 -14220 -10088
rect -14124 -9312 -14090 -9296
rect -14124 -10104 -14090 -10088
rect -13666 -9312 -13632 -9296
rect -13666 -10104 -13632 -10088
rect -13536 -9312 -13502 -9296
rect -13536 -10104 -13502 -10088
rect -13078 -9312 -13044 -9296
rect -13078 -10104 -13044 -10088
rect -12948 -9312 -12914 -9296
rect -12948 -10104 -12914 -10088
rect -12490 -9312 -12456 -9296
rect -12490 -10104 -12456 -10088
rect -12360 -9312 -12326 -9296
rect -12360 -10104 -12326 -10088
rect -11902 -9312 -11868 -9296
rect -11902 -10104 -11868 -10088
rect -11772 -9312 -11738 -9296
rect -11772 -10104 -11738 -10088
rect -11314 -9312 -11280 -9296
rect -11314 -10104 -11280 -10088
rect -11184 -9312 -11150 -9296
rect -11184 -10104 -11150 -10088
rect -10726 -9312 -10692 -9296
rect -10726 -10104 -10692 -10088
rect -10596 -9312 -10562 -9296
rect -10596 -10104 -10562 -10088
rect -10138 -9312 -10104 -9296
rect -10138 -10104 -10104 -10088
rect -10008 -9312 -9974 -9296
rect -10008 -10104 -9974 -10088
rect -9550 -9312 -9516 -9296
rect -9550 -10104 -9516 -10088
rect -9420 -9312 -9386 -9296
rect -9420 -10104 -9386 -10088
rect -8962 -9312 -8928 -9296
rect -8962 -10104 -8928 -10088
rect -8832 -9312 -8798 -9296
rect -8832 -10104 -8798 -10088
rect -8374 -9312 -8340 -9296
rect -8374 -10104 -8340 -10088
rect -8244 -9312 -8210 -9296
rect -8244 -10104 -8210 -10088
rect -7786 -9312 -7752 -9296
rect -7786 -10104 -7752 -10088
rect -7656 -9312 -7622 -9296
rect -7656 -10104 -7622 -10088
rect -7198 -9312 -7164 -9296
rect -7198 -10104 -7164 -10088
rect -7068 -9312 -7034 -9296
rect -7068 -10104 -7034 -10088
rect -6610 -9312 -6576 -9296
rect -6610 -10104 -6576 -10088
rect -6480 -9312 -6446 -9296
rect -6480 -10104 -6446 -10088
rect -6022 -9312 -5988 -9296
rect -6022 -10104 -5988 -10088
rect -5892 -9312 -5858 -9296
rect -5892 -10104 -5858 -10088
rect -5434 -9312 -5400 -9296
rect -5434 -10104 -5400 -10088
rect -5304 -9312 -5270 -9296
rect -5304 -10104 -5270 -10088
rect -4846 -9312 -4812 -9296
rect -4846 -10104 -4812 -10088
rect -4716 -9312 -4682 -9296
rect -4716 -10104 -4682 -10088
rect -4258 -9312 -4224 -9296
rect -4258 -10104 -4224 -10088
rect -4128 -9312 -4094 -9254
rect -4128 -10146 -4094 -10088
rect -3670 -9312 -3636 -9296
rect -3670 -10104 -3636 -10088
rect -3540 -9312 -3506 -9296
rect -3540 -10104 -3506 -10088
rect -3082 -9312 -3048 -9296
rect -3082 -10104 -3048 -10088
rect -2952 -9312 -2918 -9296
rect -2952 -10104 -2918 -10088
rect -2494 -9312 -2460 -9296
rect -2494 -10104 -2460 -10088
rect -2364 -9312 -2330 -9296
rect -2364 -10104 -2330 -10088
rect -1906 -9312 -1742 -9254
rect -1872 -10088 -1776 -9312
rect -1906 -10146 -1742 -10088
rect -1318 -9312 -1284 -9296
rect -1318 -10104 -1284 -10088
rect -1188 -9312 -1154 -9296
rect -1188 -10104 -1154 -10088
rect -730 -9312 -696 -9296
rect -730 -10104 -696 -10088
rect -600 -9312 -566 -9296
rect -600 -10104 -566 -10088
rect -142 -9312 -108 -9296
rect -142 -10104 -108 -10088
rect -12 -9312 22 -9296
rect -12 -10104 22 -10088
rect 446 -9312 480 -9254
rect 446 -10146 480 -10088
rect 576 -9312 610 -9296
rect 576 -10104 610 -10088
rect 1034 -9312 1068 -9296
rect 1034 -10104 1068 -10088
rect 1164 -9312 1198 -9296
rect 1164 -10104 1198 -10088
rect 1622 -9312 1656 -9296
rect 1622 -10104 1656 -10088
rect 1752 -9312 1786 -9296
rect 1752 -10104 1786 -10088
rect 2210 -9312 2244 -9296
rect 2210 -10104 2244 -10088
rect 2340 -9312 2374 -9296
rect 2340 -10104 2374 -10088
rect 2798 -9312 2832 -9296
rect 2798 -10104 2832 -10088
rect 2928 -9312 2962 -9296
rect 2928 -10104 2962 -10088
rect 3386 -9312 3420 -9296
rect 3386 -10104 3420 -10088
rect 3516 -9312 3550 -9296
rect 3516 -10104 3550 -10088
rect 3974 -9312 4008 -9296
rect 3974 -10104 4008 -10088
rect 4104 -9312 4138 -9296
rect 4104 -10104 4138 -10088
rect 4562 -9312 4596 -9296
rect 4562 -10104 4596 -10088
rect 4692 -9312 4726 -9296
rect 4692 -10104 4726 -10088
rect 5150 -9312 5184 -9296
rect 5150 -10104 5184 -10088
rect 5280 -9312 5314 -9296
rect 5280 -10104 5314 -10088
rect 5738 -9312 5772 -9296
rect 5738 -10104 5772 -10088
rect 5868 -9312 5902 -9296
rect 5868 -10104 5902 -10088
rect 6326 -9312 6360 -9296
rect 6326 -10104 6360 -10088
rect 6456 -9312 6490 -9296
rect 6456 -10104 6490 -10088
rect 6914 -9312 6948 -9296
rect 6914 -10104 6948 -10088
rect 7044 -9312 7078 -9296
rect 7044 -10104 7078 -10088
rect 7502 -9312 7536 -9296
rect 7502 -10104 7536 -10088
rect 7632 -9312 7666 -9296
rect 7632 -10104 7666 -10088
rect 8090 -9312 8124 -9296
rect 8090 -10104 8124 -10088
rect 8220 -9312 8254 -9296
rect 8220 -10104 8254 -10088
rect 8678 -9312 8712 -9296
rect 8678 -10104 8712 -10088
rect 8808 -9312 8842 -9296
rect 8808 -10104 8842 -10088
rect 9266 -9312 9300 -9296
rect 9266 -10104 9300 -10088
rect 9396 -9312 9430 -9296
rect 9396 -10104 9430 -10088
rect 9854 -9312 9888 -9296
rect 9854 -10104 9888 -10088
rect 9984 -9312 10018 -9296
rect 9984 -10104 10018 -10088
rect 10442 -9312 10476 -9296
rect 10442 -10104 10476 -10088
rect 10572 -9312 10606 -9296
rect 10572 -10104 10606 -10088
rect 11030 -9312 11064 -9296
rect 11030 -10104 11064 -10088
rect 11160 -9312 11194 -9296
rect 11160 -10104 11194 -10088
rect 11618 -9312 11652 -9296
rect 11618 -10104 11652 -10088
rect 11748 -9312 11782 -9296
rect 11748 -10104 11782 -10088
rect 12206 -9312 12240 -9296
rect 12206 -10104 12240 -10088
rect -15842 -10147 -4082 -10146
rect -3682 -10147 -3494 -10146
rect -3094 -10147 -2906 -10146
rect -2506 -10147 -2318 -10146
rect -1918 -10147 -1730 -10146
rect -1330 -10147 -1142 -10146
rect -742 -10147 -554 -10146
rect -154 -10147 34 -10146
rect 434 -10147 12194 -10146
rect -15842 -10181 -15826 -10147
rect -15458 -10181 -15238 -10147
rect -14870 -10181 -14650 -10147
rect -14282 -10181 -14062 -10147
rect -13694 -10181 -13474 -10147
rect -13106 -10181 -12886 -10147
rect -12518 -10181 -12298 -10147
rect -11930 -10181 -11710 -10147
rect -11342 -10181 -11122 -10147
rect -10754 -10181 -10534 -10147
rect -10166 -10181 -9946 -10147
rect -9578 -10181 -9358 -10147
rect -8990 -10181 -8770 -10147
rect -8402 -10181 -8182 -10147
rect -7814 -10181 -7594 -10147
rect -7226 -10181 -7006 -10147
rect -6638 -10181 -6418 -10147
rect -6050 -10181 -5830 -10147
rect -5462 -10181 -5242 -10147
rect -4874 -10181 -4654 -10147
rect -4286 -10181 -4066 -10147
rect -3698 -10181 -3478 -10147
rect -3110 -10181 -2890 -10147
rect -2522 -10181 -2302 -10147
rect -1934 -10181 -1714 -10147
rect -1346 -10181 -1126 -10147
rect -758 -10181 -538 -10147
rect -170 -10181 50 -10147
rect 418 -10181 638 -10147
rect 1006 -10181 1226 -10147
rect 1594 -10181 1814 -10147
rect 2182 -10181 2402 -10147
rect 2770 -10181 2990 -10147
rect 3358 -10181 3578 -10147
rect 3946 -10181 4166 -10147
rect 4534 -10181 4754 -10147
rect 5122 -10181 5342 -10147
rect 5710 -10181 5930 -10147
rect 6298 -10181 6518 -10147
rect 6886 -10181 7106 -10147
rect 7474 -10181 7694 -10147
rect 8062 -10181 8282 -10147
rect 8650 -10181 8870 -10147
rect 9238 -10181 9458 -10147
rect 9826 -10181 10046 -10147
rect 10414 -10181 10634 -10147
rect 11002 -10181 11222 -10147
rect 11590 -10181 11810 -10147
rect 12178 -10181 12194 -10147
rect -15842 -10219 -4082 -10181
rect -3682 -10219 -3494 -10181
rect -3094 -10182 -2906 -10181
rect -3094 -10219 -2906 -10218
rect -2506 -10219 -2318 -10181
rect -1918 -10219 -1730 -10181
rect -1330 -10219 -1142 -10181
rect -742 -10182 -554 -10181
rect -742 -10219 -554 -10218
rect -154 -10219 34 -10181
rect 434 -10219 12194 -10181
rect -15842 -10253 -15826 -10219
rect -15458 -10253 -15238 -10219
rect -14870 -10253 -14650 -10219
rect -14282 -10253 -14062 -10219
rect -13694 -10253 -13474 -10219
rect -13106 -10253 -12886 -10219
rect -12518 -10253 -12298 -10219
rect -11930 -10253 -11710 -10219
rect -11342 -10253 -11122 -10219
rect -10754 -10253 -10534 -10219
rect -10166 -10253 -9946 -10219
rect -9578 -10253 -9358 -10219
rect -8990 -10253 -8770 -10219
rect -8402 -10253 -8182 -10219
rect -7814 -10253 -7594 -10219
rect -7226 -10253 -7006 -10219
rect -6638 -10253 -6418 -10219
rect -6050 -10253 -5830 -10219
rect -5462 -10253 -5242 -10219
rect -4874 -10253 -4654 -10219
rect -4286 -10253 -4066 -10219
rect -3698 -10253 -3478 -10219
rect -3110 -10253 -2890 -10219
rect -2522 -10253 -2302 -10219
rect -1934 -10253 -1714 -10219
rect -1346 -10253 -1126 -10219
rect -758 -10253 -538 -10219
rect -170 -10253 50 -10219
rect 418 -10253 638 -10219
rect 1006 -10253 1226 -10219
rect 1594 -10253 1814 -10219
rect 2182 -10253 2402 -10219
rect 2770 -10253 2990 -10219
rect 3358 -10253 3578 -10219
rect 3946 -10253 4166 -10219
rect 4534 -10253 4754 -10219
rect 5122 -10253 5342 -10219
rect 5710 -10253 5930 -10219
rect 6298 -10253 6518 -10219
rect 6886 -10253 7106 -10219
rect 7474 -10253 7694 -10219
rect 8062 -10253 8282 -10219
rect 8650 -10253 8870 -10219
rect 9238 -10253 9458 -10219
rect 9826 -10253 10046 -10219
rect 10414 -10253 10634 -10219
rect 11002 -10253 11222 -10219
rect 11590 -10253 11810 -10219
rect 12178 -10253 12194 -10219
rect -15842 -10254 -4082 -10253
rect -3682 -10254 -3494 -10253
rect -3094 -10254 -2906 -10253
rect -2506 -10254 -2318 -10253
rect -1918 -10254 -1730 -10253
rect -1330 -10254 -1142 -10253
rect -742 -10254 -554 -10253
rect -154 -10254 34 -10253
rect 434 -10254 12194 -10253
rect -15888 -10312 -15854 -10296
rect -15888 -11104 -15854 -11088
rect -15430 -10312 -15396 -10296
rect -15430 -11104 -15396 -11088
rect -15300 -10312 -15266 -10296
rect -15300 -11104 -15266 -11088
rect -14842 -10312 -14808 -10296
rect -14842 -11104 -14808 -11088
rect -14712 -10312 -14678 -10296
rect -14712 -11104 -14678 -11088
rect -14254 -10312 -14220 -10296
rect -14254 -11104 -14220 -11088
rect -14124 -10312 -14090 -10296
rect -14124 -11104 -14090 -11088
rect -13666 -10312 -13632 -10296
rect -13666 -11104 -13632 -11088
rect -13536 -10312 -13502 -10296
rect -13536 -11104 -13502 -11088
rect -13078 -10312 -13044 -10296
rect -13078 -11104 -13044 -11088
rect -12948 -10312 -12914 -10296
rect -12948 -11104 -12914 -11088
rect -12490 -10312 -12456 -10296
rect -12490 -11104 -12456 -11088
rect -12360 -10312 -12326 -10296
rect -12360 -11104 -12326 -11088
rect -11902 -10312 -11868 -10296
rect -11902 -11104 -11868 -11088
rect -11772 -10312 -11738 -10296
rect -11772 -11104 -11738 -11088
rect -11314 -10312 -11280 -10296
rect -11314 -11104 -11280 -11088
rect -11184 -10312 -11150 -10296
rect -11184 -11104 -11150 -11088
rect -10726 -10312 -10692 -10296
rect -10726 -11104 -10692 -11088
rect -10596 -10312 -10562 -10296
rect -10596 -11104 -10562 -11088
rect -10138 -10312 -10104 -10296
rect -10138 -11104 -10104 -11088
rect -10008 -10312 -9974 -10296
rect -10008 -11104 -9974 -11088
rect -9550 -10312 -9516 -10296
rect -9550 -11104 -9516 -11088
rect -9420 -10312 -9386 -10296
rect -9420 -11104 -9386 -11088
rect -8962 -10312 -8928 -10296
rect -8962 -11104 -8928 -11088
rect -8832 -10312 -8798 -10296
rect -8832 -11104 -8798 -11088
rect -8374 -10312 -8340 -10296
rect -8374 -11104 -8340 -11088
rect -8244 -10312 -8210 -10296
rect -8244 -11104 -8210 -11088
rect -7786 -10312 -7752 -10296
rect -7786 -11104 -7752 -11088
rect -7656 -10312 -7622 -10296
rect -7656 -11104 -7622 -11088
rect -7198 -10312 -7164 -10296
rect -7198 -11104 -7164 -11088
rect -7068 -10312 -7034 -10296
rect -7068 -11104 -7034 -11088
rect -6610 -10312 -6576 -10296
rect -6610 -11104 -6576 -11088
rect -6480 -10312 -6446 -10296
rect -6480 -11104 -6446 -11088
rect -6022 -10312 -5988 -10296
rect -6022 -11104 -5988 -11088
rect -5892 -10312 -5858 -10296
rect -5892 -11104 -5858 -11088
rect -5434 -10312 -5400 -10296
rect -5434 -11104 -5400 -11088
rect -5304 -10312 -5270 -10296
rect -5304 -11104 -5270 -11088
rect -4846 -10312 -4812 -10296
rect -4846 -11104 -4812 -11088
rect -4716 -10312 -4682 -10296
rect -4716 -11104 -4682 -11088
rect -4258 -10312 -4224 -10296
rect -4258 -11104 -4224 -11088
rect -4128 -10312 -4094 -10254
rect -4128 -11104 -4094 -11088
rect -3670 -10312 -3636 -10296
rect -3670 -11104 -3636 -11088
rect -3540 -10312 -3506 -10296
rect -3540 -11104 -3506 -11088
rect -3082 -10312 -3048 -10296
rect -3082 -11104 -3048 -11088
rect -2952 -10312 -2918 -10296
rect -2952 -11104 -2918 -11088
rect -2494 -10312 -2460 -10296
rect -2494 -11104 -2460 -11088
rect -2364 -10312 -2330 -10296
rect -2364 -11104 -2330 -11088
rect -1906 -10312 -1742 -10254
rect -1872 -11088 -1776 -10312
rect -1906 -11104 -1742 -11088
rect -1318 -10312 -1284 -10296
rect -1318 -11104 -1284 -11088
rect -1188 -10312 -1154 -10296
rect -1188 -11104 -1154 -11088
rect -730 -10312 -696 -10296
rect -730 -11104 -696 -11088
rect -600 -10312 -566 -10296
rect -600 -11104 -566 -11088
rect -142 -10312 -108 -10296
rect -142 -11104 -108 -11088
rect -12 -10312 22 -10296
rect -12 -11104 22 -11088
rect 446 -10312 480 -10254
rect 446 -11104 480 -11088
rect 576 -10312 610 -10296
rect 576 -11104 610 -11088
rect 1034 -10312 1068 -10296
rect 1034 -11104 1068 -11088
rect 1164 -10312 1198 -10296
rect 1164 -11104 1198 -11088
rect 1622 -10312 1656 -10296
rect 1622 -11104 1656 -11088
rect 1752 -10312 1786 -10296
rect 1752 -11104 1786 -11088
rect 2210 -10312 2244 -10296
rect 2210 -11104 2244 -11088
rect 2340 -10312 2374 -10296
rect 2340 -11104 2374 -11088
rect 2798 -10312 2832 -10296
rect 2798 -11104 2832 -11088
rect 2928 -10312 2962 -10296
rect 2928 -11104 2962 -11088
rect 3386 -10312 3420 -10296
rect 3386 -11104 3420 -11088
rect 3516 -10312 3550 -10296
rect 3516 -11104 3550 -11088
rect 3974 -10312 4008 -10296
rect 3974 -11104 4008 -11088
rect 4104 -10312 4138 -10296
rect 4104 -11104 4138 -11088
rect 4562 -10312 4596 -10296
rect 4562 -11104 4596 -11088
rect 4692 -10312 4726 -10296
rect 4692 -11104 4726 -11088
rect 5150 -10312 5184 -10296
rect 5150 -11104 5184 -11088
rect 5280 -10312 5314 -10296
rect 5280 -11104 5314 -11088
rect 5738 -10312 5772 -10296
rect 5738 -11104 5772 -11088
rect 5868 -10312 5902 -10296
rect 5868 -11104 5902 -11088
rect 6326 -10312 6360 -10296
rect 6326 -11104 6360 -11088
rect 6456 -10312 6490 -10296
rect 6456 -11104 6490 -11088
rect 6914 -10312 6948 -10296
rect 6914 -11104 6948 -11088
rect 7044 -10312 7078 -10296
rect 7044 -11104 7078 -11088
rect 7502 -10312 7536 -10296
rect 7502 -11104 7536 -11088
rect 7632 -10312 7666 -10296
rect 7632 -11104 7666 -11088
rect 8090 -10312 8124 -10296
rect 8090 -11104 8124 -11088
rect 8220 -10312 8254 -10296
rect 8220 -11104 8254 -11088
rect 8678 -10312 8712 -10296
rect 8678 -11104 8712 -11088
rect 8808 -10312 8842 -10296
rect 8808 -11104 8842 -11088
rect 9266 -10312 9300 -10296
rect 9266 -11104 9300 -11088
rect 9396 -10312 9430 -10296
rect 9396 -11104 9430 -11088
rect 9854 -10312 9888 -10296
rect 9854 -11104 9888 -11088
rect 9984 -10312 10018 -10296
rect 9984 -11104 10018 -11088
rect 10442 -10312 10476 -10296
rect 10442 -11104 10476 -11088
rect 10572 -10312 10606 -10296
rect 10572 -11104 10606 -11088
rect 11030 -10312 11064 -10296
rect 11030 -11104 11064 -11088
rect 11160 -10312 11194 -10296
rect 11160 -11104 11194 -11088
rect 11618 -10312 11652 -10296
rect 11618 -11104 11652 -11088
rect 11748 -10312 11782 -10296
rect 11748 -11104 11782 -11088
rect 12206 -10312 12240 -10296
rect 12206 -11104 12240 -11088
rect -4128 -11146 -4082 -11104
rect -15842 -11147 -4082 -11146
rect -3682 -11147 -3494 -11146
rect -3094 -11147 -2906 -11146
rect -2506 -11147 -2318 -11146
rect -1918 -11147 -1730 -11104
rect 434 -11146 480 -11104
rect -1330 -11147 -1142 -11146
rect -742 -11147 -554 -11146
rect -154 -11147 34 -11146
rect 434 -11147 12194 -11146
rect -15842 -11181 -15826 -11147
rect -15458 -11181 -15238 -11147
rect -14870 -11181 -14650 -11147
rect -14282 -11181 -14062 -11147
rect -13694 -11181 -13474 -11147
rect -13106 -11181 -12886 -11147
rect -12518 -11181 -12298 -11147
rect -11930 -11181 -11710 -11147
rect -11342 -11181 -11122 -11147
rect -10754 -11181 -10534 -11147
rect -10166 -11181 -9946 -11147
rect -9578 -11181 -9358 -11147
rect -8990 -11181 -8770 -11147
rect -8402 -11181 -8182 -11147
rect -7814 -11181 -7594 -11147
rect -7226 -11181 -7006 -11147
rect -6638 -11181 -6418 -11147
rect -6050 -11181 -5830 -11147
rect -5462 -11181 -5242 -11147
rect -4874 -11181 -4654 -11147
rect -4286 -11181 -4066 -11147
rect -3698 -11181 -3478 -11147
rect -3110 -11181 -2890 -11147
rect -2522 -11181 -2302 -11147
rect -1934 -11181 -1714 -11147
rect -1346 -11181 -1126 -11147
rect -758 -11181 -538 -11147
rect -170 -11181 50 -11147
rect 418 -11181 638 -11147
rect 1006 -11181 1226 -11147
rect 1594 -11181 1814 -11147
rect 2182 -11181 2402 -11147
rect 2770 -11181 2990 -11147
rect 3358 -11181 3578 -11147
rect 3946 -11181 4166 -11147
rect 4534 -11181 4754 -11147
rect 5122 -11181 5342 -11147
rect 5710 -11181 5930 -11147
rect 6298 -11181 6518 -11147
rect 6886 -11181 7106 -11147
rect 7474 -11181 7694 -11147
rect 8062 -11181 8282 -11147
rect 8650 -11181 8870 -11147
rect 9238 -11181 9458 -11147
rect 9826 -11181 10046 -11147
rect 10414 -11181 10634 -11147
rect 11002 -11181 11222 -11147
rect 11590 -11181 11810 -11147
rect 12178 -11181 12194 -11147
rect -15842 -11182 -4082 -11181
rect -3682 -11182 -3494 -11181
rect -3094 -11182 -2906 -11181
rect -2506 -11182 -2318 -11181
rect -1918 -11182 -1730 -11181
rect -1330 -11182 -1142 -11181
rect -742 -11182 -554 -11181
rect -154 -11182 34 -11181
rect 434 -11182 12194 -11181
rect -16234 -11498 -16200 -11478
rect 12552 -11498 12586 -11444
rect -16234 -11532 -16116 -11498
rect 12498 -11532 12586 -11498
rect -2532 -11560 -2506 -11532
rect -2318 -11560 -2288 -11532
rect -2532 -12242 -2288 -11560
rect -1358 -11560 -1330 -11532
rect -1142 -11560 -1114 -11532
rect -1358 -12242 -1114 -11560
rect -3222 -12276 -3188 -12242
rect -460 -12276 -426 -12242
rect -2790 -12708 -2774 -12576
rect -2736 -12708 -2508 -12576
rect -2470 -12708 -2452 -12576
rect -2258 -12708 -2242 -12576
rect -2204 -12708 -1976 -12576
rect -1938 -12708 -1920 -12576
rect -1726 -12708 -1710 -12576
rect -1672 -12708 -1444 -12576
rect -1406 -12708 -1388 -12576
rect -1194 -12708 -1178 -12576
rect -1140 -12708 -912 -12576
rect -874 -12708 -856 -12576
rect -2836 -12758 -2802 -12742
rect -2836 -13550 -2802 -13534
rect -2708 -12758 -2674 -12742
rect -2708 -13550 -2674 -13534
rect -2570 -12758 -2536 -12742
rect -2570 -13550 -2536 -13534
rect -2442 -12758 -2408 -12742
rect -2442 -13550 -2408 -13534
rect -2304 -12758 -2270 -12742
rect -2304 -13550 -2270 -13534
rect -2176 -12758 -2142 -12742
rect -2176 -13550 -2142 -13534
rect -2038 -12758 -2004 -12742
rect -2038 -13550 -2004 -13534
rect -1910 -12758 -1876 -12742
rect -1910 -13550 -1876 -13534
rect -1772 -12758 -1738 -12742
rect -1772 -13550 -1738 -13534
rect -1644 -12758 -1610 -12742
rect -1644 -13550 -1610 -13534
rect -1506 -12758 -1472 -12742
rect -1506 -13550 -1472 -13534
rect -1378 -12758 -1344 -12742
rect -1378 -13550 -1344 -13534
rect -1240 -12758 -1206 -12742
rect -1240 -13550 -1206 -13534
rect -1112 -12758 -1078 -12742
rect -1112 -13550 -1078 -13534
rect -974 -12758 -940 -12742
rect -974 -13550 -940 -13534
rect -846 -12758 -812 -12742
rect -846 -13550 -812 -13534
rect -2790 -13718 -2774 -13586
rect -2736 -13718 -2508 -13586
rect -2470 -13718 -2452 -13586
rect -2258 -13718 -2242 -13586
rect -2204 -13718 -1976 -13586
rect -1938 -13718 -1920 -13586
rect -1726 -13718 -1710 -13586
rect -1672 -13718 -1444 -13586
rect -1406 -13718 -1388 -13586
rect -1194 -13718 -1178 -13586
rect -1140 -13718 -912 -13586
rect -874 -13718 -856 -13586
rect -2836 -13768 -2802 -13752
rect -2836 -14560 -2802 -14544
rect -2708 -13768 -2674 -13752
rect -2708 -14560 -2674 -14544
rect -2570 -13768 -2536 -13752
rect -2570 -14560 -2536 -14544
rect -2442 -13768 -2408 -13752
rect -2442 -14560 -2408 -14544
rect -2304 -13768 -2270 -13752
rect -2304 -14560 -2270 -14544
rect -2176 -13768 -2142 -13752
rect -2176 -14560 -2142 -14544
rect -2038 -13768 -2004 -13752
rect -2038 -14560 -2004 -14544
rect -1910 -13768 -1876 -13752
rect -1910 -14560 -1876 -14544
rect -1772 -13768 -1738 -13752
rect -1772 -14560 -1738 -14544
rect -1644 -13768 -1610 -13752
rect -1644 -14560 -1610 -14544
rect -1506 -13768 -1472 -13752
rect -1506 -14560 -1472 -14544
rect -1378 -13768 -1344 -13752
rect -1378 -14560 -1344 -14544
rect -1240 -13768 -1206 -13752
rect -1240 -14560 -1206 -14544
rect -1112 -13768 -1078 -13752
rect -1112 -14560 -1078 -14544
rect -974 -13768 -940 -13752
rect -974 -14560 -940 -14544
rect -846 -13768 -812 -13752
rect -846 -14560 -812 -14544
rect -2790 -14728 -2774 -14596
rect -2736 -14728 -2508 -14596
rect -2470 -14728 -2452 -14596
rect -2258 -14728 -2242 -14596
rect -2204 -14728 -1976 -14596
rect -1938 -14728 -1920 -14596
rect -1726 -14728 -1710 -14596
rect -1672 -14728 -1444 -14596
rect -1406 -14728 -1388 -14596
rect -1194 -14728 -1178 -14596
rect -1140 -14728 -912 -14596
rect -874 -14728 -856 -14596
rect -2836 -14778 -2802 -14762
rect -2836 -15570 -2802 -15554
rect -2708 -14778 -2674 -14762
rect -2708 -15570 -2674 -15554
rect -2570 -14778 -2536 -14762
rect -2570 -15570 -2536 -15554
rect -2442 -14778 -2408 -14762
rect -2442 -15570 -2408 -15554
rect -2304 -14778 -2270 -14762
rect -2304 -15570 -2270 -15554
rect -2176 -14778 -2142 -14762
rect -2176 -15570 -2142 -15554
rect -2038 -14778 -2004 -14762
rect -2038 -15570 -2004 -15554
rect -1910 -14778 -1876 -14762
rect -1910 -15570 -1876 -15554
rect -1772 -14778 -1738 -14762
rect -1772 -15570 -1738 -15554
rect -1644 -14778 -1610 -14762
rect -1644 -15570 -1610 -15554
rect -1506 -14778 -1472 -14762
rect -1506 -15570 -1472 -15554
rect -1378 -14778 -1344 -14762
rect -1378 -15570 -1344 -15554
rect -1240 -14778 -1206 -14762
rect -1240 -15570 -1206 -15554
rect -1112 -14778 -1078 -14762
rect -1112 -15570 -1078 -15554
rect -974 -14778 -940 -14762
rect -974 -15570 -940 -15554
rect -846 -14778 -812 -14762
rect -846 -15570 -812 -15554
rect -2790 -15738 -2774 -15606
rect -2736 -15738 -2508 -15606
rect -2470 -15738 -2452 -15606
rect -2258 -15738 -2242 -15606
rect -2204 -15738 -1976 -15606
rect -1938 -15738 -1920 -15606
rect -1726 -15738 -1710 -15606
rect -1672 -15738 -1444 -15606
rect -1406 -15738 -1388 -15606
rect -1194 -15738 -1178 -15606
rect -1140 -15738 -912 -15606
rect -874 -15738 -856 -15606
rect -3222 -16072 -3188 -16038
rect -460 -16072 -426 -16038
rect 4237 -14883 4333 -14849
rect 4471 -14858 4567 -14849
rect 4471 -14878 4792 -14858
rect 4471 -14883 4634 -14878
rect 4237 -14945 4271 -14883
rect 4533 -14945 4634 -14883
rect 4237 -16039 4271 -15977
rect 4567 -15338 4634 -14945
rect 4774 -15338 4792 -14878
rect 4567 -15360 4792 -15338
rect 4533 -16039 4567 -15977
rect 4237 -16073 4333 -16039
rect 4471 -16073 4567 -16039
rect -2610 -16468 -2464 -16434
rect -1254 -16468 -1036 -16434
rect -2264 -16774 -1382 -16768
rect -2264 -16900 -2202 -16774
rect -2164 -16900 -1962 -16774
rect -1924 -16900 -1722 -16774
rect -1684 -16900 -1482 -16774
rect -1444 -16900 -1382 -16774
rect -2264 -16950 -2230 -16900
rect -2264 -17576 -2230 -17526
rect -2136 -16950 -2102 -16934
rect -2136 -17542 -2102 -17526
rect -2024 -16950 -1990 -16934
rect -2024 -17542 -1990 -17526
rect -1896 -16950 -1862 -16934
rect -1896 -17542 -1862 -17526
rect -1784 -16950 -1750 -16934
rect -1784 -17542 -1750 -17526
rect -1656 -16950 -1622 -16934
rect -1656 -17542 -1622 -17526
rect -1544 -16950 -1510 -16934
rect -1544 -17542 -1510 -17526
rect -1416 -16950 -1382 -16900
rect -1416 -17576 -1382 -17526
rect -2264 -17708 -2202 -17576
rect -2164 -17708 -1962 -17576
rect -1924 -17708 -1722 -17576
rect -1684 -17708 -1482 -17576
rect -1444 -17708 -1382 -17576
rect -2264 -17758 -2230 -17708
rect -2264 -18384 -2230 -18334
rect -2136 -17758 -2102 -17742
rect -2136 -18350 -2102 -18334
rect -2024 -17758 -1990 -17742
rect -2024 -18350 -1990 -18334
rect -1896 -17758 -1862 -17742
rect -1896 -18350 -1862 -18334
rect -1784 -17758 -1750 -17742
rect -1784 -18350 -1750 -18334
rect -1656 -17758 -1622 -17742
rect -1656 -18350 -1622 -18334
rect -1544 -17758 -1510 -17742
rect -1544 -18350 -1510 -18334
rect -1416 -17758 -1382 -17708
rect -1416 -18384 -1382 -18334
rect -2264 -18516 -2202 -18384
rect -2164 -18516 -1962 -18384
rect -1924 -18516 -1722 -18384
rect -1684 -18516 -1482 -18384
rect -1444 -18516 -1382 -18384
rect -2610 -18850 -2512 -18816
rect -1160 -18850 -1036 -18816
<< viali >>
rect -6438 -3746 -6328 -3712
rect -5958 -3746 -5848 -3712
rect -5478 -3746 -5368 -3712
rect -4998 -3746 -4888 -3712
rect -4518 -3746 -4408 -3712
rect -4038 -3746 -3928 -3712
rect -3558 -3746 -3448 -3712
rect -3078 -3746 -2968 -3712
rect -2598 -3746 -2488 -3712
rect -2118 -3746 -2008 -3712
rect -1638 -3746 -1528 -3712
rect -1158 -3746 -1048 -3712
rect -678 -3746 -568 -3712
rect -198 -3746 -88 -3712
rect 282 -3746 392 -3712
rect 762 -3746 872 -3712
rect 1242 -3746 1352 -3712
rect 1722 -3746 1832 -3712
rect 2202 -3746 2312 -3712
rect 2682 -3746 2792 -3712
rect -6438 -3784 -6328 -3746
rect -5958 -3784 -5848 -3746
rect -5478 -3784 -5368 -3746
rect -4998 -3784 -4888 -3746
rect -4518 -3784 -4408 -3746
rect -4038 -3784 -3928 -3746
rect -3558 -3784 -3448 -3746
rect -3078 -3784 -2968 -3746
rect -2598 -3784 -2488 -3746
rect -2118 -3784 -2008 -3746
rect -1638 -3784 -1528 -3746
rect -1158 -3784 -1048 -3746
rect -678 -3784 -568 -3746
rect -198 -3784 -88 -3746
rect 282 -3784 392 -3746
rect 762 -3784 872 -3746
rect 1242 -3784 1352 -3746
rect 1722 -3784 1832 -3746
rect 2202 -3784 2312 -3746
rect 2682 -3784 2792 -3746
rect -6522 -4188 -6484 -4056
rect -6282 -4188 -6244 -4056
rect -6042 -4188 -6004 -4056
rect -5802 -4188 -5764 -4056
rect -5562 -4188 -5524 -4056
rect -5322 -4188 -5284 -4056
rect -5082 -4188 -5044 -4056
rect -4842 -4188 -4804 -4056
rect -4602 -4188 -4564 -4056
rect -4362 -4188 -4324 -4056
rect -4122 -4188 -4084 -4056
rect -3882 -4188 -3844 -4056
rect -3642 -4188 -3604 -4056
rect -3402 -4188 -3364 -4056
rect -3162 -4188 -3124 -4056
rect -2922 -4188 -2884 -4056
rect -2682 -4188 -2644 -4056
rect -2442 -4188 -2404 -4056
rect -2202 -4188 -2164 -4056
rect -1962 -4188 -1924 -4056
rect -1722 -4188 -1684 -4056
rect -1482 -4188 -1444 -4056
rect -1242 -4188 -1204 -4056
rect -1002 -4188 -964 -4056
rect -762 -4188 -724 -4056
rect -522 -4188 -484 -4056
rect -282 -4188 -244 -4056
rect -42 -4188 -4 -4056
rect 198 -4188 236 -4056
rect 438 -4188 476 -4056
rect 678 -4188 716 -4056
rect 918 -4188 956 -4056
rect 1158 -4188 1196 -4056
rect 1398 -4188 1436 -4056
rect 1638 -4188 1676 -4056
rect 1878 -4188 1916 -4056
rect 2118 -4188 2156 -4056
rect 2358 -4188 2396 -4056
rect 2598 -4188 2636 -4056
rect 2838 -4188 2876 -4056
rect -6584 -4814 -6550 -4238
rect -6456 -4814 -6422 -4238
rect -6344 -4814 -6310 -4238
rect -6216 -4814 -6182 -4238
rect -6104 -4814 -6070 -4238
rect -5976 -4814 -5942 -4238
rect -5864 -4814 -5830 -4238
rect -5736 -4814 -5702 -4238
rect -5624 -4814 -5590 -4238
rect -5496 -4814 -5462 -4238
rect -5384 -4814 -5350 -4238
rect -5256 -4814 -5222 -4238
rect -5144 -4814 -5110 -4238
rect -5016 -4814 -4982 -4238
rect -4904 -4814 -4870 -4238
rect -4776 -4814 -4742 -4238
rect -4664 -4814 -4630 -4238
rect -4536 -4814 -4502 -4238
rect -4424 -4814 -4390 -4238
rect -4296 -4814 -4262 -4238
rect -4184 -4814 -4150 -4238
rect -4056 -4814 -4022 -4238
rect -3944 -4814 -3910 -4238
rect -3816 -4814 -3782 -4238
rect -3704 -4814 -3670 -4238
rect -3576 -4814 -3542 -4238
rect -3464 -4814 -3430 -4238
rect -3336 -4814 -3302 -4238
rect -3224 -4814 -3190 -4238
rect -3096 -4814 -3062 -4238
rect -2984 -4814 -2950 -4238
rect -2856 -4814 -2822 -4238
rect -2744 -4814 -2710 -4238
rect -2616 -4814 -2582 -4238
rect -2504 -4814 -2470 -4238
rect -2376 -4814 -2342 -4238
rect -2264 -4814 -2230 -4238
rect -2136 -4814 -2102 -4238
rect -2024 -4814 -1990 -4238
rect -1896 -4814 -1862 -4238
rect -1784 -4814 -1750 -4238
rect -1656 -4814 -1622 -4238
rect -1544 -4814 -1510 -4238
rect -1416 -4814 -1382 -4238
rect -1304 -4814 -1270 -4238
rect -1176 -4814 -1142 -4238
rect -1064 -4814 -1030 -4238
rect -936 -4814 -902 -4238
rect -824 -4814 -790 -4238
rect -696 -4814 -662 -4238
rect -584 -4814 -550 -4238
rect -456 -4814 -422 -4238
rect -344 -4814 -310 -4238
rect -216 -4814 -182 -4238
rect -104 -4814 -70 -4238
rect 24 -4814 58 -4238
rect 136 -4814 170 -4238
rect 264 -4814 298 -4238
rect 376 -4814 410 -4238
rect 504 -4814 538 -4238
rect 616 -4814 650 -4238
rect 744 -4814 778 -4238
rect 856 -4814 890 -4238
rect 984 -4814 1018 -4238
rect 1096 -4814 1130 -4238
rect 1224 -4814 1258 -4238
rect 1336 -4814 1370 -4238
rect 1464 -4814 1498 -4238
rect 1576 -4814 1610 -4238
rect 1704 -4814 1738 -4238
rect 1816 -4814 1850 -4238
rect 1944 -4814 1978 -4238
rect 2056 -4814 2090 -4238
rect 2184 -4814 2218 -4238
rect 2296 -4814 2330 -4238
rect 2424 -4814 2458 -4238
rect 2536 -4814 2570 -4238
rect 2664 -4814 2698 -4238
rect 2776 -4814 2810 -4238
rect 2904 -4814 2938 -4238
rect -6522 -4996 -6484 -4864
rect -6282 -4996 -6244 -4864
rect -6042 -4996 -6004 -4864
rect -5802 -4996 -5764 -4864
rect -5562 -4996 -5524 -4864
rect -5322 -4996 -5284 -4864
rect -5082 -4996 -5044 -4864
rect -4842 -4996 -4804 -4864
rect -4602 -4996 -4564 -4864
rect -4362 -4996 -4324 -4864
rect -4122 -4996 -4084 -4864
rect -3882 -4996 -3844 -4864
rect -3642 -4996 -3604 -4864
rect -3402 -4996 -3364 -4864
rect -3162 -4996 -3124 -4864
rect -2922 -4996 -2884 -4864
rect -2682 -4996 -2644 -4864
rect -2442 -4996 -2404 -4864
rect -2202 -4996 -2164 -4864
rect -1962 -4996 -1924 -4864
rect -1722 -4996 -1684 -4864
rect -1482 -4996 -1444 -4864
rect -1242 -4996 -1204 -4864
rect -1002 -4996 -964 -4864
rect -762 -4996 -724 -4864
rect -522 -4996 -484 -4864
rect -282 -4996 -244 -4864
rect -42 -4996 -4 -4864
rect 198 -4996 236 -4864
rect 438 -4996 476 -4864
rect 678 -4996 716 -4864
rect 918 -4996 956 -4864
rect 1158 -4996 1196 -4864
rect 1398 -4996 1436 -4864
rect 1638 -4996 1676 -4864
rect 1878 -4996 1916 -4864
rect 2118 -4996 2156 -4864
rect 2358 -4996 2396 -4864
rect 2598 -4996 2636 -4864
rect 2838 -4996 2876 -4864
rect -6584 -5622 -6550 -5046
rect -6456 -5622 -6422 -5046
rect -6344 -5622 -6310 -5046
rect -6216 -5622 -6182 -5046
rect -6104 -5622 -6070 -5046
rect -5976 -5622 -5942 -5046
rect -5864 -5622 -5830 -5046
rect -5736 -5622 -5702 -5046
rect -5624 -5622 -5590 -5046
rect -5496 -5622 -5462 -5046
rect -5384 -5622 -5350 -5046
rect -5256 -5622 -5222 -5046
rect -5144 -5622 -5110 -5046
rect -5016 -5622 -4982 -5046
rect -4904 -5622 -4870 -5046
rect -4776 -5622 -4742 -5046
rect -4664 -5622 -4630 -5046
rect -4536 -5622 -4502 -5046
rect -4424 -5622 -4390 -5046
rect -4296 -5622 -4262 -5046
rect -4184 -5622 -4150 -5046
rect -4056 -5622 -4022 -5046
rect -3944 -5622 -3910 -5046
rect -3816 -5622 -3782 -5046
rect -3704 -5622 -3670 -5046
rect -3576 -5622 -3542 -5046
rect -3464 -5622 -3430 -5046
rect -3336 -5622 -3302 -5046
rect -3224 -5622 -3190 -5046
rect -3096 -5622 -3062 -5046
rect -2984 -5622 -2950 -5046
rect -2856 -5622 -2822 -5046
rect -2744 -5622 -2710 -5046
rect -2616 -5622 -2582 -5046
rect -2504 -5622 -2470 -5046
rect -2376 -5622 -2342 -5046
rect -2264 -5622 -2230 -5046
rect -2136 -5622 -2102 -5046
rect -2024 -5622 -1990 -5046
rect -1896 -5622 -1862 -5046
rect -1784 -5622 -1750 -5046
rect -1656 -5622 -1622 -5046
rect -1544 -5622 -1510 -5046
rect -1416 -5622 -1382 -5046
rect -1304 -5622 -1270 -5046
rect -1176 -5622 -1142 -5046
rect -1064 -5622 -1030 -5046
rect -936 -5622 -902 -5046
rect -824 -5622 -790 -5046
rect -696 -5622 -662 -5046
rect -584 -5622 -550 -5046
rect -456 -5622 -422 -5046
rect -344 -5622 -310 -5046
rect -216 -5622 -182 -5046
rect -104 -5622 -70 -5046
rect 24 -5622 58 -5046
rect 136 -5622 170 -5046
rect 264 -5622 298 -5046
rect 376 -5622 410 -5046
rect 504 -5622 538 -5046
rect 616 -5622 650 -5046
rect 744 -5622 778 -5046
rect 856 -5622 890 -5046
rect 984 -5622 1018 -5046
rect 1096 -5622 1130 -5046
rect 1224 -5622 1258 -5046
rect 1336 -5622 1370 -5046
rect 1464 -5622 1498 -5046
rect 1576 -5622 1610 -5046
rect 1704 -5622 1738 -5046
rect 1816 -5622 1850 -5046
rect 1944 -5622 1978 -5046
rect 2056 -5622 2090 -5046
rect 2184 -5622 2218 -5046
rect 2296 -5622 2330 -5046
rect 2424 -5622 2458 -5046
rect 2536 -5622 2570 -5046
rect 2664 -5622 2698 -5046
rect 2776 -5622 2810 -5046
rect 2904 -5622 2938 -5046
rect -6522 -5804 -6484 -5672
rect -6282 -5804 -6244 -5672
rect -6042 -5804 -6004 -5672
rect -5802 -5804 -5764 -5672
rect -5562 -5804 -5524 -5672
rect -5322 -5804 -5284 -5672
rect -5082 -5804 -5044 -5672
rect -4842 -5804 -4804 -5672
rect -4602 -5804 -4564 -5672
rect -4362 -5804 -4324 -5672
rect -4122 -5804 -4084 -5672
rect -3882 -5804 -3844 -5672
rect -3642 -5804 -3604 -5672
rect -3402 -5804 -3364 -5672
rect -3162 -5804 -3124 -5672
rect -2922 -5804 -2884 -5672
rect -2682 -5804 -2644 -5672
rect -2442 -5804 -2404 -5672
rect -2202 -5804 -2164 -5672
rect -1962 -5804 -1924 -5672
rect -1722 -5804 -1684 -5672
rect -1482 -5804 -1444 -5672
rect -1242 -5804 -1204 -5672
rect -1002 -5804 -964 -5672
rect -762 -5804 -724 -5672
rect -522 -5804 -484 -5672
rect -282 -5804 -244 -5672
rect -42 -5804 -4 -5672
rect 198 -5804 236 -5672
rect 438 -5804 476 -5672
rect 678 -5804 716 -5672
rect 918 -5804 956 -5672
rect 1158 -5804 1196 -5672
rect 1398 -5804 1436 -5672
rect 1638 -5804 1676 -5672
rect 1878 -5804 1916 -5672
rect 2118 -5804 2156 -5672
rect 2358 -5804 2396 -5672
rect 2598 -5804 2636 -5672
rect 2838 -5804 2876 -5672
rect -15826 -8253 -15458 -8219
rect -15238 -8253 -14870 -8219
rect -14650 -8253 -14282 -8219
rect -14062 -8253 -13694 -8219
rect -13474 -8253 -13106 -8219
rect -12886 -8253 -12518 -8219
rect -12298 -8253 -11930 -8219
rect -11710 -8253 -11342 -8219
rect -11122 -8253 -10754 -8219
rect -10534 -8253 -10166 -8219
rect -9946 -8253 -9578 -8219
rect -9358 -8253 -8990 -8219
rect -8770 -8253 -8402 -8219
rect -8182 -8253 -7814 -8219
rect -7594 -8253 -7226 -8219
rect -7006 -8253 -6638 -8219
rect -6418 -8253 -6050 -8219
rect -5830 -8253 -5462 -8219
rect -5242 -8253 -4874 -8219
rect -4654 -8253 -4286 -8219
rect -4066 -8253 -3698 -8219
rect -3478 -8253 -3110 -8219
rect -2890 -8253 -2522 -8219
rect -2302 -8253 -1934 -8219
rect -1714 -8253 -1346 -8219
rect -1126 -8253 -758 -8219
rect -538 -8253 -170 -8219
rect 50 -8253 418 -8219
rect 638 -8253 1006 -8219
rect 1226 -8253 1594 -8219
rect 1814 -8253 2182 -8219
rect 2402 -8253 2770 -8219
rect 2990 -8253 3358 -8219
rect 3578 -8253 3946 -8219
rect 4166 -8253 4534 -8219
rect 4754 -8253 5122 -8219
rect 5342 -8253 5710 -8219
rect 5930 -8253 6298 -8219
rect 6518 -8253 6886 -8219
rect 7106 -8253 7474 -8219
rect 7694 -8253 8062 -8219
rect 8282 -8253 8650 -8219
rect 8870 -8253 9238 -8219
rect 9458 -8253 9826 -8219
rect 10046 -8253 10414 -8219
rect 10634 -8253 11002 -8219
rect 11222 -8253 11590 -8219
rect 11810 -8253 12178 -8219
rect -15888 -9088 -15854 -8312
rect -15430 -9088 -15396 -8312
rect -15300 -9088 -15266 -8312
rect -14842 -9088 -14808 -8312
rect -14712 -9088 -14678 -8312
rect -14254 -9088 -14220 -8312
rect -14124 -9088 -14090 -8312
rect -13666 -9088 -13632 -8312
rect -13536 -9088 -13502 -8312
rect -13078 -9088 -13044 -8312
rect -12948 -9088 -12914 -8312
rect -12490 -9088 -12456 -8312
rect -12360 -9088 -12326 -8312
rect -11902 -9088 -11868 -8312
rect -11772 -9088 -11738 -8312
rect -11314 -9088 -11280 -8312
rect -11184 -9088 -11150 -8312
rect -10726 -9088 -10692 -8312
rect -10596 -9088 -10562 -8312
rect -10138 -9088 -10104 -8312
rect -10008 -9088 -9974 -8312
rect -9550 -9088 -9516 -8312
rect -9420 -9088 -9386 -8312
rect -8962 -9088 -8928 -8312
rect -8832 -9088 -8798 -8312
rect -8374 -9088 -8340 -8312
rect -8244 -9088 -8210 -8312
rect -7786 -9088 -7752 -8312
rect -7656 -9088 -7622 -8312
rect -7198 -9088 -7164 -8312
rect -7068 -9088 -7034 -8312
rect -6610 -9088 -6576 -8312
rect -6480 -9088 -6446 -8312
rect -6022 -9088 -5988 -8312
rect -5892 -9088 -5858 -8312
rect -5434 -9088 -5400 -8312
rect -5304 -9088 -5270 -8312
rect -4846 -9088 -4812 -8312
rect -4716 -9088 -4682 -8312
rect -4258 -9088 -4224 -8312
rect -4128 -9088 -4094 -8312
rect -3670 -9088 -3636 -8312
rect -3540 -9088 -3506 -8312
rect -3082 -9088 -3048 -8312
rect -2952 -9088 -2918 -8312
rect -2494 -9088 -2460 -8312
rect -2364 -9088 -2330 -8312
rect -1906 -9088 -1872 -8312
rect -1776 -9088 -1742 -8312
rect -1318 -9088 -1284 -8312
rect -1188 -9088 -1154 -8312
rect -730 -9088 -696 -8312
rect -600 -9088 -566 -8312
rect -142 -9088 -108 -8312
rect -12 -9088 22 -8312
rect 446 -9088 480 -8312
rect 576 -9088 610 -8312
rect 1034 -9088 1068 -8312
rect 1164 -9088 1198 -8312
rect 1622 -9088 1656 -8312
rect 1752 -9088 1786 -8312
rect 2210 -9088 2244 -8312
rect 2340 -9088 2374 -8312
rect 2798 -9088 2832 -8312
rect 2928 -9088 2962 -8312
rect 3386 -9088 3420 -8312
rect 3516 -9088 3550 -8312
rect 3974 -9088 4008 -8312
rect 4104 -9088 4138 -8312
rect 4562 -9088 4596 -8312
rect 4692 -9088 4726 -8312
rect 5150 -9088 5184 -8312
rect 5280 -9088 5314 -8312
rect 5738 -9088 5772 -8312
rect 5868 -9088 5902 -8312
rect 6326 -9088 6360 -8312
rect 6456 -9088 6490 -8312
rect 6914 -9088 6948 -8312
rect 7044 -9088 7078 -8312
rect 7502 -9088 7536 -8312
rect 7632 -9088 7666 -8312
rect 8090 -9088 8124 -8312
rect 8220 -9088 8254 -8312
rect 8678 -9088 8712 -8312
rect 8808 -9088 8842 -8312
rect 9266 -9088 9300 -8312
rect 9396 -9088 9430 -8312
rect 9854 -9088 9888 -8312
rect 9984 -9088 10018 -8312
rect 10442 -9088 10476 -8312
rect 10572 -9088 10606 -8312
rect 11030 -9088 11064 -8312
rect 11160 -9088 11194 -8312
rect 11618 -9088 11652 -8312
rect 11748 -9088 11782 -8312
rect 12206 -9088 12240 -8312
rect -15826 -9181 -15458 -9147
rect -15238 -9181 -14870 -9147
rect -14650 -9181 -14282 -9147
rect -14062 -9181 -13694 -9147
rect -13474 -9181 -13106 -9147
rect -12886 -9181 -12518 -9147
rect -12298 -9181 -11930 -9147
rect -11710 -9181 -11342 -9147
rect -11122 -9181 -10754 -9147
rect -10534 -9181 -10166 -9147
rect -9946 -9181 -9578 -9147
rect -9358 -9181 -8990 -9147
rect -8770 -9181 -8402 -9147
rect -8182 -9181 -7814 -9147
rect -7594 -9181 -7226 -9147
rect -7006 -9181 -6638 -9147
rect -6418 -9181 -6050 -9147
rect -5830 -9181 -5462 -9147
rect -5242 -9181 -4874 -9147
rect -4654 -9181 -4286 -9147
rect -4066 -9181 -3698 -9147
rect -3478 -9181 -3110 -9147
rect -2890 -9181 -2522 -9147
rect -2302 -9181 -1934 -9147
rect -1714 -9181 -1346 -9147
rect -1126 -9181 -758 -9147
rect -538 -9181 -170 -9147
rect 50 -9181 418 -9147
rect 638 -9181 1006 -9147
rect 1226 -9181 1594 -9147
rect 1814 -9181 2182 -9147
rect 2402 -9181 2770 -9147
rect 2990 -9181 3358 -9147
rect 3578 -9181 3946 -9147
rect 4166 -9181 4534 -9147
rect 4754 -9181 5122 -9147
rect 5342 -9181 5710 -9147
rect 5930 -9181 6298 -9147
rect 6518 -9181 6886 -9147
rect 7106 -9181 7474 -9147
rect 7694 -9181 8062 -9147
rect 8282 -9181 8650 -9147
rect 8870 -9181 9238 -9147
rect 9458 -9181 9826 -9147
rect 10046 -9181 10414 -9147
rect 10634 -9181 11002 -9147
rect 11222 -9181 11590 -9147
rect 11810 -9181 12178 -9147
rect -15826 -9253 -15458 -9219
rect -15238 -9253 -14870 -9219
rect -14650 -9253 -14282 -9219
rect -14062 -9253 -13694 -9219
rect -13474 -9253 -13106 -9219
rect -12886 -9253 -12518 -9219
rect -12298 -9253 -11930 -9219
rect -11710 -9253 -11342 -9219
rect -11122 -9253 -10754 -9219
rect -10534 -9253 -10166 -9219
rect -9946 -9253 -9578 -9219
rect -9358 -9253 -8990 -9219
rect -8770 -9253 -8402 -9219
rect -8182 -9253 -7814 -9219
rect -7594 -9253 -7226 -9219
rect -7006 -9253 -6638 -9219
rect -6418 -9253 -6050 -9219
rect -5830 -9253 -5462 -9219
rect -5242 -9253 -4874 -9219
rect -4654 -9253 -4286 -9219
rect -4066 -9253 -3698 -9219
rect -3478 -9253 -3110 -9219
rect -2890 -9253 -2522 -9219
rect -2302 -9253 -1934 -9219
rect -1714 -9253 -1346 -9219
rect -1126 -9253 -758 -9219
rect -538 -9253 -170 -9219
rect 50 -9253 418 -9219
rect 638 -9253 1006 -9219
rect 1226 -9253 1594 -9219
rect 1814 -9253 2182 -9219
rect 2402 -9253 2770 -9219
rect 2990 -9253 3358 -9219
rect 3578 -9253 3946 -9219
rect 4166 -9253 4534 -9219
rect 4754 -9253 5122 -9219
rect 5342 -9253 5710 -9219
rect 5930 -9253 6298 -9219
rect 6518 -9253 6886 -9219
rect 7106 -9253 7474 -9219
rect 7694 -9253 8062 -9219
rect 8282 -9253 8650 -9219
rect 8870 -9253 9238 -9219
rect 9458 -9253 9826 -9219
rect 10046 -9253 10414 -9219
rect 10634 -9253 11002 -9219
rect 11222 -9253 11590 -9219
rect 11810 -9253 12178 -9219
rect -15888 -10088 -15854 -9312
rect -15430 -10088 -15396 -9312
rect -15300 -10088 -15266 -9312
rect -14842 -10088 -14808 -9312
rect -14712 -10088 -14678 -9312
rect -14254 -10088 -14220 -9312
rect -14124 -10088 -14090 -9312
rect -13666 -10088 -13632 -9312
rect -13536 -10088 -13502 -9312
rect -13078 -10088 -13044 -9312
rect -12948 -10088 -12914 -9312
rect -12490 -10088 -12456 -9312
rect -12360 -10088 -12326 -9312
rect -11902 -10088 -11868 -9312
rect -11772 -10088 -11738 -9312
rect -11314 -10088 -11280 -9312
rect -11184 -10088 -11150 -9312
rect -10726 -10088 -10692 -9312
rect -10596 -10088 -10562 -9312
rect -10138 -10088 -10104 -9312
rect -10008 -10088 -9974 -9312
rect -9550 -10088 -9516 -9312
rect -9420 -10088 -9386 -9312
rect -8962 -10088 -8928 -9312
rect -8832 -10088 -8798 -9312
rect -8374 -10088 -8340 -9312
rect -8244 -10088 -8210 -9312
rect -7786 -10088 -7752 -9312
rect -7656 -10088 -7622 -9312
rect -7198 -10088 -7164 -9312
rect -7068 -10088 -7034 -9312
rect -6610 -10088 -6576 -9312
rect -6480 -10088 -6446 -9312
rect -6022 -10088 -5988 -9312
rect -5892 -10088 -5858 -9312
rect -5434 -10088 -5400 -9312
rect -5304 -10088 -5270 -9312
rect -4846 -10088 -4812 -9312
rect -4716 -10088 -4682 -9312
rect -4258 -10088 -4224 -9312
rect -4128 -10088 -4094 -9312
rect -3670 -10088 -3636 -9312
rect -3540 -10088 -3506 -9312
rect -3082 -10088 -3048 -9312
rect -2952 -10088 -2918 -9312
rect -2494 -10088 -2460 -9312
rect -2364 -10088 -2330 -9312
rect -1906 -10088 -1872 -9312
rect -1776 -10088 -1742 -9312
rect -1318 -10088 -1284 -9312
rect -1188 -10088 -1154 -9312
rect -730 -10088 -696 -9312
rect -600 -10088 -566 -9312
rect -142 -10088 -108 -9312
rect -12 -10088 22 -9312
rect 446 -10088 480 -9312
rect 576 -10088 610 -9312
rect 1034 -10088 1068 -9312
rect 1164 -10088 1198 -9312
rect 1622 -10088 1656 -9312
rect 1752 -10088 1786 -9312
rect 2210 -10088 2244 -9312
rect 2340 -10088 2374 -9312
rect 2798 -10088 2832 -9312
rect 2928 -10088 2962 -9312
rect 3386 -10088 3420 -9312
rect 3516 -10088 3550 -9312
rect 3974 -10088 4008 -9312
rect 4104 -10088 4138 -9312
rect 4562 -10088 4596 -9312
rect 4692 -10088 4726 -9312
rect 5150 -10088 5184 -9312
rect 5280 -10088 5314 -9312
rect 5738 -10088 5772 -9312
rect 5868 -10088 5902 -9312
rect 6326 -10088 6360 -9312
rect 6456 -10088 6490 -9312
rect 6914 -10088 6948 -9312
rect 7044 -10088 7078 -9312
rect 7502 -10088 7536 -9312
rect 7632 -10088 7666 -9312
rect 8090 -10088 8124 -9312
rect 8220 -10088 8254 -9312
rect 8678 -10088 8712 -9312
rect 8808 -10088 8842 -9312
rect 9266 -10088 9300 -9312
rect 9396 -10088 9430 -9312
rect 9854 -10088 9888 -9312
rect 9984 -10088 10018 -9312
rect 10442 -10088 10476 -9312
rect 10572 -10088 10606 -9312
rect 11030 -10088 11064 -9312
rect 11160 -10088 11194 -9312
rect 11618 -10088 11652 -9312
rect 11748 -10088 11782 -9312
rect 12206 -10088 12240 -9312
rect -15826 -10181 -15458 -10147
rect -15238 -10181 -14870 -10147
rect -14650 -10181 -14282 -10147
rect -14062 -10181 -13694 -10147
rect -13474 -10181 -13106 -10147
rect -12886 -10181 -12518 -10147
rect -12298 -10181 -11930 -10147
rect -11710 -10181 -11342 -10147
rect -11122 -10181 -10754 -10147
rect -10534 -10181 -10166 -10147
rect -9946 -10181 -9578 -10147
rect -9358 -10181 -8990 -10147
rect -8770 -10181 -8402 -10147
rect -8182 -10181 -7814 -10147
rect -7594 -10181 -7226 -10147
rect -7006 -10181 -6638 -10147
rect -6418 -10181 -6050 -10147
rect -5830 -10181 -5462 -10147
rect -5242 -10181 -4874 -10147
rect -4654 -10181 -4286 -10147
rect -4066 -10181 -3698 -10147
rect -3478 -10181 -3110 -10147
rect -2890 -10181 -2522 -10147
rect -2302 -10181 -1934 -10147
rect -1714 -10181 -1346 -10147
rect -1126 -10181 -758 -10147
rect -538 -10181 -170 -10147
rect 50 -10181 418 -10147
rect 638 -10181 1006 -10147
rect 1226 -10181 1594 -10147
rect 1814 -10181 2182 -10147
rect 2402 -10181 2770 -10147
rect 2990 -10181 3358 -10147
rect 3578 -10181 3946 -10147
rect 4166 -10181 4534 -10147
rect 4754 -10181 5122 -10147
rect 5342 -10181 5710 -10147
rect 5930 -10181 6298 -10147
rect 6518 -10181 6886 -10147
rect 7106 -10181 7474 -10147
rect 7694 -10181 8062 -10147
rect 8282 -10181 8650 -10147
rect 8870 -10181 9238 -10147
rect 9458 -10181 9826 -10147
rect 10046 -10181 10414 -10147
rect 10634 -10181 11002 -10147
rect 11222 -10181 11590 -10147
rect 11810 -10181 12178 -10147
rect -15826 -10253 -15458 -10219
rect -15238 -10253 -14870 -10219
rect -14650 -10253 -14282 -10219
rect -14062 -10253 -13694 -10219
rect -13474 -10253 -13106 -10219
rect -12886 -10253 -12518 -10219
rect -12298 -10253 -11930 -10219
rect -11710 -10253 -11342 -10219
rect -11122 -10253 -10754 -10219
rect -10534 -10253 -10166 -10219
rect -9946 -10253 -9578 -10219
rect -9358 -10253 -8990 -10219
rect -8770 -10253 -8402 -10219
rect -8182 -10253 -7814 -10219
rect -7594 -10253 -7226 -10219
rect -7006 -10253 -6638 -10219
rect -6418 -10253 -6050 -10219
rect -5830 -10253 -5462 -10219
rect -5242 -10253 -4874 -10219
rect -4654 -10253 -4286 -10219
rect -4066 -10253 -3698 -10219
rect -3478 -10253 -3110 -10219
rect -2890 -10253 -2522 -10219
rect -2302 -10253 -1934 -10219
rect -1714 -10253 -1346 -10219
rect -1126 -10253 -758 -10219
rect -538 -10253 -170 -10219
rect 50 -10253 418 -10219
rect 638 -10253 1006 -10219
rect 1226 -10253 1594 -10219
rect 1814 -10253 2182 -10219
rect 2402 -10253 2770 -10219
rect 2990 -10253 3358 -10219
rect 3578 -10253 3946 -10219
rect 4166 -10253 4534 -10219
rect 4754 -10253 5122 -10219
rect 5342 -10253 5710 -10219
rect 5930 -10253 6298 -10219
rect 6518 -10253 6886 -10219
rect 7106 -10253 7474 -10219
rect 7694 -10253 8062 -10219
rect 8282 -10253 8650 -10219
rect 8870 -10253 9238 -10219
rect 9458 -10253 9826 -10219
rect 10046 -10253 10414 -10219
rect 10634 -10253 11002 -10219
rect 11222 -10253 11590 -10219
rect 11810 -10253 12178 -10219
rect -15888 -11088 -15854 -10312
rect -15430 -11088 -15396 -10312
rect -15300 -11088 -15266 -10312
rect -14842 -11088 -14808 -10312
rect -14712 -11088 -14678 -10312
rect -14254 -11088 -14220 -10312
rect -14124 -11088 -14090 -10312
rect -13666 -11088 -13632 -10312
rect -13536 -11088 -13502 -10312
rect -13078 -11088 -13044 -10312
rect -12948 -11088 -12914 -10312
rect -12490 -11088 -12456 -10312
rect -12360 -11088 -12326 -10312
rect -11902 -11088 -11868 -10312
rect -11772 -11088 -11738 -10312
rect -11314 -11088 -11280 -10312
rect -11184 -11088 -11150 -10312
rect -10726 -11088 -10692 -10312
rect -10596 -11088 -10562 -10312
rect -10138 -11088 -10104 -10312
rect -10008 -11088 -9974 -10312
rect -9550 -11088 -9516 -10312
rect -9420 -11088 -9386 -10312
rect -8962 -11088 -8928 -10312
rect -8832 -11088 -8798 -10312
rect -8374 -11088 -8340 -10312
rect -8244 -11088 -8210 -10312
rect -7786 -11088 -7752 -10312
rect -7656 -11088 -7622 -10312
rect -7198 -11088 -7164 -10312
rect -7068 -11088 -7034 -10312
rect -6610 -11088 -6576 -10312
rect -6480 -11088 -6446 -10312
rect -6022 -11088 -5988 -10312
rect -5892 -11088 -5858 -10312
rect -5434 -11088 -5400 -10312
rect -5304 -11088 -5270 -10312
rect -4846 -11088 -4812 -10312
rect -4716 -11088 -4682 -10312
rect -4258 -11088 -4224 -10312
rect -4128 -11088 -4094 -10312
rect -3670 -11088 -3636 -10312
rect -3540 -11088 -3506 -10312
rect -3082 -11088 -3048 -10312
rect -2952 -11088 -2918 -10312
rect -2494 -11088 -2460 -10312
rect -2364 -11088 -2330 -10312
rect -1906 -11088 -1872 -10312
rect -1776 -11088 -1742 -10312
rect -1318 -11088 -1284 -10312
rect -1188 -11088 -1154 -10312
rect -730 -11088 -696 -10312
rect -600 -11088 -566 -10312
rect -142 -11088 -108 -10312
rect -12 -11088 22 -10312
rect 446 -11088 480 -10312
rect 576 -11088 610 -10312
rect 1034 -11088 1068 -10312
rect 1164 -11088 1198 -10312
rect 1622 -11088 1656 -10312
rect 1752 -11088 1786 -10312
rect 2210 -11088 2244 -10312
rect 2340 -11088 2374 -10312
rect 2798 -11088 2832 -10312
rect 2928 -11088 2962 -10312
rect 3386 -11088 3420 -10312
rect 3516 -11088 3550 -10312
rect 3974 -11088 4008 -10312
rect 4104 -11088 4138 -10312
rect 4562 -11088 4596 -10312
rect 4692 -11088 4726 -10312
rect 5150 -11088 5184 -10312
rect 5280 -11088 5314 -10312
rect 5738 -11088 5772 -10312
rect 5868 -11088 5902 -10312
rect 6326 -11088 6360 -10312
rect 6456 -11088 6490 -10312
rect 6914 -11088 6948 -10312
rect 7044 -11088 7078 -10312
rect 7502 -11088 7536 -10312
rect 7632 -11088 7666 -10312
rect 8090 -11088 8124 -10312
rect 8220 -11088 8254 -10312
rect 8678 -11088 8712 -10312
rect 8808 -11088 8842 -10312
rect 9266 -11088 9300 -10312
rect 9396 -11088 9430 -10312
rect 9854 -11088 9888 -10312
rect 9984 -11088 10018 -10312
rect 10442 -11088 10476 -10312
rect 10572 -11088 10606 -10312
rect 11030 -11088 11064 -10312
rect 11160 -11088 11194 -10312
rect 11618 -11088 11652 -10312
rect 11748 -11088 11782 -10312
rect 12206 -11088 12240 -10312
rect -15826 -11181 -15458 -11147
rect -15238 -11181 -14870 -11147
rect -14650 -11181 -14282 -11147
rect -14062 -11181 -13694 -11147
rect -13474 -11181 -13106 -11147
rect -12886 -11181 -12518 -11147
rect -12298 -11181 -11930 -11147
rect -11710 -11181 -11342 -11147
rect -11122 -11181 -10754 -11147
rect -10534 -11181 -10166 -11147
rect -9946 -11181 -9578 -11147
rect -9358 -11181 -8990 -11147
rect -8770 -11181 -8402 -11147
rect -8182 -11181 -7814 -11147
rect -7594 -11181 -7226 -11147
rect -7006 -11181 -6638 -11147
rect -6418 -11181 -6050 -11147
rect -5830 -11181 -5462 -11147
rect -5242 -11181 -4874 -11147
rect -4654 -11181 -4286 -11147
rect -4066 -11181 -3698 -11147
rect -3478 -11181 -3110 -11147
rect -2890 -11181 -2522 -11147
rect -2302 -11181 -1934 -11147
rect -1714 -11181 -1346 -11147
rect -1126 -11181 -758 -11147
rect -538 -11181 -170 -11147
rect 50 -11181 418 -11147
rect 638 -11181 1006 -11147
rect 1226 -11181 1594 -11147
rect 1814 -11181 2182 -11147
rect 2402 -11181 2770 -11147
rect 2990 -11181 3358 -11147
rect 3578 -11181 3946 -11147
rect 4166 -11181 4534 -11147
rect 4754 -11181 5122 -11147
rect 5342 -11181 5710 -11147
rect 5930 -11181 6298 -11147
rect 6518 -11181 6886 -11147
rect 7106 -11181 7474 -11147
rect 7694 -11181 8062 -11147
rect 8282 -11181 8650 -11147
rect 8870 -11181 9238 -11147
rect 9458 -11181 9826 -11147
rect 10046 -11181 10414 -11147
rect 10634 -11181 11002 -11147
rect 11222 -11181 11590 -11147
rect 11810 -11181 12178 -11147
rect -15442 -11498 -15254 -11450
rect -14266 -11498 -14078 -11450
rect -13090 -11498 -12902 -11450
rect -11914 -11498 -11726 -11450
rect -10738 -11498 -10550 -11450
rect -9562 -11498 -9374 -11450
rect -8386 -11498 -8198 -11450
rect -7210 -11498 -7022 -11450
rect -6034 -11498 -5846 -11450
rect -4858 -11498 -4670 -11450
rect -3682 -11498 -3494 -11450
rect -2506 -11498 -2318 -11450
rect -1330 -11498 -1142 -11450
rect -154 -11498 34 -11450
rect 1022 -11498 1210 -11450
rect 2198 -11498 2386 -11450
rect 3374 -11498 3562 -11440
rect 4550 -11498 4738 -11450
rect 5726 -11498 5914 -11450
rect 6902 -11498 7090 -11450
rect 8064 -11498 8276 -11440
rect 9254 -11498 9442 -11450
rect 10430 -11498 10618 -11450
rect 11606 -11498 11794 -11450
rect -15442 -11532 -15254 -11498
rect -14266 -11532 -14078 -11498
rect -13090 -11532 -12902 -11498
rect -11914 -11532 -11726 -11498
rect -10738 -11532 -10550 -11498
rect -9562 -11532 -9374 -11498
rect -8386 -11532 -8198 -11498
rect -7210 -11532 -7022 -11498
rect -6034 -11532 -5846 -11498
rect -4858 -11532 -4670 -11498
rect -3682 -11532 -3494 -11498
rect -2506 -11532 -2318 -11498
rect -1330 -11532 -1142 -11498
rect -154 -11532 34 -11498
rect 1022 -11532 1210 -11498
rect 2198 -11532 2386 -11498
rect 3374 -11532 3562 -11498
rect 4550 -11532 4738 -11498
rect 5726 -11532 5914 -11498
rect 6902 -11532 7090 -11498
rect 8064 -11532 8276 -11498
rect 9254 -11532 9442 -11498
rect 10430 -11532 10618 -11498
rect 11606 -11532 11794 -11498
rect -15442 -11560 -15254 -11532
rect -14266 -11560 -14078 -11532
rect -13090 -11560 -12902 -11532
rect -11914 -11560 -11726 -11532
rect -10738 -11560 -10550 -11532
rect -9562 -11560 -9374 -11532
rect -8386 -11560 -8198 -11532
rect -7210 -11560 -7022 -11532
rect -6034 -11560 -5846 -11532
rect -4858 -11560 -4670 -11532
rect -3682 -11560 -3494 -11532
rect -2506 -11560 -2318 -11532
rect -1330 -11560 -1142 -11532
rect -154 -11560 34 -11532
rect 1022 -11560 1210 -11532
rect 2198 -11560 2386 -11532
rect 3374 -11550 3562 -11532
rect 4550 -11560 4738 -11532
rect 5726 -11560 5914 -11532
rect 6902 -11560 7090 -11532
rect 8064 -11562 8276 -11532
rect 9254 -11560 9442 -11532
rect 10430 -11560 10618 -11532
rect 11606 -11560 11794 -11532
rect -2774 -12708 -2736 -12576
rect -2508 -12708 -2470 -12576
rect -2242 -12708 -2204 -12576
rect -1976 -12708 -1938 -12576
rect -1710 -12708 -1672 -12576
rect -1444 -12708 -1406 -12576
rect -1178 -12708 -1140 -12576
rect -912 -12708 -874 -12576
rect -2836 -13534 -2802 -12758
rect -2708 -13534 -2674 -12758
rect -2570 -13534 -2536 -12758
rect -2442 -13534 -2408 -12758
rect -2304 -13534 -2270 -12758
rect -2176 -13534 -2142 -12758
rect -2038 -13534 -2004 -12758
rect -1910 -13534 -1876 -12758
rect -1772 -13534 -1738 -12758
rect -1644 -13534 -1610 -12758
rect -1506 -13534 -1472 -12758
rect -1378 -13534 -1344 -12758
rect -1240 -13534 -1206 -12758
rect -1112 -13534 -1078 -12758
rect -974 -13534 -940 -12758
rect -846 -13534 -812 -12758
rect -2774 -13718 -2736 -13586
rect -2508 -13718 -2470 -13586
rect -2242 -13718 -2204 -13586
rect -1976 -13718 -1938 -13586
rect -1710 -13718 -1672 -13586
rect -1444 -13718 -1406 -13586
rect -1178 -13718 -1140 -13586
rect -912 -13718 -874 -13586
rect -2836 -14544 -2802 -13768
rect -2708 -14544 -2674 -13768
rect -2570 -14544 -2536 -13768
rect -2442 -14544 -2408 -13768
rect -2304 -14544 -2270 -13768
rect -2176 -14544 -2142 -13768
rect -2038 -14544 -2004 -13768
rect -1910 -14544 -1876 -13768
rect -1772 -14544 -1738 -13768
rect -1644 -14544 -1610 -13768
rect -1506 -14544 -1472 -13768
rect -1378 -14544 -1344 -13768
rect -1240 -14544 -1206 -13768
rect -1112 -14544 -1078 -13768
rect -974 -14544 -940 -13768
rect -846 -14544 -812 -13768
rect -2774 -14728 -2736 -14596
rect -2508 -14728 -2470 -14596
rect -2242 -14728 -2204 -14596
rect -1976 -14728 -1938 -14596
rect -1710 -14728 -1672 -14596
rect -1444 -14728 -1406 -14596
rect -1178 -14728 -1140 -14596
rect -912 -14728 -874 -14596
rect -2836 -15554 -2802 -14778
rect -2708 -15554 -2674 -14778
rect -2570 -15554 -2536 -14778
rect -2442 -15554 -2408 -14778
rect -2304 -15554 -2270 -14778
rect -2176 -15554 -2142 -14778
rect -2038 -15554 -2004 -14778
rect -1910 -15554 -1876 -14778
rect -1772 -15554 -1738 -14778
rect -1644 -15554 -1610 -14778
rect -1506 -15554 -1472 -14778
rect -1378 -15554 -1344 -14778
rect -1240 -15554 -1206 -14778
rect -1112 -15554 -1078 -14778
rect -974 -15554 -940 -14778
rect -846 -15554 -812 -14778
rect -2774 -15738 -2736 -15606
rect -2508 -15738 -2470 -15606
rect -2242 -15738 -2204 -15606
rect -1976 -15738 -1938 -15606
rect -1710 -15738 -1672 -15606
rect -1444 -15738 -1406 -15606
rect -1178 -15738 -1140 -15606
rect -912 -15738 -874 -15606
rect 4383 -15394 4421 -14997
rect 4383 -15925 4421 -15528
rect 4634 -15338 4774 -14878
rect -2202 -16900 -2164 -16774
rect -1962 -16900 -1924 -16774
rect -1722 -16900 -1684 -16774
rect -1482 -16900 -1444 -16774
rect -2264 -17526 -2230 -16950
rect -2136 -17526 -2102 -16950
rect -2024 -17526 -1990 -16950
rect -1896 -17526 -1862 -16950
rect -1784 -17526 -1750 -16950
rect -1656 -17526 -1622 -16950
rect -1544 -17526 -1510 -16950
rect -1416 -17526 -1382 -16950
rect -2202 -17708 -2164 -17576
rect -1962 -17708 -1924 -17576
rect -1722 -17708 -1684 -17576
rect -1482 -17708 -1444 -17576
rect -2264 -18334 -2230 -17758
rect -2136 -18334 -2102 -17758
rect -2024 -18334 -1990 -17758
rect -1896 -18334 -1862 -17758
rect -1784 -18334 -1750 -17758
rect -1656 -18334 -1622 -17758
rect -1544 -18334 -1510 -17758
rect -1416 -18334 -1382 -17758
rect -2202 -18516 -2164 -18384
rect -1962 -18516 -1924 -18384
rect -1722 -18516 -1684 -18384
rect -1482 -18516 -1444 -18384
rect -2512 -18816 -1160 -18768
rect -2512 -18850 -2452 -18816
rect -2452 -18850 -1242 -18816
rect -1242 -18850 -1160 -18816
rect -2512 -18880 -1160 -18850
<< metal1 >>
rect -6450 -3712 -6316 -3706
rect -6450 -3784 -6438 -3712
rect -6328 -3784 -6316 -3712
rect -6450 -3790 -6316 -3784
rect -5970 -3712 -5836 -3706
rect -5970 -3784 -5958 -3712
rect -5848 -3784 -5836 -3712
rect -5970 -3790 -5836 -3784
rect -5490 -3712 -5356 -3706
rect -5490 -3784 -5478 -3712
rect -5368 -3784 -5356 -3712
rect -5490 -3790 -5356 -3784
rect -5010 -3712 -4876 -3706
rect -5010 -3784 -4998 -3712
rect -4888 -3784 -4876 -3712
rect -5010 -3790 -4876 -3784
rect -4530 -3712 -4396 -3706
rect -4530 -3784 -4518 -3712
rect -4408 -3784 -4396 -3712
rect -4530 -3790 -4396 -3784
rect -4050 -3712 -3916 -3706
rect -4050 -3784 -4038 -3712
rect -3928 -3784 -3916 -3712
rect -4050 -3790 -3916 -3784
rect -3570 -3712 -3436 -3706
rect -3570 -3784 -3558 -3712
rect -3448 -3784 -3436 -3712
rect -3570 -3790 -3436 -3784
rect -3090 -3712 -2956 -3706
rect -3090 -3784 -3078 -3712
rect -2968 -3784 -2956 -3712
rect -3090 -3790 -2956 -3784
rect -2610 -3712 -2476 -3706
rect -2610 -3784 -2598 -3712
rect -2488 -3784 -2476 -3712
rect -2610 -3790 -2476 -3784
rect -2130 -3712 -1996 -3706
rect -2130 -3784 -2118 -3712
rect -2008 -3784 -1996 -3712
rect -2130 -3790 -1996 -3784
rect -1650 -3712 -1516 -3706
rect -1650 -3784 -1638 -3712
rect -1528 -3784 -1516 -3712
rect -1650 -3790 -1516 -3784
rect -1170 -3712 -1036 -3706
rect -1170 -3784 -1158 -3712
rect -1048 -3784 -1036 -3712
rect -1170 -3790 -1036 -3784
rect -690 -3712 -556 -3706
rect -690 -3784 -678 -3712
rect -568 -3784 -556 -3712
rect -690 -3790 -556 -3784
rect -210 -3712 -76 -3706
rect -210 -3784 -198 -3712
rect -88 -3784 -76 -3712
rect -210 -3790 -76 -3784
rect 270 -3712 404 -3706
rect 270 -3784 282 -3712
rect 392 -3784 404 -3712
rect 270 -3790 404 -3784
rect 750 -3712 884 -3706
rect 750 -3784 762 -3712
rect 872 -3784 884 -3712
rect 750 -3790 884 -3784
rect 1230 -3712 1364 -3706
rect 1230 -3784 1242 -3712
rect 1352 -3784 1364 -3712
rect 1230 -3790 1364 -3784
rect 1710 -3712 1844 -3706
rect 1710 -3784 1722 -3712
rect 1832 -3784 1844 -3712
rect 1710 -3790 1844 -3784
rect 2190 -3712 2324 -3706
rect 2190 -3784 2202 -3712
rect 2312 -3784 2324 -3712
rect 2190 -3790 2324 -3784
rect 2670 -3712 2804 -3706
rect 2670 -3784 2682 -3712
rect 2792 -3784 2804 -3712
rect 2670 -3790 2804 -3784
rect -6538 -4056 -6468 -4050
rect -6548 -4188 -6538 -4056
rect -6468 -4188 -6458 -4056
rect -6538 -4194 -6468 -4188
rect -6410 -4226 -6356 -3790
rect -6298 -4056 -6228 -4050
rect -6308 -4188 -6298 -4056
rect -6228 -4188 -6218 -4056
rect -6298 -4194 -6228 -4188
rect -6170 -4198 -6116 -4046
rect -6058 -4056 -5988 -4050
rect -6068 -4188 -6058 -4056
rect -5988 -4188 -5978 -4056
rect -6058 -4194 -5988 -4188
rect -5930 -4226 -5876 -3790
rect -5818 -4056 -5748 -4050
rect -5828 -4188 -5818 -4056
rect -5748 -4188 -5738 -4056
rect -5818 -4194 -5748 -4188
rect -5690 -4198 -5636 -4046
rect -5578 -4056 -5508 -4050
rect -5588 -4188 -5578 -4056
rect -5508 -4188 -5498 -4056
rect -5578 -4194 -5508 -4188
rect -5450 -4226 -5396 -3790
rect -5338 -4056 -5268 -4050
rect -5348 -4188 -5338 -4056
rect -5268 -4188 -5258 -4056
rect -5338 -4194 -5268 -4188
rect -5210 -4198 -5156 -4046
rect -5098 -4056 -5028 -4050
rect -5108 -4188 -5098 -4056
rect -5028 -4188 -5018 -4056
rect -5098 -4194 -5028 -4188
rect -4970 -4226 -4916 -3790
rect -4858 -4056 -4788 -4050
rect -4868 -4188 -4858 -4056
rect -4788 -4188 -4778 -4056
rect -4858 -4194 -4788 -4188
rect -4730 -4198 -4676 -4046
rect -4618 -4056 -4548 -4050
rect -4628 -4188 -4618 -4056
rect -4548 -4188 -4538 -4056
rect -4618 -4194 -4548 -4188
rect -4490 -4226 -4436 -3790
rect -4378 -4056 -4308 -4050
rect -4388 -4188 -4378 -4056
rect -4308 -4188 -4298 -4056
rect -4378 -4194 -4308 -4188
rect -4250 -4198 -4196 -4046
rect -4138 -4056 -4068 -4050
rect -4148 -4188 -4138 -4056
rect -4068 -4188 -4058 -4056
rect -4138 -4194 -4068 -4188
rect -4010 -4226 -3956 -3790
rect -3898 -4056 -3828 -4050
rect -3908 -4188 -3898 -4056
rect -3828 -4188 -3818 -4056
rect -3898 -4194 -3828 -4188
rect -3770 -4198 -3716 -4046
rect -3658 -4056 -3588 -4050
rect -3668 -4188 -3658 -4056
rect -3588 -4188 -3578 -4056
rect -3658 -4194 -3588 -4188
rect -3530 -4226 -3476 -3790
rect -3418 -4056 -3348 -4050
rect -3428 -4188 -3418 -4056
rect -3348 -4188 -3338 -4056
rect -3418 -4194 -3348 -4188
rect -3290 -4198 -3236 -4046
rect -3178 -4056 -3108 -4050
rect -3188 -4188 -3178 -4056
rect -3108 -4188 -3098 -4056
rect -3178 -4194 -3108 -4188
rect -3050 -4226 -2996 -3790
rect -2938 -4056 -2868 -4050
rect -2948 -4188 -2938 -4056
rect -2868 -4188 -2858 -4056
rect -2938 -4194 -2868 -4188
rect -2810 -4198 -2756 -4046
rect -2698 -4056 -2628 -4050
rect -2708 -4188 -2698 -4056
rect -2628 -4188 -2618 -4056
rect -2698 -4194 -2628 -4188
rect -2570 -4226 -2516 -3790
rect -2458 -4056 -2388 -4050
rect -2468 -4188 -2458 -4056
rect -2388 -4188 -2378 -4056
rect -2458 -4194 -2388 -4188
rect -2330 -4198 -2276 -4046
rect -2218 -4056 -2148 -4050
rect -2228 -4188 -2218 -4056
rect -2148 -4188 -2138 -4056
rect -2218 -4194 -2148 -4188
rect -2090 -4226 -2036 -3790
rect -1978 -4056 -1908 -4050
rect -1988 -4188 -1978 -4056
rect -1908 -4188 -1898 -4056
rect -1978 -4194 -1908 -4188
rect -1850 -4198 -1796 -4046
rect -1738 -4056 -1668 -4050
rect -1748 -4188 -1738 -4056
rect -1668 -4188 -1658 -4056
rect -1738 -4194 -1668 -4188
rect -1610 -4226 -1556 -3790
rect -1498 -4056 -1428 -4050
rect -1508 -4188 -1498 -4056
rect -1428 -4188 -1418 -4056
rect -1498 -4194 -1428 -4188
rect -1370 -4198 -1316 -4046
rect -1258 -4056 -1188 -4050
rect -1268 -4188 -1258 -4056
rect -1188 -4188 -1178 -4056
rect -1258 -4194 -1188 -4188
rect -1130 -4226 -1076 -3790
rect -1018 -4056 -948 -4050
rect -1028 -4188 -1018 -4056
rect -948 -4188 -938 -4056
rect -1018 -4194 -948 -4188
rect -890 -4198 -836 -4046
rect -778 -4056 -708 -4050
rect -788 -4188 -778 -4056
rect -708 -4188 -698 -4056
rect -778 -4194 -708 -4188
rect -650 -4226 -596 -3790
rect -538 -4056 -468 -4050
rect -548 -4188 -538 -4056
rect -468 -4188 -458 -4056
rect -538 -4194 -468 -4188
rect -410 -4198 -356 -4046
rect -298 -4056 -228 -4050
rect -308 -4188 -298 -4056
rect -228 -4188 -218 -4056
rect -298 -4194 -228 -4188
rect -170 -4226 -116 -3790
rect -58 -4056 12 -4050
rect -68 -4188 -58 -4056
rect 12 -4188 22 -4056
rect -58 -4194 12 -4188
rect 70 -4198 124 -4046
rect 182 -4056 252 -4050
rect 172 -4188 182 -4056
rect 252 -4188 262 -4056
rect 182 -4194 252 -4188
rect 310 -4226 364 -3790
rect 422 -4056 492 -4050
rect 412 -4188 422 -4056
rect 492 -4188 502 -4056
rect 422 -4194 492 -4188
rect 550 -4198 604 -4046
rect 662 -4056 732 -4050
rect 652 -4188 662 -4056
rect 732 -4188 742 -4056
rect 662 -4194 732 -4188
rect 790 -4226 844 -3790
rect 902 -4056 972 -4050
rect 892 -4188 902 -4056
rect 972 -4188 982 -4056
rect 902 -4194 972 -4188
rect 1030 -4198 1084 -4046
rect 1142 -4056 1212 -4050
rect 1132 -4188 1142 -4056
rect 1212 -4188 1222 -4056
rect 1142 -4194 1212 -4188
rect 1270 -4226 1324 -3790
rect 1382 -4056 1452 -4050
rect 1372 -4188 1382 -4056
rect 1452 -4188 1462 -4056
rect 1382 -4194 1452 -4188
rect 1510 -4198 1564 -4046
rect 1622 -4056 1692 -4050
rect 1612 -4188 1622 -4056
rect 1692 -4188 1702 -4056
rect 1622 -4194 1692 -4188
rect 1750 -4226 1804 -3790
rect 1862 -4056 1932 -4050
rect 1852 -4188 1862 -4056
rect 1932 -4188 1942 -4056
rect 1862 -4194 1932 -4188
rect 1990 -4198 2044 -4046
rect 2102 -4056 2172 -4050
rect 2092 -4188 2102 -4056
rect 2172 -4188 2182 -4056
rect 2102 -4194 2172 -4188
rect 2230 -4226 2284 -3790
rect 2342 -4056 2412 -4050
rect 2332 -4188 2342 -4056
rect 2412 -4188 2422 -4056
rect 2342 -4194 2412 -4188
rect 2470 -4198 2524 -4046
rect 2582 -4056 2652 -4050
rect 2572 -4188 2582 -4056
rect 2652 -4188 2662 -4056
rect 2582 -4194 2652 -4188
rect 2710 -4226 2764 -3790
rect 2822 -4056 2892 -4050
rect 2812 -4188 2822 -4056
rect 2892 -4188 2902 -4056
rect 2822 -4194 2892 -4188
rect -6662 -4238 -6544 -4226
rect -6662 -4814 -6584 -4238
rect -6550 -4814 -6544 -4238
rect -6662 -4826 -6544 -4814
rect -6462 -4238 -6304 -4226
rect -6462 -4814 -6456 -4238
rect -6422 -4814 -6344 -4238
rect -6310 -4814 -6304 -4238
rect -6462 -4826 -6304 -4814
rect -6222 -4238 -6064 -4226
rect -6222 -4814 -6216 -4238
rect -6182 -4814 -6104 -4238
rect -6070 -4814 -6064 -4238
rect -6222 -4826 -6064 -4814
rect -5982 -4238 -5824 -4226
rect -5982 -4814 -5976 -4238
rect -5942 -4814 -5864 -4238
rect -5830 -4814 -5824 -4238
rect -5982 -4826 -5824 -4814
rect -5742 -4238 -5584 -4226
rect -5742 -4814 -5736 -4238
rect -5702 -4814 -5624 -4238
rect -5590 -4814 -5584 -4238
rect -5742 -4826 -5584 -4814
rect -5502 -4238 -5344 -4226
rect -5502 -4814 -5496 -4238
rect -5462 -4814 -5384 -4238
rect -5350 -4814 -5344 -4238
rect -5502 -4826 -5344 -4814
rect -5262 -4238 -5104 -4226
rect -5262 -4814 -5256 -4238
rect -5222 -4814 -5144 -4238
rect -5110 -4814 -5104 -4238
rect -5262 -4826 -5104 -4814
rect -5022 -4238 -4864 -4226
rect -5022 -4814 -5016 -4238
rect -4982 -4814 -4904 -4238
rect -4870 -4814 -4864 -4238
rect -5022 -4826 -4864 -4814
rect -4782 -4238 -4624 -4226
rect -4782 -4814 -4776 -4238
rect -4742 -4814 -4664 -4238
rect -4630 -4814 -4624 -4238
rect -4782 -4826 -4624 -4814
rect -4542 -4238 -4384 -4226
rect -4542 -4814 -4536 -4238
rect -4502 -4814 -4424 -4238
rect -4390 -4814 -4384 -4238
rect -4542 -4826 -4384 -4814
rect -4302 -4238 -4144 -4226
rect -4302 -4814 -4296 -4238
rect -4262 -4814 -4184 -4238
rect -4150 -4814 -4144 -4238
rect -4302 -4826 -4144 -4814
rect -4062 -4238 -3904 -4226
rect -4062 -4814 -4056 -4238
rect -4022 -4814 -3944 -4238
rect -3910 -4814 -3904 -4238
rect -4062 -4826 -3904 -4814
rect -3822 -4238 -3664 -4226
rect -3822 -4814 -3816 -4238
rect -3782 -4814 -3704 -4238
rect -3670 -4814 -3664 -4238
rect -3822 -4826 -3664 -4814
rect -3582 -4238 -3424 -4226
rect -3582 -4814 -3576 -4238
rect -3542 -4814 -3464 -4238
rect -3430 -4814 -3424 -4238
rect -3582 -4826 -3424 -4814
rect -3342 -4238 -3184 -4226
rect -3342 -4814 -3336 -4238
rect -3302 -4814 -3224 -4238
rect -3190 -4814 -3184 -4238
rect -3342 -4826 -3184 -4814
rect -3102 -4238 -2944 -4226
rect -3102 -4814 -3096 -4238
rect -3062 -4814 -2984 -4238
rect -2950 -4814 -2944 -4238
rect -3102 -4826 -2944 -4814
rect -2862 -4238 -2704 -4226
rect -2862 -4814 -2856 -4238
rect -2822 -4814 -2744 -4238
rect -2710 -4814 -2704 -4238
rect -2862 -4826 -2704 -4814
rect -2622 -4238 -2464 -4226
rect -2622 -4814 -2616 -4238
rect -2582 -4814 -2504 -4238
rect -2470 -4814 -2464 -4238
rect -2622 -4826 -2464 -4814
rect -2382 -4238 -2224 -4226
rect -2382 -4814 -2376 -4238
rect -2342 -4814 -2264 -4238
rect -2230 -4814 -2224 -4238
rect -2382 -4826 -2224 -4814
rect -2142 -4238 -1984 -4226
rect -2142 -4814 -2136 -4238
rect -2102 -4814 -2024 -4238
rect -1990 -4814 -1984 -4238
rect -2142 -4826 -1984 -4814
rect -1902 -4238 -1744 -4226
rect -1902 -4814 -1896 -4238
rect -1862 -4814 -1784 -4238
rect -1750 -4814 -1744 -4238
rect -1902 -4826 -1744 -4814
rect -1662 -4238 -1504 -4226
rect -1662 -4814 -1656 -4238
rect -1622 -4814 -1544 -4238
rect -1510 -4814 -1504 -4238
rect -1662 -4826 -1504 -4814
rect -1422 -4238 -1264 -4226
rect -1422 -4814 -1416 -4238
rect -1382 -4814 -1304 -4238
rect -1270 -4814 -1264 -4238
rect -1422 -4826 -1264 -4814
rect -1182 -4238 -1024 -4226
rect -1182 -4814 -1176 -4238
rect -1142 -4814 -1064 -4238
rect -1030 -4814 -1024 -4238
rect -1182 -4826 -1024 -4814
rect -942 -4238 -784 -4226
rect -942 -4814 -936 -4238
rect -902 -4814 -824 -4238
rect -790 -4814 -784 -4238
rect -942 -4826 -784 -4814
rect -702 -4238 -544 -4226
rect -702 -4814 -696 -4238
rect -662 -4814 -584 -4238
rect -550 -4814 -544 -4238
rect -702 -4826 -544 -4814
rect -462 -4238 -304 -4226
rect -462 -4814 -456 -4238
rect -422 -4814 -344 -4238
rect -310 -4814 -304 -4238
rect -462 -4826 -304 -4814
rect -222 -4238 -64 -4226
rect -222 -4814 -216 -4238
rect -182 -4814 -104 -4238
rect -70 -4814 -64 -4238
rect -222 -4826 -64 -4814
rect 18 -4238 176 -4226
rect 18 -4814 24 -4238
rect 58 -4814 136 -4238
rect 170 -4814 176 -4238
rect 18 -4826 176 -4814
rect 258 -4238 416 -4226
rect 258 -4814 264 -4238
rect 298 -4814 376 -4238
rect 410 -4814 416 -4238
rect 258 -4826 416 -4814
rect 498 -4238 656 -4226
rect 498 -4814 504 -4238
rect 538 -4814 616 -4238
rect 650 -4814 656 -4238
rect 498 -4826 656 -4814
rect 738 -4238 896 -4226
rect 738 -4814 744 -4238
rect 778 -4814 856 -4238
rect 890 -4814 896 -4238
rect 738 -4826 896 -4814
rect 978 -4238 1136 -4226
rect 978 -4814 984 -4238
rect 1018 -4814 1096 -4238
rect 1130 -4814 1136 -4238
rect 978 -4826 1136 -4814
rect 1218 -4238 1376 -4226
rect 1218 -4814 1224 -4238
rect 1258 -4814 1336 -4238
rect 1370 -4814 1376 -4238
rect 1218 -4826 1376 -4814
rect 1458 -4238 1616 -4226
rect 1458 -4814 1464 -4238
rect 1498 -4814 1576 -4238
rect 1610 -4814 1616 -4238
rect 1458 -4826 1616 -4814
rect 1698 -4238 1856 -4226
rect 1698 -4814 1704 -4238
rect 1738 -4814 1816 -4238
rect 1850 -4814 1856 -4238
rect 1698 -4826 1856 -4814
rect 1938 -4238 2096 -4226
rect 1938 -4814 1944 -4238
rect 1978 -4814 2056 -4238
rect 2090 -4814 2096 -4238
rect 1938 -4826 2096 -4814
rect 2178 -4238 2336 -4226
rect 2178 -4814 2184 -4238
rect 2218 -4814 2296 -4238
rect 2330 -4814 2336 -4238
rect 2178 -4826 2336 -4814
rect 2418 -4238 2576 -4226
rect 2418 -4814 2424 -4238
rect 2458 -4814 2536 -4238
rect 2570 -4814 2576 -4238
rect 2418 -4826 2576 -4814
rect 2658 -4238 2816 -4226
rect 2658 -4814 2664 -4238
rect 2698 -4814 2776 -4238
rect 2810 -4814 2816 -4238
rect 2658 -4826 2816 -4814
rect 2898 -4238 3016 -4226
rect 2898 -4814 2904 -4238
rect 2938 -4814 3016 -4238
rect 2898 -4826 3016 -4814
rect -6662 -5034 -6584 -4826
rect -6538 -4864 -6468 -4858
rect -6548 -4996 -6538 -4864
rect -6468 -4996 -6458 -4864
rect -6538 -5002 -6468 -4996
rect -6416 -5034 -6350 -4826
rect -6298 -4864 -6228 -4858
rect -6308 -4996 -6298 -4864
rect -6228 -4996 -6218 -4864
rect -6298 -5002 -6228 -4996
rect -6176 -5034 -6110 -4826
rect -6058 -4864 -5988 -4858
rect -6068 -4996 -6058 -4864
rect -5988 -4996 -5978 -4864
rect -6058 -5002 -5988 -4996
rect -5936 -5034 -5870 -4826
rect -5818 -4864 -5748 -4858
rect -5828 -4996 -5818 -4864
rect -5748 -4996 -5738 -4864
rect -5818 -5002 -5748 -4996
rect -5702 -5034 -5624 -4826
rect -5578 -4864 -5508 -4858
rect -5588 -4996 -5578 -4864
rect -5508 -4996 -5498 -4864
rect -5578 -5002 -5508 -4996
rect -5456 -5034 -5390 -4826
rect -5338 -4864 -5268 -4858
rect -5348 -4996 -5338 -4864
rect -5268 -4996 -5258 -4864
rect -5338 -5002 -5268 -4996
rect -5216 -5034 -5150 -4826
rect -5098 -4864 -5028 -4858
rect -5108 -4996 -5098 -4864
rect -5028 -4996 -5018 -4864
rect -5098 -5002 -5028 -4996
rect -4976 -5034 -4910 -4826
rect -4858 -4864 -4788 -4858
rect -4868 -4996 -4858 -4864
rect -4788 -4996 -4778 -4864
rect -4858 -5002 -4788 -4996
rect -4742 -5034 -4664 -4826
rect -4618 -4864 -4548 -4858
rect -4628 -4996 -4618 -4864
rect -4548 -4996 -4538 -4864
rect -4618 -5002 -4548 -4996
rect -4496 -5034 -4430 -4826
rect -4378 -4864 -4308 -4858
rect -4388 -4996 -4378 -4864
rect -4308 -4996 -4298 -4864
rect -4378 -5002 -4308 -4996
rect -4256 -5034 -4190 -4826
rect -4138 -4864 -4068 -4858
rect -4148 -4996 -4138 -4864
rect -4068 -4996 -4058 -4864
rect -4138 -5002 -4068 -4996
rect -4016 -5034 -3950 -4826
rect -3898 -4864 -3828 -4858
rect -3908 -4996 -3898 -4864
rect -3828 -4996 -3818 -4864
rect -3898 -5002 -3828 -4996
rect -3782 -5034 -3704 -4826
rect -3658 -4864 -3588 -4858
rect -3668 -4996 -3658 -4864
rect -3588 -4996 -3578 -4864
rect -3658 -5002 -3588 -4996
rect -3536 -5034 -3470 -4826
rect -3418 -4864 -3348 -4858
rect -3428 -4996 -3418 -4864
rect -3348 -4996 -3338 -4864
rect -3418 -5002 -3348 -4996
rect -3296 -5034 -3230 -4826
rect -3178 -4864 -3108 -4858
rect -3188 -4996 -3178 -4864
rect -3108 -4996 -3098 -4864
rect -3178 -5002 -3108 -4996
rect -3056 -5034 -2990 -4826
rect -2938 -4864 -2868 -4858
rect -2948 -4996 -2938 -4864
rect -2868 -4996 -2858 -4864
rect -2938 -5002 -2868 -4996
rect -2822 -5034 -2744 -4826
rect -2698 -4864 -2628 -4858
rect -2708 -4996 -2698 -4864
rect -2628 -4996 -2618 -4864
rect -2698 -5002 -2628 -4996
rect -2576 -5034 -2510 -4826
rect -2458 -4864 -2388 -4858
rect -2468 -4996 -2458 -4864
rect -2388 -4996 -2378 -4864
rect -2458 -5002 -2388 -4996
rect -2336 -5034 -2270 -4826
rect -2218 -4864 -2148 -4858
rect -2228 -4996 -2218 -4864
rect -2148 -4996 -2138 -4864
rect -2218 -5002 -2148 -4996
rect -2096 -5034 -2030 -4826
rect -1978 -4864 -1908 -4858
rect -1988 -4996 -1978 -4864
rect -1908 -4996 -1898 -4864
rect -1978 -5002 -1908 -4996
rect -1862 -5034 -1784 -4826
rect -1738 -4864 -1668 -4858
rect -1748 -4996 -1738 -4864
rect -1668 -4996 -1658 -4864
rect -1738 -5002 -1668 -4996
rect -1616 -5034 -1550 -4826
rect -1498 -4864 -1428 -4858
rect -1508 -4996 -1498 -4864
rect -1428 -4996 -1418 -4864
rect -1498 -5002 -1428 -4996
rect -1376 -5034 -1310 -4826
rect -1258 -4864 -1188 -4858
rect -1268 -4996 -1258 -4864
rect -1188 -4996 -1178 -4864
rect -1258 -5002 -1188 -4996
rect -1136 -5034 -1070 -4826
rect -1018 -4864 -948 -4858
rect -1028 -4996 -1018 -4864
rect -948 -4996 -938 -4864
rect -1018 -5002 -948 -4996
rect -902 -5034 -824 -4826
rect -778 -4864 -708 -4858
rect -788 -4996 -778 -4864
rect -708 -4996 -698 -4864
rect -778 -5002 -708 -4996
rect -656 -5034 -590 -4826
rect -538 -4864 -468 -4858
rect -548 -4996 -538 -4864
rect -468 -4996 -458 -4864
rect -538 -5002 -468 -4996
rect -416 -5034 -350 -4826
rect -298 -4864 -228 -4858
rect -308 -4996 -298 -4864
rect -228 -4996 -218 -4864
rect -298 -5002 -228 -4996
rect -176 -5034 -110 -4826
rect -58 -4864 12 -4858
rect -68 -4996 -58 -4864
rect 12 -4996 22 -4864
rect -58 -5002 12 -4996
rect 58 -5034 136 -4826
rect 182 -4864 252 -4858
rect 172 -4996 182 -4864
rect 252 -4996 262 -4864
rect 182 -5002 252 -4996
rect 304 -5034 370 -4826
rect 422 -4864 492 -4858
rect 412 -4996 422 -4864
rect 492 -4996 502 -4864
rect 422 -5002 492 -4996
rect 544 -5034 610 -4826
rect 662 -4864 732 -4858
rect 652 -4996 662 -4864
rect 732 -4996 742 -4864
rect 662 -5002 732 -4996
rect 784 -5034 850 -4826
rect 902 -4864 972 -4858
rect 892 -4996 902 -4864
rect 972 -4996 982 -4864
rect 902 -5002 972 -4996
rect 1018 -5034 1096 -4826
rect 1142 -4864 1212 -4858
rect 1132 -4996 1142 -4864
rect 1212 -4996 1222 -4864
rect 1142 -5002 1212 -4996
rect 1264 -5034 1330 -4826
rect 1382 -4864 1452 -4858
rect 1372 -4996 1382 -4864
rect 1452 -4996 1462 -4864
rect 1382 -5002 1452 -4996
rect 1504 -5034 1570 -4826
rect 1622 -4864 1692 -4858
rect 1612 -4996 1622 -4864
rect 1692 -4996 1702 -4864
rect 1622 -5002 1692 -4996
rect 1744 -5034 1810 -4826
rect 1862 -4864 1932 -4858
rect 1852 -4996 1862 -4864
rect 1932 -4996 1942 -4864
rect 1862 -5002 1932 -4996
rect 1978 -5034 2056 -4826
rect 2102 -4864 2172 -4858
rect 2092 -4996 2102 -4864
rect 2172 -4996 2182 -4864
rect 2102 -5002 2172 -4996
rect 2224 -5034 2290 -4826
rect 2342 -4864 2412 -4858
rect 2332 -4996 2342 -4864
rect 2412 -4996 2422 -4864
rect 2342 -5002 2412 -4996
rect 2464 -5034 2530 -4826
rect 2582 -4864 2652 -4858
rect 2572 -4996 2582 -4864
rect 2652 -4996 2662 -4864
rect 2582 -5002 2652 -4996
rect 2704 -5034 2770 -4826
rect 2822 -4864 2892 -4858
rect 2812 -4996 2822 -4864
rect 2892 -4996 2902 -4864
rect 2822 -5002 2892 -4996
rect 2938 -5034 3016 -4826
rect -6662 -5046 -6544 -5034
rect -6662 -5622 -6584 -5046
rect -6550 -5622 -6544 -5046
rect -6662 -5634 -6544 -5622
rect -6462 -5046 -6304 -5034
rect -6462 -5622 -6456 -5046
rect -6422 -5622 -6344 -5046
rect -6310 -5622 -6304 -5046
rect -6462 -5634 -6304 -5622
rect -6222 -5046 -6064 -5034
rect -6222 -5622 -6216 -5046
rect -6182 -5622 -6104 -5046
rect -6070 -5622 -6064 -5046
rect -6222 -5634 -6064 -5622
rect -5982 -5046 -5824 -5034
rect -5982 -5622 -5976 -5046
rect -5942 -5622 -5864 -5046
rect -5830 -5622 -5824 -5046
rect -5982 -5634 -5824 -5622
rect -5742 -5046 -5584 -5034
rect -5742 -5622 -5736 -5046
rect -5702 -5622 -5624 -5046
rect -5590 -5622 -5584 -5046
rect -5742 -5634 -5584 -5622
rect -5502 -5046 -5344 -5034
rect -5502 -5622 -5496 -5046
rect -5462 -5622 -5384 -5046
rect -5350 -5622 -5344 -5046
rect -5502 -5634 -5344 -5622
rect -5262 -5046 -5104 -5034
rect -5262 -5622 -5256 -5046
rect -5222 -5622 -5144 -5046
rect -5110 -5622 -5104 -5046
rect -5262 -5634 -5104 -5622
rect -5022 -5046 -4864 -5034
rect -5022 -5622 -5016 -5046
rect -4982 -5622 -4904 -5046
rect -4870 -5622 -4864 -5046
rect -5022 -5634 -4864 -5622
rect -4782 -5046 -4624 -5034
rect -4782 -5622 -4776 -5046
rect -4742 -5622 -4664 -5046
rect -4630 -5622 -4624 -5046
rect -4782 -5634 -4624 -5622
rect -4542 -5046 -4384 -5034
rect -4542 -5622 -4536 -5046
rect -4502 -5622 -4424 -5046
rect -4390 -5622 -4384 -5046
rect -4542 -5634 -4384 -5622
rect -4302 -5046 -4144 -5034
rect -4302 -5622 -4296 -5046
rect -4262 -5622 -4184 -5046
rect -4150 -5622 -4144 -5046
rect -4302 -5634 -4144 -5622
rect -4062 -5046 -3904 -5034
rect -4062 -5622 -4056 -5046
rect -4022 -5622 -3944 -5046
rect -3910 -5622 -3904 -5046
rect -4062 -5634 -3904 -5622
rect -3822 -5046 -3664 -5034
rect -3822 -5622 -3816 -5046
rect -3782 -5622 -3704 -5046
rect -3670 -5622 -3664 -5046
rect -3822 -5634 -3664 -5622
rect -3582 -5046 -3424 -5034
rect -3582 -5622 -3576 -5046
rect -3542 -5622 -3464 -5046
rect -3430 -5622 -3424 -5046
rect -3582 -5634 -3424 -5622
rect -3342 -5046 -3184 -5034
rect -3342 -5622 -3336 -5046
rect -3302 -5622 -3224 -5046
rect -3190 -5622 -3184 -5046
rect -3342 -5634 -3184 -5622
rect -3102 -5046 -2944 -5034
rect -3102 -5622 -3096 -5046
rect -3062 -5622 -2984 -5046
rect -2950 -5622 -2944 -5046
rect -3102 -5634 -2944 -5622
rect -2862 -5046 -2704 -5034
rect -2862 -5622 -2856 -5046
rect -2822 -5622 -2744 -5046
rect -2710 -5622 -2704 -5046
rect -2862 -5634 -2704 -5622
rect -2622 -5046 -2464 -5034
rect -2622 -5622 -2616 -5046
rect -2582 -5622 -2504 -5046
rect -2470 -5622 -2464 -5046
rect -2622 -5634 -2464 -5622
rect -2382 -5046 -2224 -5034
rect -2382 -5622 -2376 -5046
rect -2342 -5622 -2264 -5046
rect -2230 -5622 -2224 -5046
rect -2382 -5634 -2224 -5622
rect -2142 -5046 -1984 -5034
rect -2142 -5622 -2136 -5046
rect -2102 -5622 -2024 -5046
rect -1990 -5622 -1984 -5046
rect -2142 -5634 -1984 -5622
rect -1902 -5046 -1744 -5034
rect -1902 -5622 -1896 -5046
rect -1862 -5622 -1784 -5046
rect -1750 -5622 -1744 -5046
rect -1902 -5634 -1744 -5622
rect -1662 -5046 -1504 -5034
rect -1662 -5622 -1656 -5046
rect -1622 -5622 -1544 -5046
rect -1510 -5622 -1504 -5046
rect -1662 -5634 -1504 -5622
rect -1422 -5046 -1264 -5034
rect -1422 -5622 -1416 -5046
rect -1382 -5622 -1304 -5046
rect -1270 -5622 -1264 -5046
rect -1422 -5634 -1264 -5622
rect -1182 -5046 -1024 -5034
rect -1182 -5622 -1176 -5046
rect -1142 -5622 -1064 -5046
rect -1030 -5622 -1024 -5046
rect -1182 -5634 -1024 -5622
rect -942 -5046 -784 -5034
rect -942 -5622 -936 -5046
rect -902 -5622 -824 -5046
rect -790 -5622 -784 -5046
rect -942 -5634 -784 -5622
rect -702 -5046 -544 -5034
rect -702 -5622 -696 -5046
rect -662 -5622 -584 -5046
rect -550 -5622 -544 -5046
rect -702 -5634 -544 -5622
rect -462 -5046 -304 -5034
rect -462 -5622 -456 -5046
rect -422 -5622 -344 -5046
rect -310 -5622 -304 -5046
rect -462 -5634 -304 -5622
rect -222 -5046 -64 -5034
rect -222 -5622 -216 -5046
rect -182 -5622 -104 -5046
rect -70 -5622 -64 -5046
rect -222 -5634 -64 -5622
rect 18 -5046 176 -5034
rect 18 -5622 24 -5046
rect 58 -5622 136 -5046
rect 170 -5622 176 -5046
rect 18 -5634 176 -5622
rect 258 -5046 416 -5034
rect 258 -5622 264 -5046
rect 298 -5622 376 -5046
rect 410 -5622 416 -5046
rect 258 -5634 416 -5622
rect 498 -5046 656 -5034
rect 498 -5622 504 -5046
rect 538 -5622 616 -5046
rect 650 -5622 656 -5046
rect 498 -5634 656 -5622
rect 738 -5046 896 -5034
rect 738 -5622 744 -5046
rect 778 -5622 856 -5046
rect 890 -5622 896 -5046
rect 738 -5634 896 -5622
rect 978 -5046 1136 -5034
rect 978 -5622 984 -5046
rect 1018 -5622 1096 -5046
rect 1130 -5622 1136 -5046
rect 978 -5634 1136 -5622
rect 1218 -5046 1376 -5034
rect 1218 -5622 1224 -5046
rect 1258 -5622 1336 -5046
rect 1370 -5622 1376 -5046
rect 1218 -5634 1376 -5622
rect 1458 -5046 1616 -5034
rect 1458 -5622 1464 -5046
rect 1498 -5622 1576 -5046
rect 1610 -5622 1616 -5046
rect 1458 -5634 1616 -5622
rect 1698 -5046 1856 -5034
rect 1698 -5622 1704 -5046
rect 1738 -5622 1816 -5046
rect 1850 -5622 1856 -5046
rect 1698 -5634 1856 -5622
rect 1938 -5046 2096 -5034
rect 1938 -5622 1944 -5046
rect 1978 -5622 2056 -5046
rect 2090 -5622 2096 -5046
rect 1938 -5634 2096 -5622
rect 2178 -5046 2336 -5034
rect 2178 -5622 2184 -5046
rect 2218 -5622 2296 -5046
rect 2330 -5622 2336 -5046
rect 2178 -5634 2336 -5622
rect 2418 -5046 2576 -5034
rect 2418 -5622 2424 -5046
rect 2458 -5622 2536 -5046
rect 2570 -5622 2576 -5046
rect 2418 -5634 2576 -5622
rect 2658 -5046 2816 -5034
rect 2658 -5622 2664 -5046
rect 2698 -5622 2776 -5046
rect 2810 -5622 2816 -5046
rect 2658 -5634 2816 -5622
rect 2898 -5046 3016 -5034
rect 2898 -5622 2904 -5046
rect 2938 -5622 3016 -5046
rect 2898 -5634 3016 -5622
rect -6662 -6500 -6596 -5634
rect -6538 -5672 -6468 -5666
rect -6298 -5672 -6228 -5666
rect -6548 -5804 -6538 -5672
rect -6468 -5804 -6458 -5672
rect -6308 -5804 -6298 -5672
rect -6228 -5804 -6218 -5672
rect -6538 -5810 -6468 -5804
rect -6298 -5810 -6228 -5804
rect -6170 -6500 -6116 -5634
rect -6058 -5672 -5988 -5666
rect -5818 -5672 -5748 -5666
rect -6068 -5804 -6058 -5672
rect -5988 -5804 -5978 -5672
rect -5828 -5804 -5818 -5672
rect -5748 -5804 -5738 -5672
rect -6058 -5810 -5988 -5804
rect -5818 -5810 -5748 -5804
rect -5690 -6500 -5636 -5634
rect -5578 -5672 -5508 -5666
rect -5338 -5672 -5268 -5666
rect -5588 -5804 -5578 -5672
rect -5508 -5804 -5498 -5672
rect -5348 -5804 -5338 -5672
rect -5268 -5804 -5258 -5672
rect -5578 -5810 -5508 -5804
rect -5338 -5810 -5268 -5804
rect -5210 -6500 -5156 -5634
rect -5098 -5672 -5028 -5666
rect -4858 -5672 -4788 -5666
rect -5108 -5804 -5098 -5672
rect -5028 -5804 -5018 -5672
rect -4868 -5804 -4858 -5672
rect -4788 -5804 -4778 -5672
rect -5098 -5810 -5028 -5804
rect -4858 -5810 -4788 -5804
rect -4730 -6500 -4676 -5634
rect -4618 -5672 -4548 -5666
rect -4378 -5672 -4308 -5666
rect -4628 -5804 -4618 -5672
rect -4548 -5804 -4538 -5672
rect -4388 -5804 -4378 -5672
rect -4308 -5804 -4298 -5672
rect -4618 -5810 -4548 -5804
rect -4378 -5810 -4308 -5804
rect -4250 -6500 -4196 -5634
rect -4138 -5672 -4068 -5666
rect -3898 -5672 -3828 -5666
rect -4148 -5804 -4138 -5672
rect -4068 -5804 -4058 -5672
rect -3908 -5804 -3898 -5672
rect -3828 -5804 -3818 -5672
rect -4138 -5810 -4068 -5804
rect -3898 -5810 -3828 -5804
rect -3770 -6500 -3716 -5634
rect -3658 -5672 -3588 -5666
rect -3418 -5672 -3348 -5666
rect -3668 -5804 -3658 -5672
rect -3588 -5804 -3578 -5672
rect -3428 -5804 -3418 -5672
rect -3348 -5804 -3338 -5672
rect -3658 -5810 -3588 -5804
rect -3418 -5810 -3348 -5804
rect -3290 -6500 -3236 -5634
rect -3178 -5672 -3108 -5666
rect -2938 -5672 -2868 -5666
rect -3188 -5804 -3178 -5672
rect -3108 -5804 -3098 -5672
rect -2948 -5804 -2938 -5672
rect -2868 -5804 -2858 -5672
rect -3178 -5810 -3108 -5804
rect -2938 -5810 -2868 -5804
rect -2810 -6500 -2756 -5634
rect -2698 -5672 -2628 -5666
rect -2458 -5672 -2388 -5666
rect -2708 -5804 -2698 -5672
rect -2628 -5804 -2618 -5672
rect -2468 -5804 -2458 -5672
rect -2388 -5804 -2378 -5672
rect -2698 -5810 -2628 -5804
rect -2458 -5810 -2388 -5804
rect -2330 -6500 -2276 -5634
rect -2218 -5672 -2148 -5666
rect -1978 -5672 -1908 -5666
rect -2228 -5804 -2218 -5672
rect -2148 -5804 -2138 -5672
rect -1988 -5804 -1978 -5672
rect -1908 -5804 -1898 -5672
rect -2218 -5810 -2148 -5804
rect -1978 -5810 -1908 -5804
rect -1850 -6500 -1796 -5634
rect -1738 -5672 -1668 -5666
rect -1498 -5672 -1428 -5666
rect -1748 -5804 -1738 -5672
rect -1668 -5804 -1658 -5672
rect -1508 -5804 -1498 -5672
rect -1428 -5804 -1418 -5672
rect -1738 -5810 -1668 -5804
rect -1498 -5810 -1428 -5804
rect -1370 -6500 -1316 -5634
rect -1258 -5672 -1188 -5666
rect -1018 -5672 -948 -5666
rect -1268 -5804 -1258 -5672
rect -1188 -5804 -1178 -5672
rect -1028 -5804 -1018 -5672
rect -948 -5804 -938 -5672
rect -1258 -5810 -1188 -5804
rect -1018 -5810 -948 -5804
rect -890 -6500 -836 -5634
rect -778 -5672 -708 -5666
rect -538 -5672 -468 -5666
rect -788 -5804 -778 -5672
rect -708 -5804 -698 -5672
rect -548 -5804 -538 -5672
rect -468 -5804 -458 -5672
rect -778 -5810 -708 -5804
rect -538 -5810 -468 -5804
rect -410 -6500 -356 -5634
rect -298 -5672 -228 -5666
rect -58 -5672 12 -5666
rect -308 -5804 -298 -5672
rect -228 -5804 -218 -5672
rect -68 -5804 -58 -5672
rect 12 -5804 22 -5672
rect -298 -5810 -228 -5804
rect -58 -5810 12 -5804
rect 70 -6500 124 -5634
rect 182 -5672 252 -5666
rect 422 -5672 492 -5666
rect 172 -5804 182 -5672
rect 252 -5804 262 -5672
rect 412 -5804 422 -5672
rect 492 -5804 502 -5672
rect 182 -5810 252 -5804
rect 422 -5810 492 -5804
rect 550 -6500 604 -5634
rect 662 -5672 732 -5666
rect 902 -5672 972 -5666
rect 652 -5804 662 -5672
rect 732 -5804 742 -5672
rect 892 -5804 902 -5672
rect 972 -5804 982 -5672
rect 662 -5810 732 -5804
rect 902 -5810 972 -5804
rect 1030 -6500 1084 -5634
rect 1142 -5672 1212 -5666
rect 1382 -5672 1452 -5666
rect 1132 -5804 1142 -5672
rect 1212 -5804 1222 -5672
rect 1372 -5804 1382 -5672
rect 1452 -5804 1462 -5672
rect 1142 -5810 1212 -5804
rect 1382 -5810 1452 -5804
rect 1510 -6500 1564 -5634
rect 1622 -5672 1692 -5666
rect 1862 -5672 1932 -5666
rect 1612 -5804 1622 -5672
rect 1692 -5804 1702 -5672
rect 1852 -5804 1862 -5672
rect 1932 -5804 1942 -5672
rect 1622 -5810 1692 -5804
rect 1862 -5810 1932 -5804
rect 1990 -6500 2044 -5634
rect 2102 -5672 2172 -5666
rect 2342 -5672 2412 -5666
rect 2092 -5804 2102 -5672
rect 2172 -5804 2182 -5672
rect 2332 -5804 2342 -5672
rect 2412 -5804 2422 -5672
rect 2102 -5810 2172 -5804
rect 2342 -5810 2412 -5804
rect 2470 -6500 2524 -5634
rect 2582 -5672 2652 -5666
rect 2822 -5672 2892 -5666
rect 2572 -5804 2582 -5672
rect 2652 -5804 2662 -5672
rect 2812 -5804 2822 -5672
rect 2892 -5804 2902 -5672
rect 2582 -5810 2652 -5804
rect 2822 -5810 2892 -5804
rect 2950 -6500 3016 -5634
rect -15978 -6698 12330 -6500
rect -15978 -7196 7404 -6698
rect 8304 -7196 12330 -6698
rect -15978 -7362 12330 -7196
rect -15978 -8300 -15900 -7362
rect -15838 -8219 -15446 -8213
rect -15838 -8253 -15826 -8219
rect -15458 -8253 -15446 -8219
rect -15838 -8259 -15446 -8253
rect -15250 -8219 -14858 -8213
rect -15250 -8253 -15238 -8219
rect -14870 -8253 -14858 -8219
rect -15250 -8259 -14858 -8253
rect -14796 -8300 -14724 -7362
rect -14662 -8219 -14270 -8213
rect -14662 -8253 -14650 -8219
rect -14282 -8253 -14270 -8219
rect -14662 -8259 -14270 -8253
rect -14074 -8219 -13682 -8213
rect -14074 -8253 -14062 -8219
rect -13694 -8253 -13682 -8219
rect -14074 -8259 -13682 -8253
rect -13620 -8300 -13548 -7362
rect -13486 -8219 -13094 -8213
rect -13486 -8253 -13474 -8219
rect -13106 -8253 -13094 -8219
rect -13486 -8259 -13094 -8253
rect -12898 -8219 -12506 -8213
rect -12898 -8253 -12886 -8219
rect -12518 -8253 -12506 -8219
rect -12898 -8259 -12506 -8253
rect -12444 -8300 -12372 -7362
rect -12310 -8219 -11918 -8213
rect -12310 -8253 -12298 -8219
rect -11930 -8253 -11918 -8219
rect -12310 -8259 -11918 -8253
rect -11722 -8219 -11330 -8213
rect -11722 -8253 -11710 -8219
rect -11342 -8253 -11330 -8219
rect -11722 -8259 -11330 -8253
rect -11268 -8300 -11196 -7362
rect -11134 -8219 -10742 -8213
rect -11134 -8253 -11122 -8219
rect -10754 -8253 -10742 -8219
rect -11134 -8259 -10742 -8253
rect -10546 -8219 -10154 -8213
rect -10546 -8253 -10534 -8219
rect -10166 -8253 -10154 -8219
rect -10546 -8259 -10154 -8253
rect -10092 -8300 -10020 -7362
rect -9958 -8219 -9566 -8213
rect -9958 -8253 -9946 -8219
rect -9578 -8253 -9566 -8219
rect -9958 -8259 -9566 -8253
rect -9370 -8219 -8978 -8213
rect -9370 -8253 -9358 -8219
rect -8990 -8253 -8978 -8219
rect -9370 -8259 -8978 -8253
rect -8916 -8300 -8844 -7362
rect -8782 -8219 -8390 -8213
rect -8782 -8253 -8770 -8219
rect -8402 -8253 -8390 -8219
rect -8782 -8259 -8390 -8253
rect -8194 -8219 -7802 -8213
rect -8194 -8253 -8182 -8219
rect -7814 -8253 -7802 -8219
rect -8194 -8259 -7802 -8253
rect -7740 -8300 -7668 -7362
rect -7606 -8219 -7214 -8213
rect -7606 -8253 -7594 -8219
rect -7226 -8253 -7214 -8219
rect -7606 -8259 -7214 -8253
rect -7018 -8219 -6626 -8213
rect -7018 -8253 -7006 -8219
rect -6638 -8253 -6626 -8219
rect -7018 -8259 -6626 -8253
rect -6564 -8300 -6492 -7362
rect -6430 -8219 -6038 -8213
rect -6430 -8253 -6418 -8219
rect -6050 -8253 -6038 -8219
rect -6430 -8259 -6038 -8253
rect -5842 -8219 -5450 -8213
rect -5842 -8253 -5830 -8219
rect -5462 -8253 -5450 -8219
rect -5842 -8259 -5450 -8253
rect -5388 -8300 -5316 -7362
rect -5254 -8219 -4862 -8213
rect -5254 -8253 -5242 -8219
rect -4874 -8253 -4862 -8219
rect -5254 -8259 -4862 -8253
rect -4666 -8219 -4274 -8213
rect -4666 -8253 -4654 -8219
rect -4286 -8253 -4274 -8219
rect -4666 -8259 -4274 -8253
rect -4240 -8300 -4168 -7362
rect -4078 -8219 -3686 -8213
rect -4078 -8253 -4066 -8219
rect -3698 -8253 -3686 -8219
rect -4078 -8259 -3686 -8253
rect -3490 -8219 -3098 -8213
rect -3490 -8253 -3478 -8219
rect -3110 -8253 -3098 -8219
rect -3490 -8259 -3098 -8253
rect -2902 -8219 -2510 -8213
rect -2902 -8253 -2890 -8219
rect -2522 -8253 -2510 -8219
rect -2902 -8259 -2510 -8253
rect -2314 -8219 -1922 -8213
rect -2314 -8253 -2302 -8219
rect -1934 -8253 -1922 -8219
rect -2314 -8259 -1922 -8253
rect -1726 -8219 -1334 -8213
rect -1726 -8253 -1714 -8219
rect -1346 -8253 -1334 -8219
rect -1726 -8259 -1334 -8253
rect -1138 -8219 -746 -8213
rect -1138 -8253 -1126 -8219
rect -758 -8253 -746 -8219
rect -1138 -8259 -746 -8253
rect -550 -8219 -158 -8213
rect -550 -8253 -538 -8219
rect -170 -8253 -158 -8219
rect -550 -8259 -158 -8253
rect 38 -8219 430 -8213
rect 38 -8253 50 -8219
rect 418 -8253 430 -8219
rect 38 -8259 430 -8253
rect 520 -8300 592 -7362
rect 626 -8219 1018 -8213
rect 626 -8253 638 -8219
rect 1006 -8253 1018 -8219
rect 626 -8259 1018 -8253
rect 1214 -8219 1606 -8213
rect 1214 -8253 1226 -8219
rect 1594 -8253 1606 -8219
rect 1214 -8259 1606 -8253
rect 1668 -8300 1740 -7362
rect 1802 -8219 2194 -8213
rect 1802 -8253 1814 -8219
rect 2182 -8253 2194 -8219
rect 1802 -8259 2194 -8253
rect 2390 -8219 2782 -8213
rect 2390 -8253 2402 -8219
rect 2770 -8253 2782 -8219
rect 2390 -8259 2782 -8253
rect 2844 -8300 2916 -7362
rect 2978 -8219 3370 -8213
rect 2978 -8253 2990 -8219
rect 3358 -8253 3370 -8219
rect 2978 -8259 3370 -8253
rect 3566 -8219 3958 -8213
rect 3566 -8253 3578 -8219
rect 3946 -8253 3958 -8219
rect 3566 -8259 3958 -8253
rect 4020 -8300 4092 -7362
rect 4154 -8219 4546 -8213
rect 4154 -8253 4166 -8219
rect 4534 -8253 4546 -8219
rect 4154 -8259 4546 -8253
rect 4742 -8219 5134 -8213
rect 4742 -8253 4754 -8219
rect 5122 -8253 5134 -8219
rect 4742 -8259 5134 -8253
rect 5196 -8300 5268 -7362
rect 5330 -8219 5722 -8213
rect 5330 -8253 5342 -8219
rect 5710 -8253 5722 -8219
rect 5330 -8259 5722 -8253
rect 5918 -8219 6310 -8213
rect 5918 -8253 5930 -8219
rect 6298 -8253 6310 -8219
rect 5918 -8259 6310 -8253
rect 6372 -8300 6444 -7362
rect 6506 -8219 6898 -8213
rect 6506 -8253 6518 -8219
rect 6886 -8253 6898 -8219
rect 6506 -8259 6898 -8253
rect 7094 -8219 7486 -8213
rect 7094 -8253 7106 -8219
rect 7474 -8253 7486 -8219
rect 7094 -8259 7486 -8253
rect 7548 -8300 7620 -7362
rect 7682 -8219 8074 -8213
rect 7682 -8253 7694 -8219
rect 8062 -8253 8074 -8219
rect 7682 -8259 8074 -8253
rect 8270 -8219 8662 -8213
rect 8270 -8253 8282 -8219
rect 8650 -8253 8662 -8219
rect 8270 -8259 8662 -8253
rect 8724 -8300 8796 -7362
rect 8858 -8219 9250 -8213
rect 8858 -8253 8870 -8219
rect 9238 -8253 9250 -8219
rect 8858 -8259 9250 -8253
rect 9446 -8219 9838 -8213
rect 9446 -8253 9458 -8219
rect 9826 -8253 9838 -8219
rect 9446 -8259 9838 -8253
rect 9900 -8300 9972 -7362
rect 10034 -8219 10426 -8213
rect 10034 -8253 10046 -8219
rect 10414 -8253 10426 -8219
rect 10034 -8259 10426 -8253
rect 10622 -8219 11014 -8213
rect 10622 -8253 10634 -8219
rect 11002 -8253 11014 -8219
rect 10622 -8259 11014 -8253
rect 11076 -8300 11148 -7362
rect 11210 -8219 11602 -8213
rect 11210 -8253 11222 -8219
rect 11590 -8253 11602 -8219
rect 11210 -8259 11602 -8253
rect 11798 -8219 12190 -8213
rect 11798 -8253 11810 -8219
rect 12178 -8253 12190 -8219
rect 11798 -8259 12190 -8253
rect 12252 -8300 12330 -7362
rect -15978 -8312 -15848 -8300
rect -15978 -9088 -15888 -8312
rect -15854 -9088 -15848 -8312
rect -15978 -9100 -15848 -9088
rect -15436 -8312 -15260 -8300
rect -15436 -9088 -15430 -8312
rect -15396 -9088 -15300 -8312
rect -15266 -9088 -15260 -8312
rect -15436 -9100 -15260 -9088
rect -14848 -8312 -14672 -8300
rect -14848 -9088 -14842 -8312
rect -14808 -9088 -14712 -8312
rect -14678 -9088 -14672 -8312
rect -14848 -9100 -14672 -9088
rect -14260 -8312 -14084 -8300
rect -14260 -9088 -14254 -8312
rect -14220 -9088 -14124 -8312
rect -14090 -9088 -14084 -8312
rect -14260 -9100 -14084 -9088
rect -13672 -8312 -13496 -8300
rect -13672 -9088 -13666 -8312
rect -13632 -9088 -13536 -8312
rect -13502 -9088 -13496 -8312
rect -13672 -9100 -13496 -9088
rect -13084 -8312 -12908 -8300
rect -13084 -9088 -13078 -8312
rect -13044 -9088 -12948 -8312
rect -12914 -9088 -12908 -8312
rect -13084 -9100 -12908 -9088
rect -12496 -8312 -12320 -8300
rect -12496 -9088 -12490 -8312
rect -12456 -9088 -12360 -8312
rect -12326 -9088 -12320 -8312
rect -12496 -9100 -12320 -9088
rect -11908 -8312 -11732 -8300
rect -11908 -9088 -11902 -8312
rect -11868 -9088 -11772 -8312
rect -11738 -9088 -11732 -8312
rect -11908 -9100 -11732 -9088
rect -11320 -8312 -11144 -8300
rect -11320 -9088 -11314 -8312
rect -11280 -9088 -11184 -8312
rect -11150 -9088 -11144 -8312
rect -11320 -9100 -11144 -9088
rect -10732 -8312 -10556 -8300
rect -10732 -9088 -10726 -8312
rect -10692 -9088 -10596 -8312
rect -10562 -9088 -10556 -8312
rect -10732 -9100 -10556 -9088
rect -10144 -8312 -9968 -8300
rect -10144 -9088 -10138 -8312
rect -10104 -9088 -10008 -8312
rect -9974 -9088 -9968 -8312
rect -10144 -9100 -9968 -9088
rect -9556 -8312 -9380 -8300
rect -9556 -9088 -9550 -8312
rect -9516 -9088 -9420 -8312
rect -9386 -9088 -9380 -8312
rect -9556 -9100 -9380 -9088
rect -8968 -8312 -8792 -8300
rect -8968 -9088 -8962 -8312
rect -8928 -9088 -8832 -8312
rect -8798 -9088 -8792 -8312
rect -8968 -9100 -8792 -9088
rect -8380 -8312 -8204 -8300
rect -8380 -9088 -8374 -8312
rect -8340 -9088 -8244 -8312
rect -8210 -9088 -8204 -8312
rect -8380 -9100 -8204 -9088
rect -7792 -8312 -7616 -8300
rect -7792 -9088 -7786 -8312
rect -7752 -9088 -7656 -8312
rect -7622 -9088 -7616 -8312
rect -7792 -9100 -7616 -9088
rect -7204 -8312 -7028 -8300
rect -7204 -9088 -7198 -8312
rect -7164 -9088 -7068 -8312
rect -7034 -9088 -7028 -8312
rect -7204 -9100 -7028 -9088
rect -6616 -8312 -6440 -8300
rect -6616 -9088 -6610 -8312
rect -6576 -9088 -6480 -8312
rect -6446 -9088 -6440 -8312
rect -6616 -9100 -6440 -9088
rect -6028 -8312 -5852 -8300
rect -6028 -9088 -6022 -8312
rect -5988 -9088 -5892 -8312
rect -5858 -9088 -5852 -8312
rect -6028 -9100 -5852 -9088
rect -5440 -8312 -5264 -8300
rect -5440 -9088 -5434 -8312
rect -5400 -9088 -5304 -8312
rect -5270 -9088 -5264 -8312
rect -5440 -9100 -5264 -9088
rect -4852 -8312 -4676 -8300
rect -4852 -9088 -4846 -8312
rect -4812 -9088 -4716 -8312
rect -4682 -9088 -4676 -8312
rect -4852 -9100 -4676 -9088
rect -4264 -8312 -4168 -8300
rect -4264 -9088 -4258 -8312
rect -4224 -9036 -4168 -8312
rect -4134 -8312 -4088 -8300
rect -4224 -9088 -4166 -9036
rect -4264 -9100 -4166 -9088
rect -4134 -9088 -4128 -8312
rect -4094 -9088 -4088 -8312
rect -4134 -9100 -4088 -9088
rect -3676 -8312 -3500 -8300
rect -3676 -9088 -3670 -8312
rect -3636 -9088 -3540 -8312
rect -3506 -9088 -3500 -8312
rect -3676 -9100 -3500 -9088
rect -3088 -8312 -2912 -8300
rect -3088 -9088 -3082 -8312
rect -3048 -9088 -2952 -8312
rect -2918 -9088 -2912 -8312
rect -3088 -9100 -2912 -9088
rect -2500 -8312 -2324 -8300
rect -2500 -9088 -2494 -8312
rect -2460 -9088 -2364 -8312
rect -2330 -9088 -2324 -8312
rect -2500 -9100 -2324 -9088
rect -1912 -8312 -1866 -8300
rect -1912 -9088 -1906 -8312
rect -1872 -9088 -1866 -8312
rect -1912 -9100 -1866 -9088
rect -1782 -8312 -1736 -8300
rect -1782 -9088 -1776 -8312
rect -1742 -9088 -1736 -8312
rect -1782 -9100 -1736 -9088
rect -1324 -8312 -1148 -8300
rect -1324 -9088 -1318 -8312
rect -1284 -9088 -1188 -8312
rect -1154 -9088 -1148 -8312
rect -1324 -9100 -1148 -9088
rect -736 -8312 -560 -8300
rect -736 -9088 -730 -8312
rect -696 -9088 -600 -8312
rect -566 -9088 -560 -8312
rect -736 -9100 -560 -9088
rect -148 -8312 28 -8300
rect -148 -9088 -142 -8312
rect -108 -9088 -12 -8312
rect 22 -9088 28 -8312
rect -148 -9100 28 -9088
rect 440 -8312 486 -8300
rect 440 -9088 446 -8312
rect 480 -9088 486 -8312
rect 440 -9100 486 -9088
rect 520 -8312 616 -8300
rect 520 -9088 576 -8312
rect 610 -9088 616 -8312
rect 520 -9100 616 -9088
rect 1028 -8312 1204 -8300
rect 1028 -9088 1034 -8312
rect 1068 -9088 1164 -8312
rect 1198 -9088 1204 -8312
rect 1028 -9100 1204 -9088
rect 1616 -8312 1792 -8300
rect 1616 -9088 1622 -8312
rect 1656 -9088 1752 -8312
rect 1786 -9088 1792 -8312
rect 1616 -9100 1792 -9088
rect 2204 -8312 2380 -8300
rect 2204 -9088 2210 -8312
rect 2244 -9088 2340 -8312
rect 2374 -9088 2380 -8312
rect 2204 -9100 2380 -9088
rect 2792 -8312 2968 -8300
rect 2792 -9088 2798 -8312
rect 2832 -9088 2928 -8312
rect 2962 -9088 2968 -8312
rect 2792 -9100 2968 -9088
rect 3380 -8312 3556 -8300
rect 3380 -9088 3386 -8312
rect 3420 -9088 3516 -8312
rect 3550 -9088 3556 -8312
rect 3380 -9100 3556 -9088
rect 3968 -8312 4144 -8300
rect 3968 -9088 3974 -8312
rect 4008 -9088 4104 -8312
rect 4138 -9088 4144 -8312
rect 3968 -9100 4144 -9088
rect 4556 -8312 4732 -8300
rect 4556 -9088 4562 -8312
rect 4596 -9088 4692 -8312
rect 4726 -9088 4732 -8312
rect 4556 -9100 4732 -9088
rect 5144 -8312 5320 -8300
rect 5144 -9088 5150 -8312
rect 5184 -9088 5280 -8312
rect 5314 -9088 5320 -8312
rect 5144 -9100 5320 -9088
rect 5732 -8312 5908 -8300
rect 5732 -9088 5738 -8312
rect 5772 -9088 5868 -8312
rect 5902 -9088 5908 -8312
rect 5732 -9100 5908 -9088
rect 6320 -8312 6496 -8300
rect 6320 -9088 6326 -8312
rect 6360 -9088 6456 -8312
rect 6490 -9088 6496 -8312
rect 6320 -9100 6496 -9088
rect 6908 -8312 7084 -8300
rect 6908 -9088 6914 -8312
rect 6948 -9088 7044 -8312
rect 7078 -9088 7084 -8312
rect 6908 -9100 7084 -9088
rect 7496 -8312 7672 -8300
rect 7496 -9088 7502 -8312
rect 7536 -9088 7632 -8312
rect 7666 -9088 7672 -8312
rect 7496 -9100 7672 -9088
rect 8084 -8312 8260 -8300
rect 8084 -9088 8090 -8312
rect 8124 -9088 8220 -8312
rect 8254 -9088 8260 -8312
rect 8084 -9100 8260 -9088
rect 8672 -8312 8848 -8300
rect 8672 -9088 8678 -8312
rect 8712 -9088 8808 -8312
rect 8842 -9088 8848 -8312
rect 8672 -9100 8848 -9088
rect 9260 -8312 9436 -8300
rect 9260 -9088 9266 -8312
rect 9300 -9088 9396 -8312
rect 9430 -9088 9436 -8312
rect 9260 -9100 9436 -9088
rect 9848 -8312 10024 -8300
rect 9848 -9088 9854 -8312
rect 9888 -9088 9984 -8312
rect 10018 -9088 10024 -8312
rect 9848 -9100 10024 -9088
rect 10436 -8312 10612 -8300
rect 10436 -9088 10442 -8312
rect 10476 -9088 10572 -8312
rect 10606 -9088 10612 -8312
rect 10436 -9100 10612 -9088
rect 11024 -8312 11200 -8300
rect 11024 -9088 11030 -8312
rect 11064 -9088 11160 -8312
rect 11194 -9088 11200 -8312
rect 11024 -9100 11200 -9088
rect 11612 -8312 11788 -8300
rect 11612 -9088 11618 -8312
rect 11652 -9088 11748 -8312
rect 11782 -9088 11788 -8312
rect 11612 -9100 11788 -9088
rect 12200 -8312 12330 -8300
rect 12200 -9088 12206 -8312
rect 12240 -9088 12330 -8312
rect 12200 -9100 12330 -9088
rect -15978 -9300 -15894 -9100
rect -15838 -9147 -15446 -9141
rect -15838 -9181 -15826 -9147
rect -15458 -9181 -15446 -9147
rect -15838 -9219 -15446 -9181
rect -15838 -9253 -15826 -9219
rect -15458 -9253 -15446 -9219
rect -15838 -9259 -15446 -9253
rect -15390 -9300 -15306 -9100
rect -15250 -9147 -14858 -9141
rect -15250 -9181 -15238 -9147
rect -14870 -9181 -14858 -9147
rect -15250 -9219 -14858 -9181
rect -15250 -9253 -15238 -9219
rect -14870 -9253 -14858 -9219
rect -15250 -9259 -14858 -9253
rect -14802 -9300 -14718 -9100
rect -14662 -9147 -14270 -9141
rect -14662 -9181 -14650 -9147
rect -14282 -9181 -14270 -9147
rect -14662 -9219 -14270 -9181
rect -14662 -9253 -14650 -9219
rect -14282 -9253 -14270 -9219
rect -14662 -9259 -14270 -9253
rect -14214 -9300 -14130 -9100
rect -14074 -9147 -13682 -9141
rect -14074 -9181 -14062 -9147
rect -13694 -9181 -13682 -9147
rect -14074 -9219 -13682 -9181
rect -14074 -9253 -14062 -9219
rect -13694 -9253 -13682 -9219
rect -14074 -9259 -13682 -9253
rect -13626 -9300 -13542 -9100
rect -13486 -9147 -13094 -9141
rect -13486 -9181 -13474 -9147
rect -13106 -9181 -13094 -9147
rect -13486 -9219 -13094 -9181
rect -13486 -9253 -13474 -9219
rect -13106 -9253 -13094 -9219
rect -13486 -9259 -13094 -9253
rect -13038 -9300 -12954 -9100
rect -12898 -9147 -12506 -9141
rect -12898 -9181 -12886 -9147
rect -12518 -9181 -12506 -9147
rect -12898 -9219 -12506 -9181
rect -12898 -9253 -12886 -9219
rect -12518 -9253 -12506 -9219
rect -12898 -9259 -12506 -9253
rect -12450 -9300 -12366 -9100
rect -12310 -9147 -11918 -9141
rect -12310 -9181 -12298 -9147
rect -11930 -9181 -11918 -9147
rect -12310 -9219 -11918 -9181
rect -12310 -9253 -12298 -9219
rect -11930 -9253 -11918 -9219
rect -12310 -9259 -11918 -9253
rect -11862 -9300 -11778 -9100
rect -11722 -9147 -11330 -9141
rect -11722 -9181 -11710 -9147
rect -11342 -9181 -11330 -9147
rect -11722 -9219 -11330 -9181
rect -11722 -9253 -11710 -9219
rect -11342 -9253 -11330 -9219
rect -11722 -9259 -11330 -9253
rect -11274 -9300 -11190 -9100
rect -11134 -9147 -10742 -9141
rect -11134 -9181 -11122 -9147
rect -10754 -9181 -10742 -9147
rect -11134 -9219 -10742 -9181
rect -11134 -9253 -11122 -9219
rect -10754 -9253 -10742 -9219
rect -11134 -9259 -10742 -9253
rect -10686 -9300 -10602 -9100
rect -10546 -9147 -10154 -9141
rect -10546 -9181 -10534 -9147
rect -10166 -9181 -10154 -9147
rect -10546 -9219 -10154 -9181
rect -10546 -9253 -10534 -9219
rect -10166 -9253 -10154 -9219
rect -10546 -9259 -10154 -9253
rect -10098 -9300 -10014 -9100
rect -9958 -9147 -9566 -9141
rect -9958 -9181 -9946 -9147
rect -9578 -9181 -9566 -9147
rect -9958 -9219 -9566 -9181
rect -9958 -9253 -9946 -9219
rect -9578 -9253 -9566 -9219
rect -9958 -9259 -9566 -9253
rect -9510 -9300 -9426 -9100
rect -9370 -9147 -8978 -9141
rect -9370 -9181 -9358 -9147
rect -8990 -9181 -8978 -9147
rect -9370 -9219 -8978 -9181
rect -9370 -9253 -9358 -9219
rect -8990 -9253 -8978 -9219
rect -9370 -9259 -8978 -9253
rect -8922 -9300 -8838 -9100
rect -8782 -9147 -8390 -9141
rect -8782 -9181 -8770 -9147
rect -8402 -9181 -8390 -9147
rect -8782 -9219 -8390 -9181
rect -8782 -9253 -8770 -9219
rect -8402 -9253 -8390 -9219
rect -8782 -9259 -8390 -9253
rect -8334 -9300 -8250 -9100
rect -8194 -9147 -7802 -9141
rect -8194 -9181 -8182 -9147
rect -7814 -9181 -7802 -9147
rect -8194 -9219 -7802 -9181
rect -8194 -9253 -8182 -9219
rect -7814 -9253 -7802 -9219
rect -8194 -9259 -7802 -9253
rect -7746 -9300 -7662 -9100
rect -7606 -9147 -7214 -9141
rect -7606 -9181 -7594 -9147
rect -7226 -9181 -7214 -9147
rect -7606 -9219 -7214 -9181
rect -7606 -9253 -7594 -9219
rect -7226 -9253 -7214 -9219
rect -7606 -9259 -7214 -9253
rect -7158 -9300 -7074 -9100
rect -7018 -9147 -6626 -9141
rect -7018 -9181 -7006 -9147
rect -6638 -9181 -6626 -9147
rect -7018 -9219 -6626 -9181
rect -7018 -9253 -7006 -9219
rect -6638 -9253 -6626 -9219
rect -7018 -9259 -6626 -9253
rect -6570 -9300 -6486 -9100
rect -6430 -9147 -6038 -9141
rect -6430 -9181 -6418 -9147
rect -6050 -9181 -6038 -9147
rect -6430 -9219 -6038 -9181
rect -6430 -9253 -6418 -9219
rect -6050 -9253 -6038 -9219
rect -6430 -9259 -6038 -9253
rect -5982 -9300 -5898 -9100
rect -5842 -9147 -5450 -9141
rect -5842 -9181 -5830 -9147
rect -5462 -9181 -5450 -9147
rect -5842 -9219 -5450 -9181
rect -5842 -9253 -5830 -9219
rect -5462 -9253 -5450 -9219
rect -5842 -9259 -5450 -9253
rect -5394 -9300 -5310 -9100
rect -5254 -9147 -4862 -9141
rect -5254 -9181 -5242 -9147
rect -4874 -9181 -4862 -9147
rect -5254 -9219 -4862 -9181
rect -5254 -9253 -5242 -9219
rect -4874 -9253 -4862 -9219
rect -5254 -9259 -4862 -9253
rect -4806 -9300 -4722 -9100
rect -4666 -9147 -4274 -9141
rect -4666 -9181 -4654 -9147
rect -4286 -9181 -4274 -9147
rect -4666 -9219 -4274 -9181
rect -4666 -9253 -4654 -9219
rect -4286 -9253 -4274 -9219
rect -4666 -9259 -4274 -9253
rect -4224 -9300 -4166 -9100
rect -4078 -9147 -3686 -9141
rect -4078 -9181 -4066 -9147
rect -3698 -9181 -3686 -9147
rect -4078 -9219 -3686 -9181
rect -4078 -9253 -4066 -9219
rect -3698 -9253 -3686 -9219
rect -4078 -9259 -3686 -9253
rect -3630 -9300 -3546 -9100
rect -3490 -9147 -3098 -9141
rect -3490 -9181 -3478 -9147
rect -3110 -9181 -3098 -9147
rect -3490 -9219 -3098 -9181
rect -3490 -9253 -3478 -9219
rect -3110 -9253 -3098 -9219
rect -3490 -9259 -3098 -9253
rect -3042 -9300 -2958 -9100
rect -2902 -9147 -2510 -9141
rect -2902 -9181 -2890 -9147
rect -2522 -9181 -2510 -9147
rect -2902 -9219 -2510 -9181
rect -2902 -9253 -2890 -9219
rect -2522 -9253 -2510 -9219
rect -2902 -9259 -2510 -9253
rect -2454 -9300 -2370 -9100
rect -2314 -9147 -1922 -9141
rect -2314 -9181 -2302 -9147
rect -1934 -9181 -1922 -9147
rect -2314 -9219 -1922 -9181
rect -2314 -9253 -2302 -9219
rect -1934 -9253 -1922 -9219
rect -2314 -9259 -1922 -9253
rect -1726 -9147 -1334 -9141
rect -1726 -9181 -1714 -9147
rect -1346 -9181 -1334 -9147
rect -1726 -9219 -1334 -9181
rect -1726 -9253 -1714 -9219
rect -1346 -9253 -1334 -9219
rect -1726 -9259 -1334 -9253
rect -1278 -9300 -1194 -9100
rect -1138 -9147 -746 -9141
rect -1138 -9181 -1126 -9147
rect -758 -9181 -746 -9147
rect -1138 -9219 -746 -9181
rect -1138 -9253 -1126 -9219
rect -758 -9253 -746 -9219
rect -1138 -9259 -746 -9253
rect -690 -9300 -606 -9100
rect -550 -9147 -158 -9141
rect -550 -9181 -538 -9147
rect -170 -9181 -158 -9147
rect -550 -9219 -158 -9181
rect -550 -9253 -538 -9219
rect -170 -9253 -158 -9219
rect -550 -9259 -158 -9253
rect -102 -9300 -18 -9100
rect 38 -9147 430 -9141
rect 38 -9181 50 -9147
rect 418 -9181 430 -9147
rect 38 -9219 430 -9181
rect 38 -9253 50 -9219
rect 418 -9253 430 -9219
rect 38 -9259 430 -9253
rect 520 -9300 576 -9100
rect 626 -9147 1018 -9141
rect 626 -9181 638 -9147
rect 1006 -9181 1018 -9147
rect 626 -9219 1018 -9181
rect 626 -9253 638 -9219
rect 1006 -9253 1018 -9219
rect 626 -9259 1018 -9253
rect 1074 -9300 1158 -9100
rect 1214 -9147 1606 -9141
rect 1214 -9181 1226 -9147
rect 1594 -9181 1606 -9147
rect 1214 -9219 1606 -9181
rect 1214 -9253 1226 -9219
rect 1594 -9253 1606 -9219
rect 1214 -9259 1606 -9253
rect 1662 -9300 1746 -9100
rect 1802 -9147 2194 -9141
rect 1802 -9181 1814 -9147
rect 2182 -9181 2194 -9147
rect 1802 -9219 2194 -9181
rect 1802 -9253 1814 -9219
rect 2182 -9253 2194 -9219
rect 1802 -9259 2194 -9253
rect 2250 -9300 2334 -9100
rect 2390 -9147 2782 -9141
rect 2390 -9181 2402 -9147
rect 2770 -9181 2782 -9147
rect 2390 -9219 2782 -9181
rect 2390 -9253 2402 -9219
rect 2770 -9253 2782 -9219
rect 2390 -9259 2782 -9253
rect 2838 -9300 2922 -9100
rect 2978 -9147 3370 -9141
rect 2978 -9181 2990 -9147
rect 3358 -9181 3370 -9147
rect 2978 -9219 3370 -9181
rect 2978 -9253 2990 -9219
rect 3358 -9253 3370 -9219
rect 2978 -9259 3370 -9253
rect 3426 -9300 3510 -9100
rect 3566 -9147 3958 -9141
rect 3566 -9181 3578 -9147
rect 3946 -9181 3958 -9147
rect 3566 -9219 3958 -9181
rect 3566 -9253 3578 -9219
rect 3946 -9253 3958 -9219
rect 3566 -9259 3958 -9253
rect 4014 -9300 4098 -9100
rect 4154 -9147 4546 -9141
rect 4154 -9181 4166 -9147
rect 4534 -9181 4546 -9147
rect 4154 -9219 4546 -9181
rect 4154 -9253 4166 -9219
rect 4534 -9253 4546 -9219
rect 4154 -9259 4546 -9253
rect 4602 -9300 4686 -9100
rect 4742 -9147 5134 -9141
rect 4742 -9181 4754 -9147
rect 5122 -9181 5134 -9147
rect 4742 -9219 5134 -9181
rect 4742 -9253 4754 -9219
rect 5122 -9253 5134 -9219
rect 4742 -9259 5134 -9253
rect 5190 -9300 5274 -9100
rect 5330 -9147 5722 -9141
rect 5330 -9181 5342 -9147
rect 5710 -9181 5722 -9147
rect 5330 -9219 5722 -9181
rect 5330 -9253 5342 -9219
rect 5710 -9253 5722 -9219
rect 5330 -9259 5722 -9253
rect 5778 -9300 5862 -9100
rect 5918 -9147 6310 -9141
rect 5918 -9181 5930 -9147
rect 6298 -9181 6310 -9147
rect 5918 -9219 6310 -9181
rect 5918 -9253 5930 -9219
rect 6298 -9253 6310 -9219
rect 5918 -9259 6310 -9253
rect 6366 -9300 6450 -9100
rect 6506 -9147 6898 -9141
rect 6506 -9181 6518 -9147
rect 6886 -9181 6898 -9147
rect 6506 -9219 6898 -9181
rect 6506 -9253 6518 -9219
rect 6886 -9253 6898 -9219
rect 6506 -9259 6898 -9253
rect 6954 -9300 7038 -9100
rect 7094 -9147 7486 -9141
rect 7094 -9181 7106 -9147
rect 7474 -9181 7486 -9147
rect 7094 -9219 7486 -9181
rect 7094 -9253 7106 -9219
rect 7474 -9253 7486 -9219
rect 7094 -9259 7486 -9253
rect 7542 -9300 7626 -9100
rect 7682 -9147 8074 -9141
rect 7682 -9181 7694 -9147
rect 8062 -9181 8074 -9147
rect 7682 -9219 8074 -9181
rect 7682 -9253 7694 -9219
rect 8062 -9253 8074 -9219
rect 7682 -9259 8074 -9253
rect 8130 -9300 8214 -9100
rect 8270 -9147 8662 -9141
rect 8270 -9181 8282 -9147
rect 8650 -9181 8662 -9147
rect 8270 -9219 8662 -9181
rect 8270 -9253 8282 -9219
rect 8650 -9253 8662 -9219
rect 8270 -9259 8662 -9253
rect 8718 -9300 8802 -9100
rect 8858 -9147 9250 -9141
rect 8858 -9181 8870 -9147
rect 9238 -9181 9250 -9147
rect 8858 -9219 9250 -9181
rect 8858 -9253 8870 -9219
rect 9238 -9253 9250 -9219
rect 8858 -9259 9250 -9253
rect 9306 -9300 9390 -9100
rect 9446 -9147 9838 -9141
rect 9446 -9181 9458 -9147
rect 9826 -9181 9838 -9147
rect 9446 -9219 9838 -9181
rect 9446 -9253 9458 -9219
rect 9826 -9253 9838 -9219
rect 9446 -9259 9838 -9253
rect 9894 -9300 9978 -9100
rect 10034 -9147 10426 -9141
rect 10034 -9181 10046 -9147
rect 10414 -9181 10426 -9147
rect 10034 -9219 10426 -9181
rect 10034 -9253 10046 -9219
rect 10414 -9253 10426 -9219
rect 10034 -9259 10426 -9253
rect 10482 -9300 10566 -9100
rect 10622 -9147 11014 -9141
rect 10622 -9181 10634 -9147
rect 11002 -9181 11014 -9147
rect 10622 -9219 11014 -9181
rect 10622 -9253 10634 -9219
rect 11002 -9253 11014 -9219
rect 10622 -9259 11014 -9253
rect 11070 -9300 11154 -9100
rect 11210 -9147 11602 -9141
rect 11210 -9181 11222 -9147
rect 11590 -9181 11602 -9147
rect 11210 -9219 11602 -9181
rect 11210 -9253 11222 -9219
rect 11590 -9253 11602 -9219
rect 11210 -9259 11602 -9253
rect 11658 -9300 11742 -9100
rect 11798 -9147 12190 -9141
rect 11798 -9181 11810 -9147
rect 12178 -9181 12190 -9147
rect 11798 -9219 12190 -9181
rect 11798 -9253 11810 -9219
rect 12178 -9253 12190 -9219
rect 11798 -9259 12190 -9253
rect 12246 -9300 12330 -9100
rect -15978 -9312 -15848 -9300
rect -15978 -10088 -15888 -9312
rect -15854 -10088 -15848 -9312
rect -15978 -10100 -15848 -10088
rect -15436 -9312 -15260 -9300
rect -15436 -10088 -15430 -9312
rect -15396 -10088 -15300 -9312
rect -15266 -10088 -15260 -9312
rect -15436 -10100 -15260 -10088
rect -14848 -9312 -14672 -9300
rect -14848 -10088 -14842 -9312
rect -14808 -10088 -14712 -9312
rect -14678 -10088 -14672 -9312
rect -14848 -10100 -14672 -10088
rect -14260 -9312 -14084 -9300
rect -14260 -10088 -14254 -9312
rect -14220 -10088 -14124 -9312
rect -14090 -10088 -14084 -9312
rect -14260 -10100 -14084 -10088
rect -13672 -9312 -13496 -9300
rect -13672 -10088 -13666 -9312
rect -13632 -10088 -13536 -9312
rect -13502 -10088 -13496 -9312
rect -13672 -10100 -13496 -10088
rect -13084 -9312 -12908 -9300
rect -13084 -10088 -13078 -9312
rect -13044 -10088 -12948 -9312
rect -12914 -10088 -12908 -9312
rect -13084 -10100 -12908 -10088
rect -12496 -9312 -12320 -9300
rect -12496 -10088 -12490 -9312
rect -12456 -10088 -12360 -9312
rect -12326 -10088 -12320 -9312
rect -12496 -10100 -12320 -10088
rect -11908 -9312 -11732 -9300
rect -11908 -10088 -11902 -9312
rect -11868 -10088 -11772 -9312
rect -11738 -10088 -11732 -9312
rect -11908 -10100 -11732 -10088
rect -11320 -9312 -11144 -9300
rect -11320 -10088 -11314 -9312
rect -11280 -10088 -11184 -9312
rect -11150 -10088 -11144 -9312
rect -11320 -10100 -11144 -10088
rect -10732 -9312 -10556 -9300
rect -10732 -10088 -10726 -9312
rect -10692 -10088 -10596 -9312
rect -10562 -10088 -10556 -9312
rect -10732 -10100 -10556 -10088
rect -10144 -9312 -9968 -9300
rect -10144 -10088 -10138 -9312
rect -10104 -10088 -10008 -9312
rect -9974 -10088 -9968 -9312
rect -10144 -10100 -9968 -10088
rect -9556 -9312 -9380 -9300
rect -9556 -10088 -9550 -9312
rect -9516 -10088 -9420 -9312
rect -9386 -10088 -9380 -9312
rect -9556 -10100 -9380 -10088
rect -8968 -9312 -8792 -9300
rect -8968 -10088 -8962 -9312
rect -8928 -10088 -8832 -9312
rect -8798 -10088 -8792 -9312
rect -8968 -10100 -8792 -10088
rect -8380 -9312 -8204 -9300
rect -8380 -10088 -8374 -9312
rect -8340 -10088 -8244 -9312
rect -8210 -10088 -8204 -9312
rect -8380 -10100 -8204 -10088
rect -7792 -9312 -7616 -9300
rect -7792 -10088 -7786 -9312
rect -7752 -10088 -7656 -9312
rect -7622 -10088 -7616 -9312
rect -7792 -10100 -7616 -10088
rect -7204 -9312 -7028 -9300
rect -7204 -10088 -7198 -9312
rect -7164 -10088 -7068 -9312
rect -7034 -10088 -7028 -9312
rect -7204 -10100 -7028 -10088
rect -6616 -9312 -6440 -9300
rect -6616 -10088 -6610 -9312
rect -6576 -10088 -6480 -9312
rect -6446 -10088 -6440 -9312
rect -6616 -10100 -6440 -10088
rect -6028 -9312 -5852 -9300
rect -6028 -10088 -6022 -9312
rect -5988 -10088 -5892 -9312
rect -5858 -10088 -5852 -9312
rect -6028 -10100 -5852 -10088
rect -5440 -9312 -5264 -9300
rect -5440 -10088 -5434 -9312
rect -5400 -10088 -5304 -9312
rect -5270 -10088 -5264 -9312
rect -5440 -10100 -5264 -10088
rect -4852 -9312 -4676 -9300
rect -4852 -10088 -4846 -9312
rect -4812 -10088 -4716 -9312
rect -4682 -10088 -4676 -9312
rect -4852 -10100 -4676 -10088
rect -4264 -9312 -4166 -9300
rect -4264 -10088 -4258 -9312
rect -4224 -10088 -4166 -9312
rect -4264 -10100 -4166 -10088
rect -4134 -9312 -4088 -9300
rect -4134 -10088 -4128 -9312
rect -4094 -10088 -4088 -9312
rect -4134 -10100 -4088 -10088
rect -3676 -9312 -3500 -9300
rect -3676 -10088 -3670 -9312
rect -3636 -10088 -3540 -9312
rect -3506 -10088 -3500 -9312
rect -3676 -10100 -3500 -10088
rect -3088 -9312 -2912 -9300
rect -3088 -10088 -3082 -9312
rect -3048 -10088 -2952 -9312
rect -2918 -10088 -2912 -9312
rect -3088 -10100 -2912 -10088
rect -2500 -9312 -2324 -9300
rect -2500 -10088 -2494 -9312
rect -2460 -10088 -2364 -9312
rect -2330 -10088 -2324 -9312
rect -2500 -10100 -2324 -10088
rect -1912 -9312 -1866 -9300
rect -1912 -10088 -1906 -9312
rect -1872 -10088 -1866 -9312
rect -1912 -10100 -1866 -10088
rect -1782 -9312 -1736 -9300
rect -1782 -10088 -1776 -9312
rect -1742 -10088 -1736 -9312
rect -1782 -10100 -1736 -10088
rect -1324 -9312 -1148 -9300
rect -1324 -10088 -1318 -9312
rect -1284 -10088 -1188 -9312
rect -1154 -10088 -1148 -9312
rect -1324 -10100 -1148 -10088
rect -736 -9312 -560 -9300
rect -736 -10088 -730 -9312
rect -696 -10088 -600 -9312
rect -566 -10088 -560 -9312
rect -736 -10100 -560 -10088
rect -148 -9312 28 -9300
rect -148 -10088 -142 -9312
rect -108 -10088 -12 -9312
rect 22 -10088 28 -9312
rect -148 -10100 28 -10088
rect 440 -9312 486 -9300
rect 440 -10088 446 -9312
rect 480 -10088 486 -9312
rect 440 -10100 486 -10088
rect 520 -9312 616 -9300
rect 520 -10088 576 -9312
rect 610 -10088 616 -9312
rect 520 -10100 616 -10088
rect 1028 -9312 1204 -9300
rect 1028 -10088 1034 -9312
rect 1068 -10088 1164 -9312
rect 1198 -10088 1204 -9312
rect 1028 -10100 1204 -10088
rect 1616 -9312 1792 -9300
rect 1616 -10088 1622 -9312
rect 1656 -10088 1752 -9312
rect 1786 -10088 1792 -9312
rect 1616 -10100 1792 -10088
rect 2204 -9312 2380 -9300
rect 2204 -10088 2210 -9312
rect 2244 -10088 2340 -9312
rect 2374 -10088 2380 -9312
rect 2204 -10100 2380 -10088
rect 2792 -9312 2968 -9300
rect 2792 -10088 2798 -9312
rect 2832 -10088 2928 -9312
rect 2962 -10088 2968 -9312
rect 2792 -10100 2968 -10088
rect 3380 -9312 3556 -9300
rect 3380 -10088 3386 -9312
rect 3420 -10088 3516 -9312
rect 3550 -10088 3556 -9312
rect 3380 -10100 3556 -10088
rect 3968 -9312 4144 -9300
rect 3968 -10088 3974 -9312
rect 4008 -10088 4104 -9312
rect 4138 -10088 4144 -9312
rect 3968 -10100 4144 -10088
rect 4556 -9312 4732 -9300
rect 4556 -10088 4562 -9312
rect 4596 -10088 4692 -9312
rect 4726 -10088 4732 -9312
rect 4556 -10100 4732 -10088
rect 5144 -9312 5320 -9300
rect 5144 -10088 5150 -9312
rect 5184 -10088 5280 -9312
rect 5314 -10088 5320 -9312
rect 5144 -10100 5320 -10088
rect 5732 -9312 5908 -9300
rect 5732 -10088 5738 -9312
rect 5772 -10088 5868 -9312
rect 5902 -10088 5908 -9312
rect 5732 -10100 5908 -10088
rect 6320 -9312 6496 -9300
rect 6320 -10088 6326 -9312
rect 6360 -10088 6456 -9312
rect 6490 -10088 6496 -9312
rect 6320 -10100 6496 -10088
rect 6908 -9312 7084 -9300
rect 6908 -10088 6914 -9312
rect 6948 -10088 7044 -9312
rect 7078 -10088 7084 -9312
rect 6908 -10100 7084 -10088
rect 7496 -9312 7672 -9300
rect 7496 -10088 7502 -9312
rect 7536 -10088 7632 -9312
rect 7666 -10088 7672 -9312
rect 7496 -10100 7672 -10088
rect 8084 -9312 8260 -9300
rect 8084 -10088 8090 -9312
rect 8124 -10088 8220 -9312
rect 8254 -10088 8260 -9312
rect 8084 -10100 8260 -10088
rect 8672 -9312 8848 -9300
rect 8672 -10088 8678 -9312
rect 8712 -10088 8808 -9312
rect 8842 -10088 8848 -9312
rect 8672 -10100 8848 -10088
rect 9260 -9312 9436 -9300
rect 9260 -10088 9266 -9312
rect 9300 -10088 9396 -9312
rect 9430 -10088 9436 -9312
rect 9260 -10100 9436 -10088
rect 9848 -9312 10024 -9300
rect 9848 -10088 9854 -9312
rect 9888 -10088 9984 -9312
rect 10018 -10088 10024 -9312
rect 9848 -10100 10024 -10088
rect 10436 -9312 10612 -9300
rect 10436 -10088 10442 -9312
rect 10476 -10088 10572 -9312
rect 10606 -10088 10612 -9312
rect 10436 -10100 10612 -10088
rect 11024 -9312 11200 -9300
rect 11024 -10088 11030 -9312
rect 11064 -10088 11160 -9312
rect 11194 -10088 11200 -9312
rect 11024 -10100 11200 -10088
rect 11612 -9312 11788 -9300
rect 11612 -10088 11618 -9312
rect 11652 -10088 11748 -9312
rect 11782 -10088 11788 -9312
rect 11612 -10100 11788 -10088
rect 12200 -9312 12330 -9300
rect 12200 -10088 12206 -9312
rect 12240 -10088 12330 -9312
rect 12200 -10100 12330 -10088
rect -15978 -10300 -15894 -10100
rect -15838 -10147 -15446 -10141
rect -15838 -10181 -15826 -10147
rect -15458 -10181 -15446 -10147
rect -15838 -10219 -15446 -10181
rect -15838 -10253 -15826 -10219
rect -15458 -10253 -15446 -10219
rect -15838 -10259 -15446 -10253
rect -15390 -10300 -15306 -10100
rect -15250 -10147 -14858 -10141
rect -15250 -10181 -15238 -10147
rect -14870 -10181 -14858 -10147
rect -15250 -10219 -14858 -10181
rect -15250 -10253 -15238 -10219
rect -14870 -10253 -14858 -10219
rect -15250 -10259 -14858 -10253
rect -14802 -10300 -14718 -10100
rect -14662 -10147 -14270 -10141
rect -14662 -10181 -14650 -10147
rect -14282 -10181 -14270 -10147
rect -14662 -10219 -14270 -10181
rect -14662 -10253 -14650 -10219
rect -14282 -10253 -14270 -10219
rect -14662 -10259 -14270 -10253
rect -14214 -10300 -14130 -10100
rect -14074 -10147 -13682 -10141
rect -14074 -10181 -14062 -10147
rect -13694 -10181 -13682 -10147
rect -14074 -10219 -13682 -10181
rect -14074 -10253 -14062 -10219
rect -13694 -10253 -13682 -10219
rect -14074 -10259 -13682 -10253
rect -13626 -10300 -13542 -10100
rect -13486 -10147 -13094 -10141
rect -13486 -10181 -13474 -10147
rect -13106 -10181 -13094 -10147
rect -13486 -10219 -13094 -10181
rect -13486 -10253 -13474 -10219
rect -13106 -10253 -13094 -10219
rect -13486 -10259 -13094 -10253
rect -13038 -10300 -12954 -10100
rect -12898 -10147 -12506 -10141
rect -12898 -10181 -12886 -10147
rect -12518 -10181 -12506 -10147
rect -12898 -10219 -12506 -10181
rect -12898 -10253 -12886 -10219
rect -12518 -10253 -12506 -10219
rect -12898 -10259 -12506 -10253
rect -12450 -10300 -12366 -10100
rect -12310 -10147 -11918 -10141
rect -12310 -10181 -12298 -10147
rect -11930 -10181 -11918 -10147
rect -12310 -10219 -11918 -10181
rect -12310 -10253 -12298 -10219
rect -11930 -10253 -11918 -10219
rect -12310 -10259 -11918 -10253
rect -11862 -10300 -11778 -10100
rect -11722 -10147 -11330 -10141
rect -11722 -10181 -11710 -10147
rect -11342 -10181 -11330 -10147
rect -11722 -10219 -11330 -10181
rect -11722 -10253 -11710 -10219
rect -11342 -10253 -11330 -10219
rect -11722 -10259 -11330 -10253
rect -11274 -10300 -11190 -10100
rect -11134 -10147 -10742 -10141
rect -11134 -10181 -11122 -10147
rect -10754 -10181 -10742 -10147
rect -11134 -10219 -10742 -10181
rect -11134 -10253 -11122 -10219
rect -10754 -10253 -10742 -10219
rect -11134 -10259 -10742 -10253
rect -10686 -10300 -10602 -10100
rect -10546 -10147 -10154 -10141
rect -10546 -10181 -10534 -10147
rect -10166 -10181 -10154 -10147
rect -10546 -10219 -10154 -10181
rect -10546 -10253 -10534 -10219
rect -10166 -10253 -10154 -10219
rect -10546 -10259 -10154 -10253
rect -10098 -10300 -10014 -10100
rect -9958 -10147 -9566 -10141
rect -9958 -10181 -9946 -10147
rect -9578 -10181 -9566 -10147
rect -9958 -10219 -9566 -10181
rect -9958 -10253 -9946 -10219
rect -9578 -10253 -9566 -10219
rect -9958 -10259 -9566 -10253
rect -9510 -10300 -9426 -10100
rect -9370 -10147 -8978 -10141
rect -9370 -10181 -9358 -10147
rect -8990 -10181 -8978 -10147
rect -9370 -10219 -8978 -10181
rect -9370 -10253 -9358 -10219
rect -8990 -10253 -8978 -10219
rect -9370 -10259 -8978 -10253
rect -8922 -10300 -8838 -10100
rect -8782 -10147 -8390 -10141
rect -8782 -10181 -8770 -10147
rect -8402 -10181 -8390 -10147
rect -8782 -10219 -8390 -10181
rect -8782 -10253 -8770 -10219
rect -8402 -10253 -8390 -10219
rect -8782 -10259 -8390 -10253
rect -8334 -10300 -8250 -10100
rect -8194 -10147 -7802 -10141
rect -8194 -10181 -8182 -10147
rect -7814 -10181 -7802 -10147
rect -8194 -10219 -7802 -10181
rect -8194 -10253 -8182 -10219
rect -7814 -10253 -7802 -10219
rect -8194 -10259 -7802 -10253
rect -7746 -10300 -7662 -10100
rect -7606 -10147 -7214 -10141
rect -7606 -10181 -7594 -10147
rect -7226 -10181 -7214 -10147
rect -7606 -10219 -7214 -10181
rect -7606 -10253 -7594 -10219
rect -7226 -10253 -7214 -10219
rect -7606 -10259 -7214 -10253
rect -7158 -10300 -7074 -10100
rect -7018 -10147 -6626 -10141
rect -7018 -10181 -7006 -10147
rect -6638 -10181 -6626 -10147
rect -7018 -10219 -6626 -10181
rect -7018 -10253 -7006 -10219
rect -6638 -10253 -6626 -10219
rect -7018 -10259 -6626 -10253
rect -6570 -10300 -6486 -10100
rect -6430 -10147 -6038 -10141
rect -6430 -10181 -6418 -10147
rect -6050 -10181 -6038 -10147
rect -6430 -10219 -6038 -10181
rect -6430 -10253 -6418 -10219
rect -6050 -10253 -6038 -10219
rect -6430 -10259 -6038 -10253
rect -5982 -10300 -5898 -10100
rect -5842 -10147 -5450 -10141
rect -5842 -10181 -5830 -10147
rect -5462 -10181 -5450 -10147
rect -5842 -10219 -5450 -10181
rect -5842 -10253 -5830 -10219
rect -5462 -10253 -5450 -10219
rect -5842 -10259 -5450 -10253
rect -5394 -10300 -5310 -10100
rect -5254 -10147 -4862 -10141
rect -5254 -10181 -5242 -10147
rect -4874 -10181 -4862 -10147
rect -5254 -10219 -4862 -10181
rect -5254 -10253 -5242 -10219
rect -4874 -10253 -4862 -10219
rect -5254 -10259 -4862 -10253
rect -4806 -10300 -4722 -10100
rect -4666 -10147 -4274 -10141
rect -4666 -10181 -4654 -10147
rect -4286 -10181 -4274 -10147
rect -4666 -10219 -4274 -10181
rect -4666 -10253 -4654 -10219
rect -4286 -10253 -4274 -10219
rect -4666 -10259 -4274 -10253
rect -4224 -10300 -4166 -10100
rect -4078 -10147 -3686 -10141
rect -4078 -10181 -4066 -10147
rect -3698 -10181 -3686 -10147
rect -4078 -10219 -3686 -10181
rect -4078 -10253 -4066 -10219
rect -3698 -10253 -3686 -10219
rect -4078 -10259 -3686 -10253
rect -3630 -10300 -3546 -10100
rect -3490 -10147 -3098 -10141
rect -3490 -10181 -3478 -10147
rect -3110 -10181 -3098 -10147
rect -3490 -10219 -3098 -10181
rect -3490 -10253 -3478 -10219
rect -3110 -10253 -3098 -10219
rect -3490 -10259 -3098 -10253
rect -3042 -10300 -2958 -10100
rect -2902 -10147 -2510 -10141
rect -2902 -10181 -2890 -10147
rect -2522 -10181 -2510 -10147
rect -2902 -10219 -2510 -10181
rect -2902 -10253 -2890 -10219
rect -2522 -10253 -2510 -10219
rect -2902 -10259 -2510 -10253
rect -2454 -10300 -2370 -10100
rect -2314 -10147 -1922 -10141
rect -2314 -10181 -2302 -10147
rect -1934 -10181 -1922 -10147
rect -2314 -10219 -1922 -10181
rect -2314 -10253 -2302 -10219
rect -1934 -10253 -1922 -10219
rect -2314 -10259 -1922 -10253
rect -1726 -10147 -1334 -10141
rect -1726 -10181 -1714 -10147
rect -1346 -10181 -1334 -10147
rect -1726 -10219 -1334 -10181
rect -1726 -10253 -1714 -10219
rect -1346 -10253 -1334 -10219
rect -1726 -10259 -1334 -10253
rect -1278 -10300 -1194 -10100
rect -1138 -10147 -746 -10141
rect -1138 -10181 -1126 -10147
rect -758 -10181 -746 -10147
rect -1138 -10219 -746 -10181
rect -1138 -10253 -1126 -10219
rect -758 -10253 -746 -10219
rect -1138 -10259 -746 -10253
rect -690 -10300 -606 -10100
rect -550 -10147 -158 -10141
rect -550 -10181 -538 -10147
rect -170 -10181 -158 -10147
rect -550 -10219 -158 -10181
rect -550 -10253 -538 -10219
rect -170 -10253 -158 -10219
rect -550 -10259 -158 -10253
rect -102 -10300 -18 -10100
rect 38 -10147 430 -10141
rect 38 -10181 50 -10147
rect 418 -10181 430 -10147
rect 38 -10219 430 -10181
rect 38 -10253 50 -10219
rect 418 -10253 430 -10219
rect 38 -10259 430 -10253
rect 520 -10300 576 -10100
rect 626 -10147 1018 -10141
rect 626 -10181 638 -10147
rect 1006 -10181 1018 -10147
rect 626 -10219 1018 -10181
rect 626 -10253 638 -10219
rect 1006 -10253 1018 -10219
rect 626 -10259 1018 -10253
rect 1074 -10300 1158 -10100
rect 1214 -10147 1606 -10141
rect 1214 -10181 1226 -10147
rect 1594 -10181 1606 -10147
rect 1214 -10219 1606 -10181
rect 1214 -10253 1226 -10219
rect 1594 -10253 1606 -10219
rect 1214 -10259 1606 -10253
rect 1662 -10300 1746 -10100
rect 1802 -10147 2194 -10141
rect 1802 -10181 1814 -10147
rect 2182 -10181 2194 -10147
rect 1802 -10219 2194 -10181
rect 1802 -10253 1814 -10219
rect 2182 -10253 2194 -10219
rect 1802 -10259 2194 -10253
rect 2250 -10300 2334 -10100
rect 2390 -10147 2782 -10141
rect 2390 -10181 2402 -10147
rect 2770 -10181 2782 -10147
rect 2390 -10219 2782 -10181
rect 2390 -10253 2402 -10219
rect 2770 -10253 2782 -10219
rect 2390 -10259 2782 -10253
rect 2838 -10300 2922 -10100
rect 2978 -10147 3370 -10141
rect 2978 -10181 2990 -10147
rect 3358 -10181 3370 -10147
rect 2978 -10219 3370 -10181
rect 2978 -10253 2990 -10219
rect 3358 -10253 3370 -10219
rect 2978 -10259 3370 -10253
rect 3426 -10300 3510 -10100
rect 3566 -10147 3958 -10141
rect 3566 -10181 3578 -10147
rect 3946 -10181 3958 -10147
rect 3566 -10219 3958 -10181
rect 3566 -10253 3578 -10219
rect 3946 -10253 3958 -10219
rect 3566 -10259 3958 -10253
rect 4014 -10300 4098 -10100
rect 4154 -10147 4546 -10141
rect 4154 -10181 4166 -10147
rect 4534 -10181 4546 -10147
rect 4154 -10219 4546 -10181
rect 4154 -10253 4166 -10219
rect 4534 -10253 4546 -10219
rect 4154 -10259 4546 -10253
rect 4602 -10300 4686 -10100
rect 4742 -10147 5134 -10141
rect 4742 -10181 4754 -10147
rect 5122 -10181 5134 -10147
rect 4742 -10219 5134 -10181
rect 4742 -10253 4754 -10219
rect 5122 -10253 5134 -10219
rect 4742 -10259 5134 -10253
rect 5190 -10300 5274 -10100
rect 5330 -10147 5722 -10141
rect 5330 -10181 5342 -10147
rect 5710 -10181 5722 -10147
rect 5330 -10219 5722 -10181
rect 5330 -10253 5342 -10219
rect 5710 -10253 5722 -10219
rect 5330 -10259 5722 -10253
rect 5778 -10300 5862 -10100
rect 5918 -10147 6310 -10141
rect 5918 -10181 5930 -10147
rect 6298 -10181 6310 -10147
rect 5918 -10219 6310 -10181
rect 5918 -10253 5930 -10219
rect 6298 -10253 6310 -10219
rect 5918 -10259 6310 -10253
rect 6366 -10300 6450 -10100
rect 6506 -10147 6898 -10141
rect 6506 -10181 6518 -10147
rect 6886 -10181 6898 -10147
rect 6506 -10219 6898 -10181
rect 6506 -10253 6518 -10219
rect 6886 -10253 6898 -10219
rect 6506 -10259 6898 -10253
rect 6954 -10300 7038 -10100
rect 7094 -10147 7486 -10141
rect 7094 -10181 7106 -10147
rect 7474 -10181 7486 -10147
rect 7094 -10219 7486 -10181
rect 7094 -10253 7106 -10219
rect 7474 -10253 7486 -10219
rect 7094 -10259 7486 -10253
rect 7542 -10300 7626 -10100
rect 7682 -10147 8074 -10141
rect 7682 -10181 7694 -10147
rect 8062 -10181 8074 -10147
rect 7682 -10219 8074 -10181
rect 7682 -10253 7694 -10219
rect 8062 -10253 8074 -10219
rect 7682 -10259 8074 -10253
rect 8130 -10300 8214 -10100
rect 8270 -10147 8662 -10141
rect 8270 -10181 8282 -10147
rect 8650 -10181 8662 -10147
rect 8270 -10219 8662 -10181
rect 8270 -10253 8282 -10219
rect 8650 -10253 8662 -10219
rect 8270 -10259 8662 -10253
rect 8718 -10300 8802 -10100
rect 8858 -10147 9250 -10141
rect 8858 -10181 8870 -10147
rect 9238 -10181 9250 -10147
rect 8858 -10219 9250 -10181
rect 8858 -10253 8870 -10219
rect 9238 -10253 9250 -10219
rect 8858 -10259 9250 -10253
rect 9306 -10300 9390 -10100
rect 9446 -10147 9838 -10141
rect 9446 -10181 9458 -10147
rect 9826 -10181 9838 -10147
rect 9446 -10219 9838 -10181
rect 9446 -10253 9458 -10219
rect 9826 -10253 9838 -10219
rect 9446 -10259 9838 -10253
rect 9894 -10300 9978 -10100
rect 10034 -10147 10426 -10141
rect 10034 -10181 10046 -10147
rect 10414 -10181 10426 -10147
rect 10034 -10219 10426 -10181
rect 10034 -10253 10046 -10219
rect 10414 -10253 10426 -10219
rect 10034 -10259 10426 -10253
rect 10482 -10300 10566 -10100
rect 10622 -10147 11014 -10141
rect 10622 -10181 10634 -10147
rect 11002 -10181 11014 -10147
rect 10622 -10219 11014 -10181
rect 10622 -10253 10634 -10219
rect 11002 -10253 11014 -10219
rect 10622 -10259 11014 -10253
rect 11070 -10300 11154 -10100
rect 11210 -10147 11602 -10141
rect 11210 -10181 11222 -10147
rect 11590 -10181 11602 -10147
rect 11210 -10219 11602 -10181
rect 11210 -10253 11222 -10219
rect 11590 -10253 11602 -10219
rect 11210 -10259 11602 -10253
rect 11658 -10300 11742 -10100
rect 11798 -10147 12190 -10141
rect 11798 -10181 11810 -10147
rect 12178 -10181 12190 -10147
rect 11798 -10219 12190 -10181
rect 11798 -10253 11810 -10219
rect 12178 -10253 12190 -10219
rect 11798 -10259 12190 -10253
rect 12246 -10300 12330 -10100
rect -15978 -10312 -15848 -10300
rect -15978 -11088 -15888 -10312
rect -15854 -11088 -15848 -10312
rect -15978 -11100 -15848 -11088
rect -15436 -10312 -15260 -10300
rect -15436 -11088 -15430 -10312
rect -15396 -11088 -15300 -10312
rect -15266 -11088 -15260 -10312
rect -15436 -11100 -15260 -11088
rect -14848 -10312 -14672 -10300
rect -14848 -11088 -14842 -10312
rect -14808 -11088 -14712 -10312
rect -14678 -11088 -14672 -10312
rect -14848 -11100 -14672 -11088
rect -14260 -10312 -14084 -10300
rect -14260 -11088 -14254 -10312
rect -14220 -11088 -14124 -10312
rect -14090 -11088 -14084 -10312
rect -14260 -11100 -14084 -11088
rect -13672 -10312 -13496 -10300
rect -13672 -11088 -13666 -10312
rect -13632 -11088 -13536 -10312
rect -13502 -11088 -13496 -10312
rect -13672 -11100 -13496 -11088
rect -13084 -10312 -12908 -10300
rect -13084 -11088 -13078 -10312
rect -13044 -11088 -12948 -10312
rect -12914 -11088 -12908 -10312
rect -13084 -11100 -12908 -11088
rect -12496 -10312 -12320 -10300
rect -12496 -11088 -12490 -10312
rect -12456 -11088 -12360 -10312
rect -12326 -11088 -12320 -10312
rect -12496 -11100 -12320 -11088
rect -11908 -10312 -11732 -10300
rect -11908 -11088 -11902 -10312
rect -11868 -11088 -11772 -10312
rect -11738 -11088 -11732 -10312
rect -11908 -11100 -11732 -11088
rect -11320 -10312 -11144 -10300
rect -11320 -11088 -11314 -10312
rect -11280 -11088 -11184 -10312
rect -11150 -11088 -11144 -10312
rect -11320 -11100 -11144 -11088
rect -10732 -10312 -10556 -10300
rect -10732 -11088 -10726 -10312
rect -10692 -11088 -10596 -10312
rect -10562 -11088 -10556 -10312
rect -10732 -11100 -10556 -11088
rect -10144 -10312 -9968 -10300
rect -10144 -11088 -10138 -10312
rect -10104 -11088 -10008 -10312
rect -9974 -11088 -9968 -10312
rect -10144 -11100 -9968 -11088
rect -9556 -10312 -9380 -10300
rect -9556 -11088 -9550 -10312
rect -9516 -11088 -9420 -10312
rect -9386 -11088 -9380 -10312
rect -9556 -11100 -9380 -11088
rect -8968 -10312 -8792 -10300
rect -8968 -11088 -8962 -10312
rect -8928 -11088 -8832 -10312
rect -8798 -11088 -8792 -10312
rect -8968 -11100 -8792 -11088
rect -8380 -10312 -8204 -10300
rect -8380 -11088 -8374 -10312
rect -8340 -11088 -8244 -10312
rect -8210 -11088 -8204 -10312
rect -8380 -11100 -8204 -11088
rect -7792 -10312 -7616 -10300
rect -7792 -11088 -7786 -10312
rect -7752 -11088 -7656 -10312
rect -7622 -11088 -7616 -10312
rect -7792 -11100 -7616 -11088
rect -7204 -10312 -7028 -10300
rect -7204 -11088 -7198 -10312
rect -7164 -11088 -7068 -10312
rect -7034 -11088 -7028 -10312
rect -7204 -11100 -7028 -11088
rect -6616 -10312 -6440 -10300
rect -6616 -11088 -6610 -10312
rect -6576 -11088 -6480 -10312
rect -6446 -11088 -6440 -10312
rect -6616 -11100 -6440 -11088
rect -6028 -10312 -5852 -10300
rect -6028 -11088 -6022 -10312
rect -5988 -11088 -5892 -10312
rect -5858 -11088 -5852 -10312
rect -6028 -11100 -5852 -11088
rect -5440 -10312 -5264 -10300
rect -5440 -11088 -5434 -10312
rect -5400 -11088 -5304 -10312
rect -5270 -11088 -5264 -10312
rect -5440 -11100 -5264 -11088
rect -4852 -10312 -4676 -10300
rect -4852 -11088 -4846 -10312
rect -4812 -11088 -4716 -10312
rect -4682 -11088 -4676 -10312
rect -4852 -11100 -4676 -11088
rect -4264 -10312 -4166 -10300
rect -4264 -11088 -4258 -10312
rect -4224 -11088 -4166 -10312
rect -4264 -11100 -4166 -11088
rect -4134 -10312 -4088 -10300
rect -4134 -11088 -4128 -10312
rect -4094 -11088 -4088 -10312
rect -4134 -11100 -4088 -11088
rect -3676 -10312 -3500 -10300
rect -3676 -11088 -3670 -10312
rect -3636 -11088 -3540 -10312
rect -3506 -11088 -3500 -10312
rect -3676 -11100 -3500 -11088
rect -3088 -10312 -2912 -10300
rect -3088 -11088 -3082 -10312
rect -3048 -11088 -2952 -10312
rect -2918 -11088 -2912 -10312
rect -3088 -11100 -2912 -11088
rect -2500 -10312 -2324 -10300
rect -2500 -11088 -2494 -10312
rect -2460 -11088 -2364 -10312
rect -2330 -11088 -2324 -10312
rect -2500 -11100 -2324 -11088
rect -1912 -10312 -1866 -10300
rect -1912 -11088 -1906 -10312
rect -1872 -11088 -1866 -10312
rect -1912 -11100 -1866 -11088
rect -1782 -10312 -1736 -10300
rect -1782 -11088 -1776 -10312
rect -1742 -11088 -1736 -10312
rect -1782 -11100 -1736 -11088
rect -1324 -10312 -1148 -10300
rect -1324 -11088 -1318 -10312
rect -1284 -11088 -1188 -10312
rect -1154 -11088 -1148 -10312
rect -1324 -11100 -1148 -11088
rect -736 -10312 -560 -10300
rect -736 -11088 -730 -10312
rect -696 -11088 -600 -10312
rect -566 -11088 -560 -10312
rect -736 -11100 -560 -11088
rect -148 -10312 28 -10300
rect -148 -11088 -142 -10312
rect -108 -11088 -12 -10312
rect 22 -11088 28 -10312
rect -148 -11100 28 -11088
rect 440 -10312 486 -10300
rect 440 -11088 446 -10312
rect 480 -11088 486 -10312
rect 440 -11100 486 -11088
rect 520 -10312 616 -10300
rect 520 -11088 576 -10312
rect 610 -11088 616 -10312
rect 520 -11100 616 -11088
rect 1028 -10312 1204 -10300
rect 1028 -11088 1034 -10312
rect 1068 -11088 1164 -10312
rect 1198 -11088 1204 -10312
rect 1028 -11100 1204 -11088
rect 1616 -10312 1792 -10300
rect 1616 -11088 1622 -10312
rect 1656 -11088 1752 -10312
rect 1786 -11088 1792 -10312
rect 1616 -11100 1792 -11088
rect 2204 -10312 2380 -10300
rect 2204 -11088 2210 -10312
rect 2244 -11088 2340 -10312
rect 2374 -11088 2380 -10312
rect 2204 -11100 2380 -11088
rect 2792 -10312 2968 -10300
rect 2792 -11088 2798 -10312
rect 2832 -11088 2928 -10312
rect 2962 -11088 2968 -10312
rect 2792 -11100 2968 -11088
rect 3380 -10312 3556 -10300
rect 3380 -11088 3386 -10312
rect 3420 -11088 3516 -10312
rect 3550 -11088 3556 -10312
rect 3380 -11100 3556 -11088
rect 3968 -10312 4144 -10300
rect 3968 -11088 3974 -10312
rect 4008 -11088 4104 -10312
rect 4138 -11088 4144 -10312
rect 3968 -11100 4144 -11088
rect 4556 -10312 4732 -10300
rect 4556 -11088 4562 -10312
rect 4596 -11088 4692 -10312
rect 4726 -11088 4732 -10312
rect 4556 -11100 4732 -11088
rect 5144 -10312 5320 -10300
rect 5144 -11088 5150 -10312
rect 5184 -11088 5280 -10312
rect 5314 -11088 5320 -10312
rect 5144 -11100 5320 -11088
rect 5732 -10312 5908 -10300
rect 5732 -11088 5738 -10312
rect 5772 -11088 5868 -10312
rect 5902 -11088 5908 -10312
rect 5732 -11100 5908 -11088
rect 6320 -10312 6496 -10300
rect 6320 -11088 6326 -10312
rect 6360 -11088 6456 -10312
rect 6490 -11088 6496 -10312
rect 6320 -11100 6496 -11088
rect 6908 -10312 7084 -10300
rect 6908 -11088 6914 -10312
rect 6948 -11088 7044 -10312
rect 7078 -11088 7084 -10312
rect 6908 -11100 7084 -11088
rect 7496 -10312 7672 -10300
rect 7496 -11088 7502 -10312
rect 7536 -11088 7632 -10312
rect 7666 -11088 7672 -10312
rect 7496 -11100 7672 -11088
rect 8084 -10312 8260 -10300
rect 8084 -11088 8090 -10312
rect 8124 -11088 8220 -10312
rect 8254 -11088 8260 -10312
rect 8084 -11100 8260 -11088
rect 8672 -10312 8848 -10300
rect 8672 -11088 8678 -10312
rect 8712 -11088 8808 -10312
rect 8842 -11088 8848 -10312
rect 8672 -11100 8848 -11088
rect 9260 -10312 9436 -10300
rect 9260 -11088 9266 -10312
rect 9300 -11088 9396 -10312
rect 9430 -11088 9436 -10312
rect 9260 -11100 9436 -11088
rect 9848 -10312 10024 -10300
rect 9848 -11088 9854 -10312
rect 9888 -11088 9984 -10312
rect 10018 -11088 10024 -10312
rect 9848 -11100 10024 -11088
rect 10436 -10312 10612 -10300
rect 10436 -11088 10442 -10312
rect 10476 -11088 10572 -10312
rect 10606 -11088 10612 -10312
rect 10436 -11100 10612 -11088
rect 11024 -10312 11200 -10300
rect 11024 -11088 11030 -10312
rect 11064 -11088 11160 -10312
rect 11194 -11088 11200 -10312
rect 11024 -11100 11200 -11088
rect 11612 -10312 11788 -10300
rect 11612 -11088 11618 -10312
rect 11652 -11088 11748 -10312
rect 11782 -11088 11788 -10312
rect 11612 -11100 11788 -11088
rect 12200 -10312 12330 -10300
rect 12200 -11088 12206 -10312
rect 12240 -11088 12330 -10312
rect 12200 -11100 12330 -11088
rect -15838 -11147 -15446 -11141
rect -15838 -11181 -15826 -11147
rect -15458 -11181 -15446 -11147
rect -15838 -11187 -15446 -11181
rect -15384 -11444 -15312 -11100
rect -15250 -11147 -14858 -11141
rect -15250 -11181 -15238 -11147
rect -14870 -11181 -14858 -11147
rect -15250 -11187 -14858 -11181
rect -14662 -11147 -14270 -11141
rect -14662 -11181 -14650 -11147
rect -14282 -11181 -14270 -11147
rect -14662 -11187 -14270 -11181
rect -14208 -11444 -14136 -11100
rect -14074 -11147 -13682 -11141
rect -14074 -11181 -14062 -11147
rect -13694 -11181 -13682 -11147
rect -14074 -11187 -13682 -11181
rect -13486 -11147 -13094 -11141
rect -13486 -11181 -13474 -11147
rect -13106 -11181 -13094 -11147
rect -13486 -11187 -13094 -11181
rect -13032 -11444 -12960 -11100
rect -12898 -11147 -12506 -11141
rect -12898 -11181 -12886 -11147
rect -12518 -11181 -12506 -11147
rect -12898 -11187 -12506 -11181
rect -12310 -11147 -11918 -11141
rect -12310 -11181 -12298 -11147
rect -11930 -11181 -11918 -11147
rect -12310 -11187 -11918 -11181
rect -11856 -11444 -11784 -11100
rect -11722 -11147 -11330 -11141
rect -11722 -11181 -11710 -11147
rect -11342 -11181 -11330 -11147
rect -11722 -11187 -11330 -11181
rect -11134 -11147 -10742 -11141
rect -11134 -11181 -11122 -11147
rect -10754 -11181 -10742 -11147
rect -11134 -11187 -10742 -11181
rect -10680 -11444 -10608 -11100
rect -10546 -11147 -10154 -11141
rect -10546 -11181 -10534 -11147
rect -10166 -11181 -10154 -11147
rect -10546 -11187 -10154 -11181
rect -9958 -11147 -9566 -11141
rect -9958 -11181 -9946 -11147
rect -9578 -11181 -9566 -11147
rect -9958 -11187 -9566 -11181
rect -9504 -11444 -9432 -11100
rect -9370 -11147 -8978 -11141
rect -9370 -11181 -9358 -11147
rect -8990 -11181 -8978 -11147
rect -9370 -11187 -8978 -11181
rect -8782 -11147 -8390 -11141
rect -8782 -11181 -8770 -11147
rect -8402 -11181 -8390 -11147
rect -8782 -11187 -8390 -11181
rect -8328 -11444 -8256 -11100
rect -8194 -11147 -7802 -11141
rect -8194 -11181 -8182 -11147
rect -7814 -11181 -7802 -11147
rect -8194 -11187 -7802 -11181
rect -7606 -11147 -7214 -11141
rect -7606 -11181 -7594 -11147
rect -7226 -11181 -7214 -11147
rect -7606 -11187 -7214 -11181
rect -7152 -11444 -7080 -11100
rect -7018 -11147 -6626 -11141
rect -7018 -11181 -7006 -11147
rect -6638 -11181 -6626 -11147
rect -7018 -11187 -6626 -11181
rect -6430 -11147 -6038 -11141
rect -6430 -11181 -6418 -11147
rect -6050 -11181 -6038 -11147
rect -6430 -11187 -6038 -11181
rect -5976 -11444 -5904 -11100
rect -5842 -11147 -5450 -11141
rect -5842 -11181 -5830 -11147
rect -5462 -11181 -5450 -11147
rect -5842 -11187 -5450 -11181
rect -5254 -11147 -4862 -11141
rect -5254 -11181 -5242 -11147
rect -4874 -11181 -4862 -11147
rect -5254 -11187 -4862 -11181
rect -4800 -11444 -4728 -11100
rect -4666 -11147 -4274 -11141
rect -4666 -11181 -4654 -11147
rect -4286 -11181 -4274 -11147
rect -4666 -11187 -4274 -11181
rect -4078 -11147 -3686 -11141
rect -4078 -11181 -4066 -11147
rect -3698 -11181 -3686 -11147
rect -4078 -11187 -3686 -11181
rect -3624 -11444 -3552 -11100
rect -3490 -11147 -3098 -11141
rect -3490 -11181 -3478 -11147
rect -3110 -11181 -3098 -11147
rect -3490 -11187 -3098 -11181
rect -15454 -11450 -15242 -11444
rect -15454 -11560 -15442 -11450
rect -15254 -11560 -15242 -11450
rect -15454 -11566 -15242 -11560
rect -14278 -11450 -14066 -11444
rect -14278 -11560 -14266 -11450
rect -14078 -11560 -14066 -11450
rect -14278 -11566 -14066 -11560
rect -13102 -11450 -12890 -11444
rect -13102 -11560 -13090 -11450
rect -12902 -11560 -12890 -11450
rect -13102 -11566 -12890 -11560
rect -11926 -11450 -11714 -11444
rect -11926 -11560 -11914 -11450
rect -11726 -11560 -11714 -11450
rect -11926 -11566 -11714 -11560
rect -10750 -11450 -10538 -11444
rect -10750 -11560 -10738 -11450
rect -10550 -11560 -10538 -11450
rect -10750 -11566 -10538 -11560
rect -9574 -11450 -9362 -11444
rect -9574 -11560 -9562 -11450
rect -9374 -11560 -9362 -11450
rect -9574 -11566 -9362 -11560
rect -8398 -11450 -8186 -11444
rect -8398 -11560 -8386 -11450
rect -8198 -11560 -8186 -11450
rect -8398 -11566 -8186 -11560
rect -7222 -11450 -7010 -11444
rect -7222 -11560 -7210 -11450
rect -7022 -11560 -7010 -11450
rect -7222 -11566 -7010 -11560
rect -6046 -11450 -5834 -11444
rect -6046 -11560 -6034 -11450
rect -5846 -11560 -5834 -11450
rect -6046 -11566 -5834 -11560
rect -4870 -11450 -4658 -11444
rect -4870 -11560 -4858 -11450
rect -4670 -11560 -4658 -11450
rect -4870 -11566 -4658 -11560
rect -3694 -11450 -3482 -11444
rect -3694 -11560 -3682 -11450
rect -3494 -11560 -3482 -11450
rect -3694 -11566 -3482 -11560
rect -3036 -11952 -2964 -11100
rect -2902 -11147 -2510 -11141
rect -2902 -11181 -2890 -11147
rect -2522 -11181 -2510 -11147
rect -2902 -11187 -2510 -11181
rect -2448 -11444 -2376 -11100
rect -2314 -11147 -1922 -11141
rect -2314 -11181 -2302 -11147
rect -1934 -11181 -1922 -11147
rect -2314 -11187 -1922 -11181
rect -1726 -11147 -1334 -11141
rect -1726 -11181 -1714 -11147
rect -1346 -11181 -1334 -11147
rect -1726 -11187 -1334 -11181
rect -1272 -11444 -1200 -11100
rect -1138 -11147 -746 -11141
rect -1138 -11181 -1126 -11147
rect -758 -11181 -746 -11147
rect -1138 -11187 -746 -11181
rect -2518 -11450 -2306 -11444
rect -2518 -11560 -2506 -11450
rect -2318 -11560 -2306 -11450
rect -2518 -11566 -2306 -11560
rect -1342 -11450 -1130 -11444
rect -1342 -11560 -1330 -11450
rect -1142 -11560 -1130 -11450
rect -1342 -11566 -1130 -11560
rect -684 -11952 -612 -11100
rect -550 -11147 -158 -11141
rect -550 -11181 -538 -11147
rect -170 -11181 -158 -11147
rect -550 -11187 -158 -11181
rect -96 -11444 -24 -11100
rect 38 -11147 430 -11141
rect 38 -11181 50 -11147
rect 418 -11181 430 -11147
rect 38 -11187 430 -11181
rect 626 -11147 1018 -11141
rect 626 -11181 638 -11147
rect 1006 -11181 1018 -11147
rect 626 -11187 1018 -11181
rect 1080 -11444 1152 -11100
rect 1214 -11147 1606 -11141
rect 1214 -11181 1226 -11147
rect 1594 -11181 1606 -11147
rect 1214 -11187 1606 -11181
rect 1802 -11147 2194 -11141
rect 1802 -11181 1814 -11147
rect 2182 -11181 2194 -11147
rect 1802 -11187 2194 -11181
rect 2256 -11444 2328 -11100
rect 2390 -11147 2782 -11141
rect 2390 -11181 2402 -11147
rect 2770 -11181 2782 -11147
rect 2390 -11187 2782 -11181
rect 2978 -11147 3370 -11141
rect 2978 -11181 2990 -11147
rect 3358 -11181 3370 -11147
rect 2978 -11187 3370 -11181
rect 3432 -11434 3504 -11100
rect 3566 -11147 3958 -11141
rect 3566 -11181 3578 -11147
rect 3946 -11181 3958 -11147
rect 3566 -11187 3958 -11181
rect 4154 -11147 4546 -11141
rect 4154 -11181 4166 -11147
rect 4534 -11181 4546 -11147
rect 4154 -11187 4546 -11181
rect 3362 -11440 3574 -11434
rect -166 -11450 46 -11444
rect -166 -11560 -154 -11450
rect 34 -11560 46 -11450
rect -166 -11566 46 -11560
rect 1010 -11450 1222 -11444
rect 1010 -11560 1022 -11450
rect 1210 -11560 1222 -11450
rect 1010 -11566 1222 -11560
rect 2186 -11450 2398 -11444
rect 2186 -11560 2198 -11450
rect 2386 -11560 2398 -11450
rect 3362 -11550 3374 -11440
rect 3562 -11550 3574 -11440
rect 4608 -11444 4680 -11100
rect 4742 -11147 5134 -11141
rect 4742 -11181 4754 -11147
rect 5122 -11181 5134 -11147
rect 4742 -11187 5134 -11181
rect 5330 -11147 5722 -11141
rect 5330 -11181 5342 -11147
rect 5710 -11181 5722 -11147
rect 5330 -11187 5722 -11181
rect 5784 -11444 5856 -11100
rect 5918 -11147 6310 -11141
rect 5918 -11181 5930 -11147
rect 6298 -11181 6310 -11147
rect 5918 -11187 6310 -11181
rect 6506 -11147 6898 -11141
rect 6506 -11181 6518 -11147
rect 6886 -11181 6898 -11147
rect 6506 -11187 6898 -11181
rect 6960 -11444 7032 -11100
rect 7094 -11147 7486 -11141
rect 7094 -11181 7106 -11147
rect 7474 -11181 7486 -11147
rect 7094 -11187 7486 -11181
rect 7682 -11147 8074 -11141
rect 7682 -11181 7694 -11147
rect 8062 -11181 8074 -11147
rect 7682 -11187 8074 -11181
rect 8136 -11434 8208 -11100
rect 8270 -11147 8662 -11141
rect 8270 -11181 8282 -11147
rect 8650 -11181 8662 -11147
rect 8270 -11187 8662 -11181
rect 8858 -11147 9250 -11141
rect 8858 -11181 8870 -11147
rect 9238 -11181 9250 -11147
rect 8858 -11187 9250 -11181
rect 8052 -11440 8288 -11434
rect 3362 -11556 3574 -11550
rect 4538 -11450 4750 -11444
rect 2186 -11566 2398 -11560
rect 4538 -11560 4550 -11450
rect 4738 -11560 4750 -11450
rect 4538 -11566 4750 -11560
rect 5714 -11450 5926 -11444
rect 5714 -11560 5726 -11450
rect 5914 -11560 5926 -11450
rect 5714 -11566 5926 -11560
rect 6890 -11450 7102 -11444
rect 6890 -11560 6902 -11450
rect 7090 -11560 7102 -11450
rect 6890 -11566 7102 -11560
rect 8052 -11562 8064 -11440
rect 8276 -11562 8288 -11440
rect 9312 -11444 9384 -11100
rect 9446 -11147 9838 -11141
rect 9446 -11181 9458 -11147
rect 9826 -11181 9838 -11147
rect 9446 -11187 9838 -11181
rect 10034 -11147 10426 -11141
rect 10034 -11181 10046 -11147
rect 10414 -11181 10426 -11147
rect 10034 -11187 10426 -11181
rect 10488 -11444 10560 -11100
rect 10622 -11147 11014 -11141
rect 10622 -11181 10634 -11147
rect 11002 -11181 11014 -11147
rect 10622 -11187 11014 -11181
rect 11210 -11147 11602 -11141
rect 11210 -11181 11222 -11147
rect 11590 -11181 11602 -11147
rect 11210 -11187 11602 -11181
rect 11664 -11444 11736 -11100
rect 11798 -11147 12190 -11141
rect 11798 -11181 11810 -11147
rect 12178 -11181 12190 -11147
rect 11798 -11187 12190 -11181
rect 8052 -11568 8288 -11562
rect 9242 -11450 9454 -11444
rect 9242 -11560 9254 -11450
rect 9442 -11560 9454 -11450
rect 9242 -11566 9454 -11560
rect 10418 -11450 10630 -11444
rect 10418 -11560 10430 -11450
rect 10618 -11560 10630 -11450
rect 10418 -11566 10630 -11560
rect 11594 -11450 11806 -11444
rect 11594 -11560 11606 -11450
rect 11794 -11560 11806 -11450
rect 11594 -11566 11806 -11560
rect -3036 -12032 -612 -11952
rect -2928 -12746 -2848 -12032
rect -2792 -12576 -2718 -12570
rect -2792 -12708 -2782 -12576
rect -2728 -12708 -2718 -12576
rect -2792 -12714 -2718 -12708
rect -2526 -12576 -2452 -12570
rect -2526 -12708 -2516 -12576
rect -2462 -12708 -2452 -12576
rect -2526 -12714 -2452 -12708
rect -2396 -12746 -2316 -12032
rect -2260 -12576 -2186 -12570
rect -2260 -12708 -2250 -12576
rect -2196 -12708 -2186 -12576
rect -2260 -12714 -2186 -12708
rect -1994 -12576 -1920 -12570
rect -1994 -12708 -1984 -12576
rect -1930 -12708 -1920 -12576
rect -1994 -12714 -1920 -12708
rect -1864 -12746 -1784 -12032
rect -1728 -12576 -1654 -12570
rect -1728 -12708 -1718 -12576
rect -1664 -12708 -1654 -12576
rect -1728 -12714 -1654 -12708
rect -1462 -12576 -1388 -12570
rect -1462 -12708 -1452 -12576
rect -1398 -12708 -1388 -12576
rect -1462 -12714 -1388 -12708
rect -1332 -12746 -1252 -12032
rect -1196 -12576 -1122 -12570
rect -1196 -12708 -1186 -12576
rect -1132 -12708 -1122 -12576
rect -1196 -12714 -1122 -12708
rect -930 -12576 -856 -12570
rect -930 -12708 -920 -12576
rect -866 -12708 -856 -12576
rect -930 -12714 -856 -12708
rect -800 -12746 -720 -12032
rect -2928 -12758 -2796 -12746
rect -2928 -13534 -2836 -12758
rect -2802 -13534 -2796 -12758
rect -2928 -13546 -2796 -13534
rect -2714 -12758 -2530 -12746
rect -2714 -13534 -2708 -12758
rect -2674 -13534 -2570 -12758
rect -2536 -13534 -2530 -12758
rect -2714 -13546 -2530 -13534
rect -2448 -12758 -2264 -12746
rect -2448 -13534 -2442 -12758
rect -2408 -13534 -2304 -12758
rect -2270 -13534 -2264 -12758
rect -2448 -13546 -2264 -13534
rect -2182 -12758 -1998 -12746
rect -2182 -13534 -2176 -12758
rect -2142 -13534 -2038 -12758
rect -2004 -13534 -1998 -12758
rect -2182 -13546 -1998 -13534
rect -1916 -12758 -1732 -12746
rect -1916 -13534 -1910 -12758
rect -1876 -13534 -1772 -12758
rect -1738 -13534 -1732 -12758
rect -1916 -13546 -1732 -13534
rect -1650 -12758 -1466 -12746
rect -1650 -13534 -1644 -12758
rect -1610 -13534 -1506 -12758
rect -1472 -13534 -1466 -12758
rect -1650 -13546 -1466 -13534
rect -1384 -12758 -1200 -12746
rect -1384 -13534 -1378 -12758
rect -1344 -13534 -1240 -12758
rect -1206 -13534 -1200 -12758
rect -1384 -13546 -1200 -13534
rect -1118 -12758 -934 -12746
rect -1118 -13534 -1112 -12758
rect -1078 -13534 -974 -12758
rect -940 -13534 -934 -12758
rect -1118 -13546 -934 -13534
rect -852 -12758 -720 -12746
rect -852 -13534 -846 -12758
rect -812 -13534 -720 -12758
rect -852 -13546 -720 -13534
rect -2928 -13756 -2842 -13546
rect -2792 -13586 -2718 -13580
rect -2792 -13718 -2782 -13586
rect -2728 -13718 -2718 -13586
rect -2792 -13724 -2718 -13718
rect -2668 -13756 -2576 -13546
rect -2526 -13586 -2452 -13580
rect -2526 -13718 -2516 -13586
rect -2462 -13718 -2452 -13586
rect -2526 -13724 -2452 -13718
rect -2402 -13756 -2310 -13546
rect -2260 -13586 -2186 -13580
rect -2260 -13718 -2250 -13586
rect -2196 -13718 -2186 -13586
rect -2260 -13724 -2186 -13718
rect -2136 -13756 -2044 -13546
rect -1994 -13586 -1920 -13580
rect -1994 -13718 -1984 -13586
rect -1930 -13718 -1920 -13586
rect -1994 -13724 -1920 -13718
rect -1870 -13756 -1778 -13546
rect -1728 -13586 -1654 -13580
rect -1728 -13718 -1718 -13586
rect -1664 -13718 -1654 -13586
rect -1728 -13724 -1654 -13718
rect -1604 -13756 -1512 -13546
rect -1462 -13586 -1388 -13580
rect -1462 -13718 -1452 -13586
rect -1398 -13718 -1388 -13586
rect -1462 -13724 -1388 -13718
rect -1338 -13756 -1246 -13546
rect -1196 -13586 -1122 -13580
rect -1196 -13718 -1186 -13586
rect -1132 -13718 -1122 -13586
rect -1196 -13724 -1122 -13718
rect -1072 -13756 -980 -13546
rect -930 -13586 -856 -13580
rect -930 -13718 -920 -13586
rect -866 -13718 -856 -13586
rect -930 -13724 -856 -13718
rect -806 -13756 -720 -13546
rect -2928 -13768 -2796 -13756
rect -2928 -14544 -2836 -13768
rect -2802 -14544 -2796 -13768
rect -2928 -14556 -2796 -14544
rect -2714 -13768 -2530 -13756
rect -2714 -14544 -2708 -13768
rect -2674 -14544 -2570 -13768
rect -2536 -14544 -2530 -13768
rect -2714 -14556 -2530 -14544
rect -2448 -13768 -2264 -13756
rect -2448 -14544 -2442 -13768
rect -2408 -14544 -2304 -13768
rect -2270 -14544 -2264 -13768
rect -2448 -14556 -2264 -14544
rect -2182 -13768 -1998 -13756
rect -2182 -14544 -2176 -13768
rect -2142 -14544 -2038 -13768
rect -2004 -14544 -1998 -13768
rect -2182 -14556 -1998 -14544
rect -1916 -13768 -1732 -13756
rect -1916 -14544 -1910 -13768
rect -1876 -14544 -1772 -13768
rect -1738 -14544 -1732 -13768
rect -1916 -14556 -1732 -14544
rect -1650 -13768 -1466 -13756
rect -1650 -14544 -1644 -13768
rect -1610 -14544 -1506 -13768
rect -1472 -14544 -1466 -13768
rect -1650 -14556 -1466 -14544
rect -1384 -13768 -1200 -13756
rect -1384 -14544 -1378 -13768
rect -1344 -14544 -1240 -13768
rect -1206 -14544 -1200 -13768
rect -1384 -14556 -1200 -14544
rect -1118 -13768 -934 -13756
rect -1118 -14544 -1112 -13768
rect -1078 -14544 -974 -13768
rect -940 -14544 -934 -13768
rect -1118 -14556 -934 -14544
rect -852 -13768 -720 -13756
rect -852 -14544 -846 -13768
rect -812 -14544 -720 -13768
rect -852 -14556 -720 -14544
rect -2928 -14766 -2842 -14556
rect -2792 -14596 -2718 -14590
rect -2792 -14728 -2782 -14596
rect -2728 -14728 -2718 -14596
rect -2792 -14734 -2718 -14728
rect -2668 -14766 -2576 -14556
rect -2526 -14596 -2452 -14590
rect -2526 -14728 -2516 -14596
rect -2462 -14728 -2452 -14596
rect -2526 -14734 -2452 -14728
rect -2402 -14766 -2310 -14556
rect -2260 -14596 -2186 -14590
rect -2260 -14728 -2250 -14596
rect -2196 -14728 -2186 -14596
rect -2260 -14734 -2186 -14728
rect -2136 -14766 -2044 -14556
rect -1994 -14596 -1920 -14590
rect -1994 -14728 -1984 -14596
rect -1930 -14728 -1920 -14596
rect -1994 -14734 -1920 -14728
rect -1870 -14766 -1778 -14556
rect -1728 -14596 -1654 -14590
rect -1728 -14728 -1718 -14596
rect -1664 -14728 -1654 -14596
rect -1728 -14734 -1654 -14728
rect -1604 -14766 -1512 -14556
rect -1462 -14596 -1388 -14590
rect -1462 -14728 -1452 -14596
rect -1398 -14728 -1388 -14596
rect -1462 -14734 -1388 -14728
rect -1338 -14766 -1246 -14556
rect -1196 -14596 -1122 -14590
rect -1196 -14728 -1186 -14596
rect -1132 -14728 -1122 -14596
rect -1196 -14734 -1122 -14728
rect -1072 -14766 -980 -14556
rect -930 -14596 -856 -14590
rect -930 -14728 -920 -14596
rect -866 -14728 -856 -14596
rect -930 -14734 -856 -14728
rect -806 -14766 -720 -14556
rect 4356 -14724 4366 -14514
rect 4570 -14724 4580 -14514
rect -2928 -14778 -2796 -14766
rect -2928 -15554 -2836 -14778
rect -2802 -15554 -2796 -14778
rect -2928 -15566 -2796 -15554
rect -2714 -14778 -2530 -14766
rect -2714 -15554 -2708 -14778
rect -2674 -15554 -2570 -14778
rect -2536 -15554 -2530 -14778
rect -2714 -15566 -2530 -15554
rect -2448 -14778 -2264 -14766
rect -2448 -15554 -2442 -14778
rect -2408 -15554 -2304 -14778
rect -2270 -15554 -2264 -14778
rect -2448 -15566 -2264 -15554
rect -2182 -14778 -1998 -14766
rect -2182 -15554 -2176 -14778
rect -2142 -15554 -2038 -14778
rect -2004 -15554 -1998 -14778
rect -2182 -15566 -1998 -15554
rect -1916 -14778 -1732 -14766
rect -1916 -15554 -1910 -14778
rect -1876 -15554 -1772 -14778
rect -1738 -15554 -1732 -14778
rect -1916 -15566 -1732 -15554
rect -1650 -14778 -1466 -14766
rect -1650 -15554 -1644 -14778
rect -1610 -15554 -1506 -14778
rect -1472 -15554 -1466 -14778
rect -1650 -15566 -1466 -15554
rect -1384 -14778 -1200 -14766
rect -1384 -15554 -1378 -14778
rect -1344 -15554 -1240 -14778
rect -1206 -15554 -1200 -14778
rect -1384 -15566 -1200 -15554
rect -1118 -14778 -934 -14766
rect -1118 -15554 -1112 -14778
rect -1078 -15554 -974 -14778
rect -940 -15554 -934 -14778
rect -1118 -15566 -934 -15554
rect -852 -14778 -720 -14766
rect -852 -15554 -846 -14778
rect -812 -15554 -720 -14778
rect 4366 -14997 4438 -14724
rect 4366 -15088 4383 -14997
rect 4377 -15394 4383 -15088
rect 4421 -15088 4438 -14997
rect 4618 -14878 4792 -14858
rect 4421 -15394 4427 -15088
rect 4377 -15406 4427 -15394
rect 4618 -15338 4634 -14878
rect 4774 -15338 4792 -14878
rect -852 -15566 -720 -15554
rect 4377 -15528 4427 -15516
rect -2792 -15606 -2718 -15600
rect -2792 -15738 -2782 -15606
rect -2728 -15738 -2718 -15606
rect -2792 -15744 -2718 -15738
rect -2662 -16938 -2582 -15566
rect -2526 -15606 -2452 -15600
rect -2526 -15738 -2516 -15606
rect -2462 -15738 -2452 -15606
rect -2526 -15744 -2452 -15738
rect -2260 -15606 -2186 -15600
rect -2260 -15738 -2250 -15606
rect -2196 -15738 -2186 -15606
rect -2260 -15744 -2186 -15738
rect -2130 -16122 -2050 -15566
rect -1994 -15606 -1920 -15600
rect -1994 -15738 -1984 -15606
rect -1930 -15738 -1920 -15606
rect -1994 -15744 -1920 -15738
rect -1728 -15606 -1654 -15600
rect -1728 -15738 -1718 -15606
rect -1664 -15738 -1654 -15606
rect -1728 -15744 -1654 -15738
rect -1598 -16122 -1518 -15566
rect -1462 -15606 -1388 -15600
rect -1462 -15738 -1452 -15606
rect -1398 -15738 -1388 -15606
rect -1462 -15744 -1388 -15738
rect -1196 -15606 -1122 -15600
rect -1196 -15738 -1186 -15606
rect -1132 -15738 -1122 -15606
rect -1196 -15744 -1122 -15738
rect -2130 -16154 -1518 -16122
rect -2130 -16282 -2084 -16154
rect -1590 -16282 -1518 -16154
rect -2130 -16312 -1518 -16282
rect -2218 -16774 -1908 -16768
rect -2218 -16900 -2202 -16774
rect -2164 -16900 -1962 -16774
rect -1924 -16900 -1908 -16774
rect -2218 -16906 -2148 -16900
rect -1978 -16906 -1908 -16900
rect -1850 -16938 -1796 -16312
rect -1738 -16774 -1428 -16768
rect -1738 -16900 -1722 -16774
rect -1684 -16900 -1482 -16774
rect -1444 -16900 -1428 -16774
rect -1738 -16906 -1668 -16900
rect -1498 -16906 -1428 -16900
rect -1066 -16938 -986 -15566
rect -930 -15606 -856 -15600
rect -930 -15738 -920 -15606
rect -866 -15738 -856 -15606
rect -930 -15744 -856 -15738
rect 4377 -15914 4383 -15528
rect 4366 -15925 4383 -15914
rect 4421 -15914 4427 -15528
rect 4421 -15925 4438 -15914
rect 4366 -16136 4438 -15925
rect 4198 -16472 4208 -16136
rect 4520 -16472 4530 -16136
rect -2662 -16950 -2224 -16938
rect -2662 -17008 -2264 -16950
rect -2314 -17526 -2264 -17008
rect -2230 -17526 -2224 -16950
rect -2314 -17538 -2224 -17526
rect -2142 -16950 -1984 -16938
rect -2142 -17526 -2136 -16950
rect -2102 -17526 -2024 -16950
rect -1990 -17526 -1984 -16950
rect -2142 -17538 -1984 -17526
rect -1902 -16950 -1744 -16938
rect -1902 -17526 -1896 -16950
rect -1862 -17526 -1784 -16950
rect -1750 -17526 -1744 -16950
rect -1902 -17538 -1744 -17526
rect -1662 -16950 -1504 -16938
rect -1662 -17526 -1656 -16950
rect -1622 -17526 -1544 -16950
rect -1510 -17526 -1504 -16950
rect -1662 -17538 -1504 -17526
rect -1422 -16950 -986 -16938
rect -1422 -17526 -1416 -16950
rect -1382 -17008 -986 -16950
rect -1382 -17526 -1326 -17008
rect -1422 -17538 -1326 -17526
rect -2314 -17746 -2264 -17538
rect -2218 -17576 -2148 -17570
rect -2218 -17708 -2202 -17576
rect -2164 -17708 -2148 -17576
rect -2218 -17714 -2148 -17708
rect -2096 -17746 -2030 -17538
rect -1978 -17576 -1908 -17570
rect -1978 -17708 -1962 -17576
rect -1924 -17708 -1908 -17576
rect -1978 -17714 -1908 -17708
rect -1856 -17746 -1790 -17538
rect -1738 -17576 -1668 -17570
rect -1738 -17708 -1722 -17576
rect -1684 -17708 -1668 -17576
rect -1738 -17714 -1668 -17708
rect -1616 -17746 -1550 -17538
rect -1498 -17576 -1428 -17570
rect -1498 -17708 -1482 -17576
rect -1444 -17708 -1428 -17576
rect -1498 -17714 -1428 -17708
rect -1376 -17746 -1326 -17538
rect -2314 -17758 -2224 -17746
rect -2314 -18334 -2264 -17758
rect -2230 -18334 -2224 -17758
rect -2314 -18346 -2224 -18334
rect -2142 -17758 -1984 -17746
rect -2142 -18334 -2136 -17758
rect -2102 -18334 -2024 -17758
rect -1990 -18334 -1984 -17758
rect -2142 -18346 -1984 -18334
rect -1902 -17758 -1744 -17746
rect -1902 -18334 -1896 -17758
rect -1862 -18334 -1784 -17758
rect -1750 -18334 -1744 -17758
rect -1902 -18346 -1744 -18334
rect -1662 -17758 -1504 -17746
rect -1662 -18334 -1656 -17758
rect -1622 -18334 -1544 -17758
rect -1510 -18334 -1504 -17758
rect -1662 -18346 -1504 -18334
rect -1422 -17758 -1326 -17746
rect -1422 -18334 -1416 -17758
rect -1382 -18334 -1326 -17758
rect 4618 -18188 4792 -15338
rect -1422 -18346 -1326 -18334
rect -2218 -18384 -2148 -18378
rect -2218 -18516 -2202 -18384
rect -2164 -18516 -2148 -18384
rect -2218 -18522 -2148 -18516
rect -2090 -18762 -2036 -18346
rect -1978 -18384 -1908 -18378
rect -1978 -18516 -1962 -18384
rect -1924 -18516 -1908 -18384
rect -1978 -18522 -1908 -18516
rect -1738 -18384 -1668 -18378
rect -1738 -18516 -1722 -18384
rect -1684 -18516 -1668 -18384
rect -1738 -18522 -1668 -18516
rect -1610 -18762 -1556 -18346
rect -1498 -18384 -1428 -18378
rect -1498 -18516 -1482 -18384
rect -1444 -18516 -1428 -18384
rect -1498 -18522 -1428 -18516
rect -2524 -18768 -1148 -18762
rect -2524 -18880 -2512 -18768
rect -1160 -18880 -1148 -18768
rect 4330 -18854 4340 -18188
rect 5096 -18854 5106 -18188
rect -2524 -18886 -1148 -18880
<< via1 >>
rect -6438 -3784 -6328 -3712
rect -5958 -3784 -5848 -3712
rect -5478 -3784 -5368 -3712
rect -4998 -3784 -4888 -3712
rect -4518 -3784 -4408 -3712
rect -4038 -3784 -3928 -3712
rect -3558 -3784 -3448 -3712
rect -3078 -3784 -2968 -3712
rect -2598 -3784 -2488 -3712
rect -2118 -3784 -2008 -3712
rect -1638 -3784 -1528 -3712
rect -1158 -3784 -1048 -3712
rect -678 -3784 -568 -3712
rect -198 -3784 -88 -3712
rect 282 -3784 392 -3712
rect 762 -3784 872 -3712
rect 1242 -3784 1352 -3712
rect 1722 -3784 1832 -3712
rect 2202 -3784 2312 -3712
rect 2682 -3784 2792 -3712
rect -6538 -4188 -6522 -4056
rect -6522 -4188 -6484 -4056
rect -6484 -4188 -6468 -4056
rect -6298 -4188 -6282 -4056
rect -6282 -4188 -6244 -4056
rect -6244 -4188 -6228 -4056
rect -6058 -4188 -6042 -4056
rect -6042 -4188 -6004 -4056
rect -6004 -4188 -5988 -4056
rect -5818 -4188 -5802 -4056
rect -5802 -4188 -5764 -4056
rect -5764 -4188 -5748 -4056
rect -5578 -4188 -5562 -4056
rect -5562 -4188 -5524 -4056
rect -5524 -4188 -5508 -4056
rect -5338 -4188 -5322 -4056
rect -5322 -4188 -5284 -4056
rect -5284 -4188 -5268 -4056
rect -5098 -4188 -5082 -4056
rect -5082 -4188 -5044 -4056
rect -5044 -4188 -5028 -4056
rect -4858 -4188 -4842 -4056
rect -4842 -4188 -4804 -4056
rect -4804 -4188 -4788 -4056
rect -4618 -4188 -4602 -4056
rect -4602 -4188 -4564 -4056
rect -4564 -4188 -4548 -4056
rect -4378 -4188 -4362 -4056
rect -4362 -4188 -4324 -4056
rect -4324 -4188 -4308 -4056
rect -4138 -4188 -4122 -4056
rect -4122 -4188 -4084 -4056
rect -4084 -4188 -4068 -4056
rect -3898 -4188 -3882 -4056
rect -3882 -4188 -3844 -4056
rect -3844 -4188 -3828 -4056
rect -3658 -4188 -3642 -4056
rect -3642 -4188 -3604 -4056
rect -3604 -4188 -3588 -4056
rect -3418 -4188 -3402 -4056
rect -3402 -4188 -3364 -4056
rect -3364 -4188 -3348 -4056
rect -3178 -4188 -3162 -4056
rect -3162 -4188 -3124 -4056
rect -3124 -4188 -3108 -4056
rect -2938 -4188 -2922 -4056
rect -2922 -4188 -2884 -4056
rect -2884 -4188 -2868 -4056
rect -2698 -4188 -2682 -4056
rect -2682 -4188 -2644 -4056
rect -2644 -4188 -2628 -4056
rect -2458 -4188 -2442 -4056
rect -2442 -4188 -2404 -4056
rect -2404 -4188 -2388 -4056
rect -2218 -4188 -2202 -4056
rect -2202 -4188 -2164 -4056
rect -2164 -4188 -2148 -4056
rect -1978 -4188 -1962 -4056
rect -1962 -4188 -1924 -4056
rect -1924 -4188 -1908 -4056
rect -1738 -4188 -1722 -4056
rect -1722 -4188 -1684 -4056
rect -1684 -4188 -1668 -4056
rect -1498 -4188 -1482 -4056
rect -1482 -4188 -1444 -4056
rect -1444 -4188 -1428 -4056
rect -1258 -4188 -1242 -4056
rect -1242 -4188 -1204 -4056
rect -1204 -4188 -1188 -4056
rect -1018 -4188 -1002 -4056
rect -1002 -4188 -964 -4056
rect -964 -4188 -948 -4056
rect -778 -4188 -762 -4056
rect -762 -4188 -724 -4056
rect -724 -4188 -708 -4056
rect -538 -4188 -522 -4056
rect -522 -4188 -484 -4056
rect -484 -4188 -468 -4056
rect -298 -4188 -282 -4056
rect -282 -4188 -244 -4056
rect -244 -4188 -228 -4056
rect -58 -4188 -42 -4056
rect -42 -4188 -4 -4056
rect -4 -4188 12 -4056
rect 182 -4188 198 -4056
rect 198 -4188 236 -4056
rect 236 -4188 252 -4056
rect 422 -4188 438 -4056
rect 438 -4188 476 -4056
rect 476 -4188 492 -4056
rect 662 -4188 678 -4056
rect 678 -4188 716 -4056
rect 716 -4188 732 -4056
rect 902 -4188 918 -4056
rect 918 -4188 956 -4056
rect 956 -4188 972 -4056
rect 1142 -4188 1158 -4056
rect 1158 -4188 1196 -4056
rect 1196 -4188 1212 -4056
rect 1382 -4188 1398 -4056
rect 1398 -4188 1436 -4056
rect 1436 -4188 1452 -4056
rect 1622 -4188 1638 -4056
rect 1638 -4188 1676 -4056
rect 1676 -4188 1692 -4056
rect 1862 -4188 1878 -4056
rect 1878 -4188 1916 -4056
rect 1916 -4188 1932 -4056
rect 2102 -4188 2118 -4056
rect 2118 -4188 2156 -4056
rect 2156 -4188 2172 -4056
rect 2342 -4188 2358 -4056
rect 2358 -4188 2396 -4056
rect 2396 -4188 2412 -4056
rect 2582 -4188 2598 -4056
rect 2598 -4188 2636 -4056
rect 2636 -4188 2652 -4056
rect 2822 -4188 2838 -4056
rect 2838 -4188 2876 -4056
rect 2876 -4188 2892 -4056
rect -6538 -4996 -6522 -4864
rect -6522 -4996 -6484 -4864
rect -6484 -4996 -6468 -4864
rect -6298 -4996 -6282 -4864
rect -6282 -4996 -6244 -4864
rect -6244 -4996 -6228 -4864
rect -6058 -4996 -6042 -4864
rect -6042 -4996 -6004 -4864
rect -6004 -4996 -5988 -4864
rect -5818 -4996 -5802 -4864
rect -5802 -4996 -5764 -4864
rect -5764 -4996 -5748 -4864
rect -5578 -4996 -5562 -4864
rect -5562 -4996 -5524 -4864
rect -5524 -4996 -5508 -4864
rect -5338 -4996 -5322 -4864
rect -5322 -4996 -5284 -4864
rect -5284 -4996 -5268 -4864
rect -5098 -4996 -5082 -4864
rect -5082 -4996 -5044 -4864
rect -5044 -4996 -5028 -4864
rect -4858 -4996 -4842 -4864
rect -4842 -4996 -4804 -4864
rect -4804 -4996 -4788 -4864
rect -4618 -4996 -4602 -4864
rect -4602 -4996 -4564 -4864
rect -4564 -4996 -4548 -4864
rect -4378 -4996 -4362 -4864
rect -4362 -4996 -4324 -4864
rect -4324 -4996 -4308 -4864
rect -4138 -4996 -4122 -4864
rect -4122 -4996 -4084 -4864
rect -4084 -4996 -4068 -4864
rect -3898 -4996 -3882 -4864
rect -3882 -4996 -3844 -4864
rect -3844 -4996 -3828 -4864
rect -3658 -4996 -3642 -4864
rect -3642 -4996 -3604 -4864
rect -3604 -4996 -3588 -4864
rect -3418 -4996 -3402 -4864
rect -3402 -4996 -3364 -4864
rect -3364 -4996 -3348 -4864
rect -3178 -4996 -3162 -4864
rect -3162 -4996 -3124 -4864
rect -3124 -4996 -3108 -4864
rect -2938 -4996 -2922 -4864
rect -2922 -4996 -2884 -4864
rect -2884 -4996 -2868 -4864
rect -2698 -4996 -2682 -4864
rect -2682 -4996 -2644 -4864
rect -2644 -4996 -2628 -4864
rect -2458 -4996 -2442 -4864
rect -2442 -4996 -2404 -4864
rect -2404 -4996 -2388 -4864
rect -2218 -4996 -2202 -4864
rect -2202 -4996 -2164 -4864
rect -2164 -4996 -2148 -4864
rect -1978 -4996 -1962 -4864
rect -1962 -4996 -1924 -4864
rect -1924 -4996 -1908 -4864
rect -1738 -4996 -1722 -4864
rect -1722 -4996 -1684 -4864
rect -1684 -4996 -1668 -4864
rect -1498 -4996 -1482 -4864
rect -1482 -4996 -1444 -4864
rect -1444 -4996 -1428 -4864
rect -1258 -4996 -1242 -4864
rect -1242 -4996 -1204 -4864
rect -1204 -4996 -1188 -4864
rect -1018 -4996 -1002 -4864
rect -1002 -4996 -964 -4864
rect -964 -4996 -948 -4864
rect -778 -4996 -762 -4864
rect -762 -4996 -724 -4864
rect -724 -4996 -708 -4864
rect -538 -4996 -522 -4864
rect -522 -4996 -484 -4864
rect -484 -4996 -468 -4864
rect -298 -4996 -282 -4864
rect -282 -4996 -244 -4864
rect -244 -4996 -228 -4864
rect -58 -4996 -42 -4864
rect -42 -4996 -4 -4864
rect -4 -4996 12 -4864
rect 182 -4996 198 -4864
rect 198 -4996 236 -4864
rect 236 -4996 252 -4864
rect 422 -4996 438 -4864
rect 438 -4996 476 -4864
rect 476 -4996 492 -4864
rect 662 -4996 678 -4864
rect 678 -4996 716 -4864
rect 716 -4996 732 -4864
rect 902 -4996 918 -4864
rect 918 -4996 956 -4864
rect 956 -4996 972 -4864
rect 1142 -4996 1158 -4864
rect 1158 -4996 1196 -4864
rect 1196 -4996 1212 -4864
rect 1382 -4996 1398 -4864
rect 1398 -4996 1436 -4864
rect 1436 -4996 1452 -4864
rect 1622 -4996 1638 -4864
rect 1638 -4996 1676 -4864
rect 1676 -4996 1692 -4864
rect 1862 -4996 1878 -4864
rect 1878 -4996 1916 -4864
rect 1916 -4996 1932 -4864
rect 2102 -4996 2118 -4864
rect 2118 -4996 2156 -4864
rect 2156 -4996 2172 -4864
rect 2342 -4996 2358 -4864
rect 2358 -4996 2396 -4864
rect 2396 -4996 2412 -4864
rect 2582 -4996 2598 -4864
rect 2598 -4996 2636 -4864
rect 2636 -4996 2652 -4864
rect 2822 -4996 2838 -4864
rect 2838 -4996 2876 -4864
rect 2876 -4996 2892 -4864
rect -6538 -5804 -6522 -5672
rect -6522 -5804 -6484 -5672
rect -6484 -5804 -6468 -5672
rect -6298 -5804 -6282 -5672
rect -6282 -5804 -6244 -5672
rect -6244 -5804 -6228 -5672
rect -6058 -5804 -6042 -5672
rect -6042 -5804 -6004 -5672
rect -6004 -5804 -5988 -5672
rect -5818 -5804 -5802 -5672
rect -5802 -5804 -5764 -5672
rect -5764 -5804 -5748 -5672
rect -5578 -5804 -5562 -5672
rect -5562 -5804 -5524 -5672
rect -5524 -5804 -5508 -5672
rect -5338 -5804 -5322 -5672
rect -5322 -5804 -5284 -5672
rect -5284 -5804 -5268 -5672
rect -5098 -5804 -5082 -5672
rect -5082 -5804 -5044 -5672
rect -5044 -5804 -5028 -5672
rect -4858 -5804 -4842 -5672
rect -4842 -5804 -4804 -5672
rect -4804 -5804 -4788 -5672
rect -4618 -5804 -4602 -5672
rect -4602 -5804 -4564 -5672
rect -4564 -5804 -4548 -5672
rect -4378 -5804 -4362 -5672
rect -4362 -5804 -4324 -5672
rect -4324 -5804 -4308 -5672
rect -4138 -5804 -4122 -5672
rect -4122 -5804 -4084 -5672
rect -4084 -5804 -4068 -5672
rect -3898 -5804 -3882 -5672
rect -3882 -5804 -3844 -5672
rect -3844 -5804 -3828 -5672
rect -3658 -5804 -3642 -5672
rect -3642 -5804 -3604 -5672
rect -3604 -5804 -3588 -5672
rect -3418 -5804 -3402 -5672
rect -3402 -5804 -3364 -5672
rect -3364 -5804 -3348 -5672
rect -3178 -5804 -3162 -5672
rect -3162 -5804 -3124 -5672
rect -3124 -5804 -3108 -5672
rect -2938 -5804 -2922 -5672
rect -2922 -5804 -2884 -5672
rect -2884 -5804 -2868 -5672
rect -2698 -5804 -2682 -5672
rect -2682 -5804 -2644 -5672
rect -2644 -5804 -2628 -5672
rect -2458 -5804 -2442 -5672
rect -2442 -5804 -2404 -5672
rect -2404 -5804 -2388 -5672
rect -2218 -5804 -2202 -5672
rect -2202 -5804 -2164 -5672
rect -2164 -5804 -2148 -5672
rect -1978 -5804 -1962 -5672
rect -1962 -5804 -1924 -5672
rect -1924 -5804 -1908 -5672
rect -1738 -5804 -1722 -5672
rect -1722 -5804 -1684 -5672
rect -1684 -5804 -1668 -5672
rect -1498 -5804 -1482 -5672
rect -1482 -5804 -1444 -5672
rect -1444 -5804 -1428 -5672
rect -1258 -5804 -1242 -5672
rect -1242 -5804 -1204 -5672
rect -1204 -5804 -1188 -5672
rect -1018 -5804 -1002 -5672
rect -1002 -5804 -964 -5672
rect -964 -5804 -948 -5672
rect -778 -5804 -762 -5672
rect -762 -5804 -724 -5672
rect -724 -5804 -708 -5672
rect -538 -5804 -522 -5672
rect -522 -5804 -484 -5672
rect -484 -5804 -468 -5672
rect -298 -5804 -282 -5672
rect -282 -5804 -244 -5672
rect -244 -5804 -228 -5672
rect -58 -5804 -42 -5672
rect -42 -5804 -4 -5672
rect -4 -5804 12 -5672
rect 182 -5804 198 -5672
rect 198 -5804 236 -5672
rect 236 -5804 252 -5672
rect 422 -5804 438 -5672
rect 438 -5804 476 -5672
rect 476 -5804 492 -5672
rect 662 -5804 678 -5672
rect 678 -5804 716 -5672
rect 716 -5804 732 -5672
rect 902 -5804 918 -5672
rect 918 -5804 956 -5672
rect 956 -5804 972 -5672
rect 1142 -5804 1158 -5672
rect 1158 -5804 1196 -5672
rect 1196 -5804 1212 -5672
rect 1382 -5804 1398 -5672
rect 1398 -5804 1436 -5672
rect 1436 -5804 1452 -5672
rect 1622 -5804 1638 -5672
rect 1638 -5804 1676 -5672
rect 1676 -5804 1692 -5672
rect 1862 -5804 1878 -5672
rect 1878 -5804 1916 -5672
rect 1916 -5804 1932 -5672
rect 2102 -5804 2118 -5672
rect 2118 -5804 2156 -5672
rect 2156 -5804 2172 -5672
rect 2342 -5804 2358 -5672
rect 2358 -5804 2396 -5672
rect 2396 -5804 2412 -5672
rect 2582 -5804 2598 -5672
rect 2598 -5804 2636 -5672
rect 2636 -5804 2652 -5672
rect 2822 -5804 2838 -5672
rect 2838 -5804 2876 -5672
rect 2876 -5804 2892 -5672
rect 7404 -7196 8304 -6698
rect -15442 -11560 -15254 -11450
rect -14266 -11560 -14078 -11450
rect -13090 -11560 -12902 -11450
rect -11914 -11560 -11726 -11450
rect -10738 -11560 -10550 -11450
rect -9562 -11560 -9374 -11450
rect -8386 -11560 -8198 -11450
rect -7210 -11560 -7022 -11450
rect -6034 -11560 -5846 -11450
rect -4858 -11560 -4670 -11450
rect -3682 -11560 -3494 -11450
rect -2506 -11560 -2318 -11450
rect -1330 -11560 -1142 -11450
rect -154 -11560 34 -11450
rect 1022 -11560 1210 -11450
rect 2198 -11560 2386 -11450
rect 4550 -11560 4738 -11450
rect 5726 -11560 5914 -11450
rect 6902 -11560 7090 -11450
rect 9254 -11560 9442 -11450
rect 10430 -11560 10618 -11450
rect 11606 -11560 11794 -11450
rect -2782 -12708 -2774 -12576
rect -2774 -12708 -2736 -12576
rect -2736 -12708 -2728 -12576
rect -2516 -12708 -2508 -12576
rect -2508 -12708 -2470 -12576
rect -2470 -12708 -2462 -12576
rect -2250 -12708 -2242 -12576
rect -2242 -12708 -2204 -12576
rect -2204 -12708 -2196 -12576
rect -1984 -12708 -1976 -12576
rect -1976 -12708 -1938 -12576
rect -1938 -12708 -1930 -12576
rect -1718 -12708 -1710 -12576
rect -1710 -12708 -1672 -12576
rect -1672 -12708 -1664 -12576
rect -1452 -12708 -1444 -12576
rect -1444 -12708 -1406 -12576
rect -1406 -12708 -1398 -12576
rect -1186 -12708 -1178 -12576
rect -1178 -12708 -1140 -12576
rect -1140 -12708 -1132 -12576
rect -920 -12708 -912 -12576
rect -912 -12708 -874 -12576
rect -874 -12708 -866 -12576
rect -2782 -13718 -2774 -13586
rect -2774 -13718 -2736 -13586
rect -2736 -13718 -2728 -13586
rect -2516 -13718 -2508 -13586
rect -2508 -13718 -2470 -13586
rect -2470 -13718 -2462 -13586
rect -2250 -13718 -2242 -13586
rect -2242 -13718 -2204 -13586
rect -2204 -13718 -2196 -13586
rect -1984 -13718 -1976 -13586
rect -1976 -13718 -1938 -13586
rect -1938 -13718 -1930 -13586
rect -1718 -13718 -1710 -13586
rect -1710 -13718 -1672 -13586
rect -1672 -13718 -1664 -13586
rect -1452 -13718 -1444 -13586
rect -1444 -13718 -1406 -13586
rect -1406 -13718 -1398 -13586
rect -1186 -13718 -1178 -13586
rect -1178 -13718 -1140 -13586
rect -1140 -13718 -1132 -13586
rect -920 -13718 -912 -13586
rect -912 -13718 -874 -13586
rect -874 -13718 -866 -13586
rect -2782 -14728 -2774 -14596
rect -2774 -14728 -2736 -14596
rect -2736 -14728 -2728 -14596
rect -2516 -14728 -2508 -14596
rect -2508 -14728 -2470 -14596
rect -2470 -14728 -2462 -14596
rect -2250 -14728 -2242 -14596
rect -2242 -14728 -2204 -14596
rect -2204 -14728 -2196 -14596
rect -1984 -14728 -1976 -14596
rect -1976 -14728 -1938 -14596
rect -1938 -14728 -1930 -14596
rect -1718 -14728 -1710 -14596
rect -1710 -14728 -1672 -14596
rect -1672 -14728 -1664 -14596
rect -1452 -14728 -1444 -14596
rect -1444 -14728 -1406 -14596
rect -1406 -14728 -1398 -14596
rect -1186 -14728 -1178 -14596
rect -1178 -14728 -1140 -14596
rect -1140 -14728 -1132 -14596
rect -920 -14728 -912 -14596
rect -912 -14728 -874 -14596
rect -874 -14728 -866 -14596
rect 4366 -14724 4570 -14514
rect -2782 -15738 -2774 -15606
rect -2774 -15738 -2736 -15606
rect -2736 -15738 -2728 -15606
rect -2516 -15738 -2508 -15606
rect -2508 -15738 -2470 -15606
rect -2470 -15738 -2462 -15606
rect -2250 -15738 -2242 -15606
rect -2242 -15738 -2204 -15606
rect -2204 -15738 -2196 -15606
rect -1984 -15738 -1976 -15606
rect -1976 -15738 -1938 -15606
rect -1938 -15738 -1930 -15606
rect -1718 -15738 -1710 -15606
rect -1710 -15738 -1672 -15606
rect -1672 -15738 -1664 -15606
rect -1452 -15738 -1444 -15606
rect -1444 -15738 -1406 -15606
rect -1406 -15738 -1398 -15606
rect -1186 -15738 -1178 -15606
rect -1178 -15738 -1140 -15606
rect -1140 -15738 -1132 -15606
rect -2084 -16282 -1590 -16154
rect -920 -15738 -912 -15606
rect -912 -15738 -874 -15606
rect -874 -15738 -866 -15606
rect 4208 -16472 4520 -16136
rect -2512 -18880 -1160 -18768
rect 4340 -18854 5096 -18188
<< metal2 >>
rect -6438 -3712 -6328 -3702
rect -6438 -3794 -6328 -3784
rect -5958 -3712 -5848 -3702
rect -5958 -3794 -5848 -3784
rect -5478 -3712 -5368 -3702
rect -5478 -3794 -5368 -3784
rect -4998 -3712 -4888 -3702
rect -4998 -3794 -4888 -3784
rect -4518 -3712 -4408 -3702
rect -4518 -3794 -4408 -3784
rect -4038 -3712 -3928 -3702
rect -4038 -3794 -3928 -3784
rect -3558 -3712 -3448 -3702
rect -3558 -3794 -3448 -3784
rect -3078 -3712 -2968 -3702
rect -3078 -3794 -2968 -3784
rect -2598 -3712 -2488 -3702
rect -2598 -3794 -2488 -3784
rect -2118 -3712 -2008 -3702
rect -2118 -3794 -2008 -3784
rect -1638 -3712 -1528 -3702
rect -1638 -3794 -1528 -3784
rect -1158 -3712 -1048 -3702
rect -1158 -3794 -1048 -3784
rect -678 -3712 -568 -3702
rect -678 -3794 -568 -3784
rect -198 -3712 -88 -3702
rect -198 -3794 -88 -3784
rect 282 -3712 392 -3702
rect 282 -3794 392 -3784
rect 762 -3712 872 -3702
rect 762 -3794 872 -3784
rect 1242 -3712 1352 -3702
rect 1242 -3794 1352 -3784
rect 1722 -3712 1832 -3702
rect 1722 -3794 1832 -3784
rect 2202 -3712 2312 -3702
rect 2202 -3794 2312 -3784
rect 2682 -3712 2792 -3702
rect 2682 -3794 2792 -3784
rect 3500 -3898 3800 -3888
rect -6548 -4056 3500 -4046
rect -6548 -4188 -6538 -4056
rect -6468 -4188 -6298 -4056
rect -6228 -4188 -6058 -4056
rect -5988 -4188 -5818 -4056
rect -5748 -4188 -5578 -4056
rect -5508 -4188 -5338 -4056
rect -5268 -4188 -5098 -4056
rect -5028 -4188 -4858 -4056
rect -4788 -4188 -4618 -4056
rect -4548 -4188 -4378 -4056
rect -4308 -4188 -4138 -4056
rect -4068 -4188 -3898 -4056
rect -3828 -4188 -3658 -4056
rect -3588 -4188 -3418 -4056
rect -3348 -4188 -3178 -4056
rect -3108 -4188 -2938 -4056
rect -2868 -4188 -2698 -4056
rect -2628 -4188 -2458 -4056
rect -2388 -4188 -2218 -4056
rect -2148 -4188 -1978 -4056
rect -1908 -4188 -1738 -4056
rect -1668 -4188 -1498 -4056
rect -1428 -4188 -1258 -4056
rect -1188 -4188 -1018 -4056
rect -948 -4188 -778 -4056
rect -708 -4188 -538 -4056
rect -468 -4188 -298 -4056
rect -228 -4188 -58 -4056
rect 12 -4188 182 -4056
rect 252 -4188 422 -4056
rect 492 -4188 662 -4056
rect 732 -4188 902 -4056
rect 972 -4188 1142 -4056
rect 1212 -4188 1382 -4056
rect 1452 -4188 1622 -4056
rect 1692 -4188 1862 -4056
rect 1932 -4188 2102 -4056
rect 2172 -4188 2342 -4056
rect 2412 -4188 2582 -4056
rect 2652 -4188 2822 -4056
rect 2892 -4188 3500 -4056
rect -6548 -4198 3500 -4188
rect 3500 -4208 3800 -4198
rect 3500 -4706 3800 -4696
rect -6548 -4864 3500 -4854
rect -6548 -4996 -6538 -4864
rect -6468 -4996 -6298 -4864
rect -6228 -4996 -6058 -4864
rect -5988 -4996 -5818 -4864
rect -5748 -4996 -5578 -4864
rect -5508 -4996 -5338 -4864
rect -5268 -4996 -5098 -4864
rect -5028 -4996 -4858 -4864
rect -4788 -4996 -4618 -4864
rect -4548 -4996 -4378 -4864
rect -4308 -4996 -4138 -4864
rect -4068 -4996 -3898 -4864
rect -3828 -4996 -3658 -4864
rect -3588 -4996 -3418 -4864
rect -3348 -4996 -3178 -4864
rect -3108 -4996 -2938 -4864
rect -2868 -4996 -2698 -4864
rect -2628 -4996 -2458 -4864
rect -2388 -4996 -2218 -4864
rect -2148 -4996 -1978 -4864
rect -1908 -4996 -1738 -4864
rect -1668 -4996 -1498 -4864
rect -1428 -4996 -1258 -4864
rect -1188 -4996 -1018 -4864
rect -948 -4996 -778 -4864
rect -708 -4996 -538 -4864
rect -468 -4996 -298 -4864
rect -228 -4996 -58 -4864
rect 12 -4996 182 -4864
rect 252 -4996 422 -4864
rect 492 -4996 662 -4864
rect 732 -4996 902 -4864
rect 972 -4996 1142 -4864
rect 1212 -4996 1382 -4864
rect 1452 -4996 1622 -4864
rect 1692 -4996 1862 -4864
rect 1932 -4996 2102 -4864
rect 2172 -4996 2342 -4864
rect 2412 -4996 2582 -4864
rect 2652 -4996 2822 -4864
rect 2892 -4996 3500 -4864
rect -6548 -5006 3500 -4996
rect 3500 -5016 3800 -5006
rect 3500 -5514 3800 -5504
rect -6548 -5672 3500 -5662
rect -6548 -5804 -6538 -5672
rect -6468 -5804 -6298 -5672
rect -6228 -5804 -6058 -5672
rect -5988 -5804 -5818 -5672
rect -5748 -5804 -5578 -5672
rect -5508 -5804 -5338 -5672
rect -5268 -5804 -5098 -5672
rect -5028 -5804 -4858 -5672
rect -4788 -5804 -4618 -5672
rect -4548 -5804 -4378 -5672
rect -4308 -5804 -4138 -5672
rect -4068 -5804 -3898 -5672
rect -3828 -5804 -3658 -5672
rect -3588 -5804 -3418 -5672
rect -3348 -5804 -3178 -5672
rect -3108 -5804 -2938 -5672
rect -2868 -5804 -2698 -5672
rect -2628 -5804 -2458 -5672
rect -2388 -5804 -2218 -5672
rect -2148 -5804 -1978 -5672
rect -1908 -5804 -1738 -5672
rect -1668 -5804 -1498 -5672
rect -1428 -5804 -1258 -5672
rect -1188 -5804 -1018 -5672
rect -948 -5804 -778 -5672
rect -708 -5804 -538 -5672
rect -468 -5804 -298 -5672
rect -228 -5804 -58 -5672
rect 12 -5804 182 -5672
rect 252 -5804 422 -5672
rect 492 -5804 662 -5672
rect 732 -5804 902 -5672
rect 972 -5804 1142 -5672
rect 1212 -5804 1382 -5672
rect 1452 -5804 1622 -5672
rect 1692 -5804 1862 -5672
rect 1932 -5804 2102 -5672
rect 2172 -5804 2342 -5672
rect 2412 -5804 2582 -5672
rect 2652 -5804 2822 -5672
rect 2892 -5804 3500 -5672
rect -6548 -5814 3500 -5804
rect 3500 -5824 3800 -5814
rect 7404 -6698 8304 -6688
rect 7404 -7206 8304 -7196
rect -15442 -11450 -15254 -11440
rect -15442 -11570 -15254 -11560
rect -14266 -11450 -14078 -11440
rect -14266 -11570 -14078 -11560
rect -13090 -11450 -12902 -11440
rect -13090 -11570 -12902 -11560
rect -11914 -11450 -11726 -11440
rect -11914 -11570 -11726 -11560
rect -10738 -11450 -10550 -11440
rect -10738 -11570 -10550 -11560
rect -9562 -11450 -9374 -11440
rect -9562 -11570 -9374 -11560
rect -8386 -11450 -8198 -11440
rect -8386 -11570 -8198 -11560
rect -7210 -11450 -7022 -11440
rect -7210 -11570 -7022 -11560
rect -6034 -11450 -5846 -11440
rect -6034 -11570 -5846 -11560
rect -4858 -11450 -4670 -11440
rect -4858 -11570 -4670 -11560
rect -3682 -11450 -3494 -11440
rect -3682 -11570 -3494 -11560
rect -2506 -11450 -2318 -11440
rect -2506 -11570 -2318 -11560
rect -1330 -11450 -1142 -11440
rect -1330 -11570 -1142 -11560
rect -154 -11450 34 -11440
rect -154 -11570 34 -11560
rect 1022 -11450 1210 -11440
rect 1022 -11570 1210 -11560
rect 2198 -11450 2386 -11440
rect 2198 -11570 2386 -11560
rect 4550 -11450 4738 -11440
rect 4550 -11570 4738 -11560
rect 5726 -11450 5914 -11440
rect 5726 -11570 5914 -11560
rect 6902 -11450 7090 -11440
rect 6902 -11570 7090 -11560
rect 9254 -11450 9442 -11440
rect 9254 -11570 9442 -11560
rect 10430 -11450 10618 -11440
rect 10430 -11570 10618 -11560
rect 11606 -11450 11794 -11440
rect 11606 -11570 11794 -11560
rect -2250 -12452 -72 -12326
rect -2250 -12566 -1930 -12452
rect -2782 -12576 -2462 -12566
rect -2728 -12708 -2516 -12576
rect -2782 -12832 -2462 -12708
rect -2250 -12576 -2196 -12566
rect -2250 -12718 -2196 -12708
rect -1984 -12576 -1930 -12566
rect -1984 -12718 -1930 -12708
rect -1718 -12576 -1398 -12452
rect -1664 -12708 -1452 -12576
rect -1718 -12714 -1398 -12708
rect -1186 -12576 -1132 -12566
rect -1186 -12714 -1132 -12708
rect -920 -12576 -866 -12566
rect -920 -12714 -866 -12708
rect -1186 -12832 -866 -12714
rect -3576 -12958 -866 -12832
rect -3576 -13842 -3328 -12958
rect -320 -13336 -72 -12452
rect -2250 -13462 -72 -13336
rect -2250 -13576 -1930 -13462
rect -1710 -13576 -1390 -13462
rect -2782 -13586 -2728 -13576
rect -2782 -13728 -2728 -13718
rect -2516 -13586 -2462 -13576
rect -2516 -13728 -2462 -13718
rect -2250 -13586 -2196 -13576
rect -2250 -13728 -2196 -13718
rect -1984 -13586 -1930 -13576
rect -1984 -13728 -1930 -13718
rect -1718 -13586 -1664 -13576
rect -1718 -13728 -1664 -13718
rect -1452 -13586 -1398 -13576
rect -1452 -13728 -1398 -13718
rect -1186 -13586 -1132 -13576
rect -1186 -13728 -1132 -13718
rect -920 -13586 -866 -13576
rect -920 -13728 -866 -13718
rect -2782 -13842 -2462 -13728
rect -1186 -13842 -866 -13728
rect -3576 -13968 -866 -13842
rect -3576 -14852 -3328 -13968
rect -320 -14346 -72 -13462
rect -2250 -14472 -72 -14346
rect -2250 -14586 -1930 -14472
rect -2782 -14596 -2728 -14586
rect -2782 -14738 -2728 -14728
rect -2516 -14596 -2462 -14586
rect -2516 -14738 -2462 -14728
rect -2250 -14596 -2196 -14586
rect -2250 -14738 -2196 -14728
rect -1984 -14596 -1930 -14586
rect -1984 -14738 -1930 -14728
rect -1718 -14590 -1398 -14472
rect -1718 -14596 -1664 -14590
rect -1718 -14738 -1664 -14728
rect -1452 -14596 -1398 -14590
rect -1452 -14738 -1398 -14728
rect -1186 -14596 -1132 -14586
rect -1186 -14738 -1132 -14728
rect -920 -14596 -866 -14586
rect -920 -14738 -866 -14728
rect -2782 -14852 -2462 -14738
rect -1186 -14852 -866 -14738
rect -3576 -14978 -866 -14852
rect -3576 -15862 -3328 -14978
rect -320 -15356 -72 -14472
rect 5594 -14382 5894 -14370
rect 4366 -14514 4570 -14504
rect 4570 -14682 5594 -14516
rect 5594 -14692 5894 -14682
rect 4366 -14734 4570 -14724
rect -2250 -15482 -72 -15356
rect -2250 -15596 -1930 -15482
rect -2782 -15606 -2728 -15596
rect -2782 -15748 -2728 -15738
rect -2516 -15606 -2462 -15596
rect -2516 -15748 -2462 -15738
rect -2250 -15606 -2196 -15596
rect -2250 -15748 -2196 -15738
rect -1984 -15606 -1930 -15596
rect -1984 -15748 -1930 -15738
rect -1718 -15596 -1398 -15482
rect -1718 -15606 -1664 -15596
rect -1718 -15748 -1664 -15738
rect -1452 -15606 -1398 -15596
rect -1452 -15748 -1398 -15738
rect -1186 -15606 -1132 -15596
rect -1186 -15748 -1132 -15738
rect -920 -15606 -866 -15596
rect -920 -15748 -866 -15738
rect -2782 -15862 -2462 -15748
rect -1186 -15862 -866 -15748
rect -3576 -15988 -866 -15862
rect 3510 -15992 3810 -15982
rect -2084 -16154 3510 -16144
rect -1590 -16282 3510 -16154
rect -2084 -16292 3510 -16282
rect 4208 -16136 4520 -16126
rect 3810 -16292 4208 -16144
rect 3510 -16302 3810 -16292
rect 4208 -16482 4520 -16472
rect 4340 -18188 5096 -18178
rect -2512 -18768 -1160 -18758
rect 4340 -18864 5096 -18854
rect -2512 -18890 -1160 -18880
<< via2 >>
rect -6438 -3784 -6328 -3712
rect -5958 -3784 -5848 -3712
rect -5478 -3784 -5368 -3712
rect -4998 -3784 -4888 -3712
rect -4518 -3784 -4408 -3712
rect -4038 -3784 -3928 -3712
rect -3558 -3784 -3448 -3712
rect -3078 -3784 -2968 -3712
rect -2598 -3784 -2488 -3712
rect -2118 -3784 -2008 -3712
rect -1638 -3784 -1528 -3712
rect -1158 -3784 -1048 -3712
rect -678 -3784 -568 -3712
rect -198 -3784 -88 -3712
rect 282 -3784 392 -3712
rect 762 -3784 872 -3712
rect 1242 -3784 1352 -3712
rect 1722 -3784 1832 -3712
rect 2202 -3784 2312 -3712
rect 2682 -3784 2792 -3712
rect 3500 -4198 3800 -3898
rect 3500 -5006 3800 -4706
rect 3500 -5814 3800 -5514
rect 7404 -7196 8304 -6698
rect -15442 -11560 -15254 -11450
rect -14266 -11560 -14078 -11450
rect -13090 -11560 -12902 -11450
rect -11914 -11560 -11726 -11450
rect -10738 -11560 -10550 -11450
rect -9562 -11560 -9374 -11450
rect -8386 -11560 -8198 -11450
rect -7210 -11560 -7022 -11450
rect -6034 -11560 -5846 -11450
rect -4858 -11560 -4670 -11450
rect -3682 -11560 -3494 -11450
rect -2506 -11560 -2318 -11450
rect -1330 -11560 -1142 -11450
rect -154 -11560 34 -11450
rect 1022 -11560 1210 -11450
rect 2198 -11560 2386 -11450
rect 4550 -11560 4738 -11450
rect 5726 -11560 5914 -11450
rect 6902 -11560 7090 -11450
rect 9254 -11560 9442 -11450
rect 10430 -11560 10618 -11450
rect 11606 -11560 11794 -11450
rect 5594 -14682 5894 -14382
rect 3510 -16292 3810 -15992
rect -2512 -18880 -1160 -18768
rect 4340 -18854 5096 -18188
<< metal3 >>
rect -6448 -3712 -6318 -3707
rect -6448 -3784 -6438 -3712
rect -6328 -3784 -6318 -3712
rect -6448 -3789 -6318 -3784
rect -5968 -3712 -5838 -3707
rect -5968 -3784 -5958 -3712
rect -5848 -3784 -5838 -3712
rect -5968 -3789 -5838 -3784
rect -5488 -3712 -5358 -3707
rect -5488 -3784 -5478 -3712
rect -5368 -3784 -5358 -3712
rect -5488 -3789 -5358 -3784
rect -5008 -3712 -4878 -3707
rect -5008 -3784 -4998 -3712
rect -4888 -3784 -4878 -3712
rect -5008 -3789 -4878 -3784
rect -4528 -3712 -4398 -3707
rect -4528 -3784 -4518 -3712
rect -4408 -3784 -4398 -3712
rect -4528 -3789 -4398 -3784
rect -4048 -3712 -3918 -3707
rect -4048 -3784 -4038 -3712
rect -3928 -3784 -3918 -3712
rect -4048 -3789 -3918 -3784
rect -3568 -3712 -3438 -3707
rect -3568 -3784 -3558 -3712
rect -3448 -3784 -3438 -3712
rect -3568 -3789 -3438 -3784
rect -3088 -3712 -2958 -3707
rect -3088 -3784 -3078 -3712
rect -2968 -3784 -2958 -3712
rect -3088 -3789 -2958 -3784
rect -2608 -3712 -2478 -3707
rect -2608 -3784 -2598 -3712
rect -2488 -3784 -2478 -3712
rect -2608 -3789 -2478 -3784
rect -2128 -3712 -1998 -3707
rect -2128 -3784 -2118 -3712
rect -2008 -3784 -1998 -3712
rect -2128 -3789 -1998 -3784
rect -1648 -3712 -1518 -3707
rect -1648 -3784 -1638 -3712
rect -1528 -3784 -1518 -3712
rect -1648 -3789 -1518 -3784
rect -1168 -3712 -1038 -3707
rect -1168 -3784 -1158 -3712
rect -1048 -3784 -1038 -3712
rect -1168 -3789 -1038 -3784
rect -688 -3712 -558 -3707
rect -688 -3784 -678 -3712
rect -568 -3784 -558 -3712
rect -688 -3789 -558 -3784
rect -208 -3712 -78 -3707
rect -208 -3784 -198 -3712
rect -88 -3784 -78 -3712
rect -208 -3789 -78 -3784
rect 272 -3712 402 -3707
rect 272 -3784 282 -3712
rect 392 -3784 402 -3712
rect 272 -3789 402 -3784
rect 752 -3712 882 -3707
rect 752 -3784 762 -3712
rect 872 -3784 882 -3712
rect 752 -3789 882 -3784
rect 1232 -3712 1362 -3707
rect 1232 -3784 1242 -3712
rect 1352 -3784 1362 -3712
rect 1232 -3789 1362 -3784
rect 1712 -3712 1842 -3707
rect 1712 -3784 1722 -3712
rect 1832 -3784 1842 -3712
rect 1712 -3789 1842 -3784
rect 2192 -3712 2322 -3707
rect 2192 -3784 2202 -3712
rect 2312 -3784 2322 -3712
rect 2192 -3789 2322 -3784
rect 2672 -3712 2802 -3707
rect 2672 -3784 2682 -3712
rect 2792 -3784 2802 -3712
rect 2672 -3789 2802 -3784
rect 3490 -3894 3810 -3893
rect 3490 -3898 3820 -3894
rect 3490 -4198 3500 -3898
rect 3800 -4198 3820 -3898
rect 3490 -4203 3820 -4198
rect 3500 -4701 3820 -4203
rect 3490 -4706 3820 -4701
rect 3490 -5006 3500 -4706
rect 3800 -5006 3820 -4706
rect 3490 -5011 3820 -5006
rect 3500 -5509 3820 -5011
rect 3490 -5514 3820 -5509
rect 3490 -5814 3500 -5514
rect 3800 -5814 3820 -5514
rect 3490 -5819 3820 -5814
rect -15452 -11450 -15244 -11445
rect -15452 -11560 -15442 -11450
rect -15254 -11560 -15244 -11450
rect -15452 -11565 -15244 -11560
rect -14276 -11450 -14068 -11445
rect -14276 -11560 -14266 -11450
rect -14078 -11560 -14068 -11450
rect -14276 -11565 -14068 -11560
rect -13100 -11450 -12892 -11445
rect -13100 -11560 -13090 -11450
rect -12902 -11560 -12892 -11450
rect -13100 -11565 -12892 -11560
rect -11924 -11450 -11716 -11445
rect -11924 -11560 -11914 -11450
rect -11726 -11560 -11716 -11450
rect -11924 -11565 -11716 -11560
rect -10748 -11450 -10540 -11445
rect -10748 -11560 -10738 -11450
rect -10550 -11560 -10540 -11450
rect -10748 -11565 -10540 -11560
rect -9572 -11450 -9364 -11445
rect -9572 -11560 -9562 -11450
rect -9374 -11560 -9364 -11450
rect -9572 -11565 -9364 -11560
rect -8396 -11450 -8188 -11445
rect -8396 -11560 -8386 -11450
rect -8198 -11560 -8188 -11450
rect -8396 -11565 -8188 -11560
rect -7220 -11450 -7012 -11445
rect -7220 -11560 -7210 -11450
rect -7022 -11560 -7012 -11450
rect -7220 -11565 -7012 -11560
rect -6044 -11450 -5836 -11445
rect -6044 -11560 -6034 -11450
rect -5846 -11560 -5836 -11450
rect -6044 -11565 -5836 -11560
rect -4868 -11450 -4660 -11445
rect -4868 -11560 -4858 -11450
rect -4670 -11560 -4660 -11450
rect -4868 -11565 -4660 -11560
rect -3692 -11450 -3484 -11445
rect -3692 -11560 -3682 -11450
rect -3494 -11560 -3484 -11450
rect -3692 -11565 -3484 -11560
rect -2516 -11450 -2308 -11445
rect -2516 -11560 -2506 -11450
rect -2318 -11560 -2308 -11450
rect -2516 -11565 -2308 -11560
rect -1340 -11450 -1132 -11445
rect -1340 -11560 -1330 -11450
rect -1142 -11560 -1132 -11450
rect -1340 -11565 -1132 -11560
rect -164 -11450 44 -11445
rect -164 -11560 -154 -11450
rect 34 -11560 44 -11450
rect -164 -11565 44 -11560
rect 1012 -11450 1220 -11445
rect 1012 -11560 1022 -11450
rect 1210 -11560 1220 -11450
rect 1012 -11565 1220 -11560
rect 2188 -11450 2396 -11445
rect 2188 -11560 2198 -11450
rect 2386 -11560 2396 -11450
rect 2188 -11565 2396 -11560
rect 3500 -15992 3820 -5819
rect 7394 -6698 8314 -6693
rect 7394 -7196 7404 -6698
rect 8304 -7196 8314 -6698
rect 7394 -7201 8314 -7196
rect 4540 -11450 4748 -11445
rect 4540 -11560 4550 -11450
rect 4738 -11560 4748 -11450
rect 4540 -11565 4748 -11560
rect 5716 -11450 5924 -11445
rect 5716 -11560 5726 -11450
rect 5914 -11560 5924 -11450
rect 5716 -11565 5924 -11560
rect 6892 -11450 7100 -11445
rect 6892 -11560 6902 -11450
rect 7090 -11560 7100 -11450
rect 6892 -11565 7100 -11560
rect 7448 -12458 8286 -7201
rect 9244 -11450 9452 -11445
rect 9244 -11560 9254 -11450
rect 9442 -11560 9452 -11450
rect 9244 -11565 9452 -11560
rect 10420 -11450 10628 -11445
rect 10420 -11560 10430 -11450
rect 10618 -11560 10628 -11450
rect 10420 -11565 10628 -11560
rect 11596 -11450 11804 -11445
rect 11596 -11560 11606 -11450
rect 11794 -11560 11804 -11450
rect 11596 -11565 11804 -11560
rect 7410 -13358 7420 -12458
rect 8320 -13358 8330 -12458
rect 6484 -14376 9384 -13508
rect 5584 -14382 9384 -14376
rect 5584 -14682 5594 -14382
rect 5894 -14682 9384 -14382
rect 5584 -14688 9384 -14682
rect 3500 -16292 3510 -15992
rect 3810 -16292 3820 -15992
rect 3500 -16297 3820 -16292
rect 6484 -16406 9384 -14688
rect 4330 -18188 5106 -18183
rect -2522 -18768 -1150 -18763
rect -2522 -18880 -2512 -18768
rect -1160 -18880 -1150 -18768
rect 4330 -18854 4340 -18188
rect 5096 -18854 5106 -18188
rect 4330 -18859 5106 -18854
rect -2522 -18885 -1150 -18880
<< via3 >>
rect -6438 -3784 -6328 -3712
rect -5958 -3784 -5848 -3712
rect -5478 -3784 -5368 -3712
rect -4998 -3784 -4888 -3712
rect -4518 -3784 -4408 -3712
rect -4038 -3784 -3928 -3712
rect -3558 -3784 -3448 -3712
rect -3078 -3784 -2968 -3712
rect -2598 -3784 -2488 -3712
rect -2118 -3784 -2008 -3712
rect -1638 -3784 -1528 -3712
rect -1158 -3784 -1048 -3712
rect -678 -3784 -568 -3712
rect -198 -3784 -88 -3712
rect 282 -3784 392 -3712
rect 762 -3784 872 -3712
rect 1242 -3784 1352 -3712
rect 1722 -3784 1832 -3712
rect 2202 -3784 2312 -3712
rect 2682 -3784 2792 -3712
rect -15442 -11560 -15254 -11450
rect -14266 -11560 -14078 -11450
rect -13090 -11560 -12902 -11450
rect -11914 -11560 -11726 -11450
rect -10738 -11560 -10550 -11450
rect -9562 -11560 -9374 -11450
rect -8386 -11560 -8198 -11450
rect -7210 -11560 -7022 -11450
rect -6034 -11560 -5846 -11450
rect -4858 -11560 -4670 -11450
rect -3682 -11560 -3494 -11450
rect -2506 -11560 -2318 -11450
rect -1330 -11560 -1142 -11450
rect -154 -11560 34 -11450
rect 1022 -11560 1210 -11450
rect 2198 -11560 2386 -11450
rect 4550 -11560 4738 -11450
rect 5726 -11560 5914 -11450
rect 6902 -11560 7090 -11450
rect 9254 -11560 9442 -11450
rect 10430 -11560 10618 -11450
rect 11606 -11560 11794 -11450
rect 7420 -13358 8320 -12458
rect -2512 -18880 -1160 -18768
rect 4340 -18854 5096 -18188
<< mimcap >>
rect 6584 -13646 9284 -13606
rect 6584 -16266 6624 -13646
rect 9244 -16266 9284 -13646
rect 6584 -16306 9284 -16266
<< mimcapcontact >>
rect 6624 -16266 9244 -13646
<< metal4 >>
rect -18126 -3080 9244 -3006
rect -19208 -3712 9244 -3080
rect -19208 -3784 -6438 -3712
rect -6328 -3784 -5958 -3712
rect -5848 -3784 -5478 -3712
rect -5368 -3784 -4998 -3712
rect -4888 -3784 -4518 -3712
rect -4408 -3784 -4038 -3712
rect -3928 -3784 -3558 -3712
rect -3448 -3784 -3078 -3712
rect -2968 -3784 -2598 -3712
rect -2488 -3784 -2118 -3712
rect -2008 -3784 -1638 -3712
rect -1528 -3784 -1158 -3712
rect -1048 -3784 -678 -3712
rect -568 -3784 -198 -3712
rect -88 -3784 282 -3712
rect 392 -3784 762 -3712
rect 872 -3784 1242 -3712
rect 1352 -3784 1722 -3712
rect 1832 -3784 2202 -3712
rect 2312 -3784 2682 -3712
rect 2792 -3784 9244 -3712
rect -19208 -4270 9244 -3784
rect -19208 -4272 -12590 -4270
rect -19208 -17874 -17826 -4272
rect -17466 -11450 12858 -10586
rect -17466 -11560 -15442 -11450
rect -15254 -11560 -14266 -11450
rect -14078 -11560 -13090 -11450
rect -12902 -11560 -11914 -11450
rect -11726 -11560 -10738 -11450
rect -10550 -11560 -9562 -11450
rect -9374 -11560 -8386 -11450
rect -8198 -11560 -7210 -11450
rect -7022 -11560 -6034 -11450
rect -5846 -11560 -4858 -11450
rect -4670 -11560 -3682 -11450
rect -3494 -11560 -2506 -11450
rect -2318 -11560 -1330 -11450
rect -1142 -11560 -154 -11450
rect 34 -11560 1022 -11450
rect 1210 -11560 2198 -11450
rect 2386 -11560 4550 -11450
rect 4738 -11560 5726 -11450
rect 5914 -11560 6902 -11450
rect 7090 -11560 9254 -11450
rect 9442 -11560 10430 -11450
rect 10618 -11560 11606 -11450
rect 11794 -11560 12858 -11450
rect -17466 -12118 12858 -11560
rect 7419 -12458 8321 -12457
rect 7419 -13358 7420 -12458
rect 8320 -13358 8321 -12458
rect 7419 -13359 8321 -13358
rect 7476 -13644 8278 -13359
rect 6622 -13646 9246 -13644
rect 6622 -16266 6624 -13646
rect 9244 -16266 9246 -13646
rect 6622 -16268 9246 -16266
rect -19208 -18188 12858 -17874
rect -19208 -18768 4340 -18188
rect -19208 -18880 -2512 -18768
rect -1160 -18854 4340 -18768
rect 5096 -18854 12858 -18188
rect -1160 -18880 12858 -18854
rect -19208 -19406 12858 -18880
rect -19208 -19408 -17826 -19406
<< labels >>
flabel metal1 10808 -7008 10808 -7008 0 FreeSans 1600 0 0 0 vout
port 5 nsew
flabel metal1 -15668 -10204 -15668 -10204 0 FreeSans 1600 0 0 0 vbias
port 3 nsew
flabel metal2 -3484 -14186 -3484 -14186 0 FreeSans 1600 0 0 0 vn
port 2 nsew
flabel metal2 -236 -13718 -236 -13718 0 FreeSans 1600 0 0 0 vp
port 1 nsew
flabel metal4 -17004 -11600 -17004 -11600 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal4 -16806 -18734 -16806 -18734 0 FreeSans 1600 0 0 0 vss
port 4 nsew
<< end >>
