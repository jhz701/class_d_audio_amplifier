magic
tech sky130A
magscale 1 2
timestamp 1629189117
<< nwell >>
rect 28625 10221 40749 12331
rect 30113 5597 33309 9943
<< pwell >>
rect 33740 6168 34142 7644
rect 30113 3375 39261 5249
<< pmoslvt >>
rect 28821 11712 29021 12112
rect 29193 11712 29393 12112
rect 29565 11712 29765 12112
rect 29937 11712 30137 12112
rect 30309 11712 30509 12112
rect 30681 11712 30881 12112
rect 31053 11712 31253 12112
rect 31425 11712 31625 12112
rect 31797 11712 31997 12112
rect 32169 11712 32369 12112
rect 32541 11712 32741 12112
rect 32913 11712 33113 12112
rect 33285 11712 33485 12112
rect 33657 11712 33857 12112
rect 34029 11712 34229 12112
rect 34401 11712 34601 12112
rect 34773 11712 34973 12112
rect 35145 11712 35345 12112
rect 35517 11712 35717 12112
rect 35889 11712 36089 12112
rect 36261 11712 36461 12112
rect 36633 11712 36833 12112
rect 37005 11712 37205 12112
rect 37377 11712 37577 12112
rect 37749 11712 37949 12112
rect 38121 11712 38321 12112
rect 38493 11712 38693 12112
rect 38865 11712 39065 12112
rect 39237 11712 39437 12112
rect 39609 11712 39809 12112
rect 39981 11712 40181 12112
rect 40353 11712 40553 12112
rect 28821 11076 29021 11476
rect 29193 11076 29393 11476
rect 29565 11076 29765 11476
rect 29937 11076 30137 11476
rect 30309 11076 30509 11476
rect 30681 11076 30881 11476
rect 31053 11076 31253 11476
rect 31425 11076 31625 11476
rect 31797 11076 31997 11476
rect 32169 11076 32369 11476
rect 32541 11076 32741 11476
rect 32913 11076 33113 11476
rect 33285 11076 33485 11476
rect 33657 11076 33857 11476
rect 34029 11076 34229 11476
rect 34401 11076 34601 11476
rect 34773 11076 34973 11476
rect 35145 11076 35345 11476
rect 35517 11076 35717 11476
rect 35889 11076 36089 11476
rect 36261 11076 36461 11476
rect 36633 11076 36833 11476
rect 37005 11076 37205 11476
rect 37377 11076 37577 11476
rect 37749 11076 37949 11476
rect 38121 11076 38321 11476
rect 38493 11076 38693 11476
rect 38865 11076 39065 11476
rect 39237 11076 39437 11476
rect 39609 11076 39809 11476
rect 39981 11076 40181 11476
rect 40353 11076 40553 11476
rect 28821 10440 29021 10840
rect 29193 10440 29393 10840
rect 29565 10440 29765 10840
rect 29937 10440 30137 10840
rect 30309 10440 30509 10840
rect 30681 10440 30881 10840
rect 31053 10440 31253 10840
rect 31425 10440 31625 10840
rect 31797 10440 31997 10840
rect 32169 10440 32369 10840
rect 32541 10440 32741 10840
rect 32913 10440 33113 10840
rect 33285 10440 33485 10840
rect 33657 10440 33857 10840
rect 34029 10440 34229 10840
rect 34401 10440 34601 10840
rect 34773 10440 34973 10840
rect 35145 10440 35345 10840
rect 35517 10440 35717 10840
rect 35889 10440 36089 10840
rect 36261 10440 36461 10840
rect 36633 10440 36833 10840
rect 37005 10440 37205 10840
rect 37377 10440 37577 10840
rect 37749 10440 37949 10840
rect 38121 10440 38321 10840
rect 38493 10440 38693 10840
rect 38865 10440 39065 10840
rect 39237 10440 39437 10840
rect 39609 10440 39809 10840
rect 39981 10440 40181 10840
rect 40353 10440 40553 10840
rect 30309 8924 30509 9724
rect 30681 8924 30881 9724
rect 31053 8924 31253 9724
rect 31425 8924 31625 9724
rect 31797 8924 31997 9724
rect 32169 8924 32369 9724
rect 32541 8924 32741 9724
rect 32913 8924 33113 9724
rect 30309 7888 30509 8688
rect 30681 7888 30881 8688
rect 31053 7888 31253 8688
rect 31425 7888 31625 8688
rect 31797 7888 31997 8688
rect 32169 7888 32369 8688
rect 32541 7888 32741 8688
rect 32913 7888 33113 8688
rect 30309 6852 30509 7652
rect 30681 6852 30881 7652
rect 31053 6852 31253 7652
rect 31425 6852 31625 7652
rect 31797 6852 31997 7652
rect 32169 6852 32369 7652
rect 32541 6852 32741 7652
rect 32913 6852 33113 7652
rect 30309 5816 30509 6616
rect 30681 5816 30881 6616
rect 31053 5816 31253 6616
rect 31425 5816 31625 6616
rect 31797 5816 31997 6616
rect 32169 5816 32369 6616
rect 32541 5816 32741 6616
rect 32913 5816 33113 6616
<< nmoslvt >>
rect 30309 4839 30509 5039
rect 30681 4839 30881 5039
rect 31053 4839 31253 5039
rect 31425 4839 31625 5039
rect 31797 4839 31997 5039
rect 32169 4839 32369 5039
rect 32541 4839 32741 5039
rect 32913 4839 33113 5039
rect 33285 4839 33485 5039
rect 33657 4839 33857 5039
rect 34029 4839 34229 5039
rect 34401 4839 34601 5039
rect 34773 4839 34973 5039
rect 35145 4839 35345 5039
rect 35517 4839 35717 5039
rect 35889 4839 36089 5039
rect 36261 4839 36461 5039
rect 36633 4839 36833 5039
rect 37005 4839 37205 5039
rect 37377 4839 37577 5039
rect 37749 4839 37949 5039
rect 38121 4839 38321 5039
rect 38493 4839 38693 5039
rect 38865 4839 39065 5039
rect 30309 4421 30509 4621
rect 30681 4421 30881 4621
rect 31053 4421 31253 4621
rect 31425 4421 31625 4621
rect 31797 4421 31997 4621
rect 32169 4421 32369 4621
rect 32541 4421 32741 4621
rect 32913 4421 33113 4621
rect 33285 4421 33485 4621
rect 33657 4421 33857 4621
rect 34029 4421 34229 4621
rect 34401 4421 34601 4621
rect 34773 4421 34973 4621
rect 35145 4421 35345 4621
rect 35517 4421 35717 4621
rect 35889 4421 36089 4621
rect 36261 4421 36461 4621
rect 36633 4421 36833 4621
rect 37005 4421 37205 4621
rect 37377 4421 37577 4621
rect 37749 4421 37949 4621
rect 38121 4421 38321 4621
rect 38493 4421 38693 4621
rect 38865 4421 39065 4621
rect 30309 4003 30509 4203
rect 30681 4003 30881 4203
rect 31053 4003 31253 4203
rect 31425 4003 31625 4203
rect 31797 4003 31997 4203
rect 32169 4003 32369 4203
rect 32541 4003 32741 4203
rect 32913 4003 33113 4203
rect 33285 4003 33485 4203
rect 33657 4003 33857 4203
rect 34029 4003 34229 4203
rect 34401 4003 34601 4203
rect 34773 4003 34973 4203
rect 35145 4003 35345 4203
rect 35517 4003 35717 4203
rect 35889 4003 36089 4203
rect 36261 4003 36461 4203
rect 36633 4003 36833 4203
rect 37005 4003 37205 4203
rect 37377 4003 37577 4203
rect 37749 4003 37949 4203
rect 38121 4003 38321 4203
rect 38493 4003 38693 4203
rect 38865 4003 39065 4203
rect 30309 3585 30509 3785
rect 30681 3585 30881 3785
rect 31053 3585 31253 3785
rect 31425 3585 31625 3785
rect 31797 3585 31997 3785
rect 32169 3585 32369 3785
rect 32541 3585 32741 3785
rect 32913 3585 33113 3785
rect 33285 3585 33485 3785
rect 33657 3585 33857 3785
rect 34029 3585 34229 3785
rect 34401 3585 34601 3785
rect 34773 3585 34973 3785
rect 35145 3585 35345 3785
rect 35517 3585 35717 3785
rect 35889 3585 36089 3785
rect 36261 3585 36461 3785
rect 36633 3585 36833 3785
rect 37005 3585 37205 3785
rect 37377 3585 37577 3785
rect 37749 3585 37949 3785
rect 38121 3585 38321 3785
rect 38493 3585 38693 3785
rect 38865 3585 39065 3785
<< ndiff >>
rect 30251 5027 30309 5039
rect 30251 4851 30263 5027
rect 30297 4851 30309 5027
rect 30251 4839 30309 4851
rect 30509 5027 30567 5039
rect 30509 4851 30521 5027
rect 30555 4851 30567 5027
rect 30509 4839 30567 4851
rect 30623 5027 30681 5039
rect 30623 4851 30635 5027
rect 30669 4851 30681 5027
rect 30623 4839 30681 4851
rect 30881 5027 30939 5039
rect 30881 4851 30893 5027
rect 30927 4851 30939 5027
rect 30881 4839 30939 4851
rect 30995 5027 31053 5039
rect 30995 4851 31007 5027
rect 31041 4851 31053 5027
rect 30995 4839 31053 4851
rect 31253 5027 31311 5039
rect 31253 4851 31265 5027
rect 31299 4851 31311 5027
rect 31253 4839 31311 4851
rect 31367 5027 31425 5039
rect 31367 4851 31379 5027
rect 31413 4851 31425 5027
rect 31367 4839 31425 4851
rect 31625 5027 31683 5039
rect 31625 4851 31637 5027
rect 31671 4851 31683 5027
rect 31625 4839 31683 4851
rect 31739 5027 31797 5039
rect 31739 4851 31751 5027
rect 31785 4851 31797 5027
rect 31739 4839 31797 4851
rect 31997 5027 32055 5039
rect 31997 4851 32009 5027
rect 32043 4851 32055 5027
rect 31997 4839 32055 4851
rect 32111 5027 32169 5039
rect 32111 4851 32123 5027
rect 32157 4851 32169 5027
rect 32111 4839 32169 4851
rect 32369 5027 32427 5039
rect 32369 4851 32381 5027
rect 32415 4851 32427 5027
rect 32369 4839 32427 4851
rect 32483 5027 32541 5039
rect 32483 4851 32495 5027
rect 32529 4851 32541 5027
rect 32483 4839 32541 4851
rect 32741 5027 32799 5039
rect 32741 4851 32753 5027
rect 32787 4851 32799 5027
rect 32741 4839 32799 4851
rect 32855 5027 32913 5039
rect 32855 4851 32867 5027
rect 32901 4851 32913 5027
rect 32855 4839 32913 4851
rect 33113 5027 33171 5039
rect 33113 4851 33125 5027
rect 33159 4851 33171 5027
rect 33113 4839 33171 4851
rect 33227 5027 33285 5039
rect 33227 4851 33239 5027
rect 33273 4851 33285 5027
rect 33227 4839 33285 4851
rect 33485 5027 33543 5039
rect 33485 4851 33497 5027
rect 33531 4851 33543 5027
rect 33485 4839 33543 4851
rect 33599 5027 33657 5039
rect 33599 4851 33611 5027
rect 33645 4851 33657 5027
rect 33599 4839 33657 4851
rect 33857 5027 33915 5039
rect 33857 4851 33869 5027
rect 33903 4851 33915 5027
rect 33857 4839 33915 4851
rect 33971 5027 34029 5039
rect 33971 4851 33983 5027
rect 34017 4851 34029 5027
rect 33971 4839 34029 4851
rect 34229 5027 34287 5039
rect 34229 4851 34241 5027
rect 34275 4851 34287 5027
rect 34229 4839 34287 4851
rect 34343 5027 34401 5039
rect 34343 4851 34355 5027
rect 34389 4851 34401 5027
rect 34343 4839 34401 4851
rect 34601 5027 34659 5039
rect 34601 4851 34613 5027
rect 34647 4851 34659 5027
rect 34601 4839 34659 4851
rect 34715 5027 34773 5039
rect 34715 4851 34727 5027
rect 34761 4851 34773 5027
rect 34715 4839 34773 4851
rect 34973 5027 35031 5039
rect 34973 4851 34985 5027
rect 35019 4851 35031 5027
rect 34973 4839 35031 4851
rect 35087 5027 35145 5039
rect 35087 4851 35099 5027
rect 35133 4851 35145 5027
rect 35087 4839 35145 4851
rect 35345 5027 35403 5039
rect 35345 4851 35357 5027
rect 35391 4851 35403 5027
rect 35345 4839 35403 4851
rect 35459 5027 35517 5039
rect 35459 4851 35471 5027
rect 35505 4851 35517 5027
rect 35459 4839 35517 4851
rect 35717 5027 35775 5039
rect 35717 4851 35729 5027
rect 35763 4851 35775 5027
rect 35717 4839 35775 4851
rect 35831 5027 35889 5039
rect 35831 4851 35843 5027
rect 35877 4851 35889 5027
rect 35831 4839 35889 4851
rect 36089 5027 36147 5039
rect 36089 4851 36101 5027
rect 36135 4851 36147 5027
rect 36089 4839 36147 4851
rect 36203 5027 36261 5039
rect 36203 4851 36215 5027
rect 36249 4851 36261 5027
rect 36203 4839 36261 4851
rect 36461 5027 36519 5039
rect 36461 4851 36473 5027
rect 36507 4851 36519 5027
rect 36461 4839 36519 4851
rect 36575 5027 36633 5039
rect 36575 4851 36587 5027
rect 36621 4851 36633 5027
rect 36575 4839 36633 4851
rect 36833 5027 36891 5039
rect 36833 4851 36845 5027
rect 36879 4851 36891 5027
rect 36833 4839 36891 4851
rect 36947 5027 37005 5039
rect 36947 4851 36959 5027
rect 36993 4851 37005 5027
rect 36947 4839 37005 4851
rect 37205 5027 37263 5039
rect 37205 4851 37217 5027
rect 37251 4851 37263 5027
rect 37205 4839 37263 4851
rect 37319 5027 37377 5039
rect 37319 4851 37331 5027
rect 37365 4851 37377 5027
rect 37319 4839 37377 4851
rect 37577 5027 37635 5039
rect 37577 4851 37589 5027
rect 37623 4851 37635 5027
rect 37577 4839 37635 4851
rect 37691 5027 37749 5039
rect 37691 4851 37703 5027
rect 37737 4851 37749 5027
rect 37691 4839 37749 4851
rect 37949 5027 38007 5039
rect 37949 4851 37961 5027
rect 37995 4851 38007 5027
rect 37949 4839 38007 4851
rect 38063 5027 38121 5039
rect 38063 4851 38075 5027
rect 38109 4851 38121 5027
rect 38063 4839 38121 4851
rect 38321 5027 38379 5039
rect 38321 4851 38333 5027
rect 38367 4851 38379 5027
rect 38321 4839 38379 4851
rect 38435 5027 38493 5039
rect 38435 4851 38447 5027
rect 38481 4851 38493 5027
rect 38435 4839 38493 4851
rect 38693 5027 38751 5039
rect 38693 4851 38705 5027
rect 38739 4851 38751 5027
rect 38693 4839 38751 4851
rect 38807 5027 38865 5039
rect 38807 4851 38819 5027
rect 38853 4851 38865 5027
rect 38807 4839 38865 4851
rect 39065 5027 39123 5039
rect 39065 4851 39077 5027
rect 39111 4851 39123 5027
rect 39065 4839 39123 4851
rect 30251 4609 30309 4621
rect 30251 4433 30263 4609
rect 30297 4433 30309 4609
rect 30251 4421 30309 4433
rect 30509 4609 30567 4621
rect 30509 4433 30521 4609
rect 30555 4433 30567 4609
rect 30509 4421 30567 4433
rect 30623 4609 30681 4621
rect 30623 4433 30635 4609
rect 30669 4433 30681 4609
rect 30623 4421 30681 4433
rect 30881 4609 30939 4621
rect 30881 4433 30893 4609
rect 30927 4433 30939 4609
rect 30881 4421 30939 4433
rect 30995 4609 31053 4621
rect 30995 4433 31007 4609
rect 31041 4433 31053 4609
rect 30995 4421 31053 4433
rect 31253 4609 31311 4621
rect 31253 4433 31265 4609
rect 31299 4433 31311 4609
rect 31253 4421 31311 4433
rect 31367 4609 31425 4621
rect 31367 4433 31379 4609
rect 31413 4433 31425 4609
rect 31367 4421 31425 4433
rect 31625 4609 31683 4621
rect 31625 4433 31637 4609
rect 31671 4433 31683 4609
rect 31625 4421 31683 4433
rect 31739 4609 31797 4621
rect 31739 4433 31751 4609
rect 31785 4433 31797 4609
rect 31739 4421 31797 4433
rect 31997 4609 32055 4621
rect 31997 4433 32009 4609
rect 32043 4433 32055 4609
rect 31997 4421 32055 4433
rect 32111 4609 32169 4621
rect 32111 4433 32123 4609
rect 32157 4433 32169 4609
rect 32111 4421 32169 4433
rect 32369 4609 32427 4621
rect 32369 4433 32381 4609
rect 32415 4433 32427 4609
rect 32369 4421 32427 4433
rect 32483 4609 32541 4621
rect 32483 4433 32495 4609
rect 32529 4433 32541 4609
rect 32483 4421 32541 4433
rect 32741 4609 32799 4621
rect 32741 4433 32753 4609
rect 32787 4433 32799 4609
rect 32741 4421 32799 4433
rect 32855 4609 32913 4621
rect 32855 4433 32867 4609
rect 32901 4433 32913 4609
rect 32855 4421 32913 4433
rect 33113 4609 33171 4621
rect 33113 4433 33125 4609
rect 33159 4433 33171 4609
rect 33113 4421 33171 4433
rect 33227 4609 33285 4621
rect 33227 4433 33239 4609
rect 33273 4433 33285 4609
rect 33227 4421 33285 4433
rect 33485 4609 33543 4621
rect 33485 4433 33497 4609
rect 33531 4433 33543 4609
rect 33485 4421 33543 4433
rect 33599 4609 33657 4621
rect 33599 4433 33611 4609
rect 33645 4433 33657 4609
rect 33599 4421 33657 4433
rect 33857 4609 33915 4621
rect 33857 4433 33869 4609
rect 33903 4433 33915 4609
rect 33857 4421 33915 4433
rect 33971 4609 34029 4621
rect 33971 4433 33983 4609
rect 34017 4433 34029 4609
rect 33971 4421 34029 4433
rect 34229 4609 34287 4621
rect 34229 4433 34241 4609
rect 34275 4433 34287 4609
rect 34229 4421 34287 4433
rect 34343 4609 34401 4621
rect 34343 4433 34355 4609
rect 34389 4433 34401 4609
rect 34343 4421 34401 4433
rect 34601 4609 34659 4621
rect 34601 4433 34613 4609
rect 34647 4433 34659 4609
rect 34601 4421 34659 4433
rect 34715 4609 34773 4621
rect 34715 4433 34727 4609
rect 34761 4433 34773 4609
rect 34715 4421 34773 4433
rect 34973 4609 35031 4621
rect 34973 4433 34985 4609
rect 35019 4433 35031 4609
rect 34973 4421 35031 4433
rect 35087 4609 35145 4621
rect 35087 4433 35099 4609
rect 35133 4433 35145 4609
rect 35087 4421 35145 4433
rect 35345 4609 35403 4621
rect 35345 4433 35357 4609
rect 35391 4433 35403 4609
rect 35345 4421 35403 4433
rect 35459 4609 35517 4621
rect 35459 4433 35471 4609
rect 35505 4433 35517 4609
rect 35459 4421 35517 4433
rect 35717 4609 35775 4621
rect 35717 4433 35729 4609
rect 35763 4433 35775 4609
rect 35717 4421 35775 4433
rect 35831 4609 35889 4621
rect 35831 4433 35843 4609
rect 35877 4433 35889 4609
rect 35831 4421 35889 4433
rect 36089 4609 36147 4621
rect 36089 4433 36101 4609
rect 36135 4433 36147 4609
rect 36089 4421 36147 4433
rect 36203 4609 36261 4621
rect 36203 4433 36215 4609
rect 36249 4433 36261 4609
rect 36203 4421 36261 4433
rect 36461 4609 36519 4621
rect 36461 4433 36473 4609
rect 36507 4433 36519 4609
rect 36461 4421 36519 4433
rect 36575 4609 36633 4621
rect 36575 4433 36587 4609
rect 36621 4433 36633 4609
rect 36575 4421 36633 4433
rect 36833 4609 36891 4621
rect 36833 4433 36845 4609
rect 36879 4433 36891 4609
rect 36833 4421 36891 4433
rect 36947 4609 37005 4621
rect 36947 4433 36959 4609
rect 36993 4433 37005 4609
rect 36947 4421 37005 4433
rect 37205 4609 37263 4621
rect 37205 4433 37217 4609
rect 37251 4433 37263 4609
rect 37205 4421 37263 4433
rect 37319 4609 37377 4621
rect 37319 4433 37331 4609
rect 37365 4433 37377 4609
rect 37319 4421 37377 4433
rect 37577 4609 37635 4621
rect 37577 4433 37589 4609
rect 37623 4433 37635 4609
rect 37577 4421 37635 4433
rect 37691 4609 37749 4621
rect 37691 4433 37703 4609
rect 37737 4433 37749 4609
rect 37691 4421 37749 4433
rect 37949 4609 38007 4621
rect 37949 4433 37961 4609
rect 37995 4433 38007 4609
rect 37949 4421 38007 4433
rect 38063 4609 38121 4621
rect 38063 4433 38075 4609
rect 38109 4433 38121 4609
rect 38063 4421 38121 4433
rect 38321 4609 38379 4621
rect 38321 4433 38333 4609
rect 38367 4433 38379 4609
rect 38321 4421 38379 4433
rect 38435 4609 38493 4621
rect 38435 4433 38447 4609
rect 38481 4433 38493 4609
rect 38435 4421 38493 4433
rect 38693 4609 38751 4621
rect 38693 4433 38705 4609
rect 38739 4433 38751 4609
rect 38693 4421 38751 4433
rect 38807 4609 38865 4621
rect 38807 4433 38819 4609
rect 38853 4433 38865 4609
rect 38807 4421 38865 4433
rect 39065 4609 39123 4621
rect 39065 4433 39077 4609
rect 39111 4433 39123 4609
rect 39065 4421 39123 4433
rect 30251 4191 30309 4203
rect 30251 4015 30263 4191
rect 30297 4015 30309 4191
rect 30251 4003 30309 4015
rect 30509 4191 30567 4203
rect 30509 4015 30521 4191
rect 30555 4015 30567 4191
rect 30509 4003 30567 4015
rect 30623 4191 30681 4203
rect 30623 4015 30635 4191
rect 30669 4015 30681 4191
rect 30623 4003 30681 4015
rect 30881 4191 30939 4203
rect 30881 4015 30893 4191
rect 30927 4015 30939 4191
rect 30881 4003 30939 4015
rect 30995 4191 31053 4203
rect 30995 4015 31007 4191
rect 31041 4015 31053 4191
rect 30995 4003 31053 4015
rect 31253 4191 31311 4203
rect 31253 4015 31265 4191
rect 31299 4015 31311 4191
rect 31253 4003 31311 4015
rect 31367 4191 31425 4203
rect 31367 4015 31379 4191
rect 31413 4015 31425 4191
rect 31367 4003 31425 4015
rect 31625 4191 31683 4203
rect 31625 4015 31637 4191
rect 31671 4015 31683 4191
rect 31625 4003 31683 4015
rect 31739 4191 31797 4203
rect 31739 4015 31751 4191
rect 31785 4015 31797 4191
rect 31739 4003 31797 4015
rect 31997 4191 32055 4203
rect 31997 4015 32009 4191
rect 32043 4015 32055 4191
rect 31997 4003 32055 4015
rect 32111 4191 32169 4203
rect 32111 4015 32123 4191
rect 32157 4015 32169 4191
rect 32111 4003 32169 4015
rect 32369 4191 32427 4203
rect 32369 4015 32381 4191
rect 32415 4015 32427 4191
rect 32369 4003 32427 4015
rect 32483 4191 32541 4203
rect 32483 4015 32495 4191
rect 32529 4015 32541 4191
rect 32483 4003 32541 4015
rect 32741 4191 32799 4203
rect 32741 4015 32753 4191
rect 32787 4015 32799 4191
rect 32741 4003 32799 4015
rect 32855 4191 32913 4203
rect 32855 4015 32867 4191
rect 32901 4015 32913 4191
rect 32855 4003 32913 4015
rect 33113 4191 33171 4203
rect 33113 4015 33125 4191
rect 33159 4015 33171 4191
rect 33113 4003 33171 4015
rect 33227 4191 33285 4203
rect 33227 4015 33239 4191
rect 33273 4015 33285 4191
rect 33227 4003 33285 4015
rect 33485 4191 33543 4203
rect 33485 4015 33497 4191
rect 33531 4015 33543 4191
rect 33485 4003 33543 4015
rect 33599 4191 33657 4203
rect 33599 4015 33611 4191
rect 33645 4015 33657 4191
rect 33599 4003 33657 4015
rect 33857 4191 33915 4203
rect 33857 4015 33869 4191
rect 33903 4015 33915 4191
rect 33857 4003 33915 4015
rect 33971 4191 34029 4203
rect 33971 4015 33983 4191
rect 34017 4015 34029 4191
rect 33971 4003 34029 4015
rect 34229 4191 34287 4203
rect 34229 4015 34241 4191
rect 34275 4015 34287 4191
rect 34229 4003 34287 4015
rect 34343 4191 34401 4203
rect 34343 4015 34355 4191
rect 34389 4015 34401 4191
rect 34343 4003 34401 4015
rect 34601 4191 34659 4203
rect 34601 4015 34613 4191
rect 34647 4015 34659 4191
rect 34601 4003 34659 4015
rect 34715 4191 34773 4203
rect 34715 4015 34727 4191
rect 34761 4015 34773 4191
rect 34715 4003 34773 4015
rect 34973 4191 35031 4203
rect 34973 4015 34985 4191
rect 35019 4015 35031 4191
rect 34973 4003 35031 4015
rect 35087 4191 35145 4203
rect 35087 4015 35099 4191
rect 35133 4015 35145 4191
rect 35087 4003 35145 4015
rect 35345 4191 35403 4203
rect 35345 4015 35357 4191
rect 35391 4015 35403 4191
rect 35345 4003 35403 4015
rect 35459 4191 35517 4203
rect 35459 4015 35471 4191
rect 35505 4015 35517 4191
rect 35459 4003 35517 4015
rect 35717 4191 35775 4203
rect 35717 4015 35729 4191
rect 35763 4015 35775 4191
rect 35717 4003 35775 4015
rect 35831 4191 35889 4203
rect 35831 4015 35843 4191
rect 35877 4015 35889 4191
rect 35831 4003 35889 4015
rect 36089 4191 36147 4203
rect 36089 4015 36101 4191
rect 36135 4015 36147 4191
rect 36089 4003 36147 4015
rect 36203 4191 36261 4203
rect 36203 4015 36215 4191
rect 36249 4015 36261 4191
rect 36203 4003 36261 4015
rect 36461 4191 36519 4203
rect 36461 4015 36473 4191
rect 36507 4015 36519 4191
rect 36461 4003 36519 4015
rect 36575 4191 36633 4203
rect 36575 4015 36587 4191
rect 36621 4015 36633 4191
rect 36575 4003 36633 4015
rect 36833 4191 36891 4203
rect 36833 4015 36845 4191
rect 36879 4015 36891 4191
rect 36833 4003 36891 4015
rect 36947 4191 37005 4203
rect 36947 4015 36959 4191
rect 36993 4015 37005 4191
rect 36947 4003 37005 4015
rect 37205 4191 37263 4203
rect 37205 4015 37217 4191
rect 37251 4015 37263 4191
rect 37205 4003 37263 4015
rect 37319 4191 37377 4203
rect 37319 4015 37331 4191
rect 37365 4015 37377 4191
rect 37319 4003 37377 4015
rect 37577 4191 37635 4203
rect 37577 4015 37589 4191
rect 37623 4015 37635 4191
rect 37577 4003 37635 4015
rect 37691 4191 37749 4203
rect 37691 4015 37703 4191
rect 37737 4015 37749 4191
rect 37691 4003 37749 4015
rect 37949 4191 38007 4203
rect 37949 4015 37961 4191
rect 37995 4015 38007 4191
rect 37949 4003 38007 4015
rect 38063 4191 38121 4203
rect 38063 4015 38075 4191
rect 38109 4015 38121 4191
rect 38063 4003 38121 4015
rect 38321 4191 38379 4203
rect 38321 4015 38333 4191
rect 38367 4015 38379 4191
rect 38321 4003 38379 4015
rect 38435 4191 38493 4203
rect 38435 4015 38447 4191
rect 38481 4015 38493 4191
rect 38435 4003 38493 4015
rect 38693 4191 38751 4203
rect 38693 4015 38705 4191
rect 38739 4015 38751 4191
rect 38693 4003 38751 4015
rect 38807 4191 38865 4203
rect 38807 4015 38819 4191
rect 38853 4015 38865 4191
rect 38807 4003 38865 4015
rect 39065 4191 39123 4203
rect 39065 4015 39077 4191
rect 39111 4015 39123 4191
rect 39065 4003 39123 4015
rect 30251 3773 30309 3785
rect 30251 3597 30263 3773
rect 30297 3597 30309 3773
rect 30251 3585 30309 3597
rect 30509 3773 30567 3785
rect 30509 3597 30521 3773
rect 30555 3597 30567 3773
rect 30509 3585 30567 3597
rect 30623 3773 30681 3785
rect 30623 3597 30635 3773
rect 30669 3597 30681 3773
rect 30623 3585 30681 3597
rect 30881 3773 30939 3785
rect 30881 3597 30893 3773
rect 30927 3597 30939 3773
rect 30881 3585 30939 3597
rect 30995 3773 31053 3785
rect 30995 3597 31007 3773
rect 31041 3597 31053 3773
rect 30995 3585 31053 3597
rect 31253 3773 31311 3785
rect 31253 3597 31265 3773
rect 31299 3597 31311 3773
rect 31253 3585 31311 3597
rect 31367 3773 31425 3785
rect 31367 3597 31379 3773
rect 31413 3597 31425 3773
rect 31367 3585 31425 3597
rect 31625 3773 31683 3785
rect 31625 3597 31637 3773
rect 31671 3597 31683 3773
rect 31625 3585 31683 3597
rect 31739 3773 31797 3785
rect 31739 3597 31751 3773
rect 31785 3597 31797 3773
rect 31739 3585 31797 3597
rect 31997 3773 32055 3785
rect 31997 3597 32009 3773
rect 32043 3597 32055 3773
rect 31997 3585 32055 3597
rect 32111 3773 32169 3785
rect 32111 3597 32123 3773
rect 32157 3597 32169 3773
rect 32111 3585 32169 3597
rect 32369 3773 32427 3785
rect 32369 3597 32381 3773
rect 32415 3597 32427 3773
rect 32369 3585 32427 3597
rect 32483 3773 32541 3785
rect 32483 3597 32495 3773
rect 32529 3597 32541 3773
rect 32483 3585 32541 3597
rect 32741 3773 32799 3785
rect 32741 3597 32753 3773
rect 32787 3597 32799 3773
rect 32741 3585 32799 3597
rect 32855 3773 32913 3785
rect 32855 3597 32867 3773
rect 32901 3597 32913 3773
rect 32855 3585 32913 3597
rect 33113 3773 33171 3785
rect 33113 3597 33125 3773
rect 33159 3597 33171 3773
rect 33113 3585 33171 3597
rect 33227 3773 33285 3785
rect 33227 3597 33239 3773
rect 33273 3597 33285 3773
rect 33227 3585 33285 3597
rect 33485 3773 33543 3785
rect 33485 3597 33497 3773
rect 33531 3597 33543 3773
rect 33485 3585 33543 3597
rect 33599 3773 33657 3785
rect 33599 3597 33611 3773
rect 33645 3597 33657 3773
rect 33599 3585 33657 3597
rect 33857 3773 33915 3785
rect 33857 3597 33869 3773
rect 33903 3597 33915 3773
rect 33857 3585 33915 3597
rect 33971 3773 34029 3785
rect 33971 3597 33983 3773
rect 34017 3597 34029 3773
rect 33971 3585 34029 3597
rect 34229 3773 34287 3785
rect 34229 3597 34241 3773
rect 34275 3597 34287 3773
rect 34229 3585 34287 3597
rect 34343 3773 34401 3785
rect 34343 3597 34355 3773
rect 34389 3597 34401 3773
rect 34343 3585 34401 3597
rect 34601 3773 34659 3785
rect 34601 3597 34613 3773
rect 34647 3597 34659 3773
rect 34601 3585 34659 3597
rect 34715 3773 34773 3785
rect 34715 3597 34727 3773
rect 34761 3597 34773 3773
rect 34715 3585 34773 3597
rect 34973 3773 35031 3785
rect 34973 3597 34985 3773
rect 35019 3597 35031 3773
rect 34973 3585 35031 3597
rect 35087 3773 35145 3785
rect 35087 3597 35099 3773
rect 35133 3597 35145 3773
rect 35087 3585 35145 3597
rect 35345 3773 35403 3785
rect 35345 3597 35357 3773
rect 35391 3597 35403 3773
rect 35345 3585 35403 3597
rect 35459 3773 35517 3785
rect 35459 3597 35471 3773
rect 35505 3597 35517 3773
rect 35459 3585 35517 3597
rect 35717 3773 35775 3785
rect 35717 3597 35729 3773
rect 35763 3597 35775 3773
rect 35717 3585 35775 3597
rect 35831 3773 35889 3785
rect 35831 3597 35843 3773
rect 35877 3597 35889 3773
rect 35831 3585 35889 3597
rect 36089 3773 36147 3785
rect 36089 3597 36101 3773
rect 36135 3597 36147 3773
rect 36089 3585 36147 3597
rect 36203 3773 36261 3785
rect 36203 3597 36215 3773
rect 36249 3597 36261 3773
rect 36203 3585 36261 3597
rect 36461 3773 36519 3785
rect 36461 3597 36473 3773
rect 36507 3597 36519 3773
rect 36461 3585 36519 3597
rect 36575 3773 36633 3785
rect 36575 3597 36587 3773
rect 36621 3597 36633 3773
rect 36575 3585 36633 3597
rect 36833 3773 36891 3785
rect 36833 3597 36845 3773
rect 36879 3597 36891 3773
rect 36833 3585 36891 3597
rect 36947 3773 37005 3785
rect 36947 3597 36959 3773
rect 36993 3597 37005 3773
rect 36947 3585 37005 3597
rect 37205 3773 37263 3785
rect 37205 3597 37217 3773
rect 37251 3597 37263 3773
rect 37205 3585 37263 3597
rect 37319 3773 37377 3785
rect 37319 3597 37331 3773
rect 37365 3597 37377 3773
rect 37319 3585 37377 3597
rect 37577 3773 37635 3785
rect 37577 3597 37589 3773
rect 37623 3597 37635 3773
rect 37577 3585 37635 3597
rect 37691 3773 37749 3785
rect 37691 3597 37703 3773
rect 37737 3597 37749 3773
rect 37691 3585 37749 3597
rect 37949 3773 38007 3785
rect 37949 3597 37961 3773
rect 37995 3597 38007 3773
rect 37949 3585 38007 3597
rect 38063 3773 38121 3785
rect 38063 3597 38075 3773
rect 38109 3597 38121 3773
rect 38063 3585 38121 3597
rect 38321 3773 38379 3785
rect 38321 3597 38333 3773
rect 38367 3597 38379 3773
rect 38321 3585 38379 3597
rect 38435 3773 38493 3785
rect 38435 3597 38447 3773
rect 38481 3597 38493 3773
rect 38435 3585 38493 3597
rect 38693 3773 38751 3785
rect 38693 3597 38705 3773
rect 38739 3597 38751 3773
rect 38693 3585 38751 3597
rect 38807 3773 38865 3785
rect 38807 3597 38819 3773
rect 38853 3597 38865 3773
rect 38807 3585 38865 3597
rect 39065 3773 39123 3785
rect 39065 3597 39077 3773
rect 39111 3597 39123 3773
rect 39065 3585 39123 3597
<< pdiff >>
rect 28763 12100 28821 12112
rect 28763 11724 28775 12100
rect 28809 11724 28821 12100
rect 28763 11712 28821 11724
rect 29021 12100 29079 12112
rect 29021 11724 29033 12100
rect 29067 11724 29079 12100
rect 29021 11712 29079 11724
rect 29135 12100 29193 12112
rect 29135 11724 29147 12100
rect 29181 11724 29193 12100
rect 29135 11712 29193 11724
rect 29393 12100 29451 12112
rect 29393 11724 29405 12100
rect 29439 11724 29451 12100
rect 29393 11712 29451 11724
rect 29507 12100 29565 12112
rect 29507 11724 29519 12100
rect 29553 11724 29565 12100
rect 29507 11712 29565 11724
rect 29765 12100 29823 12112
rect 29765 11724 29777 12100
rect 29811 11724 29823 12100
rect 29765 11712 29823 11724
rect 29879 12100 29937 12112
rect 29879 11724 29891 12100
rect 29925 11724 29937 12100
rect 29879 11712 29937 11724
rect 30137 12100 30195 12112
rect 30137 11724 30149 12100
rect 30183 11724 30195 12100
rect 30137 11712 30195 11724
rect 30251 12100 30309 12112
rect 30251 11724 30263 12100
rect 30297 11724 30309 12100
rect 30251 11712 30309 11724
rect 30509 12100 30567 12112
rect 30509 11724 30521 12100
rect 30555 11724 30567 12100
rect 30509 11712 30567 11724
rect 30623 12100 30681 12112
rect 30623 11724 30635 12100
rect 30669 11724 30681 12100
rect 30623 11712 30681 11724
rect 30881 12100 30939 12112
rect 30881 11724 30893 12100
rect 30927 11724 30939 12100
rect 30881 11712 30939 11724
rect 30995 12100 31053 12112
rect 30995 11724 31007 12100
rect 31041 11724 31053 12100
rect 30995 11712 31053 11724
rect 31253 12100 31311 12112
rect 31253 11724 31265 12100
rect 31299 11724 31311 12100
rect 31253 11712 31311 11724
rect 31367 12100 31425 12112
rect 31367 11724 31379 12100
rect 31413 11724 31425 12100
rect 31367 11712 31425 11724
rect 31625 12100 31683 12112
rect 31625 11724 31637 12100
rect 31671 11724 31683 12100
rect 31625 11712 31683 11724
rect 31739 12100 31797 12112
rect 31739 11724 31751 12100
rect 31785 11724 31797 12100
rect 31739 11712 31797 11724
rect 31997 12100 32055 12112
rect 31997 11724 32009 12100
rect 32043 11724 32055 12100
rect 31997 11712 32055 11724
rect 32111 12100 32169 12112
rect 32111 11724 32123 12100
rect 32157 11724 32169 12100
rect 32111 11712 32169 11724
rect 32369 12100 32427 12112
rect 32369 11724 32381 12100
rect 32415 11724 32427 12100
rect 32369 11712 32427 11724
rect 32483 12100 32541 12112
rect 32483 11724 32495 12100
rect 32529 11724 32541 12100
rect 32483 11712 32541 11724
rect 32741 12100 32799 12112
rect 32741 11724 32753 12100
rect 32787 11724 32799 12100
rect 32741 11712 32799 11724
rect 32855 12100 32913 12112
rect 32855 11724 32867 12100
rect 32901 11724 32913 12100
rect 32855 11712 32913 11724
rect 33113 12100 33171 12112
rect 33113 11724 33125 12100
rect 33159 11724 33171 12100
rect 33113 11712 33171 11724
rect 33227 12100 33285 12112
rect 33227 11724 33239 12100
rect 33273 11724 33285 12100
rect 33227 11712 33285 11724
rect 33485 12100 33543 12112
rect 33485 11724 33497 12100
rect 33531 11724 33543 12100
rect 33485 11712 33543 11724
rect 33599 12100 33657 12112
rect 33599 11724 33611 12100
rect 33645 11724 33657 12100
rect 33599 11712 33657 11724
rect 33857 12100 33915 12112
rect 33857 11724 33869 12100
rect 33903 11724 33915 12100
rect 33857 11712 33915 11724
rect 33971 12100 34029 12112
rect 33971 11724 33983 12100
rect 34017 11724 34029 12100
rect 33971 11712 34029 11724
rect 34229 12100 34287 12112
rect 34229 11724 34241 12100
rect 34275 11724 34287 12100
rect 34229 11712 34287 11724
rect 34343 12100 34401 12112
rect 34343 11724 34355 12100
rect 34389 11724 34401 12100
rect 34343 11712 34401 11724
rect 34601 12100 34659 12112
rect 34601 11724 34613 12100
rect 34647 11724 34659 12100
rect 34601 11712 34659 11724
rect 34715 12100 34773 12112
rect 34715 11724 34727 12100
rect 34761 11724 34773 12100
rect 34715 11712 34773 11724
rect 34973 12100 35031 12112
rect 34973 11724 34985 12100
rect 35019 11724 35031 12100
rect 34973 11712 35031 11724
rect 35087 12100 35145 12112
rect 35087 11724 35099 12100
rect 35133 11724 35145 12100
rect 35087 11712 35145 11724
rect 35345 12100 35403 12112
rect 35345 11724 35357 12100
rect 35391 11724 35403 12100
rect 35345 11712 35403 11724
rect 35459 12100 35517 12112
rect 35459 11724 35471 12100
rect 35505 11724 35517 12100
rect 35459 11712 35517 11724
rect 35717 12100 35775 12112
rect 35717 11724 35729 12100
rect 35763 11724 35775 12100
rect 35717 11712 35775 11724
rect 35831 12100 35889 12112
rect 35831 11724 35843 12100
rect 35877 11724 35889 12100
rect 35831 11712 35889 11724
rect 36089 12100 36147 12112
rect 36089 11724 36101 12100
rect 36135 11724 36147 12100
rect 36089 11712 36147 11724
rect 36203 12100 36261 12112
rect 36203 11724 36215 12100
rect 36249 11724 36261 12100
rect 36203 11712 36261 11724
rect 36461 12100 36519 12112
rect 36461 11724 36473 12100
rect 36507 11724 36519 12100
rect 36461 11712 36519 11724
rect 36575 12100 36633 12112
rect 36575 11724 36587 12100
rect 36621 11724 36633 12100
rect 36575 11712 36633 11724
rect 36833 12100 36891 12112
rect 36833 11724 36845 12100
rect 36879 11724 36891 12100
rect 36833 11712 36891 11724
rect 36947 12100 37005 12112
rect 36947 11724 36959 12100
rect 36993 11724 37005 12100
rect 36947 11712 37005 11724
rect 37205 12100 37263 12112
rect 37205 11724 37217 12100
rect 37251 11724 37263 12100
rect 37205 11712 37263 11724
rect 37319 12100 37377 12112
rect 37319 11724 37331 12100
rect 37365 11724 37377 12100
rect 37319 11712 37377 11724
rect 37577 12100 37635 12112
rect 37577 11724 37589 12100
rect 37623 11724 37635 12100
rect 37577 11712 37635 11724
rect 37691 12100 37749 12112
rect 37691 11724 37703 12100
rect 37737 11724 37749 12100
rect 37691 11712 37749 11724
rect 37949 12100 38007 12112
rect 37949 11724 37961 12100
rect 37995 11724 38007 12100
rect 37949 11712 38007 11724
rect 38063 12100 38121 12112
rect 38063 11724 38075 12100
rect 38109 11724 38121 12100
rect 38063 11712 38121 11724
rect 38321 12100 38379 12112
rect 38321 11724 38333 12100
rect 38367 11724 38379 12100
rect 38321 11712 38379 11724
rect 38435 12100 38493 12112
rect 38435 11724 38447 12100
rect 38481 11724 38493 12100
rect 38435 11712 38493 11724
rect 38693 12100 38751 12112
rect 38693 11724 38705 12100
rect 38739 11724 38751 12100
rect 38693 11712 38751 11724
rect 38807 12100 38865 12112
rect 38807 11724 38819 12100
rect 38853 11724 38865 12100
rect 38807 11712 38865 11724
rect 39065 12100 39123 12112
rect 39065 11724 39077 12100
rect 39111 11724 39123 12100
rect 39065 11712 39123 11724
rect 39179 12100 39237 12112
rect 39179 11724 39191 12100
rect 39225 11724 39237 12100
rect 39179 11712 39237 11724
rect 39437 12100 39495 12112
rect 39437 11724 39449 12100
rect 39483 11724 39495 12100
rect 39437 11712 39495 11724
rect 39551 12100 39609 12112
rect 39551 11724 39563 12100
rect 39597 11724 39609 12100
rect 39551 11712 39609 11724
rect 39809 12100 39867 12112
rect 39809 11724 39821 12100
rect 39855 11724 39867 12100
rect 39809 11712 39867 11724
rect 39923 12100 39981 12112
rect 39923 11724 39935 12100
rect 39969 11724 39981 12100
rect 39923 11712 39981 11724
rect 40181 12100 40239 12112
rect 40181 11724 40193 12100
rect 40227 11724 40239 12100
rect 40181 11712 40239 11724
rect 40295 12100 40353 12112
rect 40295 11724 40307 12100
rect 40341 11724 40353 12100
rect 40295 11712 40353 11724
rect 40553 12100 40611 12112
rect 40553 11724 40565 12100
rect 40599 11724 40611 12100
rect 40553 11712 40611 11724
rect 28763 11464 28821 11476
rect 28763 11088 28775 11464
rect 28809 11088 28821 11464
rect 28763 11076 28821 11088
rect 29021 11464 29079 11476
rect 29021 11088 29033 11464
rect 29067 11088 29079 11464
rect 29021 11076 29079 11088
rect 29135 11464 29193 11476
rect 29135 11088 29147 11464
rect 29181 11088 29193 11464
rect 29135 11076 29193 11088
rect 29393 11464 29451 11476
rect 29393 11088 29405 11464
rect 29439 11088 29451 11464
rect 29393 11076 29451 11088
rect 29507 11464 29565 11476
rect 29507 11088 29519 11464
rect 29553 11088 29565 11464
rect 29507 11076 29565 11088
rect 29765 11464 29823 11476
rect 29765 11088 29777 11464
rect 29811 11088 29823 11464
rect 29765 11076 29823 11088
rect 29879 11464 29937 11476
rect 29879 11088 29891 11464
rect 29925 11088 29937 11464
rect 29879 11076 29937 11088
rect 30137 11464 30195 11476
rect 30137 11088 30149 11464
rect 30183 11088 30195 11464
rect 30137 11076 30195 11088
rect 30251 11464 30309 11476
rect 30251 11088 30263 11464
rect 30297 11088 30309 11464
rect 30251 11076 30309 11088
rect 30509 11464 30567 11476
rect 30509 11088 30521 11464
rect 30555 11088 30567 11464
rect 30509 11076 30567 11088
rect 30623 11464 30681 11476
rect 30623 11088 30635 11464
rect 30669 11088 30681 11464
rect 30623 11076 30681 11088
rect 30881 11464 30939 11476
rect 30881 11088 30893 11464
rect 30927 11088 30939 11464
rect 30881 11076 30939 11088
rect 30995 11464 31053 11476
rect 30995 11088 31007 11464
rect 31041 11088 31053 11464
rect 30995 11076 31053 11088
rect 31253 11464 31311 11476
rect 31253 11088 31265 11464
rect 31299 11088 31311 11464
rect 31253 11076 31311 11088
rect 31367 11464 31425 11476
rect 31367 11088 31379 11464
rect 31413 11088 31425 11464
rect 31367 11076 31425 11088
rect 31625 11464 31683 11476
rect 31625 11088 31637 11464
rect 31671 11088 31683 11464
rect 31625 11076 31683 11088
rect 31739 11464 31797 11476
rect 31739 11088 31751 11464
rect 31785 11088 31797 11464
rect 31739 11076 31797 11088
rect 31997 11464 32055 11476
rect 31997 11088 32009 11464
rect 32043 11088 32055 11464
rect 31997 11076 32055 11088
rect 32111 11464 32169 11476
rect 32111 11088 32123 11464
rect 32157 11088 32169 11464
rect 32111 11076 32169 11088
rect 32369 11464 32427 11476
rect 32369 11088 32381 11464
rect 32415 11088 32427 11464
rect 32369 11076 32427 11088
rect 32483 11464 32541 11476
rect 32483 11088 32495 11464
rect 32529 11088 32541 11464
rect 32483 11076 32541 11088
rect 32741 11464 32799 11476
rect 32741 11088 32753 11464
rect 32787 11088 32799 11464
rect 32741 11076 32799 11088
rect 32855 11464 32913 11476
rect 32855 11088 32867 11464
rect 32901 11088 32913 11464
rect 32855 11076 32913 11088
rect 33113 11464 33171 11476
rect 33113 11088 33125 11464
rect 33159 11088 33171 11464
rect 33113 11076 33171 11088
rect 33227 11464 33285 11476
rect 33227 11088 33239 11464
rect 33273 11088 33285 11464
rect 33227 11076 33285 11088
rect 33485 11464 33543 11476
rect 33485 11088 33497 11464
rect 33531 11088 33543 11464
rect 33485 11076 33543 11088
rect 33599 11464 33657 11476
rect 33599 11088 33611 11464
rect 33645 11088 33657 11464
rect 33599 11076 33657 11088
rect 33857 11464 33915 11476
rect 33857 11088 33869 11464
rect 33903 11088 33915 11464
rect 33857 11076 33915 11088
rect 33971 11464 34029 11476
rect 33971 11088 33983 11464
rect 34017 11088 34029 11464
rect 33971 11076 34029 11088
rect 34229 11464 34287 11476
rect 34229 11088 34241 11464
rect 34275 11088 34287 11464
rect 34229 11076 34287 11088
rect 34343 11464 34401 11476
rect 34343 11088 34355 11464
rect 34389 11088 34401 11464
rect 34343 11076 34401 11088
rect 34601 11464 34659 11476
rect 34601 11088 34613 11464
rect 34647 11088 34659 11464
rect 34601 11076 34659 11088
rect 34715 11464 34773 11476
rect 34715 11088 34727 11464
rect 34761 11088 34773 11464
rect 34715 11076 34773 11088
rect 34973 11464 35031 11476
rect 34973 11088 34985 11464
rect 35019 11088 35031 11464
rect 34973 11076 35031 11088
rect 35087 11464 35145 11476
rect 35087 11088 35099 11464
rect 35133 11088 35145 11464
rect 35087 11076 35145 11088
rect 35345 11464 35403 11476
rect 35345 11088 35357 11464
rect 35391 11088 35403 11464
rect 35345 11076 35403 11088
rect 35459 11464 35517 11476
rect 35459 11088 35471 11464
rect 35505 11088 35517 11464
rect 35459 11076 35517 11088
rect 35717 11464 35775 11476
rect 35717 11088 35729 11464
rect 35763 11088 35775 11464
rect 35717 11076 35775 11088
rect 35831 11464 35889 11476
rect 35831 11088 35843 11464
rect 35877 11088 35889 11464
rect 35831 11076 35889 11088
rect 36089 11464 36147 11476
rect 36089 11088 36101 11464
rect 36135 11088 36147 11464
rect 36089 11076 36147 11088
rect 36203 11464 36261 11476
rect 36203 11088 36215 11464
rect 36249 11088 36261 11464
rect 36203 11076 36261 11088
rect 36461 11464 36519 11476
rect 36461 11088 36473 11464
rect 36507 11088 36519 11464
rect 36461 11076 36519 11088
rect 36575 11464 36633 11476
rect 36575 11088 36587 11464
rect 36621 11088 36633 11464
rect 36575 11076 36633 11088
rect 36833 11464 36891 11476
rect 36833 11088 36845 11464
rect 36879 11088 36891 11464
rect 36833 11076 36891 11088
rect 36947 11464 37005 11476
rect 36947 11088 36959 11464
rect 36993 11088 37005 11464
rect 36947 11076 37005 11088
rect 37205 11464 37263 11476
rect 37205 11088 37217 11464
rect 37251 11088 37263 11464
rect 37205 11076 37263 11088
rect 37319 11464 37377 11476
rect 37319 11088 37331 11464
rect 37365 11088 37377 11464
rect 37319 11076 37377 11088
rect 37577 11464 37635 11476
rect 37577 11088 37589 11464
rect 37623 11088 37635 11464
rect 37577 11076 37635 11088
rect 37691 11464 37749 11476
rect 37691 11088 37703 11464
rect 37737 11088 37749 11464
rect 37691 11076 37749 11088
rect 37949 11464 38007 11476
rect 37949 11088 37961 11464
rect 37995 11088 38007 11464
rect 37949 11076 38007 11088
rect 38063 11464 38121 11476
rect 38063 11088 38075 11464
rect 38109 11088 38121 11464
rect 38063 11076 38121 11088
rect 38321 11464 38379 11476
rect 38321 11088 38333 11464
rect 38367 11088 38379 11464
rect 38321 11076 38379 11088
rect 38435 11464 38493 11476
rect 38435 11088 38447 11464
rect 38481 11088 38493 11464
rect 38435 11076 38493 11088
rect 38693 11464 38751 11476
rect 38693 11088 38705 11464
rect 38739 11088 38751 11464
rect 38693 11076 38751 11088
rect 38807 11464 38865 11476
rect 38807 11088 38819 11464
rect 38853 11088 38865 11464
rect 38807 11076 38865 11088
rect 39065 11464 39123 11476
rect 39065 11088 39077 11464
rect 39111 11088 39123 11464
rect 39065 11076 39123 11088
rect 39179 11464 39237 11476
rect 39179 11088 39191 11464
rect 39225 11088 39237 11464
rect 39179 11076 39237 11088
rect 39437 11464 39495 11476
rect 39437 11088 39449 11464
rect 39483 11088 39495 11464
rect 39437 11076 39495 11088
rect 39551 11464 39609 11476
rect 39551 11088 39563 11464
rect 39597 11088 39609 11464
rect 39551 11076 39609 11088
rect 39809 11464 39867 11476
rect 39809 11088 39821 11464
rect 39855 11088 39867 11464
rect 39809 11076 39867 11088
rect 39923 11464 39981 11476
rect 39923 11088 39935 11464
rect 39969 11088 39981 11464
rect 39923 11076 39981 11088
rect 40181 11464 40239 11476
rect 40181 11088 40193 11464
rect 40227 11088 40239 11464
rect 40181 11076 40239 11088
rect 40295 11464 40353 11476
rect 40295 11088 40307 11464
rect 40341 11088 40353 11464
rect 40295 11076 40353 11088
rect 40553 11464 40611 11476
rect 40553 11088 40565 11464
rect 40599 11088 40611 11464
rect 40553 11076 40611 11088
rect 28763 10828 28821 10840
rect 28763 10452 28775 10828
rect 28809 10452 28821 10828
rect 28763 10440 28821 10452
rect 29021 10828 29079 10840
rect 29021 10452 29033 10828
rect 29067 10452 29079 10828
rect 29021 10440 29079 10452
rect 29135 10828 29193 10840
rect 29135 10452 29147 10828
rect 29181 10452 29193 10828
rect 29135 10440 29193 10452
rect 29393 10828 29451 10840
rect 29393 10452 29405 10828
rect 29439 10452 29451 10828
rect 29393 10440 29451 10452
rect 29507 10828 29565 10840
rect 29507 10452 29519 10828
rect 29553 10452 29565 10828
rect 29507 10440 29565 10452
rect 29765 10828 29823 10840
rect 29765 10452 29777 10828
rect 29811 10452 29823 10828
rect 29765 10440 29823 10452
rect 29879 10828 29937 10840
rect 29879 10452 29891 10828
rect 29925 10452 29937 10828
rect 29879 10440 29937 10452
rect 30137 10828 30195 10840
rect 30137 10452 30149 10828
rect 30183 10452 30195 10828
rect 30137 10440 30195 10452
rect 30251 10828 30309 10840
rect 30251 10452 30263 10828
rect 30297 10452 30309 10828
rect 30251 10440 30309 10452
rect 30509 10828 30567 10840
rect 30509 10452 30521 10828
rect 30555 10452 30567 10828
rect 30509 10440 30567 10452
rect 30623 10828 30681 10840
rect 30623 10452 30635 10828
rect 30669 10452 30681 10828
rect 30623 10440 30681 10452
rect 30881 10828 30939 10840
rect 30881 10452 30893 10828
rect 30927 10452 30939 10828
rect 30881 10440 30939 10452
rect 30995 10828 31053 10840
rect 30995 10452 31007 10828
rect 31041 10452 31053 10828
rect 30995 10440 31053 10452
rect 31253 10828 31311 10840
rect 31253 10452 31265 10828
rect 31299 10452 31311 10828
rect 31253 10440 31311 10452
rect 31367 10828 31425 10840
rect 31367 10452 31379 10828
rect 31413 10452 31425 10828
rect 31367 10440 31425 10452
rect 31625 10828 31683 10840
rect 31625 10452 31637 10828
rect 31671 10452 31683 10828
rect 31625 10440 31683 10452
rect 31739 10828 31797 10840
rect 31739 10452 31751 10828
rect 31785 10452 31797 10828
rect 31739 10440 31797 10452
rect 31997 10828 32055 10840
rect 31997 10452 32009 10828
rect 32043 10452 32055 10828
rect 31997 10440 32055 10452
rect 32111 10828 32169 10840
rect 32111 10452 32123 10828
rect 32157 10452 32169 10828
rect 32111 10440 32169 10452
rect 32369 10828 32427 10840
rect 32369 10452 32381 10828
rect 32415 10452 32427 10828
rect 32369 10440 32427 10452
rect 32483 10828 32541 10840
rect 32483 10452 32495 10828
rect 32529 10452 32541 10828
rect 32483 10440 32541 10452
rect 32741 10828 32799 10840
rect 32741 10452 32753 10828
rect 32787 10452 32799 10828
rect 32741 10440 32799 10452
rect 32855 10828 32913 10840
rect 32855 10452 32867 10828
rect 32901 10452 32913 10828
rect 32855 10440 32913 10452
rect 33113 10828 33171 10840
rect 33113 10452 33125 10828
rect 33159 10452 33171 10828
rect 33113 10440 33171 10452
rect 33227 10828 33285 10840
rect 33227 10452 33239 10828
rect 33273 10452 33285 10828
rect 33227 10440 33285 10452
rect 33485 10828 33543 10840
rect 33485 10452 33497 10828
rect 33531 10452 33543 10828
rect 33485 10440 33543 10452
rect 33599 10828 33657 10840
rect 33599 10452 33611 10828
rect 33645 10452 33657 10828
rect 33599 10440 33657 10452
rect 33857 10828 33915 10840
rect 33857 10452 33869 10828
rect 33903 10452 33915 10828
rect 33857 10440 33915 10452
rect 33971 10828 34029 10840
rect 33971 10452 33983 10828
rect 34017 10452 34029 10828
rect 33971 10440 34029 10452
rect 34229 10828 34287 10840
rect 34229 10452 34241 10828
rect 34275 10452 34287 10828
rect 34229 10440 34287 10452
rect 34343 10828 34401 10840
rect 34343 10452 34355 10828
rect 34389 10452 34401 10828
rect 34343 10440 34401 10452
rect 34601 10828 34659 10840
rect 34601 10452 34613 10828
rect 34647 10452 34659 10828
rect 34601 10440 34659 10452
rect 34715 10828 34773 10840
rect 34715 10452 34727 10828
rect 34761 10452 34773 10828
rect 34715 10440 34773 10452
rect 34973 10828 35031 10840
rect 34973 10452 34985 10828
rect 35019 10452 35031 10828
rect 34973 10440 35031 10452
rect 35087 10828 35145 10840
rect 35087 10452 35099 10828
rect 35133 10452 35145 10828
rect 35087 10440 35145 10452
rect 35345 10828 35403 10840
rect 35345 10452 35357 10828
rect 35391 10452 35403 10828
rect 35345 10440 35403 10452
rect 35459 10828 35517 10840
rect 35459 10452 35471 10828
rect 35505 10452 35517 10828
rect 35459 10440 35517 10452
rect 35717 10828 35775 10840
rect 35717 10452 35729 10828
rect 35763 10452 35775 10828
rect 35717 10440 35775 10452
rect 35831 10828 35889 10840
rect 35831 10452 35843 10828
rect 35877 10452 35889 10828
rect 35831 10440 35889 10452
rect 36089 10828 36147 10840
rect 36089 10452 36101 10828
rect 36135 10452 36147 10828
rect 36089 10440 36147 10452
rect 36203 10828 36261 10840
rect 36203 10452 36215 10828
rect 36249 10452 36261 10828
rect 36203 10440 36261 10452
rect 36461 10828 36519 10840
rect 36461 10452 36473 10828
rect 36507 10452 36519 10828
rect 36461 10440 36519 10452
rect 36575 10828 36633 10840
rect 36575 10452 36587 10828
rect 36621 10452 36633 10828
rect 36575 10440 36633 10452
rect 36833 10828 36891 10840
rect 36833 10452 36845 10828
rect 36879 10452 36891 10828
rect 36833 10440 36891 10452
rect 36947 10828 37005 10840
rect 36947 10452 36959 10828
rect 36993 10452 37005 10828
rect 36947 10440 37005 10452
rect 37205 10828 37263 10840
rect 37205 10452 37217 10828
rect 37251 10452 37263 10828
rect 37205 10440 37263 10452
rect 37319 10828 37377 10840
rect 37319 10452 37331 10828
rect 37365 10452 37377 10828
rect 37319 10440 37377 10452
rect 37577 10828 37635 10840
rect 37577 10452 37589 10828
rect 37623 10452 37635 10828
rect 37577 10440 37635 10452
rect 37691 10828 37749 10840
rect 37691 10452 37703 10828
rect 37737 10452 37749 10828
rect 37691 10440 37749 10452
rect 37949 10828 38007 10840
rect 37949 10452 37961 10828
rect 37995 10452 38007 10828
rect 37949 10440 38007 10452
rect 38063 10828 38121 10840
rect 38063 10452 38075 10828
rect 38109 10452 38121 10828
rect 38063 10440 38121 10452
rect 38321 10828 38379 10840
rect 38321 10452 38333 10828
rect 38367 10452 38379 10828
rect 38321 10440 38379 10452
rect 38435 10828 38493 10840
rect 38435 10452 38447 10828
rect 38481 10452 38493 10828
rect 38435 10440 38493 10452
rect 38693 10828 38751 10840
rect 38693 10452 38705 10828
rect 38739 10452 38751 10828
rect 38693 10440 38751 10452
rect 38807 10828 38865 10840
rect 38807 10452 38819 10828
rect 38853 10452 38865 10828
rect 38807 10440 38865 10452
rect 39065 10828 39123 10840
rect 39065 10452 39077 10828
rect 39111 10452 39123 10828
rect 39065 10440 39123 10452
rect 39179 10828 39237 10840
rect 39179 10452 39191 10828
rect 39225 10452 39237 10828
rect 39179 10440 39237 10452
rect 39437 10828 39495 10840
rect 39437 10452 39449 10828
rect 39483 10452 39495 10828
rect 39437 10440 39495 10452
rect 39551 10828 39609 10840
rect 39551 10452 39563 10828
rect 39597 10452 39609 10828
rect 39551 10440 39609 10452
rect 39809 10828 39867 10840
rect 39809 10452 39821 10828
rect 39855 10452 39867 10828
rect 39809 10440 39867 10452
rect 39923 10828 39981 10840
rect 39923 10452 39935 10828
rect 39969 10452 39981 10828
rect 39923 10440 39981 10452
rect 40181 10828 40239 10840
rect 40181 10452 40193 10828
rect 40227 10452 40239 10828
rect 40181 10440 40239 10452
rect 40295 10828 40353 10840
rect 40295 10452 40307 10828
rect 40341 10452 40353 10828
rect 40295 10440 40353 10452
rect 40553 10828 40611 10840
rect 40553 10452 40565 10828
rect 40599 10452 40611 10828
rect 40553 10440 40611 10452
rect 30251 9712 30309 9724
rect 30251 8936 30263 9712
rect 30297 8936 30309 9712
rect 30251 8924 30309 8936
rect 30509 9712 30567 9724
rect 30509 8936 30521 9712
rect 30555 8936 30567 9712
rect 30509 8924 30567 8936
rect 30623 9712 30681 9724
rect 30623 8936 30635 9712
rect 30669 8936 30681 9712
rect 30623 8924 30681 8936
rect 30881 9712 30939 9724
rect 30881 8936 30893 9712
rect 30927 8936 30939 9712
rect 30881 8924 30939 8936
rect 30995 9712 31053 9724
rect 30995 8936 31007 9712
rect 31041 8936 31053 9712
rect 30995 8924 31053 8936
rect 31253 9712 31311 9724
rect 31253 8936 31265 9712
rect 31299 8936 31311 9712
rect 31253 8924 31311 8936
rect 31367 9712 31425 9724
rect 31367 8936 31379 9712
rect 31413 8936 31425 9712
rect 31367 8924 31425 8936
rect 31625 9712 31683 9724
rect 31625 8936 31637 9712
rect 31671 8936 31683 9712
rect 31625 8924 31683 8936
rect 31739 9712 31797 9724
rect 31739 8936 31751 9712
rect 31785 8936 31797 9712
rect 31739 8924 31797 8936
rect 31997 9712 32055 9724
rect 31997 8936 32009 9712
rect 32043 8936 32055 9712
rect 31997 8924 32055 8936
rect 32111 9712 32169 9724
rect 32111 8936 32123 9712
rect 32157 8936 32169 9712
rect 32111 8924 32169 8936
rect 32369 9712 32427 9724
rect 32369 8936 32381 9712
rect 32415 8936 32427 9712
rect 32369 8924 32427 8936
rect 32483 9712 32541 9724
rect 32483 8936 32495 9712
rect 32529 8936 32541 9712
rect 32483 8924 32541 8936
rect 32741 9712 32799 9724
rect 32741 8936 32753 9712
rect 32787 8936 32799 9712
rect 32741 8924 32799 8936
rect 32855 9712 32913 9724
rect 32855 8936 32867 9712
rect 32901 8936 32913 9712
rect 32855 8924 32913 8936
rect 33113 9712 33171 9724
rect 33113 8936 33125 9712
rect 33159 8936 33171 9712
rect 33113 8924 33171 8936
rect 30251 8676 30309 8688
rect 30251 7900 30263 8676
rect 30297 7900 30309 8676
rect 30251 7888 30309 7900
rect 30509 8676 30567 8688
rect 30509 7900 30521 8676
rect 30555 7900 30567 8676
rect 30509 7888 30567 7900
rect 30623 8676 30681 8688
rect 30623 7900 30635 8676
rect 30669 7900 30681 8676
rect 30623 7888 30681 7900
rect 30881 8676 30939 8688
rect 30881 7900 30893 8676
rect 30927 7900 30939 8676
rect 30881 7888 30939 7900
rect 30995 8676 31053 8688
rect 30995 7900 31007 8676
rect 31041 7900 31053 8676
rect 30995 7888 31053 7900
rect 31253 8676 31311 8688
rect 31253 7900 31265 8676
rect 31299 7900 31311 8676
rect 31253 7888 31311 7900
rect 31367 8676 31425 8688
rect 31367 7900 31379 8676
rect 31413 7900 31425 8676
rect 31367 7888 31425 7900
rect 31625 8676 31683 8688
rect 31625 7900 31637 8676
rect 31671 7900 31683 8676
rect 31625 7888 31683 7900
rect 31739 8676 31797 8688
rect 31739 7900 31751 8676
rect 31785 7900 31797 8676
rect 31739 7888 31797 7900
rect 31997 8676 32055 8688
rect 31997 7900 32009 8676
rect 32043 7900 32055 8676
rect 31997 7888 32055 7900
rect 32111 8676 32169 8688
rect 32111 7900 32123 8676
rect 32157 7900 32169 8676
rect 32111 7888 32169 7900
rect 32369 8676 32427 8688
rect 32369 7900 32381 8676
rect 32415 7900 32427 8676
rect 32369 7888 32427 7900
rect 32483 8676 32541 8688
rect 32483 7900 32495 8676
rect 32529 7900 32541 8676
rect 32483 7888 32541 7900
rect 32741 8676 32799 8688
rect 32741 7900 32753 8676
rect 32787 7900 32799 8676
rect 32741 7888 32799 7900
rect 32855 8676 32913 8688
rect 32855 7900 32867 8676
rect 32901 7900 32913 8676
rect 32855 7888 32913 7900
rect 33113 8676 33171 8688
rect 33113 7900 33125 8676
rect 33159 7900 33171 8676
rect 33113 7888 33171 7900
rect 30251 7640 30309 7652
rect 30251 6864 30263 7640
rect 30297 6864 30309 7640
rect 30251 6852 30309 6864
rect 30509 7640 30567 7652
rect 30509 6864 30521 7640
rect 30555 6864 30567 7640
rect 30509 6852 30567 6864
rect 30623 7640 30681 7652
rect 30623 6864 30635 7640
rect 30669 6864 30681 7640
rect 30623 6852 30681 6864
rect 30881 7640 30939 7652
rect 30881 6864 30893 7640
rect 30927 6864 30939 7640
rect 30881 6852 30939 6864
rect 30995 7640 31053 7652
rect 30995 6864 31007 7640
rect 31041 6864 31053 7640
rect 30995 6852 31053 6864
rect 31253 7640 31311 7652
rect 31253 6864 31265 7640
rect 31299 6864 31311 7640
rect 31253 6852 31311 6864
rect 31367 7640 31425 7652
rect 31367 6864 31379 7640
rect 31413 6864 31425 7640
rect 31367 6852 31425 6864
rect 31625 7640 31683 7652
rect 31625 6864 31637 7640
rect 31671 6864 31683 7640
rect 31625 6852 31683 6864
rect 31739 7640 31797 7652
rect 31739 6864 31751 7640
rect 31785 6864 31797 7640
rect 31739 6852 31797 6864
rect 31997 7640 32055 7652
rect 31997 6864 32009 7640
rect 32043 6864 32055 7640
rect 31997 6852 32055 6864
rect 32111 7640 32169 7652
rect 32111 6864 32123 7640
rect 32157 6864 32169 7640
rect 32111 6852 32169 6864
rect 32369 7640 32427 7652
rect 32369 6864 32381 7640
rect 32415 6864 32427 7640
rect 32369 6852 32427 6864
rect 32483 7640 32541 7652
rect 32483 6864 32495 7640
rect 32529 6864 32541 7640
rect 32483 6852 32541 6864
rect 32741 7640 32799 7652
rect 32741 6864 32753 7640
rect 32787 6864 32799 7640
rect 32741 6852 32799 6864
rect 32855 7640 32913 7652
rect 32855 6864 32867 7640
rect 32901 6864 32913 7640
rect 32855 6852 32913 6864
rect 33113 7640 33171 7652
rect 33113 6864 33125 7640
rect 33159 6864 33171 7640
rect 33113 6852 33171 6864
rect 30251 6604 30309 6616
rect 30251 5828 30263 6604
rect 30297 5828 30309 6604
rect 30251 5816 30309 5828
rect 30509 6604 30567 6616
rect 30509 5828 30521 6604
rect 30555 5828 30567 6604
rect 30509 5816 30567 5828
rect 30623 6604 30681 6616
rect 30623 5828 30635 6604
rect 30669 5828 30681 6604
rect 30623 5816 30681 5828
rect 30881 6604 30939 6616
rect 30881 5828 30893 6604
rect 30927 5828 30939 6604
rect 30881 5816 30939 5828
rect 30995 6604 31053 6616
rect 30995 5828 31007 6604
rect 31041 5828 31053 6604
rect 30995 5816 31053 5828
rect 31253 6604 31311 6616
rect 31253 5828 31265 6604
rect 31299 5828 31311 6604
rect 31253 5816 31311 5828
rect 31367 6604 31425 6616
rect 31367 5828 31379 6604
rect 31413 5828 31425 6604
rect 31367 5816 31425 5828
rect 31625 6604 31683 6616
rect 31625 5828 31637 6604
rect 31671 5828 31683 6604
rect 31625 5816 31683 5828
rect 31739 6604 31797 6616
rect 31739 5828 31751 6604
rect 31785 5828 31797 6604
rect 31739 5816 31797 5828
rect 31997 6604 32055 6616
rect 31997 5828 32009 6604
rect 32043 5828 32055 6604
rect 31997 5816 32055 5828
rect 32111 6604 32169 6616
rect 32111 5828 32123 6604
rect 32157 5828 32169 6604
rect 32111 5816 32169 5828
rect 32369 6604 32427 6616
rect 32369 5828 32381 6604
rect 32415 5828 32427 6604
rect 32369 5816 32427 5828
rect 32483 6604 32541 6616
rect 32483 5828 32495 6604
rect 32529 5828 32541 6604
rect 32483 5816 32541 5828
rect 32741 6604 32799 6616
rect 32741 5828 32753 6604
rect 32787 5828 32799 6604
rect 32741 5816 32799 5828
rect 32855 6604 32913 6616
rect 32855 5828 32867 6604
rect 32901 5828 32913 6604
rect 32855 5816 32913 5828
rect 33113 6604 33171 6616
rect 33113 5828 33125 6604
rect 33159 5828 33171 6604
rect 33113 5816 33171 5828
<< ndiffc >>
rect 30263 4851 30297 5027
rect 30521 4851 30555 5027
rect 30635 4851 30669 5027
rect 30893 4851 30927 5027
rect 31007 4851 31041 5027
rect 31265 4851 31299 5027
rect 31379 4851 31413 5027
rect 31637 4851 31671 5027
rect 31751 4851 31785 5027
rect 32009 4851 32043 5027
rect 32123 4851 32157 5027
rect 32381 4851 32415 5027
rect 32495 4851 32529 5027
rect 32753 4851 32787 5027
rect 32867 4851 32901 5027
rect 33125 4851 33159 5027
rect 33239 4851 33273 5027
rect 33497 4851 33531 5027
rect 33611 4851 33645 5027
rect 33869 4851 33903 5027
rect 33983 4851 34017 5027
rect 34241 4851 34275 5027
rect 34355 4851 34389 5027
rect 34613 4851 34647 5027
rect 34727 4851 34761 5027
rect 34985 4851 35019 5027
rect 35099 4851 35133 5027
rect 35357 4851 35391 5027
rect 35471 4851 35505 5027
rect 35729 4851 35763 5027
rect 35843 4851 35877 5027
rect 36101 4851 36135 5027
rect 36215 4851 36249 5027
rect 36473 4851 36507 5027
rect 36587 4851 36621 5027
rect 36845 4851 36879 5027
rect 36959 4851 36993 5027
rect 37217 4851 37251 5027
rect 37331 4851 37365 5027
rect 37589 4851 37623 5027
rect 37703 4851 37737 5027
rect 37961 4851 37995 5027
rect 38075 4851 38109 5027
rect 38333 4851 38367 5027
rect 38447 4851 38481 5027
rect 38705 4851 38739 5027
rect 38819 4851 38853 5027
rect 39077 4851 39111 5027
rect 30263 4433 30297 4609
rect 30521 4433 30555 4609
rect 30635 4433 30669 4609
rect 30893 4433 30927 4609
rect 31007 4433 31041 4609
rect 31265 4433 31299 4609
rect 31379 4433 31413 4609
rect 31637 4433 31671 4609
rect 31751 4433 31785 4609
rect 32009 4433 32043 4609
rect 32123 4433 32157 4609
rect 32381 4433 32415 4609
rect 32495 4433 32529 4609
rect 32753 4433 32787 4609
rect 32867 4433 32901 4609
rect 33125 4433 33159 4609
rect 33239 4433 33273 4609
rect 33497 4433 33531 4609
rect 33611 4433 33645 4609
rect 33869 4433 33903 4609
rect 33983 4433 34017 4609
rect 34241 4433 34275 4609
rect 34355 4433 34389 4609
rect 34613 4433 34647 4609
rect 34727 4433 34761 4609
rect 34985 4433 35019 4609
rect 35099 4433 35133 4609
rect 35357 4433 35391 4609
rect 35471 4433 35505 4609
rect 35729 4433 35763 4609
rect 35843 4433 35877 4609
rect 36101 4433 36135 4609
rect 36215 4433 36249 4609
rect 36473 4433 36507 4609
rect 36587 4433 36621 4609
rect 36845 4433 36879 4609
rect 36959 4433 36993 4609
rect 37217 4433 37251 4609
rect 37331 4433 37365 4609
rect 37589 4433 37623 4609
rect 37703 4433 37737 4609
rect 37961 4433 37995 4609
rect 38075 4433 38109 4609
rect 38333 4433 38367 4609
rect 38447 4433 38481 4609
rect 38705 4433 38739 4609
rect 38819 4433 38853 4609
rect 39077 4433 39111 4609
rect 30263 4015 30297 4191
rect 30521 4015 30555 4191
rect 30635 4015 30669 4191
rect 30893 4015 30927 4191
rect 31007 4015 31041 4191
rect 31265 4015 31299 4191
rect 31379 4015 31413 4191
rect 31637 4015 31671 4191
rect 31751 4015 31785 4191
rect 32009 4015 32043 4191
rect 32123 4015 32157 4191
rect 32381 4015 32415 4191
rect 32495 4015 32529 4191
rect 32753 4015 32787 4191
rect 32867 4015 32901 4191
rect 33125 4015 33159 4191
rect 33239 4015 33273 4191
rect 33497 4015 33531 4191
rect 33611 4015 33645 4191
rect 33869 4015 33903 4191
rect 33983 4015 34017 4191
rect 34241 4015 34275 4191
rect 34355 4015 34389 4191
rect 34613 4015 34647 4191
rect 34727 4015 34761 4191
rect 34985 4015 35019 4191
rect 35099 4015 35133 4191
rect 35357 4015 35391 4191
rect 35471 4015 35505 4191
rect 35729 4015 35763 4191
rect 35843 4015 35877 4191
rect 36101 4015 36135 4191
rect 36215 4015 36249 4191
rect 36473 4015 36507 4191
rect 36587 4015 36621 4191
rect 36845 4015 36879 4191
rect 36959 4015 36993 4191
rect 37217 4015 37251 4191
rect 37331 4015 37365 4191
rect 37589 4015 37623 4191
rect 37703 4015 37737 4191
rect 37961 4015 37995 4191
rect 38075 4015 38109 4191
rect 38333 4015 38367 4191
rect 38447 4015 38481 4191
rect 38705 4015 38739 4191
rect 38819 4015 38853 4191
rect 39077 4015 39111 4191
rect 30263 3597 30297 3773
rect 30521 3597 30555 3773
rect 30635 3597 30669 3773
rect 30893 3597 30927 3773
rect 31007 3597 31041 3773
rect 31265 3597 31299 3773
rect 31379 3597 31413 3773
rect 31637 3597 31671 3773
rect 31751 3597 31785 3773
rect 32009 3597 32043 3773
rect 32123 3597 32157 3773
rect 32381 3597 32415 3773
rect 32495 3597 32529 3773
rect 32753 3597 32787 3773
rect 32867 3597 32901 3773
rect 33125 3597 33159 3773
rect 33239 3597 33273 3773
rect 33497 3597 33531 3773
rect 33611 3597 33645 3773
rect 33869 3597 33903 3773
rect 33983 3597 34017 3773
rect 34241 3597 34275 3773
rect 34355 3597 34389 3773
rect 34613 3597 34647 3773
rect 34727 3597 34761 3773
rect 34985 3597 35019 3773
rect 35099 3597 35133 3773
rect 35357 3597 35391 3773
rect 35471 3597 35505 3773
rect 35729 3597 35763 3773
rect 35843 3597 35877 3773
rect 36101 3597 36135 3773
rect 36215 3597 36249 3773
rect 36473 3597 36507 3773
rect 36587 3597 36621 3773
rect 36845 3597 36879 3773
rect 36959 3597 36993 3773
rect 37217 3597 37251 3773
rect 37331 3597 37365 3773
rect 37589 3597 37623 3773
rect 37703 3597 37737 3773
rect 37961 3597 37995 3773
rect 38075 3597 38109 3773
rect 38333 3597 38367 3773
rect 38447 3597 38481 3773
rect 38705 3597 38739 3773
rect 38819 3597 38853 3773
rect 39077 3597 39111 3773
<< pdiffc >>
rect 28775 11724 28809 12100
rect 29033 11724 29067 12100
rect 29147 11724 29181 12100
rect 29405 11724 29439 12100
rect 29519 11724 29553 12100
rect 29777 11724 29811 12100
rect 29891 11724 29925 12100
rect 30149 11724 30183 12100
rect 30263 11724 30297 12100
rect 30521 11724 30555 12100
rect 30635 11724 30669 12100
rect 30893 11724 30927 12100
rect 31007 11724 31041 12100
rect 31265 11724 31299 12100
rect 31379 11724 31413 12100
rect 31637 11724 31671 12100
rect 31751 11724 31785 12100
rect 32009 11724 32043 12100
rect 32123 11724 32157 12100
rect 32381 11724 32415 12100
rect 32495 11724 32529 12100
rect 32753 11724 32787 12100
rect 32867 11724 32901 12100
rect 33125 11724 33159 12100
rect 33239 11724 33273 12100
rect 33497 11724 33531 12100
rect 33611 11724 33645 12100
rect 33869 11724 33903 12100
rect 33983 11724 34017 12100
rect 34241 11724 34275 12100
rect 34355 11724 34389 12100
rect 34613 11724 34647 12100
rect 34727 11724 34761 12100
rect 34985 11724 35019 12100
rect 35099 11724 35133 12100
rect 35357 11724 35391 12100
rect 35471 11724 35505 12100
rect 35729 11724 35763 12100
rect 35843 11724 35877 12100
rect 36101 11724 36135 12100
rect 36215 11724 36249 12100
rect 36473 11724 36507 12100
rect 36587 11724 36621 12100
rect 36845 11724 36879 12100
rect 36959 11724 36993 12100
rect 37217 11724 37251 12100
rect 37331 11724 37365 12100
rect 37589 11724 37623 12100
rect 37703 11724 37737 12100
rect 37961 11724 37995 12100
rect 38075 11724 38109 12100
rect 38333 11724 38367 12100
rect 38447 11724 38481 12100
rect 38705 11724 38739 12100
rect 38819 11724 38853 12100
rect 39077 11724 39111 12100
rect 39191 11724 39225 12100
rect 39449 11724 39483 12100
rect 39563 11724 39597 12100
rect 39821 11724 39855 12100
rect 39935 11724 39969 12100
rect 40193 11724 40227 12100
rect 40307 11724 40341 12100
rect 40565 11724 40599 12100
rect 28775 11088 28809 11464
rect 29033 11088 29067 11464
rect 29147 11088 29181 11464
rect 29405 11088 29439 11464
rect 29519 11088 29553 11464
rect 29777 11088 29811 11464
rect 29891 11088 29925 11464
rect 30149 11088 30183 11464
rect 30263 11088 30297 11464
rect 30521 11088 30555 11464
rect 30635 11088 30669 11464
rect 30893 11088 30927 11464
rect 31007 11088 31041 11464
rect 31265 11088 31299 11464
rect 31379 11088 31413 11464
rect 31637 11088 31671 11464
rect 31751 11088 31785 11464
rect 32009 11088 32043 11464
rect 32123 11088 32157 11464
rect 32381 11088 32415 11464
rect 32495 11088 32529 11464
rect 32753 11088 32787 11464
rect 32867 11088 32901 11464
rect 33125 11088 33159 11464
rect 33239 11088 33273 11464
rect 33497 11088 33531 11464
rect 33611 11088 33645 11464
rect 33869 11088 33903 11464
rect 33983 11088 34017 11464
rect 34241 11088 34275 11464
rect 34355 11088 34389 11464
rect 34613 11088 34647 11464
rect 34727 11088 34761 11464
rect 34985 11088 35019 11464
rect 35099 11088 35133 11464
rect 35357 11088 35391 11464
rect 35471 11088 35505 11464
rect 35729 11088 35763 11464
rect 35843 11088 35877 11464
rect 36101 11088 36135 11464
rect 36215 11088 36249 11464
rect 36473 11088 36507 11464
rect 36587 11088 36621 11464
rect 36845 11088 36879 11464
rect 36959 11088 36993 11464
rect 37217 11088 37251 11464
rect 37331 11088 37365 11464
rect 37589 11088 37623 11464
rect 37703 11088 37737 11464
rect 37961 11088 37995 11464
rect 38075 11088 38109 11464
rect 38333 11088 38367 11464
rect 38447 11088 38481 11464
rect 38705 11088 38739 11464
rect 38819 11088 38853 11464
rect 39077 11088 39111 11464
rect 39191 11088 39225 11464
rect 39449 11088 39483 11464
rect 39563 11088 39597 11464
rect 39821 11088 39855 11464
rect 39935 11088 39969 11464
rect 40193 11088 40227 11464
rect 40307 11088 40341 11464
rect 40565 11088 40599 11464
rect 28775 10452 28809 10828
rect 29033 10452 29067 10828
rect 29147 10452 29181 10828
rect 29405 10452 29439 10828
rect 29519 10452 29553 10828
rect 29777 10452 29811 10828
rect 29891 10452 29925 10828
rect 30149 10452 30183 10828
rect 30263 10452 30297 10828
rect 30521 10452 30555 10828
rect 30635 10452 30669 10828
rect 30893 10452 30927 10828
rect 31007 10452 31041 10828
rect 31265 10452 31299 10828
rect 31379 10452 31413 10828
rect 31637 10452 31671 10828
rect 31751 10452 31785 10828
rect 32009 10452 32043 10828
rect 32123 10452 32157 10828
rect 32381 10452 32415 10828
rect 32495 10452 32529 10828
rect 32753 10452 32787 10828
rect 32867 10452 32901 10828
rect 33125 10452 33159 10828
rect 33239 10452 33273 10828
rect 33497 10452 33531 10828
rect 33611 10452 33645 10828
rect 33869 10452 33903 10828
rect 33983 10452 34017 10828
rect 34241 10452 34275 10828
rect 34355 10452 34389 10828
rect 34613 10452 34647 10828
rect 34727 10452 34761 10828
rect 34985 10452 35019 10828
rect 35099 10452 35133 10828
rect 35357 10452 35391 10828
rect 35471 10452 35505 10828
rect 35729 10452 35763 10828
rect 35843 10452 35877 10828
rect 36101 10452 36135 10828
rect 36215 10452 36249 10828
rect 36473 10452 36507 10828
rect 36587 10452 36621 10828
rect 36845 10452 36879 10828
rect 36959 10452 36993 10828
rect 37217 10452 37251 10828
rect 37331 10452 37365 10828
rect 37589 10452 37623 10828
rect 37703 10452 37737 10828
rect 37961 10452 37995 10828
rect 38075 10452 38109 10828
rect 38333 10452 38367 10828
rect 38447 10452 38481 10828
rect 38705 10452 38739 10828
rect 38819 10452 38853 10828
rect 39077 10452 39111 10828
rect 39191 10452 39225 10828
rect 39449 10452 39483 10828
rect 39563 10452 39597 10828
rect 39821 10452 39855 10828
rect 39935 10452 39969 10828
rect 40193 10452 40227 10828
rect 40307 10452 40341 10828
rect 40565 10452 40599 10828
rect 30263 8936 30297 9712
rect 30521 8936 30555 9712
rect 30635 8936 30669 9712
rect 30893 8936 30927 9712
rect 31007 8936 31041 9712
rect 31265 8936 31299 9712
rect 31379 8936 31413 9712
rect 31637 8936 31671 9712
rect 31751 8936 31785 9712
rect 32009 8936 32043 9712
rect 32123 8936 32157 9712
rect 32381 8936 32415 9712
rect 32495 8936 32529 9712
rect 32753 8936 32787 9712
rect 32867 8936 32901 9712
rect 33125 8936 33159 9712
rect 30263 7900 30297 8676
rect 30521 7900 30555 8676
rect 30635 7900 30669 8676
rect 30893 7900 30927 8676
rect 31007 7900 31041 8676
rect 31265 7900 31299 8676
rect 31379 7900 31413 8676
rect 31637 7900 31671 8676
rect 31751 7900 31785 8676
rect 32009 7900 32043 8676
rect 32123 7900 32157 8676
rect 32381 7900 32415 8676
rect 32495 7900 32529 8676
rect 32753 7900 32787 8676
rect 32867 7900 32901 8676
rect 33125 7900 33159 8676
rect 30263 6864 30297 7640
rect 30521 6864 30555 7640
rect 30635 6864 30669 7640
rect 30893 6864 30927 7640
rect 31007 6864 31041 7640
rect 31265 6864 31299 7640
rect 31379 6864 31413 7640
rect 31637 6864 31671 7640
rect 31751 6864 31785 7640
rect 32009 6864 32043 7640
rect 32123 6864 32157 7640
rect 32381 6864 32415 7640
rect 32495 6864 32529 7640
rect 32753 6864 32787 7640
rect 32867 6864 32901 7640
rect 33125 6864 33159 7640
rect 30263 5828 30297 6604
rect 30521 5828 30555 6604
rect 30635 5828 30669 6604
rect 30893 5828 30927 6604
rect 31007 5828 31041 6604
rect 31265 5828 31299 6604
rect 31379 5828 31413 6604
rect 31637 5828 31671 6604
rect 31751 5828 31785 6604
rect 32009 5828 32043 6604
rect 32123 5828 32157 6604
rect 32381 5828 32415 6604
rect 32495 5828 32529 6604
rect 32753 5828 32787 6604
rect 32867 5828 32901 6604
rect 33125 5828 33159 6604
<< psubdiff >>
rect 33776 7574 33872 7608
rect 34010 7574 34106 7608
rect 33776 7512 33810 7574
rect 34072 7512 34106 7574
rect 33776 6238 33810 6300
rect 34072 6238 34106 6300
rect 33776 6204 33872 6238
rect 34010 6204 34106 6238
rect 30149 5179 30245 5213
rect 39129 5179 39225 5213
rect 30149 5117 30183 5179
rect 39191 5117 39225 5179
rect 30149 3445 30183 3507
rect 39191 3445 39225 3507
rect 30149 3411 30245 3445
rect 39129 3411 39225 3445
<< nsubdiff >>
rect 28661 12261 28757 12295
rect 40617 12261 40713 12295
rect 28661 12199 28695 12261
rect 40679 12199 40713 12261
rect 28661 10291 28695 10353
rect 40679 10291 40713 10353
rect 28661 10257 28757 10291
rect 40617 10257 40713 10291
rect 30149 9873 30245 9907
rect 33177 9873 33273 9907
rect 30149 9811 30183 9873
rect 33239 9811 33273 9873
rect 30149 5667 30183 5729
rect 33239 5667 33273 5729
rect 30149 5633 30245 5667
rect 33177 5633 33273 5667
<< psubdiffcont >>
rect 33872 7574 34010 7608
rect 33776 6300 33810 7512
rect 34072 6300 34106 7512
rect 33872 6204 34010 6238
rect 30245 5179 39129 5213
rect 30149 3507 30183 5117
rect 39191 3507 39225 5117
rect 30245 3411 39129 3445
<< nsubdiffcont >>
rect 28757 12261 40617 12295
rect 28661 10353 28695 12199
rect 40679 10353 40713 12199
rect 28757 10257 40617 10291
rect 30245 9873 33177 9907
rect 30149 5729 30183 9811
rect 33239 5729 33273 9811
rect 30245 5633 33177 5667
<< poly >>
rect 28821 12193 29021 12209
rect 28821 12159 28837 12193
rect 29005 12159 29021 12193
rect 28821 12112 29021 12159
rect 29193 12193 29393 12209
rect 29193 12159 29209 12193
rect 29377 12159 29393 12193
rect 29193 12112 29393 12159
rect 29565 12193 29765 12209
rect 29565 12159 29581 12193
rect 29749 12159 29765 12193
rect 29565 12112 29765 12159
rect 29937 12193 30137 12209
rect 29937 12159 29953 12193
rect 30121 12159 30137 12193
rect 29937 12112 30137 12159
rect 30309 12193 30509 12209
rect 30309 12159 30325 12193
rect 30493 12159 30509 12193
rect 30309 12112 30509 12159
rect 30681 12193 30881 12209
rect 30681 12159 30697 12193
rect 30865 12159 30881 12193
rect 30681 12112 30881 12159
rect 31053 12193 31253 12209
rect 31053 12159 31069 12193
rect 31237 12159 31253 12193
rect 31053 12112 31253 12159
rect 31425 12193 31625 12209
rect 31425 12159 31441 12193
rect 31609 12159 31625 12193
rect 31425 12112 31625 12159
rect 31797 12193 31997 12209
rect 31797 12159 31813 12193
rect 31981 12159 31997 12193
rect 31797 12112 31997 12159
rect 32169 12193 32369 12209
rect 32169 12159 32185 12193
rect 32353 12159 32369 12193
rect 32169 12112 32369 12159
rect 32541 12193 32741 12209
rect 32541 12159 32557 12193
rect 32725 12159 32741 12193
rect 32541 12112 32741 12159
rect 32913 12193 33113 12209
rect 32913 12159 32929 12193
rect 33097 12159 33113 12193
rect 32913 12112 33113 12159
rect 33285 12193 33485 12209
rect 33285 12159 33301 12193
rect 33469 12159 33485 12193
rect 33285 12112 33485 12159
rect 33657 12193 33857 12209
rect 33657 12159 33673 12193
rect 33841 12159 33857 12193
rect 33657 12112 33857 12159
rect 34029 12193 34229 12209
rect 34029 12159 34045 12193
rect 34213 12159 34229 12193
rect 34029 12112 34229 12159
rect 34401 12193 34601 12209
rect 34401 12159 34417 12193
rect 34585 12159 34601 12193
rect 34401 12112 34601 12159
rect 34773 12193 34973 12209
rect 34773 12159 34789 12193
rect 34957 12159 34973 12193
rect 34773 12112 34973 12159
rect 35145 12193 35345 12209
rect 35145 12159 35161 12193
rect 35329 12159 35345 12193
rect 35145 12112 35345 12159
rect 35517 12193 35717 12209
rect 35517 12159 35533 12193
rect 35701 12159 35717 12193
rect 35517 12112 35717 12159
rect 35889 12193 36089 12209
rect 35889 12159 35905 12193
rect 36073 12159 36089 12193
rect 35889 12112 36089 12159
rect 36261 12193 36461 12209
rect 36261 12159 36277 12193
rect 36445 12159 36461 12193
rect 36261 12112 36461 12159
rect 36633 12193 36833 12209
rect 36633 12159 36649 12193
rect 36817 12159 36833 12193
rect 36633 12112 36833 12159
rect 37005 12193 37205 12209
rect 37005 12159 37021 12193
rect 37189 12159 37205 12193
rect 37005 12112 37205 12159
rect 37377 12193 37577 12209
rect 37377 12159 37393 12193
rect 37561 12159 37577 12193
rect 37377 12112 37577 12159
rect 37749 12193 37949 12209
rect 37749 12159 37765 12193
rect 37933 12159 37949 12193
rect 37749 12112 37949 12159
rect 38121 12193 38321 12209
rect 38121 12159 38137 12193
rect 38305 12159 38321 12193
rect 38121 12112 38321 12159
rect 38493 12193 38693 12209
rect 38493 12159 38509 12193
rect 38677 12159 38693 12193
rect 38493 12112 38693 12159
rect 38865 12193 39065 12209
rect 38865 12159 38881 12193
rect 39049 12159 39065 12193
rect 38865 12112 39065 12159
rect 39237 12193 39437 12209
rect 39237 12159 39253 12193
rect 39421 12159 39437 12193
rect 39237 12112 39437 12159
rect 39609 12193 39809 12209
rect 39609 12159 39625 12193
rect 39793 12159 39809 12193
rect 39609 12112 39809 12159
rect 39981 12193 40181 12209
rect 39981 12159 39997 12193
rect 40165 12159 40181 12193
rect 39981 12112 40181 12159
rect 40353 12193 40553 12209
rect 40353 12159 40369 12193
rect 40537 12159 40553 12193
rect 40353 12112 40553 12159
rect 28821 11665 29021 11712
rect 28821 11631 28837 11665
rect 29005 11631 29021 11665
rect 28821 11615 29021 11631
rect 29193 11665 29393 11712
rect 29193 11631 29209 11665
rect 29377 11631 29393 11665
rect 29193 11615 29393 11631
rect 29565 11665 29765 11712
rect 29565 11631 29581 11665
rect 29749 11631 29765 11665
rect 29565 11615 29765 11631
rect 29937 11665 30137 11712
rect 29937 11631 29953 11665
rect 30121 11631 30137 11665
rect 29937 11615 30137 11631
rect 30309 11665 30509 11712
rect 30309 11631 30325 11665
rect 30493 11631 30509 11665
rect 30309 11615 30509 11631
rect 30681 11665 30881 11712
rect 30681 11631 30697 11665
rect 30865 11631 30881 11665
rect 30681 11615 30881 11631
rect 31053 11665 31253 11712
rect 31053 11631 31069 11665
rect 31237 11631 31253 11665
rect 31053 11615 31253 11631
rect 31425 11665 31625 11712
rect 31425 11631 31441 11665
rect 31609 11631 31625 11665
rect 31425 11615 31625 11631
rect 31797 11665 31997 11712
rect 31797 11631 31813 11665
rect 31981 11631 31997 11665
rect 31797 11615 31997 11631
rect 32169 11665 32369 11712
rect 32169 11631 32185 11665
rect 32353 11631 32369 11665
rect 32169 11615 32369 11631
rect 32541 11665 32741 11712
rect 32541 11631 32557 11665
rect 32725 11631 32741 11665
rect 32541 11615 32741 11631
rect 32913 11665 33113 11712
rect 32913 11631 32929 11665
rect 33097 11631 33113 11665
rect 32913 11615 33113 11631
rect 33285 11665 33485 11712
rect 33285 11631 33301 11665
rect 33469 11631 33485 11665
rect 33285 11615 33485 11631
rect 33657 11665 33857 11712
rect 33657 11631 33673 11665
rect 33841 11631 33857 11665
rect 33657 11615 33857 11631
rect 34029 11665 34229 11712
rect 34029 11631 34045 11665
rect 34213 11631 34229 11665
rect 34029 11615 34229 11631
rect 34401 11665 34601 11712
rect 34401 11631 34417 11665
rect 34585 11631 34601 11665
rect 34401 11615 34601 11631
rect 34773 11665 34973 11712
rect 34773 11631 34789 11665
rect 34957 11631 34973 11665
rect 34773 11615 34973 11631
rect 35145 11665 35345 11712
rect 35145 11631 35161 11665
rect 35329 11631 35345 11665
rect 35145 11615 35345 11631
rect 35517 11665 35717 11712
rect 35517 11631 35533 11665
rect 35701 11631 35717 11665
rect 35517 11615 35717 11631
rect 35889 11665 36089 11712
rect 35889 11631 35905 11665
rect 36073 11631 36089 11665
rect 35889 11615 36089 11631
rect 36261 11665 36461 11712
rect 36261 11631 36277 11665
rect 36445 11631 36461 11665
rect 36261 11615 36461 11631
rect 36633 11665 36833 11712
rect 36633 11631 36649 11665
rect 36817 11631 36833 11665
rect 36633 11615 36833 11631
rect 37005 11665 37205 11712
rect 37005 11631 37021 11665
rect 37189 11631 37205 11665
rect 37005 11615 37205 11631
rect 37377 11665 37577 11712
rect 37377 11631 37393 11665
rect 37561 11631 37577 11665
rect 37377 11615 37577 11631
rect 37749 11665 37949 11712
rect 37749 11631 37765 11665
rect 37933 11631 37949 11665
rect 37749 11615 37949 11631
rect 38121 11665 38321 11712
rect 38121 11631 38137 11665
rect 38305 11631 38321 11665
rect 38121 11615 38321 11631
rect 38493 11665 38693 11712
rect 38493 11631 38509 11665
rect 38677 11631 38693 11665
rect 38493 11615 38693 11631
rect 38865 11665 39065 11712
rect 38865 11631 38881 11665
rect 39049 11631 39065 11665
rect 38865 11615 39065 11631
rect 39237 11665 39437 11712
rect 39237 11631 39253 11665
rect 39421 11631 39437 11665
rect 39237 11615 39437 11631
rect 39609 11665 39809 11712
rect 39609 11631 39625 11665
rect 39793 11631 39809 11665
rect 39609 11615 39809 11631
rect 39981 11665 40181 11712
rect 39981 11631 39997 11665
rect 40165 11631 40181 11665
rect 39981 11615 40181 11631
rect 40353 11665 40553 11712
rect 40353 11631 40369 11665
rect 40537 11631 40553 11665
rect 40353 11615 40553 11631
rect 28821 11557 29021 11573
rect 28821 11523 28837 11557
rect 29005 11523 29021 11557
rect 28821 11476 29021 11523
rect 29193 11557 29393 11573
rect 29193 11523 29209 11557
rect 29377 11523 29393 11557
rect 29193 11476 29393 11523
rect 29565 11557 29765 11573
rect 29565 11523 29581 11557
rect 29749 11523 29765 11557
rect 29565 11476 29765 11523
rect 29937 11557 30137 11573
rect 29937 11523 29953 11557
rect 30121 11523 30137 11557
rect 29937 11476 30137 11523
rect 30309 11557 30509 11573
rect 30309 11523 30325 11557
rect 30493 11523 30509 11557
rect 30309 11476 30509 11523
rect 30681 11557 30881 11573
rect 30681 11523 30697 11557
rect 30865 11523 30881 11557
rect 30681 11476 30881 11523
rect 31053 11557 31253 11573
rect 31053 11523 31069 11557
rect 31237 11523 31253 11557
rect 31053 11476 31253 11523
rect 31425 11557 31625 11573
rect 31425 11523 31441 11557
rect 31609 11523 31625 11557
rect 31425 11476 31625 11523
rect 31797 11557 31997 11573
rect 31797 11523 31813 11557
rect 31981 11523 31997 11557
rect 31797 11476 31997 11523
rect 32169 11557 32369 11573
rect 32169 11523 32185 11557
rect 32353 11523 32369 11557
rect 32169 11476 32369 11523
rect 32541 11557 32741 11573
rect 32541 11523 32557 11557
rect 32725 11523 32741 11557
rect 32541 11476 32741 11523
rect 32913 11557 33113 11573
rect 32913 11523 32929 11557
rect 33097 11523 33113 11557
rect 32913 11476 33113 11523
rect 33285 11557 33485 11573
rect 33285 11523 33301 11557
rect 33469 11523 33485 11557
rect 33285 11476 33485 11523
rect 33657 11557 33857 11573
rect 33657 11523 33673 11557
rect 33841 11523 33857 11557
rect 33657 11476 33857 11523
rect 34029 11557 34229 11573
rect 34029 11523 34045 11557
rect 34213 11523 34229 11557
rect 34029 11476 34229 11523
rect 34401 11557 34601 11573
rect 34401 11523 34417 11557
rect 34585 11523 34601 11557
rect 34401 11476 34601 11523
rect 34773 11557 34973 11573
rect 34773 11523 34789 11557
rect 34957 11523 34973 11557
rect 34773 11476 34973 11523
rect 35145 11557 35345 11573
rect 35145 11523 35161 11557
rect 35329 11523 35345 11557
rect 35145 11476 35345 11523
rect 35517 11557 35717 11573
rect 35517 11523 35533 11557
rect 35701 11523 35717 11557
rect 35517 11476 35717 11523
rect 35889 11557 36089 11573
rect 35889 11523 35905 11557
rect 36073 11523 36089 11557
rect 35889 11476 36089 11523
rect 36261 11557 36461 11573
rect 36261 11523 36277 11557
rect 36445 11523 36461 11557
rect 36261 11476 36461 11523
rect 36633 11557 36833 11573
rect 36633 11523 36649 11557
rect 36817 11523 36833 11557
rect 36633 11476 36833 11523
rect 37005 11557 37205 11573
rect 37005 11523 37021 11557
rect 37189 11523 37205 11557
rect 37005 11476 37205 11523
rect 37377 11557 37577 11573
rect 37377 11523 37393 11557
rect 37561 11523 37577 11557
rect 37377 11476 37577 11523
rect 37749 11557 37949 11573
rect 37749 11523 37765 11557
rect 37933 11523 37949 11557
rect 37749 11476 37949 11523
rect 38121 11557 38321 11573
rect 38121 11523 38137 11557
rect 38305 11523 38321 11557
rect 38121 11476 38321 11523
rect 38493 11557 38693 11573
rect 38493 11523 38509 11557
rect 38677 11523 38693 11557
rect 38493 11476 38693 11523
rect 38865 11557 39065 11573
rect 38865 11523 38881 11557
rect 39049 11523 39065 11557
rect 38865 11476 39065 11523
rect 39237 11557 39437 11573
rect 39237 11523 39253 11557
rect 39421 11523 39437 11557
rect 39237 11476 39437 11523
rect 39609 11557 39809 11573
rect 39609 11523 39625 11557
rect 39793 11523 39809 11557
rect 39609 11476 39809 11523
rect 39981 11557 40181 11573
rect 39981 11523 39997 11557
rect 40165 11523 40181 11557
rect 39981 11476 40181 11523
rect 40353 11557 40553 11573
rect 40353 11523 40369 11557
rect 40537 11523 40553 11557
rect 40353 11476 40553 11523
rect 28821 11029 29021 11076
rect 28821 10995 28837 11029
rect 29005 10995 29021 11029
rect 28821 10979 29021 10995
rect 29193 11029 29393 11076
rect 29193 10995 29209 11029
rect 29377 10995 29393 11029
rect 29193 10979 29393 10995
rect 29565 11029 29765 11076
rect 29565 10995 29581 11029
rect 29749 10995 29765 11029
rect 29565 10979 29765 10995
rect 29937 11029 30137 11076
rect 29937 10995 29953 11029
rect 30121 10995 30137 11029
rect 29937 10979 30137 10995
rect 30309 11029 30509 11076
rect 30309 10995 30325 11029
rect 30493 10995 30509 11029
rect 30309 10979 30509 10995
rect 30681 11029 30881 11076
rect 30681 10995 30697 11029
rect 30865 10995 30881 11029
rect 30681 10979 30881 10995
rect 31053 11029 31253 11076
rect 31053 10995 31069 11029
rect 31237 10995 31253 11029
rect 31053 10979 31253 10995
rect 31425 11029 31625 11076
rect 31425 10995 31441 11029
rect 31609 10995 31625 11029
rect 31425 10979 31625 10995
rect 31797 11029 31997 11076
rect 31797 10995 31813 11029
rect 31981 10995 31997 11029
rect 31797 10979 31997 10995
rect 32169 11029 32369 11076
rect 32169 10995 32185 11029
rect 32353 10995 32369 11029
rect 32169 10979 32369 10995
rect 32541 11029 32741 11076
rect 32541 10995 32557 11029
rect 32725 10995 32741 11029
rect 32541 10979 32741 10995
rect 32913 11029 33113 11076
rect 32913 10995 32929 11029
rect 33097 10995 33113 11029
rect 32913 10979 33113 10995
rect 33285 11029 33485 11076
rect 33285 10995 33301 11029
rect 33469 10995 33485 11029
rect 33285 10979 33485 10995
rect 33657 11029 33857 11076
rect 33657 10995 33673 11029
rect 33841 10995 33857 11029
rect 33657 10979 33857 10995
rect 34029 11029 34229 11076
rect 34029 10995 34045 11029
rect 34213 10995 34229 11029
rect 34029 10979 34229 10995
rect 34401 11029 34601 11076
rect 34401 10995 34417 11029
rect 34585 10995 34601 11029
rect 34401 10979 34601 10995
rect 34773 11029 34973 11076
rect 34773 10995 34789 11029
rect 34957 10995 34973 11029
rect 34773 10979 34973 10995
rect 35145 11029 35345 11076
rect 35145 10995 35161 11029
rect 35329 10995 35345 11029
rect 35145 10979 35345 10995
rect 35517 11029 35717 11076
rect 35517 10995 35533 11029
rect 35701 10995 35717 11029
rect 35517 10979 35717 10995
rect 35889 11029 36089 11076
rect 35889 10995 35905 11029
rect 36073 10995 36089 11029
rect 35889 10979 36089 10995
rect 36261 11029 36461 11076
rect 36261 10995 36277 11029
rect 36445 10995 36461 11029
rect 36261 10979 36461 10995
rect 36633 11029 36833 11076
rect 36633 10995 36649 11029
rect 36817 10995 36833 11029
rect 36633 10979 36833 10995
rect 37005 11029 37205 11076
rect 37005 10995 37021 11029
rect 37189 10995 37205 11029
rect 37005 10979 37205 10995
rect 37377 11029 37577 11076
rect 37377 10995 37393 11029
rect 37561 10995 37577 11029
rect 37377 10979 37577 10995
rect 37749 11029 37949 11076
rect 37749 10995 37765 11029
rect 37933 10995 37949 11029
rect 37749 10979 37949 10995
rect 38121 11029 38321 11076
rect 38121 10995 38137 11029
rect 38305 10995 38321 11029
rect 38121 10979 38321 10995
rect 38493 11029 38693 11076
rect 38493 10995 38509 11029
rect 38677 10995 38693 11029
rect 38493 10979 38693 10995
rect 38865 11029 39065 11076
rect 38865 10995 38881 11029
rect 39049 10995 39065 11029
rect 38865 10979 39065 10995
rect 39237 11029 39437 11076
rect 39237 10995 39253 11029
rect 39421 10995 39437 11029
rect 39237 10979 39437 10995
rect 39609 11029 39809 11076
rect 39609 10995 39625 11029
rect 39793 10995 39809 11029
rect 39609 10979 39809 10995
rect 39981 11029 40181 11076
rect 39981 10995 39997 11029
rect 40165 10995 40181 11029
rect 39981 10979 40181 10995
rect 40353 11029 40553 11076
rect 40353 10995 40369 11029
rect 40537 10995 40553 11029
rect 40353 10979 40553 10995
rect 28821 10921 29021 10937
rect 28821 10887 28837 10921
rect 29005 10887 29021 10921
rect 28821 10840 29021 10887
rect 29193 10921 29393 10937
rect 29193 10887 29209 10921
rect 29377 10887 29393 10921
rect 29193 10840 29393 10887
rect 29565 10921 29765 10937
rect 29565 10887 29581 10921
rect 29749 10887 29765 10921
rect 29565 10840 29765 10887
rect 29937 10921 30137 10937
rect 29937 10887 29953 10921
rect 30121 10887 30137 10921
rect 29937 10840 30137 10887
rect 30309 10921 30509 10937
rect 30309 10887 30325 10921
rect 30493 10887 30509 10921
rect 30309 10840 30509 10887
rect 30681 10921 30881 10937
rect 30681 10887 30697 10921
rect 30865 10887 30881 10921
rect 30681 10840 30881 10887
rect 31053 10921 31253 10937
rect 31053 10887 31069 10921
rect 31237 10887 31253 10921
rect 31053 10840 31253 10887
rect 31425 10921 31625 10937
rect 31425 10887 31441 10921
rect 31609 10887 31625 10921
rect 31425 10840 31625 10887
rect 31797 10921 31997 10937
rect 31797 10887 31813 10921
rect 31981 10887 31997 10921
rect 31797 10840 31997 10887
rect 32169 10921 32369 10937
rect 32169 10887 32185 10921
rect 32353 10887 32369 10921
rect 32169 10840 32369 10887
rect 32541 10921 32741 10937
rect 32541 10887 32557 10921
rect 32725 10887 32741 10921
rect 32541 10840 32741 10887
rect 32913 10921 33113 10937
rect 32913 10887 32929 10921
rect 33097 10887 33113 10921
rect 32913 10840 33113 10887
rect 33285 10921 33485 10937
rect 33285 10887 33301 10921
rect 33469 10887 33485 10921
rect 33285 10840 33485 10887
rect 33657 10921 33857 10937
rect 33657 10887 33673 10921
rect 33841 10887 33857 10921
rect 33657 10840 33857 10887
rect 34029 10921 34229 10937
rect 34029 10887 34045 10921
rect 34213 10887 34229 10921
rect 34029 10840 34229 10887
rect 34401 10921 34601 10937
rect 34401 10887 34417 10921
rect 34585 10887 34601 10921
rect 34401 10840 34601 10887
rect 34773 10921 34973 10937
rect 34773 10887 34789 10921
rect 34957 10887 34973 10921
rect 34773 10840 34973 10887
rect 35145 10921 35345 10937
rect 35145 10887 35161 10921
rect 35329 10887 35345 10921
rect 35145 10840 35345 10887
rect 35517 10921 35717 10937
rect 35517 10887 35533 10921
rect 35701 10887 35717 10921
rect 35517 10840 35717 10887
rect 35889 10921 36089 10937
rect 35889 10887 35905 10921
rect 36073 10887 36089 10921
rect 35889 10840 36089 10887
rect 36261 10921 36461 10937
rect 36261 10887 36277 10921
rect 36445 10887 36461 10921
rect 36261 10840 36461 10887
rect 36633 10921 36833 10937
rect 36633 10887 36649 10921
rect 36817 10887 36833 10921
rect 36633 10840 36833 10887
rect 37005 10921 37205 10937
rect 37005 10887 37021 10921
rect 37189 10887 37205 10921
rect 37005 10840 37205 10887
rect 37377 10921 37577 10937
rect 37377 10887 37393 10921
rect 37561 10887 37577 10921
rect 37377 10840 37577 10887
rect 37749 10921 37949 10937
rect 37749 10887 37765 10921
rect 37933 10887 37949 10921
rect 37749 10840 37949 10887
rect 38121 10921 38321 10937
rect 38121 10887 38137 10921
rect 38305 10887 38321 10921
rect 38121 10840 38321 10887
rect 38493 10921 38693 10937
rect 38493 10887 38509 10921
rect 38677 10887 38693 10921
rect 38493 10840 38693 10887
rect 38865 10921 39065 10937
rect 38865 10887 38881 10921
rect 39049 10887 39065 10921
rect 38865 10840 39065 10887
rect 39237 10921 39437 10937
rect 39237 10887 39253 10921
rect 39421 10887 39437 10921
rect 39237 10840 39437 10887
rect 39609 10921 39809 10937
rect 39609 10887 39625 10921
rect 39793 10887 39809 10921
rect 39609 10840 39809 10887
rect 39981 10921 40181 10937
rect 39981 10887 39997 10921
rect 40165 10887 40181 10921
rect 39981 10840 40181 10887
rect 40353 10921 40553 10937
rect 40353 10887 40369 10921
rect 40537 10887 40553 10921
rect 40353 10840 40553 10887
rect 28821 10393 29021 10440
rect 28821 10359 28837 10393
rect 29005 10359 29021 10393
rect 28821 10343 29021 10359
rect 29193 10393 29393 10440
rect 29193 10359 29209 10393
rect 29377 10359 29393 10393
rect 29193 10343 29393 10359
rect 29565 10393 29765 10440
rect 29565 10359 29581 10393
rect 29749 10359 29765 10393
rect 29565 10343 29765 10359
rect 29937 10393 30137 10440
rect 29937 10359 29953 10393
rect 30121 10359 30137 10393
rect 29937 10343 30137 10359
rect 30309 10393 30509 10440
rect 30309 10359 30325 10393
rect 30493 10359 30509 10393
rect 30309 10343 30509 10359
rect 30681 10393 30881 10440
rect 30681 10359 30697 10393
rect 30865 10359 30881 10393
rect 30681 10343 30881 10359
rect 31053 10393 31253 10440
rect 31053 10359 31069 10393
rect 31237 10359 31253 10393
rect 31053 10343 31253 10359
rect 31425 10393 31625 10440
rect 31425 10359 31441 10393
rect 31609 10359 31625 10393
rect 31425 10343 31625 10359
rect 31797 10393 31997 10440
rect 31797 10359 31813 10393
rect 31981 10359 31997 10393
rect 31797 10343 31997 10359
rect 32169 10393 32369 10440
rect 32169 10359 32185 10393
rect 32353 10359 32369 10393
rect 32169 10343 32369 10359
rect 32541 10393 32741 10440
rect 32541 10359 32557 10393
rect 32725 10359 32741 10393
rect 32541 10343 32741 10359
rect 32913 10393 33113 10440
rect 32913 10359 32929 10393
rect 33097 10359 33113 10393
rect 32913 10343 33113 10359
rect 33285 10393 33485 10440
rect 33285 10359 33301 10393
rect 33469 10359 33485 10393
rect 33285 10343 33485 10359
rect 33657 10393 33857 10440
rect 33657 10359 33673 10393
rect 33841 10359 33857 10393
rect 33657 10343 33857 10359
rect 34029 10393 34229 10440
rect 34029 10359 34045 10393
rect 34213 10359 34229 10393
rect 34029 10343 34229 10359
rect 34401 10393 34601 10440
rect 34401 10359 34417 10393
rect 34585 10359 34601 10393
rect 34401 10343 34601 10359
rect 34773 10393 34973 10440
rect 34773 10359 34789 10393
rect 34957 10359 34973 10393
rect 34773 10343 34973 10359
rect 35145 10393 35345 10440
rect 35145 10359 35161 10393
rect 35329 10359 35345 10393
rect 35145 10343 35345 10359
rect 35517 10393 35717 10440
rect 35517 10359 35533 10393
rect 35701 10359 35717 10393
rect 35517 10343 35717 10359
rect 35889 10393 36089 10440
rect 35889 10359 35905 10393
rect 36073 10359 36089 10393
rect 35889 10343 36089 10359
rect 36261 10393 36461 10440
rect 36261 10359 36277 10393
rect 36445 10359 36461 10393
rect 36261 10343 36461 10359
rect 36633 10393 36833 10440
rect 36633 10359 36649 10393
rect 36817 10359 36833 10393
rect 36633 10343 36833 10359
rect 37005 10393 37205 10440
rect 37005 10359 37021 10393
rect 37189 10359 37205 10393
rect 37005 10343 37205 10359
rect 37377 10393 37577 10440
rect 37377 10359 37393 10393
rect 37561 10359 37577 10393
rect 37377 10343 37577 10359
rect 37749 10393 37949 10440
rect 37749 10359 37765 10393
rect 37933 10359 37949 10393
rect 37749 10343 37949 10359
rect 38121 10393 38321 10440
rect 38121 10359 38137 10393
rect 38305 10359 38321 10393
rect 38121 10343 38321 10359
rect 38493 10393 38693 10440
rect 38493 10359 38509 10393
rect 38677 10359 38693 10393
rect 38493 10343 38693 10359
rect 38865 10393 39065 10440
rect 38865 10359 38881 10393
rect 39049 10359 39065 10393
rect 38865 10343 39065 10359
rect 39237 10393 39437 10440
rect 39237 10359 39253 10393
rect 39421 10359 39437 10393
rect 39237 10343 39437 10359
rect 39609 10393 39809 10440
rect 39609 10359 39625 10393
rect 39793 10359 39809 10393
rect 39609 10343 39809 10359
rect 39981 10393 40181 10440
rect 39981 10359 39997 10393
rect 40165 10359 40181 10393
rect 39981 10343 40181 10359
rect 40353 10393 40553 10440
rect 40353 10359 40369 10393
rect 40537 10359 40553 10393
rect 40353 10343 40553 10359
rect 30309 9805 30509 9821
rect 30309 9771 30325 9805
rect 30493 9771 30509 9805
rect 30309 9724 30509 9771
rect 30681 9805 30881 9821
rect 30681 9771 30697 9805
rect 30865 9771 30881 9805
rect 30681 9724 30881 9771
rect 31053 9805 31253 9821
rect 31053 9771 31069 9805
rect 31237 9771 31253 9805
rect 31053 9724 31253 9771
rect 31425 9805 31625 9821
rect 31425 9771 31441 9805
rect 31609 9771 31625 9805
rect 31425 9724 31625 9771
rect 31797 9805 31997 9821
rect 31797 9771 31813 9805
rect 31981 9771 31997 9805
rect 31797 9724 31997 9771
rect 32169 9805 32369 9821
rect 32169 9771 32185 9805
rect 32353 9771 32369 9805
rect 32169 9724 32369 9771
rect 32541 9805 32741 9821
rect 32541 9771 32557 9805
rect 32725 9771 32741 9805
rect 32541 9724 32741 9771
rect 32913 9805 33113 9821
rect 32913 9771 32929 9805
rect 33097 9771 33113 9805
rect 32913 9724 33113 9771
rect 30309 8877 30509 8924
rect 30309 8843 30325 8877
rect 30493 8843 30509 8877
rect 30309 8827 30509 8843
rect 30681 8877 30881 8924
rect 30681 8843 30697 8877
rect 30865 8843 30881 8877
rect 30681 8827 30881 8843
rect 31053 8877 31253 8924
rect 31053 8843 31069 8877
rect 31237 8843 31253 8877
rect 31053 8827 31253 8843
rect 31425 8877 31625 8924
rect 31425 8843 31441 8877
rect 31609 8843 31625 8877
rect 31425 8827 31625 8843
rect 31797 8877 31997 8924
rect 31797 8843 31813 8877
rect 31981 8843 31997 8877
rect 31797 8827 31997 8843
rect 32169 8877 32369 8924
rect 32169 8843 32185 8877
rect 32353 8843 32369 8877
rect 32169 8827 32369 8843
rect 32541 8877 32741 8924
rect 32541 8843 32557 8877
rect 32725 8843 32741 8877
rect 32541 8827 32741 8843
rect 32913 8877 33113 8924
rect 32913 8843 32929 8877
rect 33097 8843 33113 8877
rect 32913 8827 33113 8843
rect 30309 8769 30509 8785
rect 30309 8735 30325 8769
rect 30493 8735 30509 8769
rect 30309 8688 30509 8735
rect 30681 8769 30881 8785
rect 30681 8735 30697 8769
rect 30865 8735 30881 8769
rect 30681 8688 30881 8735
rect 31053 8769 31253 8785
rect 31053 8735 31069 8769
rect 31237 8735 31253 8769
rect 31053 8688 31253 8735
rect 31425 8769 31625 8785
rect 31425 8735 31441 8769
rect 31609 8735 31625 8769
rect 31425 8688 31625 8735
rect 31797 8769 31997 8785
rect 31797 8735 31813 8769
rect 31981 8735 31997 8769
rect 31797 8688 31997 8735
rect 32169 8769 32369 8785
rect 32169 8735 32185 8769
rect 32353 8735 32369 8769
rect 32169 8688 32369 8735
rect 32541 8769 32741 8785
rect 32541 8735 32557 8769
rect 32725 8735 32741 8769
rect 32541 8688 32741 8735
rect 32913 8769 33113 8785
rect 32913 8735 32929 8769
rect 33097 8735 33113 8769
rect 32913 8688 33113 8735
rect 30309 7841 30509 7888
rect 30309 7807 30325 7841
rect 30493 7807 30509 7841
rect 30309 7791 30509 7807
rect 30681 7841 30881 7888
rect 30681 7807 30697 7841
rect 30865 7807 30881 7841
rect 30681 7791 30881 7807
rect 31053 7841 31253 7888
rect 31053 7807 31069 7841
rect 31237 7807 31253 7841
rect 31053 7791 31253 7807
rect 31425 7841 31625 7888
rect 31425 7807 31441 7841
rect 31609 7807 31625 7841
rect 31425 7791 31625 7807
rect 31797 7841 31997 7888
rect 31797 7807 31813 7841
rect 31981 7807 31997 7841
rect 31797 7791 31997 7807
rect 32169 7841 32369 7888
rect 32169 7807 32185 7841
rect 32353 7807 32369 7841
rect 32169 7791 32369 7807
rect 32541 7841 32741 7888
rect 32541 7807 32557 7841
rect 32725 7807 32741 7841
rect 32541 7791 32741 7807
rect 32913 7841 33113 7888
rect 32913 7807 32929 7841
rect 33097 7807 33113 7841
rect 32913 7791 33113 7807
rect 30309 7733 30509 7749
rect 30309 7699 30325 7733
rect 30493 7699 30509 7733
rect 30309 7652 30509 7699
rect 30681 7733 30881 7749
rect 30681 7699 30697 7733
rect 30865 7699 30881 7733
rect 30681 7652 30881 7699
rect 31053 7733 31253 7749
rect 31053 7699 31069 7733
rect 31237 7699 31253 7733
rect 31053 7652 31253 7699
rect 31425 7733 31625 7749
rect 31425 7699 31441 7733
rect 31609 7699 31625 7733
rect 31425 7652 31625 7699
rect 31797 7733 31997 7749
rect 31797 7699 31813 7733
rect 31981 7699 31997 7733
rect 31797 7652 31997 7699
rect 32169 7733 32369 7749
rect 32169 7699 32185 7733
rect 32353 7699 32369 7733
rect 32169 7652 32369 7699
rect 32541 7733 32741 7749
rect 32541 7699 32557 7733
rect 32725 7699 32741 7733
rect 32541 7652 32741 7699
rect 32913 7733 33113 7749
rect 32913 7699 32929 7733
rect 33097 7699 33113 7733
rect 32913 7652 33113 7699
rect 30309 6805 30509 6852
rect 30309 6771 30325 6805
rect 30493 6771 30509 6805
rect 30309 6755 30509 6771
rect 30681 6805 30881 6852
rect 30681 6771 30697 6805
rect 30865 6771 30881 6805
rect 30681 6755 30881 6771
rect 31053 6805 31253 6852
rect 31053 6771 31069 6805
rect 31237 6771 31253 6805
rect 31053 6755 31253 6771
rect 31425 6805 31625 6852
rect 31425 6771 31441 6805
rect 31609 6771 31625 6805
rect 31425 6755 31625 6771
rect 31797 6805 31997 6852
rect 31797 6771 31813 6805
rect 31981 6771 31997 6805
rect 31797 6755 31997 6771
rect 32169 6805 32369 6852
rect 32169 6771 32185 6805
rect 32353 6771 32369 6805
rect 32169 6755 32369 6771
rect 32541 6805 32741 6852
rect 32541 6771 32557 6805
rect 32725 6771 32741 6805
rect 32541 6755 32741 6771
rect 32913 6805 33113 6852
rect 32913 6771 32929 6805
rect 33097 6771 33113 6805
rect 32913 6755 33113 6771
rect 30309 6697 30509 6713
rect 30309 6663 30325 6697
rect 30493 6663 30509 6697
rect 30309 6616 30509 6663
rect 30681 6697 30881 6713
rect 30681 6663 30697 6697
rect 30865 6663 30881 6697
rect 30681 6616 30881 6663
rect 31053 6697 31253 6713
rect 31053 6663 31069 6697
rect 31237 6663 31253 6697
rect 31053 6616 31253 6663
rect 31425 6697 31625 6713
rect 31425 6663 31441 6697
rect 31609 6663 31625 6697
rect 31425 6616 31625 6663
rect 31797 6697 31997 6713
rect 31797 6663 31813 6697
rect 31981 6663 31997 6697
rect 31797 6616 31997 6663
rect 32169 6697 32369 6713
rect 32169 6663 32185 6697
rect 32353 6663 32369 6697
rect 32169 6616 32369 6663
rect 32541 6697 32741 6713
rect 32541 6663 32557 6697
rect 32725 6663 32741 6697
rect 32541 6616 32741 6663
rect 32913 6697 33113 6713
rect 32913 6663 32929 6697
rect 33097 6663 33113 6697
rect 32913 6616 33113 6663
rect 30309 5769 30509 5816
rect 30309 5735 30325 5769
rect 30493 5735 30509 5769
rect 30309 5719 30509 5735
rect 30681 5769 30881 5816
rect 30681 5735 30697 5769
rect 30865 5735 30881 5769
rect 30681 5719 30881 5735
rect 31053 5769 31253 5816
rect 31053 5735 31069 5769
rect 31237 5735 31253 5769
rect 31053 5719 31253 5735
rect 31425 5769 31625 5816
rect 31425 5735 31441 5769
rect 31609 5735 31625 5769
rect 31425 5719 31625 5735
rect 31797 5769 31997 5816
rect 31797 5735 31813 5769
rect 31981 5735 31997 5769
rect 31797 5719 31997 5735
rect 32169 5769 32369 5816
rect 32169 5735 32185 5769
rect 32353 5735 32369 5769
rect 32169 5719 32369 5735
rect 32541 5769 32741 5816
rect 32541 5735 32557 5769
rect 32725 5735 32741 5769
rect 32541 5719 32741 5735
rect 32913 5769 33113 5816
rect 32913 5735 32929 5769
rect 33097 5735 33113 5769
rect 32913 5719 33113 5735
rect 30309 5111 30509 5127
rect 30309 5077 30325 5111
rect 30493 5077 30509 5111
rect 30309 5039 30509 5077
rect 30681 5111 30881 5127
rect 30681 5077 30697 5111
rect 30865 5077 30881 5111
rect 30681 5039 30881 5077
rect 31053 5111 31253 5127
rect 31053 5077 31069 5111
rect 31237 5077 31253 5111
rect 31053 5039 31253 5077
rect 31425 5111 31625 5127
rect 31425 5077 31441 5111
rect 31609 5077 31625 5111
rect 31425 5039 31625 5077
rect 31797 5111 31997 5127
rect 31797 5077 31813 5111
rect 31981 5077 31997 5111
rect 31797 5039 31997 5077
rect 32169 5111 32369 5127
rect 32169 5077 32185 5111
rect 32353 5077 32369 5111
rect 32169 5039 32369 5077
rect 32541 5111 32741 5127
rect 32541 5077 32557 5111
rect 32725 5077 32741 5111
rect 32541 5039 32741 5077
rect 32913 5111 33113 5127
rect 32913 5077 32929 5111
rect 33097 5077 33113 5111
rect 32913 5039 33113 5077
rect 33285 5111 33485 5127
rect 33285 5077 33301 5111
rect 33469 5077 33485 5111
rect 33285 5039 33485 5077
rect 33657 5111 33857 5127
rect 33657 5077 33673 5111
rect 33841 5077 33857 5111
rect 33657 5039 33857 5077
rect 34029 5111 34229 5127
rect 34029 5077 34045 5111
rect 34213 5077 34229 5111
rect 34029 5039 34229 5077
rect 34401 5111 34601 5127
rect 34401 5077 34417 5111
rect 34585 5077 34601 5111
rect 34401 5039 34601 5077
rect 34773 5111 34973 5127
rect 34773 5077 34789 5111
rect 34957 5077 34973 5111
rect 34773 5039 34973 5077
rect 35145 5111 35345 5127
rect 35145 5077 35161 5111
rect 35329 5077 35345 5111
rect 35145 5039 35345 5077
rect 35517 5111 35717 5127
rect 35517 5077 35533 5111
rect 35701 5077 35717 5111
rect 35517 5039 35717 5077
rect 35889 5111 36089 5127
rect 35889 5077 35905 5111
rect 36073 5077 36089 5111
rect 35889 5039 36089 5077
rect 36261 5111 36461 5127
rect 36261 5077 36277 5111
rect 36445 5077 36461 5111
rect 36261 5039 36461 5077
rect 36633 5111 36833 5127
rect 36633 5077 36649 5111
rect 36817 5077 36833 5111
rect 36633 5039 36833 5077
rect 37005 5111 37205 5127
rect 37005 5077 37021 5111
rect 37189 5077 37205 5111
rect 37005 5039 37205 5077
rect 37377 5111 37577 5127
rect 37377 5077 37393 5111
rect 37561 5077 37577 5111
rect 37377 5039 37577 5077
rect 37749 5111 37949 5127
rect 37749 5077 37765 5111
rect 37933 5077 37949 5111
rect 37749 5039 37949 5077
rect 38121 5111 38321 5127
rect 38121 5077 38137 5111
rect 38305 5077 38321 5111
rect 38121 5039 38321 5077
rect 38493 5111 38693 5127
rect 38493 5077 38509 5111
rect 38677 5077 38693 5111
rect 38493 5039 38693 5077
rect 38865 5111 39065 5127
rect 38865 5077 38881 5111
rect 39049 5077 39065 5111
rect 38865 5039 39065 5077
rect 30309 4801 30509 4839
rect 30309 4767 30325 4801
rect 30493 4767 30509 4801
rect 30309 4751 30509 4767
rect 30681 4801 30881 4839
rect 30681 4767 30697 4801
rect 30865 4767 30881 4801
rect 30681 4751 30881 4767
rect 31053 4801 31253 4839
rect 31053 4767 31069 4801
rect 31237 4767 31253 4801
rect 31053 4751 31253 4767
rect 31425 4801 31625 4839
rect 31425 4767 31441 4801
rect 31609 4767 31625 4801
rect 31425 4751 31625 4767
rect 31797 4801 31997 4839
rect 31797 4767 31813 4801
rect 31981 4767 31997 4801
rect 31797 4751 31997 4767
rect 32169 4801 32369 4839
rect 32169 4767 32185 4801
rect 32353 4767 32369 4801
rect 32169 4751 32369 4767
rect 32541 4801 32741 4839
rect 32541 4767 32557 4801
rect 32725 4767 32741 4801
rect 32541 4751 32741 4767
rect 32913 4801 33113 4839
rect 32913 4767 32929 4801
rect 33097 4767 33113 4801
rect 32913 4751 33113 4767
rect 33285 4801 33485 4839
rect 33285 4767 33301 4801
rect 33469 4767 33485 4801
rect 33285 4751 33485 4767
rect 33657 4801 33857 4839
rect 33657 4767 33673 4801
rect 33841 4767 33857 4801
rect 33657 4751 33857 4767
rect 34029 4801 34229 4839
rect 34029 4767 34045 4801
rect 34213 4767 34229 4801
rect 34029 4751 34229 4767
rect 34401 4801 34601 4839
rect 34401 4767 34417 4801
rect 34585 4767 34601 4801
rect 34401 4751 34601 4767
rect 34773 4801 34973 4839
rect 34773 4767 34789 4801
rect 34957 4767 34973 4801
rect 34773 4751 34973 4767
rect 35145 4801 35345 4839
rect 35145 4767 35161 4801
rect 35329 4767 35345 4801
rect 35145 4751 35345 4767
rect 35517 4801 35717 4839
rect 35517 4767 35533 4801
rect 35701 4767 35717 4801
rect 35517 4751 35717 4767
rect 35889 4801 36089 4839
rect 35889 4767 35905 4801
rect 36073 4767 36089 4801
rect 35889 4751 36089 4767
rect 36261 4801 36461 4839
rect 36261 4767 36277 4801
rect 36445 4767 36461 4801
rect 36261 4751 36461 4767
rect 36633 4801 36833 4839
rect 36633 4767 36649 4801
rect 36817 4767 36833 4801
rect 36633 4751 36833 4767
rect 37005 4801 37205 4839
rect 37005 4767 37021 4801
rect 37189 4767 37205 4801
rect 37005 4751 37205 4767
rect 37377 4801 37577 4839
rect 37377 4767 37393 4801
rect 37561 4767 37577 4801
rect 37377 4751 37577 4767
rect 37749 4801 37949 4839
rect 37749 4767 37765 4801
rect 37933 4767 37949 4801
rect 37749 4751 37949 4767
rect 38121 4801 38321 4839
rect 38121 4767 38137 4801
rect 38305 4767 38321 4801
rect 38121 4751 38321 4767
rect 38493 4801 38693 4839
rect 38493 4767 38509 4801
rect 38677 4767 38693 4801
rect 38493 4751 38693 4767
rect 38865 4801 39065 4839
rect 38865 4767 38881 4801
rect 39049 4767 39065 4801
rect 38865 4751 39065 4767
rect 30309 4693 30509 4709
rect 30309 4659 30325 4693
rect 30493 4659 30509 4693
rect 30309 4621 30509 4659
rect 30681 4693 30881 4709
rect 30681 4659 30697 4693
rect 30865 4659 30881 4693
rect 30681 4621 30881 4659
rect 31053 4693 31253 4709
rect 31053 4659 31069 4693
rect 31237 4659 31253 4693
rect 31053 4621 31253 4659
rect 31425 4693 31625 4709
rect 31425 4659 31441 4693
rect 31609 4659 31625 4693
rect 31425 4621 31625 4659
rect 31797 4693 31997 4709
rect 31797 4659 31813 4693
rect 31981 4659 31997 4693
rect 31797 4621 31997 4659
rect 32169 4693 32369 4709
rect 32169 4659 32185 4693
rect 32353 4659 32369 4693
rect 32169 4621 32369 4659
rect 32541 4693 32741 4709
rect 32541 4659 32557 4693
rect 32725 4659 32741 4693
rect 32541 4621 32741 4659
rect 32913 4693 33113 4709
rect 32913 4659 32929 4693
rect 33097 4659 33113 4693
rect 32913 4621 33113 4659
rect 33285 4693 33485 4709
rect 33285 4659 33301 4693
rect 33469 4659 33485 4693
rect 33285 4621 33485 4659
rect 33657 4693 33857 4709
rect 33657 4659 33673 4693
rect 33841 4659 33857 4693
rect 33657 4621 33857 4659
rect 34029 4693 34229 4709
rect 34029 4659 34045 4693
rect 34213 4659 34229 4693
rect 34029 4621 34229 4659
rect 34401 4693 34601 4709
rect 34401 4659 34417 4693
rect 34585 4659 34601 4693
rect 34401 4621 34601 4659
rect 34773 4693 34973 4709
rect 34773 4659 34789 4693
rect 34957 4659 34973 4693
rect 34773 4621 34973 4659
rect 35145 4693 35345 4709
rect 35145 4659 35161 4693
rect 35329 4659 35345 4693
rect 35145 4621 35345 4659
rect 35517 4693 35717 4709
rect 35517 4659 35533 4693
rect 35701 4659 35717 4693
rect 35517 4621 35717 4659
rect 35889 4693 36089 4709
rect 35889 4659 35905 4693
rect 36073 4659 36089 4693
rect 35889 4621 36089 4659
rect 36261 4693 36461 4709
rect 36261 4659 36277 4693
rect 36445 4659 36461 4693
rect 36261 4621 36461 4659
rect 36633 4693 36833 4709
rect 36633 4659 36649 4693
rect 36817 4659 36833 4693
rect 36633 4621 36833 4659
rect 37005 4693 37205 4709
rect 37005 4659 37021 4693
rect 37189 4659 37205 4693
rect 37005 4621 37205 4659
rect 37377 4693 37577 4709
rect 37377 4659 37393 4693
rect 37561 4659 37577 4693
rect 37377 4621 37577 4659
rect 37749 4693 37949 4709
rect 37749 4659 37765 4693
rect 37933 4659 37949 4693
rect 37749 4621 37949 4659
rect 38121 4693 38321 4709
rect 38121 4659 38137 4693
rect 38305 4659 38321 4693
rect 38121 4621 38321 4659
rect 38493 4693 38693 4709
rect 38493 4659 38509 4693
rect 38677 4659 38693 4693
rect 38493 4621 38693 4659
rect 38865 4693 39065 4709
rect 38865 4659 38881 4693
rect 39049 4659 39065 4693
rect 38865 4621 39065 4659
rect 30309 4383 30509 4421
rect 30309 4349 30325 4383
rect 30493 4349 30509 4383
rect 30309 4333 30509 4349
rect 30681 4383 30881 4421
rect 30681 4349 30697 4383
rect 30865 4349 30881 4383
rect 30681 4333 30881 4349
rect 31053 4383 31253 4421
rect 31053 4349 31069 4383
rect 31237 4349 31253 4383
rect 31053 4333 31253 4349
rect 31425 4383 31625 4421
rect 31425 4349 31441 4383
rect 31609 4349 31625 4383
rect 31425 4333 31625 4349
rect 31797 4383 31997 4421
rect 31797 4349 31813 4383
rect 31981 4349 31997 4383
rect 31797 4333 31997 4349
rect 32169 4383 32369 4421
rect 32169 4349 32185 4383
rect 32353 4349 32369 4383
rect 32169 4333 32369 4349
rect 32541 4383 32741 4421
rect 32541 4349 32557 4383
rect 32725 4349 32741 4383
rect 32541 4333 32741 4349
rect 32913 4383 33113 4421
rect 32913 4349 32929 4383
rect 33097 4349 33113 4383
rect 32913 4333 33113 4349
rect 33285 4383 33485 4421
rect 33285 4349 33301 4383
rect 33469 4349 33485 4383
rect 33285 4333 33485 4349
rect 33657 4383 33857 4421
rect 33657 4349 33673 4383
rect 33841 4349 33857 4383
rect 33657 4333 33857 4349
rect 34029 4383 34229 4421
rect 34029 4349 34045 4383
rect 34213 4349 34229 4383
rect 34029 4333 34229 4349
rect 34401 4383 34601 4421
rect 34401 4349 34417 4383
rect 34585 4349 34601 4383
rect 34401 4333 34601 4349
rect 34773 4383 34973 4421
rect 34773 4349 34789 4383
rect 34957 4349 34973 4383
rect 34773 4333 34973 4349
rect 35145 4383 35345 4421
rect 35145 4349 35161 4383
rect 35329 4349 35345 4383
rect 35145 4333 35345 4349
rect 35517 4383 35717 4421
rect 35517 4349 35533 4383
rect 35701 4349 35717 4383
rect 35517 4333 35717 4349
rect 35889 4383 36089 4421
rect 35889 4349 35905 4383
rect 36073 4349 36089 4383
rect 35889 4333 36089 4349
rect 36261 4383 36461 4421
rect 36261 4349 36277 4383
rect 36445 4349 36461 4383
rect 36261 4333 36461 4349
rect 36633 4383 36833 4421
rect 36633 4349 36649 4383
rect 36817 4349 36833 4383
rect 36633 4333 36833 4349
rect 37005 4383 37205 4421
rect 37005 4349 37021 4383
rect 37189 4349 37205 4383
rect 37005 4333 37205 4349
rect 37377 4383 37577 4421
rect 37377 4349 37393 4383
rect 37561 4349 37577 4383
rect 37377 4333 37577 4349
rect 37749 4383 37949 4421
rect 37749 4349 37765 4383
rect 37933 4349 37949 4383
rect 37749 4333 37949 4349
rect 38121 4383 38321 4421
rect 38121 4349 38137 4383
rect 38305 4349 38321 4383
rect 38121 4333 38321 4349
rect 38493 4383 38693 4421
rect 38493 4349 38509 4383
rect 38677 4349 38693 4383
rect 38493 4333 38693 4349
rect 38865 4383 39065 4421
rect 38865 4349 38881 4383
rect 39049 4349 39065 4383
rect 38865 4333 39065 4349
rect 30309 4275 30509 4291
rect 30309 4241 30325 4275
rect 30493 4241 30509 4275
rect 30309 4203 30509 4241
rect 30681 4275 30881 4291
rect 30681 4241 30697 4275
rect 30865 4241 30881 4275
rect 30681 4203 30881 4241
rect 31053 4275 31253 4291
rect 31053 4241 31069 4275
rect 31237 4241 31253 4275
rect 31053 4203 31253 4241
rect 31425 4275 31625 4291
rect 31425 4241 31441 4275
rect 31609 4241 31625 4275
rect 31425 4203 31625 4241
rect 31797 4275 31997 4291
rect 31797 4241 31813 4275
rect 31981 4241 31997 4275
rect 31797 4203 31997 4241
rect 32169 4275 32369 4291
rect 32169 4241 32185 4275
rect 32353 4241 32369 4275
rect 32169 4203 32369 4241
rect 32541 4275 32741 4291
rect 32541 4241 32557 4275
rect 32725 4241 32741 4275
rect 32541 4203 32741 4241
rect 32913 4275 33113 4291
rect 32913 4241 32929 4275
rect 33097 4241 33113 4275
rect 32913 4203 33113 4241
rect 33285 4275 33485 4291
rect 33285 4241 33301 4275
rect 33469 4241 33485 4275
rect 33285 4203 33485 4241
rect 33657 4275 33857 4291
rect 33657 4241 33673 4275
rect 33841 4241 33857 4275
rect 33657 4203 33857 4241
rect 34029 4275 34229 4291
rect 34029 4241 34045 4275
rect 34213 4241 34229 4275
rect 34029 4203 34229 4241
rect 34401 4275 34601 4291
rect 34401 4241 34417 4275
rect 34585 4241 34601 4275
rect 34401 4203 34601 4241
rect 34773 4275 34973 4291
rect 34773 4241 34789 4275
rect 34957 4241 34973 4275
rect 34773 4203 34973 4241
rect 35145 4275 35345 4291
rect 35145 4241 35161 4275
rect 35329 4241 35345 4275
rect 35145 4203 35345 4241
rect 35517 4275 35717 4291
rect 35517 4241 35533 4275
rect 35701 4241 35717 4275
rect 35517 4203 35717 4241
rect 35889 4275 36089 4291
rect 35889 4241 35905 4275
rect 36073 4241 36089 4275
rect 35889 4203 36089 4241
rect 36261 4275 36461 4291
rect 36261 4241 36277 4275
rect 36445 4241 36461 4275
rect 36261 4203 36461 4241
rect 36633 4275 36833 4291
rect 36633 4241 36649 4275
rect 36817 4241 36833 4275
rect 36633 4203 36833 4241
rect 37005 4275 37205 4291
rect 37005 4241 37021 4275
rect 37189 4241 37205 4275
rect 37005 4203 37205 4241
rect 37377 4275 37577 4291
rect 37377 4241 37393 4275
rect 37561 4241 37577 4275
rect 37377 4203 37577 4241
rect 37749 4275 37949 4291
rect 37749 4241 37765 4275
rect 37933 4241 37949 4275
rect 37749 4203 37949 4241
rect 38121 4275 38321 4291
rect 38121 4241 38137 4275
rect 38305 4241 38321 4275
rect 38121 4203 38321 4241
rect 38493 4275 38693 4291
rect 38493 4241 38509 4275
rect 38677 4241 38693 4275
rect 38493 4203 38693 4241
rect 38865 4275 39065 4291
rect 38865 4241 38881 4275
rect 39049 4241 39065 4275
rect 38865 4203 39065 4241
rect 30309 3965 30509 4003
rect 30309 3931 30325 3965
rect 30493 3931 30509 3965
rect 30309 3915 30509 3931
rect 30681 3965 30881 4003
rect 30681 3931 30697 3965
rect 30865 3931 30881 3965
rect 30681 3915 30881 3931
rect 31053 3965 31253 4003
rect 31053 3931 31069 3965
rect 31237 3931 31253 3965
rect 31053 3915 31253 3931
rect 31425 3965 31625 4003
rect 31425 3931 31441 3965
rect 31609 3931 31625 3965
rect 31425 3915 31625 3931
rect 31797 3965 31997 4003
rect 31797 3931 31813 3965
rect 31981 3931 31997 3965
rect 31797 3915 31997 3931
rect 32169 3965 32369 4003
rect 32169 3931 32185 3965
rect 32353 3931 32369 3965
rect 32169 3915 32369 3931
rect 32541 3965 32741 4003
rect 32541 3931 32557 3965
rect 32725 3931 32741 3965
rect 32541 3915 32741 3931
rect 32913 3965 33113 4003
rect 32913 3931 32929 3965
rect 33097 3931 33113 3965
rect 32913 3915 33113 3931
rect 33285 3965 33485 4003
rect 33285 3931 33301 3965
rect 33469 3931 33485 3965
rect 33285 3915 33485 3931
rect 33657 3965 33857 4003
rect 33657 3931 33673 3965
rect 33841 3931 33857 3965
rect 33657 3915 33857 3931
rect 34029 3965 34229 4003
rect 34029 3931 34045 3965
rect 34213 3931 34229 3965
rect 34029 3915 34229 3931
rect 34401 3965 34601 4003
rect 34401 3931 34417 3965
rect 34585 3931 34601 3965
rect 34401 3915 34601 3931
rect 34773 3965 34973 4003
rect 34773 3931 34789 3965
rect 34957 3931 34973 3965
rect 34773 3915 34973 3931
rect 35145 3965 35345 4003
rect 35145 3931 35161 3965
rect 35329 3931 35345 3965
rect 35145 3915 35345 3931
rect 35517 3965 35717 4003
rect 35517 3931 35533 3965
rect 35701 3931 35717 3965
rect 35517 3915 35717 3931
rect 35889 3965 36089 4003
rect 35889 3931 35905 3965
rect 36073 3931 36089 3965
rect 35889 3915 36089 3931
rect 36261 3965 36461 4003
rect 36261 3931 36277 3965
rect 36445 3931 36461 3965
rect 36261 3915 36461 3931
rect 36633 3965 36833 4003
rect 36633 3931 36649 3965
rect 36817 3931 36833 3965
rect 36633 3915 36833 3931
rect 37005 3965 37205 4003
rect 37005 3931 37021 3965
rect 37189 3931 37205 3965
rect 37005 3915 37205 3931
rect 37377 3965 37577 4003
rect 37377 3931 37393 3965
rect 37561 3931 37577 3965
rect 37377 3915 37577 3931
rect 37749 3965 37949 4003
rect 37749 3931 37765 3965
rect 37933 3931 37949 3965
rect 37749 3915 37949 3931
rect 38121 3965 38321 4003
rect 38121 3931 38137 3965
rect 38305 3931 38321 3965
rect 38121 3915 38321 3931
rect 38493 3965 38693 4003
rect 38493 3931 38509 3965
rect 38677 3931 38693 3965
rect 38493 3915 38693 3931
rect 38865 3965 39065 4003
rect 38865 3931 38881 3965
rect 39049 3931 39065 3965
rect 38865 3915 39065 3931
rect 30309 3857 30509 3873
rect 30309 3823 30325 3857
rect 30493 3823 30509 3857
rect 30309 3785 30509 3823
rect 30681 3857 30881 3873
rect 30681 3823 30697 3857
rect 30865 3823 30881 3857
rect 30681 3785 30881 3823
rect 31053 3857 31253 3873
rect 31053 3823 31069 3857
rect 31237 3823 31253 3857
rect 31053 3785 31253 3823
rect 31425 3857 31625 3873
rect 31425 3823 31441 3857
rect 31609 3823 31625 3857
rect 31425 3785 31625 3823
rect 31797 3857 31997 3873
rect 31797 3823 31813 3857
rect 31981 3823 31997 3857
rect 31797 3785 31997 3823
rect 32169 3857 32369 3873
rect 32169 3823 32185 3857
rect 32353 3823 32369 3857
rect 32169 3785 32369 3823
rect 32541 3857 32741 3873
rect 32541 3823 32557 3857
rect 32725 3823 32741 3857
rect 32541 3785 32741 3823
rect 32913 3857 33113 3873
rect 32913 3823 32929 3857
rect 33097 3823 33113 3857
rect 32913 3785 33113 3823
rect 33285 3857 33485 3873
rect 33285 3823 33301 3857
rect 33469 3823 33485 3857
rect 33285 3785 33485 3823
rect 33657 3857 33857 3873
rect 33657 3823 33673 3857
rect 33841 3823 33857 3857
rect 33657 3785 33857 3823
rect 34029 3857 34229 3873
rect 34029 3823 34045 3857
rect 34213 3823 34229 3857
rect 34029 3785 34229 3823
rect 34401 3857 34601 3873
rect 34401 3823 34417 3857
rect 34585 3823 34601 3857
rect 34401 3785 34601 3823
rect 34773 3857 34973 3873
rect 34773 3823 34789 3857
rect 34957 3823 34973 3857
rect 34773 3785 34973 3823
rect 35145 3857 35345 3873
rect 35145 3823 35161 3857
rect 35329 3823 35345 3857
rect 35145 3785 35345 3823
rect 35517 3857 35717 3873
rect 35517 3823 35533 3857
rect 35701 3823 35717 3857
rect 35517 3785 35717 3823
rect 35889 3857 36089 3873
rect 35889 3823 35905 3857
rect 36073 3823 36089 3857
rect 35889 3785 36089 3823
rect 36261 3857 36461 3873
rect 36261 3823 36277 3857
rect 36445 3823 36461 3857
rect 36261 3785 36461 3823
rect 36633 3857 36833 3873
rect 36633 3823 36649 3857
rect 36817 3823 36833 3857
rect 36633 3785 36833 3823
rect 37005 3857 37205 3873
rect 37005 3823 37021 3857
rect 37189 3823 37205 3857
rect 37005 3785 37205 3823
rect 37377 3857 37577 3873
rect 37377 3823 37393 3857
rect 37561 3823 37577 3857
rect 37377 3785 37577 3823
rect 37749 3857 37949 3873
rect 37749 3823 37765 3857
rect 37933 3823 37949 3857
rect 37749 3785 37949 3823
rect 38121 3857 38321 3873
rect 38121 3823 38137 3857
rect 38305 3823 38321 3857
rect 38121 3785 38321 3823
rect 38493 3857 38693 3873
rect 38493 3823 38509 3857
rect 38677 3823 38693 3857
rect 38493 3785 38693 3823
rect 38865 3857 39065 3873
rect 38865 3823 38881 3857
rect 39049 3823 39065 3857
rect 38865 3785 39065 3823
rect 30309 3547 30509 3585
rect 30309 3513 30325 3547
rect 30493 3513 30509 3547
rect 30309 3497 30509 3513
rect 30681 3547 30881 3585
rect 30681 3513 30697 3547
rect 30865 3513 30881 3547
rect 30681 3497 30881 3513
rect 31053 3547 31253 3585
rect 31053 3513 31069 3547
rect 31237 3513 31253 3547
rect 31053 3497 31253 3513
rect 31425 3547 31625 3585
rect 31425 3513 31441 3547
rect 31609 3513 31625 3547
rect 31425 3497 31625 3513
rect 31797 3547 31997 3585
rect 31797 3513 31813 3547
rect 31981 3513 31997 3547
rect 31797 3497 31997 3513
rect 32169 3547 32369 3585
rect 32169 3513 32185 3547
rect 32353 3513 32369 3547
rect 32169 3497 32369 3513
rect 32541 3547 32741 3585
rect 32541 3513 32557 3547
rect 32725 3513 32741 3547
rect 32541 3497 32741 3513
rect 32913 3547 33113 3585
rect 32913 3513 32929 3547
rect 33097 3513 33113 3547
rect 32913 3497 33113 3513
rect 33285 3547 33485 3585
rect 33285 3513 33301 3547
rect 33469 3513 33485 3547
rect 33285 3497 33485 3513
rect 33657 3547 33857 3585
rect 33657 3513 33673 3547
rect 33841 3513 33857 3547
rect 33657 3497 33857 3513
rect 34029 3547 34229 3585
rect 34029 3513 34045 3547
rect 34213 3513 34229 3547
rect 34029 3497 34229 3513
rect 34401 3547 34601 3585
rect 34401 3513 34417 3547
rect 34585 3513 34601 3547
rect 34401 3497 34601 3513
rect 34773 3547 34973 3585
rect 34773 3513 34789 3547
rect 34957 3513 34973 3547
rect 34773 3497 34973 3513
rect 35145 3547 35345 3585
rect 35145 3513 35161 3547
rect 35329 3513 35345 3547
rect 35145 3497 35345 3513
rect 35517 3547 35717 3585
rect 35517 3513 35533 3547
rect 35701 3513 35717 3547
rect 35517 3497 35717 3513
rect 35889 3547 36089 3585
rect 35889 3513 35905 3547
rect 36073 3513 36089 3547
rect 35889 3497 36089 3513
rect 36261 3547 36461 3585
rect 36261 3513 36277 3547
rect 36445 3513 36461 3547
rect 36261 3497 36461 3513
rect 36633 3547 36833 3585
rect 36633 3513 36649 3547
rect 36817 3513 36833 3547
rect 36633 3497 36833 3513
rect 37005 3547 37205 3585
rect 37005 3513 37021 3547
rect 37189 3513 37205 3547
rect 37005 3497 37205 3513
rect 37377 3547 37577 3585
rect 37377 3513 37393 3547
rect 37561 3513 37577 3547
rect 37377 3497 37577 3513
rect 37749 3547 37949 3585
rect 37749 3513 37765 3547
rect 37933 3513 37949 3547
rect 37749 3497 37949 3513
rect 38121 3547 38321 3585
rect 38121 3513 38137 3547
rect 38305 3513 38321 3547
rect 38121 3497 38321 3513
rect 38493 3547 38693 3585
rect 38493 3513 38509 3547
rect 38677 3513 38693 3547
rect 38493 3497 38693 3513
rect 38865 3547 39065 3585
rect 38865 3513 38881 3547
rect 39049 3513 39065 3547
rect 38865 3497 39065 3513
<< polycont >>
rect 28837 12159 29005 12193
rect 29209 12159 29377 12193
rect 29581 12159 29749 12193
rect 29953 12159 30121 12193
rect 30325 12159 30493 12193
rect 30697 12159 30865 12193
rect 31069 12159 31237 12193
rect 31441 12159 31609 12193
rect 31813 12159 31981 12193
rect 32185 12159 32353 12193
rect 32557 12159 32725 12193
rect 32929 12159 33097 12193
rect 33301 12159 33469 12193
rect 33673 12159 33841 12193
rect 34045 12159 34213 12193
rect 34417 12159 34585 12193
rect 34789 12159 34957 12193
rect 35161 12159 35329 12193
rect 35533 12159 35701 12193
rect 35905 12159 36073 12193
rect 36277 12159 36445 12193
rect 36649 12159 36817 12193
rect 37021 12159 37189 12193
rect 37393 12159 37561 12193
rect 37765 12159 37933 12193
rect 38137 12159 38305 12193
rect 38509 12159 38677 12193
rect 38881 12159 39049 12193
rect 39253 12159 39421 12193
rect 39625 12159 39793 12193
rect 39997 12159 40165 12193
rect 40369 12159 40537 12193
rect 28837 11631 29005 11665
rect 29209 11631 29377 11665
rect 29581 11631 29749 11665
rect 29953 11631 30121 11665
rect 30325 11631 30493 11665
rect 30697 11631 30865 11665
rect 31069 11631 31237 11665
rect 31441 11631 31609 11665
rect 31813 11631 31981 11665
rect 32185 11631 32353 11665
rect 32557 11631 32725 11665
rect 32929 11631 33097 11665
rect 33301 11631 33469 11665
rect 33673 11631 33841 11665
rect 34045 11631 34213 11665
rect 34417 11631 34585 11665
rect 34789 11631 34957 11665
rect 35161 11631 35329 11665
rect 35533 11631 35701 11665
rect 35905 11631 36073 11665
rect 36277 11631 36445 11665
rect 36649 11631 36817 11665
rect 37021 11631 37189 11665
rect 37393 11631 37561 11665
rect 37765 11631 37933 11665
rect 38137 11631 38305 11665
rect 38509 11631 38677 11665
rect 38881 11631 39049 11665
rect 39253 11631 39421 11665
rect 39625 11631 39793 11665
rect 39997 11631 40165 11665
rect 40369 11631 40537 11665
rect 28837 11523 29005 11557
rect 29209 11523 29377 11557
rect 29581 11523 29749 11557
rect 29953 11523 30121 11557
rect 30325 11523 30493 11557
rect 30697 11523 30865 11557
rect 31069 11523 31237 11557
rect 31441 11523 31609 11557
rect 31813 11523 31981 11557
rect 32185 11523 32353 11557
rect 32557 11523 32725 11557
rect 32929 11523 33097 11557
rect 33301 11523 33469 11557
rect 33673 11523 33841 11557
rect 34045 11523 34213 11557
rect 34417 11523 34585 11557
rect 34789 11523 34957 11557
rect 35161 11523 35329 11557
rect 35533 11523 35701 11557
rect 35905 11523 36073 11557
rect 36277 11523 36445 11557
rect 36649 11523 36817 11557
rect 37021 11523 37189 11557
rect 37393 11523 37561 11557
rect 37765 11523 37933 11557
rect 38137 11523 38305 11557
rect 38509 11523 38677 11557
rect 38881 11523 39049 11557
rect 39253 11523 39421 11557
rect 39625 11523 39793 11557
rect 39997 11523 40165 11557
rect 40369 11523 40537 11557
rect 28837 10995 29005 11029
rect 29209 10995 29377 11029
rect 29581 10995 29749 11029
rect 29953 10995 30121 11029
rect 30325 10995 30493 11029
rect 30697 10995 30865 11029
rect 31069 10995 31237 11029
rect 31441 10995 31609 11029
rect 31813 10995 31981 11029
rect 32185 10995 32353 11029
rect 32557 10995 32725 11029
rect 32929 10995 33097 11029
rect 33301 10995 33469 11029
rect 33673 10995 33841 11029
rect 34045 10995 34213 11029
rect 34417 10995 34585 11029
rect 34789 10995 34957 11029
rect 35161 10995 35329 11029
rect 35533 10995 35701 11029
rect 35905 10995 36073 11029
rect 36277 10995 36445 11029
rect 36649 10995 36817 11029
rect 37021 10995 37189 11029
rect 37393 10995 37561 11029
rect 37765 10995 37933 11029
rect 38137 10995 38305 11029
rect 38509 10995 38677 11029
rect 38881 10995 39049 11029
rect 39253 10995 39421 11029
rect 39625 10995 39793 11029
rect 39997 10995 40165 11029
rect 40369 10995 40537 11029
rect 28837 10887 29005 10921
rect 29209 10887 29377 10921
rect 29581 10887 29749 10921
rect 29953 10887 30121 10921
rect 30325 10887 30493 10921
rect 30697 10887 30865 10921
rect 31069 10887 31237 10921
rect 31441 10887 31609 10921
rect 31813 10887 31981 10921
rect 32185 10887 32353 10921
rect 32557 10887 32725 10921
rect 32929 10887 33097 10921
rect 33301 10887 33469 10921
rect 33673 10887 33841 10921
rect 34045 10887 34213 10921
rect 34417 10887 34585 10921
rect 34789 10887 34957 10921
rect 35161 10887 35329 10921
rect 35533 10887 35701 10921
rect 35905 10887 36073 10921
rect 36277 10887 36445 10921
rect 36649 10887 36817 10921
rect 37021 10887 37189 10921
rect 37393 10887 37561 10921
rect 37765 10887 37933 10921
rect 38137 10887 38305 10921
rect 38509 10887 38677 10921
rect 38881 10887 39049 10921
rect 39253 10887 39421 10921
rect 39625 10887 39793 10921
rect 39997 10887 40165 10921
rect 40369 10887 40537 10921
rect 28837 10359 29005 10393
rect 29209 10359 29377 10393
rect 29581 10359 29749 10393
rect 29953 10359 30121 10393
rect 30325 10359 30493 10393
rect 30697 10359 30865 10393
rect 31069 10359 31237 10393
rect 31441 10359 31609 10393
rect 31813 10359 31981 10393
rect 32185 10359 32353 10393
rect 32557 10359 32725 10393
rect 32929 10359 33097 10393
rect 33301 10359 33469 10393
rect 33673 10359 33841 10393
rect 34045 10359 34213 10393
rect 34417 10359 34585 10393
rect 34789 10359 34957 10393
rect 35161 10359 35329 10393
rect 35533 10359 35701 10393
rect 35905 10359 36073 10393
rect 36277 10359 36445 10393
rect 36649 10359 36817 10393
rect 37021 10359 37189 10393
rect 37393 10359 37561 10393
rect 37765 10359 37933 10393
rect 38137 10359 38305 10393
rect 38509 10359 38677 10393
rect 38881 10359 39049 10393
rect 39253 10359 39421 10393
rect 39625 10359 39793 10393
rect 39997 10359 40165 10393
rect 40369 10359 40537 10393
rect 30325 9771 30493 9805
rect 30697 9771 30865 9805
rect 31069 9771 31237 9805
rect 31441 9771 31609 9805
rect 31813 9771 31981 9805
rect 32185 9771 32353 9805
rect 32557 9771 32725 9805
rect 32929 9771 33097 9805
rect 30325 8843 30493 8877
rect 30697 8843 30865 8877
rect 31069 8843 31237 8877
rect 31441 8843 31609 8877
rect 31813 8843 31981 8877
rect 32185 8843 32353 8877
rect 32557 8843 32725 8877
rect 32929 8843 33097 8877
rect 30325 8735 30493 8769
rect 30697 8735 30865 8769
rect 31069 8735 31237 8769
rect 31441 8735 31609 8769
rect 31813 8735 31981 8769
rect 32185 8735 32353 8769
rect 32557 8735 32725 8769
rect 32929 8735 33097 8769
rect 30325 7807 30493 7841
rect 30697 7807 30865 7841
rect 31069 7807 31237 7841
rect 31441 7807 31609 7841
rect 31813 7807 31981 7841
rect 32185 7807 32353 7841
rect 32557 7807 32725 7841
rect 32929 7807 33097 7841
rect 30325 7699 30493 7733
rect 30697 7699 30865 7733
rect 31069 7699 31237 7733
rect 31441 7699 31609 7733
rect 31813 7699 31981 7733
rect 32185 7699 32353 7733
rect 32557 7699 32725 7733
rect 32929 7699 33097 7733
rect 30325 6771 30493 6805
rect 30697 6771 30865 6805
rect 31069 6771 31237 6805
rect 31441 6771 31609 6805
rect 31813 6771 31981 6805
rect 32185 6771 32353 6805
rect 32557 6771 32725 6805
rect 32929 6771 33097 6805
rect 30325 6663 30493 6697
rect 30697 6663 30865 6697
rect 31069 6663 31237 6697
rect 31441 6663 31609 6697
rect 31813 6663 31981 6697
rect 32185 6663 32353 6697
rect 32557 6663 32725 6697
rect 32929 6663 33097 6697
rect 30325 5735 30493 5769
rect 30697 5735 30865 5769
rect 31069 5735 31237 5769
rect 31441 5735 31609 5769
rect 31813 5735 31981 5769
rect 32185 5735 32353 5769
rect 32557 5735 32725 5769
rect 32929 5735 33097 5769
rect 30325 5077 30493 5111
rect 30697 5077 30865 5111
rect 31069 5077 31237 5111
rect 31441 5077 31609 5111
rect 31813 5077 31981 5111
rect 32185 5077 32353 5111
rect 32557 5077 32725 5111
rect 32929 5077 33097 5111
rect 33301 5077 33469 5111
rect 33673 5077 33841 5111
rect 34045 5077 34213 5111
rect 34417 5077 34585 5111
rect 34789 5077 34957 5111
rect 35161 5077 35329 5111
rect 35533 5077 35701 5111
rect 35905 5077 36073 5111
rect 36277 5077 36445 5111
rect 36649 5077 36817 5111
rect 37021 5077 37189 5111
rect 37393 5077 37561 5111
rect 37765 5077 37933 5111
rect 38137 5077 38305 5111
rect 38509 5077 38677 5111
rect 38881 5077 39049 5111
rect 30325 4767 30493 4801
rect 30697 4767 30865 4801
rect 31069 4767 31237 4801
rect 31441 4767 31609 4801
rect 31813 4767 31981 4801
rect 32185 4767 32353 4801
rect 32557 4767 32725 4801
rect 32929 4767 33097 4801
rect 33301 4767 33469 4801
rect 33673 4767 33841 4801
rect 34045 4767 34213 4801
rect 34417 4767 34585 4801
rect 34789 4767 34957 4801
rect 35161 4767 35329 4801
rect 35533 4767 35701 4801
rect 35905 4767 36073 4801
rect 36277 4767 36445 4801
rect 36649 4767 36817 4801
rect 37021 4767 37189 4801
rect 37393 4767 37561 4801
rect 37765 4767 37933 4801
rect 38137 4767 38305 4801
rect 38509 4767 38677 4801
rect 38881 4767 39049 4801
rect 30325 4659 30493 4693
rect 30697 4659 30865 4693
rect 31069 4659 31237 4693
rect 31441 4659 31609 4693
rect 31813 4659 31981 4693
rect 32185 4659 32353 4693
rect 32557 4659 32725 4693
rect 32929 4659 33097 4693
rect 33301 4659 33469 4693
rect 33673 4659 33841 4693
rect 34045 4659 34213 4693
rect 34417 4659 34585 4693
rect 34789 4659 34957 4693
rect 35161 4659 35329 4693
rect 35533 4659 35701 4693
rect 35905 4659 36073 4693
rect 36277 4659 36445 4693
rect 36649 4659 36817 4693
rect 37021 4659 37189 4693
rect 37393 4659 37561 4693
rect 37765 4659 37933 4693
rect 38137 4659 38305 4693
rect 38509 4659 38677 4693
rect 38881 4659 39049 4693
rect 30325 4349 30493 4383
rect 30697 4349 30865 4383
rect 31069 4349 31237 4383
rect 31441 4349 31609 4383
rect 31813 4349 31981 4383
rect 32185 4349 32353 4383
rect 32557 4349 32725 4383
rect 32929 4349 33097 4383
rect 33301 4349 33469 4383
rect 33673 4349 33841 4383
rect 34045 4349 34213 4383
rect 34417 4349 34585 4383
rect 34789 4349 34957 4383
rect 35161 4349 35329 4383
rect 35533 4349 35701 4383
rect 35905 4349 36073 4383
rect 36277 4349 36445 4383
rect 36649 4349 36817 4383
rect 37021 4349 37189 4383
rect 37393 4349 37561 4383
rect 37765 4349 37933 4383
rect 38137 4349 38305 4383
rect 38509 4349 38677 4383
rect 38881 4349 39049 4383
rect 30325 4241 30493 4275
rect 30697 4241 30865 4275
rect 31069 4241 31237 4275
rect 31441 4241 31609 4275
rect 31813 4241 31981 4275
rect 32185 4241 32353 4275
rect 32557 4241 32725 4275
rect 32929 4241 33097 4275
rect 33301 4241 33469 4275
rect 33673 4241 33841 4275
rect 34045 4241 34213 4275
rect 34417 4241 34585 4275
rect 34789 4241 34957 4275
rect 35161 4241 35329 4275
rect 35533 4241 35701 4275
rect 35905 4241 36073 4275
rect 36277 4241 36445 4275
rect 36649 4241 36817 4275
rect 37021 4241 37189 4275
rect 37393 4241 37561 4275
rect 37765 4241 37933 4275
rect 38137 4241 38305 4275
rect 38509 4241 38677 4275
rect 38881 4241 39049 4275
rect 30325 3931 30493 3965
rect 30697 3931 30865 3965
rect 31069 3931 31237 3965
rect 31441 3931 31609 3965
rect 31813 3931 31981 3965
rect 32185 3931 32353 3965
rect 32557 3931 32725 3965
rect 32929 3931 33097 3965
rect 33301 3931 33469 3965
rect 33673 3931 33841 3965
rect 34045 3931 34213 3965
rect 34417 3931 34585 3965
rect 34789 3931 34957 3965
rect 35161 3931 35329 3965
rect 35533 3931 35701 3965
rect 35905 3931 36073 3965
rect 36277 3931 36445 3965
rect 36649 3931 36817 3965
rect 37021 3931 37189 3965
rect 37393 3931 37561 3965
rect 37765 3931 37933 3965
rect 38137 3931 38305 3965
rect 38509 3931 38677 3965
rect 38881 3931 39049 3965
rect 30325 3823 30493 3857
rect 30697 3823 30865 3857
rect 31069 3823 31237 3857
rect 31441 3823 31609 3857
rect 31813 3823 31981 3857
rect 32185 3823 32353 3857
rect 32557 3823 32725 3857
rect 32929 3823 33097 3857
rect 33301 3823 33469 3857
rect 33673 3823 33841 3857
rect 34045 3823 34213 3857
rect 34417 3823 34585 3857
rect 34789 3823 34957 3857
rect 35161 3823 35329 3857
rect 35533 3823 35701 3857
rect 35905 3823 36073 3857
rect 36277 3823 36445 3857
rect 36649 3823 36817 3857
rect 37021 3823 37189 3857
rect 37393 3823 37561 3857
rect 37765 3823 37933 3857
rect 38137 3823 38305 3857
rect 38509 3823 38677 3857
rect 38881 3823 39049 3857
rect 30325 3513 30493 3547
rect 30697 3513 30865 3547
rect 31069 3513 31237 3547
rect 31441 3513 31609 3547
rect 31813 3513 31981 3547
rect 32185 3513 32353 3547
rect 32557 3513 32725 3547
rect 32929 3513 33097 3547
rect 33301 3513 33469 3547
rect 33673 3513 33841 3547
rect 34045 3513 34213 3547
rect 34417 3513 34585 3547
rect 34789 3513 34957 3547
rect 35161 3513 35329 3547
rect 35533 3513 35701 3547
rect 35905 3513 36073 3547
rect 36277 3513 36445 3547
rect 36649 3513 36817 3547
rect 37021 3513 37189 3547
rect 37393 3513 37561 3547
rect 37765 3513 37933 3547
rect 38137 3513 38305 3547
rect 38509 3513 38677 3547
rect 38881 3513 39049 3547
<< xpolycontact >>
rect 33906 7046 33976 7478
rect 33906 6334 33976 6766
<< xpolyres >>
rect 33906 6766 33976 7046
<< locali >>
rect 28661 12261 28757 12295
rect 40620 12261 40713 12295
rect 28661 12199 28695 12261
rect 40679 12199 40713 12261
rect 28821 12159 28837 12193
rect 29005 12159 29021 12193
rect 29193 12159 29209 12193
rect 29377 12159 29393 12193
rect 29565 12159 29581 12193
rect 29749 12159 29765 12193
rect 29937 12159 29953 12193
rect 30121 12159 30137 12193
rect 30309 12159 30325 12193
rect 30493 12159 30509 12193
rect 30681 12159 30697 12193
rect 30865 12159 30881 12193
rect 31053 12159 31069 12193
rect 31237 12159 31253 12193
rect 31425 12159 31441 12193
rect 31609 12159 31625 12193
rect 31797 12159 31813 12193
rect 31981 12159 31997 12193
rect 32169 12159 32185 12193
rect 32353 12159 32369 12193
rect 32541 12159 32557 12193
rect 32725 12159 32741 12193
rect 32913 12159 32929 12193
rect 33097 12159 33113 12193
rect 33285 12159 33301 12193
rect 33469 12159 33485 12193
rect 33657 12159 33673 12193
rect 33841 12159 33857 12193
rect 34029 12159 34045 12193
rect 34213 12159 34229 12193
rect 34401 12159 34417 12193
rect 34585 12159 34601 12193
rect 34773 12159 34789 12193
rect 34957 12159 34973 12193
rect 35145 12159 35161 12193
rect 35329 12159 35345 12193
rect 35517 12159 35533 12193
rect 35701 12159 35717 12193
rect 35889 12159 35905 12193
rect 36073 12159 36089 12193
rect 36261 12159 36277 12193
rect 36445 12159 36461 12193
rect 36633 12159 36649 12193
rect 36817 12159 36833 12193
rect 37005 12159 37021 12193
rect 37189 12159 37205 12193
rect 37377 12159 37393 12193
rect 37561 12159 37577 12193
rect 37749 12159 37765 12193
rect 37933 12159 37949 12193
rect 38121 12159 38137 12193
rect 38305 12159 38321 12193
rect 38493 12159 38509 12193
rect 38677 12159 38693 12193
rect 38865 12159 38881 12193
rect 39049 12159 39065 12193
rect 39237 12159 39253 12193
rect 39421 12159 39437 12193
rect 39609 12159 39625 12193
rect 39793 12159 39809 12193
rect 39981 12159 39997 12193
rect 40165 12159 40181 12193
rect 40353 12159 40369 12193
rect 40537 12159 40553 12193
rect 28775 12100 28809 12116
rect 28775 11708 28809 11724
rect 29033 12100 29067 12116
rect 29033 11708 29067 11724
rect 29147 12100 29181 12116
rect 29147 11708 29181 11724
rect 29405 12100 29439 12116
rect 29405 11708 29439 11724
rect 29519 12100 29553 12116
rect 29519 11708 29553 11724
rect 29777 12100 29811 12116
rect 29777 11708 29811 11724
rect 29891 12100 29925 12116
rect 29891 11708 29925 11724
rect 30149 12100 30183 12116
rect 30149 11708 30183 11724
rect 30263 12100 30297 12116
rect 30263 11708 30297 11724
rect 30521 12100 30555 12116
rect 30521 11708 30555 11724
rect 30635 12100 30669 12116
rect 30635 11708 30669 11724
rect 30893 12100 30927 12116
rect 30893 11708 30927 11724
rect 31007 12100 31041 12116
rect 31007 11708 31041 11724
rect 31265 12100 31299 12116
rect 31265 11708 31299 11724
rect 31379 12100 31413 12116
rect 31379 11708 31413 11724
rect 31637 12100 31671 12116
rect 31637 11708 31671 11724
rect 31751 12100 31785 12116
rect 31751 11708 31785 11724
rect 32009 12100 32043 12116
rect 32009 11708 32043 11724
rect 32123 12100 32157 12116
rect 32123 11708 32157 11724
rect 32381 12100 32415 12116
rect 32381 11708 32415 11724
rect 32495 12100 32529 12116
rect 32495 11708 32529 11724
rect 32753 12100 32787 12116
rect 32753 11708 32787 11724
rect 32867 12100 32901 12116
rect 32867 11708 32901 11724
rect 33125 12100 33159 12116
rect 33125 11708 33159 11724
rect 33239 12100 33273 12116
rect 33239 11708 33273 11724
rect 33497 12100 33531 12116
rect 33497 11708 33531 11724
rect 33611 12100 33645 12116
rect 33611 11708 33645 11724
rect 33869 12100 33903 12116
rect 33869 11708 33903 11724
rect 33983 12100 34017 12116
rect 33983 11708 34017 11724
rect 34241 12100 34275 12116
rect 34241 11708 34275 11724
rect 34355 12100 34389 12116
rect 34355 11708 34389 11724
rect 34613 12100 34647 12116
rect 34613 11708 34647 11724
rect 34727 12100 34761 12116
rect 34727 11708 34761 11724
rect 34985 12100 35019 12116
rect 34985 11708 35019 11724
rect 35099 12100 35133 12116
rect 35099 11708 35133 11724
rect 35357 12100 35391 12116
rect 35357 11708 35391 11724
rect 35471 12100 35505 12116
rect 35471 11708 35505 11724
rect 35729 12100 35763 12116
rect 35729 11708 35763 11724
rect 35843 12100 35877 12116
rect 35843 11708 35877 11724
rect 36101 12100 36135 12116
rect 36101 11708 36135 11724
rect 36215 12100 36249 12116
rect 36215 11708 36249 11724
rect 36473 12100 36507 12116
rect 36473 11708 36507 11724
rect 36587 12100 36621 12116
rect 36587 11708 36621 11724
rect 36845 12100 36879 12116
rect 36845 11708 36879 11724
rect 36959 12100 36993 12116
rect 36959 11708 36993 11724
rect 37217 12100 37251 12116
rect 37217 11708 37251 11724
rect 37331 12100 37365 12116
rect 37331 11708 37365 11724
rect 37589 12100 37623 12116
rect 37589 11708 37623 11724
rect 37703 12100 37737 12116
rect 37703 11708 37737 11724
rect 37961 12100 37995 12116
rect 37961 11708 37995 11724
rect 38075 12100 38109 12116
rect 38075 11708 38109 11724
rect 38333 12100 38367 12116
rect 38333 11708 38367 11724
rect 38447 12100 38481 12116
rect 38447 11708 38481 11724
rect 38705 12100 38739 12116
rect 38705 11708 38739 11724
rect 38819 12100 38853 12116
rect 38819 11708 38853 11724
rect 39077 12100 39111 12116
rect 39077 11708 39111 11724
rect 39191 12100 39225 12116
rect 39191 11708 39225 11724
rect 39449 12100 39483 12116
rect 39449 11708 39483 11724
rect 39563 12100 39597 12116
rect 39563 11708 39597 11724
rect 39821 12100 39855 12116
rect 39821 11708 39855 11724
rect 39935 12100 39969 12116
rect 39935 11708 39969 11724
rect 40193 12100 40227 12116
rect 40193 11708 40227 11724
rect 40307 12100 40341 12116
rect 40307 11708 40341 11724
rect 40565 12100 40599 12116
rect 40565 11708 40599 11724
rect 28821 11631 28837 11665
rect 29005 11631 29021 11665
rect 29193 11631 29209 11665
rect 29377 11631 29393 11665
rect 29565 11631 29581 11665
rect 29749 11631 29765 11665
rect 29937 11631 29953 11665
rect 30121 11631 30137 11665
rect 30309 11631 30325 11665
rect 30493 11631 30509 11665
rect 30681 11631 30697 11665
rect 30865 11631 30881 11665
rect 31053 11631 31069 11665
rect 31237 11631 31253 11665
rect 31425 11631 31441 11665
rect 31609 11631 31625 11665
rect 31797 11631 31813 11665
rect 31981 11631 31997 11665
rect 32169 11631 32185 11665
rect 32353 11631 32369 11665
rect 32541 11631 32557 11665
rect 32725 11631 32741 11665
rect 32913 11631 32929 11665
rect 33097 11631 33113 11665
rect 33285 11631 33301 11665
rect 33469 11631 33485 11665
rect 33657 11631 33673 11665
rect 33841 11631 33857 11665
rect 34029 11631 34045 11665
rect 34213 11631 34229 11665
rect 34401 11631 34417 11665
rect 34585 11631 34601 11665
rect 34773 11631 34789 11665
rect 34957 11631 34973 11665
rect 35145 11631 35161 11665
rect 35329 11631 35345 11665
rect 35517 11631 35533 11665
rect 35701 11631 35717 11665
rect 35889 11631 35905 11665
rect 36073 11631 36089 11665
rect 36261 11631 36277 11665
rect 36445 11631 36461 11665
rect 36633 11631 36649 11665
rect 36817 11631 36833 11665
rect 37005 11631 37021 11665
rect 37189 11631 37205 11665
rect 37377 11631 37393 11665
rect 37561 11631 37577 11665
rect 37749 11631 37765 11665
rect 37933 11631 37949 11665
rect 38121 11631 38137 11665
rect 38305 11631 38321 11665
rect 38493 11631 38509 11665
rect 38677 11631 38693 11665
rect 38865 11631 38881 11665
rect 39049 11631 39065 11665
rect 39237 11631 39253 11665
rect 39421 11631 39437 11665
rect 39609 11631 39625 11665
rect 39793 11631 39809 11665
rect 39981 11631 39997 11665
rect 40165 11631 40181 11665
rect 40353 11631 40369 11665
rect 40537 11631 40553 11665
rect 28821 11523 28837 11557
rect 29005 11523 29021 11557
rect 29193 11523 29209 11557
rect 29377 11523 29393 11557
rect 29565 11523 29581 11557
rect 29749 11523 29765 11557
rect 29937 11523 29953 11557
rect 30121 11523 30137 11557
rect 30309 11523 30325 11557
rect 30493 11523 30509 11557
rect 30681 11523 30697 11557
rect 30865 11523 30881 11557
rect 31053 11523 31069 11557
rect 31237 11523 31253 11557
rect 31425 11523 31441 11557
rect 31609 11523 31625 11557
rect 31797 11523 31813 11557
rect 31981 11523 31997 11557
rect 32169 11523 32185 11557
rect 32353 11523 32369 11557
rect 32541 11523 32557 11557
rect 32725 11523 32741 11557
rect 32913 11523 32929 11557
rect 33097 11523 33113 11557
rect 33285 11523 33301 11557
rect 33469 11523 33485 11557
rect 33657 11523 33673 11557
rect 33841 11523 33857 11557
rect 34029 11523 34045 11557
rect 34213 11523 34229 11557
rect 34401 11523 34417 11557
rect 34585 11523 34601 11557
rect 34773 11523 34789 11557
rect 34957 11523 34973 11557
rect 35145 11523 35161 11557
rect 35329 11523 35345 11557
rect 35517 11523 35533 11557
rect 35701 11523 35717 11557
rect 35889 11523 35905 11557
rect 36073 11523 36089 11557
rect 36261 11523 36277 11557
rect 36445 11523 36461 11557
rect 36633 11523 36649 11557
rect 36817 11523 36833 11557
rect 37005 11523 37021 11557
rect 37189 11523 37205 11557
rect 37377 11523 37393 11557
rect 37561 11523 37577 11557
rect 37749 11523 37765 11557
rect 37933 11523 37949 11557
rect 38121 11523 38137 11557
rect 38305 11523 38321 11557
rect 38493 11523 38509 11557
rect 38677 11523 38693 11557
rect 38865 11523 38881 11557
rect 39049 11523 39065 11557
rect 39237 11523 39253 11557
rect 39421 11523 39437 11557
rect 39609 11523 39625 11557
rect 39793 11523 39809 11557
rect 39981 11523 39997 11557
rect 40165 11523 40181 11557
rect 40353 11523 40369 11557
rect 40537 11523 40553 11557
rect 28775 11464 28809 11480
rect 28775 11072 28809 11088
rect 29033 11464 29067 11480
rect 29033 11072 29067 11088
rect 29147 11464 29181 11480
rect 29147 11072 29181 11088
rect 29405 11464 29439 11480
rect 29405 11072 29439 11088
rect 29519 11464 29553 11480
rect 29519 11072 29553 11088
rect 29777 11464 29811 11480
rect 29777 11072 29811 11088
rect 29891 11464 29925 11480
rect 29891 11072 29925 11088
rect 30149 11464 30183 11480
rect 30149 11072 30183 11088
rect 30263 11464 30297 11480
rect 30263 11072 30297 11088
rect 30521 11464 30555 11480
rect 30521 11072 30555 11088
rect 30635 11464 30669 11480
rect 30635 11072 30669 11088
rect 30893 11464 30927 11480
rect 30893 11072 30927 11088
rect 31007 11464 31041 11480
rect 31007 11072 31041 11088
rect 31265 11464 31299 11480
rect 31265 11072 31299 11088
rect 31379 11464 31413 11480
rect 31379 11072 31413 11088
rect 31637 11464 31671 11480
rect 31637 11072 31671 11088
rect 31751 11464 31785 11480
rect 31751 11072 31785 11088
rect 32009 11464 32043 11480
rect 32009 11072 32043 11088
rect 32123 11464 32157 11480
rect 32123 11072 32157 11088
rect 32381 11464 32415 11480
rect 32381 11072 32415 11088
rect 32495 11464 32529 11480
rect 32495 11072 32529 11088
rect 32753 11464 32787 11480
rect 32753 11072 32787 11088
rect 32867 11464 32901 11480
rect 32867 11072 32901 11088
rect 33125 11464 33159 11480
rect 33125 11072 33159 11088
rect 33239 11464 33273 11480
rect 33239 11072 33273 11088
rect 33497 11464 33531 11480
rect 33497 11072 33531 11088
rect 33611 11464 33645 11480
rect 33611 11072 33645 11088
rect 33869 11464 33903 11480
rect 33869 11072 33903 11088
rect 33983 11464 34017 11480
rect 33983 11072 34017 11088
rect 34241 11464 34275 11480
rect 34241 11072 34275 11088
rect 34355 11464 34389 11480
rect 34355 11072 34389 11088
rect 34613 11464 34647 11480
rect 34613 11072 34647 11088
rect 34727 11464 34761 11480
rect 34727 11072 34761 11088
rect 34985 11464 35019 11480
rect 34985 11072 35019 11088
rect 35099 11464 35133 11480
rect 35099 11072 35133 11088
rect 35357 11464 35391 11480
rect 35357 11072 35391 11088
rect 35471 11464 35505 11480
rect 35471 11072 35505 11088
rect 35729 11464 35763 11480
rect 35729 11072 35763 11088
rect 35843 11464 35877 11480
rect 35843 11072 35877 11088
rect 36101 11464 36135 11480
rect 36101 11072 36135 11088
rect 36215 11464 36249 11480
rect 36215 11072 36249 11088
rect 36473 11464 36507 11480
rect 36473 11072 36507 11088
rect 36587 11464 36621 11480
rect 36587 11072 36621 11088
rect 36845 11464 36879 11480
rect 36845 11072 36879 11088
rect 36959 11464 36993 11480
rect 36959 11072 36993 11088
rect 37217 11464 37251 11480
rect 37217 11072 37251 11088
rect 37331 11464 37365 11480
rect 37331 11072 37365 11088
rect 37589 11464 37623 11480
rect 37589 11072 37623 11088
rect 37703 11464 37737 11480
rect 37703 11072 37737 11088
rect 37961 11464 37995 11480
rect 37961 11072 37995 11088
rect 38075 11464 38109 11480
rect 38075 11072 38109 11088
rect 38333 11464 38367 11480
rect 38333 11072 38367 11088
rect 38447 11464 38481 11480
rect 38447 11072 38481 11088
rect 38705 11464 38739 11480
rect 38705 11072 38739 11088
rect 38819 11464 38853 11480
rect 38819 11072 38853 11088
rect 39077 11464 39111 11480
rect 39077 11072 39111 11088
rect 39191 11464 39225 11480
rect 39191 11072 39225 11088
rect 39449 11464 39483 11480
rect 39449 11072 39483 11088
rect 39563 11464 39597 11480
rect 39563 11072 39597 11088
rect 39821 11464 39855 11480
rect 39821 11072 39855 11088
rect 39935 11464 39969 11480
rect 39935 11072 39969 11088
rect 40193 11464 40227 11480
rect 40193 11072 40227 11088
rect 40307 11464 40341 11480
rect 40307 11072 40341 11088
rect 40565 11464 40599 11480
rect 40565 11072 40599 11088
rect 28821 10995 28837 11029
rect 29005 10995 29021 11029
rect 29193 10995 29209 11029
rect 29377 10995 29393 11029
rect 29565 10995 29581 11029
rect 29749 10995 29765 11029
rect 29937 10995 29953 11029
rect 30121 10995 30137 11029
rect 30309 10995 30325 11029
rect 30493 10995 30509 11029
rect 30681 10995 30697 11029
rect 30865 10995 30881 11029
rect 31053 10995 31069 11029
rect 31237 10995 31253 11029
rect 31425 10995 31441 11029
rect 31609 10995 31625 11029
rect 31797 10995 31813 11029
rect 31981 10995 31997 11029
rect 32169 10995 32185 11029
rect 32353 10995 32369 11029
rect 32541 10995 32557 11029
rect 32725 10995 32741 11029
rect 32913 10995 32929 11029
rect 33097 10995 33113 11029
rect 33285 10995 33301 11029
rect 33469 10995 33485 11029
rect 33657 10995 33673 11029
rect 33841 10995 33857 11029
rect 34029 10995 34045 11029
rect 34213 10995 34229 11029
rect 34401 10995 34417 11029
rect 34585 10995 34601 11029
rect 34773 10995 34789 11029
rect 34957 10995 34973 11029
rect 35145 10995 35161 11029
rect 35329 10995 35345 11029
rect 35517 10995 35533 11029
rect 35701 10995 35717 11029
rect 35889 10995 35905 11029
rect 36073 10995 36089 11029
rect 36261 10995 36277 11029
rect 36445 10995 36461 11029
rect 36633 10995 36649 11029
rect 36817 10995 36833 11029
rect 37005 10995 37021 11029
rect 37189 10995 37205 11029
rect 37377 10995 37393 11029
rect 37561 10995 37577 11029
rect 37749 10995 37765 11029
rect 37933 10995 37949 11029
rect 38121 10995 38137 11029
rect 38305 10995 38321 11029
rect 38493 10995 38509 11029
rect 38677 10995 38693 11029
rect 38865 10995 38881 11029
rect 39049 10995 39065 11029
rect 39237 10995 39253 11029
rect 39421 10995 39437 11029
rect 39609 10995 39625 11029
rect 39793 10995 39809 11029
rect 39981 10995 39997 11029
rect 40165 10995 40181 11029
rect 40353 10995 40369 11029
rect 40537 10995 40553 11029
rect 28821 10887 28837 10921
rect 29005 10887 29021 10921
rect 29193 10887 29209 10921
rect 29377 10887 29393 10921
rect 29565 10887 29581 10921
rect 29749 10887 29765 10921
rect 29937 10887 29953 10921
rect 30121 10887 30137 10921
rect 30309 10887 30325 10921
rect 30493 10887 30509 10921
rect 30681 10887 30697 10921
rect 30865 10887 30881 10921
rect 31053 10887 31069 10921
rect 31237 10887 31253 10921
rect 31425 10887 31441 10921
rect 31609 10887 31625 10921
rect 31797 10887 31813 10921
rect 31981 10887 31997 10921
rect 32169 10887 32185 10921
rect 32353 10887 32369 10921
rect 32541 10887 32557 10921
rect 32725 10887 32741 10921
rect 32913 10887 32929 10921
rect 33097 10887 33113 10921
rect 33285 10887 33301 10921
rect 33469 10887 33485 10921
rect 33657 10887 33673 10921
rect 33841 10887 33857 10921
rect 34029 10887 34045 10921
rect 34213 10887 34229 10921
rect 34401 10887 34417 10921
rect 34585 10887 34601 10921
rect 34773 10887 34789 10921
rect 34957 10887 34973 10921
rect 35145 10887 35161 10921
rect 35329 10887 35345 10921
rect 35517 10887 35533 10921
rect 35701 10887 35717 10921
rect 35889 10887 35905 10921
rect 36073 10887 36089 10921
rect 36261 10887 36277 10921
rect 36445 10887 36461 10921
rect 36633 10887 36649 10921
rect 36817 10887 36833 10921
rect 37005 10887 37021 10921
rect 37189 10887 37205 10921
rect 37377 10887 37393 10921
rect 37561 10887 37577 10921
rect 37749 10887 37765 10921
rect 37933 10887 37949 10921
rect 38121 10887 38137 10921
rect 38305 10887 38321 10921
rect 38493 10887 38509 10921
rect 38677 10887 38693 10921
rect 38865 10887 38881 10921
rect 39049 10887 39065 10921
rect 39237 10887 39253 10921
rect 39421 10887 39437 10921
rect 39609 10887 39625 10921
rect 39793 10887 39809 10921
rect 39981 10887 39997 10921
rect 40165 10887 40181 10921
rect 40353 10887 40369 10921
rect 40537 10887 40553 10921
rect 28775 10828 28809 10844
rect 28775 10436 28809 10452
rect 29033 10828 29067 10844
rect 29033 10436 29067 10452
rect 29147 10828 29181 10844
rect 29147 10436 29181 10452
rect 29405 10828 29439 10844
rect 29405 10436 29439 10452
rect 29519 10828 29553 10844
rect 29519 10436 29553 10452
rect 29777 10828 29811 10844
rect 29777 10436 29811 10452
rect 29891 10828 29925 10844
rect 29891 10436 29925 10452
rect 30149 10828 30183 10844
rect 30149 10436 30183 10452
rect 30263 10828 30297 10844
rect 30263 10436 30297 10452
rect 30521 10828 30555 10844
rect 30521 10436 30555 10452
rect 30635 10828 30669 10844
rect 30635 10436 30669 10452
rect 30893 10828 30927 10844
rect 30893 10436 30927 10452
rect 31007 10828 31041 10844
rect 31007 10436 31041 10452
rect 31265 10828 31299 10844
rect 31265 10436 31299 10452
rect 31379 10828 31413 10844
rect 31379 10436 31413 10452
rect 31637 10828 31671 10844
rect 31637 10436 31671 10452
rect 31751 10828 31785 10844
rect 31751 10436 31785 10452
rect 32009 10828 32043 10844
rect 32009 10436 32043 10452
rect 32123 10828 32157 10844
rect 32123 10436 32157 10452
rect 32381 10828 32415 10844
rect 32381 10436 32415 10452
rect 32495 10828 32529 10844
rect 32495 10436 32529 10452
rect 32753 10828 32787 10844
rect 32753 10436 32787 10452
rect 32867 10828 32901 10844
rect 32867 10436 32901 10452
rect 33125 10828 33159 10844
rect 33125 10436 33159 10452
rect 33239 10828 33273 10844
rect 33239 10436 33273 10452
rect 33497 10828 33531 10844
rect 33497 10436 33531 10452
rect 33611 10828 33645 10844
rect 33611 10436 33645 10452
rect 33869 10828 33903 10844
rect 33869 10436 33903 10452
rect 33983 10828 34017 10844
rect 33983 10436 34017 10452
rect 34241 10828 34275 10844
rect 34241 10436 34275 10452
rect 34355 10828 34389 10844
rect 34355 10436 34389 10452
rect 34613 10828 34647 10844
rect 34613 10436 34647 10452
rect 34727 10828 34761 10844
rect 34727 10436 34761 10452
rect 34985 10828 35019 10844
rect 34985 10436 35019 10452
rect 35099 10828 35133 10844
rect 35099 10436 35133 10452
rect 35357 10828 35391 10844
rect 35357 10436 35391 10452
rect 35471 10828 35505 10844
rect 35471 10436 35505 10452
rect 35729 10828 35763 10844
rect 35729 10436 35763 10452
rect 35843 10828 35877 10844
rect 35843 10436 35877 10452
rect 36101 10828 36135 10844
rect 36101 10436 36135 10452
rect 36215 10828 36249 10844
rect 36215 10436 36249 10452
rect 36473 10828 36507 10844
rect 36473 10436 36507 10452
rect 36587 10828 36621 10844
rect 36587 10436 36621 10452
rect 36845 10828 36879 10844
rect 36845 10436 36879 10452
rect 36959 10828 36993 10844
rect 36959 10436 36993 10452
rect 37217 10828 37251 10844
rect 37217 10436 37251 10452
rect 37331 10828 37365 10844
rect 37331 10436 37365 10452
rect 37589 10828 37623 10844
rect 37589 10436 37623 10452
rect 37703 10828 37737 10844
rect 37703 10436 37737 10452
rect 37961 10828 37995 10844
rect 37961 10436 37995 10452
rect 38075 10828 38109 10844
rect 38075 10436 38109 10452
rect 38333 10828 38367 10844
rect 38333 10436 38367 10452
rect 38447 10828 38481 10844
rect 38447 10436 38481 10452
rect 38705 10828 38739 10844
rect 38705 10436 38739 10452
rect 38819 10828 38853 10844
rect 38819 10436 38853 10452
rect 39077 10828 39111 10844
rect 39077 10436 39111 10452
rect 39191 10828 39225 10844
rect 39191 10436 39225 10452
rect 39449 10828 39483 10844
rect 39449 10436 39483 10452
rect 39563 10828 39597 10844
rect 39563 10436 39597 10452
rect 39821 10828 39855 10844
rect 39821 10436 39855 10452
rect 39935 10828 39969 10844
rect 39935 10436 39969 10452
rect 40193 10828 40227 10844
rect 40193 10436 40227 10452
rect 40307 10828 40341 10844
rect 40307 10436 40341 10452
rect 40565 10828 40599 10844
rect 40565 10436 40599 10452
rect 28821 10359 28837 10393
rect 29005 10359 29021 10393
rect 29193 10359 29209 10393
rect 29377 10359 29393 10393
rect 29565 10359 29581 10393
rect 29749 10359 29765 10393
rect 29937 10359 29953 10393
rect 30121 10359 30137 10393
rect 30309 10359 30325 10393
rect 30493 10359 30509 10393
rect 30681 10359 30697 10393
rect 30865 10359 30881 10393
rect 31053 10359 31069 10393
rect 31237 10359 31253 10393
rect 31425 10359 31441 10393
rect 31609 10359 31625 10393
rect 31797 10359 31813 10393
rect 31981 10359 31997 10393
rect 32169 10359 32185 10393
rect 32353 10359 32369 10393
rect 32541 10359 32557 10393
rect 32725 10359 32741 10393
rect 32913 10359 32929 10393
rect 33097 10359 33113 10393
rect 33285 10359 33301 10393
rect 33469 10359 33485 10393
rect 33657 10359 33673 10393
rect 33841 10359 33857 10393
rect 34029 10359 34045 10393
rect 34213 10359 34229 10393
rect 34401 10359 34417 10393
rect 34585 10359 34601 10393
rect 34773 10359 34789 10393
rect 34957 10359 34973 10393
rect 35145 10359 35161 10393
rect 35329 10359 35345 10393
rect 35517 10359 35533 10393
rect 35701 10359 35717 10393
rect 35889 10359 35905 10393
rect 36073 10359 36089 10393
rect 36261 10359 36277 10393
rect 36445 10359 36461 10393
rect 36633 10359 36649 10393
rect 36817 10359 36833 10393
rect 37005 10359 37021 10393
rect 37189 10359 37205 10393
rect 37377 10359 37393 10393
rect 37561 10359 37577 10393
rect 37749 10359 37765 10393
rect 37933 10359 37949 10393
rect 38121 10359 38137 10393
rect 38305 10359 38321 10393
rect 38493 10359 38509 10393
rect 38677 10359 38693 10393
rect 38865 10359 38881 10393
rect 39049 10359 39065 10393
rect 39237 10359 39253 10393
rect 39421 10359 39437 10393
rect 39609 10359 39625 10393
rect 39793 10359 39809 10393
rect 39981 10359 39997 10393
rect 40165 10359 40181 10393
rect 40353 10359 40369 10393
rect 40537 10359 40553 10393
rect 28661 10291 28695 10353
rect 40679 10291 40713 10353
rect 28661 10257 28757 10291
rect 40617 10257 40713 10291
rect 30149 9873 30234 9907
rect 33177 9873 33273 9907
rect 30149 9811 30183 9873
rect 33239 9811 33273 9873
rect 30309 9771 30325 9805
rect 30493 9771 30509 9805
rect 30681 9771 30697 9805
rect 30865 9771 30881 9805
rect 31053 9771 31069 9805
rect 31237 9771 31253 9805
rect 31425 9771 31441 9805
rect 31609 9771 31625 9805
rect 31797 9771 31813 9805
rect 31981 9771 31997 9805
rect 32169 9771 32185 9805
rect 32353 9771 32369 9805
rect 32541 9771 32557 9805
rect 32725 9771 32741 9805
rect 32913 9771 32929 9805
rect 33097 9771 33113 9805
rect 30263 9712 30297 9728
rect 30263 8920 30297 8936
rect 30521 9712 30555 9728
rect 30521 8920 30555 8936
rect 30635 9712 30669 9728
rect 30635 8920 30669 8936
rect 30893 9712 30927 9728
rect 30893 8920 30927 8936
rect 31007 9712 31041 9728
rect 31007 8920 31041 8936
rect 31265 9712 31299 9728
rect 31265 8920 31299 8936
rect 31379 9712 31413 9728
rect 31379 8920 31413 8936
rect 31637 9712 31671 9728
rect 31637 8920 31671 8936
rect 31751 9712 31785 9728
rect 31751 8920 31785 8936
rect 32009 9712 32043 9728
rect 32009 8920 32043 8936
rect 32123 9712 32157 9728
rect 32123 8920 32157 8936
rect 32381 9712 32415 9728
rect 32381 8920 32415 8936
rect 32495 9712 32529 9728
rect 32495 8920 32529 8936
rect 32753 9712 32787 9728
rect 32753 8920 32787 8936
rect 32867 9712 32901 9728
rect 32867 8920 32901 8936
rect 33125 9712 33159 9728
rect 33125 8920 33159 8936
rect 30309 8843 30325 8877
rect 30493 8843 30509 8877
rect 30681 8843 30697 8877
rect 30865 8843 30881 8877
rect 31053 8843 31069 8877
rect 31237 8843 31253 8877
rect 31425 8843 31441 8877
rect 31609 8843 31625 8877
rect 31797 8843 31813 8877
rect 31981 8843 31997 8877
rect 32169 8843 32185 8877
rect 32353 8843 32369 8877
rect 32541 8843 32557 8877
rect 32725 8843 32741 8877
rect 32913 8843 32929 8877
rect 33097 8843 33113 8877
rect 30309 8735 30325 8769
rect 30493 8735 30509 8769
rect 30681 8735 30697 8769
rect 30865 8735 30881 8769
rect 31053 8735 31069 8769
rect 31237 8735 31253 8769
rect 31425 8735 31441 8769
rect 31609 8735 31625 8769
rect 31797 8735 31813 8769
rect 31981 8735 31997 8769
rect 32169 8735 32185 8769
rect 32353 8735 32369 8769
rect 32541 8735 32557 8769
rect 32725 8735 32741 8769
rect 32913 8735 32929 8769
rect 33097 8735 33113 8769
rect 30263 8676 30297 8692
rect 30263 7884 30297 7900
rect 30521 8676 30555 8692
rect 30521 7884 30555 7900
rect 30635 8676 30669 8692
rect 30635 7884 30669 7900
rect 30893 8676 30927 8692
rect 30893 7884 30927 7900
rect 31007 8676 31041 8692
rect 31007 7884 31041 7900
rect 31265 8676 31299 8692
rect 31265 7884 31299 7900
rect 31379 8676 31413 8692
rect 31379 7884 31413 7900
rect 31637 8676 31671 8692
rect 31637 7884 31671 7900
rect 31751 8676 31785 8692
rect 31751 7884 31785 7900
rect 32009 8676 32043 8692
rect 32009 7884 32043 7900
rect 32123 8676 32157 8692
rect 32123 7884 32157 7900
rect 32381 8676 32415 8692
rect 32381 7884 32415 7900
rect 32495 8676 32529 8692
rect 32495 7884 32529 7900
rect 32753 8676 32787 8692
rect 32753 7884 32787 7900
rect 32867 8676 32901 8692
rect 32867 7884 32901 7900
rect 33125 8676 33159 8692
rect 33125 7884 33159 7900
rect 30309 7807 30325 7841
rect 30493 7807 30509 7841
rect 30681 7807 30697 7841
rect 30865 7807 30881 7841
rect 31053 7807 31069 7841
rect 31237 7807 31253 7841
rect 31425 7807 31441 7841
rect 31609 7807 31625 7841
rect 31797 7807 31813 7841
rect 31981 7807 31997 7841
rect 32169 7807 32185 7841
rect 32353 7807 32369 7841
rect 32541 7807 32557 7841
rect 32725 7807 32741 7841
rect 32913 7807 32929 7841
rect 33097 7807 33113 7841
rect 30309 7699 30325 7733
rect 30493 7699 30509 7733
rect 30681 7699 30697 7733
rect 30865 7699 30881 7733
rect 31053 7699 31069 7733
rect 31237 7699 31253 7733
rect 31425 7699 31441 7733
rect 31609 7699 31625 7733
rect 31797 7699 31813 7733
rect 31981 7699 31997 7733
rect 32169 7699 32185 7733
rect 32353 7699 32369 7733
rect 32541 7699 32557 7733
rect 32725 7699 32741 7733
rect 32913 7699 32929 7733
rect 33097 7699 33113 7733
rect 30263 7640 30297 7656
rect 30263 6848 30297 6864
rect 30521 7640 30555 7656
rect 30521 6848 30555 6864
rect 30635 7640 30669 7656
rect 30635 6848 30669 6864
rect 30893 7640 30927 7656
rect 30893 6848 30927 6864
rect 31007 7640 31041 7656
rect 31007 6848 31041 6864
rect 31265 7640 31299 7656
rect 31265 6848 31299 6864
rect 31379 7640 31413 7656
rect 31379 6848 31413 6864
rect 31637 7640 31671 7656
rect 31637 6848 31671 6864
rect 31751 7640 31785 7656
rect 31751 6848 31785 6864
rect 32009 7640 32043 7656
rect 32009 6848 32043 6864
rect 32123 7640 32157 7656
rect 32123 6848 32157 6864
rect 32381 7640 32415 7656
rect 32381 6848 32415 6864
rect 32495 7640 32529 7656
rect 32495 6848 32529 6864
rect 32753 7640 32787 7656
rect 32753 6848 32787 6864
rect 32867 7640 32901 7656
rect 32867 6848 32901 6864
rect 33125 7640 33159 7656
rect 33125 6848 33159 6864
rect 30309 6771 30325 6805
rect 30493 6771 30509 6805
rect 30681 6771 30697 6805
rect 30865 6771 30881 6805
rect 31053 6771 31069 6805
rect 31237 6771 31253 6805
rect 31425 6771 31441 6805
rect 31609 6771 31625 6805
rect 31797 6771 31813 6805
rect 31981 6771 31997 6805
rect 32169 6771 32185 6805
rect 32353 6771 32369 6805
rect 32541 6771 32557 6805
rect 32725 6771 32741 6805
rect 32913 6771 32929 6805
rect 33097 6771 33113 6805
rect 30309 6663 30325 6697
rect 30493 6663 30509 6697
rect 30681 6663 30697 6697
rect 30865 6663 30881 6697
rect 31053 6663 31069 6697
rect 31237 6663 31253 6697
rect 31425 6663 31441 6697
rect 31609 6663 31625 6697
rect 31797 6663 31813 6697
rect 31981 6663 31997 6697
rect 32169 6663 32185 6697
rect 32353 6663 32369 6697
rect 32541 6663 32557 6697
rect 32725 6663 32741 6697
rect 32913 6663 32929 6697
rect 33097 6663 33113 6697
rect 30263 6604 30297 6620
rect 30263 5812 30297 5828
rect 30521 6604 30555 6620
rect 30521 5812 30555 5828
rect 30635 6604 30669 6620
rect 30635 5812 30669 5828
rect 30893 6604 30927 6620
rect 30893 5812 30927 5828
rect 31007 6604 31041 6620
rect 31007 5812 31041 5828
rect 31265 6604 31299 6620
rect 31265 5812 31299 5828
rect 31379 6604 31413 6620
rect 31379 5812 31413 5828
rect 31637 6604 31671 6620
rect 31637 5812 31671 5828
rect 31751 6604 31785 6620
rect 31751 5812 31785 5828
rect 32009 6604 32043 6620
rect 32009 5812 32043 5828
rect 32123 6604 32157 6620
rect 32123 5812 32157 5828
rect 32381 6604 32415 6620
rect 32381 5812 32415 5828
rect 32495 6604 32529 6620
rect 32495 5812 32529 5828
rect 32753 6604 32787 6620
rect 32753 5812 32787 5828
rect 32867 6604 32901 6620
rect 32867 5812 32901 5828
rect 33125 6604 33159 6620
rect 33125 5812 33159 5828
rect 30309 5735 30325 5769
rect 30493 5735 30509 5769
rect 30681 5735 30697 5769
rect 30865 5735 30881 5769
rect 31053 5735 31069 5769
rect 31237 5735 31253 5769
rect 31425 5735 31441 5769
rect 31609 5735 31625 5769
rect 31797 5735 31813 5769
rect 31981 5735 31997 5769
rect 32169 5735 32185 5769
rect 32353 5735 32369 5769
rect 32541 5735 32557 5769
rect 32725 5735 32741 5769
rect 32913 5735 32929 5769
rect 33097 5735 33113 5769
rect 30149 5667 30183 5729
rect 33776 7574 33872 7608
rect 34010 7574 34106 7608
rect 33776 7512 33810 7574
rect 34072 7512 34106 7574
rect 33776 6238 33810 6300
rect 34072 6238 34106 6300
rect 33776 6204 33872 6238
rect 34010 6204 34106 6238
rect 33239 5667 33273 5729
rect 30149 5633 30245 5667
rect 33177 5633 33273 5667
rect 30149 5179 30245 5213
rect 39129 5179 39225 5213
rect 30149 5117 30183 5179
rect 39191 5117 39225 5179
rect 30309 5077 30325 5111
rect 30493 5077 30509 5111
rect 30681 5077 30697 5111
rect 30865 5077 30881 5111
rect 31053 5077 31069 5111
rect 31237 5077 31253 5111
rect 31425 5077 31441 5111
rect 31609 5077 31625 5111
rect 31797 5077 31813 5111
rect 31981 5077 31997 5111
rect 32169 5077 32185 5111
rect 32353 5077 32369 5111
rect 32541 5077 32557 5111
rect 32725 5077 32741 5111
rect 32913 5077 32929 5111
rect 33097 5077 33113 5111
rect 33285 5077 33301 5111
rect 33469 5077 33485 5111
rect 33657 5077 33673 5111
rect 33841 5077 33857 5111
rect 34029 5077 34045 5111
rect 34213 5077 34229 5111
rect 34401 5077 34417 5111
rect 34585 5077 34601 5111
rect 34773 5077 34789 5111
rect 34957 5077 34973 5111
rect 35145 5077 35161 5111
rect 35329 5077 35345 5111
rect 35517 5077 35533 5111
rect 35701 5077 35717 5111
rect 35889 5077 35905 5111
rect 36073 5077 36089 5111
rect 36261 5077 36277 5111
rect 36445 5077 36461 5111
rect 36633 5077 36649 5111
rect 36817 5077 36833 5111
rect 37005 5077 37021 5111
rect 37189 5077 37205 5111
rect 37377 5077 37393 5111
rect 37561 5077 37577 5111
rect 37749 5077 37765 5111
rect 37933 5077 37949 5111
rect 38121 5077 38137 5111
rect 38305 5077 38321 5111
rect 38493 5077 38509 5111
rect 38677 5077 38693 5111
rect 38865 5077 38881 5111
rect 39049 5077 39065 5111
rect 30263 5027 30297 5043
rect 30263 4835 30297 4851
rect 30521 5027 30555 5043
rect 30521 4835 30555 4851
rect 30635 5027 30669 5043
rect 30635 4835 30669 4851
rect 30893 5027 30927 5043
rect 30893 4835 30927 4851
rect 31007 5027 31041 5043
rect 31007 4835 31041 4851
rect 31265 5027 31299 5043
rect 31265 4835 31299 4851
rect 31379 5027 31413 5043
rect 31379 4835 31413 4851
rect 31637 5027 31671 5043
rect 31637 4835 31671 4851
rect 31751 5027 31785 5043
rect 31751 4835 31785 4851
rect 32009 5027 32043 5043
rect 32009 4835 32043 4851
rect 32123 5027 32157 5043
rect 32123 4835 32157 4851
rect 32381 5027 32415 5043
rect 32381 4835 32415 4851
rect 32495 5027 32529 5043
rect 32495 4835 32529 4851
rect 32753 5027 32787 5043
rect 32753 4835 32787 4851
rect 32867 5027 32901 5043
rect 32867 4835 32901 4851
rect 33125 5027 33159 5043
rect 33125 4835 33159 4851
rect 33239 5027 33273 5043
rect 33239 4835 33273 4851
rect 33497 5027 33531 5043
rect 33497 4835 33531 4851
rect 33611 5027 33645 5043
rect 33611 4835 33645 4851
rect 33869 5027 33903 5043
rect 33869 4835 33903 4851
rect 33983 5027 34017 5043
rect 33983 4835 34017 4851
rect 34241 5027 34275 5043
rect 34241 4835 34275 4851
rect 34355 5027 34389 5043
rect 34355 4835 34389 4851
rect 34613 5027 34647 5043
rect 34613 4835 34647 4851
rect 34727 5027 34761 5043
rect 34727 4835 34761 4851
rect 34985 5027 35019 5043
rect 34985 4835 35019 4851
rect 35099 5027 35133 5043
rect 35099 4835 35133 4851
rect 35357 5027 35391 5043
rect 35357 4835 35391 4851
rect 35471 5027 35505 5043
rect 35471 4835 35505 4851
rect 35729 5027 35763 5043
rect 35729 4835 35763 4851
rect 35843 5027 35877 5043
rect 35843 4835 35877 4851
rect 36101 5027 36135 5043
rect 36101 4835 36135 4851
rect 36215 5027 36249 5043
rect 36215 4835 36249 4851
rect 36473 5027 36507 5043
rect 36473 4835 36507 4851
rect 36587 5027 36621 5043
rect 36587 4835 36621 4851
rect 36845 5027 36879 5043
rect 36845 4835 36879 4851
rect 36959 5027 36993 5043
rect 36959 4835 36993 4851
rect 37217 5027 37251 5043
rect 37217 4835 37251 4851
rect 37331 5027 37365 5043
rect 37331 4835 37365 4851
rect 37589 5027 37623 5043
rect 37589 4835 37623 4851
rect 37703 5027 37737 5043
rect 37703 4835 37737 4851
rect 37961 5027 37995 5043
rect 37961 4835 37995 4851
rect 38075 5027 38109 5043
rect 38075 4835 38109 4851
rect 38333 5027 38367 5043
rect 38333 4835 38367 4851
rect 38447 5027 38481 5043
rect 38447 4835 38481 4851
rect 38705 5027 38739 5043
rect 38705 4835 38739 4851
rect 38819 5027 38853 5043
rect 38819 4835 38853 4851
rect 39077 5027 39111 5043
rect 39077 4835 39111 4851
rect 30309 4767 30325 4801
rect 30493 4767 30509 4801
rect 30681 4767 30697 4801
rect 30865 4767 30881 4801
rect 31053 4767 31069 4801
rect 31237 4767 31253 4801
rect 31425 4767 31441 4801
rect 31609 4767 31625 4801
rect 31797 4767 31813 4801
rect 31981 4767 31997 4801
rect 32169 4767 32185 4801
rect 32353 4767 32369 4801
rect 32541 4767 32557 4801
rect 32725 4767 32741 4801
rect 32913 4767 32929 4801
rect 33097 4767 33113 4801
rect 33285 4767 33301 4801
rect 33469 4767 33485 4801
rect 33657 4767 33673 4801
rect 33841 4767 33857 4801
rect 34029 4767 34045 4801
rect 34213 4767 34229 4801
rect 34401 4767 34417 4801
rect 34585 4767 34601 4801
rect 34773 4767 34789 4801
rect 34957 4767 34973 4801
rect 35145 4767 35161 4801
rect 35329 4767 35345 4801
rect 35517 4767 35533 4801
rect 35701 4767 35717 4801
rect 35889 4767 35905 4801
rect 36073 4767 36089 4801
rect 36261 4767 36277 4801
rect 36445 4767 36461 4801
rect 36633 4767 36649 4801
rect 36817 4767 36833 4801
rect 37005 4767 37021 4801
rect 37189 4767 37205 4801
rect 37377 4767 37393 4801
rect 37561 4767 37577 4801
rect 37749 4767 37765 4801
rect 37933 4767 37949 4801
rect 38121 4767 38137 4801
rect 38305 4767 38321 4801
rect 38493 4767 38509 4801
rect 38677 4767 38693 4801
rect 38865 4767 38881 4801
rect 39049 4767 39065 4801
rect 30309 4659 30325 4693
rect 30493 4659 30509 4693
rect 30681 4659 30697 4693
rect 30865 4659 30881 4693
rect 31053 4659 31069 4693
rect 31237 4659 31253 4693
rect 31425 4659 31441 4693
rect 31609 4659 31625 4693
rect 31797 4659 31813 4693
rect 31981 4659 31997 4693
rect 32169 4659 32185 4693
rect 32353 4659 32369 4693
rect 32541 4659 32557 4693
rect 32725 4659 32741 4693
rect 32913 4659 32929 4693
rect 33097 4659 33113 4693
rect 33285 4659 33301 4693
rect 33469 4659 33485 4693
rect 33657 4659 33673 4693
rect 33841 4659 33857 4693
rect 34029 4659 34045 4693
rect 34213 4659 34229 4693
rect 34401 4659 34417 4693
rect 34585 4659 34601 4693
rect 34773 4659 34789 4693
rect 34957 4659 34973 4693
rect 35145 4659 35161 4693
rect 35329 4659 35345 4693
rect 35517 4659 35533 4693
rect 35701 4659 35717 4693
rect 35889 4659 35905 4693
rect 36073 4659 36089 4693
rect 36261 4659 36277 4693
rect 36445 4659 36461 4693
rect 36633 4659 36649 4693
rect 36817 4659 36833 4693
rect 37005 4659 37021 4693
rect 37189 4659 37205 4693
rect 37377 4659 37393 4693
rect 37561 4659 37577 4693
rect 37749 4659 37765 4693
rect 37933 4659 37949 4693
rect 38121 4659 38137 4693
rect 38305 4659 38321 4693
rect 38493 4659 38509 4693
rect 38677 4659 38693 4693
rect 38865 4659 38881 4693
rect 39049 4659 39065 4693
rect 30263 4609 30297 4625
rect 30263 4417 30297 4433
rect 30521 4609 30555 4625
rect 30521 4417 30555 4433
rect 30635 4609 30669 4625
rect 30635 4417 30669 4433
rect 30893 4609 30927 4625
rect 30893 4417 30927 4433
rect 31007 4609 31041 4625
rect 31007 4417 31041 4433
rect 31265 4609 31299 4625
rect 31265 4417 31299 4433
rect 31379 4609 31413 4625
rect 31379 4417 31413 4433
rect 31637 4609 31671 4625
rect 31637 4417 31671 4433
rect 31751 4609 31785 4625
rect 31751 4417 31785 4433
rect 32009 4609 32043 4625
rect 32009 4417 32043 4433
rect 32123 4609 32157 4625
rect 32123 4417 32157 4433
rect 32381 4609 32415 4625
rect 32381 4417 32415 4433
rect 32495 4609 32529 4625
rect 32495 4417 32529 4433
rect 32753 4609 32787 4625
rect 32753 4417 32787 4433
rect 32867 4609 32901 4625
rect 32867 4417 32901 4433
rect 33125 4609 33159 4625
rect 33125 4417 33159 4433
rect 33239 4609 33273 4625
rect 33239 4417 33273 4433
rect 33497 4609 33531 4625
rect 33497 4417 33531 4433
rect 33611 4609 33645 4625
rect 33611 4417 33645 4433
rect 33869 4609 33903 4625
rect 33869 4417 33903 4433
rect 33983 4609 34017 4625
rect 33983 4417 34017 4433
rect 34241 4609 34275 4625
rect 34241 4417 34275 4433
rect 34355 4609 34389 4625
rect 34355 4417 34389 4433
rect 34613 4609 34647 4625
rect 34613 4417 34647 4433
rect 34727 4609 34761 4625
rect 34727 4417 34761 4433
rect 34985 4609 35019 4625
rect 34985 4417 35019 4433
rect 35099 4609 35133 4625
rect 35099 4417 35133 4433
rect 35357 4609 35391 4625
rect 35357 4417 35391 4433
rect 35471 4609 35505 4625
rect 35471 4417 35505 4433
rect 35729 4609 35763 4625
rect 35729 4417 35763 4433
rect 35843 4609 35877 4625
rect 35843 4417 35877 4433
rect 36101 4609 36135 4625
rect 36101 4417 36135 4433
rect 36215 4609 36249 4625
rect 36215 4417 36249 4433
rect 36473 4609 36507 4625
rect 36473 4417 36507 4433
rect 36587 4609 36621 4625
rect 36587 4417 36621 4433
rect 36845 4609 36879 4625
rect 36845 4417 36879 4433
rect 36959 4609 36993 4625
rect 36959 4417 36993 4433
rect 37217 4609 37251 4625
rect 37217 4417 37251 4433
rect 37331 4609 37365 4625
rect 37331 4417 37365 4433
rect 37589 4609 37623 4625
rect 37589 4417 37623 4433
rect 37703 4609 37737 4625
rect 37703 4417 37737 4433
rect 37961 4609 37995 4625
rect 37961 4417 37995 4433
rect 38075 4609 38109 4625
rect 38075 4417 38109 4433
rect 38333 4609 38367 4625
rect 38333 4417 38367 4433
rect 38447 4609 38481 4625
rect 38447 4417 38481 4433
rect 38705 4609 38739 4625
rect 38705 4417 38739 4433
rect 38819 4609 38853 4625
rect 38819 4417 38853 4433
rect 39077 4609 39111 4625
rect 39077 4417 39111 4433
rect 30309 4349 30325 4383
rect 30493 4349 30509 4383
rect 30681 4349 30697 4383
rect 30865 4349 30881 4383
rect 31053 4349 31069 4383
rect 31237 4349 31253 4383
rect 31425 4349 31441 4383
rect 31609 4349 31625 4383
rect 31797 4349 31813 4383
rect 31981 4349 31997 4383
rect 32169 4349 32185 4383
rect 32353 4349 32369 4383
rect 32541 4349 32557 4383
rect 32725 4349 32741 4383
rect 32913 4349 32929 4383
rect 33097 4349 33113 4383
rect 33285 4349 33301 4383
rect 33469 4349 33485 4383
rect 33657 4349 33673 4383
rect 33841 4349 33857 4383
rect 34029 4349 34045 4383
rect 34213 4349 34229 4383
rect 34401 4349 34417 4383
rect 34585 4349 34601 4383
rect 34773 4349 34789 4383
rect 34957 4349 34973 4383
rect 35145 4349 35161 4383
rect 35329 4349 35345 4383
rect 35517 4349 35533 4383
rect 35701 4349 35717 4383
rect 35889 4349 35905 4383
rect 36073 4349 36089 4383
rect 36261 4349 36277 4383
rect 36445 4349 36461 4383
rect 36633 4349 36649 4383
rect 36817 4349 36833 4383
rect 37005 4349 37021 4383
rect 37189 4349 37205 4383
rect 37377 4349 37393 4383
rect 37561 4349 37577 4383
rect 37749 4349 37765 4383
rect 37933 4349 37949 4383
rect 38121 4349 38137 4383
rect 38305 4349 38321 4383
rect 38493 4349 38509 4383
rect 38677 4349 38693 4383
rect 38865 4349 38881 4383
rect 39049 4349 39065 4383
rect 30309 4241 30325 4275
rect 30493 4241 30509 4275
rect 30681 4241 30697 4275
rect 30865 4241 30881 4275
rect 31053 4241 31069 4275
rect 31237 4241 31253 4275
rect 31425 4241 31441 4275
rect 31609 4241 31625 4275
rect 31797 4241 31813 4275
rect 31981 4241 31997 4275
rect 32169 4241 32185 4275
rect 32353 4241 32369 4275
rect 32541 4241 32557 4275
rect 32725 4241 32741 4275
rect 32913 4241 32929 4275
rect 33097 4241 33113 4275
rect 33285 4241 33301 4275
rect 33469 4241 33485 4275
rect 33657 4241 33673 4275
rect 33841 4241 33857 4275
rect 34029 4241 34045 4275
rect 34213 4241 34229 4275
rect 34401 4241 34417 4275
rect 34585 4241 34601 4275
rect 34773 4241 34789 4275
rect 34957 4241 34973 4275
rect 35145 4241 35161 4275
rect 35329 4241 35345 4275
rect 35517 4241 35533 4275
rect 35701 4241 35717 4275
rect 35889 4241 35905 4275
rect 36073 4241 36089 4275
rect 36261 4241 36277 4275
rect 36445 4241 36461 4275
rect 36633 4241 36649 4275
rect 36817 4241 36833 4275
rect 37005 4241 37021 4275
rect 37189 4241 37205 4275
rect 37377 4241 37393 4275
rect 37561 4241 37577 4275
rect 37749 4241 37765 4275
rect 37933 4241 37949 4275
rect 38121 4241 38137 4275
rect 38305 4241 38321 4275
rect 38493 4241 38509 4275
rect 38677 4241 38693 4275
rect 38865 4241 38881 4275
rect 39049 4241 39065 4275
rect 30263 4191 30297 4207
rect 30263 3999 30297 4015
rect 30521 4191 30555 4207
rect 30521 3999 30555 4015
rect 30635 4191 30669 4207
rect 30635 3999 30669 4015
rect 30893 4191 30927 4207
rect 30893 3999 30927 4015
rect 31007 4191 31041 4207
rect 31007 3999 31041 4015
rect 31265 4191 31299 4207
rect 31265 3999 31299 4015
rect 31379 4191 31413 4207
rect 31379 3999 31413 4015
rect 31637 4191 31671 4207
rect 31637 3999 31671 4015
rect 31751 4191 31785 4207
rect 31751 3999 31785 4015
rect 32009 4191 32043 4207
rect 32009 3999 32043 4015
rect 32123 4191 32157 4207
rect 32123 3999 32157 4015
rect 32381 4191 32415 4207
rect 32381 3999 32415 4015
rect 32495 4191 32529 4207
rect 32495 3999 32529 4015
rect 32753 4191 32787 4207
rect 32753 3999 32787 4015
rect 32867 4191 32901 4207
rect 32867 3999 32901 4015
rect 33125 4191 33159 4207
rect 33125 3999 33159 4015
rect 33239 4191 33273 4207
rect 33239 3999 33273 4015
rect 33497 4191 33531 4207
rect 33497 3999 33531 4015
rect 33611 4191 33645 4207
rect 33611 3999 33645 4015
rect 33869 4191 33903 4207
rect 33869 3999 33903 4015
rect 33983 4191 34017 4207
rect 33983 3999 34017 4015
rect 34241 4191 34275 4207
rect 34241 3999 34275 4015
rect 34355 4191 34389 4207
rect 34355 3999 34389 4015
rect 34613 4191 34647 4207
rect 34613 3999 34647 4015
rect 34727 4191 34761 4207
rect 34727 3999 34761 4015
rect 34985 4191 35019 4207
rect 34985 3999 35019 4015
rect 35099 4191 35133 4207
rect 35099 3999 35133 4015
rect 35357 4191 35391 4207
rect 35357 3999 35391 4015
rect 35471 4191 35505 4207
rect 35471 3999 35505 4015
rect 35729 4191 35763 4207
rect 35729 3999 35763 4015
rect 35843 4191 35877 4207
rect 35843 3999 35877 4015
rect 36101 4191 36135 4207
rect 36101 3999 36135 4015
rect 36215 4191 36249 4207
rect 36215 3999 36249 4015
rect 36473 4191 36507 4207
rect 36473 3999 36507 4015
rect 36587 4191 36621 4207
rect 36587 3999 36621 4015
rect 36845 4191 36879 4207
rect 36845 3999 36879 4015
rect 36959 4191 36993 4207
rect 36959 3999 36993 4015
rect 37217 4191 37251 4207
rect 37217 3999 37251 4015
rect 37331 4191 37365 4207
rect 37331 3999 37365 4015
rect 37589 4191 37623 4207
rect 37589 3999 37623 4015
rect 37703 4191 37737 4207
rect 37703 3999 37737 4015
rect 37961 4191 37995 4207
rect 37961 3999 37995 4015
rect 38075 4191 38109 4207
rect 38075 3999 38109 4015
rect 38333 4191 38367 4207
rect 38333 3999 38367 4015
rect 38447 4191 38481 4207
rect 38447 3999 38481 4015
rect 38705 4191 38739 4207
rect 38705 3999 38739 4015
rect 38819 4191 38853 4207
rect 38819 3999 38853 4015
rect 39077 4191 39111 4207
rect 39077 3999 39111 4015
rect 30309 3931 30325 3965
rect 30493 3931 30509 3965
rect 30681 3931 30697 3965
rect 30865 3931 30881 3965
rect 31053 3931 31069 3965
rect 31237 3931 31253 3965
rect 31425 3931 31441 3965
rect 31609 3931 31625 3965
rect 31797 3931 31813 3965
rect 31981 3931 31997 3965
rect 32169 3931 32185 3965
rect 32353 3931 32369 3965
rect 32541 3931 32557 3965
rect 32725 3931 32741 3965
rect 32913 3931 32929 3965
rect 33097 3931 33113 3965
rect 33285 3931 33301 3965
rect 33469 3931 33485 3965
rect 33657 3931 33673 3965
rect 33841 3931 33857 3965
rect 34029 3931 34045 3965
rect 34213 3931 34229 3965
rect 34401 3931 34417 3965
rect 34585 3931 34601 3965
rect 34773 3931 34789 3965
rect 34957 3931 34973 3965
rect 35145 3931 35161 3965
rect 35329 3931 35345 3965
rect 35517 3931 35533 3965
rect 35701 3931 35717 3965
rect 35889 3931 35905 3965
rect 36073 3931 36089 3965
rect 36261 3931 36277 3965
rect 36445 3931 36461 3965
rect 36633 3931 36649 3965
rect 36817 3931 36833 3965
rect 37005 3931 37021 3965
rect 37189 3931 37205 3965
rect 37377 3931 37393 3965
rect 37561 3931 37577 3965
rect 37749 3931 37765 3965
rect 37933 3931 37949 3965
rect 38121 3931 38137 3965
rect 38305 3931 38321 3965
rect 38493 3931 38509 3965
rect 38677 3931 38693 3965
rect 38865 3931 38881 3965
rect 39049 3931 39065 3965
rect 30309 3823 30325 3857
rect 30493 3823 30509 3857
rect 30681 3823 30697 3857
rect 30865 3823 30881 3857
rect 31053 3823 31069 3857
rect 31237 3823 31253 3857
rect 31425 3823 31441 3857
rect 31609 3823 31625 3857
rect 31797 3823 31813 3857
rect 31981 3823 31997 3857
rect 32169 3823 32185 3857
rect 32353 3823 32369 3857
rect 32541 3823 32557 3857
rect 32725 3823 32741 3857
rect 32913 3823 32929 3857
rect 33097 3823 33113 3857
rect 33285 3823 33301 3857
rect 33469 3823 33485 3857
rect 33657 3823 33673 3857
rect 33841 3823 33857 3857
rect 34029 3823 34045 3857
rect 34213 3823 34229 3857
rect 34401 3823 34417 3857
rect 34585 3823 34601 3857
rect 34773 3823 34789 3857
rect 34957 3823 34973 3857
rect 35145 3823 35161 3857
rect 35329 3823 35345 3857
rect 35517 3823 35533 3857
rect 35701 3823 35717 3857
rect 35889 3823 35905 3857
rect 36073 3823 36089 3857
rect 36261 3823 36277 3857
rect 36445 3823 36461 3857
rect 36633 3823 36649 3857
rect 36817 3823 36833 3857
rect 37005 3823 37021 3857
rect 37189 3823 37205 3857
rect 37377 3823 37393 3857
rect 37561 3823 37577 3857
rect 37749 3823 37765 3857
rect 37933 3823 37949 3857
rect 38121 3823 38137 3857
rect 38305 3823 38321 3857
rect 38493 3823 38509 3857
rect 38677 3823 38693 3857
rect 38865 3823 38881 3857
rect 39049 3823 39065 3857
rect 30263 3773 30297 3789
rect 30263 3581 30297 3597
rect 30521 3773 30555 3789
rect 30521 3581 30555 3597
rect 30635 3773 30669 3789
rect 30635 3581 30669 3597
rect 30893 3773 30927 3789
rect 30893 3581 30927 3597
rect 31007 3773 31041 3789
rect 31007 3581 31041 3597
rect 31265 3773 31299 3789
rect 31265 3581 31299 3597
rect 31379 3773 31413 3789
rect 31379 3581 31413 3597
rect 31637 3773 31671 3789
rect 31637 3581 31671 3597
rect 31751 3773 31785 3789
rect 31751 3581 31785 3597
rect 32009 3773 32043 3789
rect 32009 3581 32043 3597
rect 32123 3773 32157 3789
rect 32123 3581 32157 3597
rect 32381 3773 32415 3789
rect 32381 3581 32415 3597
rect 32495 3773 32529 3789
rect 32495 3581 32529 3597
rect 32753 3773 32787 3789
rect 32753 3581 32787 3597
rect 32867 3773 32901 3789
rect 32867 3581 32901 3597
rect 33125 3773 33159 3789
rect 33125 3581 33159 3597
rect 33239 3773 33273 3789
rect 33239 3581 33273 3597
rect 33497 3773 33531 3789
rect 33497 3581 33531 3597
rect 33611 3773 33645 3789
rect 33611 3581 33645 3597
rect 33869 3773 33903 3789
rect 33869 3581 33903 3597
rect 33983 3773 34017 3789
rect 33983 3581 34017 3597
rect 34241 3773 34275 3789
rect 34241 3581 34275 3597
rect 34355 3773 34389 3789
rect 34355 3581 34389 3597
rect 34613 3773 34647 3789
rect 34613 3581 34647 3597
rect 34727 3773 34761 3789
rect 34727 3581 34761 3597
rect 34985 3773 35019 3789
rect 34985 3581 35019 3597
rect 35099 3773 35133 3789
rect 35099 3581 35133 3597
rect 35357 3773 35391 3789
rect 35357 3581 35391 3597
rect 35471 3773 35505 3789
rect 35471 3581 35505 3597
rect 35729 3773 35763 3789
rect 35729 3581 35763 3597
rect 35843 3773 35877 3789
rect 35843 3581 35877 3597
rect 36101 3773 36135 3789
rect 36101 3581 36135 3597
rect 36215 3773 36249 3789
rect 36215 3581 36249 3597
rect 36473 3773 36507 3789
rect 36473 3581 36507 3597
rect 36587 3773 36621 3789
rect 36587 3581 36621 3597
rect 36845 3773 36879 3789
rect 36845 3581 36879 3597
rect 36959 3773 36993 3789
rect 36959 3581 36993 3597
rect 37217 3773 37251 3789
rect 37217 3581 37251 3597
rect 37331 3773 37365 3789
rect 37331 3581 37365 3597
rect 37589 3773 37623 3789
rect 37589 3581 37623 3597
rect 37703 3773 37737 3789
rect 37703 3581 37737 3597
rect 37961 3773 37995 3789
rect 37961 3581 37995 3597
rect 38075 3773 38109 3789
rect 38075 3581 38109 3597
rect 38333 3773 38367 3789
rect 38333 3581 38367 3597
rect 38447 3773 38481 3789
rect 38447 3581 38481 3597
rect 38705 3773 38739 3789
rect 38705 3581 38739 3597
rect 38819 3773 38853 3789
rect 38819 3581 38853 3597
rect 39077 3773 39111 3789
rect 39077 3581 39111 3597
rect 30309 3513 30325 3547
rect 30493 3513 30509 3547
rect 30681 3513 30697 3547
rect 30865 3513 30881 3547
rect 31053 3513 31069 3547
rect 31237 3513 31253 3547
rect 31425 3513 31441 3547
rect 31609 3513 31625 3547
rect 31797 3513 31813 3547
rect 31981 3513 31997 3547
rect 32169 3513 32185 3547
rect 32353 3513 32369 3547
rect 32541 3513 32557 3547
rect 32725 3513 32741 3547
rect 32913 3513 32929 3547
rect 33097 3513 33113 3547
rect 33285 3513 33301 3547
rect 33469 3513 33485 3547
rect 33657 3513 33673 3547
rect 33841 3513 33857 3547
rect 34029 3513 34045 3547
rect 34213 3513 34229 3547
rect 34401 3513 34417 3547
rect 34585 3513 34601 3547
rect 34773 3513 34789 3547
rect 34957 3513 34973 3547
rect 35145 3513 35161 3547
rect 35329 3513 35345 3547
rect 35517 3513 35533 3547
rect 35701 3513 35717 3547
rect 35889 3513 35905 3547
rect 36073 3513 36089 3547
rect 36261 3513 36277 3547
rect 36445 3513 36461 3547
rect 36633 3513 36649 3547
rect 36817 3513 36833 3547
rect 37005 3513 37021 3547
rect 37189 3513 37205 3547
rect 37377 3513 37393 3547
rect 37561 3513 37577 3547
rect 37749 3513 37765 3547
rect 37933 3513 37949 3547
rect 38121 3513 38137 3547
rect 38305 3513 38321 3547
rect 38493 3513 38509 3547
rect 38677 3513 38693 3547
rect 38865 3513 38881 3547
rect 39049 3513 39065 3547
rect 30149 3445 30183 3507
rect 39191 3445 39225 3507
rect 30149 3411 30245 3445
rect 39129 3411 39225 3445
<< viali >>
rect 29072 12295 29142 12312
rect 29816 12295 29886 12312
rect 30560 12295 30630 12312
rect 31304 12295 31374 12312
rect 32048 12295 32118 12312
rect 32792 12295 32862 12312
rect 33536 12295 33606 12312
rect 34280 12295 34350 12312
rect 34652 12295 34722 12312
rect 35396 12295 35466 12312
rect 36140 12295 36210 12312
rect 36884 12295 36954 12312
rect 37628 12295 37698 12312
rect 38372 12295 38442 12312
rect 39116 12295 39186 12312
rect 39860 12295 39930 12312
rect 40550 12295 40620 12312
rect 29072 12261 29142 12295
rect 29816 12261 29886 12295
rect 30560 12261 30630 12295
rect 31304 12261 31374 12295
rect 32048 12261 32118 12295
rect 32792 12261 32862 12295
rect 33536 12261 33606 12295
rect 34280 12261 34350 12295
rect 34652 12261 34722 12295
rect 35396 12261 35466 12295
rect 36140 12261 36210 12295
rect 36884 12261 36954 12295
rect 37628 12261 37698 12295
rect 38372 12261 38442 12295
rect 39116 12261 39186 12295
rect 39860 12261 39930 12295
rect 40550 12261 40617 12295
rect 40617 12261 40620 12295
rect 29072 12242 29142 12261
rect 29816 12242 29886 12261
rect 30560 12242 30630 12261
rect 31304 12242 31374 12261
rect 32048 12242 32118 12261
rect 32792 12242 32862 12261
rect 33536 12242 33606 12261
rect 34280 12242 34350 12261
rect 34652 12242 34722 12261
rect 35396 12242 35466 12261
rect 36140 12242 36210 12261
rect 36884 12242 36954 12261
rect 37628 12242 37698 12261
rect 38372 12242 38442 12261
rect 39116 12242 39186 12261
rect 39860 12242 39930 12261
rect 40550 12242 40620 12261
rect 28837 12159 29005 12193
rect 29209 12159 29377 12193
rect 29581 12159 29749 12193
rect 29953 12159 30121 12193
rect 30325 12159 30493 12193
rect 30697 12159 30865 12193
rect 31069 12159 31237 12193
rect 31441 12159 31609 12193
rect 31813 12159 31981 12193
rect 32185 12159 32353 12193
rect 32557 12159 32725 12193
rect 32929 12159 33097 12193
rect 33301 12159 33469 12193
rect 33673 12159 33841 12193
rect 34045 12159 34213 12193
rect 34417 12159 34585 12193
rect 34789 12159 34957 12193
rect 35161 12159 35329 12193
rect 35533 12159 35701 12193
rect 35905 12159 36073 12193
rect 36277 12159 36445 12193
rect 36649 12159 36817 12193
rect 37021 12159 37189 12193
rect 37393 12159 37561 12193
rect 37765 12159 37933 12193
rect 38137 12159 38305 12193
rect 38509 12159 38677 12193
rect 38881 12159 39049 12193
rect 39253 12159 39421 12193
rect 39625 12159 39793 12193
rect 39997 12159 40165 12193
rect 40369 12159 40537 12193
rect 28775 11724 28809 12100
rect 29033 11724 29067 12100
rect 29147 11724 29181 12100
rect 29405 11724 29439 12100
rect 29519 11724 29553 12100
rect 29777 11724 29811 12100
rect 29891 11724 29925 12100
rect 30149 11724 30183 12100
rect 30263 11724 30297 12100
rect 30521 11724 30555 12100
rect 30635 11724 30669 12100
rect 30893 11724 30927 12100
rect 31007 11724 31041 12100
rect 31265 11724 31299 12100
rect 31379 11724 31413 12100
rect 31637 11724 31671 12100
rect 31751 11724 31785 12100
rect 32009 11724 32043 12100
rect 32123 11724 32157 12100
rect 32381 11724 32415 12100
rect 32495 11724 32529 12100
rect 32753 11724 32787 12100
rect 32867 11724 32901 12100
rect 33125 11724 33159 12100
rect 33239 11724 33273 12100
rect 33497 11724 33531 12100
rect 33611 11724 33645 12100
rect 33869 11724 33903 12100
rect 33983 11724 34017 12100
rect 34241 11724 34275 12100
rect 34355 11724 34389 12100
rect 34613 11724 34647 12100
rect 34727 11724 34761 12100
rect 34985 11724 35019 12100
rect 35099 11724 35133 12100
rect 35357 11724 35391 12100
rect 35471 11724 35505 12100
rect 35729 11724 35763 12100
rect 35843 11724 35877 12100
rect 36101 11724 36135 12100
rect 36215 11724 36249 12100
rect 36473 11724 36507 12100
rect 36587 11724 36621 12100
rect 36845 11724 36879 12100
rect 36959 11724 36993 12100
rect 37217 11724 37251 12100
rect 37331 11724 37365 12100
rect 37589 11724 37623 12100
rect 37703 11724 37737 12100
rect 37961 11724 37995 12100
rect 38075 11724 38109 12100
rect 38333 11724 38367 12100
rect 38447 11724 38481 12100
rect 38705 11724 38739 12100
rect 38819 11724 38853 12100
rect 39077 11724 39111 12100
rect 39191 11724 39225 12100
rect 39449 11724 39483 12100
rect 39563 11724 39597 12100
rect 39821 11724 39855 12100
rect 39935 11724 39969 12100
rect 40193 11724 40227 12100
rect 40307 11724 40341 12100
rect 40565 11724 40599 12100
rect 28837 11631 29005 11665
rect 29209 11631 29377 11665
rect 29581 11631 29749 11665
rect 29953 11631 30121 11665
rect 30325 11631 30493 11665
rect 30697 11631 30865 11665
rect 31069 11631 31237 11665
rect 31441 11631 31609 11665
rect 31813 11631 31981 11665
rect 32185 11631 32353 11665
rect 32557 11631 32725 11665
rect 32929 11631 33097 11665
rect 33301 11631 33469 11665
rect 33673 11631 33841 11665
rect 34045 11631 34213 11665
rect 34417 11631 34585 11665
rect 34789 11631 34957 11665
rect 35161 11631 35329 11665
rect 35533 11631 35701 11665
rect 35905 11631 36073 11665
rect 36277 11631 36445 11665
rect 36649 11631 36817 11665
rect 37021 11631 37189 11665
rect 37393 11631 37561 11665
rect 37765 11631 37933 11665
rect 38137 11631 38305 11665
rect 38509 11631 38677 11665
rect 38881 11631 39049 11665
rect 39253 11631 39421 11665
rect 39625 11631 39793 11665
rect 39997 11631 40165 11665
rect 40369 11631 40537 11665
rect 28837 11523 29005 11557
rect 29209 11523 29377 11557
rect 29581 11523 29749 11557
rect 29953 11523 30121 11557
rect 30325 11523 30493 11557
rect 30697 11523 30865 11557
rect 31069 11523 31237 11557
rect 31441 11523 31609 11557
rect 31813 11523 31981 11557
rect 32185 11523 32353 11557
rect 32557 11523 32725 11557
rect 32929 11523 33097 11557
rect 33301 11523 33469 11557
rect 33673 11523 33841 11557
rect 34045 11523 34213 11557
rect 34417 11523 34585 11557
rect 34789 11523 34957 11557
rect 35161 11523 35329 11557
rect 35533 11523 35701 11557
rect 35905 11523 36073 11557
rect 36277 11523 36445 11557
rect 36649 11523 36817 11557
rect 37021 11523 37189 11557
rect 37393 11523 37561 11557
rect 37765 11523 37933 11557
rect 38137 11523 38305 11557
rect 38509 11523 38677 11557
rect 38881 11523 39049 11557
rect 39253 11523 39421 11557
rect 39625 11523 39793 11557
rect 39997 11523 40165 11557
rect 40369 11523 40537 11557
rect 28775 11088 28809 11464
rect 29033 11088 29067 11464
rect 29147 11088 29181 11464
rect 29405 11088 29439 11464
rect 29519 11088 29553 11464
rect 29777 11088 29811 11464
rect 29891 11088 29925 11464
rect 30149 11088 30183 11464
rect 30263 11088 30297 11464
rect 30521 11088 30555 11464
rect 30635 11088 30669 11464
rect 30893 11088 30927 11464
rect 31007 11088 31041 11464
rect 31265 11088 31299 11464
rect 31379 11088 31413 11464
rect 31637 11088 31671 11464
rect 31751 11088 31785 11464
rect 32009 11088 32043 11464
rect 32123 11088 32157 11464
rect 32381 11088 32415 11464
rect 32495 11088 32529 11464
rect 32753 11088 32787 11464
rect 32867 11088 32901 11464
rect 33125 11088 33159 11464
rect 33239 11088 33273 11464
rect 33497 11088 33531 11464
rect 33611 11088 33645 11464
rect 33869 11088 33903 11464
rect 33983 11088 34017 11464
rect 34241 11088 34275 11464
rect 34355 11088 34389 11464
rect 34613 11088 34647 11464
rect 34727 11088 34761 11464
rect 34985 11088 35019 11464
rect 35099 11088 35133 11464
rect 35357 11088 35391 11464
rect 35471 11088 35505 11464
rect 35729 11088 35763 11464
rect 35843 11088 35877 11464
rect 36101 11088 36135 11464
rect 36215 11088 36249 11464
rect 36473 11088 36507 11464
rect 36587 11088 36621 11464
rect 36845 11088 36879 11464
rect 36959 11088 36993 11464
rect 37217 11088 37251 11464
rect 37331 11088 37365 11464
rect 37589 11088 37623 11464
rect 37703 11088 37737 11464
rect 37961 11088 37995 11464
rect 38075 11088 38109 11464
rect 38333 11088 38367 11464
rect 38447 11088 38481 11464
rect 38705 11088 38739 11464
rect 38819 11088 38853 11464
rect 39077 11088 39111 11464
rect 39191 11088 39225 11464
rect 39449 11088 39483 11464
rect 39563 11088 39597 11464
rect 39821 11088 39855 11464
rect 39935 11088 39969 11464
rect 40193 11088 40227 11464
rect 40307 11088 40341 11464
rect 40565 11088 40599 11464
rect 28837 10995 29005 11029
rect 29209 10995 29377 11029
rect 29581 10995 29749 11029
rect 29953 10995 30121 11029
rect 30325 10995 30493 11029
rect 30697 10995 30865 11029
rect 31069 10995 31237 11029
rect 31441 10995 31609 11029
rect 31813 10995 31981 11029
rect 32185 10995 32353 11029
rect 32557 10995 32725 11029
rect 32929 10995 33097 11029
rect 33301 10995 33469 11029
rect 33673 10995 33841 11029
rect 34045 10995 34213 11029
rect 34417 10995 34585 11029
rect 34789 10995 34957 11029
rect 35161 10995 35329 11029
rect 35533 10995 35701 11029
rect 35905 10995 36073 11029
rect 36277 10995 36445 11029
rect 36649 10995 36817 11029
rect 37021 10995 37189 11029
rect 37393 10995 37561 11029
rect 37765 10995 37933 11029
rect 38137 10995 38305 11029
rect 38509 10995 38677 11029
rect 38881 10995 39049 11029
rect 39253 10995 39421 11029
rect 39625 10995 39793 11029
rect 39997 10995 40165 11029
rect 40369 10995 40537 11029
rect 28837 10887 29005 10921
rect 29209 10887 29377 10921
rect 29581 10887 29749 10921
rect 29953 10887 30121 10921
rect 30325 10887 30493 10921
rect 30697 10887 30865 10921
rect 31069 10887 31237 10921
rect 31441 10887 31609 10921
rect 31813 10887 31981 10921
rect 32185 10887 32353 10921
rect 32557 10887 32725 10921
rect 32929 10887 33097 10921
rect 33301 10887 33469 10921
rect 33673 10887 33841 10921
rect 34045 10887 34213 10921
rect 34417 10887 34585 10921
rect 34789 10887 34957 10921
rect 35161 10887 35329 10921
rect 35533 10887 35701 10921
rect 35905 10887 36073 10921
rect 36277 10887 36445 10921
rect 36649 10887 36817 10921
rect 37021 10887 37189 10921
rect 37393 10887 37561 10921
rect 37765 10887 37933 10921
rect 38137 10887 38305 10921
rect 38509 10887 38677 10921
rect 38881 10887 39049 10921
rect 39253 10887 39421 10921
rect 39625 10887 39793 10921
rect 39997 10887 40165 10921
rect 40369 10887 40537 10921
rect 28775 10452 28809 10828
rect 29033 10452 29067 10828
rect 29147 10452 29181 10828
rect 29405 10452 29439 10828
rect 29519 10452 29553 10828
rect 29777 10452 29811 10828
rect 29891 10452 29925 10828
rect 30149 10452 30183 10828
rect 30263 10452 30297 10828
rect 30521 10452 30555 10828
rect 30635 10452 30669 10828
rect 30893 10452 30927 10828
rect 31007 10452 31041 10828
rect 31265 10452 31299 10828
rect 31379 10452 31413 10828
rect 31637 10452 31671 10828
rect 31751 10452 31785 10828
rect 32009 10452 32043 10828
rect 32123 10452 32157 10828
rect 32381 10452 32415 10828
rect 32495 10452 32529 10828
rect 32753 10452 32787 10828
rect 32867 10452 32901 10828
rect 33125 10452 33159 10828
rect 33239 10452 33273 10828
rect 33497 10452 33531 10828
rect 33611 10452 33645 10828
rect 33869 10452 33903 10828
rect 33983 10452 34017 10828
rect 34241 10452 34275 10828
rect 34355 10452 34389 10828
rect 34613 10452 34647 10828
rect 34727 10452 34761 10828
rect 34985 10452 35019 10828
rect 35099 10452 35133 10828
rect 35357 10452 35391 10828
rect 35471 10452 35505 10828
rect 35729 10452 35763 10828
rect 35843 10452 35877 10828
rect 36101 10452 36135 10828
rect 36215 10452 36249 10828
rect 36473 10452 36507 10828
rect 36587 10452 36621 10828
rect 36845 10452 36879 10828
rect 36959 10452 36993 10828
rect 37217 10452 37251 10828
rect 37331 10452 37365 10828
rect 37589 10452 37623 10828
rect 37703 10452 37737 10828
rect 37961 10452 37995 10828
rect 38075 10452 38109 10828
rect 38333 10452 38367 10828
rect 38447 10452 38481 10828
rect 38705 10452 38739 10828
rect 38819 10452 38853 10828
rect 39077 10452 39111 10828
rect 39191 10452 39225 10828
rect 39449 10452 39483 10828
rect 39563 10452 39597 10828
rect 39821 10452 39855 10828
rect 39935 10452 39969 10828
rect 40193 10452 40227 10828
rect 40307 10452 40341 10828
rect 40565 10452 40599 10828
rect 28837 10359 29005 10393
rect 29209 10359 29377 10393
rect 29581 10359 29749 10393
rect 29953 10359 30121 10393
rect 30325 10359 30493 10393
rect 30697 10359 30865 10393
rect 31069 10359 31237 10393
rect 31441 10359 31609 10393
rect 31813 10359 31981 10393
rect 32185 10359 32353 10393
rect 32557 10359 32725 10393
rect 32929 10359 33097 10393
rect 33301 10359 33469 10393
rect 33673 10359 33841 10393
rect 34045 10359 34213 10393
rect 34417 10359 34585 10393
rect 34789 10359 34957 10393
rect 35161 10359 35329 10393
rect 35533 10359 35701 10393
rect 35905 10359 36073 10393
rect 36277 10359 36445 10393
rect 36649 10359 36817 10393
rect 37021 10359 37189 10393
rect 37393 10359 37561 10393
rect 37765 10359 37933 10393
rect 38137 10359 38305 10393
rect 38509 10359 38677 10393
rect 38881 10359 39049 10393
rect 39253 10359 39421 10393
rect 39625 10359 39793 10393
rect 39997 10359 40165 10393
rect 40369 10359 40537 10393
rect 30234 9907 30304 9924
rect 30606 9907 30676 9924
rect 30978 9907 31048 9924
rect 31350 9907 31420 9924
rect 31722 9907 31792 9924
rect 32094 9907 32164 9924
rect 32466 9907 32536 9924
rect 32838 9907 32908 9924
rect 33100 9907 33170 9924
rect 30234 9873 30245 9907
rect 30245 9873 30304 9907
rect 30606 9873 30676 9907
rect 30978 9873 31048 9907
rect 31350 9873 31420 9907
rect 31722 9873 31792 9907
rect 32094 9873 32164 9907
rect 32466 9873 32536 9907
rect 32838 9873 32908 9907
rect 33100 9873 33170 9907
rect 30234 9854 30304 9873
rect 30606 9854 30676 9873
rect 30978 9854 31048 9873
rect 31350 9854 31420 9873
rect 31722 9854 31792 9873
rect 32094 9854 32164 9873
rect 32466 9854 32536 9873
rect 32838 9854 32908 9873
rect 33100 9854 33170 9873
rect 30325 9771 30493 9805
rect 30697 9771 30865 9805
rect 31069 9771 31237 9805
rect 31441 9771 31609 9805
rect 31813 9771 31981 9805
rect 32185 9771 32353 9805
rect 32557 9771 32725 9805
rect 32929 9771 33097 9805
rect 30263 8936 30297 9712
rect 30521 8936 30555 9712
rect 30635 8936 30669 9712
rect 30893 8936 30927 9712
rect 31007 8936 31041 9712
rect 31265 8936 31299 9712
rect 31379 8936 31413 9712
rect 31637 8936 31671 9712
rect 31751 8936 31785 9712
rect 32009 8936 32043 9712
rect 32123 8936 32157 9712
rect 32381 8936 32415 9712
rect 32495 8936 32529 9712
rect 32753 8936 32787 9712
rect 32867 8936 32901 9712
rect 33125 8936 33159 9712
rect 30325 8843 30493 8877
rect 30697 8843 30865 8877
rect 31069 8843 31237 8877
rect 31441 8843 31609 8877
rect 31813 8843 31981 8877
rect 32185 8843 32353 8877
rect 32557 8843 32725 8877
rect 32929 8843 33097 8877
rect 30325 8735 30493 8769
rect 30697 8735 30865 8769
rect 31069 8735 31237 8769
rect 31441 8735 31609 8769
rect 31813 8735 31981 8769
rect 32185 8735 32353 8769
rect 32557 8735 32725 8769
rect 32929 8735 33097 8769
rect 30263 7900 30297 8676
rect 30521 7900 30555 8676
rect 30635 7900 30669 8676
rect 30893 7900 30927 8676
rect 31007 7900 31041 8676
rect 31265 7900 31299 8676
rect 31379 7900 31413 8676
rect 31637 7900 31671 8676
rect 31751 7900 31785 8676
rect 32009 7900 32043 8676
rect 32123 7900 32157 8676
rect 32381 7900 32415 8676
rect 32495 7900 32529 8676
rect 32753 7900 32787 8676
rect 32867 7900 32901 8676
rect 33125 7900 33159 8676
rect 30325 7807 30493 7841
rect 30697 7807 30865 7841
rect 31069 7807 31237 7841
rect 31441 7807 31609 7841
rect 31813 7807 31981 7841
rect 32185 7807 32353 7841
rect 32557 7807 32725 7841
rect 32929 7807 33097 7841
rect 30325 7699 30493 7733
rect 30697 7699 30865 7733
rect 31069 7699 31237 7733
rect 31441 7699 31609 7733
rect 31813 7699 31981 7733
rect 32185 7699 32353 7733
rect 32557 7699 32725 7733
rect 32929 7699 33097 7733
rect 30263 6864 30297 7640
rect 30521 6864 30555 7640
rect 30635 6864 30669 7640
rect 30893 6864 30927 7640
rect 31007 6864 31041 7640
rect 31265 6864 31299 7640
rect 31379 6864 31413 7640
rect 31637 6864 31671 7640
rect 31751 6864 31785 7640
rect 32009 6864 32043 7640
rect 32123 6864 32157 7640
rect 32381 6864 32415 7640
rect 32495 6864 32529 7640
rect 32753 6864 32787 7640
rect 32867 6864 32901 7640
rect 33125 6864 33159 7640
rect 30325 6771 30493 6805
rect 30697 6771 30865 6805
rect 31069 6771 31237 6805
rect 31441 6771 31609 6805
rect 31813 6771 31981 6805
rect 32185 6771 32353 6805
rect 32557 6771 32725 6805
rect 32929 6771 33097 6805
rect 30325 6663 30493 6697
rect 30697 6663 30865 6697
rect 31069 6663 31237 6697
rect 31441 6663 31609 6697
rect 31813 6663 31981 6697
rect 32185 6663 32353 6697
rect 32557 6663 32725 6697
rect 32929 6663 33097 6697
rect 30263 5828 30297 6604
rect 30521 5828 30555 6604
rect 30635 5828 30669 6604
rect 30893 5828 30927 6604
rect 31007 5828 31041 6604
rect 31265 5828 31299 6604
rect 31379 5828 31413 6604
rect 31637 5828 31671 6604
rect 31751 5828 31785 6604
rect 32009 5828 32043 6604
rect 32123 5828 32157 6604
rect 32381 5828 32415 6604
rect 32495 5828 32529 6604
rect 32753 5828 32787 6604
rect 32867 5828 32901 6604
rect 33125 5828 33159 6604
rect 30325 5735 30493 5769
rect 30697 5735 30865 5769
rect 31069 5735 31237 5769
rect 31441 5735 31609 5769
rect 31813 5735 31981 5769
rect 32185 5735 32353 5769
rect 32557 5735 32725 5769
rect 32929 5735 33097 5769
rect 33922 7063 33960 7460
rect 34060 7132 34072 7178
rect 34072 7132 34106 7178
rect 34106 7132 34116 7178
rect 33922 6352 33960 6749
rect 34060 6732 34072 6778
rect 34072 6732 34106 6778
rect 34106 6732 34116 6778
rect 34060 6332 34072 6378
rect 34072 6332 34106 6378
rect 34106 6332 34116 6378
rect 30325 5077 30493 5111
rect 30697 5077 30865 5111
rect 31069 5077 31237 5111
rect 31441 5077 31609 5111
rect 31813 5077 31981 5111
rect 32185 5077 32353 5111
rect 32557 5077 32725 5111
rect 32929 5077 33097 5111
rect 33301 5077 33469 5111
rect 33673 5077 33841 5111
rect 34045 5077 34213 5111
rect 34417 5077 34585 5111
rect 34789 5077 34957 5111
rect 35161 5077 35329 5111
rect 35533 5077 35701 5111
rect 35905 5077 36073 5111
rect 36277 5077 36445 5111
rect 36649 5077 36817 5111
rect 37021 5077 37189 5111
rect 37393 5077 37561 5111
rect 37765 5077 37933 5111
rect 38137 5077 38305 5111
rect 38509 5077 38677 5111
rect 38881 5077 39049 5111
rect 30263 4851 30297 5027
rect 30521 4851 30555 5027
rect 30635 4851 30669 5027
rect 30893 4851 30927 5027
rect 31007 4851 31041 5027
rect 31265 4851 31299 5027
rect 31379 4851 31413 5027
rect 31637 4851 31671 5027
rect 31751 4851 31785 5027
rect 32009 4851 32043 5027
rect 32123 4851 32157 5027
rect 32381 4851 32415 5027
rect 32495 4851 32529 5027
rect 32753 4851 32787 5027
rect 32867 4851 32901 5027
rect 33125 4851 33159 5027
rect 33239 4851 33273 5027
rect 33497 4851 33531 5027
rect 33611 4851 33645 5027
rect 33869 4851 33903 5027
rect 33983 4851 34017 5027
rect 34241 4851 34275 5027
rect 34355 4851 34389 5027
rect 34613 4851 34647 5027
rect 34727 4851 34761 5027
rect 34985 4851 35019 5027
rect 35099 4851 35133 5027
rect 35357 4851 35391 5027
rect 35471 4851 35505 5027
rect 35729 4851 35763 5027
rect 35843 4851 35877 5027
rect 36101 4851 36135 5027
rect 36215 4851 36249 5027
rect 36473 4851 36507 5027
rect 36587 4851 36621 5027
rect 36845 4851 36879 5027
rect 36959 4851 36993 5027
rect 37217 4851 37251 5027
rect 37331 4851 37365 5027
rect 37589 4851 37623 5027
rect 37703 4851 37737 5027
rect 37961 4851 37995 5027
rect 38075 4851 38109 5027
rect 38333 4851 38367 5027
rect 38447 4851 38481 5027
rect 38705 4851 38739 5027
rect 38819 4851 38853 5027
rect 39077 4851 39111 5027
rect 30325 4767 30493 4801
rect 30697 4767 30865 4801
rect 31069 4767 31237 4801
rect 31441 4767 31609 4801
rect 31813 4767 31981 4801
rect 32185 4767 32353 4801
rect 32557 4767 32725 4801
rect 32929 4767 33097 4801
rect 33301 4767 33469 4801
rect 33673 4767 33841 4801
rect 34045 4767 34213 4801
rect 34417 4767 34585 4801
rect 34789 4767 34957 4801
rect 35161 4767 35329 4801
rect 35533 4767 35701 4801
rect 35905 4767 36073 4801
rect 36277 4767 36445 4801
rect 36649 4767 36817 4801
rect 37021 4767 37189 4801
rect 37393 4767 37561 4801
rect 37765 4767 37933 4801
rect 38137 4767 38305 4801
rect 38509 4767 38677 4801
rect 38881 4767 39049 4801
rect 30325 4659 30493 4693
rect 30697 4659 30865 4693
rect 31069 4659 31237 4693
rect 31441 4659 31609 4693
rect 31813 4659 31981 4693
rect 32185 4659 32353 4693
rect 32557 4659 32725 4693
rect 32929 4659 33097 4693
rect 33301 4659 33469 4693
rect 33673 4659 33841 4693
rect 34045 4659 34213 4693
rect 34417 4659 34585 4693
rect 34789 4659 34957 4693
rect 35161 4659 35329 4693
rect 35533 4659 35701 4693
rect 35905 4659 36073 4693
rect 36277 4659 36445 4693
rect 36649 4659 36817 4693
rect 37021 4659 37189 4693
rect 37393 4659 37561 4693
rect 37765 4659 37933 4693
rect 38137 4659 38305 4693
rect 38509 4659 38677 4693
rect 38881 4659 39049 4693
rect 30263 4433 30297 4609
rect 30521 4433 30555 4609
rect 30635 4433 30669 4609
rect 30893 4433 30927 4609
rect 31007 4433 31041 4609
rect 31265 4433 31299 4609
rect 31379 4433 31413 4609
rect 31637 4433 31671 4609
rect 31751 4433 31785 4609
rect 32009 4433 32043 4609
rect 32123 4433 32157 4609
rect 32381 4433 32415 4609
rect 32495 4433 32529 4609
rect 32753 4433 32787 4609
rect 32867 4433 32901 4609
rect 33125 4433 33159 4609
rect 33239 4433 33273 4609
rect 33497 4433 33531 4609
rect 33611 4433 33645 4609
rect 33869 4433 33903 4609
rect 33983 4433 34017 4609
rect 34241 4433 34275 4609
rect 34355 4433 34389 4609
rect 34613 4433 34647 4609
rect 34727 4433 34761 4609
rect 34985 4433 35019 4609
rect 35099 4433 35133 4609
rect 35357 4433 35391 4609
rect 35471 4433 35505 4609
rect 35729 4433 35763 4609
rect 35843 4433 35877 4609
rect 36101 4433 36135 4609
rect 36215 4433 36249 4609
rect 36473 4433 36507 4609
rect 36587 4433 36621 4609
rect 36845 4433 36879 4609
rect 36959 4433 36993 4609
rect 37217 4433 37251 4609
rect 37331 4433 37365 4609
rect 37589 4433 37623 4609
rect 37703 4433 37737 4609
rect 37961 4433 37995 4609
rect 38075 4433 38109 4609
rect 38333 4433 38367 4609
rect 38447 4433 38481 4609
rect 38705 4433 38739 4609
rect 38819 4433 38853 4609
rect 39077 4433 39111 4609
rect 30325 4349 30493 4383
rect 30697 4349 30865 4383
rect 31069 4349 31237 4383
rect 31441 4349 31609 4383
rect 31813 4349 31981 4383
rect 32185 4349 32353 4383
rect 32557 4349 32725 4383
rect 32929 4349 33097 4383
rect 33301 4349 33469 4383
rect 33673 4349 33841 4383
rect 34045 4349 34213 4383
rect 34417 4349 34585 4383
rect 34789 4349 34957 4383
rect 35161 4349 35329 4383
rect 35533 4349 35701 4383
rect 35905 4349 36073 4383
rect 36277 4349 36445 4383
rect 36649 4349 36817 4383
rect 37021 4349 37189 4383
rect 37393 4349 37561 4383
rect 37765 4349 37933 4383
rect 38137 4349 38305 4383
rect 38509 4349 38677 4383
rect 38881 4349 39049 4383
rect 30325 4241 30493 4275
rect 30697 4241 30865 4275
rect 31069 4241 31237 4275
rect 31441 4241 31609 4275
rect 31813 4241 31981 4275
rect 32185 4241 32353 4275
rect 32557 4241 32725 4275
rect 32929 4241 33097 4275
rect 33301 4241 33469 4275
rect 33673 4241 33841 4275
rect 34045 4241 34213 4275
rect 34417 4241 34585 4275
rect 34789 4241 34957 4275
rect 35161 4241 35329 4275
rect 35533 4241 35701 4275
rect 35905 4241 36073 4275
rect 36277 4241 36445 4275
rect 36649 4241 36817 4275
rect 37021 4241 37189 4275
rect 37393 4241 37561 4275
rect 37765 4241 37933 4275
rect 38137 4241 38305 4275
rect 38509 4241 38677 4275
rect 38881 4241 39049 4275
rect 30263 4015 30297 4191
rect 30521 4015 30555 4191
rect 30635 4015 30669 4191
rect 30893 4015 30927 4191
rect 31007 4015 31041 4191
rect 31265 4015 31299 4191
rect 31379 4015 31413 4191
rect 31637 4015 31671 4191
rect 31751 4015 31785 4191
rect 32009 4015 32043 4191
rect 32123 4015 32157 4191
rect 32381 4015 32415 4191
rect 32495 4015 32529 4191
rect 32753 4015 32787 4191
rect 32867 4015 32901 4191
rect 33125 4015 33159 4191
rect 33239 4015 33273 4191
rect 33497 4015 33531 4191
rect 33611 4015 33645 4191
rect 33869 4015 33903 4191
rect 33983 4015 34017 4191
rect 34241 4015 34275 4191
rect 34355 4015 34389 4191
rect 34613 4015 34647 4191
rect 34727 4015 34761 4191
rect 34985 4015 35019 4191
rect 35099 4015 35133 4191
rect 35357 4015 35391 4191
rect 35471 4015 35505 4191
rect 35729 4015 35763 4191
rect 35843 4015 35877 4191
rect 36101 4015 36135 4191
rect 36215 4015 36249 4191
rect 36473 4015 36507 4191
rect 36587 4015 36621 4191
rect 36845 4015 36879 4191
rect 36959 4015 36993 4191
rect 37217 4015 37251 4191
rect 37331 4015 37365 4191
rect 37589 4015 37623 4191
rect 37703 4015 37737 4191
rect 37961 4015 37995 4191
rect 38075 4015 38109 4191
rect 38333 4015 38367 4191
rect 38447 4015 38481 4191
rect 38705 4015 38739 4191
rect 38819 4015 38853 4191
rect 39077 4015 39111 4191
rect 30325 3931 30493 3965
rect 30697 3931 30865 3965
rect 31069 3931 31237 3965
rect 31441 3931 31609 3965
rect 31813 3931 31981 3965
rect 32185 3931 32353 3965
rect 32557 3931 32725 3965
rect 32929 3931 33097 3965
rect 33301 3931 33469 3965
rect 33673 3931 33841 3965
rect 34045 3931 34213 3965
rect 34417 3931 34585 3965
rect 34789 3931 34957 3965
rect 35161 3931 35329 3965
rect 35533 3931 35701 3965
rect 35905 3931 36073 3965
rect 36277 3931 36445 3965
rect 36649 3931 36817 3965
rect 37021 3931 37189 3965
rect 37393 3931 37561 3965
rect 37765 3931 37933 3965
rect 38137 3931 38305 3965
rect 38509 3931 38677 3965
rect 38881 3931 39049 3965
rect 30325 3823 30493 3857
rect 30697 3823 30865 3857
rect 31069 3823 31237 3857
rect 31441 3823 31609 3857
rect 31813 3823 31981 3857
rect 32185 3823 32353 3857
rect 32557 3823 32725 3857
rect 32929 3823 33097 3857
rect 33301 3823 33469 3857
rect 33673 3823 33841 3857
rect 34045 3823 34213 3857
rect 34417 3823 34585 3857
rect 34789 3823 34957 3857
rect 35161 3823 35329 3857
rect 35533 3823 35701 3857
rect 35905 3823 36073 3857
rect 36277 3823 36445 3857
rect 36649 3823 36817 3857
rect 37021 3823 37189 3857
rect 37393 3823 37561 3857
rect 37765 3823 37933 3857
rect 38137 3823 38305 3857
rect 38509 3823 38677 3857
rect 38881 3823 39049 3857
rect 30263 3597 30297 3773
rect 30521 3597 30555 3773
rect 30635 3597 30669 3773
rect 30893 3597 30927 3773
rect 31007 3597 31041 3773
rect 31265 3597 31299 3773
rect 31379 3597 31413 3773
rect 31637 3597 31671 3773
rect 31751 3597 31785 3773
rect 32009 3597 32043 3773
rect 32123 3597 32157 3773
rect 32381 3597 32415 3773
rect 32495 3597 32529 3773
rect 32753 3597 32787 3773
rect 32867 3597 32901 3773
rect 33125 3597 33159 3773
rect 33239 3597 33273 3773
rect 33497 3597 33531 3773
rect 33611 3597 33645 3773
rect 33869 3597 33903 3773
rect 33983 3597 34017 3773
rect 34241 3597 34275 3773
rect 34355 3597 34389 3773
rect 34613 3597 34647 3773
rect 34727 3597 34761 3773
rect 34985 3597 35019 3773
rect 35099 3597 35133 3773
rect 35357 3597 35391 3773
rect 35471 3597 35505 3773
rect 35729 3597 35763 3773
rect 35843 3597 35877 3773
rect 36101 3597 36135 3773
rect 36215 3597 36249 3773
rect 36473 3597 36507 3773
rect 36587 3597 36621 3773
rect 36845 3597 36879 3773
rect 36959 3597 36993 3773
rect 37217 3597 37251 3773
rect 37331 3597 37365 3773
rect 37589 3597 37623 3773
rect 37703 3597 37737 3773
rect 37961 3597 37995 3773
rect 38075 3597 38109 3773
rect 38333 3597 38367 3773
rect 38447 3597 38481 3773
rect 38705 3597 38739 3773
rect 38819 3597 38853 3773
rect 39077 3597 39111 3773
rect 30325 3513 30493 3547
rect 30697 3513 30865 3547
rect 31069 3513 31237 3547
rect 31441 3513 31609 3547
rect 31813 3513 31981 3547
rect 32185 3513 32353 3547
rect 32557 3513 32725 3547
rect 32929 3513 33097 3547
rect 33301 3513 33469 3547
rect 33673 3513 33841 3547
rect 34045 3513 34213 3547
rect 34417 3513 34585 3547
rect 34789 3513 34957 3547
rect 35161 3513 35329 3547
rect 35533 3513 35701 3547
rect 35905 3513 36073 3547
rect 36277 3513 36445 3547
rect 36649 3513 36817 3547
rect 37021 3513 37189 3547
rect 37393 3513 37561 3547
rect 37765 3513 37933 3547
rect 38137 3513 38305 3547
rect 38509 3513 38677 3547
rect 38881 3513 39049 3547
rect 30264 3445 30334 3456
rect 30932 3445 31002 3464
rect 31676 3445 31746 3464
rect 32420 3445 32490 3464
rect 33164 3445 33234 3464
rect 33908 3445 33978 3464
rect 34652 3445 34722 3464
rect 35396 3445 35466 3464
rect 36140 3445 36210 3464
rect 36884 3445 36954 3464
rect 37628 3445 37698 3464
rect 38372 3445 38442 3464
rect 39034 3445 39104 3460
rect 30264 3411 30334 3445
rect 30932 3411 31002 3445
rect 31676 3411 31746 3445
rect 32420 3411 32490 3445
rect 33164 3411 33234 3445
rect 33908 3411 33978 3445
rect 34652 3411 34722 3445
rect 35396 3411 35466 3445
rect 36140 3411 36210 3445
rect 36884 3411 36954 3445
rect 37628 3411 37698 3445
rect 38372 3411 38442 3445
rect 39034 3411 39104 3445
rect 30264 3386 30334 3411
rect 30932 3394 31002 3411
rect 31676 3394 31746 3411
rect 32420 3394 32490 3411
rect 33164 3394 33234 3411
rect 33908 3394 33978 3411
rect 34652 3394 34722 3411
rect 35396 3394 35466 3411
rect 36140 3394 36210 3411
rect 36884 3394 36954 3411
rect 37628 3394 37698 3411
rect 38372 3394 38442 3411
rect 39034 3390 39104 3411
<< metal1 >>
rect 28996 12394 29006 12594
rect 29206 12394 29216 12594
rect 29740 12394 29750 12594
rect 29950 12394 29960 12594
rect 30484 12394 30494 12594
rect 30694 12394 30704 12594
rect 31228 12394 31238 12594
rect 31438 12394 31448 12594
rect 31972 12394 31982 12594
rect 32182 12394 32192 12594
rect 32716 12394 32726 12594
rect 32926 12394 32936 12594
rect 33460 12394 33470 12594
rect 33670 12394 33680 12594
rect 34204 12394 34214 12594
rect 34414 12394 34424 12594
rect 34576 12394 34586 12594
rect 34786 12394 34796 12594
rect 35320 12394 35330 12594
rect 35530 12394 35540 12594
rect 36064 12394 36074 12594
rect 36274 12394 36284 12594
rect 36808 12394 36818 12594
rect 37018 12394 37028 12594
rect 37552 12394 37562 12594
rect 37762 12394 37772 12594
rect 38296 12394 38306 12594
rect 38506 12394 38516 12594
rect 39040 12394 39050 12594
rect 39250 12394 39260 12594
rect 39784 12394 39794 12594
rect 39994 12394 40004 12594
rect 40528 12394 40538 12594
rect 40738 12394 40748 12594
rect 29078 12318 29136 12394
rect 29822 12318 29880 12394
rect 30566 12318 30624 12394
rect 31310 12318 31368 12394
rect 32054 12318 32112 12394
rect 32798 12318 32856 12394
rect 33542 12318 33600 12394
rect 34266 12384 34344 12394
rect 34286 12318 34344 12384
rect 34696 12318 34748 12394
rect 35402 12318 35460 12394
rect 36146 12318 36204 12394
rect 36890 12318 36948 12394
rect 37634 12318 37692 12394
rect 38378 12318 38436 12394
rect 39122 12318 39180 12394
rect 39866 12318 39924 12394
rect 40592 12378 40668 12394
rect 40592 12318 40650 12378
rect 29060 12312 29154 12318
rect 29060 12242 29072 12312
rect 29142 12242 29154 12312
rect 29060 12236 29154 12242
rect 29804 12312 29898 12318
rect 29804 12242 29816 12312
rect 29886 12242 29898 12312
rect 29804 12236 29898 12242
rect 30548 12312 30642 12318
rect 30548 12242 30560 12312
rect 30630 12242 30642 12312
rect 30548 12236 30642 12242
rect 31292 12312 31386 12318
rect 31292 12242 31304 12312
rect 31374 12242 31386 12312
rect 31292 12236 31386 12242
rect 32036 12312 32130 12318
rect 32036 12242 32048 12312
rect 32118 12242 32130 12312
rect 32036 12236 32130 12242
rect 32780 12312 32874 12318
rect 32780 12242 32792 12312
rect 32862 12242 32874 12312
rect 32780 12236 32874 12242
rect 33524 12312 33618 12318
rect 33524 12242 33536 12312
rect 33606 12242 33618 12312
rect 33524 12236 33618 12242
rect 34268 12312 34362 12318
rect 34268 12242 34280 12312
rect 34350 12242 34362 12312
rect 34268 12236 34362 12242
rect 34640 12312 34748 12318
rect 34640 12242 34652 12312
rect 34722 12242 34748 12312
rect 34640 12236 34748 12242
rect 35384 12312 35478 12318
rect 35384 12242 35396 12312
rect 35466 12242 35478 12312
rect 35384 12236 35478 12242
rect 36128 12312 36222 12318
rect 36128 12242 36140 12312
rect 36210 12242 36222 12312
rect 36128 12236 36222 12242
rect 36872 12312 36966 12318
rect 36872 12242 36884 12312
rect 36954 12242 36966 12312
rect 36872 12236 36966 12242
rect 37616 12312 37710 12318
rect 37616 12242 37628 12312
rect 37698 12242 37710 12312
rect 37616 12236 37710 12242
rect 38360 12312 38454 12318
rect 38360 12242 38372 12312
rect 38442 12242 38454 12312
rect 38360 12236 38454 12242
rect 39104 12312 39198 12318
rect 39104 12242 39116 12312
rect 39186 12242 39198 12312
rect 39104 12236 39198 12242
rect 39848 12312 39942 12318
rect 39848 12242 39860 12312
rect 39930 12242 39942 12312
rect 39848 12236 39942 12242
rect 40538 12312 40650 12318
rect 40538 12242 40550 12312
rect 40620 12242 40650 12312
rect 40538 12236 40650 12242
rect 28768 12146 28836 12206
rect 29006 12199 29016 12206
rect 29006 12153 29017 12199
rect 29006 12146 29016 12153
rect 28768 12100 28816 12146
rect 29078 12112 29136 12236
rect 29198 12199 29208 12206
rect 29197 12153 29208 12199
rect 29378 12199 29388 12206
rect 29570 12199 29580 12206
rect 29198 12146 29208 12153
rect 29378 12153 29389 12199
rect 29569 12153 29580 12199
rect 29750 12199 29760 12206
rect 29378 12146 29388 12153
rect 29570 12146 29580 12153
rect 29750 12153 29761 12199
rect 29750 12146 29760 12153
rect 29822 12112 29880 12236
rect 29942 12199 29952 12206
rect 29941 12153 29952 12199
rect 29942 12146 29952 12153
rect 30122 12146 30324 12206
rect 30494 12199 30504 12206
rect 30494 12153 30505 12199
rect 30494 12146 30504 12153
rect 30194 12112 30252 12146
rect 30566 12112 30624 12236
rect 30686 12199 30696 12206
rect 30685 12153 30696 12199
rect 30866 12199 30876 12206
rect 31058 12199 31068 12206
rect 30686 12146 30696 12153
rect 30866 12153 30877 12199
rect 31057 12153 31068 12199
rect 31238 12199 31248 12206
rect 30866 12146 30876 12153
rect 31058 12146 31068 12153
rect 31238 12153 31249 12199
rect 31238 12146 31248 12153
rect 31310 12112 31368 12236
rect 31430 12199 31440 12206
rect 31429 12153 31440 12199
rect 31430 12146 31440 12153
rect 31610 12146 31812 12206
rect 31982 12199 31992 12206
rect 31982 12153 31993 12199
rect 31982 12146 31992 12153
rect 31682 12112 31740 12146
rect 32054 12112 32112 12236
rect 32174 12199 32184 12206
rect 32173 12153 32184 12199
rect 32354 12199 32364 12206
rect 32546 12199 32556 12206
rect 32174 12146 32184 12153
rect 32354 12153 32365 12199
rect 32545 12153 32556 12199
rect 32726 12199 32736 12206
rect 32354 12146 32364 12153
rect 32546 12146 32556 12153
rect 32726 12153 32737 12199
rect 32726 12146 32736 12153
rect 32798 12112 32856 12236
rect 32918 12199 32928 12206
rect 32917 12153 32928 12199
rect 32918 12146 32928 12153
rect 33098 12146 33300 12206
rect 33470 12199 33480 12206
rect 33470 12153 33481 12199
rect 33470 12146 33480 12153
rect 33170 12112 33228 12146
rect 33542 12112 33600 12236
rect 33662 12199 33672 12206
rect 33661 12153 33672 12199
rect 33842 12199 33852 12206
rect 34034 12199 34044 12206
rect 33662 12146 33672 12153
rect 33842 12153 33853 12199
rect 34033 12153 34044 12199
rect 34214 12199 34224 12206
rect 33842 12146 33852 12153
rect 34034 12146 34044 12153
rect 34214 12153 34225 12199
rect 34214 12146 34224 12153
rect 34286 12112 34344 12236
rect 34406 12199 34416 12206
rect 34405 12153 34416 12199
rect 34406 12146 34416 12153
rect 34586 12146 34658 12206
rect 28768 11724 28775 12100
rect 28809 11724 28816 12100
rect 28768 11672 28816 11724
rect 29027 12100 29187 12112
rect 29027 11724 29033 12100
rect 29067 11724 29147 12100
rect 29181 11724 29187 12100
rect 29027 11712 29187 11724
rect 29399 12100 29559 12112
rect 29399 11724 29405 12100
rect 29439 11724 29519 12100
rect 29553 11724 29559 12100
rect 29399 11712 29559 11724
rect 29771 12100 29931 12112
rect 29771 11724 29777 12100
rect 29811 11724 29891 12100
rect 29925 11724 29931 12100
rect 29771 11712 29931 11724
rect 30143 12100 30303 12112
rect 30143 11724 30149 12100
rect 30183 11724 30263 12100
rect 30297 11724 30303 12100
rect 30143 11712 30303 11724
rect 30515 12100 30675 12112
rect 30515 11724 30521 12100
rect 30555 11724 30635 12100
rect 30669 11724 30675 12100
rect 30515 11712 30675 11724
rect 30887 12100 31047 12112
rect 30887 11724 30893 12100
rect 30927 11724 31007 12100
rect 31041 11724 31047 12100
rect 30887 11712 31047 11724
rect 31259 12100 31419 12112
rect 31259 11724 31265 12100
rect 31299 11724 31379 12100
rect 31413 11724 31419 12100
rect 31259 11712 31419 11724
rect 31631 12100 31791 12112
rect 31631 11724 31637 12100
rect 31671 11724 31751 12100
rect 31785 11724 31791 12100
rect 31631 11712 31791 11724
rect 32003 12100 32163 12112
rect 32003 11724 32009 12100
rect 32043 11724 32123 12100
rect 32157 11724 32163 12100
rect 32003 11712 32163 11724
rect 32375 12100 32535 12112
rect 32375 11724 32381 12100
rect 32415 11724 32495 12100
rect 32529 11724 32535 12100
rect 32375 11712 32535 11724
rect 32747 12100 32907 12112
rect 32747 11724 32753 12100
rect 32787 11724 32867 12100
rect 32901 11724 32907 12100
rect 32747 11712 32907 11724
rect 33119 12100 33279 12112
rect 33119 11724 33125 12100
rect 33159 11724 33239 12100
rect 33273 11724 33279 12100
rect 33119 11712 33279 11724
rect 33491 12100 33651 12112
rect 33491 11724 33497 12100
rect 33531 11724 33611 12100
rect 33645 11724 33651 12100
rect 33491 11712 33651 11724
rect 33863 12100 34023 12112
rect 33863 11724 33869 12100
rect 33903 11724 33983 12100
rect 34017 11724 34023 12100
rect 33863 11712 34023 11724
rect 34235 12100 34395 12112
rect 34235 11724 34241 12100
rect 34275 11724 34355 12100
rect 34389 11724 34395 12100
rect 34235 11712 34395 11724
rect 34606 12100 34658 12146
rect 34606 11724 34613 12100
rect 34647 11724 34658 12100
rect 28768 11671 28856 11672
rect 28768 11666 29017 11671
rect 28768 11522 28836 11666
rect 29006 11625 29017 11666
rect 29006 11563 29016 11625
rect 29006 11522 29017 11563
rect 28768 11517 29017 11522
rect 28768 11516 28854 11517
rect 28768 11464 28816 11516
rect 29072 11476 29142 11712
rect 29197 11666 29389 11671
rect 29197 11625 29208 11666
rect 29198 11563 29208 11625
rect 29197 11522 29208 11563
rect 29378 11625 29389 11666
rect 29378 11563 29388 11625
rect 29378 11522 29389 11563
rect 29197 11517 29389 11522
rect 29444 11476 29514 11712
rect 29569 11666 29761 11671
rect 29569 11625 29580 11666
rect 29570 11563 29580 11625
rect 29569 11522 29580 11563
rect 29750 11625 29761 11666
rect 29750 11563 29760 11625
rect 29750 11522 29761 11563
rect 29569 11517 29761 11522
rect 29816 11476 29886 11712
rect 29941 11670 30133 11671
rect 30188 11670 30258 11712
rect 30313 11670 30505 11671
rect 29941 11666 30505 11670
rect 29941 11625 29952 11666
rect 29942 11563 29952 11625
rect 29941 11522 29952 11563
rect 30122 11522 30324 11666
rect 30494 11625 30505 11666
rect 30494 11563 30504 11625
rect 30494 11522 30505 11563
rect 29941 11518 30505 11522
rect 29941 11517 30133 11518
rect 30188 11476 30258 11518
rect 30313 11517 30505 11518
rect 30560 11476 30630 11712
rect 30685 11666 30877 11671
rect 30685 11625 30696 11666
rect 30686 11563 30696 11625
rect 30685 11522 30696 11563
rect 30866 11625 30877 11666
rect 30866 11563 30876 11625
rect 30866 11522 30877 11563
rect 30685 11517 30877 11522
rect 30932 11476 31002 11712
rect 31057 11666 31249 11671
rect 31057 11625 31068 11666
rect 31058 11563 31068 11625
rect 31057 11522 31068 11563
rect 31238 11625 31249 11666
rect 31238 11563 31248 11625
rect 31238 11522 31249 11563
rect 31057 11517 31249 11522
rect 31304 11476 31374 11712
rect 31676 11672 31746 11712
rect 31484 11671 31902 11672
rect 31429 11666 31993 11671
rect 31429 11625 31440 11666
rect 31430 11563 31440 11625
rect 31429 11522 31440 11563
rect 31610 11522 31812 11666
rect 31982 11625 31993 11666
rect 31982 11563 31992 11625
rect 31982 11522 31993 11563
rect 31429 11517 31993 11522
rect 31484 11516 31902 11517
rect 31676 11476 31746 11516
rect 32048 11476 32118 11712
rect 32173 11666 32365 11671
rect 32173 11625 32184 11666
rect 32174 11563 32184 11625
rect 32173 11522 32184 11563
rect 32354 11625 32365 11666
rect 32354 11563 32364 11625
rect 32354 11522 32365 11563
rect 32173 11517 32365 11522
rect 32420 11476 32490 11712
rect 32545 11666 32737 11671
rect 32545 11625 32556 11666
rect 32546 11563 32556 11625
rect 32545 11522 32556 11563
rect 32726 11625 32737 11666
rect 32726 11563 32736 11625
rect 32726 11522 32737 11563
rect 32545 11517 32737 11522
rect 32792 11476 32862 11712
rect 33164 11672 33234 11712
rect 33012 11671 33388 11672
rect 32917 11666 33481 11671
rect 32917 11625 32928 11666
rect 32918 11563 32928 11625
rect 32917 11522 32928 11563
rect 33098 11522 33300 11666
rect 33470 11625 33481 11666
rect 33470 11563 33480 11625
rect 33470 11522 33481 11563
rect 32917 11517 33481 11522
rect 33012 11516 33388 11517
rect 33164 11476 33234 11516
rect 33536 11476 33606 11712
rect 33661 11666 33853 11671
rect 33661 11625 33672 11666
rect 33662 11563 33672 11625
rect 33661 11522 33672 11563
rect 33842 11625 33853 11666
rect 33842 11563 33852 11625
rect 33842 11522 33853 11563
rect 33661 11517 33853 11522
rect 33908 11476 33978 11712
rect 34033 11666 34225 11671
rect 34033 11625 34044 11666
rect 34034 11563 34044 11625
rect 34033 11522 34044 11563
rect 34214 11625 34225 11666
rect 34214 11563 34224 11625
rect 34214 11522 34225 11563
rect 34033 11517 34225 11522
rect 34280 11476 34350 11712
rect 34606 11672 34658 11724
rect 34500 11671 34658 11672
rect 34405 11666 34658 11671
rect 34405 11625 34416 11666
rect 34406 11563 34416 11625
rect 34405 11522 34416 11563
rect 34586 11522 34658 11666
rect 34405 11517 34658 11522
rect 34500 11516 34658 11517
rect 28768 11088 28775 11464
rect 28809 11088 28816 11464
rect 28768 11036 28816 11088
rect 29027 11464 29187 11476
rect 29027 11088 29033 11464
rect 29067 11088 29147 11464
rect 29181 11088 29187 11464
rect 29027 11076 29187 11088
rect 29399 11464 29559 11476
rect 29399 11088 29405 11464
rect 29439 11088 29519 11464
rect 29553 11088 29559 11464
rect 29399 11076 29559 11088
rect 29771 11464 29931 11476
rect 29771 11088 29777 11464
rect 29811 11088 29891 11464
rect 29925 11088 29931 11464
rect 29771 11076 29931 11088
rect 30143 11464 30303 11476
rect 30143 11088 30149 11464
rect 30183 11088 30263 11464
rect 30297 11088 30303 11464
rect 30143 11076 30303 11088
rect 30515 11464 30675 11476
rect 30515 11088 30521 11464
rect 30555 11088 30635 11464
rect 30669 11088 30675 11464
rect 30515 11076 30675 11088
rect 30887 11464 31047 11476
rect 30887 11088 30893 11464
rect 30927 11088 31007 11464
rect 31041 11088 31047 11464
rect 30887 11076 31047 11088
rect 31259 11464 31419 11476
rect 31259 11088 31265 11464
rect 31299 11088 31379 11464
rect 31413 11088 31419 11464
rect 31259 11076 31419 11088
rect 31631 11464 31791 11476
rect 31631 11088 31637 11464
rect 31671 11088 31751 11464
rect 31785 11088 31791 11464
rect 31631 11076 31791 11088
rect 32003 11464 32163 11476
rect 32003 11088 32009 11464
rect 32043 11088 32123 11464
rect 32157 11088 32163 11464
rect 32003 11076 32163 11088
rect 32375 11464 32535 11476
rect 32375 11088 32381 11464
rect 32415 11088 32495 11464
rect 32529 11088 32535 11464
rect 32375 11076 32535 11088
rect 32747 11464 32907 11476
rect 32747 11088 32753 11464
rect 32787 11088 32867 11464
rect 32901 11088 32907 11464
rect 32747 11076 32907 11088
rect 33119 11464 33279 11476
rect 33119 11088 33125 11464
rect 33159 11088 33239 11464
rect 33273 11088 33279 11464
rect 33119 11076 33279 11088
rect 33491 11464 33651 11476
rect 33491 11088 33497 11464
rect 33531 11088 33611 11464
rect 33645 11088 33651 11464
rect 33491 11076 33651 11088
rect 33863 11464 34023 11476
rect 33863 11088 33869 11464
rect 33903 11088 33983 11464
rect 34017 11088 34023 11464
rect 33863 11076 34023 11088
rect 34235 11464 34395 11476
rect 34235 11088 34241 11464
rect 34275 11088 34355 11464
rect 34389 11088 34395 11464
rect 34235 11076 34395 11088
rect 34606 11464 34658 11516
rect 34606 11088 34613 11464
rect 34647 11088 34658 11464
rect 28768 11035 28858 11036
rect 28768 11030 29017 11035
rect 28768 10886 28836 11030
rect 29006 10989 29017 11030
rect 29006 10927 29016 10989
rect 29006 10886 29017 10927
rect 28768 10881 29017 10886
rect 28768 10876 28858 10881
rect 28768 10828 28816 10876
rect 29072 10840 29142 11076
rect 29197 11030 29389 11035
rect 29197 10989 29208 11030
rect 29198 10927 29208 10989
rect 29197 10886 29208 10927
rect 29378 10989 29389 11030
rect 29378 10927 29388 10989
rect 29378 10886 29389 10927
rect 29197 10881 29389 10886
rect 29444 10840 29514 11076
rect 29569 11030 29761 11035
rect 29569 10989 29580 11030
rect 29570 10927 29580 10989
rect 29569 10886 29580 10927
rect 29750 10989 29761 11030
rect 29750 10927 29760 10989
rect 29750 10886 29761 10927
rect 29569 10881 29761 10886
rect 29816 10840 29886 11076
rect 29941 11032 30133 11035
rect 30188 11032 30258 11076
rect 30313 11032 30505 11035
rect 29941 11030 30505 11032
rect 29941 10989 29952 11030
rect 29942 10927 29952 10989
rect 29941 10886 29952 10927
rect 30122 10886 30324 11030
rect 30494 10989 30505 11030
rect 30494 10927 30504 10989
rect 30494 10886 30505 10927
rect 29941 10881 30505 10886
rect 29982 10880 30458 10881
rect 30188 10840 30258 10880
rect 30560 10840 30630 11076
rect 30685 11030 30877 11035
rect 30685 10989 30696 11030
rect 30686 10927 30696 10989
rect 30685 10886 30696 10927
rect 30866 10989 30877 11030
rect 30866 10927 30876 10989
rect 30866 10886 30877 10927
rect 30685 10881 30877 10886
rect 30932 10840 31002 11076
rect 31057 11030 31249 11035
rect 31057 10989 31068 11030
rect 31058 10927 31068 10989
rect 31057 10886 31068 10927
rect 31238 10989 31249 11030
rect 31238 10927 31248 10989
rect 31238 10886 31249 10927
rect 31057 10881 31249 10886
rect 31304 10840 31374 11076
rect 31676 11036 31746 11076
rect 31504 11035 31922 11036
rect 31429 11030 31993 11035
rect 31429 10989 31440 11030
rect 31430 10927 31440 10989
rect 31429 10886 31440 10927
rect 31610 10886 31812 11030
rect 31982 10989 31993 11030
rect 31982 10927 31992 10989
rect 31982 10886 31993 10927
rect 31429 10881 31993 10886
rect 31504 10880 31922 10881
rect 31676 10840 31746 10880
rect 32048 10840 32118 11076
rect 32173 11030 32365 11035
rect 32173 10989 32184 11030
rect 32174 10927 32184 10989
rect 32173 10886 32184 10927
rect 32354 10989 32365 11030
rect 32354 10927 32364 10989
rect 32354 10886 32365 10927
rect 32173 10881 32365 10886
rect 32420 10840 32490 11076
rect 32545 11030 32737 11035
rect 32545 10989 32556 11030
rect 32546 10927 32556 10989
rect 32545 10886 32556 10927
rect 32726 10989 32737 11030
rect 32726 10927 32736 10989
rect 32726 10886 32737 10927
rect 32545 10881 32737 10886
rect 32792 10840 32862 11076
rect 33164 11036 33234 11076
rect 33000 11035 33376 11036
rect 32917 11030 33481 11035
rect 32917 10989 32928 11030
rect 32918 10927 32928 10989
rect 32917 10886 32928 10927
rect 33098 10886 33300 11030
rect 33470 10989 33481 11030
rect 33470 10927 33480 10989
rect 33470 10886 33481 10927
rect 32917 10881 33481 10886
rect 33000 10880 33376 10881
rect 33164 10840 33234 10880
rect 33536 10840 33606 11076
rect 33661 11030 33853 11035
rect 33661 10989 33672 11030
rect 33662 10927 33672 10989
rect 33661 10886 33672 10927
rect 33842 10989 33853 11030
rect 33842 10927 33852 10989
rect 33842 10886 33853 10927
rect 33661 10881 33853 10886
rect 33908 10840 33978 11076
rect 34033 11030 34225 11035
rect 34033 10989 34044 11030
rect 34034 10927 34044 10989
rect 34033 10886 34044 10927
rect 34214 10989 34225 11030
rect 34214 10927 34224 10989
rect 34214 10886 34225 10927
rect 34033 10881 34225 10886
rect 34280 10840 34350 11076
rect 34606 11036 34658 11088
rect 34516 11035 34658 11036
rect 34405 11030 34658 11035
rect 34405 10989 34416 11030
rect 34406 10927 34416 10989
rect 34405 10886 34416 10927
rect 34586 10886 34658 11030
rect 34405 10881 34658 10886
rect 34516 10880 34658 10881
rect 28768 10452 28775 10828
rect 28809 10452 28816 10828
rect 28768 10406 28816 10452
rect 29027 10828 29187 10840
rect 29027 10452 29033 10828
rect 29067 10452 29147 10828
rect 29181 10452 29187 10828
rect 29027 10440 29187 10452
rect 29399 10828 29559 10840
rect 29399 10452 29405 10828
rect 29439 10452 29519 10828
rect 29553 10452 29559 10828
rect 29399 10440 29559 10452
rect 29771 10828 29931 10840
rect 29771 10452 29777 10828
rect 29811 10452 29891 10828
rect 29925 10452 29931 10828
rect 29771 10440 29931 10452
rect 30143 10828 30303 10840
rect 30143 10452 30149 10828
rect 30183 10452 30263 10828
rect 30297 10452 30303 10828
rect 30143 10440 30303 10452
rect 30515 10828 30675 10840
rect 30515 10452 30521 10828
rect 30555 10452 30635 10828
rect 30669 10452 30675 10828
rect 30515 10440 30675 10452
rect 30887 10828 31047 10840
rect 30887 10452 30893 10828
rect 30927 10452 31007 10828
rect 31041 10452 31047 10828
rect 30887 10440 31047 10452
rect 31259 10828 31419 10840
rect 31259 10452 31265 10828
rect 31299 10452 31379 10828
rect 31413 10452 31419 10828
rect 31259 10440 31419 10452
rect 31631 10828 31791 10840
rect 31631 10452 31637 10828
rect 31671 10452 31751 10828
rect 31785 10452 31791 10828
rect 31631 10440 31791 10452
rect 32003 10828 32163 10840
rect 32003 10452 32009 10828
rect 32043 10452 32123 10828
rect 32157 10452 32163 10828
rect 32003 10440 32163 10452
rect 32375 10828 32535 10840
rect 32375 10452 32381 10828
rect 32415 10452 32495 10828
rect 32529 10452 32535 10828
rect 32375 10440 32535 10452
rect 32747 10828 32907 10840
rect 32747 10452 32753 10828
rect 32787 10452 32867 10828
rect 32901 10452 32907 10828
rect 32747 10440 32907 10452
rect 33119 10828 33279 10840
rect 33119 10452 33125 10828
rect 33159 10452 33239 10828
rect 33273 10452 33279 10828
rect 33119 10440 33279 10452
rect 33491 10828 33651 10840
rect 33491 10452 33497 10828
rect 33531 10452 33611 10828
rect 33645 10452 33651 10828
rect 33491 10440 33651 10452
rect 33863 10828 34023 10840
rect 33863 10452 33869 10828
rect 33903 10452 33983 10828
rect 34017 10452 34023 10828
rect 33863 10440 34023 10452
rect 34235 10828 34395 10840
rect 34235 10452 34241 10828
rect 34275 10452 34355 10828
rect 34389 10452 34395 10828
rect 34235 10440 34395 10452
rect 34606 10828 34658 10880
rect 34606 10452 34613 10828
rect 34647 10452 34658 10828
rect 28768 10346 28836 10406
rect 29006 10399 29016 10406
rect 29198 10399 29208 10406
rect 29006 10353 29017 10399
rect 29197 10353 29208 10399
rect 29378 10399 29388 10406
rect 29006 10346 29016 10353
rect 29198 10346 29208 10353
rect 29378 10353 29389 10399
rect 29378 10346 29388 10353
rect 29450 10098 29508 10440
rect 30194 10406 30252 10440
rect 29570 10399 29580 10406
rect 29569 10353 29580 10399
rect 29750 10399 29760 10406
rect 29942 10399 29952 10406
rect 29570 10346 29580 10353
rect 29750 10353 29761 10399
rect 29941 10353 29952 10399
rect 29750 10346 29760 10353
rect 29942 10346 29952 10353
rect 30122 10346 30324 10406
rect 30494 10399 30504 10406
rect 30686 10399 30696 10406
rect 30494 10353 30505 10399
rect 30685 10353 30696 10399
rect 30866 10399 30876 10406
rect 30494 10346 30504 10353
rect 30686 10346 30696 10353
rect 30866 10353 30877 10399
rect 30866 10346 30876 10353
rect 30068 10344 30398 10346
rect 30938 10098 30996 10440
rect 31682 10406 31740 10440
rect 31058 10399 31068 10406
rect 31057 10353 31068 10399
rect 31238 10399 31248 10406
rect 31430 10399 31440 10406
rect 31058 10346 31068 10353
rect 31238 10353 31249 10399
rect 31429 10353 31440 10399
rect 31238 10346 31248 10353
rect 31430 10346 31440 10353
rect 31610 10346 31812 10406
rect 31982 10399 31992 10406
rect 32174 10399 32184 10406
rect 31982 10353 31993 10399
rect 32173 10353 32184 10399
rect 32354 10399 32364 10406
rect 31982 10346 31992 10353
rect 32174 10346 32184 10353
rect 32354 10353 32365 10399
rect 32354 10346 32364 10353
rect 32426 10098 32484 10440
rect 33170 10406 33228 10440
rect 32546 10399 32556 10406
rect 32545 10353 32556 10399
rect 32726 10399 32736 10406
rect 32918 10399 32928 10406
rect 32546 10346 32556 10353
rect 32726 10353 32737 10399
rect 32917 10353 32928 10399
rect 32726 10346 32736 10353
rect 32918 10346 32928 10353
rect 33098 10346 33300 10406
rect 33470 10399 33480 10406
rect 33662 10399 33672 10406
rect 33470 10353 33481 10399
rect 33661 10353 33672 10399
rect 33842 10399 33852 10406
rect 33470 10346 33480 10353
rect 33662 10346 33672 10353
rect 33842 10353 33853 10399
rect 33842 10346 33852 10353
rect 33914 10098 33972 10440
rect 34606 10406 34658 10452
rect 34696 12112 34748 12236
rect 34782 12146 34788 12206
rect 34958 12199 34968 12206
rect 35150 12199 35160 12206
rect 34958 12153 34969 12199
rect 35149 12153 35160 12199
rect 35330 12199 35340 12206
rect 34958 12146 34968 12153
rect 35150 12146 35160 12153
rect 35330 12153 35341 12199
rect 35330 12146 35340 12153
rect 35402 12112 35460 12236
rect 35522 12199 35532 12206
rect 35521 12153 35532 12199
rect 35702 12199 35712 12206
rect 35894 12199 35904 12206
rect 35522 12146 35532 12153
rect 35702 12153 35713 12199
rect 35893 12153 35904 12199
rect 36074 12199 36084 12206
rect 35702 12146 35712 12153
rect 35894 12146 35904 12153
rect 36074 12153 36085 12199
rect 36074 12146 36084 12153
rect 36146 12112 36204 12236
rect 36266 12199 36276 12206
rect 36265 12153 36276 12199
rect 36446 12199 36456 12206
rect 36638 12199 36648 12206
rect 36266 12146 36276 12153
rect 36446 12153 36457 12199
rect 36637 12153 36648 12199
rect 36818 12199 36828 12206
rect 36446 12146 36456 12153
rect 36638 12146 36648 12153
rect 36818 12153 36829 12199
rect 36818 12146 36828 12153
rect 36890 12112 36948 12236
rect 37010 12199 37020 12206
rect 37009 12153 37020 12199
rect 37190 12199 37200 12206
rect 37382 12199 37392 12206
rect 37010 12146 37020 12153
rect 37190 12153 37201 12199
rect 37381 12153 37392 12199
rect 37562 12199 37572 12206
rect 37190 12146 37200 12153
rect 37382 12146 37392 12153
rect 37562 12153 37573 12199
rect 37562 12146 37572 12153
rect 37634 12112 37692 12236
rect 37754 12199 37764 12206
rect 37753 12153 37764 12199
rect 37934 12199 37944 12206
rect 38126 12199 38136 12206
rect 37754 12146 37764 12153
rect 37934 12153 37945 12199
rect 38125 12153 38136 12199
rect 38306 12199 38316 12206
rect 37934 12146 37944 12153
rect 38126 12146 38136 12153
rect 38306 12153 38317 12199
rect 38306 12146 38316 12153
rect 38378 12112 38436 12236
rect 38498 12199 38508 12206
rect 38497 12153 38508 12199
rect 38678 12199 38688 12206
rect 38870 12199 38880 12206
rect 38498 12146 38508 12153
rect 38678 12153 38689 12199
rect 38869 12153 38880 12199
rect 39050 12199 39060 12206
rect 38678 12146 38688 12153
rect 38870 12146 38880 12153
rect 39050 12153 39061 12199
rect 39050 12146 39060 12153
rect 39122 12112 39180 12236
rect 39242 12199 39252 12206
rect 39241 12153 39252 12199
rect 39422 12199 39432 12206
rect 39614 12199 39624 12206
rect 39242 12146 39252 12153
rect 39422 12153 39433 12199
rect 39613 12153 39624 12199
rect 39794 12199 39804 12206
rect 39422 12146 39432 12153
rect 39614 12146 39624 12153
rect 39794 12153 39805 12199
rect 39794 12146 39804 12153
rect 39866 12112 39924 12236
rect 39986 12199 39996 12206
rect 39985 12153 39996 12199
rect 40166 12199 40176 12206
rect 40358 12199 40368 12206
rect 39986 12146 39996 12153
rect 40166 12153 40177 12199
rect 40357 12153 40368 12199
rect 40538 12199 40548 12206
rect 40166 12146 40176 12153
rect 40358 12146 40368 12153
rect 40538 12153 40549 12199
rect 40538 12146 40548 12153
rect 40592 12112 40650 12236
rect 34696 12100 34767 12112
rect 34696 11724 34727 12100
rect 34761 11724 34767 12100
rect 34696 11712 34767 11724
rect 34979 12100 35139 12112
rect 34979 11724 34985 12100
rect 35019 11724 35099 12100
rect 35133 11724 35139 12100
rect 34979 11712 35139 11724
rect 35351 12100 35511 12112
rect 35351 11724 35357 12100
rect 35391 11724 35471 12100
rect 35505 11724 35511 12100
rect 35351 11712 35511 11724
rect 35723 12100 35883 12112
rect 35723 11724 35729 12100
rect 35763 11724 35843 12100
rect 35877 11724 35883 12100
rect 35723 11712 35883 11724
rect 36095 12100 36255 12112
rect 36095 11724 36101 12100
rect 36135 11724 36215 12100
rect 36249 11724 36255 12100
rect 36095 11712 36255 11724
rect 36467 12100 36627 12112
rect 36467 11724 36473 12100
rect 36507 11724 36587 12100
rect 36621 11724 36627 12100
rect 36467 11712 36627 11724
rect 36839 12100 36999 12112
rect 36839 11724 36845 12100
rect 36879 11724 36959 12100
rect 36993 11724 36999 12100
rect 36839 11712 36999 11724
rect 37211 12100 37371 12112
rect 37211 11724 37217 12100
rect 37251 11724 37331 12100
rect 37365 11724 37371 12100
rect 37211 11712 37371 11724
rect 37583 12100 37743 12112
rect 37583 11724 37589 12100
rect 37623 11724 37703 12100
rect 37737 11724 37743 12100
rect 37583 11712 37743 11724
rect 37955 12100 38115 12112
rect 37955 11724 37961 12100
rect 37995 11724 38075 12100
rect 38109 11724 38115 12100
rect 37955 11712 38115 11724
rect 38327 12100 38487 12112
rect 38327 11724 38333 12100
rect 38367 11724 38447 12100
rect 38481 11724 38487 12100
rect 38327 11712 38487 11724
rect 38699 12100 38859 12112
rect 38699 11724 38705 12100
rect 38739 11724 38819 12100
rect 38853 11724 38859 12100
rect 38699 11712 38859 11724
rect 39071 12100 39231 12112
rect 39071 11724 39077 12100
rect 39111 11724 39191 12100
rect 39225 11724 39231 12100
rect 39071 11712 39231 11724
rect 39443 12100 39603 12112
rect 39443 11724 39449 12100
rect 39483 11724 39563 12100
rect 39597 11724 39603 12100
rect 39443 11712 39603 11724
rect 39815 12100 39975 12112
rect 39815 11724 39821 12100
rect 39855 11724 39935 12100
rect 39969 11724 39975 12100
rect 39815 11712 39975 11724
rect 40187 12100 40347 12112
rect 40187 11724 40193 12100
rect 40227 11724 40307 12100
rect 40341 11724 40347 12100
rect 40187 11712 40347 11724
rect 40559 12100 40650 12112
rect 40559 11724 40565 12100
rect 40599 11724 40650 12100
rect 40559 11712 40650 11724
rect 34696 11476 34748 11712
rect 34776 11671 34902 11672
rect 34776 11666 34969 11671
rect 34776 11522 34788 11666
rect 34958 11625 34969 11666
rect 34958 11563 34968 11625
rect 34958 11522 34969 11563
rect 34776 11517 34969 11522
rect 34776 11516 34902 11517
rect 35024 11476 35094 11712
rect 35149 11666 35341 11671
rect 35149 11625 35160 11666
rect 35150 11563 35160 11625
rect 35149 11522 35160 11563
rect 35330 11625 35341 11666
rect 35330 11563 35340 11625
rect 35330 11522 35341 11563
rect 35149 11517 35341 11522
rect 35396 11476 35466 11712
rect 35521 11666 35713 11671
rect 35521 11625 35532 11666
rect 35522 11563 35532 11625
rect 35521 11522 35532 11563
rect 35702 11625 35713 11666
rect 35702 11563 35712 11625
rect 35702 11522 35713 11563
rect 35521 11517 35713 11522
rect 35768 11476 35838 11712
rect 35893 11666 36085 11671
rect 35893 11625 35904 11666
rect 35894 11563 35904 11625
rect 35893 11522 35904 11563
rect 36074 11625 36085 11666
rect 36074 11563 36084 11625
rect 36074 11522 36085 11563
rect 35893 11517 36085 11522
rect 36140 11476 36210 11712
rect 36265 11666 36457 11671
rect 36265 11625 36276 11666
rect 36266 11563 36276 11625
rect 36265 11522 36276 11563
rect 36446 11625 36457 11666
rect 36446 11563 36456 11625
rect 36446 11522 36457 11563
rect 36265 11517 36457 11522
rect 36512 11476 36582 11712
rect 36637 11666 36829 11671
rect 36637 11625 36648 11666
rect 36638 11563 36648 11625
rect 36637 11522 36648 11563
rect 36818 11625 36829 11666
rect 36818 11563 36828 11625
rect 36818 11522 36829 11563
rect 36637 11517 36829 11522
rect 36884 11476 36954 11712
rect 37009 11666 37201 11671
rect 37009 11625 37020 11666
rect 37010 11563 37020 11625
rect 37009 11522 37020 11563
rect 37190 11625 37201 11666
rect 37190 11563 37200 11625
rect 37190 11522 37201 11563
rect 37009 11517 37201 11522
rect 37256 11476 37326 11712
rect 37381 11666 37573 11671
rect 37381 11625 37392 11666
rect 37382 11563 37392 11625
rect 37381 11522 37392 11563
rect 37562 11625 37573 11666
rect 37562 11563 37572 11625
rect 37562 11522 37573 11563
rect 37381 11517 37573 11522
rect 37628 11476 37698 11712
rect 37753 11666 37945 11671
rect 37753 11625 37764 11666
rect 37754 11563 37764 11625
rect 37753 11522 37764 11563
rect 37934 11625 37945 11666
rect 37934 11563 37944 11625
rect 37934 11522 37945 11563
rect 37753 11517 37945 11522
rect 38000 11476 38070 11712
rect 38125 11666 38317 11671
rect 38125 11625 38136 11666
rect 38126 11563 38136 11625
rect 38125 11522 38136 11563
rect 38306 11625 38317 11666
rect 38306 11563 38316 11625
rect 38306 11522 38317 11563
rect 38125 11517 38317 11522
rect 38372 11476 38442 11712
rect 38497 11666 38689 11671
rect 38497 11625 38508 11666
rect 38498 11563 38508 11625
rect 38497 11522 38508 11563
rect 38678 11625 38689 11666
rect 38678 11563 38688 11625
rect 38678 11522 38689 11563
rect 38497 11517 38689 11522
rect 38744 11476 38814 11712
rect 38869 11666 39061 11671
rect 38869 11625 38880 11666
rect 38870 11563 38880 11625
rect 38869 11522 38880 11563
rect 39050 11625 39061 11666
rect 39050 11563 39060 11625
rect 39050 11522 39061 11563
rect 38869 11517 39061 11522
rect 39116 11476 39186 11712
rect 39241 11666 39433 11671
rect 39241 11625 39252 11666
rect 39242 11563 39252 11625
rect 39241 11522 39252 11563
rect 39422 11625 39433 11666
rect 39422 11563 39432 11625
rect 39422 11522 39433 11563
rect 39241 11517 39433 11522
rect 39488 11476 39558 11712
rect 39613 11666 39805 11671
rect 39613 11625 39624 11666
rect 39614 11563 39624 11625
rect 39613 11522 39624 11563
rect 39794 11625 39805 11666
rect 39794 11563 39804 11625
rect 39794 11522 39805 11563
rect 39613 11517 39805 11522
rect 39860 11476 39930 11712
rect 39985 11666 40177 11671
rect 39985 11625 39996 11666
rect 39986 11563 39996 11625
rect 39985 11522 39996 11563
rect 40166 11625 40177 11666
rect 40166 11563 40176 11625
rect 40166 11522 40177 11563
rect 39985 11517 40177 11522
rect 40232 11476 40302 11712
rect 40357 11666 40549 11671
rect 40357 11625 40368 11666
rect 40358 11563 40368 11625
rect 40357 11522 40368 11563
rect 40538 11625 40549 11666
rect 40538 11563 40548 11625
rect 40538 11522 40549 11563
rect 40357 11517 40549 11522
rect 40592 11476 40650 11712
rect 34696 11464 34767 11476
rect 34696 11088 34727 11464
rect 34761 11088 34767 11464
rect 34696 11076 34767 11088
rect 34979 11464 35139 11476
rect 34979 11088 34985 11464
rect 35019 11088 35099 11464
rect 35133 11088 35139 11464
rect 34979 11076 35139 11088
rect 35351 11464 35511 11476
rect 35351 11088 35357 11464
rect 35391 11088 35471 11464
rect 35505 11088 35511 11464
rect 35351 11076 35511 11088
rect 35723 11464 35883 11476
rect 35723 11088 35729 11464
rect 35763 11088 35843 11464
rect 35877 11088 35883 11464
rect 35723 11076 35883 11088
rect 36095 11464 36255 11476
rect 36095 11088 36101 11464
rect 36135 11088 36215 11464
rect 36249 11088 36255 11464
rect 36095 11076 36255 11088
rect 36467 11464 36627 11476
rect 36467 11088 36473 11464
rect 36507 11088 36587 11464
rect 36621 11088 36627 11464
rect 36467 11076 36627 11088
rect 36839 11464 36999 11476
rect 36839 11088 36845 11464
rect 36879 11088 36959 11464
rect 36993 11088 36999 11464
rect 36839 11076 36999 11088
rect 37211 11464 37371 11476
rect 37211 11088 37217 11464
rect 37251 11088 37331 11464
rect 37365 11088 37371 11464
rect 37211 11076 37371 11088
rect 37583 11464 37743 11476
rect 37583 11088 37589 11464
rect 37623 11088 37703 11464
rect 37737 11088 37743 11464
rect 37583 11076 37743 11088
rect 37955 11464 38115 11476
rect 37955 11088 37961 11464
rect 37995 11088 38075 11464
rect 38109 11088 38115 11464
rect 37955 11076 38115 11088
rect 38327 11464 38487 11476
rect 38327 11088 38333 11464
rect 38367 11088 38447 11464
rect 38481 11088 38487 11464
rect 38327 11076 38487 11088
rect 38699 11464 38859 11476
rect 38699 11088 38705 11464
rect 38739 11088 38819 11464
rect 38853 11088 38859 11464
rect 38699 11076 38859 11088
rect 39071 11464 39231 11476
rect 39071 11088 39077 11464
rect 39111 11088 39191 11464
rect 39225 11088 39231 11464
rect 39071 11076 39231 11088
rect 39443 11464 39603 11476
rect 39443 11088 39449 11464
rect 39483 11088 39563 11464
rect 39597 11088 39603 11464
rect 39443 11076 39603 11088
rect 39815 11464 39975 11476
rect 39815 11088 39821 11464
rect 39855 11088 39935 11464
rect 39969 11088 39975 11464
rect 39815 11076 39975 11088
rect 40187 11464 40347 11476
rect 40187 11088 40193 11464
rect 40227 11088 40307 11464
rect 40341 11088 40347 11464
rect 40187 11076 40347 11088
rect 40559 11464 40650 11476
rect 40559 11088 40565 11464
rect 40599 11088 40650 11464
rect 40559 11076 40650 11088
rect 34696 10840 34748 11076
rect 34776 11035 34918 11036
rect 34776 11030 34969 11035
rect 34776 10886 34788 11030
rect 34958 10989 34969 11030
rect 34958 10927 34968 10989
rect 34958 10886 34969 10927
rect 34776 10881 34969 10886
rect 34776 10880 34918 10881
rect 35024 10840 35094 11076
rect 35149 11030 35341 11035
rect 35149 10989 35160 11030
rect 35150 10927 35160 10989
rect 35149 10886 35160 10927
rect 35330 10989 35341 11030
rect 35330 10927 35340 10989
rect 35330 10886 35341 10927
rect 35149 10881 35341 10886
rect 35396 10840 35466 11076
rect 35521 11030 35713 11035
rect 35521 10989 35532 11030
rect 35522 10927 35532 10989
rect 35521 10886 35532 10927
rect 35702 10989 35713 11030
rect 35702 10927 35712 10989
rect 35702 10886 35713 10927
rect 35521 10881 35713 10886
rect 35768 10840 35838 11076
rect 35893 11030 36085 11035
rect 35893 10989 35904 11030
rect 35894 10927 35904 10989
rect 35893 10886 35904 10927
rect 36074 10989 36085 11030
rect 36074 10927 36084 10989
rect 36074 10886 36085 10927
rect 35893 10881 36085 10886
rect 36140 10840 36210 11076
rect 36265 11030 36457 11035
rect 36265 10989 36276 11030
rect 36266 10927 36276 10989
rect 36265 10886 36276 10927
rect 36446 10989 36457 11030
rect 36446 10927 36456 10989
rect 36446 10886 36457 10927
rect 36265 10881 36457 10886
rect 36512 10840 36582 11076
rect 36637 11030 36829 11035
rect 36637 10989 36648 11030
rect 36638 10927 36648 10989
rect 36637 10886 36648 10927
rect 36818 10989 36829 11030
rect 36818 10927 36828 10989
rect 36818 10886 36829 10927
rect 36637 10881 36829 10886
rect 36884 10840 36954 11076
rect 37009 11030 37201 11035
rect 37009 10989 37020 11030
rect 37010 10927 37020 10989
rect 37009 10886 37020 10927
rect 37190 10989 37201 11030
rect 37190 10927 37200 10989
rect 37190 10886 37201 10927
rect 37009 10881 37201 10886
rect 37256 10840 37326 11076
rect 37381 11030 37573 11035
rect 37381 10989 37392 11030
rect 37382 10927 37392 10989
rect 37381 10886 37392 10927
rect 37562 10989 37573 11030
rect 37562 10927 37572 10989
rect 37562 10886 37573 10927
rect 37381 10881 37573 10886
rect 37628 10840 37698 11076
rect 37753 11030 37945 11035
rect 37753 10989 37764 11030
rect 37754 10927 37764 10989
rect 37753 10886 37764 10927
rect 37934 10989 37945 11030
rect 37934 10927 37944 10989
rect 37934 10886 37945 10927
rect 37753 10881 37945 10886
rect 38000 10840 38070 11076
rect 38125 11030 38317 11035
rect 38125 10989 38136 11030
rect 38126 10927 38136 10989
rect 38125 10886 38136 10927
rect 38306 10989 38317 11030
rect 38306 10927 38316 10989
rect 38306 10886 38317 10927
rect 38125 10881 38317 10886
rect 38372 10840 38442 11076
rect 38497 11030 38689 11035
rect 38497 10989 38508 11030
rect 38498 10927 38508 10989
rect 38497 10886 38508 10927
rect 38678 10989 38689 11030
rect 38678 10927 38688 10989
rect 38678 10886 38689 10927
rect 38497 10881 38689 10886
rect 38744 10840 38814 11076
rect 38869 11030 39061 11035
rect 38869 10989 38880 11030
rect 38870 10927 38880 10989
rect 38869 10886 38880 10927
rect 39050 10989 39061 11030
rect 39050 10927 39060 10989
rect 39050 10886 39061 10927
rect 38869 10881 39061 10886
rect 39116 10840 39186 11076
rect 39241 11030 39433 11035
rect 39241 10989 39252 11030
rect 39242 10927 39252 10989
rect 39241 10886 39252 10927
rect 39422 10989 39433 11030
rect 39422 10927 39432 10989
rect 39422 10886 39433 10927
rect 39241 10881 39433 10886
rect 39488 10840 39558 11076
rect 39613 11030 39805 11035
rect 39613 10989 39624 11030
rect 39614 10927 39624 10989
rect 39613 10886 39624 10927
rect 39794 10989 39805 11030
rect 39794 10927 39804 10989
rect 39794 10886 39805 10927
rect 39613 10881 39805 10886
rect 39860 10840 39930 11076
rect 39985 11030 40177 11035
rect 39985 10989 39996 11030
rect 39986 10927 39996 10989
rect 39985 10886 39996 10927
rect 40166 10989 40177 11030
rect 40166 10927 40176 10989
rect 40166 10886 40177 10927
rect 39985 10881 40177 10886
rect 40232 10840 40302 11076
rect 40357 11030 40549 11035
rect 40357 10989 40368 11030
rect 40358 10927 40368 10989
rect 40357 10886 40368 10927
rect 40538 10989 40549 11030
rect 40538 10927 40548 10989
rect 40538 10886 40549 10927
rect 40357 10881 40549 10886
rect 40592 10840 40650 11076
rect 34696 10828 34767 10840
rect 34696 10452 34727 10828
rect 34761 10452 34767 10828
rect 34696 10440 34767 10452
rect 34979 10828 35139 10840
rect 34979 10452 34985 10828
rect 35019 10452 35099 10828
rect 35133 10452 35139 10828
rect 34979 10440 35139 10452
rect 35351 10828 35511 10840
rect 35351 10452 35357 10828
rect 35391 10452 35471 10828
rect 35505 10452 35511 10828
rect 35351 10440 35511 10452
rect 35723 10828 35883 10840
rect 35723 10452 35729 10828
rect 35763 10452 35843 10828
rect 35877 10452 35883 10828
rect 35723 10440 35883 10452
rect 36095 10828 36255 10840
rect 36095 10452 36101 10828
rect 36135 10452 36215 10828
rect 36249 10452 36255 10828
rect 36095 10440 36255 10452
rect 36467 10828 36627 10840
rect 36467 10452 36473 10828
rect 36507 10452 36587 10828
rect 36621 10452 36627 10828
rect 36467 10440 36627 10452
rect 36839 10828 36999 10840
rect 36839 10452 36845 10828
rect 36879 10452 36959 10828
rect 36993 10452 36999 10828
rect 36839 10440 36999 10452
rect 37211 10828 37371 10840
rect 37211 10452 37217 10828
rect 37251 10452 37331 10828
rect 37365 10452 37371 10828
rect 37211 10440 37371 10452
rect 37583 10828 37743 10840
rect 37583 10452 37589 10828
rect 37623 10452 37703 10828
rect 37737 10452 37743 10828
rect 37583 10440 37743 10452
rect 37955 10828 38115 10840
rect 37955 10452 37961 10828
rect 37995 10452 38075 10828
rect 38109 10452 38115 10828
rect 37955 10440 38115 10452
rect 38327 10828 38487 10840
rect 38327 10452 38333 10828
rect 38367 10452 38447 10828
rect 38481 10452 38487 10828
rect 38327 10440 38487 10452
rect 38699 10828 38859 10840
rect 38699 10452 38705 10828
rect 38739 10452 38819 10828
rect 38853 10452 38859 10828
rect 38699 10440 38859 10452
rect 39071 10828 39231 10840
rect 39071 10452 39077 10828
rect 39111 10452 39191 10828
rect 39225 10452 39231 10828
rect 39071 10440 39231 10452
rect 39443 10828 39603 10840
rect 39443 10452 39449 10828
rect 39483 10452 39563 10828
rect 39597 10452 39603 10828
rect 39443 10440 39603 10452
rect 39815 10828 39975 10840
rect 39815 10452 39821 10828
rect 39855 10452 39935 10828
rect 39969 10452 39975 10828
rect 39815 10440 39975 10452
rect 40187 10828 40347 10840
rect 40187 10452 40193 10828
rect 40227 10452 40307 10828
rect 40341 10452 40347 10828
rect 40187 10440 40347 10452
rect 40559 10828 40650 10840
rect 40559 10452 40565 10828
rect 40599 10452 40650 10828
rect 40559 10440 40650 10452
rect 34034 10399 34044 10406
rect 34033 10353 34044 10399
rect 34214 10399 34224 10406
rect 34406 10399 34416 10406
rect 34034 10346 34044 10353
rect 34214 10353 34225 10399
rect 34405 10353 34416 10399
rect 34214 10346 34224 10353
rect 34406 10346 34416 10353
rect 34586 10346 34658 10406
rect 34774 10346 34788 10406
rect 34958 10399 34968 10406
rect 34958 10353 34969 10399
rect 34958 10346 34968 10353
rect 29450 10034 33972 10098
rect 35024 10038 35094 10440
rect 35150 10399 35160 10406
rect 35149 10353 35160 10399
rect 35330 10399 35340 10406
rect 35522 10399 35532 10406
rect 35150 10346 35160 10353
rect 35330 10353 35341 10399
rect 35521 10353 35532 10399
rect 35702 10399 35712 10406
rect 35330 10346 35340 10353
rect 35522 10346 35532 10353
rect 35702 10353 35713 10399
rect 35702 10346 35712 10353
rect 35768 10038 35838 10440
rect 35894 10399 35904 10406
rect 35893 10353 35904 10399
rect 36074 10399 36084 10406
rect 36266 10399 36276 10406
rect 35894 10346 35904 10353
rect 36074 10353 36085 10399
rect 36265 10353 36276 10399
rect 36446 10399 36456 10406
rect 36074 10346 36084 10353
rect 36266 10346 36276 10353
rect 36446 10353 36457 10399
rect 36446 10346 36456 10353
rect 36512 10038 36582 10440
rect 36638 10399 36648 10406
rect 36637 10353 36648 10399
rect 36818 10399 36828 10406
rect 37010 10399 37020 10406
rect 36638 10346 36648 10353
rect 36818 10353 36829 10399
rect 37009 10353 37020 10399
rect 37190 10399 37200 10406
rect 36818 10346 36828 10353
rect 37010 10346 37020 10353
rect 37190 10353 37201 10399
rect 37190 10346 37200 10353
rect 37256 10038 37326 10440
rect 37382 10399 37392 10406
rect 37381 10353 37392 10399
rect 37562 10399 37572 10406
rect 37754 10399 37764 10406
rect 37382 10346 37392 10353
rect 37562 10353 37573 10399
rect 37753 10353 37764 10399
rect 37934 10399 37944 10406
rect 37562 10346 37572 10353
rect 37754 10346 37764 10353
rect 37934 10353 37945 10399
rect 37934 10346 37944 10353
rect 38000 10038 38070 10440
rect 38126 10399 38136 10406
rect 38125 10353 38136 10399
rect 38306 10399 38316 10406
rect 38498 10399 38508 10406
rect 38126 10346 38136 10353
rect 38306 10353 38317 10399
rect 38497 10353 38508 10399
rect 38678 10399 38688 10406
rect 38306 10346 38316 10353
rect 38498 10346 38508 10353
rect 38678 10353 38689 10399
rect 38678 10346 38688 10353
rect 38744 10038 38814 10440
rect 38870 10399 38880 10406
rect 38869 10353 38880 10399
rect 39050 10399 39060 10406
rect 39242 10399 39252 10406
rect 38870 10346 38880 10353
rect 39050 10353 39061 10399
rect 39241 10353 39252 10399
rect 39422 10399 39432 10406
rect 39050 10346 39060 10353
rect 39242 10346 39252 10353
rect 39422 10353 39433 10399
rect 39422 10346 39432 10353
rect 39488 10038 39558 10440
rect 39614 10399 39624 10406
rect 39613 10353 39624 10399
rect 39794 10399 39804 10406
rect 39986 10399 39996 10406
rect 39614 10346 39624 10353
rect 39794 10353 39805 10399
rect 39985 10353 39996 10399
rect 40166 10399 40176 10406
rect 39794 10346 39804 10353
rect 39986 10346 39996 10353
rect 40166 10353 40177 10399
rect 40166 10346 40176 10353
rect 40232 10038 40302 10440
rect 40358 10399 40368 10406
rect 40357 10353 40368 10399
rect 40538 10399 40548 10406
rect 40358 10346 40368 10353
rect 40538 10353 40549 10399
rect 40538 10346 40548 10353
rect 30210 9930 30264 10034
rect 30606 9930 30676 10034
rect 30938 9930 30996 10034
rect 31350 9930 31420 10034
rect 31682 9930 31740 10034
rect 32094 9930 32164 10034
rect 32426 9930 32484 10034
rect 32838 9930 32908 10034
rect 33158 9930 33212 10034
rect 30210 9924 30316 9930
rect 30210 9854 30234 9924
rect 30304 9854 30316 9924
rect 30210 9848 30316 9854
rect 30594 9924 30688 9930
rect 30594 9854 30606 9924
rect 30676 9854 30688 9924
rect 30594 9848 30688 9854
rect 30938 9924 31060 9930
rect 30938 9854 30978 9924
rect 31048 9854 31060 9924
rect 30938 9848 31060 9854
rect 31338 9924 31432 9930
rect 31338 9854 31350 9924
rect 31420 9854 31432 9924
rect 31338 9848 31432 9854
rect 31682 9924 31804 9930
rect 31682 9854 31722 9924
rect 31792 9854 31804 9924
rect 31682 9848 31804 9854
rect 32082 9924 32176 9930
rect 32082 9854 32094 9924
rect 32164 9854 32176 9924
rect 32082 9848 32176 9854
rect 32426 9924 32548 9930
rect 32426 9854 32466 9924
rect 32536 9854 32548 9924
rect 32426 9848 32548 9854
rect 32826 9924 32920 9930
rect 32826 9854 32838 9924
rect 32908 9854 32920 9924
rect 32826 9848 32920 9854
rect 33088 9924 33212 9930
rect 33088 9854 33100 9924
rect 33170 9854 33212 9924
rect 33088 9848 33212 9854
rect 30210 9724 30264 9848
rect 30314 9811 30324 9820
rect 30313 9765 30324 9811
rect 30494 9811 30504 9820
rect 30686 9811 30696 9820
rect 30314 9756 30324 9765
rect 30494 9765 30505 9811
rect 30685 9765 30696 9811
rect 30866 9811 30876 9820
rect 30494 9756 30504 9765
rect 30686 9756 30696 9765
rect 30866 9765 30877 9811
rect 30866 9756 30876 9765
rect 30938 9724 30996 9848
rect 31058 9811 31068 9820
rect 31057 9765 31068 9811
rect 31238 9811 31248 9820
rect 31430 9811 31440 9820
rect 31058 9756 31068 9765
rect 31238 9765 31249 9811
rect 31429 9765 31440 9811
rect 31610 9811 31620 9820
rect 31238 9756 31248 9765
rect 31430 9756 31440 9765
rect 31610 9765 31621 9811
rect 31610 9756 31620 9765
rect 31682 9724 31740 9848
rect 31802 9811 31812 9820
rect 31801 9765 31812 9811
rect 31982 9811 31992 9820
rect 32174 9811 32184 9820
rect 31802 9756 31812 9765
rect 31982 9765 31993 9811
rect 32173 9765 32184 9811
rect 32354 9811 32364 9820
rect 31982 9756 31992 9765
rect 32174 9756 32184 9765
rect 32354 9765 32365 9811
rect 32354 9756 32364 9765
rect 32426 9724 32484 9848
rect 32546 9811 32556 9820
rect 32545 9765 32556 9811
rect 32726 9811 32736 9820
rect 32918 9811 32928 9820
rect 32546 9756 32556 9765
rect 32726 9765 32737 9811
rect 32917 9765 32928 9811
rect 33098 9811 33108 9820
rect 32726 9756 32736 9765
rect 32918 9756 32928 9765
rect 33098 9765 33109 9811
rect 33098 9756 33108 9765
rect 33158 9724 33212 9848
rect 34910 9766 34920 10038
rect 35202 9766 35212 10038
rect 35654 9766 35664 10038
rect 35946 9766 35956 10038
rect 36398 9766 36408 10038
rect 36690 9766 36700 10038
rect 37142 9766 37152 10038
rect 37434 9766 37444 10038
rect 37886 9766 37896 10038
rect 38178 9766 38188 10038
rect 38630 9766 38640 10038
rect 38922 9766 38932 10038
rect 39374 9766 39384 10038
rect 39666 9766 39676 10038
rect 40118 9766 40128 10038
rect 40410 9766 40420 10038
rect 30210 9712 30303 9724
rect 30210 8936 30263 9712
rect 30297 8936 30303 9712
rect 30210 8924 30303 8936
rect 30515 9712 30675 9724
rect 30515 8936 30521 9712
rect 30555 8936 30635 9712
rect 30669 8936 30675 9712
rect 30515 8924 30675 8936
rect 30887 9712 31047 9724
rect 30887 8936 30893 9712
rect 30927 8936 31007 9712
rect 31041 8936 31047 9712
rect 30887 8924 31047 8936
rect 31259 9712 31419 9724
rect 31259 8936 31265 9712
rect 31299 8936 31379 9712
rect 31413 8936 31419 9712
rect 31259 8924 31419 8936
rect 31631 9712 31791 9724
rect 31631 8936 31637 9712
rect 31671 8936 31751 9712
rect 31785 8936 31791 9712
rect 31631 8924 31791 8936
rect 32003 9712 32163 9724
rect 32003 8936 32009 9712
rect 32043 8936 32123 9712
rect 32157 8936 32163 9712
rect 32003 8924 32163 8936
rect 32375 9712 32535 9724
rect 32375 8936 32381 9712
rect 32415 8936 32495 9712
rect 32529 8936 32535 9712
rect 32375 8924 32535 8936
rect 32747 9712 32907 9724
rect 32747 8936 32753 9712
rect 32787 8936 32867 9712
rect 32901 8936 32907 9712
rect 32747 8924 32907 8936
rect 33119 9712 33212 9724
rect 33119 8936 33125 9712
rect 33159 8936 33212 9712
rect 33119 8924 33212 8936
rect 30210 8688 30258 8924
rect 30313 8878 30505 8883
rect 30313 8837 30324 8878
rect 30314 8775 30324 8837
rect 30313 8734 30324 8775
rect 30494 8837 30505 8878
rect 30494 8775 30504 8837
rect 30494 8734 30505 8775
rect 30313 8729 30505 8734
rect 30560 8688 30630 8924
rect 30685 8878 30877 8883
rect 30685 8837 30696 8878
rect 30686 8775 30696 8837
rect 30685 8734 30696 8775
rect 30866 8837 30877 8878
rect 30866 8775 30876 8837
rect 30866 8734 30877 8775
rect 30685 8729 30877 8734
rect 30932 8688 31002 8924
rect 31057 8878 31249 8883
rect 31057 8837 31068 8878
rect 31058 8775 31068 8837
rect 31057 8734 31068 8775
rect 31238 8837 31249 8878
rect 31238 8775 31248 8837
rect 31238 8734 31249 8775
rect 31057 8729 31249 8734
rect 31304 8688 31374 8924
rect 31429 8878 31621 8883
rect 31429 8837 31440 8878
rect 31430 8775 31440 8837
rect 31429 8734 31440 8775
rect 31610 8837 31621 8878
rect 31610 8775 31620 8837
rect 31610 8734 31621 8775
rect 31429 8729 31621 8734
rect 31676 8688 31746 8924
rect 31801 8878 31993 8883
rect 31801 8837 31812 8878
rect 31802 8775 31812 8837
rect 31801 8734 31812 8775
rect 31982 8837 31993 8878
rect 31982 8775 31992 8837
rect 31982 8734 31993 8775
rect 31801 8729 31993 8734
rect 32048 8688 32118 8924
rect 32173 8878 32365 8883
rect 32173 8837 32184 8878
rect 32174 8775 32184 8837
rect 32173 8734 32184 8775
rect 32354 8837 32365 8878
rect 32354 8775 32364 8837
rect 32354 8734 32365 8775
rect 32173 8729 32365 8734
rect 32420 8688 32490 8924
rect 32545 8878 32737 8883
rect 32545 8837 32556 8878
rect 32546 8775 32556 8837
rect 32545 8734 32556 8775
rect 32726 8837 32737 8878
rect 32726 8775 32736 8837
rect 32726 8734 32737 8775
rect 32545 8729 32737 8734
rect 32792 8688 32862 8924
rect 32917 8878 33109 8883
rect 32917 8837 32928 8878
rect 32918 8775 32928 8837
rect 32917 8734 32928 8775
rect 33098 8837 33109 8878
rect 33098 8775 33108 8837
rect 33098 8734 33109 8775
rect 32917 8729 33109 8734
rect 33158 8688 33212 8924
rect 30210 8676 30303 8688
rect 30210 7900 30263 8676
rect 30297 7900 30303 8676
rect 30210 7888 30303 7900
rect 30515 8676 30675 8688
rect 30515 7900 30521 8676
rect 30555 7900 30635 8676
rect 30669 7900 30675 8676
rect 30515 7888 30675 7900
rect 30887 8676 31047 8688
rect 30887 7900 30893 8676
rect 30927 7900 31007 8676
rect 31041 7900 31047 8676
rect 30887 7888 31047 7900
rect 31259 8676 31419 8688
rect 31259 7900 31265 8676
rect 31299 7900 31379 8676
rect 31413 7900 31419 8676
rect 31259 7888 31419 7900
rect 31631 8676 31791 8688
rect 31631 7900 31637 8676
rect 31671 7900 31751 8676
rect 31785 7900 31791 8676
rect 31631 7888 31791 7900
rect 32003 8676 32163 8688
rect 32003 7900 32009 8676
rect 32043 7900 32123 8676
rect 32157 7900 32163 8676
rect 32003 7888 32163 7900
rect 32375 8676 32535 8688
rect 32375 7900 32381 8676
rect 32415 7900 32495 8676
rect 32529 7900 32535 8676
rect 32375 7888 32535 7900
rect 32747 8676 32907 8688
rect 32747 7900 32753 8676
rect 32787 7900 32867 8676
rect 32901 7900 32907 8676
rect 32747 7888 32907 7900
rect 33119 8676 33212 8688
rect 33119 7900 33125 8676
rect 33159 7900 33212 8676
rect 33792 8050 33802 8322
rect 34084 8050 34094 8322
rect 33119 7888 33212 7900
rect 30210 7652 30258 7888
rect 30313 7842 30505 7847
rect 30313 7801 30324 7842
rect 30314 7739 30324 7801
rect 30313 7698 30324 7739
rect 30494 7801 30505 7842
rect 30494 7739 30504 7801
rect 30494 7698 30505 7739
rect 30313 7693 30505 7698
rect 30560 7652 30630 7888
rect 30685 7842 30877 7847
rect 30685 7801 30696 7842
rect 30686 7739 30696 7801
rect 30685 7698 30696 7739
rect 30866 7801 30877 7842
rect 30866 7739 30876 7801
rect 30866 7698 30877 7739
rect 30685 7693 30877 7698
rect 30932 7652 31002 7888
rect 31057 7842 31249 7847
rect 31057 7801 31068 7842
rect 31058 7739 31068 7801
rect 31057 7698 31068 7739
rect 31238 7801 31249 7842
rect 31238 7739 31248 7801
rect 31238 7698 31249 7739
rect 31057 7693 31249 7698
rect 31304 7652 31374 7888
rect 31429 7842 31621 7847
rect 31429 7801 31440 7842
rect 31430 7739 31440 7801
rect 31429 7698 31440 7739
rect 31610 7801 31621 7842
rect 31610 7739 31620 7801
rect 31610 7698 31621 7739
rect 31429 7693 31621 7698
rect 31676 7652 31746 7888
rect 31801 7842 31993 7847
rect 31801 7801 31812 7842
rect 31802 7739 31812 7801
rect 31801 7698 31812 7739
rect 31982 7801 31993 7842
rect 31982 7739 31992 7801
rect 31982 7698 31993 7739
rect 31801 7693 31993 7698
rect 32048 7652 32118 7888
rect 32173 7842 32365 7847
rect 32173 7801 32184 7842
rect 32174 7739 32184 7801
rect 32173 7698 32184 7739
rect 32354 7801 32365 7842
rect 32354 7739 32364 7801
rect 32354 7698 32365 7739
rect 32173 7693 32365 7698
rect 32420 7652 32490 7888
rect 32545 7842 32737 7847
rect 32545 7801 32556 7842
rect 32546 7739 32556 7801
rect 32545 7698 32556 7739
rect 32726 7801 32737 7842
rect 32726 7739 32736 7801
rect 32726 7698 32737 7739
rect 32545 7693 32737 7698
rect 32792 7652 32862 7888
rect 32917 7842 33109 7847
rect 32917 7801 32928 7842
rect 32918 7739 32928 7801
rect 32917 7698 32928 7739
rect 33098 7801 33109 7842
rect 33098 7739 33108 7801
rect 33098 7698 33109 7739
rect 32917 7693 33109 7698
rect 33158 7652 33212 7888
rect 30210 7640 30303 7652
rect 30210 6864 30263 7640
rect 30297 6864 30303 7640
rect 30210 6852 30303 6864
rect 30515 7640 30675 7652
rect 30515 6864 30521 7640
rect 30555 6864 30635 7640
rect 30669 6864 30675 7640
rect 30515 6852 30675 6864
rect 30887 7640 31047 7652
rect 30887 6864 30893 7640
rect 30927 6864 31007 7640
rect 31041 6864 31047 7640
rect 30887 6852 31047 6864
rect 31259 7640 31419 7652
rect 31259 6864 31265 7640
rect 31299 6864 31379 7640
rect 31413 6864 31419 7640
rect 31259 6852 31419 6864
rect 31631 7640 31791 7652
rect 31631 6864 31637 7640
rect 31671 6864 31751 7640
rect 31785 6864 31791 7640
rect 31631 6852 31791 6864
rect 32003 7640 32163 7652
rect 32003 6864 32009 7640
rect 32043 6864 32123 7640
rect 32157 6864 32163 7640
rect 32003 6852 32163 6864
rect 32375 7640 32535 7652
rect 32375 6864 32381 7640
rect 32415 6864 32495 7640
rect 32529 6864 32535 7640
rect 32375 6852 32535 6864
rect 32747 7640 32907 7652
rect 32747 6864 32753 7640
rect 32787 6864 32867 7640
rect 32901 6864 32907 7640
rect 32747 6852 32907 6864
rect 33119 7640 33212 7652
rect 33119 6864 33125 7640
rect 33159 6864 33212 7640
rect 33904 7460 33976 8050
rect 33904 7063 33922 7460
rect 33960 7063 33976 7460
rect 34202 7184 34212 7228
rect 34048 7178 34212 7184
rect 34048 7132 34060 7178
rect 34116 7132 34212 7178
rect 34048 7126 34212 7132
rect 34202 7082 34212 7126
rect 34356 7082 34366 7228
rect 33904 7046 33976 7063
rect 33119 6852 33212 6864
rect 30210 6616 30258 6852
rect 30313 6806 30505 6811
rect 30313 6765 30324 6806
rect 30314 6703 30324 6765
rect 30313 6662 30324 6703
rect 30494 6765 30505 6806
rect 30494 6703 30504 6765
rect 30494 6662 30505 6703
rect 30313 6657 30505 6662
rect 30560 6616 30630 6852
rect 30685 6806 30877 6811
rect 30685 6765 30696 6806
rect 30686 6703 30696 6765
rect 30685 6662 30696 6703
rect 30866 6765 30877 6806
rect 30866 6703 30876 6765
rect 30866 6662 30877 6703
rect 30685 6657 30877 6662
rect 30932 6616 31002 6852
rect 31057 6806 31249 6811
rect 31057 6765 31068 6806
rect 31058 6703 31068 6765
rect 31057 6662 31068 6703
rect 31238 6765 31249 6806
rect 31238 6703 31248 6765
rect 31238 6662 31249 6703
rect 31057 6657 31249 6662
rect 31304 6616 31374 6852
rect 31429 6806 31621 6811
rect 31429 6765 31440 6806
rect 31430 6703 31440 6765
rect 31429 6662 31440 6703
rect 31610 6765 31621 6806
rect 31610 6703 31620 6765
rect 31610 6662 31621 6703
rect 31429 6657 31621 6662
rect 31676 6616 31746 6852
rect 31801 6806 31993 6811
rect 31801 6765 31812 6806
rect 31802 6703 31812 6765
rect 31801 6662 31812 6703
rect 31982 6765 31993 6806
rect 31982 6703 31992 6765
rect 31982 6662 31993 6703
rect 31801 6657 31993 6662
rect 32048 6616 32118 6852
rect 32173 6806 32365 6811
rect 32173 6765 32184 6806
rect 32174 6703 32184 6765
rect 32173 6662 32184 6703
rect 32354 6765 32365 6806
rect 32354 6703 32364 6765
rect 32354 6662 32365 6703
rect 32173 6657 32365 6662
rect 32420 6616 32490 6852
rect 32545 6806 32737 6811
rect 32545 6765 32556 6806
rect 32546 6703 32556 6765
rect 32545 6662 32556 6703
rect 32726 6765 32737 6806
rect 32726 6703 32736 6765
rect 32726 6662 32737 6703
rect 32545 6657 32737 6662
rect 32792 6616 32862 6852
rect 32917 6806 33109 6811
rect 32917 6765 32928 6806
rect 32918 6703 32928 6765
rect 32917 6662 32928 6703
rect 33098 6765 33109 6806
rect 33098 6703 33108 6765
rect 33098 6662 33109 6703
rect 32917 6657 33109 6662
rect 33158 6616 33212 6852
rect 34202 6784 34212 6828
rect 34048 6778 34212 6784
rect 30210 6604 30303 6616
rect 30210 5828 30263 6604
rect 30297 5828 30303 6604
rect 30210 5816 30303 5828
rect 30515 6604 30675 6616
rect 30515 5828 30521 6604
rect 30555 5828 30635 6604
rect 30669 5828 30675 6604
rect 30515 5816 30675 5828
rect 30887 6604 31047 6616
rect 30887 5828 30893 6604
rect 30927 5828 31007 6604
rect 31041 5828 31047 6604
rect 30887 5816 31047 5828
rect 31259 6604 31419 6616
rect 31259 5828 31265 6604
rect 31299 5828 31379 6604
rect 31413 5828 31419 6604
rect 31259 5816 31419 5828
rect 31631 6604 31791 6616
rect 31631 5828 31637 6604
rect 31671 5828 31751 6604
rect 31785 5828 31791 6604
rect 31631 5816 31791 5828
rect 32003 6604 32163 6616
rect 32003 5828 32009 6604
rect 32043 5828 32123 6604
rect 32157 5828 32163 6604
rect 32003 5816 32163 5828
rect 32375 6604 32535 6616
rect 32375 5828 32381 6604
rect 32415 5828 32495 6604
rect 32529 5828 32535 6604
rect 32375 5816 32535 5828
rect 32747 6604 32907 6616
rect 32747 5828 32753 6604
rect 32787 5828 32867 6604
rect 32901 5828 32907 6604
rect 32747 5816 32907 5828
rect 33119 6604 33212 6616
rect 33119 5828 33125 6604
rect 33159 5828 33212 6604
rect 33904 6749 33976 6766
rect 33904 6352 33922 6749
rect 33960 6352 33976 6749
rect 34048 6732 34060 6778
rect 34116 6732 34212 6778
rect 34048 6726 34212 6732
rect 34202 6682 34212 6726
rect 34356 6682 34366 6828
rect 34202 6384 34212 6428
rect 33119 5816 33212 5828
rect 30314 5775 30324 5780
rect 30313 5729 30324 5775
rect 30494 5775 30504 5780
rect 30314 5726 30324 5729
rect 30494 5729 30505 5775
rect 30494 5726 30504 5729
rect 30560 5132 30630 5816
rect 30686 5775 30696 5780
rect 30685 5729 30696 5775
rect 30866 5775 30876 5780
rect 31058 5775 31068 5780
rect 30686 5726 30696 5729
rect 30866 5729 30877 5775
rect 31057 5729 31068 5775
rect 31238 5775 31248 5780
rect 30866 5726 30876 5729
rect 31058 5726 31068 5729
rect 31238 5729 31249 5775
rect 31238 5726 31248 5729
rect 31304 5440 31374 5816
rect 31430 5775 31440 5780
rect 31429 5729 31440 5775
rect 31610 5775 31620 5780
rect 31802 5775 31812 5780
rect 31430 5726 31440 5729
rect 31610 5729 31621 5775
rect 31801 5729 31812 5775
rect 31982 5775 31992 5780
rect 31610 5726 31620 5729
rect 31802 5726 31812 5729
rect 31982 5729 31993 5775
rect 31982 5726 31992 5729
rect 32048 5440 32118 5816
rect 32174 5775 32184 5780
rect 32173 5729 32184 5775
rect 32354 5775 32364 5780
rect 32546 5775 32556 5780
rect 32174 5726 32184 5729
rect 32354 5729 32365 5775
rect 32545 5729 32556 5775
rect 32726 5775 32736 5780
rect 32354 5726 32364 5729
rect 32546 5726 32556 5729
rect 32726 5729 32737 5775
rect 32726 5726 32736 5729
rect 31294 5260 31304 5440
rect 32118 5260 32128 5440
rect 30312 5122 30878 5132
rect 30312 5076 30324 5122
rect 30313 5071 30324 5076
rect 30314 5066 30324 5071
rect 30494 5076 30696 5122
rect 30494 5071 30505 5076
rect 30494 5066 30504 5071
rect 30208 5039 30282 5040
rect 30560 5039 30630 5076
rect 30685 5071 30696 5076
rect 30686 5066 30696 5071
rect 30866 5076 30878 5122
rect 31058 5117 31068 5122
rect 30866 5071 30877 5076
rect 31057 5071 31068 5117
rect 31238 5117 31248 5122
rect 30866 5066 30876 5071
rect 31058 5066 31068 5071
rect 31238 5071 31249 5117
rect 31238 5066 31248 5071
rect 30932 5039 31002 5040
rect 31304 5039 31374 5260
rect 31430 5117 31440 5122
rect 31429 5071 31440 5117
rect 31610 5117 31620 5122
rect 31802 5117 31812 5122
rect 31430 5066 31440 5071
rect 31610 5071 31621 5117
rect 31801 5071 31812 5117
rect 31982 5117 31992 5122
rect 31610 5066 31620 5071
rect 31802 5066 31812 5071
rect 31982 5071 31993 5117
rect 31982 5066 31992 5071
rect 31676 5039 31746 5040
rect 32048 5039 32118 5260
rect 32792 5132 32862 5816
rect 32918 5775 32928 5780
rect 32917 5729 32928 5775
rect 33098 5775 33108 5780
rect 32918 5726 32928 5729
rect 33098 5729 33109 5775
rect 33098 5726 33108 5729
rect 33420 5584 33430 5856
rect 33712 5584 33722 5856
rect 32544 5122 33110 5132
rect 32174 5117 32184 5122
rect 32173 5071 32184 5117
rect 32354 5117 32364 5122
rect 32174 5066 32184 5071
rect 32354 5071 32365 5117
rect 32544 5076 32556 5122
rect 32545 5071 32556 5076
rect 32354 5066 32364 5071
rect 32546 5066 32556 5071
rect 32726 5076 32928 5122
rect 32726 5071 32737 5076
rect 32726 5066 32736 5071
rect 32420 5039 32490 5040
rect 32792 5039 32862 5076
rect 32917 5071 32928 5076
rect 32918 5066 32928 5071
rect 33098 5076 33110 5122
rect 33290 5117 33300 5122
rect 33098 5071 33109 5076
rect 33289 5071 33300 5117
rect 33470 5117 33480 5122
rect 33098 5066 33108 5071
rect 33290 5066 33300 5071
rect 33470 5071 33481 5117
rect 33470 5066 33480 5071
rect 33164 5039 33234 5040
rect 33536 5039 33606 5584
rect 33904 5510 33976 6352
rect 34048 6378 34212 6384
rect 34048 6332 34060 6378
rect 34116 6332 34212 6378
rect 34048 6326 34212 6332
rect 34202 6282 34212 6326
rect 34356 6282 34366 6428
rect 34164 5584 34174 5856
rect 34456 5584 34466 5856
rect 34908 5584 34918 5856
rect 35200 5584 35210 5856
rect 35652 5584 35662 5856
rect 35944 5584 35954 5856
rect 36396 5584 36406 5856
rect 36688 5584 36698 5856
rect 37140 5584 37150 5856
rect 37432 5584 37442 5856
rect 37884 5584 37894 5856
rect 38176 5584 38186 5856
rect 38628 5584 38638 5856
rect 38920 5584 38930 5856
rect 33800 5260 33810 5510
rect 34060 5260 34070 5510
rect 33662 5117 33672 5122
rect 33661 5071 33672 5117
rect 33842 5117 33852 5122
rect 34034 5117 34044 5122
rect 33662 5066 33672 5071
rect 33842 5071 33853 5117
rect 34033 5071 34044 5117
rect 34214 5117 34224 5122
rect 33842 5066 33852 5071
rect 34034 5066 34044 5071
rect 34214 5071 34225 5117
rect 34214 5066 34224 5071
rect 33908 5039 33978 5040
rect 34280 5039 34350 5584
rect 34406 5117 34416 5122
rect 34405 5071 34416 5117
rect 34586 5117 34596 5122
rect 34778 5117 34788 5122
rect 34406 5066 34416 5071
rect 34586 5071 34597 5117
rect 34777 5071 34788 5117
rect 34958 5117 34968 5122
rect 34586 5066 34596 5071
rect 34778 5066 34788 5071
rect 34958 5071 34969 5117
rect 34958 5066 34968 5071
rect 34652 5039 34722 5040
rect 35024 5039 35094 5584
rect 35150 5117 35160 5122
rect 35149 5071 35160 5117
rect 35330 5117 35340 5122
rect 35522 5117 35532 5122
rect 35150 5066 35160 5071
rect 35330 5071 35341 5117
rect 35521 5071 35532 5117
rect 35702 5117 35712 5122
rect 35330 5066 35340 5071
rect 35522 5066 35532 5071
rect 35702 5071 35713 5117
rect 35702 5066 35712 5071
rect 35396 5039 35466 5040
rect 35768 5039 35838 5584
rect 35894 5117 35904 5122
rect 35893 5071 35904 5117
rect 36074 5117 36084 5122
rect 36266 5117 36276 5122
rect 35894 5066 35904 5071
rect 36074 5071 36085 5117
rect 36265 5071 36276 5117
rect 36446 5117 36456 5122
rect 36074 5066 36084 5071
rect 36266 5066 36276 5071
rect 36446 5071 36457 5117
rect 36446 5066 36456 5071
rect 36140 5039 36210 5040
rect 36512 5039 36582 5584
rect 36638 5117 36648 5122
rect 36637 5071 36648 5117
rect 36818 5117 36828 5122
rect 37010 5117 37020 5122
rect 36638 5066 36648 5071
rect 36818 5071 36829 5117
rect 37009 5071 37020 5117
rect 37190 5117 37200 5122
rect 36818 5066 36828 5071
rect 37010 5066 37020 5071
rect 37190 5071 37201 5117
rect 37190 5066 37200 5071
rect 36884 5039 36954 5040
rect 37256 5039 37326 5584
rect 37382 5117 37392 5122
rect 37381 5071 37392 5117
rect 37562 5117 37572 5122
rect 37754 5117 37764 5122
rect 37382 5066 37392 5071
rect 37562 5071 37573 5117
rect 37753 5071 37764 5117
rect 37934 5117 37944 5122
rect 37562 5066 37572 5071
rect 37754 5066 37764 5071
rect 37934 5071 37945 5117
rect 37934 5066 37944 5071
rect 37628 5039 37698 5040
rect 38000 5039 38070 5584
rect 38126 5117 38136 5122
rect 38125 5071 38136 5117
rect 38306 5117 38316 5122
rect 38498 5117 38508 5122
rect 38126 5066 38136 5071
rect 38306 5071 38317 5117
rect 38497 5071 38508 5117
rect 38678 5117 38688 5122
rect 38306 5066 38316 5071
rect 38498 5066 38508 5071
rect 38678 5071 38689 5117
rect 38678 5066 38688 5071
rect 38372 5039 38442 5040
rect 38744 5039 38814 5584
rect 38870 5117 38880 5122
rect 38869 5071 38880 5117
rect 39050 5117 39060 5122
rect 38870 5066 38880 5071
rect 39050 5071 39061 5117
rect 39050 5066 39060 5071
rect 39092 5039 39166 5052
rect 30208 5027 30303 5039
rect 30208 4851 30263 5027
rect 30297 4851 30303 5027
rect 30208 4839 30303 4851
rect 30515 5027 30675 5039
rect 30515 4851 30521 5027
rect 30555 4851 30635 5027
rect 30669 4851 30675 5027
rect 30515 4839 30675 4851
rect 30887 5027 31047 5039
rect 30887 4851 30893 5027
rect 30927 4851 31007 5027
rect 31041 4851 31047 5027
rect 30887 4839 31047 4851
rect 31259 5027 31419 5039
rect 31259 4851 31265 5027
rect 31299 4851 31379 5027
rect 31413 4851 31419 5027
rect 31259 4839 31419 4851
rect 31631 5027 31791 5039
rect 31631 4851 31637 5027
rect 31671 4851 31751 5027
rect 31785 4851 31791 5027
rect 31631 4839 31791 4851
rect 32003 5027 32163 5039
rect 32003 4851 32009 5027
rect 32043 4851 32123 5027
rect 32157 4851 32163 5027
rect 32003 4839 32163 4851
rect 32375 5027 32535 5039
rect 32375 4851 32381 5027
rect 32415 4851 32495 5027
rect 32529 4851 32535 5027
rect 32375 4839 32535 4851
rect 32747 5027 32907 5039
rect 32747 4851 32753 5027
rect 32787 4851 32867 5027
rect 32901 4851 32907 5027
rect 32747 4839 32907 4851
rect 33119 5027 33279 5039
rect 33119 4851 33125 5027
rect 33159 4851 33239 5027
rect 33273 4851 33279 5027
rect 33119 4839 33279 4851
rect 33491 5027 33651 5039
rect 33491 4851 33497 5027
rect 33531 4851 33611 5027
rect 33645 4851 33651 5027
rect 33491 4839 33651 4851
rect 33863 5027 34023 5039
rect 33863 4851 33869 5027
rect 33903 4851 33983 5027
rect 34017 4851 34023 5027
rect 33863 4839 34023 4851
rect 34235 5027 34395 5039
rect 34235 4851 34241 5027
rect 34275 4851 34355 5027
rect 34389 4851 34395 5027
rect 34235 4839 34395 4851
rect 34607 5027 34767 5039
rect 34607 4851 34613 5027
rect 34647 4851 34727 5027
rect 34761 4851 34767 5027
rect 34607 4839 34767 4851
rect 34979 5027 35139 5039
rect 34979 4851 34985 5027
rect 35019 4851 35099 5027
rect 35133 4851 35139 5027
rect 34979 4839 35139 4851
rect 35351 5027 35511 5039
rect 35351 4851 35357 5027
rect 35391 4851 35471 5027
rect 35505 4851 35511 5027
rect 35351 4839 35511 4851
rect 35723 5027 35883 5039
rect 35723 4851 35729 5027
rect 35763 4851 35843 5027
rect 35877 4851 35883 5027
rect 35723 4839 35883 4851
rect 36095 5027 36255 5039
rect 36095 4851 36101 5027
rect 36135 4851 36215 5027
rect 36249 4851 36255 5027
rect 36095 4839 36255 4851
rect 36467 5027 36627 5039
rect 36467 4851 36473 5027
rect 36507 4851 36587 5027
rect 36621 4851 36627 5027
rect 36467 4839 36627 4851
rect 36839 5027 36999 5039
rect 36839 4851 36845 5027
rect 36879 4851 36959 5027
rect 36993 4851 36999 5027
rect 36839 4839 36999 4851
rect 37211 5027 37371 5039
rect 37211 4851 37217 5027
rect 37251 4851 37331 5027
rect 37365 4851 37371 5027
rect 37211 4839 37371 4851
rect 37583 5027 37743 5039
rect 37583 4851 37589 5027
rect 37623 4851 37703 5027
rect 37737 4851 37743 5027
rect 37583 4839 37743 4851
rect 37955 5027 38115 5039
rect 37955 4851 37961 5027
rect 37995 4851 38075 5027
rect 38109 4851 38115 5027
rect 37955 4839 38115 4851
rect 38327 5027 38487 5039
rect 38327 4851 38333 5027
rect 38367 4851 38447 5027
rect 38481 4851 38487 5027
rect 38327 4839 38487 4851
rect 38699 5027 38859 5039
rect 38699 4851 38705 5027
rect 38739 4851 38819 5027
rect 38853 4851 38859 5027
rect 38699 4839 38859 4851
rect 39071 5027 39166 5039
rect 39071 4851 39077 5027
rect 39111 4851 39166 5027
rect 39071 4839 39166 4851
rect 30208 4621 30282 4839
rect 30560 4808 30630 4839
rect 30312 4802 30878 4808
rect 30312 4658 30324 4802
rect 30494 4658 30696 4802
rect 30866 4658 30878 4802
rect 30312 4652 30878 4658
rect 30560 4621 30630 4652
rect 30932 4621 31002 4839
rect 31057 4802 31249 4807
rect 31057 4761 31068 4802
rect 31058 4699 31068 4761
rect 31057 4658 31068 4699
rect 31238 4761 31249 4802
rect 31238 4699 31248 4761
rect 31238 4658 31249 4699
rect 31057 4653 31249 4658
rect 31304 4621 31374 4839
rect 31429 4802 31621 4807
rect 31429 4761 31440 4802
rect 31430 4699 31440 4761
rect 31429 4658 31440 4699
rect 31610 4761 31621 4802
rect 31610 4699 31620 4761
rect 31610 4658 31621 4699
rect 31429 4653 31621 4658
rect 31676 4621 31746 4839
rect 31801 4802 31993 4807
rect 31801 4761 31812 4802
rect 31802 4699 31812 4761
rect 31801 4658 31812 4699
rect 31982 4761 31993 4802
rect 31982 4699 31992 4761
rect 31982 4658 31993 4699
rect 31801 4653 31993 4658
rect 32048 4621 32118 4839
rect 32173 4802 32365 4807
rect 32173 4761 32184 4802
rect 32174 4699 32184 4761
rect 32173 4658 32184 4699
rect 32354 4761 32365 4802
rect 32354 4699 32364 4761
rect 32354 4658 32365 4699
rect 32173 4653 32365 4658
rect 32420 4621 32490 4839
rect 32792 4808 32862 4839
rect 32544 4802 33110 4808
rect 32544 4658 32556 4802
rect 32726 4658 32928 4802
rect 33098 4658 33110 4802
rect 32544 4652 33110 4658
rect 32792 4621 32862 4652
rect 33164 4621 33234 4839
rect 33289 4802 33481 4807
rect 33289 4761 33300 4802
rect 33290 4699 33300 4761
rect 33289 4658 33300 4699
rect 33470 4761 33481 4802
rect 33470 4699 33480 4761
rect 33470 4658 33481 4699
rect 33289 4653 33481 4658
rect 33536 4621 33606 4839
rect 33661 4802 33853 4807
rect 33661 4761 33672 4802
rect 33662 4699 33672 4761
rect 33661 4658 33672 4699
rect 33842 4761 33853 4802
rect 33842 4699 33852 4761
rect 33842 4658 33853 4699
rect 33661 4653 33853 4658
rect 33908 4621 33978 4839
rect 34033 4802 34225 4807
rect 34033 4761 34044 4802
rect 34034 4699 34044 4761
rect 34033 4658 34044 4699
rect 34214 4761 34225 4802
rect 34214 4699 34224 4761
rect 34214 4658 34225 4699
rect 34033 4653 34225 4658
rect 34280 4621 34350 4839
rect 34405 4802 34597 4807
rect 34405 4761 34416 4802
rect 34406 4699 34416 4761
rect 34405 4658 34416 4699
rect 34586 4761 34597 4802
rect 34586 4699 34596 4761
rect 34586 4658 34597 4699
rect 34405 4653 34597 4658
rect 34652 4621 34722 4839
rect 34777 4802 34969 4807
rect 34777 4761 34788 4802
rect 34778 4699 34788 4761
rect 34777 4658 34788 4699
rect 34958 4761 34969 4802
rect 34958 4699 34968 4761
rect 34958 4658 34969 4699
rect 34777 4653 34969 4658
rect 35024 4621 35094 4839
rect 35149 4802 35341 4807
rect 35149 4761 35160 4802
rect 35150 4699 35160 4761
rect 35149 4658 35160 4699
rect 35330 4761 35341 4802
rect 35330 4699 35340 4761
rect 35330 4658 35341 4699
rect 35149 4653 35341 4658
rect 35396 4621 35466 4839
rect 35521 4802 35713 4807
rect 35521 4761 35532 4802
rect 35522 4699 35532 4761
rect 35521 4658 35532 4699
rect 35702 4761 35713 4802
rect 35702 4699 35712 4761
rect 35702 4658 35713 4699
rect 35521 4653 35713 4658
rect 35768 4621 35838 4839
rect 35893 4802 36085 4807
rect 35893 4761 35904 4802
rect 35894 4699 35904 4761
rect 35893 4658 35904 4699
rect 36074 4761 36085 4802
rect 36074 4699 36084 4761
rect 36074 4658 36085 4699
rect 35893 4653 36085 4658
rect 36140 4621 36210 4839
rect 36265 4802 36457 4807
rect 36265 4761 36276 4802
rect 36266 4699 36276 4761
rect 36265 4658 36276 4699
rect 36446 4761 36457 4802
rect 36446 4699 36456 4761
rect 36446 4658 36457 4699
rect 36265 4653 36457 4658
rect 36512 4621 36582 4839
rect 36637 4802 36829 4807
rect 36637 4761 36648 4802
rect 36638 4699 36648 4761
rect 36637 4658 36648 4699
rect 36818 4761 36829 4802
rect 36818 4699 36828 4761
rect 36818 4658 36829 4699
rect 36637 4653 36829 4658
rect 36884 4621 36954 4839
rect 37009 4802 37201 4807
rect 37009 4761 37020 4802
rect 37010 4699 37020 4761
rect 37009 4658 37020 4699
rect 37190 4761 37201 4802
rect 37190 4699 37200 4761
rect 37190 4658 37201 4699
rect 37009 4653 37201 4658
rect 37256 4621 37326 4839
rect 37381 4802 37573 4807
rect 37381 4761 37392 4802
rect 37382 4699 37392 4761
rect 37381 4658 37392 4699
rect 37562 4761 37573 4802
rect 37562 4699 37572 4761
rect 37562 4658 37573 4699
rect 37381 4653 37573 4658
rect 37628 4621 37698 4839
rect 37753 4802 37945 4807
rect 37753 4761 37764 4802
rect 37754 4699 37764 4761
rect 37753 4658 37764 4699
rect 37934 4761 37945 4802
rect 37934 4699 37944 4761
rect 37934 4658 37945 4699
rect 37753 4653 37945 4658
rect 38000 4621 38070 4839
rect 38125 4802 38317 4807
rect 38125 4761 38136 4802
rect 38126 4699 38136 4761
rect 38125 4658 38136 4699
rect 38306 4761 38317 4802
rect 38306 4699 38316 4761
rect 38306 4658 38317 4699
rect 38125 4653 38317 4658
rect 38372 4621 38442 4839
rect 38497 4802 38689 4807
rect 38497 4761 38508 4802
rect 38498 4699 38508 4761
rect 38497 4658 38508 4699
rect 38678 4761 38689 4802
rect 38678 4699 38688 4761
rect 38678 4658 38689 4699
rect 38497 4653 38689 4658
rect 38744 4621 38814 4839
rect 38869 4802 39061 4807
rect 38869 4761 38880 4802
rect 38870 4699 38880 4761
rect 38869 4658 38880 4699
rect 39050 4761 39061 4802
rect 39050 4699 39060 4761
rect 39050 4658 39061 4699
rect 38869 4653 39061 4658
rect 39092 4621 39166 4839
rect 30208 4609 30303 4621
rect 30208 4433 30263 4609
rect 30297 4433 30303 4609
rect 30208 4421 30303 4433
rect 30515 4609 30675 4621
rect 30515 4433 30521 4609
rect 30555 4433 30635 4609
rect 30669 4433 30675 4609
rect 30515 4421 30675 4433
rect 30887 4609 31047 4621
rect 30887 4433 30893 4609
rect 30927 4433 31007 4609
rect 31041 4433 31047 4609
rect 30887 4421 31047 4433
rect 31259 4609 31419 4621
rect 31259 4433 31265 4609
rect 31299 4433 31379 4609
rect 31413 4433 31419 4609
rect 31259 4421 31419 4433
rect 31631 4609 31791 4621
rect 31631 4433 31637 4609
rect 31671 4433 31751 4609
rect 31785 4433 31791 4609
rect 31631 4421 31791 4433
rect 32003 4609 32163 4621
rect 32003 4433 32009 4609
rect 32043 4433 32123 4609
rect 32157 4433 32163 4609
rect 32003 4421 32163 4433
rect 32375 4609 32535 4621
rect 32375 4433 32381 4609
rect 32415 4433 32495 4609
rect 32529 4433 32535 4609
rect 32375 4421 32535 4433
rect 32747 4609 32907 4621
rect 32747 4433 32753 4609
rect 32787 4433 32867 4609
rect 32901 4433 32907 4609
rect 32747 4421 32907 4433
rect 33119 4609 33279 4621
rect 33119 4433 33125 4609
rect 33159 4433 33239 4609
rect 33273 4433 33279 4609
rect 33119 4421 33279 4433
rect 33491 4609 33651 4621
rect 33491 4433 33497 4609
rect 33531 4433 33611 4609
rect 33645 4433 33651 4609
rect 33491 4421 33651 4433
rect 33863 4609 34023 4621
rect 33863 4433 33869 4609
rect 33903 4433 33983 4609
rect 34017 4433 34023 4609
rect 33863 4421 34023 4433
rect 34235 4609 34395 4621
rect 34235 4433 34241 4609
rect 34275 4433 34355 4609
rect 34389 4433 34395 4609
rect 34235 4421 34395 4433
rect 34607 4609 34767 4621
rect 34607 4433 34613 4609
rect 34647 4433 34727 4609
rect 34761 4433 34767 4609
rect 34607 4421 34767 4433
rect 34979 4609 35139 4621
rect 34979 4433 34985 4609
rect 35019 4433 35099 4609
rect 35133 4433 35139 4609
rect 34979 4421 35139 4433
rect 35351 4609 35511 4621
rect 35351 4433 35357 4609
rect 35391 4433 35471 4609
rect 35505 4433 35511 4609
rect 35351 4421 35511 4433
rect 35723 4609 35883 4621
rect 35723 4433 35729 4609
rect 35763 4433 35843 4609
rect 35877 4433 35883 4609
rect 35723 4421 35883 4433
rect 36095 4609 36255 4621
rect 36095 4433 36101 4609
rect 36135 4433 36215 4609
rect 36249 4433 36255 4609
rect 36095 4421 36255 4433
rect 36467 4609 36627 4621
rect 36467 4433 36473 4609
rect 36507 4433 36587 4609
rect 36621 4433 36627 4609
rect 36467 4421 36627 4433
rect 36839 4609 36999 4621
rect 36839 4433 36845 4609
rect 36879 4433 36959 4609
rect 36993 4433 36999 4609
rect 36839 4421 36999 4433
rect 37211 4609 37371 4621
rect 37211 4433 37217 4609
rect 37251 4433 37331 4609
rect 37365 4433 37371 4609
rect 37211 4421 37371 4433
rect 37583 4609 37743 4621
rect 37583 4433 37589 4609
rect 37623 4433 37703 4609
rect 37737 4433 37743 4609
rect 37583 4421 37743 4433
rect 37955 4609 38115 4621
rect 37955 4433 37961 4609
rect 37995 4433 38075 4609
rect 38109 4433 38115 4609
rect 37955 4421 38115 4433
rect 38327 4609 38487 4621
rect 38327 4433 38333 4609
rect 38367 4433 38447 4609
rect 38481 4433 38487 4609
rect 38327 4421 38487 4433
rect 38699 4609 38859 4621
rect 38699 4433 38705 4609
rect 38739 4433 38819 4609
rect 38853 4433 38859 4609
rect 38699 4421 38859 4433
rect 39071 4609 39166 4621
rect 39071 4433 39077 4609
rect 39111 4433 39166 4609
rect 39071 4421 39166 4433
rect 30208 4203 30282 4421
rect 30560 4390 30630 4421
rect 30312 4384 30878 4390
rect 30312 4240 30324 4384
rect 30494 4240 30696 4384
rect 30866 4240 30878 4384
rect 30312 4234 30878 4240
rect 30560 4203 30630 4234
rect 30932 4203 31002 4421
rect 31057 4384 31249 4389
rect 31057 4343 31068 4384
rect 31058 4281 31068 4343
rect 31057 4240 31068 4281
rect 31238 4343 31249 4384
rect 31238 4281 31248 4343
rect 31238 4240 31249 4281
rect 31057 4235 31249 4240
rect 31304 4203 31374 4421
rect 31429 4384 31621 4389
rect 31429 4343 31440 4384
rect 31430 4281 31440 4343
rect 31429 4240 31440 4281
rect 31610 4343 31621 4384
rect 31610 4281 31620 4343
rect 31610 4240 31621 4281
rect 31429 4235 31621 4240
rect 31676 4203 31746 4421
rect 31801 4384 31993 4389
rect 31801 4343 31812 4384
rect 31802 4281 31812 4343
rect 31801 4240 31812 4281
rect 31982 4343 31993 4384
rect 31982 4281 31992 4343
rect 31982 4240 31993 4281
rect 31801 4235 31993 4240
rect 32048 4203 32118 4421
rect 32173 4384 32365 4389
rect 32173 4343 32184 4384
rect 32174 4281 32184 4343
rect 32173 4240 32184 4281
rect 32354 4343 32365 4384
rect 32354 4281 32364 4343
rect 32354 4240 32365 4281
rect 32173 4235 32365 4240
rect 32420 4203 32490 4421
rect 32792 4390 32862 4421
rect 32544 4384 33110 4390
rect 32544 4240 32556 4384
rect 32726 4240 32928 4384
rect 33098 4240 33110 4384
rect 32544 4234 33110 4240
rect 32792 4203 32862 4234
rect 33164 4203 33234 4421
rect 33289 4384 33481 4389
rect 33289 4343 33300 4384
rect 33290 4281 33300 4343
rect 33289 4240 33300 4281
rect 33470 4343 33481 4384
rect 33470 4281 33480 4343
rect 33470 4240 33481 4281
rect 33289 4235 33481 4240
rect 33536 4203 33606 4421
rect 33661 4384 33853 4389
rect 33661 4343 33672 4384
rect 33662 4281 33672 4343
rect 33661 4240 33672 4281
rect 33842 4343 33853 4384
rect 33842 4281 33852 4343
rect 33842 4240 33853 4281
rect 33661 4235 33853 4240
rect 33908 4203 33978 4421
rect 34033 4384 34225 4389
rect 34033 4343 34044 4384
rect 34034 4281 34044 4343
rect 34033 4240 34044 4281
rect 34214 4343 34225 4384
rect 34214 4281 34224 4343
rect 34214 4240 34225 4281
rect 34033 4235 34225 4240
rect 34280 4203 34350 4421
rect 34405 4384 34597 4389
rect 34405 4343 34416 4384
rect 34406 4281 34416 4343
rect 34405 4240 34416 4281
rect 34586 4343 34597 4384
rect 34586 4281 34596 4343
rect 34586 4240 34597 4281
rect 34405 4235 34597 4240
rect 34652 4203 34722 4421
rect 34777 4384 34969 4389
rect 34777 4343 34788 4384
rect 34778 4281 34788 4343
rect 34777 4240 34788 4281
rect 34958 4343 34969 4384
rect 34958 4281 34968 4343
rect 34958 4240 34969 4281
rect 34777 4235 34969 4240
rect 35024 4203 35094 4421
rect 35149 4384 35341 4389
rect 35149 4343 35160 4384
rect 35150 4281 35160 4343
rect 35149 4240 35160 4281
rect 35330 4343 35341 4384
rect 35330 4281 35340 4343
rect 35330 4240 35341 4281
rect 35149 4235 35341 4240
rect 35396 4203 35466 4421
rect 35521 4384 35713 4389
rect 35521 4343 35532 4384
rect 35522 4281 35532 4343
rect 35521 4240 35532 4281
rect 35702 4343 35713 4384
rect 35702 4281 35712 4343
rect 35702 4240 35713 4281
rect 35521 4235 35713 4240
rect 35768 4203 35838 4421
rect 35893 4384 36085 4389
rect 35893 4343 35904 4384
rect 35894 4281 35904 4343
rect 35893 4240 35904 4281
rect 36074 4343 36085 4384
rect 36074 4281 36084 4343
rect 36074 4240 36085 4281
rect 35893 4235 36085 4240
rect 36140 4203 36210 4421
rect 36265 4384 36457 4389
rect 36265 4343 36276 4384
rect 36266 4281 36276 4343
rect 36265 4240 36276 4281
rect 36446 4343 36457 4384
rect 36446 4281 36456 4343
rect 36446 4240 36457 4281
rect 36265 4235 36457 4240
rect 36512 4203 36582 4421
rect 36637 4384 36829 4389
rect 36637 4343 36648 4384
rect 36638 4281 36648 4343
rect 36637 4240 36648 4281
rect 36818 4343 36829 4384
rect 36818 4281 36828 4343
rect 36818 4240 36829 4281
rect 36637 4235 36829 4240
rect 36884 4203 36954 4421
rect 37009 4384 37201 4389
rect 37009 4343 37020 4384
rect 37010 4281 37020 4343
rect 37009 4240 37020 4281
rect 37190 4343 37201 4384
rect 37190 4281 37200 4343
rect 37190 4240 37201 4281
rect 37009 4235 37201 4240
rect 37256 4203 37326 4421
rect 37381 4384 37573 4389
rect 37381 4343 37392 4384
rect 37382 4281 37392 4343
rect 37381 4240 37392 4281
rect 37562 4343 37573 4384
rect 37562 4281 37572 4343
rect 37562 4240 37573 4281
rect 37381 4235 37573 4240
rect 37628 4203 37698 4421
rect 37753 4384 37945 4389
rect 37753 4343 37764 4384
rect 37754 4281 37764 4343
rect 37753 4240 37764 4281
rect 37934 4343 37945 4384
rect 37934 4281 37944 4343
rect 37934 4240 37945 4281
rect 37753 4235 37945 4240
rect 38000 4203 38070 4421
rect 38125 4384 38317 4389
rect 38125 4343 38136 4384
rect 38126 4281 38136 4343
rect 38125 4240 38136 4281
rect 38306 4343 38317 4384
rect 38306 4281 38316 4343
rect 38306 4240 38317 4281
rect 38125 4235 38317 4240
rect 38372 4203 38442 4421
rect 38497 4384 38689 4389
rect 38497 4343 38508 4384
rect 38498 4281 38508 4343
rect 38497 4240 38508 4281
rect 38678 4343 38689 4384
rect 38678 4281 38688 4343
rect 38678 4240 38689 4281
rect 38497 4235 38689 4240
rect 38744 4203 38814 4421
rect 38869 4384 39061 4389
rect 38869 4343 38880 4384
rect 38870 4281 38880 4343
rect 38869 4240 38880 4281
rect 39050 4343 39061 4384
rect 39050 4281 39060 4343
rect 39050 4240 39061 4281
rect 38869 4235 39061 4240
rect 39092 4203 39166 4421
rect 30208 4191 30303 4203
rect 30208 4015 30263 4191
rect 30297 4015 30303 4191
rect 30208 4003 30303 4015
rect 30515 4191 30675 4203
rect 30515 4015 30521 4191
rect 30555 4015 30635 4191
rect 30669 4015 30675 4191
rect 30515 4003 30675 4015
rect 30887 4191 31047 4203
rect 30887 4015 30893 4191
rect 30927 4015 31007 4191
rect 31041 4015 31047 4191
rect 30887 4003 31047 4015
rect 31259 4191 31419 4203
rect 31259 4015 31265 4191
rect 31299 4015 31379 4191
rect 31413 4015 31419 4191
rect 31259 4003 31419 4015
rect 31631 4191 31791 4203
rect 31631 4015 31637 4191
rect 31671 4015 31751 4191
rect 31785 4015 31791 4191
rect 31631 4003 31791 4015
rect 32003 4191 32163 4203
rect 32003 4015 32009 4191
rect 32043 4015 32123 4191
rect 32157 4015 32163 4191
rect 32003 4003 32163 4015
rect 32375 4191 32535 4203
rect 32375 4015 32381 4191
rect 32415 4015 32495 4191
rect 32529 4015 32535 4191
rect 32375 4003 32535 4015
rect 32747 4191 32907 4203
rect 32747 4015 32753 4191
rect 32787 4015 32867 4191
rect 32901 4015 32907 4191
rect 32747 4003 32907 4015
rect 33119 4191 33279 4203
rect 33119 4015 33125 4191
rect 33159 4015 33239 4191
rect 33273 4015 33279 4191
rect 33119 4003 33279 4015
rect 33491 4191 33651 4203
rect 33491 4015 33497 4191
rect 33531 4015 33611 4191
rect 33645 4015 33651 4191
rect 33491 4003 33651 4015
rect 33863 4191 34023 4203
rect 33863 4015 33869 4191
rect 33903 4015 33983 4191
rect 34017 4015 34023 4191
rect 33863 4003 34023 4015
rect 34235 4191 34395 4203
rect 34235 4015 34241 4191
rect 34275 4015 34355 4191
rect 34389 4015 34395 4191
rect 34235 4003 34395 4015
rect 34607 4191 34767 4203
rect 34607 4015 34613 4191
rect 34647 4015 34727 4191
rect 34761 4015 34767 4191
rect 34607 4003 34767 4015
rect 34979 4191 35139 4203
rect 34979 4015 34985 4191
rect 35019 4015 35099 4191
rect 35133 4015 35139 4191
rect 34979 4003 35139 4015
rect 35351 4191 35511 4203
rect 35351 4015 35357 4191
rect 35391 4015 35471 4191
rect 35505 4015 35511 4191
rect 35351 4003 35511 4015
rect 35723 4191 35883 4203
rect 35723 4015 35729 4191
rect 35763 4015 35843 4191
rect 35877 4015 35883 4191
rect 35723 4003 35883 4015
rect 36095 4191 36255 4203
rect 36095 4015 36101 4191
rect 36135 4015 36215 4191
rect 36249 4015 36255 4191
rect 36095 4003 36255 4015
rect 36467 4191 36627 4203
rect 36467 4015 36473 4191
rect 36507 4015 36587 4191
rect 36621 4015 36627 4191
rect 36467 4003 36627 4015
rect 36839 4191 36999 4203
rect 36839 4015 36845 4191
rect 36879 4015 36959 4191
rect 36993 4015 36999 4191
rect 36839 4003 36999 4015
rect 37211 4191 37371 4203
rect 37211 4015 37217 4191
rect 37251 4015 37331 4191
rect 37365 4015 37371 4191
rect 37211 4003 37371 4015
rect 37583 4191 37743 4203
rect 37583 4015 37589 4191
rect 37623 4015 37703 4191
rect 37737 4015 37743 4191
rect 37583 4003 37743 4015
rect 37955 4191 38115 4203
rect 37955 4015 37961 4191
rect 37995 4015 38075 4191
rect 38109 4015 38115 4191
rect 37955 4003 38115 4015
rect 38327 4191 38487 4203
rect 38327 4015 38333 4191
rect 38367 4015 38447 4191
rect 38481 4015 38487 4191
rect 38327 4003 38487 4015
rect 38699 4191 38859 4203
rect 38699 4015 38705 4191
rect 38739 4015 38819 4191
rect 38853 4015 38859 4191
rect 38699 4003 38859 4015
rect 39071 4191 39166 4203
rect 39071 4015 39077 4191
rect 39111 4015 39166 4191
rect 39071 4003 39166 4015
rect 30208 3785 30282 4003
rect 30560 3972 30630 4003
rect 30312 3966 30878 3972
rect 30312 3822 30324 3966
rect 30494 3822 30696 3966
rect 30866 3822 30878 3966
rect 30312 3816 30878 3822
rect 30560 3785 30630 3816
rect 30932 3785 31002 4003
rect 31057 3966 31249 3971
rect 31057 3925 31068 3966
rect 31058 3863 31068 3925
rect 31057 3822 31068 3863
rect 31238 3925 31249 3966
rect 31238 3863 31248 3925
rect 31238 3822 31249 3863
rect 31057 3817 31249 3822
rect 31304 3785 31374 4003
rect 31429 3966 31621 3971
rect 31429 3925 31440 3966
rect 31430 3863 31440 3925
rect 31429 3822 31440 3863
rect 31610 3925 31621 3966
rect 31610 3863 31620 3925
rect 31610 3822 31621 3863
rect 31429 3817 31621 3822
rect 31676 3785 31746 4003
rect 31801 3966 31993 3971
rect 31801 3925 31812 3966
rect 31802 3863 31812 3925
rect 31801 3822 31812 3863
rect 31982 3925 31993 3966
rect 31982 3863 31992 3925
rect 31982 3822 31993 3863
rect 31801 3817 31993 3822
rect 32048 3785 32118 4003
rect 32173 3966 32365 3971
rect 32173 3925 32184 3966
rect 32174 3863 32184 3925
rect 32173 3822 32184 3863
rect 32354 3925 32365 3966
rect 32354 3863 32364 3925
rect 32354 3822 32365 3863
rect 32173 3817 32365 3822
rect 32420 3785 32490 4003
rect 32792 3972 32862 4003
rect 32544 3966 33110 3972
rect 32544 3822 32556 3966
rect 32726 3822 32928 3966
rect 33098 3822 33110 3966
rect 32544 3816 33110 3822
rect 32792 3785 32862 3816
rect 33164 3785 33234 4003
rect 33289 3966 33481 3971
rect 33289 3925 33300 3966
rect 33290 3863 33300 3925
rect 33289 3822 33300 3863
rect 33470 3925 33481 3966
rect 33470 3863 33480 3925
rect 33470 3822 33481 3863
rect 33289 3817 33481 3822
rect 33536 3785 33606 4003
rect 33661 3966 33853 3971
rect 33661 3925 33672 3966
rect 33662 3863 33672 3925
rect 33661 3822 33672 3863
rect 33842 3925 33853 3966
rect 33842 3863 33852 3925
rect 33842 3822 33853 3863
rect 33661 3817 33853 3822
rect 33908 3785 33978 4003
rect 34033 3966 34225 3971
rect 34033 3925 34044 3966
rect 34034 3863 34044 3925
rect 34033 3822 34044 3863
rect 34214 3925 34225 3966
rect 34214 3863 34224 3925
rect 34214 3822 34225 3863
rect 34033 3817 34225 3822
rect 34280 3785 34350 4003
rect 34405 3966 34597 3971
rect 34405 3925 34416 3966
rect 34406 3863 34416 3925
rect 34405 3822 34416 3863
rect 34586 3925 34597 3966
rect 34586 3863 34596 3925
rect 34586 3822 34597 3863
rect 34405 3817 34597 3822
rect 34652 3785 34722 4003
rect 34777 3966 34969 3971
rect 34777 3925 34788 3966
rect 34778 3863 34788 3925
rect 34777 3822 34788 3863
rect 34958 3925 34969 3966
rect 34958 3863 34968 3925
rect 34958 3822 34969 3863
rect 34777 3817 34969 3822
rect 35024 3785 35094 4003
rect 35149 3966 35341 3971
rect 35149 3925 35160 3966
rect 35150 3863 35160 3925
rect 35149 3822 35160 3863
rect 35330 3925 35341 3966
rect 35330 3863 35340 3925
rect 35330 3822 35341 3863
rect 35149 3817 35341 3822
rect 35396 3785 35466 4003
rect 35521 3966 35713 3971
rect 35521 3925 35532 3966
rect 35522 3863 35532 3925
rect 35521 3822 35532 3863
rect 35702 3925 35713 3966
rect 35702 3863 35712 3925
rect 35702 3822 35713 3863
rect 35521 3817 35713 3822
rect 35768 3785 35838 4003
rect 35893 3966 36085 3971
rect 35893 3925 35904 3966
rect 35894 3863 35904 3925
rect 35893 3822 35904 3863
rect 36074 3925 36085 3966
rect 36074 3863 36084 3925
rect 36074 3822 36085 3863
rect 35893 3817 36085 3822
rect 36140 3785 36210 4003
rect 36265 3966 36457 3971
rect 36265 3925 36276 3966
rect 36266 3863 36276 3925
rect 36265 3822 36276 3863
rect 36446 3925 36457 3966
rect 36446 3863 36456 3925
rect 36446 3822 36457 3863
rect 36265 3817 36457 3822
rect 36512 3785 36582 4003
rect 36637 3966 36829 3971
rect 36637 3925 36648 3966
rect 36638 3863 36648 3925
rect 36637 3822 36648 3863
rect 36818 3925 36829 3966
rect 36818 3863 36828 3925
rect 36818 3822 36829 3863
rect 36637 3817 36829 3822
rect 36884 3785 36954 4003
rect 37009 3966 37201 3971
rect 37009 3925 37020 3966
rect 37010 3863 37020 3925
rect 37009 3822 37020 3863
rect 37190 3925 37201 3966
rect 37190 3863 37200 3925
rect 37190 3822 37201 3863
rect 37009 3817 37201 3822
rect 37256 3785 37326 4003
rect 37381 3966 37573 3971
rect 37381 3925 37392 3966
rect 37382 3863 37392 3925
rect 37381 3822 37392 3863
rect 37562 3925 37573 3966
rect 37562 3863 37572 3925
rect 37562 3822 37573 3863
rect 37381 3817 37573 3822
rect 37628 3785 37698 4003
rect 37753 3966 37945 3971
rect 37753 3925 37764 3966
rect 37754 3863 37764 3925
rect 37753 3822 37764 3863
rect 37934 3925 37945 3966
rect 37934 3863 37944 3925
rect 37934 3822 37945 3863
rect 37753 3817 37945 3822
rect 38000 3785 38070 4003
rect 38125 3966 38317 3971
rect 38125 3925 38136 3966
rect 38126 3863 38136 3925
rect 38125 3822 38136 3863
rect 38306 3925 38317 3966
rect 38306 3863 38316 3925
rect 38306 3822 38317 3863
rect 38125 3817 38317 3822
rect 38372 3785 38442 4003
rect 38497 3966 38689 3971
rect 38497 3925 38508 3966
rect 38498 3863 38508 3925
rect 38497 3822 38508 3863
rect 38678 3925 38689 3966
rect 38678 3863 38688 3925
rect 38678 3822 38689 3863
rect 38497 3817 38689 3822
rect 38744 3785 38814 4003
rect 38869 3966 39061 3971
rect 38869 3925 38880 3966
rect 38870 3863 38880 3925
rect 38869 3822 38880 3863
rect 39050 3925 39061 3966
rect 39050 3863 39060 3925
rect 39050 3822 39061 3863
rect 38869 3817 39061 3822
rect 39092 3785 39166 4003
rect 30208 3773 30303 3785
rect 30208 3597 30263 3773
rect 30297 3597 30303 3773
rect 30208 3585 30303 3597
rect 30515 3773 30675 3785
rect 30515 3597 30521 3773
rect 30555 3597 30635 3773
rect 30669 3597 30675 3773
rect 30515 3585 30675 3597
rect 30887 3773 31047 3785
rect 30887 3597 30893 3773
rect 30927 3597 31007 3773
rect 31041 3597 31047 3773
rect 30887 3585 31047 3597
rect 31259 3773 31419 3785
rect 31259 3597 31265 3773
rect 31299 3597 31379 3773
rect 31413 3597 31419 3773
rect 31259 3585 31419 3597
rect 31631 3773 31791 3785
rect 31631 3597 31637 3773
rect 31671 3597 31751 3773
rect 31785 3597 31791 3773
rect 31631 3585 31791 3597
rect 32003 3773 32163 3785
rect 32003 3597 32009 3773
rect 32043 3597 32123 3773
rect 32157 3597 32163 3773
rect 32003 3585 32163 3597
rect 32375 3773 32535 3785
rect 32375 3597 32381 3773
rect 32415 3597 32495 3773
rect 32529 3597 32535 3773
rect 32375 3585 32535 3597
rect 32747 3773 32907 3785
rect 32747 3597 32753 3773
rect 32787 3597 32867 3773
rect 32901 3597 32907 3773
rect 32747 3585 32907 3597
rect 33119 3773 33279 3785
rect 33119 3597 33125 3773
rect 33159 3597 33239 3773
rect 33273 3597 33279 3773
rect 33119 3585 33279 3597
rect 33491 3773 33651 3785
rect 33491 3597 33497 3773
rect 33531 3597 33611 3773
rect 33645 3597 33651 3773
rect 33491 3585 33651 3597
rect 33863 3773 34023 3785
rect 33863 3597 33869 3773
rect 33903 3597 33983 3773
rect 34017 3597 34023 3773
rect 33863 3585 34023 3597
rect 34235 3773 34395 3785
rect 34235 3597 34241 3773
rect 34275 3597 34355 3773
rect 34389 3597 34395 3773
rect 34235 3585 34395 3597
rect 34607 3773 34767 3785
rect 34607 3597 34613 3773
rect 34647 3597 34727 3773
rect 34761 3597 34767 3773
rect 34607 3585 34767 3597
rect 34979 3773 35139 3785
rect 34979 3597 34985 3773
rect 35019 3597 35099 3773
rect 35133 3597 35139 3773
rect 34979 3585 35139 3597
rect 35351 3773 35511 3785
rect 35351 3597 35357 3773
rect 35391 3597 35471 3773
rect 35505 3597 35511 3773
rect 35351 3585 35511 3597
rect 35723 3773 35883 3785
rect 35723 3597 35729 3773
rect 35763 3597 35843 3773
rect 35877 3597 35883 3773
rect 35723 3585 35883 3597
rect 36095 3773 36255 3785
rect 36095 3597 36101 3773
rect 36135 3597 36215 3773
rect 36249 3597 36255 3773
rect 36095 3585 36255 3597
rect 36467 3773 36627 3785
rect 36467 3597 36473 3773
rect 36507 3597 36587 3773
rect 36621 3597 36627 3773
rect 36467 3585 36627 3597
rect 36839 3773 36999 3785
rect 36839 3597 36845 3773
rect 36879 3597 36959 3773
rect 36993 3597 36999 3773
rect 36839 3585 36999 3597
rect 37211 3773 37371 3785
rect 37211 3597 37217 3773
rect 37251 3597 37331 3773
rect 37365 3597 37371 3773
rect 37211 3585 37371 3597
rect 37583 3773 37743 3785
rect 37583 3597 37589 3773
rect 37623 3597 37703 3773
rect 37737 3597 37743 3773
rect 37583 3585 37743 3597
rect 37955 3773 38115 3785
rect 37955 3597 37961 3773
rect 37995 3597 38075 3773
rect 38109 3597 38115 3773
rect 37955 3585 38115 3597
rect 38327 3773 38487 3785
rect 38327 3597 38333 3773
rect 38367 3597 38447 3773
rect 38481 3597 38487 3773
rect 38327 3585 38487 3597
rect 38699 3773 38859 3785
rect 38699 3597 38705 3773
rect 38739 3597 38819 3773
rect 38853 3597 38859 3773
rect 38699 3585 38859 3597
rect 39071 3773 39166 3785
rect 39071 3597 39077 3773
rect 39111 3597 39166 3773
rect 39071 3585 39166 3597
rect 30208 3462 30282 3585
rect 30314 3553 30324 3558
rect 30313 3548 30324 3553
rect 30312 3502 30324 3548
rect 30494 3553 30504 3558
rect 30494 3548 30505 3553
rect 30560 3548 30630 3585
rect 30932 3584 31002 3585
rect 31304 3584 31374 3585
rect 31676 3584 31746 3585
rect 32048 3584 32118 3585
rect 32420 3584 32490 3585
rect 30686 3553 30696 3558
rect 30685 3548 30696 3553
rect 30494 3502 30696 3548
rect 30866 3553 30876 3558
rect 30866 3548 30877 3553
rect 30866 3502 30878 3548
rect 30312 3490 30878 3502
rect 30938 3470 30996 3584
rect 31058 3553 31068 3558
rect 31057 3507 31068 3553
rect 31238 3553 31248 3558
rect 31430 3553 31440 3558
rect 31058 3502 31068 3507
rect 31238 3507 31249 3553
rect 31429 3507 31440 3553
rect 31610 3553 31620 3558
rect 31238 3502 31248 3507
rect 31430 3502 31440 3507
rect 31610 3507 31621 3553
rect 31610 3502 31620 3507
rect 31682 3470 31740 3584
rect 31802 3553 31812 3558
rect 31801 3507 31812 3553
rect 31982 3553 31992 3558
rect 32174 3553 32184 3558
rect 31802 3502 31812 3507
rect 31982 3507 31993 3553
rect 32173 3507 32184 3553
rect 32354 3553 32364 3558
rect 31982 3502 31992 3507
rect 32174 3502 32184 3507
rect 32354 3507 32365 3553
rect 32354 3502 32364 3507
rect 32426 3470 32484 3584
rect 32546 3553 32556 3558
rect 32545 3548 32556 3553
rect 32544 3502 32556 3548
rect 32726 3553 32736 3558
rect 32726 3548 32737 3553
rect 32792 3548 32862 3585
rect 33164 3584 33234 3585
rect 33536 3584 33606 3585
rect 33908 3584 33978 3585
rect 34280 3584 34350 3585
rect 34652 3584 34722 3585
rect 35024 3584 35094 3585
rect 35396 3584 35466 3585
rect 35768 3584 35838 3585
rect 36140 3584 36210 3585
rect 36512 3584 36582 3585
rect 36884 3584 36954 3585
rect 37256 3584 37326 3585
rect 37628 3584 37698 3585
rect 38000 3584 38070 3585
rect 38372 3584 38442 3585
rect 38744 3584 38814 3585
rect 32918 3553 32928 3558
rect 32917 3548 32928 3553
rect 32726 3502 32928 3548
rect 33098 3553 33108 3558
rect 33098 3548 33109 3553
rect 33098 3502 33110 3548
rect 32544 3490 33110 3502
rect 33170 3470 33228 3584
rect 33290 3553 33300 3558
rect 33289 3507 33300 3553
rect 33470 3553 33480 3558
rect 33662 3553 33672 3558
rect 33290 3502 33300 3507
rect 33470 3507 33481 3553
rect 33661 3507 33672 3553
rect 33842 3553 33852 3558
rect 33470 3502 33480 3507
rect 33662 3502 33672 3507
rect 33842 3507 33853 3553
rect 33842 3502 33852 3507
rect 33914 3470 33972 3584
rect 34034 3553 34044 3558
rect 34033 3507 34044 3553
rect 34214 3553 34224 3558
rect 34406 3553 34416 3558
rect 34034 3502 34044 3507
rect 34214 3507 34225 3553
rect 34405 3507 34416 3553
rect 34586 3553 34596 3558
rect 34214 3502 34224 3507
rect 34406 3502 34416 3507
rect 34586 3507 34597 3553
rect 34586 3502 34596 3507
rect 34658 3470 34716 3584
rect 34778 3553 34788 3558
rect 34777 3507 34788 3553
rect 34958 3553 34968 3558
rect 35150 3553 35160 3558
rect 34778 3502 34788 3507
rect 34958 3507 34969 3553
rect 35149 3507 35160 3553
rect 35330 3553 35340 3558
rect 34958 3502 34968 3507
rect 35150 3502 35160 3507
rect 35330 3507 35341 3553
rect 35330 3502 35340 3507
rect 35402 3470 35460 3584
rect 35522 3553 35532 3558
rect 35521 3507 35532 3553
rect 35702 3553 35712 3558
rect 35894 3553 35904 3558
rect 35522 3502 35532 3507
rect 35702 3507 35713 3553
rect 35893 3507 35904 3553
rect 36074 3553 36084 3558
rect 35702 3502 35712 3507
rect 35894 3502 35904 3507
rect 36074 3507 36085 3553
rect 36074 3502 36084 3507
rect 36146 3470 36204 3584
rect 36266 3553 36276 3558
rect 36265 3507 36276 3553
rect 36446 3553 36456 3558
rect 36638 3553 36648 3558
rect 36266 3502 36276 3507
rect 36446 3507 36457 3553
rect 36637 3507 36648 3553
rect 36818 3553 36828 3558
rect 36446 3502 36456 3507
rect 36638 3502 36648 3507
rect 36818 3507 36829 3553
rect 36818 3502 36828 3507
rect 36890 3470 36948 3584
rect 37010 3553 37020 3558
rect 37009 3507 37020 3553
rect 37190 3553 37200 3558
rect 37382 3553 37392 3558
rect 37010 3502 37020 3507
rect 37190 3507 37201 3553
rect 37381 3507 37392 3553
rect 37562 3553 37572 3558
rect 37190 3502 37200 3507
rect 37382 3502 37392 3507
rect 37562 3507 37573 3553
rect 37562 3502 37572 3507
rect 37634 3470 37692 3584
rect 37754 3553 37764 3558
rect 37753 3507 37764 3553
rect 37934 3553 37944 3558
rect 38126 3553 38136 3558
rect 37754 3502 37764 3507
rect 37934 3507 37945 3553
rect 38125 3507 38136 3553
rect 38306 3553 38316 3558
rect 37934 3502 37944 3507
rect 38126 3502 38136 3507
rect 38306 3507 38317 3553
rect 38306 3502 38316 3507
rect 38378 3470 38436 3584
rect 38498 3553 38508 3558
rect 38497 3507 38508 3553
rect 38678 3553 38688 3558
rect 38870 3553 38880 3558
rect 38498 3502 38508 3507
rect 38678 3507 38689 3553
rect 38869 3507 38880 3553
rect 39050 3553 39060 3558
rect 38678 3502 38688 3507
rect 38870 3502 38880 3507
rect 39050 3507 39061 3553
rect 39050 3502 39060 3507
rect 30920 3464 31014 3470
rect 30208 3456 30346 3462
rect 30208 3386 30264 3456
rect 30334 3386 30346 3456
rect 30920 3394 30932 3464
rect 31002 3394 31014 3464
rect 30920 3388 31014 3394
rect 31664 3464 31758 3470
rect 31664 3394 31676 3464
rect 31746 3394 31758 3464
rect 31664 3388 31758 3394
rect 32408 3464 32502 3470
rect 32408 3394 32420 3464
rect 32490 3394 32502 3464
rect 32408 3388 32502 3394
rect 33152 3464 33246 3470
rect 33152 3394 33164 3464
rect 33234 3394 33246 3464
rect 33152 3388 33246 3394
rect 33896 3464 33990 3470
rect 33896 3394 33908 3464
rect 33978 3394 33990 3464
rect 33896 3388 33990 3394
rect 34640 3464 34734 3470
rect 34640 3394 34652 3464
rect 34722 3394 34734 3464
rect 34640 3388 34734 3394
rect 35384 3464 35478 3470
rect 35384 3394 35396 3464
rect 35466 3394 35478 3464
rect 35384 3388 35478 3394
rect 36128 3464 36222 3470
rect 36128 3394 36140 3464
rect 36210 3394 36222 3464
rect 36128 3388 36222 3394
rect 36872 3464 36966 3470
rect 36872 3394 36884 3464
rect 36954 3394 36966 3464
rect 36872 3388 36966 3394
rect 37616 3464 37710 3470
rect 37616 3394 37628 3464
rect 37698 3394 37710 3464
rect 37616 3388 37710 3394
rect 38360 3464 38454 3470
rect 39092 3466 39166 3585
rect 38360 3394 38372 3464
rect 38442 3394 38454 3464
rect 38360 3388 38454 3394
rect 39022 3460 39166 3466
rect 39022 3390 39034 3460
rect 39104 3390 39166 3460
rect 30208 3380 30346 3386
rect 30208 3348 30282 3380
rect 30938 3348 30996 3388
rect 31682 3348 31740 3388
rect 32426 3348 32484 3388
rect 33170 3348 33228 3388
rect 33914 3348 33972 3388
rect 34658 3348 34716 3388
rect 35402 3348 35460 3388
rect 36146 3348 36204 3388
rect 36890 3348 36948 3388
rect 37634 3348 37692 3388
rect 38378 3348 38436 3388
rect 39022 3384 39166 3390
rect 39092 3360 39166 3384
rect 39092 3348 39180 3360
rect 30134 3148 30144 3348
rect 30344 3148 30354 3348
rect 30858 3148 30868 3348
rect 31068 3148 31078 3348
rect 31602 3148 31612 3348
rect 31812 3148 31822 3348
rect 32346 3148 32356 3348
rect 32556 3148 32566 3348
rect 33090 3148 33100 3348
rect 33300 3148 33310 3348
rect 33834 3148 33844 3348
rect 34044 3148 34054 3348
rect 34578 3148 34588 3348
rect 34788 3148 34798 3348
rect 35322 3148 35332 3348
rect 35532 3148 35542 3348
rect 36066 3148 36076 3348
rect 36276 3148 36286 3348
rect 36810 3148 36820 3348
rect 37020 3148 37030 3348
rect 37554 3148 37564 3348
rect 37764 3148 37774 3348
rect 38298 3148 38308 3348
rect 38508 3148 38518 3348
rect 39042 3148 39052 3348
rect 39252 3148 39262 3348
<< via1 >>
rect 29006 12394 29206 12594
rect 29750 12394 29950 12594
rect 30494 12394 30694 12594
rect 31238 12394 31438 12594
rect 31982 12394 32182 12594
rect 32726 12394 32926 12594
rect 33470 12394 33670 12594
rect 34214 12394 34414 12594
rect 34586 12394 34786 12594
rect 35330 12394 35530 12594
rect 36074 12394 36274 12594
rect 36818 12394 37018 12594
rect 37562 12394 37762 12594
rect 38306 12394 38506 12594
rect 39050 12394 39250 12594
rect 39794 12394 39994 12594
rect 40538 12394 40738 12594
rect 28836 12193 29006 12206
rect 28836 12159 28837 12193
rect 28837 12159 29005 12193
rect 29005 12159 29006 12193
rect 28836 12146 29006 12159
rect 29208 12193 29378 12206
rect 29208 12159 29209 12193
rect 29209 12159 29377 12193
rect 29377 12159 29378 12193
rect 29208 12146 29378 12159
rect 29580 12193 29750 12206
rect 29580 12159 29581 12193
rect 29581 12159 29749 12193
rect 29749 12159 29750 12193
rect 29580 12146 29750 12159
rect 29952 12193 30122 12206
rect 29952 12159 29953 12193
rect 29953 12159 30121 12193
rect 30121 12159 30122 12193
rect 29952 12146 30122 12159
rect 30324 12193 30494 12206
rect 30324 12159 30325 12193
rect 30325 12159 30493 12193
rect 30493 12159 30494 12193
rect 30324 12146 30494 12159
rect 30696 12193 30866 12206
rect 30696 12159 30697 12193
rect 30697 12159 30865 12193
rect 30865 12159 30866 12193
rect 30696 12146 30866 12159
rect 31068 12193 31238 12206
rect 31068 12159 31069 12193
rect 31069 12159 31237 12193
rect 31237 12159 31238 12193
rect 31068 12146 31238 12159
rect 31440 12193 31610 12206
rect 31440 12159 31441 12193
rect 31441 12159 31609 12193
rect 31609 12159 31610 12193
rect 31440 12146 31610 12159
rect 31812 12193 31982 12206
rect 31812 12159 31813 12193
rect 31813 12159 31981 12193
rect 31981 12159 31982 12193
rect 31812 12146 31982 12159
rect 32184 12193 32354 12206
rect 32184 12159 32185 12193
rect 32185 12159 32353 12193
rect 32353 12159 32354 12193
rect 32184 12146 32354 12159
rect 32556 12193 32726 12206
rect 32556 12159 32557 12193
rect 32557 12159 32725 12193
rect 32725 12159 32726 12193
rect 32556 12146 32726 12159
rect 32928 12193 33098 12206
rect 32928 12159 32929 12193
rect 32929 12159 33097 12193
rect 33097 12159 33098 12193
rect 32928 12146 33098 12159
rect 33300 12193 33470 12206
rect 33300 12159 33301 12193
rect 33301 12159 33469 12193
rect 33469 12159 33470 12193
rect 33300 12146 33470 12159
rect 33672 12193 33842 12206
rect 33672 12159 33673 12193
rect 33673 12159 33841 12193
rect 33841 12159 33842 12193
rect 33672 12146 33842 12159
rect 34044 12193 34214 12206
rect 34044 12159 34045 12193
rect 34045 12159 34213 12193
rect 34213 12159 34214 12193
rect 34044 12146 34214 12159
rect 34416 12193 34586 12206
rect 34416 12159 34417 12193
rect 34417 12159 34585 12193
rect 34585 12159 34586 12193
rect 34416 12146 34586 12159
rect 28836 11665 29006 11666
rect 28836 11631 28837 11665
rect 28837 11631 29005 11665
rect 29005 11631 29006 11665
rect 28836 11557 29006 11631
rect 28836 11523 28837 11557
rect 28837 11523 29005 11557
rect 29005 11523 29006 11557
rect 28836 11522 29006 11523
rect 29208 11665 29378 11666
rect 29208 11631 29209 11665
rect 29209 11631 29377 11665
rect 29377 11631 29378 11665
rect 29208 11557 29378 11631
rect 29208 11523 29209 11557
rect 29209 11523 29377 11557
rect 29377 11523 29378 11557
rect 29208 11522 29378 11523
rect 29580 11665 29750 11666
rect 29580 11631 29581 11665
rect 29581 11631 29749 11665
rect 29749 11631 29750 11665
rect 29580 11557 29750 11631
rect 29580 11523 29581 11557
rect 29581 11523 29749 11557
rect 29749 11523 29750 11557
rect 29580 11522 29750 11523
rect 29952 11665 30122 11666
rect 29952 11631 29953 11665
rect 29953 11631 30121 11665
rect 30121 11631 30122 11665
rect 29952 11557 30122 11631
rect 29952 11523 29953 11557
rect 29953 11523 30121 11557
rect 30121 11523 30122 11557
rect 29952 11522 30122 11523
rect 30324 11665 30494 11666
rect 30324 11631 30325 11665
rect 30325 11631 30493 11665
rect 30493 11631 30494 11665
rect 30324 11557 30494 11631
rect 30324 11523 30325 11557
rect 30325 11523 30493 11557
rect 30493 11523 30494 11557
rect 30324 11522 30494 11523
rect 30696 11665 30866 11666
rect 30696 11631 30697 11665
rect 30697 11631 30865 11665
rect 30865 11631 30866 11665
rect 30696 11557 30866 11631
rect 30696 11523 30697 11557
rect 30697 11523 30865 11557
rect 30865 11523 30866 11557
rect 30696 11522 30866 11523
rect 31068 11665 31238 11666
rect 31068 11631 31069 11665
rect 31069 11631 31237 11665
rect 31237 11631 31238 11665
rect 31068 11557 31238 11631
rect 31068 11523 31069 11557
rect 31069 11523 31237 11557
rect 31237 11523 31238 11557
rect 31068 11522 31238 11523
rect 31440 11665 31610 11666
rect 31440 11631 31441 11665
rect 31441 11631 31609 11665
rect 31609 11631 31610 11665
rect 31440 11557 31610 11631
rect 31440 11523 31441 11557
rect 31441 11523 31609 11557
rect 31609 11523 31610 11557
rect 31440 11522 31610 11523
rect 31812 11665 31982 11666
rect 31812 11631 31813 11665
rect 31813 11631 31981 11665
rect 31981 11631 31982 11665
rect 31812 11557 31982 11631
rect 31812 11523 31813 11557
rect 31813 11523 31981 11557
rect 31981 11523 31982 11557
rect 31812 11522 31982 11523
rect 32184 11665 32354 11666
rect 32184 11631 32185 11665
rect 32185 11631 32353 11665
rect 32353 11631 32354 11665
rect 32184 11557 32354 11631
rect 32184 11523 32185 11557
rect 32185 11523 32353 11557
rect 32353 11523 32354 11557
rect 32184 11522 32354 11523
rect 32556 11665 32726 11666
rect 32556 11631 32557 11665
rect 32557 11631 32725 11665
rect 32725 11631 32726 11665
rect 32556 11557 32726 11631
rect 32556 11523 32557 11557
rect 32557 11523 32725 11557
rect 32725 11523 32726 11557
rect 32556 11522 32726 11523
rect 32928 11665 33098 11666
rect 32928 11631 32929 11665
rect 32929 11631 33097 11665
rect 33097 11631 33098 11665
rect 32928 11557 33098 11631
rect 32928 11523 32929 11557
rect 32929 11523 33097 11557
rect 33097 11523 33098 11557
rect 32928 11522 33098 11523
rect 33300 11665 33470 11666
rect 33300 11631 33301 11665
rect 33301 11631 33469 11665
rect 33469 11631 33470 11665
rect 33300 11557 33470 11631
rect 33300 11523 33301 11557
rect 33301 11523 33469 11557
rect 33469 11523 33470 11557
rect 33300 11522 33470 11523
rect 33672 11665 33842 11666
rect 33672 11631 33673 11665
rect 33673 11631 33841 11665
rect 33841 11631 33842 11665
rect 33672 11557 33842 11631
rect 33672 11523 33673 11557
rect 33673 11523 33841 11557
rect 33841 11523 33842 11557
rect 33672 11522 33842 11523
rect 34044 11665 34214 11666
rect 34044 11631 34045 11665
rect 34045 11631 34213 11665
rect 34213 11631 34214 11665
rect 34044 11557 34214 11631
rect 34044 11523 34045 11557
rect 34045 11523 34213 11557
rect 34213 11523 34214 11557
rect 34044 11522 34214 11523
rect 34416 11665 34586 11666
rect 34416 11631 34417 11665
rect 34417 11631 34585 11665
rect 34585 11631 34586 11665
rect 34416 11557 34586 11631
rect 34416 11523 34417 11557
rect 34417 11523 34585 11557
rect 34585 11523 34586 11557
rect 34416 11522 34586 11523
rect 28836 11029 29006 11030
rect 28836 10995 28837 11029
rect 28837 10995 29005 11029
rect 29005 10995 29006 11029
rect 28836 10921 29006 10995
rect 28836 10887 28837 10921
rect 28837 10887 29005 10921
rect 29005 10887 29006 10921
rect 28836 10886 29006 10887
rect 29208 11029 29378 11030
rect 29208 10995 29209 11029
rect 29209 10995 29377 11029
rect 29377 10995 29378 11029
rect 29208 10921 29378 10995
rect 29208 10887 29209 10921
rect 29209 10887 29377 10921
rect 29377 10887 29378 10921
rect 29208 10886 29378 10887
rect 29580 11029 29750 11030
rect 29580 10995 29581 11029
rect 29581 10995 29749 11029
rect 29749 10995 29750 11029
rect 29580 10921 29750 10995
rect 29580 10887 29581 10921
rect 29581 10887 29749 10921
rect 29749 10887 29750 10921
rect 29580 10886 29750 10887
rect 29952 11029 30122 11030
rect 29952 10995 29953 11029
rect 29953 10995 30121 11029
rect 30121 10995 30122 11029
rect 29952 10921 30122 10995
rect 29952 10887 29953 10921
rect 29953 10887 30121 10921
rect 30121 10887 30122 10921
rect 29952 10886 30122 10887
rect 30324 11029 30494 11030
rect 30324 10995 30325 11029
rect 30325 10995 30493 11029
rect 30493 10995 30494 11029
rect 30324 10921 30494 10995
rect 30324 10887 30325 10921
rect 30325 10887 30493 10921
rect 30493 10887 30494 10921
rect 30324 10886 30494 10887
rect 30696 11029 30866 11030
rect 30696 10995 30697 11029
rect 30697 10995 30865 11029
rect 30865 10995 30866 11029
rect 30696 10921 30866 10995
rect 30696 10887 30697 10921
rect 30697 10887 30865 10921
rect 30865 10887 30866 10921
rect 30696 10886 30866 10887
rect 31068 11029 31238 11030
rect 31068 10995 31069 11029
rect 31069 10995 31237 11029
rect 31237 10995 31238 11029
rect 31068 10921 31238 10995
rect 31068 10887 31069 10921
rect 31069 10887 31237 10921
rect 31237 10887 31238 10921
rect 31068 10886 31238 10887
rect 31440 11029 31610 11030
rect 31440 10995 31441 11029
rect 31441 10995 31609 11029
rect 31609 10995 31610 11029
rect 31440 10921 31610 10995
rect 31440 10887 31441 10921
rect 31441 10887 31609 10921
rect 31609 10887 31610 10921
rect 31440 10886 31610 10887
rect 31812 11029 31982 11030
rect 31812 10995 31813 11029
rect 31813 10995 31981 11029
rect 31981 10995 31982 11029
rect 31812 10921 31982 10995
rect 31812 10887 31813 10921
rect 31813 10887 31981 10921
rect 31981 10887 31982 10921
rect 31812 10886 31982 10887
rect 32184 11029 32354 11030
rect 32184 10995 32185 11029
rect 32185 10995 32353 11029
rect 32353 10995 32354 11029
rect 32184 10921 32354 10995
rect 32184 10887 32185 10921
rect 32185 10887 32353 10921
rect 32353 10887 32354 10921
rect 32184 10886 32354 10887
rect 32556 11029 32726 11030
rect 32556 10995 32557 11029
rect 32557 10995 32725 11029
rect 32725 10995 32726 11029
rect 32556 10921 32726 10995
rect 32556 10887 32557 10921
rect 32557 10887 32725 10921
rect 32725 10887 32726 10921
rect 32556 10886 32726 10887
rect 32928 11029 33098 11030
rect 32928 10995 32929 11029
rect 32929 10995 33097 11029
rect 33097 10995 33098 11029
rect 32928 10921 33098 10995
rect 32928 10887 32929 10921
rect 32929 10887 33097 10921
rect 33097 10887 33098 10921
rect 32928 10886 33098 10887
rect 33300 11029 33470 11030
rect 33300 10995 33301 11029
rect 33301 10995 33469 11029
rect 33469 10995 33470 11029
rect 33300 10921 33470 10995
rect 33300 10887 33301 10921
rect 33301 10887 33469 10921
rect 33469 10887 33470 10921
rect 33300 10886 33470 10887
rect 33672 11029 33842 11030
rect 33672 10995 33673 11029
rect 33673 10995 33841 11029
rect 33841 10995 33842 11029
rect 33672 10921 33842 10995
rect 33672 10887 33673 10921
rect 33673 10887 33841 10921
rect 33841 10887 33842 10921
rect 33672 10886 33842 10887
rect 34044 11029 34214 11030
rect 34044 10995 34045 11029
rect 34045 10995 34213 11029
rect 34213 10995 34214 11029
rect 34044 10921 34214 10995
rect 34044 10887 34045 10921
rect 34045 10887 34213 10921
rect 34213 10887 34214 10921
rect 34044 10886 34214 10887
rect 34416 11029 34586 11030
rect 34416 10995 34417 11029
rect 34417 10995 34585 11029
rect 34585 10995 34586 11029
rect 34416 10921 34586 10995
rect 34416 10887 34417 10921
rect 34417 10887 34585 10921
rect 34585 10887 34586 10921
rect 34416 10886 34586 10887
rect 28836 10393 29006 10406
rect 28836 10359 28837 10393
rect 28837 10359 29005 10393
rect 29005 10359 29006 10393
rect 28836 10346 29006 10359
rect 29208 10393 29378 10406
rect 29208 10359 29209 10393
rect 29209 10359 29377 10393
rect 29377 10359 29378 10393
rect 29208 10346 29378 10359
rect 29580 10393 29750 10406
rect 29580 10359 29581 10393
rect 29581 10359 29749 10393
rect 29749 10359 29750 10393
rect 29580 10346 29750 10359
rect 29952 10393 30122 10406
rect 29952 10359 29953 10393
rect 29953 10359 30121 10393
rect 30121 10359 30122 10393
rect 29952 10346 30122 10359
rect 30324 10393 30494 10406
rect 30324 10359 30325 10393
rect 30325 10359 30493 10393
rect 30493 10359 30494 10393
rect 30324 10346 30494 10359
rect 30696 10393 30866 10406
rect 30696 10359 30697 10393
rect 30697 10359 30865 10393
rect 30865 10359 30866 10393
rect 30696 10346 30866 10359
rect 31068 10393 31238 10406
rect 31068 10359 31069 10393
rect 31069 10359 31237 10393
rect 31237 10359 31238 10393
rect 31068 10346 31238 10359
rect 31440 10393 31610 10406
rect 31440 10359 31441 10393
rect 31441 10359 31609 10393
rect 31609 10359 31610 10393
rect 31440 10346 31610 10359
rect 31812 10393 31982 10406
rect 31812 10359 31813 10393
rect 31813 10359 31981 10393
rect 31981 10359 31982 10393
rect 31812 10346 31982 10359
rect 32184 10393 32354 10406
rect 32184 10359 32185 10393
rect 32185 10359 32353 10393
rect 32353 10359 32354 10393
rect 32184 10346 32354 10359
rect 32556 10393 32726 10406
rect 32556 10359 32557 10393
rect 32557 10359 32725 10393
rect 32725 10359 32726 10393
rect 32556 10346 32726 10359
rect 32928 10393 33098 10406
rect 32928 10359 32929 10393
rect 32929 10359 33097 10393
rect 33097 10359 33098 10393
rect 32928 10346 33098 10359
rect 33300 10393 33470 10406
rect 33300 10359 33301 10393
rect 33301 10359 33469 10393
rect 33469 10359 33470 10393
rect 33300 10346 33470 10359
rect 33672 10393 33842 10406
rect 33672 10359 33673 10393
rect 33673 10359 33841 10393
rect 33841 10359 33842 10393
rect 33672 10346 33842 10359
rect 34788 12193 34958 12206
rect 34788 12159 34789 12193
rect 34789 12159 34957 12193
rect 34957 12159 34958 12193
rect 34788 12146 34958 12159
rect 35160 12193 35330 12206
rect 35160 12159 35161 12193
rect 35161 12159 35329 12193
rect 35329 12159 35330 12193
rect 35160 12146 35330 12159
rect 35532 12193 35702 12206
rect 35532 12159 35533 12193
rect 35533 12159 35701 12193
rect 35701 12159 35702 12193
rect 35532 12146 35702 12159
rect 35904 12193 36074 12206
rect 35904 12159 35905 12193
rect 35905 12159 36073 12193
rect 36073 12159 36074 12193
rect 35904 12146 36074 12159
rect 36276 12193 36446 12206
rect 36276 12159 36277 12193
rect 36277 12159 36445 12193
rect 36445 12159 36446 12193
rect 36276 12146 36446 12159
rect 36648 12193 36818 12206
rect 36648 12159 36649 12193
rect 36649 12159 36817 12193
rect 36817 12159 36818 12193
rect 36648 12146 36818 12159
rect 37020 12193 37190 12206
rect 37020 12159 37021 12193
rect 37021 12159 37189 12193
rect 37189 12159 37190 12193
rect 37020 12146 37190 12159
rect 37392 12193 37562 12206
rect 37392 12159 37393 12193
rect 37393 12159 37561 12193
rect 37561 12159 37562 12193
rect 37392 12146 37562 12159
rect 37764 12193 37934 12206
rect 37764 12159 37765 12193
rect 37765 12159 37933 12193
rect 37933 12159 37934 12193
rect 37764 12146 37934 12159
rect 38136 12193 38306 12206
rect 38136 12159 38137 12193
rect 38137 12159 38305 12193
rect 38305 12159 38306 12193
rect 38136 12146 38306 12159
rect 38508 12193 38678 12206
rect 38508 12159 38509 12193
rect 38509 12159 38677 12193
rect 38677 12159 38678 12193
rect 38508 12146 38678 12159
rect 38880 12193 39050 12206
rect 38880 12159 38881 12193
rect 38881 12159 39049 12193
rect 39049 12159 39050 12193
rect 38880 12146 39050 12159
rect 39252 12193 39422 12206
rect 39252 12159 39253 12193
rect 39253 12159 39421 12193
rect 39421 12159 39422 12193
rect 39252 12146 39422 12159
rect 39624 12193 39794 12206
rect 39624 12159 39625 12193
rect 39625 12159 39793 12193
rect 39793 12159 39794 12193
rect 39624 12146 39794 12159
rect 39996 12193 40166 12206
rect 39996 12159 39997 12193
rect 39997 12159 40165 12193
rect 40165 12159 40166 12193
rect 39996 12146 40166 12159
rect 40368 12193 40538 12206
rect 40368 12159 40369 12193
rect 40369 12159 40537 12193
rect 40537 12159 40538 12193
rect 40368 12146 40538 12159
rect 34788 11665 34958 11666
rect 34788 11631 34789 11665
rect 34789 11631 34957 11665
rect 34957 11631 34958 11665
rect 34788 11557 34958 11631
rect 34788 11523 34789 11557
rect 34789 11523 34957 11557
rect 34957 11523 34958 11557
rect 34788 11522 34958 11523
rect 35160 11665 35330 11666
rect 35160 11631 35161 11665
rect 35161 11631 35329 11665
rect 35329 11631 35330 11665
rect 35160 11557 35330 11631
rect 35160 11523 35161 11557
rect 35161 11523 35329 11557
rect 35329 11523 35330 11557
rect 35160 11522 35330 11523
rect 35532 11665 35702 11666
rect 35532 11631 35533 11665
rect 35533 11631 35701 11665
rect 35701 11631 35702 11665
rect 35532 11557 35702 11631
rect 35532 11523 35533 11557
rect 35533 11523 35701 11557
rect 35701 11523 35702 11557
rect 35532 11522 35702 11523
rect 35904 11665 36074 11666
rect 35904 11631 35905 11665
rect 35905 11631 36073 11665
rect 36073 11631 36074 11665
rect 35904 11557 36074 11631
rect 35904 11523 35905 11557
rect 35905 11523 36073 11557
rect 36073 11523 36074 11557
rect 35904 11522 36074 11523
rect 36276 11665 36446 11666
rect 36276 11631 36277 11665
rect 36277 11631 36445 11665
rect 36445 11631 36446 11665
rect 36276 11557 36446 11631
rect 36276 11523 36277 11557
rect 36277 11523 36445 11557
rect 36445 11523 36446 11557
rect 36276 11522 36446 11523
rect 36648 11665 36818 11666
rect 36648 11631 36649 11665
rect 36649 11631 36817 11665
rect 36817 11631 36818 11665
rect 36648 11557 36818 11631
rect 36648 11523 36649 11557
rect 36649 11523 36817 11557
rect 36817 11523 36818 11557
rect 36648 11522 36818 11523
rect 37020 11665 37190 11666
rect 37020 11631 37021 11665
rect 37021 11631 37189 11665
rect 37189 11631 37190 11665
rect 37020 11557 37190 11631
rect 37020 11523 37021 11557
rect 37021 11523 37189 11557
rect 37189 11523 37190 11557
rect 37020 11522 37190 11523
rect 37392 11665 37562 11666
rect 37392 11631 37393 11665
rect 37393 11631 37561 11665
rect 37561 11631 37562 11665
rect 37392 11557 37562 11631
rect 37392 11523 37393 11557
rect 37393 11523 37561 11557
rect 37561 11523 37562 11557
rect 37392 11522 37562 11523
rect 37764 11665 37934 11666
rect 37764 11631 37765 11665
rect 37765 11631 37933 11665
rect 37933 11631 37934 11665
rect 37764 11557 37934 11631
rect 37764 11523 37765 11557
rect 37765 11523 37933 11557
rect 37933 11523 37934 11557
rect 37764 11522 37934 11523
rect 38136 11665 38306 11666
rect 38136 11631 38137 11665
rect 38137 11631 38305 11665
rect 38305 11631 38306 11665
rect 38136 11557 38306 11631
rect 38136 11523 38137 11557
rect 38137 11523 38305 11557
rect 38305 11523 38306 11557
rect 38136 11522 38306 11523
rect 38508 11665 38678 11666
rect 38508 11631 38509 11665
rect 38509 11631 38677 11665
rect 38677 11631 38678 11665
rect 38508 11557 38678 11631
rect 38508 11523 38509 11557
rect 38509 11523 38677 11557
rect 38677 11523 38678 11557
rect 38508 11522 38678 11523
rect 38880 11665 39050 11666
rect 38880 11631 38881 11665
rect 38881 11631 39049 11665
rect 39049 11631 39050 11665
rect 38880 11557 39050 11631
rect 38880 11523 38881 11557
rect 38881 11523 39049 11557
rect 39049 11523 39050 11557
rect 38880 11522 39050 11523
rect 39252 11665 39422 11666
rect 39252 11631 39253 11665
rect 39253 11631 39421 11665
rect 39421 11631 39422 11665
rect 39252 11557 39422 11631
rect 39252 11523 39253 11557
rect 39253 11523 39421 11557
rect 39421 11523 39422 11557
rect 39252 11522 39422 11523
rect 39624 11665 39794 11666
rect 39624 11631 39625 11665
rect 39625 11631 39793 11665
rect 39793 11631 39794 11665
rect 39624 11557 39794 11631
rect 39624 11523 39625 11557
rect 39625 11523 39793 11557
rect 39793 11523 39794 11557
rect 39624 11522 39794 11523
rect 39996 11665 40166 11666
rect 39996 11631 39997 11665
rect 39997 11631 40165 11665
rect 40165 11631 40166 11665
rect 39996 11557 40166 11631
rect 39996 11523 39997 11557
rect 39997 11523 40165 11557
rect 40165 11523 40166 11557
rect 39996 11522 40166 11523
rect 40368 11665 40538 11666
rect 40368 11631 40369 11665
rect 40369 11631 40537 11665
rect 40537 11631 40538 11665
rect 40368 11557 40538 11631
rect 40368 11523 40369 11557
rect 40369 11523 40537 11557
rect 40537 11523 40538 11557
rect 40368 11522 40538 11523
rect 34788 11029 34958 11030
rect 34788 10995 34789 11029
rect 34789 10995 34957 11029
rect 34957 10995 34958 11029
rect 34788 10921 34958 10995
rect 34788 10887 34789 10921
rect 34789 10887 34957 10921
rect 34957 10887 34958 10921
rect 34788 10886 34958 10887
rect 35160 11029 35330 11030
rect 35160 10995 35161 11029
rect 35161 10995 35329 11029
rect 35329 10995 35330 11029
rect 35160 10921 35330 10995
rect 35160 10887 35161 10921
rect 35161 10887 35329 10921
rect 35329 10887 35330 10921
rect 35160 10886 35330 10887
rect 35532 11029 35702 11030
rect 35532 10995 35533 11029
rect 35533 10995 35701 11029
rect 35701 10995 35702 11029
rect 35532 10921 35702 10995
rect 35532 10887 35533 10921
rect 35533 10887 35701 10921
rect 35701 10887 35702 10921
rect 35532 10886 35702 10887
rect 35904 11029 36074 11030
rect 35904 10995 35905 11029
rect 35905 10995 36073 11029
rect 36073 10995 36074 11029
rect 35904 10921 36074 10995
rect 35904 10887 35905 10921
rect 35905 10887 36073 10921
rect 36073 10887 36074 10921
rect 35904 10886 36074 10887
rect 36276 11029 36446 11030
rect 36276 10995 36277 11029
rect 36277 10995 36445 11029
rect 36445 10995 36446 11029
rect 36276 10921 36446 10995
rect 36276 10887 36277 10921
rect 36277 10887 36445 10921
rect 36445 10887 36446 10921
rect 36276 10886 36446 10887
rect 36648 11029 36818 11030
rect 36648 10995 36649 11029
rect 36649 10995 36817 11029
rect 36817 10995 36818 11029
rect 36648 10921 36818 10995
rect 36648 10887 36649 10921
rect 36649 10887 36817 10921
rect 36817 10887 36818 10921
rect 36648 10886 36818 10887
rect 37020 11029 37190 11030
rect 37020 10995 37021 11029
rect 37021 10995 37189 11029
rect 37189 10995 37190 11029
rect 37020 10921 37190 10995
rect 37020 10887 37021 10921
rect 37021 10887 37189 10921
rect 37189 10887 37190 10921
rect 37020 10886 37190 10887
rect 37392 11029 37562 11030
rect 37392 10995 37393 11029
rect 37393 10995 37561 11029
rect 37561 10995 37562 11029
rect 37392 10921 37562 10995
rect 37392 10887 37393 10921
rect 37393 10887 37561 10921
rect 37561 10887 37562 10921
rect 37392 10886 37562 10887
rect 37764 11029 37934 11030
rect 37764 10995 37765 11029
rect 37765 10995 37933 11029
rect 37933 10995 37934 11029
rect 37764 10921 37934 10995
rect 37764 10887 37765 10921
rect 37765 10887 37933 10921
rect 37933 10887 37934 10921
rect 37764 10886 37934 10887
rect 38136 11029 38306 11030
rect 38136 10995 38137 11029
rect 38137 10995 38305 11029
rect 38305 10995 38306 11029
rect 38136 10921 38306 10995
rect 38136 10887 38137 10921
rect 38137 10887 38305 10921
rect 38305 10887 38306 10921
rect 38136 10886 38306 10887
rect 38508 11029 38678 11030
rect 38508 10995 38509 11029
rect 38509 10995 38677 11029
rect 38677 10995 38678 11029
rect 38508 10921 38678 10995
rect 38508 10887 38509 10921
rect 38509 10887 38677 10921
rect 38677 10887 38678 10921
rect 38508 10886 38678 10887
rect 38880 11029 39050 11030
rect 38880 10995 38881 11029
rect 38881 10995 39049 11029
rect 39049 10995 39050 11029
rect 38880 10921 39050 10995
rect 38880 10887 38881 10921
rect 38881 10887 39049 10921
rect 39049 10887 39050 10921
rect 38880 10886 39050 10887
rect 39252 11029 39422 11030
rect 39252 10995 39253 11029
rect 39253 10995 39421 11029
rect 39421 10995 39422 11029
rect 39252 10921 39422 10995
rect 39252 10887 39253 10921
rect 39253 10887 39421 10921
rect 39421 10887 39422 10921
rect 39252 10886 39422 10887
rect 39624 11029 39794 11030
rect 39624 10995 39625 11029
rect 39625 10995 39793 11029
rect 39793 10995 39794 11029
rect 39624 10921 39794 10995
rect 39624 10887 39625 10921
rect 39625 10887 39793 10921
rect 39793 10887 39794 10921
rect 39624 10886 39794 10887
rect 39996 11029 40166 11030
rect 39996 10995 39997 11029
rect 39997 10995 40165 11029
rect 40165 10995 40166 11029
rect 39996 10921 40166 10995
rect 39996 10887 39997 10921
rect 39997 10887 40165 10921
rect 40165 10887 40166 10921
rect 39996 10886 40166 10887
rect 40368 11029 40538 11030
rect 40368 10995 40369 11029
rect 40369 10995 40537 11029
rect 40537 10995 40538 11029
rect 40368 10921 40538 10995
rect 40368 10887 40369 10921
rect 40369 10887 40537 10921
rect 40537 10887 40538 10921
rect 40368 10886 40538 10887
rect 34044 10393 34214 10406
rect 34044 10359 34045 10393
rect 34045 10359 34213 10393
rect 34213 10359 34214 10393
rect 34044 10346 34214 10359
rect 34416 10393 34586 10406
rect 34416 10359 34417 10393
rect 34417 10359 34585 10393
rect 34585 10359 34586 10393
rect 34416 10346 34586 10359
rect 34788 10393 34958 10406
rect 34788 10359 34789 10393
rect 34789 10359 34957 10393
rect 34957 10359 34958 10393
rect 34788 10346 34958 10359
rect 35160 10393 35330 10406
rect 35160 10359 35161 10393
rect 35161 10359 35329 10393
rect 35329 10359 35330 10393
rect 35160 10346 35330 10359
rect 35532 10393 35702 10406
rect 35532 10359 35533 10393
rect 35533 10359 35701 10393
rect 35701 10359 35702 10393
rect 35532 10346 35702 10359
rect 35904 10393 36074 10406
rect 35904 10359 35905 10393
rect 35905 10359 36073 10393
rect 36073 10359 36074 10393
rect 35904 10346 36074 10359
rect 36276 10393 36446 10406
rect 36276 10359 36277 10393
rect 36277 10359 36445 10393
rect 36445 10359 36446 10393
rect 36276 10346 36446 10359
rect 36648 10393 36818 10406
rect 36648 10359 36649 10393
rect 36649 10359 36817 10393
rect 36817 10359 36818 10393
rect 36648 10346 36818 10359
rect 37020 10393 37190 10406
rect 37020 10359 37021 10393
rect 37021 10359 37189 10393
rect 37189 10359 37190 10393
rect 37020 10346 37190 10359
rect 37392 10393 37562 10406
rect 37392 10359 37393 10393
rect 37393 10359 37561 10393
rect 37561 10359 37562 10393
rect 37392 10346 37562 10359
rect 37764 10393 37934 10406
rect 37764 10359 37765 10393
rect 37765 10359 37933 10393
rect 37933 10359 37934 10393
rect 37764 10346 37934 10359
rect 38136 10393 38306 10406
rect 38136 10359 38137 10393
rect 38137 10359 38305 10393
rect 38305 10359 38306 10393
rect 38136 10346 38306 10359
rect 38508 10393 38678 10406
rect 38508 10359 38509 10393
rect 38509 10359 38677 10393
rect 38677 10359 38678 10393
rect 38508 10346 38678 10359
rect 38880 10393 39050 10406
rect 38880 10359 38881 10393
rect 38881 10359 39049 10393
rect 39049 10359 39050 10393
rect 38880 10346 39050 10359
rect 39252 10393 39422 10406
rect 39252 10359 39253 10393
rect 39253 10359 39421 10393
rect 39421 10359 39422 10393
rect 39252 10346 39422 10359
rect 39624 10393 39794 10406
rect 39624 10359 39625 10393
rect 39625 10359 39793 10393
rect 39793 10359 39794 10393
rect 39624 10346 39794 10359
rect 39996 10393 40166 10406
rect 39996 10359 39997 10393
rect 39997 10359 40165 10393
rect 40165 10359 40166 10393
rect 39996 10346 40166 10359
rect 40368 10393 40538 10406
rect 40368 10359 40369 10393
rect 40369 10359 40537 10393
rect 40537 10359 40538 10393
rect 40368 10346 40538 10359
rect 30324 9805 30494 9820
rect 30324 9771 30325 9805
rect 30325 9771 30493 9805
rect 30493 9771 30494 9805
rect 30324 9756 30494 9771
rect 30696 9805 30866 9820
rect 30696 9771 30697 9805
rect 30697 9771 30865 9805
rect 30865 9771 30866 9805
rect 30696 9756 30866 9771
rect 31068 9805 31238 9820
rect 31068 9771 31069 9805
rect 31069 9771 31237 9805
rect 31237 9771 31238 9805
rect 31068 9756 31238 9771
rect 31440 9805 31610 9820
rect 31440 9771 31441 9805
rect 31441 9771 31609 9805
rect 31609 9771 31610 9805
rect 31440 9756 31610 9771
rect 31812 9805 31982 9820
rect 31812 9771 31813 9805
rect 31813 9771 31981 9805
rect 31981 9771 31982 9805
rect 31812 9756 31982 9771
rect 32184 9805 32354 9820
rect 32184 9771 32185 9805
rect 32185 9771 32353 9805
rect 32353 9771 32354 9805
rect 32184 9756 32354 9771
rect 32556 9805 32726 9820
rect 32556 9771 32557 9805
rect 32557 9771 32725 9805
rect 32725 9771 32726 9805
rect 32556 9756 32726 9771
rect 32928 9805 33098 9820
rect 32928 9771 32929 9805
rect 32929 9771 33097 9805
rect 33097 9771 33098 9805
rect 32928 9756 33098 9771
rect 34920 9766 35202 10038
rect 35664 9766 35946 10038
rect 36408 9766 36690 10038
rect 37152 9766 37434 10038
rect 37896 9766 38178 10038
rect 38640 9766 38922 10038
rect 39384 9766 39666 10038
rect 40128 9766 40410 10038
rect 30324 8877 30494 8878
rect 30324 8843 30325 8877
rect 30325 8843 30493 8877
rect 30493 8843 30494 8877
rect 30324 8769 30494 8843
rect 30324 8735 30325 8769
rect 30325 8735 30493 8769
rect 30493 8735 30494 8769
rect 30324 8734 30494 8735
rect 30696 8877 30866 8878
rect 30696 8843 30697 8877
rect 30697 8843 30865 8877
rect 30865 8843 30866 8877
rect 30696 8769 30866 8843
rect 30696 8735 30697 8769
rect 30697 8735 30865 8769
rect 30865 8735 30866 8769
rect 30696 8734 30866 8735
rect 31068 8877 31238 8878
rect 31068 8843 31069 8877
rect 31069 8843 31237 8877
rect 31237 8843 31238 8877
rect 31068 8769 31238 8843
rect 31068 8735 31069 8769
rect 31069 8735 31237 8769
rect 31237 8735 31238 8769
rect 31068 8734 31238 8735
rect 31440 8877 31610 8878
rect 31440 8843 31441 8877
rect 31441 8843 31609 8877
rect 31609 8843 31610 8877
rect 31440 8769 31610 8843
rect 31440 8735 31441 8769
rect 31441 8735 31609 8769
rect 31609 8735 31610 8769
rect 31440 8734 31610 8735
rect 31812 8877 31982 8878
rect 31812 8843 31813 8877
rect 31813 8843 31981 8877
rect 31981 8843 31982 8877
rect 31812 8769 31982 8843
rect 31812 8735 31813 8769
rect 31813 8735 31981 8769
rect 31981 8735 31982 8769
rect 31812 8734 31982 8735
rect 32184 8877 32354 8878
rect 32184 8843 32185 8877
rect 32185 8843 32353 8877
rect 32353 8843 32354 8877
rect 32184 8769 32354 8843
rect 32184 8735 32185 8769
rect 32185 8735 32353 8769
rect 32353 8735 32354 8769
rect 32184 8734 32354 8735
rect 32556 8877 32726 8878
rect 32556 8843 32557 8877
rect 32557 8843 32725 8877
rect 32725 8843 32726 8877
rect 32556 8769 32726 8843
rect 32556 8735 32557 8769
rect 32557 8735 32725 8769
rect 32725 8735 32726 8769
rect 32556 8734 32726 8735
rect 32928 8877 33098 8878
rect 32928 8843 32929 8877
rect 32929 8843 33097 8877
rect 33097 8843 33098 8877
rect 32928 8769 33098 8843
rect 32928 8735 32929 8769
rect 32929 8735 33097 8769
rect 33097 8735 33098 8769
rect 32928 8734 33098 8735
rect 33802 8050 34084 8322
rect 30324 7841 30494 7842
rect 30324 7807 30325 7841
rect 30325 7807 30493 7841
rect 30493 7807 30494 7841
rect 30324 7733 30494 7807
rect 30324 7699 30325 7733
rect 30325 7699 30493 7733
rect 30493 7699 30494 7733
rect 30324 7698 30494 7699
rect 30696 7841 30866 7842
rect 30696 7807 30697 7841
rect 30697 7807 30865 7841
rect 30865 7807 30866 7841
rect 30696 7733 30866 7807
rect 30696 7699 30697 7733
rect 30697 7699 30865 7733
rect 30865 7699 30866 7733
rect 30696 7698 30866 7699
rect 31068 7841 31238 7842
rect 31068 7807 31069 7841
rect 31069 7807 31237 7841
rect 31237 7807 31238 7841
rect 31068 7733 31238 7807
rect 31068 7699 31069 7733
rect 31069 7699 31237 7733
rect 31237 7699 31238 7733
rect 31068 7698 31238 7699
rect 31440 7841 31610 7842
rect 31440 7807 31441 7841
rect 31441 7807 31609 7841
rect 31609 7807 31610 7841
rect 31440 7733 31610 7807
rect 31440 7699 31441 7733
rect 31441 7699 31609 7733
rect 31609 7699 31610 7733
rect 31440 7698 31610 7699
rect 31812 7841 31982 7842
rect 31812 7807 31813 7841
rect 31813 7807 31981 7841
rect 31981 7807 31982 7841
rect 31812 7733 31982 7807
rect 31812 7699 31813 7733
rect 31813 7699 31981 7733
rect 31981 7699 31982 7733
rect 31812 7698 31982 7699
rect 32184 7841 32354 7842
rect 32184 7807 32185 7841
rect 32185 7807 32353 7841
rect 32353 7807 32354 7841
rect 32184 7733 32354 7807
rect 32184 7699 32185 7733
rect 32185 7699 32353 7733
rect 32353 7699 32354 7733
rect 32184 7698 32354 7699
rect 32556 7841 32726 7842
rect 32556 7807 32557 7841
rect 32557 7807 32725 7841
rect 32725 7807 32726 7841
rect 32556 7733 32726 7807
rect 32556 7699 32557 7733
rect 32557 7699 32725 7733
rect 32725 7699 32726 7733
rect 32556 7698 32726 7699
rect 32928 7841 33098 7842
rect 32928 7807 32929 7841
rect 32929 7807 33097 7841
rect 33097 7807 33098 7841
rect 32928 7733 33098 7807
rect 32928 7699 32929 7733
rect 32929 7699 33097 7733
rect 33097 7699 33098 7733
rect 32928 7698 33098 7699
rect 34212 7082 34356 7228
rect 30324 6805 30494 6806
rect 30324 6771 30325 6805
rect 30325 6771 30493 6805
rect 30493 6771 30494 6805
rect 30324 6697 30494 6771
rect 30324 6663 30325 6697
rect 30325 6663 30493 6697
rect 30493 6663 30494 6697
rect 30324 6662 30494 6663
rect 30696 6805 30866 6806
rect 30696 6771 30697 6805
rect 30697 6771 30865 6805
rect 30865 6771 30866 6805
rect 30696 6697 30866 6771
rect 30696 6663 30697 6697
rect 30697 6663 30865 6697
rect 30865 6663 30866 6697
rect 30696 6662 30866 6663
rect 31068 6805 31238 6806
rect 31068 6771 31069 6805
rect 31069 6771 31237 6805
rect 31237 6771 31238 6805
rect 31068 6697 31238 6771
rect 31068 6663 31069 6697
rect 31069 6663 31237 6697
rect 31237 6663 31238 6697
rect 31068 6662 31238 6663
rect 31440 6805 31610 6806
rect 31440 6771 31441 6805
rect 31441 6771 31609 6805
rect 31609 6771 31610 6805
rect 31440 6697 31610 6771
rect 31440 6663 31441 6697
rect 31441 6663 31609 6697
rect 31609 6663 31610 6697
rect 31440 6662 31610 6663
rect 31812 6805 31982 6806
rect 31812 6771 31813 6805
rect 31813 6771 31981 6805
rect 31981 6771 31982 6805
rect 31812 6697 31982 6771
rect 31812 6663 31813 6697
rect 31813 6663 31981 6697
rect 31981 6663 31982 6697
rect 31812 6662 31982 6663
rect 32184 6805 32354 6806
rect 32184 6771 32185 6805
rect 32185 6771 32353 6805
rect 32353 6771 32354 6805
rect 32184 6697 32354 6771
rect 32184 6663 32185 6697
rect 32185 6663 32353 6697
rect 32353 6663 32354 6697
rect 32184 6662 32354 6663
rect 32556 6805 32726 6806
rect 32556 6771 32557 6805
rect 32557 6771 32725 6805
rect 32725 6771 32726 6805
rect 32556 6697 32726 6771
rect 32556 6663 32557 6697
rect 32557 6663 32725 6697
rect 32725 6663 32726 6697
rect 32556 6662 32726 6663
rect 32928 6805 33098 6806
rect 32928 6771 32929 6805
rect 32929 6771 33097 6805
rect 33097 6771 33098 6805
rect 32928 6697 33098 6771
rect 32928 6663 32929 6697
rect 32929 6663 33097 6697
rect 33097 6663 33098 6697
rect 32928 6662 33098 6663
rect 34212 6682 34356 6828
rect 30324 5769 30494 5780
rect 30324 5735 30325 5769
rect 30325 5735 30493 5769
rect 30493 5735 30494 5769
rect 30324 5726 30494 5735
rect 30696 5769 30866 5780
rect 30696 5735 30697 5769
rect 30697 5735 30865 5769
rect 30865 5735 30866 5769
rect 30696 5726 30866 5735
rect 31068 5769 31238 5780
rect 31068 5735 31069 5769
rect 31069 5735 31237 5769
rect 31237 5735 31238 5769
rect 31068 5726 31238 5735
rect 31440 5769 31610 5780
rect 31440 5735 31441 5769
rect 31441 5735 31609 5769
rect 31609 5735 31610 5769
rect 31440 5726 31610 5735
rect 31812 5769 31982 5780
rect 31812 5735 31813 5769
rect 31813 5735 31981 5769
rect 31981 5735 31982 5769
rect 31812 5726 31982 5735
rect 32184 5769 32354 5780
rect 32184 5735 32185 5769
rect 32185 5735 32353 5769
rect 32353 5735 32354 5769
rect 32184 5726 32354 5735
rect 32556 5769 32726 5780
rect 32556 5735 32557 5769
rect 32557 5735 32725 5769
rect 32725 5735 32726 5769
rect 32556 5726 32726 5735
rect 31304 5260 32118 5440
rect 30324 5111 30494 5122
rect 30324 5077 30325 5111
rect 30325 5077 30493 5111
rect 30493 5077 30494 5111
rect 30324 5066 30494 5077
rect 30696 5111 30866 5122
rect 30696 5077 30697 5111
rect 30697 5077 30865 5111
rect 30865 5077 30866 5111
rect 30696 5066 30866 5077
rect 31068 5111 31238 5122
rect 31068 5077 31069 5111
rect 31069 5077 31237 5111
rect 31237 5077 31238 5111
rect 31068 5066 31238 5077
rect 31440 5111 31610 5122
rect 31440 5077 31441 5111
rect 31441 5077 31609 5111
rect 31609 5077 31610 5111
rect 31440 5066 31610 5077
rect 31812 5111 31982 5122
rect 31812 5077 31813 5111
rect 31813 5077 31981 5111
rect 31981 5077 31982 5111
rect 31812 5066 31982 5077
rect 32928 5769 33098 5780
rect 32928 5735 32929 5769
rect 32929 5735 33097 5769
rect 33097 5735 33098 5769
rect 32928 5726 33098 5735
rect 33430 5584 33712 5856
rect 32184 5111 32354 5122
rect 32184 5077 32185 5111
rect 32185 5077 32353 5111
rect 32353 5077 32354 5111
rect 32184 5066 32354 5077
rect 32556 5111 32726 5122
rect 32556 5077 32557 5111
rect 32557 5077 32725 5111
rect 32725 5077 32726 5111
rect 32556 5066 32726 5077
rect 32928 5111 33098 5122
rect 32928 5077 32929 5111
rect 32929 5077 33097 5111
rect 33097 5077 33098 5111
rect 32928 5066 33098 5077
rect 33300 5111 33470 5122
rect 33300 5077 33301 5111
rect 33301 5077 33469 5111
rect 33469 5077 33470 5111
rect 33300 5066 33470 5077
rect 34212 6282 34356 6428
rect 34174 5584 34456 5856
rect 34918 5584 35200 5856
rect 35662 5584 35944 5856
rect 36406 5584 36688 5856
rect 37150 5584 37432 5856
rect 37894 5584 38176 5856
rect 38638 5584 38920 5856
rect 33810 5260 34060 5510
rect 33672 5111 33842 5122
rect 33672 5077 33673 5111
rect 33673 5077 33841 5111
rect 33841 5077 33842 5111
rect 33672 5066 33842 5077
rect 34044 5111 34214 5122
rect 34044 5077 34045 5111
rect 34045 5077 34213 5111
rect 34213 5077 34214 5111
rect 34044 5066 34214 5077
rect 34416 5111 34586 5122
rect 34416 5077 34417 5111
rect 34417 5077 34585 5111
rect 34585 5077 34586 5111
rect 34416 5066 34586 5077
rect 34788 5111 34958 5122
rect 34788 5077 34789 5111
rect 34789 5077 34957 5111
rect 34957 5077 34958 5111
rect 34788 5066 34958 5077
rect 35160 5111 35330 5122
rect 35160 5077 35161 5111
rect 35161 5077 35329 5111
rect 35329 5077 35330 5111
rect 35160 5066 35330 5077
rect 35532 5111 35702 5122
rect 35532 5077 35533 5111
rect 35533 5077 35701 5111
rect 35701 5077 35702 5111
rect 35532 5066 35702 5077
rect 35904 5111 36074 5122
rect 35904 5077 35905 5111
rect 35905 5077 36073 5111
rect 36073 5077 36074 5111
rect 35904 5066 36074 5077
rect 36276 5111 36446 5122
rect 36276 5077 36277 5111
rect 36277 5077 36445 5111
rect 36445 5077 36446 5111
rect 36276 5066 36446 5077
rect 36648 5111 36818 5122
rect 36648 5077 36649 5111
rect 36649 5077 36817 5111
rect 36817 5077 36818 5111
rect 36648 5066 36818 5077
rect 37020 5111 37190 5122
rect 37020 5077 37021 5111
rect 37021 5077 37189 5111
rect 37189 5077 37190 5111
rect 37020 5066 37190 5077
rect 37392 5111 37562 5122
rect 37392 5077 37393 5111
rect 37393 5077 37561 5111
rect 37561 5077 37562 5111
rect 37392 5066 37562 5077
rect 37764 5111 37934 5122
rect 37764 5077 37765 5111
rect 37765 5077 37933 5111
rect 37933 5077 37934 5111
rect 37764 5066 37934 5077
rect 38136 5111 38306 5122
rect 38136 5077 38137 5111
rect 38137 5077 38305 5111
rect 38305 5077 38306 5111
rect 38136 5066 38306 5077
rect 38508 5111 38678 5122
rect 38508 5077 38509 5111
rect 38509 5077 38677 5111
rect 38677 5077 38678 5111
rect 38508 5066 38678 5077
rect 38880 5111 39050 5122
rect 38880 5077 38881 5111
rect 38881 5077 39049 5111
rect 39049 5077 39050 5111
rect 38880 5066 39050 5077
rect 30324 4801 30494 4802
rect 30324 4767 30325 4801
rect 30325 4767 30493 4801
rect 30493 4767 30494 4801
rect 30324 4693 30494 4767
rect 30324 4659 30325 4693
rect 30325 4659 30493 4693
rect 30493 4659 30494 4693
rect 30324 4658 30494 4659
rect 30696 4801 30866 4802
rect 30696 4767 30697 4801
rect 30697 4767 30865 4801
rect 30865 4767 30866 4801
rect 30696 4693 30866 4767
rect 30696 4659 30697 4693
rect 30697 4659 30865 4693
rect 30865 4659 30866 4693
rect 30696 4658 30866 4659
rect 31068 4801 31238 4802
rect 31068 4767 31069 4801
rect 31069 4767 31237 4801
rect 31237 4767 31238 4801
rect 31068 4693 31238 4767
rect 31068 4659 31069 4693
rect 31069 4659 31237 4693
rect 31237 4659 31238 4693
rect 31068 4658 31238 4659
rect 31440 4801 31610 4802
rect 31440 4767 31441 4801
rect 31441 4767 31609 4801
rect 31609 4767 31610 4801
rect 31440 4693 31610 4767
rect 31440 4659 31441 4693
rect 31441 4659 31609 4693
rect 31609 4659 31610 4693
rect 31440 4658 31610 4659
rect 31812 4801 31982 4802
rect 31812 4767 31813 4801
rect 31813 4767 31981 4801
rect 31981 4767 31982 4801
rect 31812 4693 31982 4767
rect 31812 4659 31813 4693
rect 31813 4659 31981 4693
rect 31981 4659 31982 4693
rect 31812 4658 31982 4659
rect 32184 4801 32354 4802
rect 32184 4767 32185 4801
rect 32185 4767 32353 4801
rect 32353 4767 32354 4801
rect 32184 4693 32354 4767
rect 32184 4659 32185 4693
rect 32185 4659 32353 4693
rect 32353 4659 32354 4693
rect 32184 4658 32354 4659
rect 32556 4801 32726 4802
rect 32556 4767 32557 4801
rect 32557 4767 32725 4801
rect 32725 4767 32726 4801
rect 32556 4693 32726 4767
rect 32556 4659 32557 4693
rect 32557 4659 32725 4693
rect 32725 4659 32726 4693
rect 32556 4658 32726 4659
rect 32928 4801 33098 4802
rect 32928 4767 32929 4801
rect 32929 4767 33097 4801
rect 33097 4767 33098 4801
rect 32928 4693 33098 4767
rect 32928 4659 32929 4693
rect 32929 4659 33097 4693
rect 33097 4659 33098 4693
rect 32928 4658 33098 4659
rect 33300 4801 33470 4802
rect 33300 4767 33301 4801
rect 33301 4767 33469 4801
rect 33469 4767 33470 4801
rect 33300 4693 33470 4767
rect 33300 4659 33301 4693
rect 33301 4659 33469 4693
rect 33469 4659 33470 4693
rect 33300 4658 33470 4659
rect 33672 4801 33842 4802
rect 33672 4767 33673 4801
rect 33673 4767 33841 4801
rect 33841 4767 33842 4801
rect 33672 4693 33842 4767
rect 33672 4659 33673 4693
rect 33673 4659 33841 4693
rect 33841 4659 33842 4693
rect 33672 4658 33842 4659
rect 34044 4801 34214 4802
rect 34044 4767 34045 4801
rect 34045 4767 34213 4801
rect 34213 4767 34214 4801
rect 34044 4693 34214 4767
rect 34044 4659 34045 4693
rect 34045 4659 34213 4693
rect 34213 4659 34214 4693
rect 34044 4658 34214 4659
rect 34416 4801 34586 4802
rect 34416 4767 34417 4801
rect 34417 4767 34585 4801
rect 34585 4767 34586 4801
rect 34416 4693 34586 4767
rect 34416 4659 34417 4693
rect 34417 4659 34585 4693
rect 34585 4659 34586 4693
rect 34416 4658 34586 4659
rect 34788 4801 34958 4802
rect 34788 4767 34789 4801
rect 34789 4767 34957 4801
rect 34957 4767 34958 4801
rect 34788 4693 34958 4767
rect 34788 4659 34789 4693
rect 34789 4659 34957 4693
rect 34957 4659 34958 4693
rect 34788 4658 34958 4659
rect 35160 4801 35330 4802
rect 35160 4767 35161 4801
rect 35161 4767 35329 4801
rect 35329 4767 35330 4801
rect 35160 4693 35330 4767
rect 35160 4659 35161 4693
rect 35161 4659 35329 4693
rect 35329 4659 35330 4693
rect 35160 4658 35330 4659
rect 35532 4801 35702 4802
rect 35532 4767 35533 4801
rect 35533 4767 35701 4801
rect 35701 4767 35702 4801
rect 35532 4693 35702 4767
rect 35532 4659 35533 4693
rect 35533 4659 35701 4693
rect 35701 4659 35702 4693
rect 35532 4658 35702 4659
rect 35904 4801 36074 4802
rect 35904 4767 35905 4801
rect 35905 4767 36073 4801
rect 36073 4767 36074 4801
rect 35904 4693 36074 4767
rect 35904 4659 35905 4693
rect 35905 4659 36073 4693
rect 36073 4659 36074 4693
rect 35904 4658 36074 4659
rect 36276 4801 36446 4802
rect 36276 4767 36277 4801
rect 36277 4767 36445 4801
rect 36445 4767 36446 4801
rect 36276 4693 36446 4767
rect 36276 4659 36277 4693
rect 36277 4659 36445 4693
rect 36445 4659 36446 4693
rect 36276 4658 36446 4659
rect 36648 4801 36818 4802
rect 36648 4767 36649 4801
rect 36649 4767 36817 4801
rect 36817 4767 36818 4801
rect 36648 4693 36818 4767
rect 36648 4659 36649 4693
rect 36649 4659 36817 4693
rect 36817 4659 36818 4693
rect 36648 4658 36818 4659
rect 37020 4801 37190 4802
rect 37020 4767 37021 4801
rect 37021 4767 37189 4801
rect 37189 4767 37190 4801
rect 37020 4693 37190 4767
rect 37020 4659 37021 4693
rect 37021 4659 37189 4693
rect 37189 4659 37190 4693
rect 37020 4658 37190 4659
rect 37392 4801 37562 4802
rect 37392 4767 37393 4801
rect 37393 4767 37561 4801
rect 37561 4767 37562 4801
rect 37392 4693 37562 4767
rect 37392 4659 37393 4693
rect 37393 4659 37561 4693
rect 37561 4659 37562 4693
rect 37392 4658 37562 4659
rect 37764 4801 37934 4802
rect 37764 4767 37765 4801
rect 37765 4767 37933 4801
rect 37933 4767 37934 4801
rect 37764 4693 37934 4767
rect 37764 4659 37765 4693
rect 37765 4659 37933 4693
rect 37933 4659 37934 4693
rect 37764 4658 37934 4659
rect 38136 4801 38306 4802
rect 38136 4767 38137 4801
rect 38137 4767 38305 4801
rect 38305 4767 38306 4801
rect 38136 4693 38306 4767
rect 38136 4659 38137 4693
rect 38137 4659 38305 4693
rect 38305 4659 38306 4693
rect 38136 4658 38306 4659
rect 38508 4801 38678 4802
rect 38508 4767 38509 4801
rect 38509 4767 38677 4801
rect 38677 4767 38678 4801
rect 38508 4693 38678 4767
rect 38508 4659 38509 4693
rect 38509 4659 38677 4693
rect 38677 4659 38678 4693
rect 38508 4658 38678 4659
rect 38880 4801 39050 4802
rect 38880 4767 38881 4801
rect 38881 4767 39049 4801
rect 39049 4767 39050 4801
rect 38880 4693 39050 4767
rect 38880 4659 38881 4693
rect 38881 4659 39049 4693
rect 39049 4659 39050 4693
rect 38880 4658 39050 4659
rect 30324 4383 30494 4384
rect 30324 4349 30325 4383
rect 30325 4349 30493 4383
rect 30493 4349 30494 4383
rect 30324 4275 30494 4349
rect 30324 4241 30325 4275
rect 30325 4241 30493 4275
rect 30493 4241 30494 4275
rect 30324 4240 30494 4241
rect 30696 4383 30866 4384
rect 30696 4349 30697 4383
rect 30697 4349 30865 4383
rect 30865 4349 30866 4383
rect 30696 4275 30866 4349
rect 30696 4241 30697 4275
rect 30697 4241 30865 4275
rect 30865 4241 30866 4275
rect 30696 4240 30866 4241
rect 31068 4383 31238 4384
rect 31068 4349 31069 4383
rect 31069 4349 31237 4383
rect 31237 4349 31238 4383
rect 31068 4275 31238 4349
rect 31068 4241 31069 4275
rect 31069 4241 31237 4275
rect 31237 4241 31238 4275
rect 31068 4240 31238 4241
rect 31440 4383 31610 4384
rect 31440 4349 31441 4383
rect 31441 4349 31609 4383
rect 31609 4349 31610 4383
rect 31440 4275 31610 4349
rect 31440 4241 31441 4275
rect 31441 4241 31609 4275
rect 31609 4241 31610 4275
rect 31440 4240 31610 4241
rect 31812 4383 31982 4384
rect 31812 4349 31813 4383
rect 31813 4349 31981 4383
rect 31981 4349 31982 4383
rect 31812 4275 31982 4349
rect 31812 4241 31813 4275
rect 31813 4241 31981 4275
rect 31981 4241 31982 4275
rect 31812 4240 31982 4241
rect 32184 4383 32354 4384
rect 32184 4349 32185 4383
rect 32185 4349 32353 4383
rect 32353 4349 32354 4383
rect 32184 4275 32354 4349
rect 32184 4241 32185 4275
rect 32185 4241 32353 4275
rect 32353 4241 32354 4275
rect 32184 4240 32354 4241
rect 32556 4383 32726 4384
rect 32556 4349 32557 4383
rect 32557 4349 32725 4383
rect 32725 4349 32726 4383
rect 32556 4275 32726 4349
rect 32556 4241 32557 4275
rect 32557 4241 32725 4275
rect 32725 4241 32726 4275
rect 32556 4240 32726 4241
rect 32928 4383 33098 4384
rect 32928 4349 32929 4383
rect 32929 4349 33097 4383
rect 33097 4349 33098 4383
rect 32928 4275 33098 4349
rect 32928 4241 32929 4275
rect 32929 4241 33097 4275
rect 33097 4241 33098 4275
rect 32928 4240 33098 4241
rect 33300 4383 33470 4384
rect 33300 4349 33301 4383
rect 33301 4349 33469 4383
rect 33469 4349 33470 4383
rect 33300 4275 33470 4349
rect 33300 4241 33301 4275
rect 33301 4241 33469 4275
rect 33469 4241 33470 4275
rect 33300 4240 33470 4241
rect 33672 4383 33842 4384
rect 33672 4349 33673 4383
rect 33673 4349 33841 4383
rect 33841 4349 33842 4383
rect 33672 4275 33842 4349
rect 33672 4241 33673 4275
rect 33673 4241 33841 4275
rect 33841 4241 33842 4275
rect 33672 4240 33842 4241
rect 34044 4383 34214 4384
rect 34044 4349 34045 4383
rect 34045 4349 34213 4383
rect 34213 4349 34214 4383
rect 34044 4275 34214 4349
rect 34044 4241 34045 4275
rect 34045 4241 34213 4275
rect 34213 4241 34214 4275
rect 34044 4240 34214 4241
rect 34416 4383 34586 4384
rect 34416 4349 34417 4383
rect 34417 4349 34585 4383
rect 34585 4349 34586 4383
rect 34416 4275 34586 4349
rect 34416 4241 34417 4275
rect 34417 4241 34585 4275
rect 34585 4241 34586 4275
rect 34416 4240 34586 4241
rect 34788 4383 34958 4384
rect 34788 4349 34789 4383
rect 34789 4349 34957 4383
rect 34957 4349 34958 4383
rect 34788 4275 34958 4349
rect 34788 4241 34789 4275
rect 34789 4241 34957 4275
rect 34957 4241 34958 4275
rect 34788 4240 34958 4241
rect 35160 4383 35330 4384
rect 35160 4349 35161 4383
rect 35161 4349 35329 4383
rect 35329 4349 35330 4383
rect 35160 4275 35330 4349
rect 35160 4241 35161 4275
rect 35161 4241 35329 4275
rect 35329 4241 35330 4275
rect 35160 4240 35330 4241
rect 35532 4383 35702 4384
rect 35532 4349 35533 4383
rect 35533 4349 35701 4383
rect 35701 4349 35702 4383
rect 35532 4275 35702 4349
rect 35532 4241 35533 4275
rect 35533 4241 35701 4275
rect 35701 4241 35702 4275
rect 35532 4240 35702 4241
rect 35904 4383 36074 4384
rect 35904 4349 35905 4383
rect 35905 4349 36073 4383
rect 36073 4349 36074 4383
rect 35904 4275 36074 4349
rect 35904 4241 35905 4275
rect 35905 4241 36073 4275
rect 36073 4241 36074 4275
rect 35904 4240 36074 4241
rect 36276 4383 36446 4384
rect 36276 4349 36277 4383
rect 36277 4349 36445 4383
rect 36445 4349 36446 4383
rect 36276 4275 36446 4349
rect 36276 4241 36277 4275
rect 36277 4241 36445 4275
rect 36445 4241 36446 4275
rect 36276 4240 36446 4241
rect 36648 4383 36818 4384
rect 36648 4349 36649 4383
rect 36649 4349 36817 4383
rect 36817 4349 36818 4383
rect 36648 4275 36818 4349
rect 36648 4241 36649 4275
rect 36649 4241 36817 4275
rect 36817 4241 36818 4275
rect 36648 4240 36818 4241
rect 37020 4383 37190 4384
rect 37020 4349 37021 4383
rect 37021 4349 37189 4383
rect 37189 4349 37190 4383
rect 37020 4275 37190 4349
rect 37020 4241 37021 4275
rect 37021 4241 37189 4275
rect 37189 4241 37190 4275
rect 37020 4240 37190 4241
rect 37392 4383 37562 4384
rect 37392 4349 37393 4383
rect 37393 4349 37561 4383
rect 37561 4349 37562 4383
rect 37392 4275 37562 4349
rect 37392 4241 37393 4275
rect 37393 4241 37561 4275
rect 37561 4241 37562 4275
rect 37392 4240 37562 4241
rect 37764 4383 37934 4384
rect 37764 4349 37765 4383
rect 37765 4349 37933 4383
rect 37933 4349 37934 4383
rect 37764 4275 37934 4349
rect 37764 4241 37765 4275
rect 37765 4241 37933 4275
rect 37933 4241 37934 4275
rect 37764 4240 37934 4241
rect 38136 4383 38306 4384
rect 38136 4349 38137 4383
rect 38137 4349 38305 4383
rect 38305 4349 38306 4383
rect 38136 4275 38306 4349
rect 38136 4241 38137 4275
rect 38137 4241 38305 4275
rect 38305 4241 38306 4275
rect 38136 4240 38306 4241
rect 38508 4383 38678 4384
rect 38508 4349 38509 4383
rect 38509 4349 38677 4383
rect 38677 4349 38678 4383
rect 38508 4275 38678 4349
rect 38508 4241 38509 4275
rect 38509 4241 38677 4275
rect 38677 4241 38678 4275
rect 38508 4240 38678 4241
rect 38880 4383 39050 4384
rect 38880 4349 38881 4383
rect 38881 4349 39049 4383
rect 39049 4349 39050 4383
rect 38880 4275 39050 4349
rect 38880 4241 38881 4275
rect 38881 4241 39049 4275
rect 39049 4241 39050 4275
rect 38880 4240 39050 4241
rect 30324 3965 30494 3966
rect 30324 3931 30325 3965
rect 30325 3931 30493 3965
rect 30493 3931 30494 3965
rect 30324 3857 30494 3931
rect 30324 3823 30325 3857
rect 30325 3823 30493 3857
rect 30493 3823 30494 3857
rect 30324 3822 30494 3823
rect 30696 3965 30866 3966
rect 30696 3931 30697 3965
rect 30697 3931 30865 3965
rect 30865 3931 30866 3965
rect 30696 3857 30866 3931
rect 30696 3823 30697 3857
rect 30697 3823 30865 3857
rect 30865 3823 30866 3857
rect 30696 3822 30866 3823
rect 31068 3965 31238 3966
rect 31068 3931 31069 3965
rect 31069 3931 31237 3965
rect 31237 3931 31238 3965
rect 31068 3857 31238 3931
rect 31068 3823 31069 3857
rect 31069 3823 31237 3857
rect 31237 3823 31238 3857
rect 31068 3822 31238 3823
rect 31440 3965 31610 3966
rect 31440 3931 31441 3965
rect 31441 3931 31609 3965
rect 31609 3931 31610 3965
rect 31440 3857 31610 3931
rect 31440 3823 31441 3857
rect 31441 3823 31609 3857
rect 31609 3823 31610 3857
rect 31440 3822 31610 3823
rect 31812 3965 31982 3966
rect 31812 3931 31813 3965
rect 31813 3931 31981 3965
rect 31981 3931 31982 3965
rect 31812 3857 31982 3931
rect 31812 3823 31813 3857
rect 31813 3823 31981 3857
rect 31981 3823 31982 3857
rect 31812 3822 31982 3823
rect 32184 3965 32354 3966
rect 32184 3931 32185 3965
rect 32185 3931 32353 3965
rect 32353 3931 32354 3965
rect 32184 3857 32354 3931
rect 32184 3823 32185 3857
rect 32185 3823 32353 3857
rect 32353 3823 32354 3857
rect 32184 3822 32354 3823
rect 32556 3965 32726 3966
rect 32556 3931 32557 3965
rect 32557 3931 32725 3965
rect 32725 3931 32726 3965
rect 32556 3857 32726 3931
rect 32556 3823 32557 3857
rect 32557 3823 32725 3857
rect 32725 3823 32726 3857
rect 32556 3822 32726 3823
rect 32928 3965 33098 3966
rect 32928 3931 32929 3965
rect 32929 3931 33097 3965
rect 33097 3931 33098 3965
rect 32928 3857 33098 3931
rect 32928 3823 32929 3857
rect 32929 3823 33097 3857
rect 33097 3823 33098 3857
rect 32928 3822 33098 3823
rect 33300 3965 33470 3966
rect 33300 3931 33301 3965
rect 33301 3931 33469 3965
rect 33469 3931 33470 3965
rect 33300 3857 33470 3931
rect 33300 3823 33301 3857
rect 33301 3823 33469 3857
rect 33469 3823 33470 3857
rect 33300 3822 33470 3823
rect 33672 3965 33842 3966
rect 33672 3931 33673 3965
rect 33673 3931 33841 3965
rect 33841 3931 33842 3965
rect 33672 3857 33842 3931
rect 33672 3823 33673 3857
rect 33673 3823 33841 3857
rect 33841 3823 33842 3857
rect 33672 3822 33842 3823
rect 34044 3965 34214 3966
rect 34044 3931 34045 3965
rect 34045 3931 34213 3965
rect 34213 3931 34214 3965
rect 34044 3857 34214 3931
rect 34044 3823 34045 3857
rect 34045 3823 34213 3857
rect 34213 3823 34214 3857
rect 34044 3822 34214 3823
rect 34416 3965 34586 3966
rect 34416 3931 34417 3965
rect 34417 3931 34585 3965
rect 34585 3931 34586 3965
rect 34416 3857 34586 3931
rect 34416 3823 34417 3857
rect 34417 3823 34585 3857
rect 34585 3823 34586 3857
rect 34416 3822 34586 3823
rect 34788 3965 34958 3966
rect 34788 3931 34789 3965
rect 34789 3931 34957 3965
rect 34957 3931 34958 3965
rect 34788 3857 34958 3931
rect 34788 3823 34789 3857
rect 34789 3823 34957 3857
rect 34957 3823 34958 3857
rect 34788 3822 34958 3823
rect 35160 3965 35330 3966
rect 35160 3931 35161 3965
rect 35161 3931 35329 3965
rect 35329 3931 35330 3965
rect 35160 3857 35330 3931
rect 35160 3823 35161 3857
rect 35161 3823 35329 3857
rect 35329 3823 35330 3857
rect 35160 3822 35330 3823
rect 35532 3965 35702 3966
rect 35532 3931 35533 3965
rect 35533 3931 35701 3965
rect 35701 3931 35702 3965
rect 35532 3857 35702 3931
rect 35532 3823 35533 3857
rect 35533 3823 35701 3857
rect 35701 3823 35702 3857
rect 35532 3822 35702 3823
rect 35904 3965 36074 3966
rect 35904 3931 35905 3965
rect 35905 3931 36073 3965
rect 36073 3931 36074 3965
rect 35904 3857 36074 3931
rect 35904 3823 35905 3857
rect 35905 3823 36073 3857
rect 36073 3823 36074 3857
rect 35904 3822 36074 3823
rect 36276 3965 36446 3966
rect 36276 3931 36277 3965
rect 36277 3931 36445 3965
rect 36445 3931 36446 3965
rect 36276 3857 36446 3931
rect 36276 3823 36277 3857
rect 36277 3823 36445 3857
rect 36445 3823 36446 3857
rect 36276 3822 36446 3823
rect 36648 3965 36818 3966
rect 36648 3931 36649 3965
rect 36649 3931 36817 3965
rect 36817 3931 36818 3965
rect 36648 3857 36818 3931
rect 36648 3823 36649 3857
rect 36649 3823 36817 3857
rect 36817 3823 36818 3857
rect 36648 3822 36818 3823
rect 37020 3965 37190 3966
rect 37020 3931 37021 3965
rect 37021 3931 37189 3965
rect 37189 3931 37190 3965
rect 37020 3857 37190 3931
rect 37020 3823 37021 3857
rect 37021 3823 37189 3857
rect 37189 3823 37190 3857
rect 37020 3822 37190 3823
rect 37392 3965 37562 3966
rect 37392 3931 37393 3965
rect 37393 3931 37561 3965
rect 37561 3931 37562 3965
rect 37392 3857 37562 3931
rect 37392 3823 37393 3857
rect 37393 3823 37561 3857
rect 37561 3823 37562 3857
rect 37392 3822 37562 3823
rect 37764 3965 37934 3966
rect 37764 3931 37765 3965
rect 37765 3931 37933 3965
rect 37933 3931 37934 3965
rect 37764 3857 37934 3931
rect 37764 3823 37765 3857
rect 37765 3823 37933 3857
rect 37933 3823 37934 3857
rect 37764 3822 37934 3823
rect 38136 3965 38306 3966
rect 38136 3931 38137 3965
rect 38137 3931 38305 3965
rect 38305 3931 38306 3965
rect 38136 3857 38306 3931
rect 38136 3823 38137 3857
rect 38137 3823 38305 3857
rect 38305 3823 38306 3857
rect 38136 3822 38306 3823
rect 38508 3965 38678 3966
rect 38508 3931 38509 3965
rect 38509 3931 38677 3965
rect 38677 3931 38678 3965
rect 38508 3857 38678 3931
rect 38508 3823 38509 3857
rect 38509 3823 38677 3857
rect 38677 3823 38678 3857
rect 38508 3822 38678 3823
rect 38880 3965 39050 3966
rect 38880 3931 38881 3965
rect 38881 3931 39049 3965
rect 39049 3931 39050 3965
rect 38880 3857 39050 3931
rect 38880 3823 38881 3857
rect 38881 3823 39049 3857
rect 39049 3823 39050 3857
rect 38880 3822 39050 3823
rect 30324 3547 30494 3558
rect 30324 3513 30325 3547
rect 30325 3513 30493 3547
rect 30493 3513 30494 3547
rect 30324 3502 30494 3513
rect 30696 3547 30866 3558
rect 30696 3513 30697 3547
rect 30697 3513 30865 3547
rect 30865 3513 30866 3547
rect 30696 3502 30866 3513
rect 31068 3547 31238 3558
rect 31068 3513 31069 3547
rect 31069 3513 31237 3547
rect 31237 3513 31238 3547
rect 31068 3502 31238 3513
rect 31440 3547 31610 3558
rect 31440 3513 31441 3547
rect 31441 3513 31609 3547
rect 31609 3513 31610 3547
rect 31440 3502 31610 3513
rect 31812 3547 31982 3558
rect 31812 3513 31813 3547
rect 31813 3513 31981 3547
rect 31981 3513 31982 3547
rect 31812 3502 31982 3513
rect 32184 3547 32354 3558
rect 32184 3513 32185 3547
rect 32185 3513 32353 3547
rect 32353 3513 32354 3547
rect 32184 3502 32354 3513
rect 32556 3547 32726 3558
rect 32556 3513 32557 3547
rect 32557 3513 32725 3547
rect 32725 3513 32726 3547
rect 32556 3502 32726 3513
rect 32928 3547 33098 3558
rect 32928 3513 32929 3547
rect 32929 3513 33097 3547
rect 33097 3513 33098 3547
rect 32928 3502 33098 3513
rect 33300 3547 33470 3558
rect 33300 3513 33301 3547
rect 33301 3513 33469 3547
rect 33469 3513 33470 3547
rect 33300 3502 33470 3513
rect 33672 3547 33842 3558
rect 33672 3513 33673 3547
rect 33673 3513 33841 3547
rect 33841 3513 33842 3547
rect 33672 3502 33842 3513
rect 34044 3547 34214 3558
rect 34044 3513 34045 3547
rect 34045 3513 34213 3547
rect 34213 3513 34214 3547
rect 34044 3502 34214 3513
rect 34416 3547 34586 3558
rect 34416 3513 34417 3547
rect 34417 3513 34585 3547
rect 34585 3513 34586 3547
rect 34416 3502 34586 3513
rect 34788 3547 34958 3558
rect 34788 3513 34789 3547
rect 34789 3513 34957 3547
rect 34957 3513 34958 3547
rect 34788 3502 34958 3513
rect 35160 3547 35330 3558
rect 35160 3513 35161 3547
rect 35161 3513 35329 3547
rect 35329 3513 35330 3547
rect 35160 3502 35330 3513
rect 35532 3547 35702 3558
rect 35532 3513 35533 3547
rect 35533 3513 35701 3547
rect 35701 3513 35702 3547
rect 35532 3502 35702 3513
rect 35904 3547 36074 3558
rect 35904 3513 35905 3547
rect 35905 3513 36073 3547
rect 36073 3513 36074 3547
rect 35904 3502 36074 3513
rect 36276 3547 36446 3558
rect 36276 3513 36277 3547
rect 36277 3513 36445 3547
rect 36445 3513 36446 3547
rect 36276 3502 36446 3513
rect 36648 3547 36818 3558
rect 36648 3513 36649 3547
rect 36649 3513 36817 3547
rect 36817 3513 36818 3547
rect 36648 3502 36818 3513
rect 37020 3547 37190 3558
rect 37020 3513 37021 3547
rect 37021 3513 37189 3547
rect 37189 3513 37190 3547
rect 37020 3502 37190 3513
rect 37392 3547 37562 3558
rect 37392 3513 37393 3547
rect 37393 3513 37561 3547
rect 37561 3513 37562 3547
rect 37392 3502 37562 3513
rect 37764 3547 37934 3558
rect 37764 3513 37765 3547
rect 37765 3513 37933 3547
rect 37933 3513 37934 3547
rect 37764 3502 37934 3513
rect 38136 3547 38306 3558
rect 38136 3513 38137 3547
rect 38137 3513 38305 3547
rect 38305 3513 38306 3547
rect 38136 3502 38306 3513
rect 38508 3547 38678 3558
rect 38508 3513 38509 3547
rect 38509 3513 38677 3547
rect 38677 3513 38678 3547
rect 38508 3502 38678 3513
rect 38880 3547 39050 3558
rect 38880 3513 38881 3547
rect 38881 3513 39049 3547
rect 39049 3513 39050 3547
rect 38880 3502 39050 3513
rect 30144 3148 30344 3348
rect 30868 3148 31068 3348
rect 31612 3148 31812 3348
rect 32356 3148 32556 3348
rect 33100 3148 33300 3348
rect 33844 3148 34044 3348
rect 34588 3148 34788 3348
rect 35332 3148 35532 3348
rect 36076 3148 36276 3348
rect 36820 3148 37020 3348
rect 37564 3148 37764 3348
rect 38308 3148 38508 3348
rect 39052 3148 39252 3348
<< metal2 >>
rect 29006 12594 29206 12604
rect 29006 12384 29206 12394
rect 29750 12594 29950 12604
rect 29750 12384 29950 12394
rect 30494 12594 30694 12604
rect 30494 12384 30694 12394
rect 31238 12594 31438 12604
rect 31238 12384 31438 12394
rect 31982 12594 32182 12604
rect 31982 12384 32182 12394
rect 32726 12594 32926 12604
rect 32726 12384 32926 12394
rect 33470 12594 33670 12604
rect 33470 12384 33670 12394
rect 34214 12594 34414 12604
rect 34214 12384 34414 12394
rect 34586 12594 34786 12604
rect 34586 12384 34786 12394
rect 35330 12594 35530 12604
rect 35330 12384 35530 12394
rect 36074 12594 36274 12604
rect 36074 12384 36274 12394
rect 36818 12594 37018 12604
rect 36818 12384 37018 12394
rect 37562 12594 37762 12604
rect 37562 12384 37762 12394
rect 38306 12594 38506 12604
rect 38306 12384 38506 12394
rect 39050 12594 39250 12604
rect 39050 12384 39250 12394
rect 39794 12594 39994 12604
rect 39794 12384 39994 12394
rect 40538 12594 40738 12604
rect 40538 12384 40738 12394
rect 28836 12206 40548 12216
rect 29006 12146 29208 12206
rect 29378 12146 29580 12206
rect 29750 12146 29952 12206
rect 30122 12146 30324 12206
rect 30494 12146 30696 12206
rect 30866 12146 31068 12206
rect 31238 12146 31440 12206
rect 31610 12146 31812 12206
rect 31982 12146 32184 12206
rect 32354 12146 32556 12206
rect 32726 12146 32928 12206
rect 33098 12146 33300 12206
rect 33470 12146 33672 12206
rect 33842 12146 34044 12206
rect 34214 12146 34416 12206
rect 34586 12146 34788 12206
rect 34958 12146 35160 12206
rect 35330 12146 35532 12206
rect 35702 12146 35904 12206
rect 36074 12146 36276 12206
rect 36446 12146 36648 12206
rect 36818 12146 37020 12206
rect 37190 12146 37392 12206
rect 37562 12146 37764 12206
rect 37934 12146 38136 12206
rect 38306 12146 38508 12206
rect 38678 12146 38880 12206
rect 39050 12146 39252 12206
rect 39422 12146 39624 12206
rect 39794 12146 39996 12206
rect 40166 12146 40368 12206
rect 40538 12146 40548 12206
rect 28836 12136 40548 12146
rect 28836 11666 40538 11676
rect 29006 11522 29208 11666
rect 29378 11522 29580 11666
rect 29750 11522 29952 11666
rect 30122 11522 30324 11666
rect 30494 11522 30696 11666
rect 30866 11522 31068 11666
rect 31238 11522 31440 11666
rect 31610 11522 31812 11666
rect 31982 11522 32184 11666
rect 32354 11522 32556 11666
rect 32726 11522 32928 11666
rect 33098 11522 33300 11666
rect 33470 11522 33672 11666
rect 33842 11522 34044 11666
rect 34214 11522 34416 11666
rect 34586 11522 34788 11666
rect 34958 11522 35160 11666
rect 35330 11522 35532 11666
rect 35702 11522 35904 11666
rect 36074 11522 36276 11666
rect 36446 11522 36648 11666
rect 36818 11522 37020 11666
rect 37190 11522 37392 11666
rect 37562 11522 37764 11666
rect 37934 11522 38136 11666
rect 38306 11522 38508 11666
rect 38678 11522 38880 11666
rect 39050 11522 39252 11666
rect 39422 11522 39624 11666
rect 39794 11522 39996 11666
rect 40166 11522 40368 11666
rect 28836 11512 40538 11522
rect 28836 11030 40538 11040
rect 29006 10886 29208 11030
rect 29378 10886 29580 11030
rect 29750 10886 29952 11030
rect 30122 10886 30324 11030
rect 30494 10886 30696 11030
rect 30866 10886 31068 11030
rect 31238 10886 31440 11030
rect 31610 10886 31812 11030
rect 31982 10886 32184 11030
rect 32354 10886 32556 11030
rect 32726 10886 32928 11030
rect 33098 10886 33300 11030
rect 33470 10886 33672 11030
rect 33842 10886 34044 11030
rect 34214 10886 34416 11030
rect 34586 10886 34788 11030
rect 34958 10886 35160 11030
rect 35330 10886 35532 11030
rect 35702 10886 35904 11030
rect 36074 10886 36276 11030
rect 36446 10886 36648 11030
rect 36818 10886 37020 11030
rect 37190 10886 37392 11030
rect 37562 10886 37764 11030
rect 37934 10886 38136 11030
rect 38306 10886 38508 11030
rect 38678 10886 38880 11030
rect 39050 10886 39252 11030
rect 39422 10886 39624 11030
rect 39794 10886 39996 11030
rect 40166 10886 40368 11030
rect 28836 10876 40538 10886
rect 28836 10406 40538 10416
rect 29006 10346 29208 10406
rect 29378 10346 29580 10406
rect 29750 10346 29952 10406
rect 30122 10346 30324 10406
rect 30494 10346 30696 10406
rect 30866 10346 31068 10406
rect 31238 10346 31440 10406
rect 31610 10346 31812 10406
rect 31982 10346 32184 10406
rect 32354 10346 32556 10406
rect 32726 10346 32928 10406
rect 33098 10346 33300 10406
rect 33470 10346 33672 10406
rect 33842 10346 34044 10406
rect 34214 10346 34416 10406
rect 34586 10346 34788 10406
rect 34958 10346 35160 10406
rect 35330 10346 35532 10406
rect 35702 10346 35904 10406
rect 36074 10346 36276 10406
rect 36446 10346 36648 10406
rect 36818 10346 37020 10406
rect 37190 10346 37392 10406
rect 37562 10346 37764 10406
rect 37934 10346 38136 10406
rect 38306 10346 38508 10406
rect 38678 10346 38880 10406
rect 39050 10346 39252 10406
rect 39422 10346 39624 10406
rect 39794 10346 39996 10406
rect 40166 10346 40368 10406
rect 28836 10336 40538 10346
rect 34920 10038 40410 10048
rect 29844 9920 32912 10018
rect 30510 9830 30680 9920
rect 32742 9830 32912 9920
rect 30324 9820 30866 9830
rect 30494 9756 30696 9820
rect 30324 9746 30866 9756
rect 31068 9820 32354 9830
rect 31238 9756 31440 9820
rect 31610 9756 31812 9820
rect 31982 9756 32184 9820
rect 31068 9746 32354 9756
rect 32556 9820 33098 9830
rect 32726 9756 32928 9820
rect 35202 9766 35664 10038
rect 35946 9766 36408 10038
rect 36690 9766 37152 10038
rect 37434 9766 37896 10038
rect 38178 9766 38640 10038
rect 38922 9766 39384 10038
rect 39666 9766 40128 10038
rect 34920 9756 40410 9766
rect 32556 9746 33098 9756
rect 30568 8888 30622 9746
rect 31312 8888 31366 9746
rect 32056 8888 32110 9746
rect 32800 8888 32854 9746
rect 30324 8878 30866 8888
rect 30494 8734 30696 8878
rect 30324 8724 30866 8734
rect 31068 8878 32354 8888
rect 31238 8734 31440 8878
rect 31610 8734 31812 8878
rect 31982 8734 32184 8878
rect 31068 8724 32354 8734
rect 32556 8878 33098 8888
rect 32726 8734 32928 8878
rect 32556 8724 33098 8734
rect 30568 7852 30622 8724
rect 31312 7852 31366 8724
rect 32056 7852 32110 8724
rect 32800 7852 32854 8724
rect 33802 8322 34084 8332
rect 33802 8040 34084 8050
rect 30324 7842 30866 7852
rect 30494 7698 30696 7842
rect 30324 7688 30866 7698
rect 31068 7842 32354 7852
rect 31238 7698 31440 7842
rect 31610 7698 31812 7842
rect 31982 7698 32184 7842
rect 31068 7688 32354 7698
rect 32556 7842 33098 7852
rect 32726 7698 32928 7842
rect 32556 7688 33098 7698
rect 30568 6816 30622 7688
rect 31312 6816 31366 7688
rect 32056 6816 32110 7688
rect 32800 6816 32854 7688
rect 34212 7228 34356 7238
rect 34212 7072 34356 7082
rect 34212 6828 34356 6838
rect 30324 6806 30866 6816
rect 30494 6662 30696 6806
rect 30324 6652 30866 6662
rect 31068 6806 32354 6816
rect 31238 6662 31440 6806
rect 31610 6662 31812 6806
rect 31982 6662 32184 6806
rect 31068 6652 32354 6662
rect 32556 6806 33098 6816
rect 32726 6662 32928 6806
rect 34212 6672 34356 6682
rect 32556 6652 33098 6662
rect 30568 5790 30622 6652
rect 31312 5790 31366 6652
rect 32056 5790 32110 6652
rect 32800 5790 32854 6652
rect 34212 6428 34356 6438
rect 34212 6272 34356 6282
rect 33430 5856 38930 5866
rect 30324 5780 30866 5790
rect 30494 5726 30696 5780
rect 30324 5716 30866 5726
rect 31068 5780 32354 5790
rect 31238 5726 31440 5780
rect 31610 5726 31812 5780
rect 31982 5726 32184 5780
rect 31068 5716 32354 5726
rect 32556 5780 33098 5790
rect 32726 5726 32928 5780
rect 32556 5716 33098 5726
rect 31254 5616 31424 5716
rect 31998 5616 32168 5716
rect 29844 5518 32168 5616
rect 33712 5692 34174 5856
rect 33430 5574 33712 5584
rect 34456 5692 34918 5856
rect 34174 5574 34456 5584
rect 35200 5692 35662 5856
rect 34918 5574 35200 5584
rect 35944 5692 36406 5856
rect 35662 5574 35944 5584
rect 36688 5692 37150 5856
rect 36406 5574 36688 5584
rect 37432 5692 37894 5856
rect 37150 5574 37432 5584
rect 38176 5692 38638 5856
rect 37894 5574 38176 5584
rect 38920 5692 38930 5856
rect 38638 5574 38920 5584
rect 33810 5510 34060 5520
rect 31304 5440 33810 5450
rect 32118 5306 33810 5440
rect 32118 5260 33284 5306
rect 31304 5250 33284 5260
rect 33810 5250 34060 5260
rect 33158 5132 33284 5250
rect 30324 5122 33110 5132
rect 30494 5066 30696 5122
rect 30866 5066 31068 5122
rect 31238 5066 31440 5122
rect 31610 5066 31812 5122
rect 31982 5066 32184 5122
rect 32354 5066 32556 5122
rect 32726 5066 32928 5122
rect 33098 5066 33110 5122
rect 30324 5056 33110 5066
rect 33158 5122 39050 5132
rect 33158 5066 33300 5122
rect 33470 5066 33672 5122
rect 33842 5066 34044 5122
rect 34214 5066 34416 5122
rect 34586 5066 34788 5122
rect 34958 5066 35160 5122
rect 35330 5066 35532 5122
rect 35702 5066 35904 5122
rect 36074 5066 36276 5122
rect 36446 5066 36648 5122
rect 36818 5066 37020 5122
rect 37190 5066 37392 5122
rect 37562 5066 37764 5122
rect 37934 5066 38136 5122
rect 38306 5066 38508 5122
rect 38678 5066 38880 5122
rect 33158 5056 39050 5066
rect 33158 4812 33284 5056
rect 30324 4802 33110 4812
rect 30494 4658 30696 4802
rect 30866 4658 31068 4802
rect 31238 4658 31440 4802
rect 31610 4658 31812 4802
rect 31982 4658 32184 4802
rect 32354 4658 32556 4802
rect 32726 4658 32928 4802
rect 33098 4658 33110 4802
rect 30324 4648 33110 4658
rect 33158 4802 39050 4812
rect 33158 4658 33300 4802
rect 33470 4658 33672 4802
rect 33842 4658 34044 4802
rect 34214 4658 34416 4802
rect 34586 4658 34788 4802
rect 34958 4658 35160 4802
rect 35330 4658 35532 4802
rect 35702 4658 35904 4802
rect 36074 4658 36276 4802
rect 36446 4658 36648 4802
rect 36818 4658 37020 4802
rect 37190 4658 37392 4802
rect 37562 4658 37764 4802
rect 37934 4658 38136 4802
rect 38306 4658 38508 4802
rect 38678 4658 38880 4802
rect 33158 4648 39050 4658
rect 33158 4394 33284 4648
rect 30324 4384 33110 4394
rect 30494 4240 30696 4384
rect 30866 4240 31068 4384
rect 31238 4240 31440 4384
rect 31610 4240 31812 4384
rect 31982 4240 32184 4384
rect 32354 4240 32556 4384
rect 32726 4240 32928 4384
rect 33098 4240 33110 4384
rect 30324 4230 33110 4240
rect 33158 4384 39050 4394
rect 33158 4240 33300 4384
rect 33470 4240 33672 4384
rect 33842 4240 34044 4384
rect 34214 4240 34416 4384
rect 34586 4240 34788 4384
rect 34958 4240 35160 4384
rect 35330 4240 35532 4384
rect 35702 4240 35904 4384
rect 36074 4240 36276 4384
rect 36446 4240 36648 4384
rect 36818 4240 37020 4384
rect 37190 4240 37392 4384
rect 37562 4240 37764 4384
rect 37934 4240 38136 4384
rect 38306 4240 38508 4384
rect 38678 4240 38880 4384
rect 33158 4230 39050 4240
rect 33158 3976 33284 4230
rect 30324 3966 33110 3976
rect 30494 3822 30696 3966
rect 30866 3822 31068 3966
rect 31238 3822 31440 3966
rect 31610 3822 31812 3966
rect 31982 3822 32184 3966
rect 32354 3822 32556 3966
rect 32726 3822 32928 3966
rect 33098 3822 33110 3966
rect 30324 3812 33110 3822
rect 33158 3966 39050 3976
rect 33158 3822 33300 3966
rect 33470 3822 33672 3966
rect 33842 3822 34044 3966
rect 34214 3822 34416 3966
rect 34586 3822 34788 3966
rect 34958 3822 35160 3966
rect 35330 3822 35532 3966
rect 35702 3822 35904 3966
rect 36074 3822 36276 3966
rect 36446 3822 36648 3966
rect 36818 3822 37020 3966
rect 37190 3822 37392 3966
rect 37562 3822 37764 3966
rect 37934 3822 38136 3966
rect 38306 3822 38508 3966
rect 38678 3822 38880 3966
rect 33158 3812 39050 3822
rect 33158 3568 33284 3812
rect 30324 3558 33110 3568
rect 30494 3502 30696 3558
rect 30866 3502 31068 3558
rect 31238 3502 31440 3558
rect 31610 3502 31812 3558
rect 31982 3502 32184 3558
rect 32354 3502 32556 3558
rect 32726 3502 32928 3558
rect 33098 3502 33110 3558
rect 30324 3492 33110 3502
rect 33158 3558 39050 3568
rect 33158 3502 33300 3558
rect 33470 3502 33672 3558
rect 33842 3502 34044 3558
rect 34214 3502 34416 3558
rect 34586 3502 34788 3558
rect 34958 3502 35160 3558
rect 35330 3502 35532 3558
rect 35702 3502 35904 3558
rect 36074 3502 36276 3558
rect 36446 3502 36648 3558
rect 36818 3502 37020 3558
rect 37190 3502 37392 3558
rect 37562 3502 37764 3558
rect 37934 3502 38136 3558
rect 38306 3502 38508 3558
rect 38678 3502 38880 3558
rect 33158 3492 39050 3502
rect 30144 3348 30344 3358
rect 30144 3138 30344 3148
rect 30868 3348 31068 3358
rect 30868 3138 31068 3148
rect 31612 3348 31812 3358
rect 31612 3138 31812 3148
rect 32356 3348 32556 3358
rect 32356 3138 32556 3148
rect 33100 3348 33300 3358
rect 33100 3138 33300 3148
rect 33844 3348 34044 3358
rect 33844 3138 34044 3148
rect 34588 3348 34788 3358
rect 34588 3138 34788 3148
rect 35332 3348 35532 3358
rect 35332 3138 35532 3148
rect 36076 3348 36276 3358
rect 36076 3138 36276 3148
rect 36820 3348 37020 3358
rect 36820 3138 37020 3148
rect 37564 3348 37764 3358
rect 37564 3138 37764 3148
rect 38308 3348 38508 3358
rect 38308 3138 38508 3148
rect 39052 3348 39252 3358
rect 39052 3138 39252 3148
<< via2 >>
rect 29006 12394 29206 12594
rect 29750 12394 29950 12594
rect 30494 12394 30694 12594
rect 31238 12394 31438 12594
rect 31982 12394 32182 12594
rect 32726 12394 32926 12594
rect 33470 12394 33670 12594
rect 34214 12394 34414 12594
rect 34586 12394 34786 12594
rect 35330 12394 35530 12594
rect 36074 12394 36274 12594
rect 36818 12394 37018 12594
rect 37562 12394 37762 12594
rect 38306 12394 38506 12594
rect 39050 12394 39250 12594
rect 39794 12394 39994 12594
rect 40538 12394 40738 12594
rect 36408 9766 36690 10038
rect 37152 9766 37434 10038
rect 37896 9766 38178 10038
rect 38640 9766 38922 10038
rect 33802 8050 34084 8322
rect 34212 7082 34356 7228
rect 34212 6682 34356 6828
rect 34212 6282 34356 6428
rect 36406 5584 36688 5856
rect 37150 5584 37432 5856
rect 37894 5584 38176 5856
rect 38638 5584 38920 5856
rect 30144 3148 30344 3348
rect 30868 3148 31068 3348
rect 31612 3148 31812 3348
rect 32356 3148 32556 3348
rect 33100 3148 33300 3348
rect 33844 3148 34044 3348
rect 34588 3148 34788 3348
rect 35332 3148 35532 3348
rect 36076 3148 36276 3348
rect 36820 3148 37020 3348
rect 37564 3148 37764 3348
rect 38308 3148 38508 3348
rect 39052 3148 39252 3348
<< metal3 >>
rect 28996 12594 29216 12599
rect 28996 12394 29006 12594
rect 29206 12394 29216 12594
rect 28996 12389 29216 12394
rect 29740 12594 29960 12599
rect 29740 12394 29750 12594
rect 29950 12394 29960 12594
rect 29740 12389 29960 12394
rect 30484 12594 30704 12599
rect 30484 12394 30494 12594
rect 30694 12394 30704 12594
rect 30484 12389 30704 12394
rect 31228 12594 31448 12599
rect 31228 12394 31238 12594
rect 31438 12394 31448 12594
rect 31228 12389 31448 12394
rect 31972 12594 32192 12599
rect 31972 12394 31982 12594
rect 32182 12394 32192 12594
rect 31972 12389 32192 12394
rect 32716 12594 32936 12599
rect 32716 12394 32726 12594
rect 32926 12394 32936 12594
rect 32716 12389 32936 12394
rect 33460 12594 33680 12599
rect 33460 12394 33470 12594
rect 33670 12394 33680 12594
rect 33460 12389 33680 12394
rect 34204 12594 34424 12599
rect 34204 12394 34214 12594
rect 34414 12394 34424 12594
rect 34204 12389 34424 12394
rect 34576 12594 34796 12599
rect 34576 12394 34586 12594
rect 34786 12394 34796 12594
rect 34576 12389 34796 12394
rect 35320 12594 35540 12599
rect 35320 12394 35330 12594
rect 35530 12394 35540 12594
rect 35320 12389 35540 12394
rect 36064 12594 36284 12599
rect 36064 12394 36074 12594
rect 36274 12394 36284 12594
rect 36064 12389 36284 12394
rect 36808 12594 37028 12599
rect 36808 12394 36818 12594
rect 37018 12394 37028 12594
rect 36808 12389 37028 12394
rect 37552 12594 37772 12599
rect 37552 12394 37562 12594
rect 37762 12394 37772 12594
rect 37552 12389 37772 12394
rect 38296 12594 38516 12599
rect 38296 12394 38306 12594
rect 38506 12394 38516 12594
rect 38296 12389 38516 12394
rect 39040 12594 39260 12599
rect 39040 12394 39050 12594
rect 39250 12394 39260 12594
rect 39040 12389 39260 12394
rect 39784 12594 40004 12599
rect 39784 12394 39794 12594
rect 39994 12394 40004 12594
rect 39784 12389 40004 12394
rect 40528 12594 40748 12599
rect 40528 12394 40538 12594
rect 40738 12394 40748 12594
rect 40528 12389 40748 12394
rect 36398 10038 36700 10043
rect 36398 9766 36408 10038
rect 36690 9766 36700 10038
rect 36398 9704 36700 9766
rect 37142 10038 37444 10043
rect 37142 9766 37152 10038
rect 37434 9766 37444 10038
rect 37142 9704 37444 9766
rect 37886 10038 38188 10043
rect 37886 9766 37896 10038
rect 38178 9766 38188 10038
rect 37886 9704 38188 9766
rect 38630 10038 38932 10043
rect 38630 9766 38640 10038
rect 38922 9766 38932 10038
rect 38630 9704 38932 9766
rect 33792 8322 34094 8327
rect 33792 8050 33802 8322
rect 34084 8050 34094 8322
rect 33792 8045 34094 8050
rect 34520 7930 40094 9704
rect 34202 7228 34366 7233
rect 34202 7082 34212 7228
rect 34356 7082 34366 7228
rect 34202 7077 34366 7082
rect 34520 7160 40774 7930
rect 34202 6828 34366 6833
rect 34202 6682 34212 6828
rect 34356 6682 34366 6828
rect 34202 6677 34366 6682
rect 34202 6428 34366 6433
rect 34202 6282 34212 6428
rect 34356 6282 34366 6428
rect 34202 6277 34366 6282
rect 34520 5904 40094 7160
rect 36396 5856 36698 5904
rect 36396 5584 36406 5856
rect 36688 5584 36698 5856
rect 36396 5579 36698 5584
rect 37140 5856 37442 5904
rect 37140 5584 37150 5856
rect 37432 5584 37442 5856
rect 37140 5579 37442 5584
rect 37884 5856 38186 5904
rect 37884 5584 37894 5856
rect 38176 5584 38186 5856
rect 37884 5579 38186 5584
rect 38628 5856 38930 5904
rect 38628 5584 38638 5856
rect 38920 5584 38930 5856
rect 38628 5579 38930 5584
rect 30134 3348 30354 3353
rect 30134 3148 30144 3348
rect 30344 3148 30354 3348
rect 30134 3143 30354 3148
rect 30858 3348 31078 3353
rect 30858 3148 30868 3348
rect 31068 3148 31078 3348
rect 30858 3143 31078 3148
rect 31602 3348 31822 3353
rect 31602 3148 31612 3348
rect 31812 3148 31822 3348
rect 31602 3143 31822 3148
rect 32346 3348 32566 3353
rect 32346 3148 32356 3348
rect 32556 3148 32566 3348
rect 32346 3143 32566 3148
rect 33090 3348 33310 3353
rect 33090 3148 33100 3348
rect 33300 3148 33310 3348
rect 33090 3143 33310 3148
rect 33834 3348 34054 3353
rect 33834 3148 33844 3348
rect 34044 3148 34054 3348
rect 33834 3143 34054 3148
rect 34578 3348 34798 3353
rect 34578 3148 34588 3348
rect 34788 3148 34798 3348
rect 34578 3143 34798 3148
rect 35322 3348 35542 3353
rect 35322 3148 35332 3348
rect 35532 3148 35542 3348
rect 35322 3143 35542 3148
rect 36066 3348 36286 3353
rect 36066 3148 36076 3348
rect 36276 3148 36286 3348
rect 36066 3143 36286 3148
rect 36810 3348 37030 3353
rect 36810 3148 36820 3348
rect 37020 3148 37030 3348
rect 36810 3143 37030 3148
rect 37554 3348 37774 3353
rect 37554 3148 37564 3348
rect 37764 3148 37774 3348
rect 37554 3143 37774 3148
rect 38298 3348 38518 3353
rect 38298 3148 38308 3348
rect 38508 3148 38518 3348
rect 38298 3143 38518 3148
rect 39042 3348 39262 3353
rect 39042 3148 39052 3348
rect 39252 3148 39262 3348
rect 39042 3143 39262 3148
<< via3 >>
rect 29006 12394 29206 12594
rect 29750 12394 29950 12594
rect 30494 12394 30694 12594
rect 31238 12394 31438 12594
rect 31982 12394 32182 12594
rect 32726 12394 32926 12594
rect 33470 12394 33670 12594
rect 34214 12394 34414 12594
rect 34586 12394 34786 12594
rect 35330 12394 35530 12594
rect 36074 12394 36274 12594
rect 36818 12394 37018 12594
rect 37562 12394 37762 12594
rect 38306 12394 38506 12594
rect 39050 12394 39250 12594
rect 39794 12394 39994 12594
rect 40538 12394 40738 12594
rect 33802 8050 34084 8322
rect 34212 7082 34356 7228
rect 34212 6682 34356 6828
rect 34212 6282 34356 6428
rect 30144 3148 30344 3348
rect 30868 3148 31068 3348
rect 31612 3148 31812 3348
rect 32356 3148 32556 3348
rect 33100 3148 33300 3348
rect 33844 3148 34044 3348
rect 34588 3148 34788 3348
rect 35332 3148 35532 3348
rect 36076 3148 36276 3348
rect 36820 3148 37020 3348
rect 37564 3148 37764 3348
rect 38308 3148 38508 3348
rect 39052 3148 39252 3348
<< mimcap >>
rect 34620 9564 40020 9604
rect 34620 6044 34660 9564
rect 39980 6044 40020 9564
rect 34620 6004 40020 6044
<< mimcapcontact >>
rect 34660 6044 39980 9564
<< metal4 >>
rect 28400 12594 40924 13372
rect 28400 12394 29006 12594
rect 29206 12394 29750 12594
rect 29950 12394 30494 12594
rect 30694 12394 31238 12594
rect 31438 12394 31982 12594
rect 32182 12394 32726 12594
rect 32926 12394 33470 12594
rect 33670 12394 34214 12594
rect 34414 12394 34586 12594
rect 34786 12394 35330 12594
rect 35530 12394 36074 12594
rect 36274 12394 36818 12594
rect 37018 12394 37562 12594
rect 37762 12394 38306 12594
rect 38506 12394 39050 12594
rect 39250 12394 39794 12594
rect 39994 12394 40538 12594
rect 40738 12394 40924 12594
rect 28400 12368 40924 12394
rect 34659 9564 39981 9565
rect 33801 8322 34085 8323
rect 33801 8050 33802 8322
rect 34084 8294 34085 8322
rect 34659 8294 34660 9564
rect 34084 8076 34660 8294
rect 34084 8050 34085 8076
rect 33801 8049 34085 8050
rect 34186 7228 34386 7254
rect 34186 7082 34212 7228
rect 34356 7082 34386 7228
rect 34186 6828 34386 7082
rect 34186 6682 34212 6828
rect 34356 6682 34386 6828
rect 34186 6428 34386 6682
rect 34186 6282 34212 6428
rect 34356 6282 34386 6428
rect 34186 3372 34386 6282
rect 34659 6044 34660 8076
rect 39980 6044 39981 9564
rect 34659 6043 39981 6044
rect 28400 3348 40924 3372
rect 28400 3148 30144 3348
rect 30344 3148 30868 3348
rect 31068 3148 31612 3348
rect 31812 3148 32356 3348
rect 32556 3148 33100 3348
rect 33300 3148 33844 3348
rect 34044 3148 34588 3348
rect 34788 3148 35332 3348
rect 35532 3148 36076 3348
rect 36276 3148 36820 3348
rect 37020 3148 37564 3348
rect 37764 3148 38308 3348
rect 38508 3148 39052 3348
rect 39252 3148 40924 3348
rect 28400 2368 40924 3148
<< labels >>
flabel metal4 29596 13046 29596 13046 0 FreeSans 8000 0 0 0 vdd
port 0 nsew
flabel metal4 29162 2532 29162 2532 0 FreeSans 8000 0 0 0 vss
port 4 nsew
flabel metal2 29874 9950 29874 9950 0 FreeSans 8000 0 0 0 vn
port 2 nsew
flabel metal2 29910 5550 29910 5550 0 FreeSans 8000 0 0 0 vp
port 1 nsew
flabel metal1 28786 10950 28786 10950 0 FreeSans 8000 0 0 0 vbias
port 3 nsew
flabel metal3 40604 7618 40604 7618 0 FreeSans 8000 0 0 0 vout
port 5 nsew
<< end >>
