magic
tech sky130A
magscale 1 2
timestamp 1630301600
<< nwell >>
rect -4199 244029 27521 254720
<< pwell >>
rect -4199 264246 27520 264248
rect -4199 262194 27521 264246
rect -4199 262128 -4017 262194
rect 27192 262128 27521 262194
rect -4199 262006 27521 262128
<< nmos >>
rect -3999 263238 -3969 264038
rect -3789 263238 -3759 264038
rect -3579 263238 -3549 264038
rect -3369 263238 -3339 264038
rect -3159 263238 -3129 264038
rect -2949 263238 -2919 264038
rect -2739 263238 -2709 264038
rect -2529 263238 -2499 264038
rect -2319 263238 -2289 264038
rect -2109 263238 -2079 264038
rect -1899 263238 -1869 264038
rect -1689 263238 -1659 264038
rect -1479 263238 -1449 264038
rect -1269 263238 -1239 264038
rect -1059 263238 -1029 264038
rect -849 263238 -819 264038
rect -639 263238 -609 264038
rect -429 263238 -399 264038
rect -219 263238 -189 264038
rect -9 263238 21 264038
rect 201 263238 231 264038
rect 411 263238 441 264038
rect 621 263238 651 264038
rect 831 263238 861 264038
rect 1041 263238 1071 264038
rect 1251 263238 1281 264038
rect 1461 263238 1491 264038
rect 1671 263238 1701 264038
rect 1881 263238 1911 264038
rect 2091 263238 2121 264038
rect 2301 263238 2331 264038
rect 2511 263238 2541 264038
rect 2721 263238 2751 264038
rect 2931 263238 2961 264038
rect 3141 263238 3171 264038
rect 3351 263238 3381 264038
rect 3561 263238 3591 264038
rect 3771 263238 3801 264038
rect 3981 263238 4011 264038
rect 4191 263238 4221 264038
rect 4401 263238 4431 264038
rect 4611 263238 4641 264038
rect 4821 263238 4851 264038
rect 5031 263238 5061 264038
rect 5241 263238 5271 264038
rect 5451 263238 5481 264038
rect 5661 263238 5691 264038
rect 5871 263238 5901 264038
rect 6081 263238 6111 264038
rect 6291 263238 6321 264038
rect 6501 263238 6531 264038
rect 6711 263238 6741 264038
rect 6921 263238 6951 264038
rect 7131 263238 7161 264038
rect 7341 263238 7371 264038
rect 7551 263238 7581 264038
rect 7761 263238 7791 264038
rect 7971 263238 8001 264038
rect 8181 263238 8211 264038
rect 8391 263238 8421 264038
rect 8601 263238 8631 264038
rect 8811 263238 8841 264038
rect 9021 263238 9051 264038
rect 9231 263238 9261 264038
rect 9441 263238 9471 264038
rect 9651 263238 9681 264038
rect 9861 263238 9891 264038
rect 10071 263238 10101 264038
rect 10281 263238 10311 264038
rect 10491 263238 10521 264038
rect 10701 263238 10731 264038
rect 10911 263238 10941 264038
rect 11121 263238 11151 264038
rect 11331 263238 11361 264038
rect 11541 263238 11571 264038
rect 11751 263238 11781 264038
rect 11961 263238 11991 264038
rect 12171 263238 12201 264038
rect 12381 263238 12411 264038
rect 12591 263238 12621 264038
rect 12801 263238 12831 264038
rect 13011 263238 13041 264038
rect 13221 263238 13251 264038
rect 13431 263238 13461 264038
rect 13641 263238 13671 264038
rect 13851 263238 13881 264038
rect 14061 263238 14091 264038
rect 14271 263238 14301 264038
rect 14481 263238 14511 264038
rect 14691 263238 14721 264038
rect 14901 263238 14931 264038
rect 15111 263238 15141 264038
rect 15321 263238 15351 264038
rect 15531 263238 15561 264038
rect 15741 263238 15771 264038
rect 15951 263238 15981 264038
rect 16161 263238 16191 264038
rect 16371 263238 16401 264038
rect 16581 263238 16611 264038
rect 16791 263238 16821 264038
rect 17001 263238 17031 264038
rect 17211 263238 17241 264038
rect 17421 263238 17451 264038
rect 17631 263238 17661 264038
rect 17841 263238 17871 264038
rect 18051 263238 18081 264038
rect 18261 263238 18291 264038
rect 18471 263238 18501 264038
rect 18681 263238 18711 264038
rect 18891 263238 18921 264038
rect 19101 263238 19131 264038
rect 19311 263238 19341 264038
rect 19521 263238 19551 264038
rect 19731 263238 19761 264038
rect 19941 263238 19971 264038
rect 20151 263238 20181 264038
rect 20361 263238 20391 264038
rect 20571 263238 20601 264038
rect 20781 263238 20811 264038
rect 20991 263238 21021 264038
rect 21201 263238 21231 264038
rect 21411 263238 21441 264038
rect 21621 263238 21651 264038
rect 21831 263238 21861 264038
rect 22041 263238 22071 264038
rect 22251 263238 22281 264038
rect 22461 263238 22491 264038
rect 22671 263238 22701 264038
rect 22881 263238 22911 264038
rect 23091 263238 23121 264038
rect 23301 263238 23331 264038
rect 23511 263238 23541 264038
rect 23721 263238 23751 264038
rect 23931 263238 23961 264038
rect 24141 263238 24171 264038
rect 24351 263238 24381 264038
rect 24561 263238 24591 264038
rect 24771 263238 24801 264038
rect 24981 263238 25011 264038
rect 25191 263238 25221 264038
rect 25401 263238 25431 264038
rect 25611 263238 25641 264038
rect 25821 263238 25851 264038
rect 26031 263238 26061 264038
rect 26241 263238 26271 264038
rect 26451 263238 26481 264038
rect 26661 263238 26691 264038
rect 26871 263238 26901 264038
rect 27081 263238 27111 264038
rect 27291 263238 27321 264038
rect -3999 262216 -3969 263016
rect -3789 262216 -3759 263016
rect -3579 262216 -3549 263016
rect -3369 262216 -3339 263016
rect -3159 262216 -3129 263016
rect -2949 262216 -2919 263016
rect -2739 262216 -2709 263016
rect -2529 262216 -2499 263016
rect -2319 262216 -2289 263016
rect -2109 262216 -2079 263016
rect -1899 262216 -1869 263016
rect -1689 262216 -1659 263016
rect -1479 262216 -1449 263016
rect -1269 262216 -1239 263016
rect -1059 262216 -1029 263016
rect -849 262216 -819 263016
rect -639 262216 -609 263016
rect -429 262216 -399 263016
rect -219 262216 -189 263016
rect -9 262216 21 263016
rect 201 262216 231 263016
rect 411 262216 441 263016
rect 621 262216 651 263016
rect 831 262216 861 263016
rect 1041 262216 1071 263016
rect 1251 262216 1281 263016
rect 1461 262216 1491 263016
rect 1671 262216 1701 263016
rect 1881 262216 1911 263016
rect 2091 262216 2121 263016
rect 2301 262216 2331 263016
rect 2511 262216 2541 263016
rect 2721 262216 2751 263016
rect 2931 262216 2961 263016
rect 3141 262216 3171 263016
rect 3351 262216 3381 263016
rect 3561 262216 3591 263016
rect 3771 262216 3801 263016
rect 3981 262216 4011 263016
rect 4191 262216 4221 263016
rect 4401 262216 4431 263016
rect 4611 262216 4641 263016
rect 4821 262216 4851 263016
rect 5031 262216 5061 263016
rect 5241 262216 5271 263016
rect 5451 262216 5481 263016
rect 5661 262216 5691 263016
rect 5871 262216 5901 263016
rect 6081 262216 6111 263016
rect 6291 262216 6321 263016
rect 6501 262216 6531 263016
rect 6711 262216 6741 263016
rect 6921 262216 6951 263016
rect 7131 262216 7161 263016
rect 7341 262216 7371 263016
rect 7551 262216 7581 263016
rect 7761 262216 7791 263016
rect 7971 262216 8001 263016
rect 8181 262216 8211 263016
rect 8391 262216 8421 263016
rect 8601 262216 8631 263016
rect 8811 262216 8841 263016
rect 9021 262216 9051 263016
rect 9231 262216 9261 263016
rect 9441 262216 9471 263016
rect 9651 262216 9681 263016
rect 9861 262216 9891 263016
rect 10071 262216 10101 263016
rect 10281 262216 10311 263016
rect 10491 262216 10521 263016
rect 10701 262216 10731 263016
rect 10911 262216 10941 263016
rect 11121 262216 11151 263016
rect 11331 262216 11361 263016
rect 11541 262216 11571 263016
rect 11751 262216 11781 263016
rect 11961 262216 11991 263016
rect 12171 262216 12201 263016
rect 12381 262216 12411 263016
rect 12591 262216 12621 263016
rect 12801 262216 12831 263016
rect 13011 262216 13041 263016
rect 13221 262216 13251 263016
rect 13431 262216 13461 263016
rect 13641 262216 13671 263016
rect 13851 262216 13881 263016
rect 14061 262216 14091 263016
rect 14271 262216 14301 263016
rect 14481 262216 14511 263016
rect 14691 262216 14721 263016
rect 14901 262216 14931 263016
rect 15111 262216 15141 263016
rect 15321 262216 15351 263016
rect 15531 262216 15561 263016
rect 15741 262216 15771 263016
rect 15951 262216 15981 263016
rect 16161 262216 16191 263016
rect 16371 262216 16401 263016
rect 16581 262216 16611 263016
rect 16791 262216 16821 263016
rect 17001 262216 17031 263016
rect 17211 262216 17241 263016
rect 17421 262216 17451 263016
rect 17631 262216 17661 263016
rect 17841 262216 17871 263016
rect 18051 262216 18081 263016
rect 18261 262216 18291 263016
rect 18471 262216 18501 263016
rect 18681 262216 18711 263016
rect 18891 262216 18921 263016
rect 19101 262216 19131 263016
rect 19311 262216 19341 263016
rect 19521 262216 19551 263016
rect 19731 262216 19761 263016
rect 19941 262216 19971 263016
rect 20151 262216 20181 263016
rect 20361 262216 20391 263016
rect 20571 262216 20601 263016
rect 20781 262216 20811 263016
rect 20991 262216 21021 263016
rect 21201 262216 21231 263016
rect 21411 262216 21441 263016
rect 21621 262216 21651 263016
rect 21831 262216 21861 263016
rect 22041 262216 22071 263016
rect 22251 262216 22281 263016
rect 22461 262216 22491 263016
rect 22671 262216 22701 263016
rect 22881 262216 22911 263016
rect 23091 262216 23121 263016
rect 23301 262216 23331 263016
rect 23511 262216 23541 263016
rect 23721 262216 23751 263016
rect 23931 262216 23961 263016
rect 24141 262216 24171 263016
rect 24351 262216 24381 263016
rect 24561 262216 24591 263016
rect 24771 262216 24801 263016
rect 24981 262216 25011 263016
rect 25191 262216 25221 263016
rect 25401 262216 25431 263016
rect 25611 262216 25641 263016
rect 25821 262216 25851 263016
rect 26031 262216 26061 263016
rect 26241 262216 26271 263016
rect 26451 262216 26481 263016
rect 26661 262216 26691 263016
rect 26871 262216 26901 263016
rect 27081 262216 27111 263016
rect 27291 262216 27321 263016
<< pmos >>
rect -3999 253701 -3969 254501
rect -3789 253701 -3759 254501
rect -3579 253701 -3549 254501
rect -3369 253701 -3339 254501
rect -3159 253701 -3129 254501
rect -2949 253701 -2919 254501
rect -2739 253701 -2709 254501
rect -2529 253701 -2499 254501
rect -2319 253701 -2289 254501
rect -2109 253701 -2079 254501
rect -1899 253701 -1869 254501
rect -1689 253701 -1659 254501
rect -1479 253701 -1449 254501
rect -1269 253701 -1239 254501
rect -1059 253701 -1029 254501
rect -849 253701 -819 254501
rect -639 253701 -609 254501
rect -429 253701 -399 254501
rect -219 253701 -189 254501
rect -9 253701 21 254501
rect 201 253701 231 254501
rect 411 253701 441 254501
rect 621 253701 651 254501
rect 831 253701 861 254501
rect 1041 253701 1071 254501
rect 1251 253701 1281 254501
rect 1461 253701 1491 254501
rect 1671 253701 1701 254501
rect 1881 253701 1911 254501
rect 2091 253701 2121 254501
rect 2301 253701 2331 254501
rect 2511 253701 2541 254501
rect 2721 253701 2751 254501
rect 2931 253701 2961 254501
rect 3141 253701 3171 254501
rect 3351 253701 3381 254501
rect 3561 253701 3591 254501
rect 3771 253701 3801 254501
rect 3981 253701 4011 254501
rect 4191 253701 4221 254501
rect 4401 253701 4431 254501
rect 4611 253701 4641 254501
rect 4821 253701 4851 254501
rect 5031 253701 5061 254501
rect 5241 253701 5271 254501
rect 5451 253701 5481 254501
rect 5661 253701 5691 254501
rect 5871 253701 5901 254501
rect 6081 253701 6111 254501
rect 6291 253701 6321 254501
rect 6501 253701 6531 254501
rect 6711 253701 6741 254501
rect 6921 253701 6951 254501
rect 7131 253701 7161 254501
rect 7341 253701 7371 254501
rect 7551 253701 7581 254501
rect 7761 253701 7791 254501
rect 7971 253701 8001 254501
rect 8181 253701 8211 254501
rect 8391 253701 8421 254501
rect 8601 253701 8631 254501
rect 8811 253701 8841 254501
rect 9021 253701 9051 254501
rect 9231 253701 9261 254501
rect 9441 253701 9471 254501
rect 9651 253701 9681 254501
rect 9861 253701 9891 254501
rect 10071 253701 10101 254501
rect 10281 253701 10311 254501
rect 10491 253701 10521 254501
rect 10701 253701 10731 254501
rect 10911 253701 10941 254501
rect 11121 253701 11151 254501
rect 11331 253701 11361 254501
rect 11541 253701 11571 254501
rect 11751 253701 11781 254501
rect 11961 253701 11991 254501
rect 12171 253701 12201 254501
rect 12381 253701 12411 254501
rect 12591 253701 12621 254501
rect 12801 253701 12831 254501
rect 13011 253701 13041 254501
rect 13221 253701 13251 254501
rect 13431 253701 13461 254501
rect 13641 253701 13671 254501
rect 13851 253701 13881 254501
rect 14061 253701 14091 254501
rect 14271 253701 14301 254501
rect 14481 253701 14511 254501
rect 14691 253701 14721 254501
rect 14901 253701 14931 254501
rect 15111 253701 15141 254501
rect 15321 253701 15351 254501
rect 15531 253701 15561 254501
rect 15741 253701 15771 254501
rect 15951 253701 15981 254501
rect 16161 253701 16191 254501
rect 16371 253701 16401 254501
rect 16581 253701 16611 254501
rect 16791 253701 16821 254501
rect 17001 253701 17031 254501
rect 17211 253701 17241 254501
rect 17421 253701 17451 254501
rect 17631 253701 17661 254501
rect 17841 253701 17871 254501
rect 18051 253701 18081 254501
rect 18261 253701 18291 254501
rect 18471 253701 18501 254501
rect 18681 253701 18711 254501
rect 18891 253701 18921 254501
rect 19101 253701 19131 254501
rect 19311 253701 19341 254501
rect 19521 253701 19551 254501
rect 19731 253701 19761 254501
rect 19941 253701 19971 254501
rect 20151 253701 20181 254501
rect 20361 253701 20391 254501
rect 20571 253701 20601 254501
rect 20781 253701 20811 254501
rect 20991 253701 21021 254501
rect 21201 253701 21231 254501
rect 21411 253701 21441 254501
rect 21621 253701 21651 254501
rect 21831 253701 21861 254501
rect 22041 253701 22071 254501
rect 22251 253701 22281 254501
rect 22461 253701 22491 254501
rect 22671 253701 22701 254501
rect 22881 253701 22911 254501
rect 23091 253701 23121 254501
rect 23301 253701 23331 254501
rect 23511 253701 23541 254501
rect 23721 253701 23751 254501
rect 23931 253701 23961 254501
rect 24141 253701 24171 254501
rect 24351 253701 24381 254501
rect 24561 253701 24591 254501
rect 24771 253701 24801 254501
rect 24981 253701 25011 254501
rect 25191 253701 25221 254501
rect 25401 253701 25431 254501
rect 25611 253701 25641 254501
rect 25821 253701 25851 254501
rect 26031 253701 26061 254501
rect 26241 253701 26271 254501
rect 26451 253701 26481 254501
rect 26661 253701 26691 254501
rect 26871 253701 26901 254501
rect 27081 253701 27111 254501
rect 27291 253701 27321 254501
rect -3999 252665 -3969 253465
rect -3789 252665 -3759 253465
rect -3579 252665 -3549 253465
rect -3369 252665 -3339 253465
rect -3159 252665 -3129 253465
rect -2949 252665 -2919 253465
rect -2739 252665 -2709 253465
rect -2529 252665 -2499 253465
rect -2319 252665 -2289 253465
rect -2109 252665 -2079 253465
rect -1899 252665 -1869 253465
rect -1689 252665 -1659 253465
rect -1479 252665 -1449 253465
rect -1269 252665 -1239 253465
rect -1059 252665 -1029 253465
rect -849 252665 -819 253465
rect -639 252665 -609 253465
rect -429 252665 -399 253465
rect -219 252665 -189 253465
rect -9 252665 21 253465
rect 201 252665 231 253465
rect 411 252665 441 253465
rect 621 252665 651 253465
rect 831 252665 861 253465
rect 1041 252665 1071 253465
rect 1251 252665 1281 253465
rect 1461 252665 1491 253465
rect 1671 252665 1701 253465
rect 1881 252665 1911 253465
rect 2091 252665 2121 253465
rect 2301 252665 2331 253465
rect 2511 252665 2541 253465
rect 2721 252665 2751 253465
rect 2931 252665 2961 253465
rect 3141 252665 3171 253465
rect 3351 252665 3381 253465
rect 3561 252665 3591 253465
rect 3771 252665 3801 253465
rect 3981 252665 4011 253465
rect 4191 252665 4221 253465
rect 4401 252665 4431 253465
rect 4611 252665 4641 253465
rect 4821 252665 4851 253465
rect 5031 252665 5061 253465
rect 5241 252665 5271 253465
rect 5451 252665 5481 253465
rect 5661 252665 5691 253465
rect 5871 252665 5901 253465
rect 6081 252665 6111 253465
rect 6291 252665 6321 253465
rect 6501 252665 6531 253465
rect 6711 252665 6741 253465
rect 6921 252665 6951 253465
rect 7131 252665 7161 253465
rect 7341 252665 7371 253465
rect 7551 252665 7581 253465
rect 7761 252665 7791 253465
rect 7971 252665 8001 253465
rect 8181 252665 8211 253465
rect 8391 252665 8421 253465
rect 8601 252665 8631 253465
rect 8811 252665 8841 253465
rect 9021 252665 9051 253465
rect 9231 252665 9261 253465
rect 9441 252665 9471 253465
rect 9651 252665 9681 253465
rect 9861 252665 9891 253465
rect 10071 252665 10101 253465
rect 10281 252665 10311 253465
rect 10491 252665 10521 253465
rect 10701 252665 10731 253465
rect 10911 252665 10941 253465
rect 11121 252665 11151 253465
rect 11331 252665 11361 253465
rect 11541 252665 11571 253465
rect 11751 252665 11781 253465
rect 11961 252665 11991 253465
rect 12171 252665 12201 253465
rect 12381 252665 12411 253465
rect 12591 252665 12621 253465
rect 12801 252665 12831 253465
rect 13011 252665 13041 253465
rect 13221 252665 13251 253465
rect 13431 252665 13461 253465
rect 13641 252665 13671 253465
rect 13851 252665 13881 253465
rect 14061 252665 14091 253465
rect 14271 252665 14301 253465
rect 14481 252665 14511 253465
rect 14691 252665 14721 253465
rect 14901 252665 14931 253465
rect 15111 252665 15141 253465
rect 15321 252665 15351 253465
rect 15531 252665 15561 253465
rect 15741 252665 15771 253465
rect 15951 252665 15981 253465
rect 16161 252665 16191 253465
rect 16371 252665 16401 253465
rect 16581 252665 16611 253465
rect 16791 252665 16821 253465
rect 17001 252665 17031 253465
rect 17211 252665 17241 253465
rect 17421 252665 17451 253465
rect 17631 252665 17661 253465
rect 17841 252665 17871 253465
rect 18051 252665 18081 253465
rect 18261 252665 18291 253465
rect 18471 252665 18501 253465
rect 18681 252665 18711 253465
rect 18891 252665 18921 253465
rect 19101 252665 19131 253465
rect 19311 252665 19341 253465
rect 19521 252665 19551 253465
rect 19731 252665 19761 253465
rect 19941 252665 19971 253465
rect 20151 252665 20181 253465
rect 20361 252665 20391 253465
rect 20571 252665 20601 253465
rect 20781 252665 20811 253465
rect 20991 252665 21021 253465
rect 21201 252665 21231 253465
rect 21411 252665 21441 253465
rect 21621 252665 21651 253465
rect 21831 252665 21861 253465
rect 22041 252665 22071 253465
rect 22251 252665 22281 253465
rect 22461 252665 22491 253465
rect 22671 252665 22701 253465
rect 22881 252665 22911 253465
rect 23091 252665 23121 253465
rect 23301 252665 23331 253465
rect 23511 252665 23541 253465
rect 23721 252665 23751 253465
rect 23931 252665 23961 253465
rect 24141 252665 24171 253465
rect 24351 252665 24381 253465
rect 24561 252665 24591 253465
rect 24771 252665 24801 253465
rect 24981 252665 25011 253465
rect 25191 252665 25221 253465
rect 25401 252665 25431 253465
rect 25611 252665 25641 253465
rect 25821 252665 25851 253465
rect 26031 252665 26061 253465
rect 26241 252665 26271 253465
rect 26451 252665 26481 253465
rect 26661 252665 26691 253465
rect 26871 252665 26901 253465
rect 27081 252665 27111 253465
rect 27291 252665 27321 253465
rect -3999 251629 -3969 252429
rect -3789 251629 -3759 252429
rect -3579 251629 -3549 252429
rect -3369 251629 -3339 252429
rect -3159 251629 -3129 252429
rect -2949 251629 -2919 252429
rect -2739 251629 -2709 252429
rect -2529 251629 -2499 252429
rect -2319 251629 -2289 252429
rect -2109 251629 -2079 252429
rect -1899 251629 -1869 252429
rect -1689 251629 -1659 252429
rect -1479 251629 -1449 252429
rect -1269 251629 -1239 252429
rect -1059 251629 -1029 252429
rect -849 251629 -819 252429
rect -639 251629 -609 252429
rect -429 251629 -399 252429
rect -219 251629 -189 252429
rect -9 251629 21 252429
rect 201 251629 231 252429
rect 411 251629 441 252429
rect 621 251629 651 252429
rect 831 251629 861 252429
rect 1041 251629 1071 252429
rect 1251 251629 1281 252429
rect 1461 251629 1491 252429
rect 1671 251629 1701 252429
rect 1881 251629 1911 252429
rect 2091 251629 2121 252429
rect 2301 251629 2331 252429
rect 2511 251629 2541 252429
rect 2721 251629 2751 252429
rect 2931 251629 2961 252429
rect 3141 251629 3171 252429
rect 3351 251629 3381 252429
rect 3561 251629 3591 252429
rect 3771 251629 3801 252429
rect 3981 251629 4011 252429
rect 4191 251629 4221 252429
rect 4401 251629 4431 252429
rect 4611 251629 4641 252429
rect 4821 251629 4851 252429
rect 5031 251629 5061 252429
rect 5241 251629 5271 252429
rect 5451 251629 5481 252429
rect 5661 251629 5691 252429
rect 5871 251629 5901 252429
rect 6081 251629 6111 252429
rect 6291 251629 6321 252429
rect 6501 251629 6531 252429
rect 6711 251629 6741 252429
rect 6921 251629 6951 252429
rect 7131 251629 7161 252429
rect 7341 251629 7371 252429
rect 7551 251629 7581 252429
rect 7761 251629 7791 252429
rect 7971 251629 8001 252429
rect 8181 251629 8211 252429
rect 8391 251629 8421 252429
rect 8601 251629 8631 252429
rect 8811 251629 8841 252429
rect 9021 251629 9051 252429
rect 9231 251629 9261 252429
rect 9441 251629 9471 252429
rect 9651 251629 9681 252429
rect 9861 251629 9891 252429
rect 10071 251629 10101 252429
rect 10281 251629 10311 252429
rect 10491 251629 10521 252429
rect 10701 251629 10731 252429
rect 10911 251629 10941 252429
rect 11121 251629 11151 252429
rect 11331 251629 11361 252429
rect 11541 251629 11571 252429
rect 11751 251629 11781 252429
rect 11961 251629 11991 252429
rect 12171 251629 12201 252429
rect 12381 251629 12411 252429
rect 12591 251629 12621 252429
rect 12801 251629 12831 252429
rect 13011 251629 13041 252429
rect 13221 251629 13251 252429
rect 13431 251629 13461 252429
rect 13641 251629 13671 252429
rect 13851 251629 13881 252429
rect 14061 251629 14091 252429
rect 14271 251629 14301 252429
rect 14481 251629 14511 252429
rect 14691 251629 14721 252429
rect 14901 251629 14931 252429
rect 15111 251629 15141 252429
rect 15321 251629 15351 252429
rect 15531 251629 15561 252429
rect 15741 251629 15771 252429
rect 15951 251629 15981 252429
rect 16161 251629 16191 252429
rect 16371 251629 16401 252429
rect 16581 251629 16611 252429
rect 16791 251629 16821 252429
rect 17001 251629 17031 252429
rect 17211 251629 17241 252429
rect 17421 251629 17451 252429
rect 17631 251629 17661 252429
rect 17841 251629 17871 252429
rect 18051 251629 18081 252429
rect 18261 251629 18291 252429
rect 18471 251629 18501 252429
rect 18681 251629 18711 252429
rect 18891 251629 18921 252429
rect 19101 251629 19131 252429
rect 19311 251629 19341 252429
rect 19521 251629 19551 252429
rect 19731 251629 19761 252429
rect 19941 251629 19971 252429
rect 20151 251629 20181 252429
rect 20361 251629 20391 252429
rect 20571 251629 20601 252429
rect 20781 251629 20811 252429
rect 20991 251629 21021 252429
rect 21201 251629 21231 252429
rect 21411 251629 21441 252429
rect 21621 251629 21651 252429
rect 21831 251629 21861 252429
rect 22041 251629 22071 252429
rect 22251 251629 22281 252429
rect 22461 251629 22491 252429
rect 22671 251629 22701 252429
rect 22881 251629 22911 252429
rect 23091 251629 23121 252429
rect 23301 251629 23331 252429
rect 23511 251629 23541 252429
rect 23721 251629 23751 252429
rect 23931 251629 23961 252429
rect 24141 251629 24171 252429
rect 24351 251629 24381 252429
rect 24561 251629 24591 252429
rect 24771 251629 24801 252429
rect 24981 251629 25011 252429
rect 25191 251629 25221 252429
rect 25401 251629 25431 252429
rect 25611 251629 25641 252429
rect 25821 251629 25851 252429
rect 26031 251629 26061 252429
rect 26241 251629 26271 252429
rect 26451 251629 26481 252429
rect 26661 251629 26691 252429
rect 26871 251629 26901 252429
rect 27081 251629 27111 252429
rect 27291 251629 27321 252429
rect -3999 250593 -3969 251393
rect -3789 250593 -3759 251393
rect -3579 250593 -3549 251393
rect -3369 250593 -3339 251393
rect -3159 250593 -3129 251393
rect -2949 250593 -2919 251393
rect -2739 250593 -2709 251393
rect -2529 250593 -2499 251393
rect -2319 250593 -2289 251393
rect -2109 250593 -2079 251393
rect -1899 250593 -1869 251393
rect -1689 250593 -1659 251393
rect -1479 250593 -1449 251393
rect -1269 250593 -1239 251393
rect -1059 250593 -1029 251393
rect -849 250593 -819 251393
rect -639 250593 -609 251393
rect -429 250593 -399 251393
rect -219 250593 -189 251393
rect -9 250593 21 251393
rect 201 250593 231 251393
rect 411 250593 441 251393
rect 621 250593 651 251393
rect 831 250593 861 251393
rect 1041 250593 1071 251393
rect 1251 250593 1281 251393
rect 1461 250593 1491 251393
rect 1671 250593 1701 251393
rect 1881 250593 1911 251393
rect 2091 250593 2121 251393
rect 2301 250593 2331 251393
rect 2511 250593 2541 251393
rect 2721 250593 2751 251393
rect 2931 250593 2961 251393
rect 3141 250593 3171 251393
rect 3351 250593 3381 251393
rect 3561 250593 3591 251393
rect 3771 250593 3801 251393
rect 3981 250593 4011 251393
rect 4191 250593 4221 251393
rect 4401 250593 4431 251393
rect 4611 250593 4641 251393
rect 4821 250593 4851 251393
rect 5031 250593 5061 251393
rect 5241 250593 5271 251393
rect 5451 250593 5481 251393
rect 5661 250593 5691 251393
rect 5871 250593 5901 251393
rect 6081 250593 6111 251393
rect 6291 250593 6321 251393
rect 6501 250593 6531 251393
rect 6711 250593 6741 251393
rect 6921 250593 6951 251393
rect 7131 250593 7161 251393
rect 7341 250593 7371 251393
rect 7551 250593 7581 251393
rect 7761 250593 7791 251393
rect 7971 250593 8001 251393
rect 8181 250593 8211 251393
rect 8391 250593 8421 251393
rect 8601 250593 8631 251393
rect 8811 250593 8841 251393
rect 9021 250593 9051 251393
rect 9231 250593 9261 251393
rect 9441 250593 9471 251393
rect 9651 250593 9681 251393
rect 9861 250593 9891 251393
rect 10071 250593 10101 251393
rect 10281 250593 10311 251393
rect 10491 250593 10521 251393
rect 10701 250593 10731 251393
rect 10911 250593 10941 251393
rect 11121 250593 11151 251393
rect 11331 250593 11361 251393
rect 11541 250593 11571 251393
rect 11751 250593 11781 251393
rect 11961 250593 11991 251393
rect 12171 250593 12201 251393
rect 12381 250593 12411 251393
rect 12591 250593 12621 251393
rect 12801 250593 12831 251393
rect 13011 250593 13041 251393
rect 13221 250593 13251 251393
rect 13431 250593 13461 251393
rect 13641 250593 13671 251393
rect 13851 250593 13881 251393
rect 14061 250593 14091 251393
rect 14271 250593 14301 251393
rect 14481 250593 14511 251393
rect 14691 250593 14721 251393
rect 14901 250593 14931 251393
rect 15111 250593 15141 251393
rect 15321 250593 15351 251393
rect 15531 250593 15561 251393
rect 15741 250593 15771 251393
rect 15951 250593 15981 251393
rect 16161 250593 16191 251393
rect 16371 250593 16401 251393
rect 16581 250593 16611 251393
rect 16791 250593 16821 251393
rect 17001 250593 17031 251393
rect 17211 250593 17241 251393
rect 17421 250593 17451 251393
rect 17631 250593 17661 251393
rect 17841 250593 17871 251393
rect 18051 250593 18081 251393
rect 18261 250593 18291 251393
rect 18471 250593 18501 251393
rect 18681 250593 18711 251393
rect 18891 250593 18921 251393
rect 19101 250593 19131 251393
rect 19311 250593 19341 251393
rect 19521 250593 19551 251393
rect 19731 250593 19761 251393
rect 19941 250593 19971 251393
rect 20151 250593 20181 251393
rect 20361 250593 20391 251393
rect 20571 250593 20601 251393
rect 20781 250593 20811 251393
rect 20991 250593 21021 251393
rect 21201 250593 21231 251393
rect 21411 250593 21441 251393
rect 21621 250593 21651 251393
rect 21831 250593 21861 251393
rect 22041 250593 22071 251393
rect 22251 250593 22281 251393
rect 22461 250593 22491 251393
rect 22671 250593 22701 251393
rect 22881 250593 22911 251393
rect 23091 250593 23121 251393
rect 23301 250593 23331 251393
rect 23511 250593 23541 251393
rect 23721 250593 23751 251393
rect 23931 250593 23961 251393
rect 24141 250593 24171 251393
rect 24351 250593 24381 251393
rect 24561 250593 24591 251393
rect 24771 250593 24801 251393
rect 24981 250593 25011 251393
rect 25191 250593 25221 251393
rect 25401 250593 25431 251393
rect 25611 250593 25641 251393
rect 25821 250593 25851 251393
rect 26031 250593 26061 251393
rect 26241 250593 26271 251393
rect 26451 250593 26481 251393
rect 26661 250593 26691 251393
rect 26871 250593 26901 251393
rect 27081 250593 27111 251393
rect 27291 250593 27321 251393
rect -3999 249557 -3969 250357
rect -3789 249557 -3759 250357
rect -3579 249557 -3549 250357
rect -3369 249557 -3339 250357
rect -3159 249557 -3129 250357
rect -2949 249557 -2919 250357
rect -2739 249557 -2709 250357
rect -2529 249557 -2499 250357
rect -2319 249557 -2289 250357
rect -2109 249557 -2079 250357
rect -1899 249557 -1869 250357
rect -1689 249557 -1659 250357
rect -1479 249557 -1449 250357
rect -1269 249557 -1239 250357
rect -1059 249557 -1029 250357
rect -849 249557 -819 250357
rect -639 249557 -609 250357
rect -429 249557 -399 250357
rect -219 249557 -189 250357
rect -9 249557 21 250357
rect 201 249557 231 250357
rect 411 249557 441 250357
rect 621 249557 651 250357
rect 831 249557 861 250357
rect 1041 249557 1071 250357
rect 1251 249557 1281 250357
rect 1461 249557 1491 250357
rect 1671 249557 1701 250357
rect 1881 249557 1911 250357
rect 2091 249557 2121 250357
rect 2301 249557 2331 250357
rect 2511 249557 2541 250357
rect 2721 249557 2751 250357
rect 2931 249557 2961 250357
rect 3141 249557 3171 250357
rect 3351 249557 3381 250357
rect 3561 249557 3591 250357
rect 3771 249557 3801 250357
rect 3981 249557 4011 250357
rect 4191 249557 4221 250357
rect 4401 249557 4431 250357
rect 4611 249557 4641 250357
rect 4821 249557 4851 250357
rect 5031 249557 5061 250357
rect 5241 249557 5271 250357
rect 5451 249557 5481 250357
rect 5661 249557 5691 250357
rect 5871 249557 5901 250357
rect 6081 249557 6111 250357
rect 6291 249557 6321 250357
rect 6501 249557 6531 250357
rect 6711 249557 6741 250357
rect 6921 249557 6951 250357
rect 7131 249557 7161 250357
rect 7341 249557 7371 250357
rect 7551 249557 7581 250357
rect 7761 249557 7791 250357
rect 7971 249557 8001 250357
rect 8181 249557 8211 250357
rect 8391 249557 8421 250357
rect 8601 249557 8631 250357
rect 8811 249557 8841 250357
rect 9021 249557 9051 250357
rect 9231 249557 9261 250357
rect 9441 249557 9471 250357
rect 9651 249557 9681 250357
rect 9861 249557 9891 250357
rect 10071 249557 10101 250357
rect 10281 249557 10311 250357
rect 10491 249557 10521 250357
rect 10701 249557 10731 250357
rect 10911 249557 10941 250357
rect 11121 249557 11151 250357
rect 11331 249557 11361 250357
rect 11541 249557 11571 250357
rect 11751 249557 11781 250357
rect 11961 249557 11991 250357
rect 12171 249557 12201 250357
rect 12381 249557 12411 250357
rect 12591 249557 12621 250357
rect 12801 249557 12831 250357
rect 13011 249557 13041 250357
rect 13221 249557 13251 250357
rect 13431 249557 13461 250357
rect 13641 249557 13671 250357
rect 13851 249557 13881 250357
rect 14061 249557 14091 250357
rect 14271 249557 14301 250357
rect 14481 249557 14511 250357
rect 14691 249557 14721 250357
rect 14901 249557 14931 250357
rect 15111 249557 15141 250357
rect 15321 249557 15351 250357
rect 15531 249557 15561 250357
rect 15741 249557 15771 250357
rect 15951 249557 15981 250357
rect 16161 249557 16191 250357
rect 16371 249557 16401 250357
rect 16581 249557 16611 250357
rect 16791 249557 16821 250357
rect 17001 249557 17031 250357
rect 17211 249557 17241 250357
rect 17421 249557 17451 250357
rect 17631 249557 17661 250357
rect 17841 249557 17871 250357
rect 18051 249557 18081 250357
rect 18261 249557 18291 250357
rect 18471 249557 18501 250357
rect 18681 249557 18711 250357
rect 18891 249557 18921 250357
rect 19101 249557 19131 250357
rect 19311 249557 19341 250357
rect 19521 249557 19551 250357
rect 19731 249557 19761 250357
rect 19941 249557 19971 250357
rect 20151 249557 20181 250357
rect 20361 249557 20391 250357
rect 20571 249557 20601 250357
rect 20781 249557 20811 250357
rect 20991 249557 21021 250357
rect 21201 249557 21231 250357
rect 21411 249557 21441 250357
rect 21621 249557 21651 250357
rect 21831 249557 21861 250357
rect 22041 249557 22071 250357
rect 22251 249557 22281 250357
rect 22461 249557 22491 250357
rect 22671 249557 22701 250357
rect 22881 249557 22911 250357
rect 23091 249557 23121 250357
rect 23301 249557 23331 250357
rect 23511 249557 23541 250357
rect 23721 249557 23751 250357
rect 23931 249557 23961 250357
rect 24141 249557 24171 250357
rect 24351 249557 24381 250357
rect 24561 249557 24591 250357
rect 24771 249557 24801 250357
rect 24981 249557 25011 250357
rect 25191 249557 25221 250357
rect 25401 249557 25431 250357
rect 25611 249557 25641 250357
rect 25821 249557 25851 250357
rect 26031 249557 26061 250357
rect 26241 249557 26271 250357
rect 26451 249557 26481 250357
rect 26661 249557 26691 250357
rect 26871 249557 26901 250357
rect 27081 249557 27111 250357
rect 27291 249557 27321 250357
rect -3999 248392 -3969 249192
rect -3789 248392 -3759 249192
rect -3579 248392 -3549 249192
rect -3369 248392 -3339 249192
rect -3159 248392 -3129 249192
rect -2949 248392 -2919 249192
rect -2739 248392 -2709 249192
rect -2529 248392 -2499 249192
rect -2319 248392 -2289 249192
rect -2109 248392 -2079 249192
rect -1899 248392 -1869 249192
rect -1689 248392 -1659 249192
rect -1479 248392 -1449 249192
rect -1269 248392 -1239 249192
rect -1059 248392 -1029 249192
rect -849 248392 -819 249192
rect -639 248392 -609 249192
rect -429 248392 -399 249192
rect -219 248392 -189 249192
rect -9 248392 21 249192
rect 201 248392 231 249192
rect 411 248392 441 249192
rect 621 248392 651 249192
rect 831 248392 861 249192
rect 1041 248392 1071 249192
rect 1251 248392 1281 249192
rect 1461 248392 1491 249192
rect 1671 248392 1701 249192
rect 1881 248392 1911 249192
rect 2091 248392 2121 249192
rect 2301 248392 2331 249192
rect 2511 248392 2541 249192
rect 2721 248392 2751 249192
rect 2931 248392 2961 249192
rect 3141 248392 3171 249192
rect 3351 248392 3381 249192
rect 3561 248392 3591 249192
rect 3771 248392 3801 249192
rect 3981 248392 4011 249192
rect 4191 248392 4221 249192
rect 4401 248392 4431 249192
rect 4611 248392 4641 249192
rect 4821 248392 4851 249192
rect 5031 248392 5061 249192
rect 5241 248392 5271 249192
rect 5451 248392 5481 249192
rect 5661 248392 5691 249192
rect 5871 248392 5901 249192
rect 6081 248392 6111 249192
rect 6291 248392 6321 249192
rect 6501 248392 6531 249192
rect 6711 248392 6741 249192
rect 6921 248392 6951 249192
rect 7131 248392 7161 249192
rect 7341 248392 7371 249192
rect 7551 248392 7581 249192
rect 7761 248392 7791 249192
rect 7971 248392 8001 249192
rect 8181 248392 8211 249192
rect 8391 248392 8421 249192
rect 8601 248392 8631 249192
rect 8811 248392 8841 249192
rect 9021 248392 9051 249192
rect 9231 248392 9261 249192
rect 9441 248392 9471 249192
rect 9651 248392 9681 249192
rect 9861 248392 9891 249192
rect 10071 248392 10101 249192
rect 10281 248392 10311 249192
rect 10491 248392 10521 249192
rect 10701 248392 10731 249192
rect 10911 248392 10941 249192
rect 11121 248392 11151 249192
rect 11331 248392 11361 249192
rect 11541 248392 11571 249192
rect 11751 248392 11781 249192
rect 11961 248392 11991 249192
rect 12171 248392 12201 249192
rect 12381 248392 12411 249192
rect 12591 248392 12621 249192
rect 12801 248392 12831 249192
rect 13011 248392 13041 249192
rect 13221 248392 13251 249192
rect 13431 248392 13461 249192
rect 13641 248392 13671 249192
rect 13851 248392 13881 249192
rect 14061 248392 14091 249192
rect 14271 248392 14301 249192
rect 14481 248392 14511 249192
rect 14691 248392 14721 249192
rect 14901 248392 14931 249192
rect 15111 248392 15141 249192
rect 15321 248392 15351 249192
rect 15531 248392 15561 249192
rect 15741 248392 15771 249192
rect 15951 248392 15981 249192
rect 16161 248392 16191 249192
rect 16371 248392 16401 249192
rect 16581 248392 16611 249192
rect 16791 248392 16821 249192
rect 17001 248392 17031 249192
rect 17211 248392 17241 249192
rect 17421 248392 17451 249192
rect 17631 248392 17661 249192
rect 17841 248392 17871 249192
rect 18051 248392 18081 249192
rect 18261 248392 18291 249192
rect 18471 248392 18501 249192
rect 18681 248392 18711 249192
rect 18891 248392 18921 249192
rect 19101 248392 19131 249192
rect 19311 248392 19341 249192
rect 19521 248392 19551 249192
rect 19731 248392 19761 249192
rect 19941 248392 19971 249192
rect 20151 248392 20181 249192
rect 20361 248392 20391 249192
rect 20571 248392 20601 249192
rect 20781 248392 20811 249192
rect 20991 248392 21021 249192
rect 21201 248392 21231 249192
rect 21411 248392 21441 249192
rect 21621 248392 21651 249192
rect 21831 248392 21861 249192
rect 22041 248392 22071 249192
rect 22251 248392 22281 249192
rect 22461 248392 22491 249192
rect 22671 248392 22701 249192
rect 22881 248392 22911 249192
rect 23091 248392 23121 249192
rect 23301 248392 23331 249192
rect 23511 248392 23541 249192
rect 23721 248392 23751 249192
rect 23931 248392 23961 249192
rect 24141 248392 24171 249192
rect 24351 248392 24381 249192
rect 24561 248392 24591 249192
rect 24771 248392 24801 249192
rect 24981 248392 25011 249192
rect 25191 248392 25221 249192
rect 25401 248392 25431 249192
rect 25611 248392 25641 249192
rect 25821 248392 25851 249192
rect 26031 248392 26061 249192
rect 26241 248392 26271 249192
rect 26451 248392 26481 249192
rect 26661 248392 26691 249192
rect 26871 248392 26901 249192
rect 27081 248392 27111 249192
rect 27291 248392 27321 249192
rect -3999 247356 -3969 248156
rect -3789 247356 -3759 248156
rect -3579 247356 -3549 248156
rect -3369 247356 -3339 248156
rect -3159 247356 -3129 248156
rect -2949 247356 -2919 248156
rect -2739 247356 -2709 248156
rect -2529 247356 -2499 248156
rect -2319 247356 -2289 248156
rect -2109 247356 -2079 248156
rect -1899 247356 -1869 248156
rect -1689 247356 -1659 248156
rect -1479 247356 -1449 248156
rect -1269 247356 -1239 248156
rect -1059 247356 -1029 248156
rect -849 247356 -819 248156
rect -639 247356 -609 248156
rect -429 247356 -399 248156
rect -219 247356 -189 248156
rect -9 247356 21 248156
rect 201 247356 231 248156
rect 411 247356 441 248156
rect 621 247356 651 248156
rect 831 247356 861 248156
rect 1041 247356 1071 248156
rect 1251 247356 1281 248156
rect 1461 247356 1491 248156
rect 1671 247356 1701 248156
rect 1881 247356 1911 248156
rect 2091 247356 2121 248156
rect 2301 247356 2331 248156
rect 2511 247356 2541 248156
rect 2721 247356 2751 248156
rect 2931 247356 2961 248156
rect 3141 247356 3171 248156
rect 3351 247356 3381 248156
rect 3561 247356 3591 248156
rect 3771 247356 3801 248156
rect 3981 247356 4011 248156
rect 4191 247356 4221 248156
rect 4401 247356 4431 248156
rect 4611 247356 4641 248156
rect 4821 247356 4851 248156
rect 5031 247356 5061 248156
rect 5241 247356 5271 248156
rect 5451 247356 5481 248156
rect 5661 247356 5691 248156
rect 5871 247356 5901 248156
rect 6081 247356 6111 248156
rect 6291 247356 6321 248156
rect 6501 247356 6531 248156
rect 6711 247356 6741 248156
rect 6921 247356 6951 248156
rect 7131 247356 7161 248156
rect 7341 247356 7371 248156
rect 7551 247356 7581 248156
rect 7761 247356 7791 248156
rect 7971 247356 8001 248156
rect 8181 247356 8211 248156
rect 8391 247356 8421 248156
rect 8601 247356 8631 248156
rect 8811 247356 8841 248156
rect 9021 247356 9051 248156
rect 9231 247356 9261 248156
rect 9441 247356 9471 248156
rect 9651 247356 9681 248156
rect 9861 247356 9891 248156
rect 10071 247356 10101 248156
rect 10281 247356 10311 248156
rect 10491 247356 10521 248156
rect 10701 247356 10731 248156
rect 10911 247356 10941 248156
rect 11121 247356 11151 248156
rect 11331 247356 11361 248156
rect 11541 247356 11571 248156
rect 11751 247356 11781 248156
rect 11961 247356 11991 248156
rect 12171 247356 12201 248156
rect 12381 247356 12411 248156
rect 12591 247356 12621 248156
rect 12801 247356 12831 248156
rect 13011 247356 13041 248156
rect 13221 247356 13251 248156
rect 13431 247356 13461 248156
rect 13641 247356 13671 248156
rect 13851 247356 13881 248156
rect 14061 247356 14091 248156
rect 14271 247356 14301 248156
rect 14481 247356 14511 248156
rect 14691 247356 14721 248156
rect 14901 247356 14931 248156
rect 15111 247356 15141 248156
rect 15321 247356 15351 248156
rect 15531 247356 15561 248156
rect 15741 247356 15771 248156
rect 15951 247356 15981 248156
rect 16161 247356 16191 248156
rect 16371 247356 16401 248156
rect 16581 247356 16611 248156
rect 16791 247356 16821 248156
rect 17001 247356 17031 248156
rect 17211 247356 17241 248156
rect 17421 247356 17451 248156
rect 17631 247356 17661 248156
rect 17841 247356 17871 248156
rect 18051 247356 18081 248156
rect 18261 247356 18291 248156
rect 18471 247356 18501 248156
rect 18681 247356 18711 248156
rect 18891 247356 18921 248156
rect 19101 247356 19131 248156
rect 19311 247356 19341 248156
rect 19521 247356 19551 248156
rect 19731 247356 19761 248156
rect 19941 247356 19971 248156
rect 20151 247356 20181 248156
rect 20361 247356 20391 248156
rect 20571 247356 20601 248156
rect 20781 247356 20811 248156
rect 20991 247356 21021 248156
rect 21201 247356 21231 248156
rect 21411 247356 21441 248156
rect 21621 247356 21651 248156
rect 21831 247356 21861 248156
rect 22041 247356 22071 248156
rect 22251 247356 22281 248156
rect 22461 247356 22491 248156
rect 22671 247356 22701 248156
rect 22881 247356 22911 248156
rect 23091 247356 23121 248156
rect 23301 247356 23331 248156
rect 23511 247356 23541 248156
rect 23721 247356 23751 248156
rect 23931 247356 23961 248156
rect 24141 247356 24171 248156
rect 24351 247356 24381 248156
rect 24561 247356 24591 248156
rect 24771 247356 24801 248156
rect 24981 247356 25011 248156
rect 25191 247356 25221 248156
rect 25401 247356 25431 248156
rect 25611 247356 25641 248156
rect 25821 247356 25851 248156
rect 26031 247356 26061 248156
rect 26241 247356 26271 248156
rect 26451 247356 26481 248156
rect 26661 247356 26691 248156
rect 26871 247356 26901 248156
rect 27081 247356 27111 248156
rect 27291 247356 27321 248156
rect -3999 246320 -3969 247120
rect -3789 246320 -3759 247120
rect -3579 246320 -3549 247120
rect -3369 246320 -3339 247120
rect -3159 246320 -3129 247120
rect -2949 246320 -2919 247120
rect -2739 246320 -2709 247120
rect -2529 246320 -2499 247120
rect -2319 246320 -2289 247120
rect -2109 246320 -2079 247120
rect -1899 246320 -1869 247120
rect -1689 246320 -1659 247120
rect -1479 246320 -1449 247120
rect -1269 246320 -1239 247120
rect -1059 246320 -1029 247120
rect -849 246320 -819 247120
rect -639 246320 -609 247120
rect -429 246320 -399 247120
rect -219 246320 -189 247120
rect -9 246320 21 247120
rect 201 246320 231 247120
rect 411 246320 441 247120
rect 621 246320 651 247120
rect 831 246320 861 247120
rect 1041 246320 1071 247120
rect 1251 246320 1281 247120
rect 1461 246320 1491 247120
rect 1671 246320 1701 247120
rect 1881 246320 1911 247120
rect 2091 246320 2121 247120
rect 2301 246320 2331 247120
rect 2511 246320 2541 247120
rect 2721 246320 2751 247120
rect 2931 246320 2961 247120
rect 3141 246320 3171 247120
rect 3351 246320 3381 247120
rect 3561 246320 3591 247120
rect 3771 246320 3801 247120
rect 3981 246320 4011 247120
rect 4191 246320 4221 247120
rect 4401 246320 4431 247120
rect 4611 246320 4641 247120
rect 4821 246320 4851 247120
rect 5031 246320 5061 247120
rect 5241 246320 5271 247120
rect 5451 246320 5481 247120
rect 5661 246320 5691 247120
rect 5871 246320 5901 247120
rect 6081 246320 6111 247120
rect 6291 246320 6321 247120
rect 6501 246320 6531 247120
rect 6711 246320 6741 247120
rect 6921 246320 6951 247120
rect 7131 246320 7161 247120
rect 7341 246320 7371 247120
rect 7551 246320 7581 247120
rect 7761 246320 7791 247120
rect 7971 246320 8001 247120
rect 8181 246320 8211 247120
rect 8391 246320 8421 247120
rect 8601 246320 8631 247120
rect 8811 246320 8841 247120
rect 9021 246320 9051 247120
rect 9231 246320 9261 247120
rect 9441 246320 9471 247120
rect 9651 246320 9681 247120
rect 9861 246320 9891 247120
rect 10071 246320 10101 247120
rect 10281 246320 10311 247120
rect 10491 246320 10521 247120
rect 10701 246320 10731 247120
rect 10911 246320 10941 247120
rect 11121 246320 11151 247120
rect 11331 246320 11361 247120
rect 11541 246320 11571 247120
rect 11751 246320 11781 247120
rect 11961 246320 11991 247120
rect 12171 246320 12201 247120
rect 12381 246320 12411 247120
rect 12591 246320 12621 247120
rect 12801 246320 12831 247120
rect 13011 246320 13041 247120
rect 13221 246320 13251 247120
rect 13431 246320 13461 247120
rect 13641 246320 13671 247120
rect 13851 246320 13881 247120
rect 14061 246320 14091 247120
rect 14271 246320 14301 247120
rect 14481 246320 14511 247120
rect 14691 246320 14721 247120
rect 14901 246320 14931 247120
rect 15111 246320 15141 247120
rect 15321 246320 15351 247120
rect 15531 246320 15561 247120
rect 15741 246320 15771 247120
rect 15951 246320 15981 247120
rect 16161 246320 16191 247120
rect 16371 246320 16401 247120
rect 16581 246320 16611 247120
rect 16791 246320 16821 247120
rect 17001 246320 17031 247120
rect 17211 246320 17241 247120
rect 17421 246320 17451 247120
rect 17631 246320 17661 247120
rect 17841 246320 17871 247120
rect 18051 246320 18081 247120
rect 18261 246320 18291 247120
rect 18471 246320 18501 247120
rect 18681 246320 18711 247120
rect 18891 246320 18921 247120
rect 19101 246320 19131 247120
rect 19311 246320 19341 247120
rect 19521 246320 19551 247120
rect 19731 246320 19761 247120
rect 19941 246320 19971 247120
rect 20151 246320 20181 247120
rect 20361 246320 20391 247120
rect 20571 246320 20601 247120
rect 20781 246320 20811 247120
rect 20991 246320 21021 247120
rect 21201 246320 21231 247120
rect 21411 246320 21441 247120
rect 21621 246320 21651 247120
rect 21831 246320 21861 247120
rect 22041 246320 22071 247120
rect 22251 246320 22281 247120
rect 22461 246320 22491 247120
rect 22671 246320 22701 247120
rect 22881 246320 22911 247120
rect 23091 246320 23121 247120
rect 23301 246320 23331 247120
rect 23511 246320 23541 247120
rect 23721 246320 23751 247120
rect 23931 246320 23961 247120
rect 24141 246320 24171 247120
rect 24351 246320 24381 247120
rect 24561 246320 24591 247120
rect 24771 246320 24801 247120
rect 24981 246320 25011 247120
rect 25191 246320 25221 247120
rect 25401 246320 25431 247120
rect 25611 246320 25641 247120
rect 25821 246320 25851 247120
rect 26031 246320 26061 247120
rect 26241 246320 26271 247120
rect 26451 246320 26481 247120
rect 26661 246320 26691 247120
rect 26871 246320 26901 247120
rect 27081 246320 27111 247120
rect 27291 246320 27321 247120
rect -3999 245284 -3969 246084
rect -3789 245284 -3759 246084
rect -3579 245284 -3549 246084
rect -3369 245284 -3339 246084
rect -3159 245284 -3129 246084
rect -2949 245284 -2919 246084
rect -2739 245284 -2709 246084
rect -2529 245284 -2499 246084
rect -2319 245284 -2289 246084
rect -2109 245284 -2079 246084
rect -1899 245284 -1869 246084
rect -1689 245284 -1659 246084
rect -1479 245284 -1449 246084
rect -1269 245284 -1239 246084
rect -1059 245284 -1029 246084
rect -849 245284 -819 246084
rect -639 245284 -609 246084
rect -429 245284 -399 246084
rect -219 245284 -189 246084
rect -9 245284 21 246084
rect 201 245284 231 246084
rect 411 245284 441 246084
rect 621 245284 651 246084
rect 831 245284 861 246084
rect 1041 245284 1071 246084
rect 1251 245284 1281 246084
rect 1461 245284 1491 246084
rect 1671 245284 1701 246084
rect 1881 245284 1911 246084
rect 2091 245284 2121 246084
rect 2301 245284 2331 246084
rect 2511 245284 2541 246084
rect 2721 245284 2751 246084
rect 2931 245284 2961 246084
rect 3141 245284 3171 246084
rect 3351 245284 3381 246084
rect 3561 245284 3591 246084
rect 3771 245284 3801 246084
rect 3981 245284 4011 246084
rect 4191 245284 4221 246084
rect 4401 245284 4431 246084
rect 4611 245284 4641 246084
rect 4821 245284 4851 246084
rect 5031 245284 5061 246084
rect 5241 245284 5271 246084
rect 5451 245284 5481 246084
rect 5661 245284 5691 246084
rect 5871 245284 5901 246084
rect 6081 245284 6111 246084
rect 6291 245284 6321 246084
rect 6501 245284 6531 246084
rect 6711 245284 6741 246084
rect 6921 245284 6951 246084
rect 7131 245284 7161 246084
rect 7341 245284 7371 246084
rect 7551 245284 7581 246084
rect 7761 245284 7791 246084
rect 7971 245284 8001 246084
rect 8181 245284 8211 246084
rect 8391 245284 8421 246084
rect 8601 245284 8631 246084
rect 8811 245284 8841 246084
rect 9021 245284 9051 246084
rect 9231 245284 9261 246084
rect 9441 245284 9471 246084
rect 9651 245284 9681 246084
rect 9861 245284 9891 246084
rect 10071 245284 10101 246084
rect 10281 245284 10311 246084
rect 10491 245284 10521 246084
rect 10701 245284 10731 246084
rect 10911 245284 10941 246084
rect 11121 245284 11151 246084
rect 11331 245284 11361 246084
rect 11541 245284 11571 246084
rect 11751 245284 11781 246084
rect 11961 245284 11991 246084
rect 12171 245284 12201 246084
rect 12381 245284 12411 246084
rect 12591 245284 12621 246084
rect 12801 245284 12831 246084
rect 13011 245284 13041 246084
rect 13221 245284 13251 246084
rect 13431 245284 13461 246084
rect 13641 245284 13671 246084
rect 13851 245284 13881 246084
rect 14061 245284 14091 246084
rect 14271 245284 14301 246084
rect 14481 245284 14511 246084
rect 14691 245284 14721 246084
rect 14901 245284 14931 246084
rect 15111 245284 15141 246084
rect 15321 245284 15351 246084
rect 15531 245284 15561 246084
rect 15741 245284 15771 246084
rect 15951 245284 15981 246084
rect 16161 245284 16191 246084
rect 16371 245284 16401 246084
rect 16581 245284 16611 246084
rect 16791 245284 16821 246084
rect 17001 245284 17031 246084
rect 17211 245284 17241 246084
rect 17421 245284 17451 246084
rect 17631 245284 17661 246084
rect 17841 245284 17871 246084
rect 18051 245284 18081 246084
rect 18261 245284 18291 246084
rect 18471 245284 18501 246084
rect 18681 245284 18711 246084
rect 18891 245284 18921 246084
rect 19101 245284 19131 246084
rect 19311 245284 19341 246084
rect 19521 245284 19551 246084
rect 19731 245284 19761 246084
rect 19941 245284 19971 246084
rect 20151 245284 20181 246084
rect 20361 245284 20391 246084
rect 20571 245284 20601 246084
rect 20781 245284 20811 246084
rect 20991 245284 21021 246084
rect 21201 245284 21231 246084
rect 21411 245284 21441 246084
rect 21621 245284 21651 246084
rect 21831 245284 21861 246084
rect 22041 245284 22071 246084
rect 22251 245284 22281 246084
rect 22461 245284 22491 246084
rect 22671 245284 22701 246084
rect 22881 245284 22911 246084
rect 23091 245284 23121 246084
rect 23301 245284 23331 246084
rect 23511 245284 23541 246084
rect 23721 245284 23751 246084
rect 23931 245284 23961 246084
rect 24141 245284 24171 246084
rect 24351 245284 24381 246084
rect 24561 245284 24591 246084
rect 24771 245284 24801 246084
rect 24981 245284 25011 246084
rect 25191 245284 25221 246084
rect 25401 245284 25431 246084
rect 25611 245284 25641 246084
rect 25821 245284 25851 246084
rect 26031 245284 26061 246084
rect 26241 245284 26271 246084
rect 26451 245284 26481 246084
rect 26661 245284 26691 246084
rect 26871 245284 26901 246084
rect 27081 245284 27111 246084
rect 27291 245284 27321 246084
rect -3999 244248 -3969 245048
rect -3789 244248 -3759 245048
rect -3579 244248 -3549 245048
rect -3369 244248 -3339 245048
rect -3159 244248 -3129 245048
rect -2949 244248 -2919 245048
rect -2739 244248 -2709 245048
rect -2529 244248 -2499 245048
rect -2319 244248 -2289 245048
rect -2109 244248 -2079 245048
rect -1899 244248 -1869 245048
rect -1689 244248 -1659 245048
rect -1479 244248 -1449 245048
rect -1269 244248 -1239 245048
rect -1059 244248 -1029 245048
rect -849 244248 -819 245048
rect -639 244248 -609 245048
rect -429 244248 -399 245048
rect -219 244248 -189 245048
rect -9 244248 21 245048
rect 201 244248 231 245048
rect 411 244248 441 245048
rect 621 244248 651 245048
rect 831 244248 861 245048
rect 1041 244248 1071 245048
rect 1251 244248 1281 245048
rect 1461 244248 1491 245048
rect 1671 244248 1701 245048
rect 1881 244248 1911 245048
rect 2091 244248 2121 245048
rect 2301 244248 2331 245048
rect 2511 244248 2541 245048
rect 2721 244248 2751 245048
rect 2931 244248 2961 245048
rect 3141 244248 3171 245048
rect 3351 244248 3381 245048
rect 3561 244248 3591 245048
rect 3771 244248 3801 245048
rect 3981 244248 4011 245048
rect 4191 244248 4221 245048
rect 4401 244248 4431 245048
rect 4611 244248 4641 245048
rect 4821 244248 4851 245048
rect 5031 244248 5061 245048
rect 5241 244248 5271 245048
rect 5451 244248 5481 245048
rect 5661 244248 5691 245048
rect 5871 244248 5901 245048
rect 6081 244248 6111 245048
rect 6291 244248 6321 245048
rect 6501 244248 6531 245048
rect 6711 244248 6741 245048
rect 6921 244248 6951 245048
rect 7131 244248 7161 245048
rect 7341 244248 7371 245048
rect 7551 244248 7581 245048
rect 7761 244248 7791 245048
rect 7971 244248 8001 245048
rect 8181 244248 8211 245048
rect 8391 244248 8421 245048
rect 8601 244248 8631 245048
rect 8811 244248 8841 245048
rect 9021 244248 9051 245048
rect 9231 244248 9261 245048
rect 9441 244248 9471 245048
rect 9651 244248 9681 245048
rect 9861 244248 9891 245048
rect 10071 244248 10101 245048
rect 10281 244248 10311 245048
rect 10491 244248 10521 245048
rect 10701 244248 10731 245048
rect 10911 244248 10941 245048
rect 11121 244248 11151 245048
rect 11331 244248 11361 245048
rect 11541 244248 11571 245048
rect 11751 244248 11781 245048
rect 11961 244248 11991 245048
rect 12171 244248 12201 245048
rect 12381 244248 12411 245048
rect 12591 244248 12621 245048
rect 12801 244248 12831 245048
rect 13011 244248 13041 245048
rect 13221 244248 13251 245048
rect 13431 244248 13461 245048
rect 13641 244248 13671 245048
rect 13851 244248 13881 245048
rect 14061 244248 14091 245048
rect 14271 244248 14301 245048
rect 14481 244248 14511 245048
rect 14691 244248 14721 245048
rect 14901 244248 14931 245048
rect 15111 244248 15141 245048
rect 15321 244248 15351 245048
rect 15531 244248 15561 245048
rect 15741 244248 15771 245048
rect 15951 244248 15981 245048
rect 16161 244248 16191 245048
rect 16371 244248 16401 245048
rect 16581 244248 16611 245048
rect 16791 244248 16821 245048
rect 17001 244248 17031 245048
rect 17211 244248 17241 245048
rect 17421 244248 17451 245048
rect 17631 244248 17661 245048
rect 17841 244248 17871 245048
rect 18051 244248 18081 245048
rect 18261 244248 18291 245048
rect 18471 244248 18501 245048
rect 18681 244248 18711 245048
rect 18891 244248 18921 245048
rect 19101 244248 19131 245048
rect 19311 244248 19341 245048
rect 19521 244248 19551 245048
rect 19731 244248 19761 245048
rect 19941 244248 19971 245048
rect 20151 244248 20181 245048
rect 20361 244248 20391 245048
rect 20571 244248 20601 245048
rect 20781 244248 20811 245048
rect 20991 244248 21021 245048
rect 21201 244248 21231 245048
rect 21411 244248 21441 245048
rect 21621 244248 21651 245048
rect 21831 244248 21861 245048
rect 22041 244248 22071 245048
rect 22251 244248 22281 245048
rect 22461 244248 22491 245048
rect 22671 244248 22701 245048
rect 22881 244248 22911 245048
rect 23091 244248 23121 245048
rect 23301 244248 23331 245048
rect 23511 244248 23541 245048
rect 23721 244248 23751 245048
rect 23931 244248 23961 245048
rect 24141 244248 24171 245048
rect 24351 244248 24381 245048
rect 24561 244248 24591 245048
rect 24771 244248 24801 245048
rect 24981 244248 25011 245048
rect 25191 244248 25221 245048
rect 25401 244248 25431 245048
rect 25611 244248 25641 245048
rect 25821 244248 25851 245048
rect 26031 244248 26061 245048
rect 26241 244248 26271 245048
rect 26451 244248 26481 245048
rect 26661 244248 26691 245048
rect 26871 244248 26901 245048
rect 27081 244248 27111 245048
rect 27291 244248 27321 245048
<< ndiff >>
rect -4061 264026 -3999 264038
rect -4061 263250 -4049 264026
rect -4015 263250 -3999 264026
rect -4061 263238 -3999 263250
rect -3969 264026 -3907 264038
rect -3969 263250 -3953 264026
rect -3919 263250 -3907 264026
rect -3969 263238 -3907 263250
rect -3851 264026 -3789 264038
rect -3851 263250 -3839 264026
rect -3805 263250 -3789 264026
rect -3851 263238 -3789 263250
rect -3759 264026 -3697 264038
rect -3759 263250 -3743 264026
rect -3709 263250 -3697 264026
rect -3759 263238 -3697 263250
rect -3641 264026 -3579 264038
rect -3641 263250 -3629 264026
rect -3595 263250 -3579 264026
rect -3641 263238 -3579 263250
rect -3549 264026 -3487 264038
rect -3549 263250 -3533 264026
rect -3499 263250 -3487 264026
rect -3549 263238 -3487 263250
rect -3431 264026 -3369 264038
rect -3431 263250 -3419 264026
rect -3385 263250 -3369 264026
rect -3431 263238 -3369 263250
rect -3339 264026 -3277 264038
rect -3339 263250 -3323 264026
rect -3289 263250 -3277 264026
rect -3339 263238 -3277 263250
rect -3221 264026 -3159 264038
rect -3221 263250 -3209 264026
rect -3175 263250 -3159 264026
rect -3221 263238 -3159 263250
rect -3129 264026 -3067 264038
rect -3129 263250 -3113 264026
rect -3079 263250 -3067 264026
rect -3129 263238 -3067 263250
rect -3011 264026 -2949 264038
rect -3011 263250 -2999 264026
rect -2965 263250 -2949 264026
rect -3011 263238 -2949 263250
rect -2919 264026 -2857 264038
rect -2919 263250 -2903 264026
rect -2869 263250 -2857 264026
rect -2919 263238 -2857 263250
rect -2801 264026 -2739 264038
rect -2801 263250 -2789 264026
rect -2755 263250 -2739 264026
rect -2801 263238 -2739 263250
rect -2709 264026 -2647 264038
rect -2709 263250 -2693 264026
rect -2659 263250 -2647 264026
rect -2709 263238 -2647 263250
rect -2591 264026 -2529 264038
rect -2591 263250 -2579 264026
rect -2545 263250 -2529 264026
rect -2591 263238 -2529 263250
rect -2499 264026 -2437 264038
rect -2499 263250 -2483 264026
rect -2449 263250 -2437 264026
rect -2499 263238 -2437 263250
rect -2381 264026 -2319 264038
rect -2381 263250 -2369 264026
rect -2335 263250 -2319 264026
rect -2381 263238 -2319 263250
rect -2289 264026 -2227 264038
rect -2289 263250 -2273 264026
rect -2239 263250 -2227 264026
rect -2289 263238 -2227 263250
rect -2171 264026 -2109 264038
rect -2171 263250 -2159 264026
rect -2125 263250 -2109 264026
rect -2171 263238 -2109 263250
rect -2079 264026 -2017 264038
rect -2079 263250 -2063 264026
rect -2029 263250 -2017 264026
rect -2079 263238 -2017 263250
rect -1961 264026 -1899 264038
rect -1961 263250 -1949 264026
rect -1915 263250 -1899 264026
rect -1961 263238 -1899 263250
rect -1869 264026 -1807 264038
rect -1869 263250 -1853 264026
rect -1819 263250 -1807 264026
rect -1869 263238 -1807 263250
rect -1751 264026 -1689 264038
rect -1751 263250 -1739 264026
rect -1705 263250 -1689 264026
rect -1751 263238 -1689 263250
rect -1659 264026 -1597 264038
rect -1659 263250 -1643 264026
rect -1609 263250 -1597 264026
rect -1659 263238 -1597 263250
rect -1541 264026 -1479 264038
rect -1541 263250 -1529 264026
rect -1495 263250 -1479 264026
rect -1541 263238 -1479 263250
rect -1449 264026 -1387 264038
rect -1449 263250 -1433 264026
rect -1399 263250 -1387 264026
rect -1449 263238 -1387 263250
rect -1331 264026 -1269 264038
rect -1331 263250 -1319 264026
rect -1285 263250 -1269 264026
rect -1331 263238 -1269 263250
rect -1239 264026 -1177 264038
rect -1239 263250 -1223 264026
rect -1189 263250 -1177 264026
rect -1239 263238 -1177 263250
rect -1121 264026 -1059 264038
rect -1121 263250 -1109 264026
rect -1075 263250 -1059 264026
rect -1121 263238 -1059 263250
rect -1029 264026 -967 264038
rect -1029 263250 -1013 264026
rect -979 263250 -967 264026
rect -1029 263238 -967 263250
rect -911 264026 -849 264038
rect -911 263250 -899 264026
rect -865 263250 -849 264026
rect -911 263238 -849 263250
rect -819 264026 -757 264038
rect -819 263250 -803 264026
rect -769 263250 -757 264026
rect -819 263238 -757 263250
rect -701 264026 -639 264038
rect -701 263250 -689 264026
rect -655 263250 -639 264026
rect -701 263238 -639 263250
rect -609 264026 -547 264038
rect -609 263250 -593 264026
rect -559 263250 -547 264026
rect -609 263238 -547 263250
rect -491 264026 -429 264038
rect -491 263250 -479 264026
rect -445 263250 -429 264026
rect -491 263238 -429 263250
rect -399 264026 -337 264038
rect -399 263250 -383 264026
rect -349 263250 -337 264026
rect -399 263238 -337 263250
rect -281 264026 -219 264038
rect -281 263250 -269 264026
rect -235 263250 -219 264026
rect -281 263238 -219 263250
rect -189 264026 -127 264038
rect -189 263250 -173 264026
rect -139 263250 -127 264026
rect -189 263238 -127 263250
rect -71 264026 -9 264038
rect -71 263250 -59 264026
rect -25 263250 -9 264026
rect -71 263238 -9 263250
rect 21 264026 83 264038
rect 21 263250 37 264026
rect 71 263250 83 264026
rect 21 263238 83 263250
rect 139 264026 201 264038
rect 139 263250 151 264026
rect 185 263250 201 264026
rect 139 263238 201 263250
rect 231 264026 293 264038
rect 231 263250 247 264026
rect 281 263250 293 264026
rect 231 263238 293 263250
rect 349 264026 411 264038
rect 349 263250 361 264026
rect 395 263250 411 264026
rect 349 263238 411 263250
rect 441 264026 503 264038
rect 441 263250 457 264026
rect 491 263250 503 264026
rect 441 263238 503 263250
rect 559 264026 621 264038
rect 559 263250 571 264026
rect 605 263250 621 264026
rect 559 263238 621 263250
rect 651 264026 713 264038
rect 651 263250 667 264026
rect 701 263250 713 264026
rect 651 263238 713 263250
rect 769 264026 831 264038
rect 769 263250 781 264026
rect 815 263250 831 264026
rect 769 263238 831 263250
rect 861 264026 923 264038
rect 861 263250 877 264026
rect 911 263250 923 264026
rect 861 263238 923 263250
rect 979 264026 1041 264038
rect 979 263250 991 264026
rect 1025 263250 1041 264026
rect 979 263238 1041 263250
rect 1071 264026 1133 264038
rect 1071 263250 1087 264026
rect 1121 263250 1133 264026
rect 1071 263238 1133 263250
rect 1189 264026 1251 264038
rect 1189 263250 1201 264026
rect 1235 263250 1251 264026
rect 1189 263238 1251 263250
rect 1281 264026 1343 264038
rect 1281 263250 1297 264026
rect 1331 263250 1343 264026
rect 1281 263238 1343 263250
rect 1399 264026 1461 264038
rect 1399 263250 1411 264026
rect 1445 263250 1461 264026
rect 1399 263238 1461 263250
rect 1491 264026 1553 264038
rect 1491 263250 1507 264026
rect 1541 263250 1553 264026
rect 1491 263238 1553 263250
rect 1609 264026 1671 264038
rect 1609 263250 1621 264026
rect 1655 263250 1671 264026
rect 1609 263238 1671 263250
rect 1701 264026 1763 264038
rect 1701 263250 1717 264026
rect 1751 263250 1763 264026
rect 1701 263238 1763 263250
rect 1819 264026 1881 264038
rect 1819 263250 1831 264026
rect 1865 263250 1881 264026
rect 1819 263238 1881 263250
rect 1911 264026 1973 264038
rect 1911 263250 1927 264026
rect 1961 263250 1973 264026
rect 1911 263238 1973 263250
rect 2029 264026 2091 264038
rect 2029 263250 2041 264026
rect 2075 263250 2091 264026
rect 2029 263238 2091 263250
rect 2121 264026 2183 264038
rect 2121 263250 2137 264026
rect 2171 263250 2183 264026
rect 2121 263238 2183 263250
rect 2239 264026 2301 264038
rect 2239 263250 2251 264026
rect 2285 263250 2301 264026
rect 2239 263238 2301 263250
rect 2331 264026 2393 264038
rect 2331 263250 2347 264026
rect 2381 263250 2393 264026
rect 2331 263238 2393 263250
rect 2449 264026 2511 264038
rect 2449 263250 2461 264026
rect 2495 263250 2511 264026
rect 2449 263238 2511 263250
rect 2541 264026 2603 264038
rect 2541 263250 2557 264026
rect 2591 263250 2603 264026
rect 2541 263238 2603 263250
rect 2659 264026 2721 264038
rect 2659 263250 2671 264026
rect 2705 263250 2721 264026
rect 2659 263238 2721 263250
rect 2751 264026 2813 264038
rect 2751 263250 2767 264026
rect 2801 263250 2813 264026
rect 2751 263238 2813 263250
rect 2869 264026 2931 264038
rect 2869 263250 2881 264026
rect 2915 263250 2931 264026
rect 2869 263238 2931 263250
rect 2961 264026 3023 264038
rect 2961 263250 2977 264026
rect 3011 263250 3023 264026
rect 2961 263238 3023 263250
rect 3079 264026 3141 264038
rect 3079 263250 3091 264026
rect 3125 263250 3141 264026
rect 3079 263238 3141 263250
rect 3171 264026 3233 264038
rect 3171 263250 3187 264026
rect 3221 263250 3233 264026
rect 3171 263238 3233 263250
rect 3289 264026 3351 264038
rect 3289 263250 3301 264026
rect 3335 263250 3351 264026
rect 3289 263238 3351 263250
rect 3381 264026 3443 264038
rect 3381 263250 3397 264026
rect 3431 263250 3443 264026
rect 3381 263238 3443 263250
rect 3499 264026 3561 264038
rect 3499 263250 3511 264026
rect 3545 263250 3561 264026
rect 3499 263238 3561 263250
rect 3591 264026 3653 264038
rect 3591 263250 3607 264026
rect 3641 263250 3653 264026
rect 3591 263238 3653 263250
rect 3709 264026 3771 264038
rect 3709 263250 3721 264026
rect 3755 263250 3771 264026
rect 3709 263238 3771 263250
rect 3801 264026 3863 264038
rect 3801 263250 3817 264026
rect 3851 263250 3863 264026
rect 3801 263238 3863 263250
rect 3919 264026 3981 264038
rect 3919 263250 3931 264026
rect 3965 263250 3981 264026
rect 3919 263238 3981 263250
rect 4011 264026 4073 264038
rect 4011 263250 4027 264026
rect 4061 263250 4073 264026
rect 4011 263238 4073 263250
rect 4129 264026 4191 264038
rect 4129 263250 4141 264026
rect 4175 263250 4191 264026
rect 4129 263238 4191 263250
rect 4221 264026 4283 264038
rect 4221 263250 4237 264026
rect 4271 263250 4283 264026
rect 4221 263238 4283 263250
rect 4339 264026 4401 264038
rect 4339 263250 4351 264026
rect 4385 263250 4401 264026
rect 4339 263238 4401 263250
rect 4431 264026 4493 264038
rect 4431 263250 4447 264026
rect 4481 263250 4493 264026
rect 4431 263238 4493 263250
rect 4549 264026 4611 264038
rect 4549 263250 4561 264026
rect 4595 263250 4611 264026
rect 4549 263238 4611 263250
rect 4641 264026 4703 264038
rect 4641 263250 4657 264026
rect 4691 263250 4703 264026
rect 4641 263238 4703 263250
rect 4759 264026 4821 264038
rect 4759 263250 4771 264026
rect 4805 263250 4821 264026
rect 4759 263238 4821 263250
rect 4851 264026 4913 264038
rect 4851 263250 4867 264026
rect 4901 263250 4913 264026
rect 4851 263238 4913 263250
rect 4969 264026 5031 264038
rect 4969 263250 4981 264026
rect 5015 263250 5031 264026
rect 4969 263238 5031 263250
rect 5061 264026 5123 264038
rect 5061 263250 5077 264026
rect 5111 263250 5123 264026
rect 5061 263238 5123 263250
rect 5179 264026 5241 264038
rect 5179 263250 5191 264026
rect 5225 263250 5241 264026
rect 5179 263238 5241 263250
rect 5271 264026 5333 264038
rect 5271 263250 5287 264026
rect 5321 263250 5333 264026
rect 5271 263238 5333 263250
rect 5389 264026 5451 264038
rect 5389 263250 5401 264026
rect 5435 263250 5451 264026
rect 5389 263238 5451 263250
rect 5481 264026 5543 264038
rect 5481 263250 5497 264026
rect 5531 263250 5543 264026
rect 5481 263238 5543 263250
rect 5599 264026 5661 264038
rect 5599 263250 5611 264026
rect 5645 263250 5661 264026
rect 5599 263238 5661 263250
rect 5691 264026 5753 264038
rect 5691 263250 5707 264026
rect 5741 263250 5753 264026
rect 5691 263238 5753 263250
rect 5809 264026 5871 264038
rect 5809 263250 5821 264026
rect 5855 263250 5871 264026
rect 5809 263238 5871 263250
rect 5901 264026 5963 264038
rect 5901 263250 5917 264026
rect 5951 263250 5963 264026
rect 5901 263238 5963 263250
rect 6019 264026 6081 264038
rect 6019 263250 6031 264026
rect 6065 263250 6081 264026
rect 6019 263238 6081 263250
rect 6111 264026 6173 264038
rect 6111 263250 6127 264026
rect 6161 263250 6173 264026
rect 6111 263238 6173 263250
rect 6229 264026 6291 264038
rect 6229 263250 6241 264026
rect 6275 263250 6291 264026
rect 6229 263238 6291 263250
rect 6321 264026 6383 264038
rect 6321 263250 6337 264026
rect 6371 263250 6383 264026
rect 6321 263238 6383 263250
rect 6439 264026 6501 264038
rect 6439 263250 6451 264026
rect 6485 263250 6501 264026
rect 6439 263238 6501 263250
rect 6531 264026 6593 264038
rect 6531 263250 6547 264026
rect 6581 263250 6593 264026
rect 6531 263238 6593 263250
rect 6649 264026 6711 264038
rect 6649 263250 6661 264026
rect 6695 263250 6711 264026
rect 6649 263238 6711 263250
rect 6741 264026 6803 264038
rect 6741 263250 6757 264026
rect 6791 263250 6803 264026
rect 6741 263238 6803 263250
rect 6859 264026 6921 264038
rect 6859 263250 6871 264026
rect 6905 263250 6921 264026
rect 6859 263238 6921 263250
rect 6951 264026 7013 264038
rect 6951 263250 6967 264026
rect 7001 263250 7013 264026
rect 6951 263238 7013 263250
rect 7069 264026 7131 264038
rect 7069 263250 7081 264026
rect 7115 263250 7131 264026
rect 7069 263238 7131 263250
rect 7161 264026 7223 264038
rect 7161 263250 7177 264026
rect 7211 263250 7223 264026
rect 7161 263238 7223 263250
rect 7279 264026 7341 264038
rect 7279 263250 7291 264026
rect 7325 263250 7341 264026
rect 7279 263238 7341 263250
rect 7371 264026 7433 264038
rect 7371 263250 7387 264026
rect 7421 263250 7433 264026
rect 7371 263238 7433 263250
rect 7489 264026 7551 264038
rect 7489 263250 7501 264026
rect 7535 263250 7551 264026
rect 7489 263238 7551 263250
rect 7581 264026 7643 264038
rect 7581 263250 7597 264026
rect 7631 263250 7643 264026
rect 7581 263238 7643 263250
rect 7699 264026 7761 264038
rect 7699 263250 7711 264026
rect 7745 263250 7761 264026
rect 7699 263238 7761 263250
rect 7791 264026 7853 264038
rect 7791 263250 7807 264026
rect 7841 263250 7853 264026
rect 7791 263238 7853 263250
rect 7909 264026 7971 264038
rect 7909 263250 7921 264026
rect 7955 263250 7971 264026
rect 7909 263238 7971 263250
rect 8001 264026 8063 264038
rect 8001 263250 8017 264026
rect 8051 263250 8063 264026
rect 8001 263238 8063 263250
rect 8119 264026 8181 264038
rect 8119 263250 8131 264026
rect 8165 263250 8181 264026
rect 8119 263238 8181 263250
rect 8211 264026 8273 264038
rect 8211 263250 8227 264026
rect 8261 263250 8273 264026
rect 8211 263238 8273 263250
rect 8329 264026 8391 264038
rect 8329 263250 8341 264026
rect 8375 263250 8391 264026
rect 8329 263238 8391 263250
rect 8421 264026 8483 264038
rect 8421 263250 8437 264026
rect 8471 263250 8483 264026
rect 8421 263238 8483 263250
rect 8539 264026 8601 264038
rect 8539 263250 8551 264026
rect 8585 263250 8601 264026
rect 8539 263238 8601 263250
rect 8631 264026 8693 264038
rect 8631 263250 8647 264026
rect 8681 263250 8693 264026
rect 8631 263238 8693 263250
rect 8749 264026 8811 264038
rect 8749 263250 8761 264026
rect 8795 263250 8811 264026
rect 8749 263238 8811 263250
rect 8841 264026 8903 264038
rect 8841 263250 8857 264026
rect 8891 263250 8903 264026
rect 8841 263238 8903 263250
rect 8959 264026 9021 264038
rect 8959 263250 8971 264026
rect 9005 263250 9021 264026
rect 8959 263238 9021 263250
rect 9051 264026 9113 264038
rect 9051 263250 9067 264026
rect 9101 263250 9113 264026
rect 9051 263238 9113 263250
rect 9169 264026 9231 264038
rect 9169 263250 9181 264026
rect 9215 263250 9231 264026
rect 9169 263238 9231 263250
rect 9261 264026 9323 264038
rect 9261 263250 9277 264026
rect 9311 263250 9323 264026
rect 9261 263238 9323 263250
rect 9379 264026 9441 264038
rect 9379 263250 9391 264026
rect 9425 263250 9441 264026
rect 9379 263238 9441 263250
rect 9471 264026 9533 264038
rect 9471 263250 9487 264026
rect 9521 263250 9533 264026
rect 9471 263238 9533 263250
rect 9589 264026 9651 264038
rect 9589 263250 9601 264026
rect 9635 263250 9651 264026
rect 9589 263238 9651 263250
rect 9681 264026 9743 264038
rect 9681 263250 9697 264026
rect 9731 263250 9743 264026
rect 9681 263238 9743 263250
rect 9799 264026 9861 264038
rect 9799 263250 9811 264026
rect 9845 263250 9861 264026
rect 9799 263238 9861 263250
rect 9891 264026 9953 264038
rect 9891 263250 9907 264026
rect 9941 263250 9953 264026
rect 9891 263238 9953 263250
rect 10009 264026 10071 264038
rect 10009 263250 10021 264026
rect 10055 263250 10071 264026
rect 10009 263238 10071 263250
rect 10101 264026 10163 264038
rect 10101 263250 10117 264026
rect 10151 263250 10163 264026
rect 10101 263238 10163 263250
rect 10219 264026 10281 264038
rect 10219 263250 10231 264026
rect 10265 263250 10281 264026
rect 10219 263238 10281 263250
rect 10311 264026 10373 264038
rect 10311 263250 10327 264026
rect 10361 263250 10373 264026
rect 10311 263238 10373 263250
rect 10429 264026 10491 264038
rect 10429 263250 10441 264026
rect 10475 263250 10491 264026
rect 10429 263238 10491 263250
rect 10521 264026 10583 264038
rect 10521 263250 10537 264026
rect 10571 263250 10583 264026
rect 10521 263238 10583 263250
rect 10639 264026 10701 264038
rect 10639 263250 10651 264026
rect 10685 263250 10701 264026
rect 10639 263238 10701 263250
rect 10731 264026 10793 264038
rect 10731 263250 10747 264026
rect 10781 263250 10793 264026
rect 10731 263238 10793 263250
rect 10849 264026 10911 264038
rect 10849 263250 10861 264026
rect 10895 263250 10911 264026
rect 10849 263238 10911 263250
rect 10941 264026 11003 264038
rect 10941 263250 10957 264026
rect 10991 263250 11003 264026
rect 10941 263238 11003 263250
rect 11059 264026 11121 264038
rect 11059 263250 11071 264026
rect 11105 263250 11121 264026
rect 11059 263238 11121 263250
rect 11151 264026 11213 264038
rect 11151 263250 11167 264026
rect 11201 263250 11213 264026
rect 11151 263238 11213 263250
rect 11269 264026 11331 264038
rect 11269 263250 11281 264026
rect 11315 263250 11331 264026
rect 11269 263238 11331 263250
rect 11361 264026 11423 264038
rect 11361 263250 11377 264026
rect 11411 263250 11423 264026
rect 11361 263238 11423 263250
rect 11479 264026 11541 264038
rect 11479 263250 11491 264026
rect 11525 263250 11541 264026
rect 11479 263238 11541 263250
rect 11571 264026 11633 264038
rect 11571 263250 11587 264026
rect 11621 263250 11633 264026
rect 11571 263238 11633 263250
rect 11689 264026 11751 264038
rect 11689 263250 11701 264026
rect 11735 263250 11751 264026
rect 11689 263238 11751 263250
rect 11781 264026 11843 264038
rect 11781 263250 11797 264026
rect 11831 263250 11843 264026
rect 11781 263238 11843 263250
rect 11899 264026 11961 264038
rect 11899 263250 11911 264026
rect 11945 263250 11961 264026
rect 11899 263238 11961 263250
rect 11991 264026 12053 264038
rect 11991 263250 12007 264026
rect 12041 263250 12053 264026
rect 11991 263238 12053 263250
rect 12109 264026 12171 264038
rect 12109 263250 12121 264026
rect 12155 263250 12171 264026
rect 12109 263238 12171 263250
rect 12201 264026 12263 264038
rect 12201 263250 12217 264026
rect 12251 263250 12263 264026
rect 12201 263238 12263 263250
rect 12319 264026 12381 264038
rect 12319 263250 12331 264026
rect 12365 263250 12381 264026
rect 12319 263238 12381 263250
rect 12411 264026 12473 264038
rect 12411 263250 12427 264026
rect 12461 263250 12473 264026
rect 12411 263238 12473 263250
rect 12529 264026 12591 264038
rect 12529 263250 12541 264026
rect 12575 263250 12591 264026
rect 12529 263238 12591 263250
rect 12621 264026 12683 264038
rect 12621 263250 12637 264026
rect 12671 263250 12683 264026
rect 12621 263238 12683 263250
rect 12739 264026 12801 264038
rect 12739 263250 12751 264026
rect 12785 263250 12801 264026
rect 12739 263238 12801 263250
rect 12831 264026 12893 264038
rect 12831 263250 12847 264026
rect 12881 263250 12893 264026
rect 12831 263238 12893 263250
rect 12949 264026 13011 264038
rect 12949 263250 12961 264026
rect 12995 263250 13011 264026
rect 12949 263238 13011 263250
rect 13041 264026 13103 264038
rect 13041 263250 13057 264026
rect 13091 263250 13103 264026
rect 13041 263238 13103 263250
rect 13159 264026 13221 264038
rect 13159 263250 13171 264026
rect 13205 263250 13221 264026
rect 13159 263238 13221 263250
rect 13251 264026 13313 264038
rect 13251 263250 13267 264026
rect 13301 263250 13313 264026
rect 13251 263238 13313 263250
rect 13369 264026 13431 264038
rect 13369 263250 13381 264026
rect 13415 263250 13431 264026
rect 13369 263238 13431 263250
rect 13461 264026 13523 264038
rect 13461 263250 13477 264026
rect 13511 263250 13523 264026
rect 13461 263238 13523 263250
rect 13579 264026 13641 264038
rect 13579 263250 13591 264026
rect 13625 263250 13641 264026
rect 13579 263238 13641 263250
rect 13671 264026 13733 264038
rect 13671 263250 13687 264026
rect 13721 263250 13733 264026
rect 13671 263238 13733 263250
rect 13789 264026 13851 264038
rect 13789 263250 13801 264026
rect 13835 263250 13851 264026
rect 13789 263238 13851 263250
rect 13881 264026 13943 264038
rect 13881 263250 13897 264026
rect 13931 263250 13943 264026
rect 13881 263238 13943 263250
rect 13999 264026 14061 264038
rect 13999 263250 14011 264026
rect 14045 263250 14061 264026
rect 13999 263238 14061 263250
rect 14091 264026 14153 264038
rect 14091 263250 14107 264026
rect 14141 263250 14153 264026
rect 14091 263238 14153 263250
rect 14209 264026 14271 264038
rect 14209 263250 14221 264026
rect 14255 263250 14271 264026
rect 14209 263238 14271 263250
rect 14301 264026 14363 264038
rect 14301 263250 14317 264026
rect 14351 263250 14363 264026
rect 14301 263238 14363 263250
rect 14419 264026 14481 264038
rect 14419 263250 14431 264026
rect 14465 263250 14481 264026
rect 14419 263238 14481 263250
rect 14511 264026 14573 264038
rect 14511 263250 14527 264026
rect 14561 263250 14573 264026
rect 14511 263238 14573 263250
rect 14629 264026 14691 264038
rect 14629 263250 14641 264026
rect 14675 263250 14691 264026
rect 14629 263238 14691 263250
rect 14721 264026 14783 264038
rect 14721 263250 14737 264026
rect 14771 263250 14783 264026
rect 14721 263238 14783 263250
rect 14839 264026 14901 264038
rect 14839 263250 14851 264026
rect 14885 263250 14901 264026
rect 14839 263238 14901 263250
rect 14931 264026 14993 264038
rect 14931 263250 14947 264026
rect 14981 263250 14993 264026
rect 14931 263238 14993 263250
rect 15049 264026 15111 264038
rect 15049 263250 15061 264026
rect 15095 263250 15111 264026
rect 15049 263238 15111 263250
rect 15141 264026 15203 264038
rect 15141 263250 15157 264026
rect 15191 263250 15203 264026
rect 15141 263238 15203 263250
rect 15259 264026 15321 264038
rect 15259 263250 15271 264026
rect 15305 263250 15321 264026
rect 15259 263238 15321 263250
rect 15351 264026 15413 264038
rect 15351 263250 15367 264026
rect 15401 263250 15413 264026
rect 15351 263238 15413 263250
rect 15469 264026 15531 264038
rect 15469 263250 15481 264026
rect 15515 263250 15531 264026
rect 15469 263238 15531 263250
rect 15561 264026 15623 264038
rect 15561 263250 15577 264026
rect 15611 263250 15623 264026
rect 15561 263238 15623 263250
rect 15679 264026 15741 264038
rect 15679 263250 15691 264026
rect 15725 263250 15741 264026
rect 15679 263238 15741 263250
rect 15771 264026 15833 264038
rect 15771 263250 15787 264026
rect 15821 263250 15833 264026
rect 15771 263238 15833 263250
rect 15889 264026 15951 264038
rect 15889 263250 15901 264026
rect 15935 263250 15951 264026
rect 15889 263238 15951 263250
rect 15981 264026 16043 264038
rect 15981 263250 15997 264026
rect 16031 263250 16043 264026
rect 15981 263238 16043 263250
rect 16099 264026 16161 264038
rect 16099 263250 16111 264026
rect 16145 263250 16161 264026
rect 16099 263238 16161 263250
rect 16191 264026 16253 264038
rect 16191 263250 16207 264026
rect 16241 263250 16253 264026
rect 16191 263238 16253 263250
rect 16309 264026 16371 264038
rect 16309 263250 16321 264026
rect 16355 263250 16371 264026
rect 16309 263238 16371 263250
rect 16401 264026 16463 264038
rect 16401 263250 16417 264026
rect 16451 263250 16463 264026
rect 16401 263238 16463 263250
rect 16519 264026 16581 264038
rect 16519 263250 16531 264026
rect 16565 263250 16581 264026
rect 16519 263238 16581 263250
rect 16611 264026 16673 264038
rect 16611 263250 16627 264026
rect 16661 263250 16673 264026
rect 16611 263238 16673 263250
rect 16729 264026 16791 264038
rect 16729 263250 16741 264026
rect 16775 263250 16791 264026
rect 16729 263238 16791 263250
rect 16821 264026 16883 264038
rect 16821 263250 16837 264026
rect 16871 263250 16883 264026
rect 16821 263238 16883 263250
rect 16939 264026 17001 264038
rect 16939 263250 16951 264026
rect 16985 263250 17001 264026
rect 16939 263238 17001 263250
rect 17031 264026 17093 264038
rect 17031 263250 17047 264026
rect 17081 263250 17093 264026
rect 17031 263238 17093 263250
rect 17149 264026 17211 264038
rect 17149 263250 17161 264026
rect 17195 263250 17211 264026
rect 17149 263238 17211 263250
rect 17241 264026 17303 264038
rect 17241 263250 17257 264026
rect 17291 263250 17303 264026
rect 17241 263238 17303 263250
rect 17359 264026 17421 264038
rect 17359 263250 17371 264026
rect 17405 263250 17421 264026
rect 17359 263238 17421 263250
rect 17451 264026 17513 264038
rect 17451 263250 17467 264026
rect 17501 263250 17513 264026
rect 17451 263238 17513 263250
rect 17569 264026 17631 264038
rect 17569 263250 17581 264026
rect 17615 263250 17631 264026
rect 17569 263238 17631 263250
rect 17661 264026 17723 264038
rect 17661 263250 17677 264026
rect 17711 263250 17723 264026
rect 17661 263238 17723 263250
rect 17779 264026 17841 264038
rect 17779 263250 17791 264026
rect 17825 263250 17841 264026
rect 17779 263238 17841 263250
rect 17871 264026 17933 264038
rect 17871 263250 17887 264026
rect 17921 263250 17933 264026
rect 17871 263238 17933 263250
rect 17989 264026 18051 264038
rect 17989 263250 18001 264026
rect 18035 263250 18051 264026
rect 17989 263238 18051 263250
rect 18081 264026 18143 264038
rect 18081 263250 18097 264026
rect 18131 263250 18143 264026
rect 18081 263238 18143 263250
rect 18199 264026 18261 264038
rect 18199 263250 18211 264026
rect 18245 263250 18261 264026
rect 18199 263238 18261 263250
rect 18291 264026 18353 264038
rect 18291 263250 18307 264026
rect 18341 263250 18353 264026
rect 18291 263238 18353 263250
rect 18409 264026 18471 264038
rect 18409 263250 18421 264026
rect 18455 263250 18471 264026
rect 18409 263238 18471 263250
rect 18501 264026 18563 264038
rect 18501 263250 18517 264026
rect 18551 263250 18563 264026
rect 18501 263238 18563 263250
rect 18619 264026 18681 264038
rect 18619 263250 18631 264026
rect 18665 263250 18681 264026
rect 18619 263238 18681 263250
rect 18711 264026 18773 264038
rect 18711 263250 18727 264026
rect 18761 263250 18773 264026
rect 18711 263238 18773 263250
rect 18829 264026 18891 264038
rect 18829 263250 18841 264026
rect 18875 263250 18891 264026
rect 18829 263238 18891 263250
rect 18921 264026 18983 264038
rect 18921 263250 18937 264026
rect 18971 263250 18983 264026
rect 18921 263238 18983 263250
rect 19039 264026 19101 264038
rect 19039 263250 19051 264026
rect 19085 263250 19101 264026
rect 19039 263238 19101 263250
rect 19131 264026 19193 264038
rect 19131 263250 19147 264026
rect 19181 263250 19193 264026
rect 19131 263238 19193 263250
rect 19249 264026 19311 264038
rect 19249 263250 19261 264026
rect 19295 263250 19311 264026
rect 19249 263238 19311 263250
rect 19341 264026 19403 264038
rect 19341 263250 19357 264026
rect 19391 263250 19403 264026
rect 19341 263238 19403 263250
rect 19459 264026 19521 264038
rect 19459 263250 19471 264026
rect 19505 263250 19521 264026
rect 19459 263238 19521 263250
rect 19551 264026 19613 264038
rect 19551 263250 19567 264026
rect 19601 263250 19613 264026
rect 19551 263238 19613 263250
rect 19669 264026 19731 264038
rect 19669 263250 19681 264026
rect 19715 263250 19731 264026
rect 19669 263238 19731 263250
rect 19761 264026 19823 264038
rect 19761 263250 19777 264026
rect 19811 263250 19823 264026
rect 19761 263238 19823 263250
rect 19879 264026 19941 264038
rect 19879 263250 19891 264026
rect 19925 263250 19941 264026
rect 19879 263238 19941 263250
rect 19971 264026 20033 264038
rect 19971 263250 19987 264026
rect 20021 263250 20033 264026
rect 19971 263238 20033 263250
rect 20089 264026 20151 264038
rect 20089 263250 20101 264026
rect 20135 263250 20151 264026
rect 20089 263238 20151 263250
rect 20181 264026 20243 264038
rect 20181 263250 20197 264026
rect 20231 263250 20243 264026
rect 20181 263238 20243 263250
rect 20299 264026 20361 264038
rect 20299 263250 20311 264026
rect 20345 263250 20361 264026
rect 20299 263238 20361 263250
rect 20391 264026 20453 264038
rect 20391 263250 20407 264026
rect 20441 263250 20453 264026
rect 20391 263238 20453 263250
rect 20509 264026 20571 264038
rect 20509 263250 20521 264026
rect 20555 263250 20571 264026
rect 20509 263238 20571 263250
rect 20601 264026 20663 264038
rect 20601 263250 20617 264026
rect 20651 263250 20663 264026
rect 20601 263238 20663 263250
rect 20719 264026 20781 264038
rect 20719 263250 20731 264026
rect 20765 263250 20781 264026
rect 20719 263238 20781 263250
rect 20811 264026 20873 264038
rect 20811 263250 20827 264026
rect 20861 263250 20873 264026
rect 20811 263238 20873 263250
rect 20929 264026 20991 264038
rect 20929 263250 20941 264026
rect 20975 263250 20991 264026
rect 20929 263238 20991 263250
rect 21021 264026 21083 264038
rect 21021 263250 21037 264026
rect 21071 263250 21083 264026
rect 21021 263238 21083 263250
rect 21139 264026 21201 264038
rect 21139 263250 21151 264026
rect 21185 263250 21201 264026
rect 21139 263238 21201 263250
rect 21231 264026 21293 264038
rect 21231 263250 21247 264026
rect 21281 263250 21293 264026
rect 21231 263238 21293 263250
rect 21349 264026 21411 264038
rect 21349 263250 21361 264026
rect 21395 263250 21411 264026
rect 21349 263238 21411 263250
rect 21441 264026 21503 264038
rect 21441 263250 21457 264026
rect 21491 263250 21503 264026
rect 21441 263238 21503 263250
rect 21559 264026 21621 264038
rect 21559 263250 21571 264026
rect 21605 263250 21621 264026
rect 21559 263238 21621 263250
rect 21651 264026 21713 264038
rect 21651 263250 21667 264026
rect 21701 263250 21713 264026
rect 21651 263238 21713 263250
rect 21769 264026 21831 264038
rect 21769 263250 21781 264026
rect 21815 263250 21831 264026
rect 21769 263238 21831 263250
rect 21861 264026 21923 264038
rect 21861 263250 21877 264026
rect 21911 263250 21923 264026
rect 21861 263238 21923 263250
rect 21979 264026 22041 264038
rect 21979 263250 21991 264026
rect 22025 263250 22041 264026
rect 21979 263238 22041 263250
rect 22071 264026 22133 264038
rect 22071 263250 22087 264026
rect 22121 263250 22133 264026
rect 22071 263238 22133 263250
rect 22189 264026 22251 264038
rect 22189 263250 22201 264026
rect 22235 263250 22251 264026
rect 22189 263238 22251 263250
rect 22281 264026 22343 264038
rect 22281 263250 22297 264026
rect 22331 263250 22343 264026
rect 22281 263238 22343 263250
rect 22399 264026 22461 264038
rect 22399 263250 22411 264026
rect 22445 263250 22461 264026
rect 22399 263238 22461 263250
rect 22491 264026 22553 264038
rect 22491 263250 22507 264026
rect 22541 263250 22553 264026
rect 22491 263238 22553 263250
rect 22609 264026 22671 264038
rect 22609 263250 22621 264026
rect 22655 263250 22671 264026
rect 22609 263238 22671 263250
rect 22701 264026 22763 264038
rect 22701 263250 22717 264026
rect 22751 263250 22763 264026
rect 22701 263238 22763 263250
rect 22819 264026 22881 264038
rect 22819 263250 22831 264026
rect 22865 263250 22881 264026
rect 22819 263238 22881 263250
rect 22911 264026 22973 264038
rect 22911 263250 22927 264026
rect 22961 263250 22973 264026
rect 22911 263238 22973 263250
rect 23029 264026 23091 264038
rect 23029 263250 23041 264026
rect 23075 263250 23091 264026
rect 23029 263238 23091 263250
rect 23121 264026 23183 264038
rect 23121 263250 23137 264026
rect 23171 263250 23183 264026
rect 23121 263238 23183 263250
rect 23239 264026 23301 264038
rect 23239 263250 23251 264026
rect 23285 263250 23301 264026
rect 23239 263238 23301 263250
rect 23331 264026 23393 264038
rect 23331 263250 23347 264026
rect 23381 263250 23393 264026
rect 23331 263238 23393 263250
rect 23449 264026 23511 264038
rect 23449 263250 23461 264026
rect 23495 263250 23511 264026
rect 23449 263238 23511 263250
rect 23541 264026 23603 264038
rect 23541 263250 23557 264026
rect 23591 263250 23603 264026
rect 23541 263238 23603 263250
rect 23659 264026 23721 264038
rect 23659 263250 23671 264026
rect 23705 263250 23721 264026
rect 23659 263238 23721 263250
rect 23751 264026 23813 264038
rect 23751 263250 23767 264026
rect 23801 263250 23813 264026
rect 23751 263238 23813 263250
rect 23869 264026 23931 264038
rect 23869 263250 23881 264026
rect 23915 263250 23931 264026
rect 23869 263238 23931 263250
rect 23961 264026 24023 264038
rect 23961 263250 23977 264026
rect 24011 263250 24023 264026
rect 23961 263238 24023 263250
rect 24079 264026 24141 264038
rect 24079 263250 24091 264026
rect 24125 263250 24141 264026
rect 24079 263238 24141 263250
rect 24171 264026 24233 264038
rect 24171 263250 24187 264026
rect 24221 263250 24233 264026
rect 24171 263238 24233 263250
rect 24289 264026 24351 264038
rect 24289 263250 24301 264026
rect 24335 263250 24351 264026
rect 24289 263238 24351 263250
rect 24381 264026 24443 264038
rect 24381 263250 24397 264026
rect 24431 263250 24443 264026
rect 24381 263238 24443 263250
rect 24499 264026 24561 264038
rect 24499 263250 24511 264026
rect 24545 263250 24561 264026
rect 24499 263238 24561 263250
rect 24591 264026 24653 264038
rect 24591 263250 24607 264026
rect 24641 263250 24653 264026
rect 24591 263238 24653 263250
rect 24709 264026 24771 264038
rect 24709 263250 24721 264026
rect 24755 263250 24771 264026
rect 24709 263238 24771 263250
rect 24801 264026 24863 264038
rect 24801 263250 24817 264026
rect 24851 263250 24863 264026
rect 24801 263238 24863 263250
rect 24919 264026 24981 264038
rect 24919 263250 24931 264026
rect 24965 263250 24981 264026
rect 24919 263238 24981 263250
rect 25011 264026 25073 264038
rect 25011 263250 25027 264026
rect 25061 263250 25073 264026
rect 25011 263238 25073 263250
rect 25129 264026 25191 264038
rect 25129 263250 25141 264026
rect 25175 263250 25191 264026
rect 25129 263238 25191 263250
rect 25221 264026 25283 264038
rect 25221 263250 25237 264026
rect 25271 263250 25283 264026
rect 25221 263238 25283 263250
rect 25339 264026 25401 264038
rect 25339 263250 25351 264026
rect 25385 263250 25401 264026
rect 25339 263238 25401 263250
rect 25431 264026 25493 264038
rect 25431 263250 25447 264026
rect 25481 263250 25493 264026
rect 25431 263238 25493 263250
rect 25549 264026 25611 264038
rect 25549 263250 25561 264026
rect 25595 263250 25611 264026
rect 25549 263238 25611 263250
rect 25641 264026 25703 264038
rect 25641 263250 25657 264026
rect 25691 263250 25703 264026
rect 25641 263238 25703 263250
rect 25759 264026 25821 264038
rect 25759 263250 25771 264026
rect 25805 263250 25821 264026
rect 25759 263238 25821 263250
rect 25851 264026 25913 264038
rect 25851 263250 25867 264026
rect 25901 263250 25913 264026
rect 25851 263238 25913 263250
rect 25969 264026 26031 264038
rect 25969 263250 25981 264026
rect 26015 263250 26031 264026
rect 25969 263238 26031 263250
rect 26061 264026 26123 264038
rect 26061 263250 26077 264026
rect 26111 263250 26123 264026
rect 26061 263238 26123 263250
rect 26179 264026 26241 264038
rect 26179 263250 26191 264026
rect 26225 263250 26241 264026
rect 26179 263238 26241 263250
rect 26271 264026 26333 264038
rect 26271 263250 26287 264026
rect 26321 263250 26333 264026
rect 26271 263238 26333 263250
rect 26389 264026 26451 264038
rect 26389 263250 26401 264026
rect 26435 263250 26451 264026
rect 26389 263238 26451 263250
rect 26481 264026 26543 264038
rect 26481 263250 26497 264026
rect 26531 263250 26543 264026
rect 26481 263238 26543 263250
rect 26599 264026 26661 264038
rect 26599 263250 26611 264026
rect 26645 263250 26661 264026
rect 26599 263238 26661 263250
rect 26691 264026 26753 264038
rect 26691 263250 26707 264026
rect 26741 263250 26753 264026
rect 26691 263238 26753 263250
rect 26809 264026 26871 264038
rect 26809 263250 26821 264026
rect 26855 263250 26871 264026
rect 26809 263238 26871 263250
rect 26901 264026 26963 264038
rect 26901 263250 26917 264026
rect 26951 263250 26963 264026
rect 26901 263238 26963 263250
rect 27019 264026 27081 264038
rect 27019 263250 27031 264026
rect 27065 263250 27081 264026
rect 27019 263238 27081 263250
rect 27111 264026 27173 264038
rect 27111 263250 27127 264026
rect 27161 263250 27173 264026
rect 27111 263238 27173 263250
rect 27229 264026 27291 264038
rect 27229 263250 27241 264026
rect 27275 263250 27291 264026
rect 27229 263238 27291 263250
rect 27321 264026 27383 264038
rect 27321 263250 27337 264026
rect 27371 263250 27383 264026
rect 27321 263238 27383 263250
rect -4061 263004 -3999 263016
rect -4061 262228 -4049 263004
rect -4015 262228 -3999 263004
rect -4061 262216 -3999 262228
rect -3969 263004 -3907 263016
rect -3969 262228 -3953 263004
rect -3919 262228 -3907 263004
rect -3969 262216 -3907 262228
rect -3851 263004 -3789 263016
rect -3851 262228 -3839 263004
rect -3805 262228 -3789 263004
rect -3851 262216 -3789 262228
rect -3759 263004 -3697 263016
rect -3759 262228 -3743 263004
rect -3709 262228 -3697 263004
rect -3759 262216 -3697 262228
rect -3641 263004 -3579 263016
rect -3641 262228 -3629 263004
rect -3595 262228 -3579 263004
rect -3641 262216 -3579 262228
rect -3549 263004 -3487 263016
rect -3549 262228 -3533 263004
rect -3499 262228 -3487 263004
rect -3549 262216 -3487 262228
rect -3431 263004 -3369 263016
rect -3431 262228 -3419 263004
rect -3385 262228 -3369 263004
rect -3431 262216 -3369 262228
rect -3339 263004 -3277 263016
rect -3339 262228 -3323 263004
rect -3289 262228 -3277 263004
rect -3339 262216 -3277 262228
rect -3221 263004 -3159 263016
rect -3221 262228 -3209 263004
rect -3175 262228 -3159 263004
rect -3221 262216 -3159 262228
rect -3129 263004 -3067 263016
rect -3129 262228 -3113 263004
rect -3079 262228 -3067 263004
rect -3129 262216 -3067 262228
rect -3011 263004 -2949 263016
rect -3011 262228 -2999 263004
rect -2965 262228 -2949 263004
rect -3011 262216 -2949 262228
rect -2919 263004 -2857 263016
rect -2919 262228 -2903 263004
rect -2869 262228 -2857 263004
rect -2919 262216 -2857 262228
rect -2801 263004 -2739 263016
rect -2801 262228 -2789 263004
rect -2755 262228 -2739 263004
rect -2801 262216 -2739 262228
rect -2709 263004 -2647 263016
rect -2709 262228 -2693 263004
rect -2659 262228 -2647 263004
rect -2709 262216 -2647 262228
rect -2591 263004 -2529 263016
rect -2591 262228 -2579 263004
rect -2545 262228 -2529 263004
rect -2591 262216 -2529 262228
rect -2499 263004 -2437 263016
rect -2499 262228 -2483 263004
rect -2449 262228 -2437 263004
rect -2499 262216 -2437 262228
rect -2381 263004 -2319 263016
rect -2381 262228 -2369 263004
rect -2335 262228 -2319 263004
rect -2381 262216 -2319 262228
rect -2289 263004 -2227 263016
rect -2289 262228 -2273 263004
rect -2239 262228 -2227 263004
rect -2289 262216 -2227 262228
rect -2171 263004 -2109 263016
rect -2171 262228 -2159 263004
rect -2125 262228 -2109 263004
rect -2171 262216 -2109 262228
rect -2079 263004 -2017 263016
rect -2079 262228 -2063 263004
rect -2029 262228 -2017 263004
rect -2079 262216 -2017 262228
rect -1961 263004 -1899 263016
rect -1961 262228 -1949 263004
rect -1915 262228 -1899 263004
rect -1961 262216 -1899 262228
rect -1869 263004 -1807 263016
rect -1869 262228 -1853 263004
rect -1819 262228 -1807 263004
rect -1869 262216 -1807 262228
rect -1751 263004 -1689 263016
rect -1751 262228 -1739 263004
rect -1705 262228 -1689 263004
rect -1751 262216 -1689 262228
rect -1659 263004 -1597 263016
rect -1659 262228 -1643 263004
rect -1609 262228 -1597 263004
rect -1659 262216 -1597 262228
rect -1541 263004 -1479 263016
rect -1541 262228 -1529 263004
rect -1495 262228 -1479 263004
rect -1541 262216 -1479 262228
rect -1449 263004 -1387 263016
rect -1449 262228 -1433 263004
rect -1399 262228 -1387 263004
rect -1449 262216 -1387 262228
rect -1331 263004 -1269 263016
rect -1331 262228 -1319 263004
rect -1285 262228 -1269 263004
rect -1331 262216 -1269 262228
rect -1239 263004 -1177 263016
rect -1239 262228 -1223 263004
rect -1189 262228 -1177 263004
rect -1239 262216 -1177 262228
rect -1121 263004 -1059 263016
rect -1121 262228 -1109 263004
rect -1075 262228 -1059 263004
rect -1121 262216 -1059 262228
rect -1029 263004 -967 263016
rect -1029 262228 -1013 263004
rect -979 262228 -967 263004
rect -1029 262216 -967 262228
rect -911 263004 -849 263016
rect -911 262228 -899 263004
rect -865 262228 -849 263004
rect -911 262216 -849 262228
rect -819 263004 -757 263016
rect -819 262228 -803 263004
rect -769 262228 -757 263004
rect -819 262216 -757 262228
rect -701 263004 -639 263016
rect -701 262228 -689 263004
rect -655 262228 -639 263004
rect -701 262216 -639 262228
rect -609 263004 -547 263016
rect -609 262228 -593 263004
rect -559 262228 -547 263004
rect -609 262216 -547 262228
rect -491 263004 -429 263016
rect -491 262228 -479 263004
rect -445 262228 -429 263004
rect -491 262216 -429 262228
rect -399 263004 -337 263016
rect -399 262228 -383 263004
rect -349 262228 -337 263004
rect -399 262216 -337 262228
rect -281 263004 -219 263016
rect -281 262228 -269 263004
rect -235 262228 -219 263004
rect -281 262216 -219 262228
rect -189 263004 -127 263016
rect -189 262228 -173 263004
rect -139 262228 -127 263004
rect -189 262216 -127 262228
rect -71 263004 -9 263016
rect -71 262228 -59 263004
rect -25 262228 -9 263004
rect -71 262216 -9 262228
rect 21 263004 83 263016
rect 21 262228 37 263004
rect 71 262228 83 263004
rect 21 262216 83 262228
rect 139 263004 201 263016
rect 139 262228 151 263004
rect 185 262228 201 263004
rect 139 262216 201 262228
rect 231 263004 293 263016
rect 231 262228 247 263004
rect 281 262228 293 263004
rect 231 262216 293 262228
rect 349 263004 411 263016
rect 349 262228 361 263004
rect 395 262228 411 263004
rect 349 262216 411 262228
rect 441 263004 503 263016
rect 441 262228 457 263004
rect 491 262228 503 263004
rect 441 262216 503 262228
rect 559 263004 621 263016
rect 559 262228 571 263004
rect 605 262228 621 263004
rect 559 262216 621 262228
rect 651 263004 713 263016
rect 651 262228 667 263004
rect 701 262228 713 263004
rect 651 262216 713 262228
rect 769 263004 831 263016
rect 769 262228 781 263004
rect 815 262228 831 263004
rect 769 262216 831 262228
rect 861 263004 923 263016
rect 861 262228 877 263004
rect 911 262228 923 263004
rect 861 262216 923 262228
rect 979 263004 1041 263016
rect 979 262228 991 263004
rect 1025 262228 1041 263004
rect 979 262216 1041 262228
rect 1071 263004 1133 263016
rect 1071 262228 1087 263004
rect 1121 262228 1133 263004
rect 1071 262216 1133 262228
rect 1189 263004 1251 263016
rect 1189 262228 1201 263004
rect 1235 262228 1251 263004
rect 1189 262216 1251 262228
rect 1281 263004 1343 263016
rect 1281 262228 1297 263004
rect 1331 262228 1343 263004
rect 1281 262216 1343 262228
rect 1399 263004 1461 263016
rect 1399 262228 1411 263004
rect 1445 262228 1461 263004
rect 1399 262216 1461 262228
rect 1491 263004 1553 263016
rect 1491 262228 1507 263004
rect 1541 262228 1553 263004
rect 1491 262216 1553 262228
rect 1609 263004 1671 263016
rect 1609 262228 1621 263004
rect 1655 262228 1671 263004
rect 1609 262216 1671 262228
rect 1701 263004 1763 263016
rect 1701 262228 1717 263004
rect 1751 262228 1763 263004
rect 1701 262216 1763 262228
rect 1819 263004 1881 263016
rect 1819 262228 1831 263004
rect 1865 262228 1881 263004
rect 1819 262216 1881 262228
rect 1911 263004 1973 263016
rect 1911 262228 1927 263004
rect 1961 262228 1973 263004
rect 1911 262216 1973 262228
rect 2029 263004 2091 263016
rect 2029 262228 2041 263004
rect 2075 262228 2091 263004
rect 2029 262216 2091 262228
rect 2121 263004 2183 263016
rect 2121 262228 2137 263004
rect 2171 262228 2183 263004
rect 2121 262216 2183 262228
rect 2239 263004 2301 263016
rect 2239 262228 2251 263004
rect 2285 262228 2301 263004
rect 2239 262216 2301 262228
rect 2331 263004 2393 263016
rect 2331 262228 2347 263004
rect 2381 262228 2393 263004
rect 2331 262216 2393 262228
rect 2449 263004 2511 263016
rect 2449 262228 2461 263004
rect 2495 262228 2511 263004
rect 2449 262216 2511 262228
rect 2541 263004 2603 263016
rect 2541 262228 2557 263004
rect 2591 262228 2603 263004
rect 2541 262216 2603 262228
rect 2659 263004 2721 263016
rect 2659 262228 2671 263004
rect 2705 262228 2721 263004
rect 2659 262216 2721 262228
rect 2751 263004 2813 263016
rect 2751 262228 2767 263004
rect 2801 262228 2813 263004
rect 2751 262216 2813 262228
rect 2869 263004 2931 263016
rect 2869 262228 2881 263004
rect 2915 262228 2931 263004
rect 2869 262216 2931 262228
rect 2961 263004 3023 263016
rect 2961 262228 2977 263004
rect 3011 262228 3023 263004
rect 2961 262216 3023 262228
rect 3079 263004 3141 263016
rect 3079 262228 3091 263004
rect 3125 262228 3141 263004
rect 3079 262216 3141 262228
rect 3171 263004 3233 263016
rect 3171 262228 3187 263004
rect 3221 262228 3233 263004
rect 3171 262216 3233 262228
rect 3289 263004 3351 263016
rect 3289 262228 3301 263004
rect 3335 262228 3351 263004
rect 3289 262216 3351 262228
rect 3381 263004 3443 263016
rect 3381 262228 3397 263004
rect 3431 262228 3443 263004
rect 3381 262216 3443 262228
rect 3499 263004 3561 263016
rect 3499 262228 3511 263004
rect 3545 262228 3561 263004
rect 3499 262216 3561 262228
rect 3591 263004 3653 263016
rect 3591 262228 3607 263004
rect 3641 262228 3653 263004
rect 3591 262216 3653 262228
rect 3709 263004 3771 263016
rect 3709 262228 3721 263004
rect 3755 262228 3771 263004
rect 3709 262216 3771 262228
rect 3801 263004 3863 263016
rect 3801 262228 3817 263004
rect 3851 262228 3863 263004
rect 3801 262216 3863 262228
rect 3919 263004 3981 263016
rect 3919 262228 3931 263004
rect 3965 262228 3981 263004
rect 3919 262216 3981 262228
rect 4011 263004 4073 263016
rect 4011 262228 4027 263004
rect 4061 262228 4073 263004
rect 4011 262216 4073 262228
rect 4129 263004 4191 263016
rect 4129 262228 4141 263004
rect 4175 262228 4191 263004
rect 4129 262216 4191 262228
rect 4221 263004 4283 263016
rect 4221 262228 4237 263004
rect 4271 262228 4283 263004
rect 4221 262216 4283 262228
rect 4339 263004 4401 263016
rect 4339 262228 4351 263004
rect 4385 262228 4401 263004
rect 4339 262216 4401 262228
rect 4431 263004 4493 263016
rect 4431 262228 4447 263004
rect 4481 262228 4493 263004
rect 4431 262216 4493 262228
rect 4549 263004 4611 263016
rect 4549 262228 4561 263004
rect 4595 262228 4611 263004
rect 4549 262216 4611 262228
rect 4641 263004 4703 263016
rect 4641 262228 4657 263004
rect 4691 262228 4703 263004
rect 4641 262216 4703 262228
rect 4759 263004 4821 263016
rect 4759 262228 4771 263004
rect 4805 262228 4821 263004
rect 4759 262216 4821 262228
rect 4851 263004 4913 263016
rect 4851 262228 4867 263004
rect 4901 262228 4913 263004
rect 4851 262216 4913 262228
rect 4969 263004 5031 263016
rect 4969 262228 4981 263004
rect 5015 262228 5031 263004
rect 4969 262216 5031 262228
rect 5061 263004 5123 263016
rect 5061 262228 5077 263004
rect 5111 262228 5123 263004
rect 5061 262216 5123 262228
rect 5179 263004 5241 263016
rect 5179 262228 5191 263004
rect 5225 262228 5241 263004
rect 5179 262216 5241 262228
rect 5271 263004 5333 263016
rect 5271 262228 5287 263004
rect 5321 262228 5333 263004
rect 5271 262216 5333 262228
rect 5389 263004 5451 263016
rect 5389 262228 5401 263004
rect 5435 262228 5451 263004
rect 5389 262216 5451 262228
rect 5481 263004 5543 263016
rect 5481 262228 5497 263004
rect 5531 262228 5543 263004
rect 5481 262216 5543 262228
rect 5599 263004 5661 263016
rect 5599 262228 5611 263004
rect 5645 262228 5661 263004
rect 5599 262216 5661 262228
rect 5691 263004 5753 263016
rect 5691 262228 5707 263004
rect 5741 262228 5753 263004
rect 5691 262216 5753 262228
rect 5809 263004 5871 263016
rect 5809 262228 5821 263004
rect 5855 262228 5871 263004
rect 5809 262216 5871 262228
rect 5901 263004 5963 263016
rect 5901 262228 5917 263004
rect 5951 262228 5963 263004
rect 5901 262216 5963 262228
rect 6019 263004 6081 263016
rect 6019 262228 6031 263004
rect 6065 262228 6081 263004
rect 6019 262216 6081 262228
rect 6111 263004 6173 263016
rect 6111 262228 6127 263004
rect 6161 262228 6173 263004
rect 6111 262216 6173 262228
rect 6229 263004 6291 263016
rect 6229 262228 6241 263004
rect 6275 262228 6291 263004
rect 6229 262216 6291 262228
rect 6321 263004 6383 263016
rect 6321 262228 6337 263004
rect 6371 262228 6383 263004
rect 6321 262216 6383 262228
rect 6439 263004 6501 263016
rect 6439 262228 6451 263004
rect 6485 262228 6501 263004
rect 6439 262216 6501 262228
rect 6531 263004 6593 263016
rect 6531 262228 6547 263004
rect 6581 262228 6593 263004
rect 6531 262216 6593 262228
rect 6649 263004 6711 263016
rect 6649 262228 6661 263004
rect 6695 262228 6711 263004
rect 6649 262216 6711 262228
rect 6741 263004 6803 263016
rect 6741 262228 6757 263004
rect 6791 262228 6803 263004
rect 6741 262216 6803 262228
rect 6859 263004 6921 263016
rect 6859 262228 6871 263004
rect 6905 262228 6921 263004
rect 6859 262216 6921 262228
rect 6951 263004 7013 263016
rect 6951 262228 6967 263004
rect 7001 262228 7013 263004
rect 6951 262216 7013 262228
rect 7069 263004 7131 263016
rect 7069 262228 7081 263004
rect 7115 262228 7131 263004
rect 7069 262216 7131 262228
rect 7161 263004 7223 263016
rect 7161 262228 7177 263004
rect 7211 262228 7223 263004
rect 7161 262216 7223 262228
rect 7279 263004 7341 263016
rect 7279 262228 7291 263004
rect 7325 262228 7341 263004
rect 7279 262216 7341 262228
rect 7371 263004 7433 263016
rect 7371 262228 7387 263004
rect 7421 262228 7433 263004
rect 7371 262216 7433 262228
rect 7489 263004 7551 263016
rect 7489 262228 7501 263004
rect 7535 262228 7551 263004
rect 7489 262216 7551 262228
rect 7581 263004 7643 263016
rect 7581 262228 7597 263004
rect 7631 262228 7643 263004
rect 7581 262216 7643 262228
rect 7699 263004 7761 263016
rect 7699 262228 7711 263004
rect 7745 262228 7761 263004
rect 7699 262216 7761 262228
rect 7791 263004 7853 263016
rect 7791 262228 7807 263004
rect 7841 262228 7853 263004
rect 7791 262216 7853 262228
rect 7909 263004 7971 263016
rect 7909 262228 7921 263004
rect 7955 262228 7971 263004
rect 7909 262216 7971 262228
rect 8001 263004 8063 263016
rect 8001 262228 8017 263004
rect 8051 262228 8063 263004
rect 8001 262216 8063 262228
rect 8119 263004 8181 263016
rect 8119 262228 8131 263004
rect 8165 262228 8181 263004
rect 8119 262216 8181 262228
rect 8211 263004 8273 263016
rect 8211 262228 8227 263004
rect 8261 262228 8273 263004
rect 8211 262216 8273 262228
rect 8329 263004 8391 263016
rect 8329 262228 8341 263004
rect 8375 262228 8391 263004
rect 8329 262216 8391 262228
rect 8421 263004 8483 263016
rect 8421 262228 8437 263004
rect 8471 262228 8483 263004
rect 8421 262216 8483 262228
rect 8539 263004 8601 263016
rect 8539 262228 8551 263004
rect 8585 262228 8601 263004
rect 8539 262216 8601 262228
rect 8631 263004 8693 263016
rect 8631 262228 8647 263004
rect 8681 262228 8693 263004
rect 8631 262216 8693 262228
rect 8749 263004 8811 263016
rect 8749 262228 8761 263004
rect 8795 262228 8811 263004
rect 8749 262216 8811 262228
rect 8841 263004 8903 263016
rect 8841 262228 8857 263004
rect 8891 262228 8903 263004
rect 8841 262216 8903 262228
rect 8959 263004 9021 263016
rect 8959 262228 8971 263004
rect 9005 262228 9021 263004
rect 8959 262216 9021 262228
rect 9051 263004 9113 263016
rect 9051 262228 9067 263004
rect 9101 262228 9113 263004
rect 9051 262216 9113 262228
rect 9169 263004 9231 263016
rect 9169 262228 9181 263004
rect 9215 262228 9231 263004
rect 9169 262216 9231 262228
rect 9261 263004 9323 263016
rect 9261 262228 9277 263004
rect 9311 262228 9323 263004
rect 9261 262216 9323 262228
rect 9379 263004 9441 263016
rect 9379 262228 9391 263004
rect 9425 262228 9441 263004
rect 9379 262216 9441 262228
rect 9471 263004 9533 263016
rect 9471 262228 9487 263004
rect 9521 262228 9533 263004
rect 9471 262216 9533 262228
rect 9589 263004 9651 263016
rect 9589 262228 9601 263004
rect 9635 262228 9651 263004
rect 9589 262216 9651 262228
rect 9681 263004 9743 263016
rect 9681 262228 9697 263004
rect 9731 262228 9743 263004
rect 9681 262216 9743 262228
rect 9799 263004 9861 263016
rect 9799 262228 9811 263004
rect 9845 262228 9861 263004
rect 9799 262216 9861 262228
rect 9891 263004 9953 263016
rect 9891 262228 9907 263004
rect 9941 262228 9953 263004
rect 9891 262216 9953 262228
rect 10009 263004 10071 263016
rect 10009 262228 10021 263004
rect 10055 262228 10071 263004
rect 10009 262216 10071 262228
rect 10101 263004 10163 263016
rect 10101 262228 10117 263004
rect 10151 262228 10163 263004
rect 10101 262216 10163 262228
rect 10219 263004 10281 263016
rect 10219 262228 10231 263004
rect 10265 262228 10281 263004
rect 10219 262216 10281 262228
rect 10311 263004 10373 263016
rect 10311 262228 10327 263004
rect 10361 262228 10373 263004
rect 10311 262216 10373 262228
rect 10429 263004 10491 263016
rect 10429 262228 10441 263004
rect 10475 262228 10491 263004
rect 10429 262216 10491 262228
rect 10521 263004 10583 263016
rect 10521 262228 10537 263004
rect 10571 262228 10583 263004
rect 10521 262216 10583 262228
rect 10639 263004 10701 263016
rect 10639 262228 10651 263004
rect 10685 262228 10701 263004
rect 10639 262216 10701 262228
rect 10731 263004 10793 263016
rect 10731 262228 10747 263004
rect 10781 262228 10793 263004
rect 10731 262216 10793 262228
rect 10849 263004 10911 263016
rect 10849 262228 10861 263004
rect 10895 262228 10911 263004
rect 10849 262216 10911 262228
rect 10941 263004 11003 263016
rect 10941 262228 10957 263004
rect 10991 262228 11003 263004
rect 10941 262216 11003 262228
rect 11059 263004 11121 263016
rect 11059 262228 11071 263004
rect 11105 262228 11121 263004
rect 11059 262216 11121 262228
rect 11151 263004 11213 263016
rect 11151 262228 11167 263004
rect 11201 262228 11213 263004
rect 11151 262216 11213 262228
rect 11269 263004 11331 263016
rect 11269 262228 11281 263004
rect 11315 262228 11331 263004
rect 11269 262216 11331 262228
rect 11361 263004 11423 263016
rect 11361 262228 11377 263004
rect 11411 262228 11423 263004
rect 11361 262216 11423 262228
rect 11479 263004 11541 263016
rect 11479 262228 11491 263004
rect 11525 262228 11541 263004
rect 11479 262216 11541 262228
rect 11571 263004 11633 263016
rect 11571 262228 11587 263004
rect 11621 262228 11633 263004
rect 11571 262216 11633 262228
rect 11689 263004 11751 263016
rect 11689 262228 11701 263004
rect 11735 262228 11751 263004
rect 11689 262216 11751 262228
rect 11781 263004 11843 263016
rect 11781 262228 11797 263004
rect 11831 262228 11843 263004
rect 11781 262216 11843 262228
rect 11899 263004 11961 263016
rect 11899 262228 11911 263004
rect 11945 262228 11961 263004
rect 11899 262216 11961 262228
rect 11991 263004 12053 263016
rect 11991 262228 12007 263004
rect 12041 262228 12053 263004
rect 11991 262216 12053 262228
rect 12109 263004 12171 263016
rect 12109 262228 12121 263004
rect 12155 262228 12171 263004
rect 12109 262216 12171 262228
rect 12201 263004 12263 263016
rect 12201 262228 12217 263004
rect 12251 262228 12263 263004
rect 12201 262216 12263 262228
rect 12319 263004 12381 263016
rect 12319 262228 12331 263004
rect 12365 262228 12381 263004
rect 12319 262216 12381 262228
rect 12411 263004 12473 263016
rect 12411 262228 12427 263004
rect 12461 262228 12473 263004
rect 12411 262216 12473 262228
rect 12529 263004 12591 263016
rect 12529 262228 12541 263004
rect 12575 262228 12591 263004
rect 12529 262216 12591 262228
rect 12621 263004 12683 263016
rect 12621 262228 12637 263004
rect 12671 262228 12683 263004
rect 12621 262216 12683 262228
rect 12739 263004 12801 263016
rect 12739 262228 12751 263004
rect 12785 262228 12801 263004
rect 12739 262216 12801 262228
rect 12831 263004 12893 263016
rect 12831 262228 12847 263004
rect 12881 262228 12893 263004
rect 12831 262216 12893 262228
rect 12949 263004 13011 263016
rect 12949 262228 12961 263004
rect 12995 262228 13011 263004
rect 12949 262216 13011 262228
rect 13041 263004 13103 263016
rect 13041 262228 13057 263004
rect 13091 262228 13103 263004
rect 13041 262216 13103 262228
rect 13159 263004 13221 263016
rect 13159 262228 13171 263004
rect 13205 262228 13221 263004
rect 13159 262216 13221 262228
rect 13251 263004 13313 263016
rect 13251 262228 13267 263004
rect 13301 262228 13313 263004
rect 13251 262216 13313 262228
rect 13369 263004 13431 263016
rect 13369 262228 13381 263004
rect 13415 262228 13431 263004
rect 13369 262216 13431 262228
rect 13461 263004 13523 263016
rect 13461 262228 13477 263004
rect 13511 262228 13523 263004
rect 13461 262216 13523 262228
rect 13579 263004 13641 263016
rect 13579 262228 13591 263004
rect 13625 262228 13641 263004
rect 13579 262216 13641 262228
rect 13671 263004 13733 263016
rect 13671 262228 13687 263004
rect 13721 262228 13733 263004
rect 13671 262216 13733 262228
rect 13789 263004 13851 263016
rect 13789 262228 13801 263004
rect 13835 262228 13851 263004
rect 13789 262216 13851 262228
rect 13881 263004 13943 263016
rect 13881 262228 13897 263004
rect 13931 262228 13943 263004
rect 13881 262216 13943 262228
rect 13999 263004 14061 263016
rect 13999 262228 14011 263004
rect 14045 262228 14061 263004
rect 13999 262216 14061 262228
rect 14091 263004 14153 263016
rect 14091 262228 14107 263004
rect 14141 262228 14153 263004
rect 14091 262216 14153 262228
rect 14209 263004 14271 263016
rect 14209 262228 14221 263004
rect 14255 262228 14271 263004
rect 14209 262216 14271 262228
rect 14301 263004 14363 263016
rect 14301 262228 14317 263004
rect 14351 262228 14363 263004
rect 14301 262216 14363 262228
rect 14419 263004 14481 263016
rect 14419 262228 14431 263004
rect 14465 262228 14481 263004
rect 14419 262216 14481 262228
rect 14511 263004 14573 263016
rect 14511 262228 14527 263004
rect 14561 262228 14573 263004
rect 14511 262216 14573 262228
rect 14629 263004 14691 263016
rect 14629 262228 14641 263004
rect 14675 262228 14691 263004
rect 14629 262216 14691 262228
rect 14721 263004 14783 263016
rect 14721 262228 14737 263004
rect 14771 262228 14783 263004
rect 14721 262216 14783 262228
rect 14839 263004 14901 263016
rect 14839 262228 14851 263004
rect 14885 262228 14901 263004
rect 14839 262216 14901 262228
rect 14931 263004 14993 263016
rect 14931 262228 14947 263004
rect 14981 262228 14993 263004
rect 14931 262216 14993 262228
rect 15049 263004 15111 263016
rect 15049 262228 15061 263004
rect 15095 262228 15111 263004
rect 15049 262216 15111 262228
rect 15141 263004 15203 263016
rect 15141 262228 15157 263004
rect 15191 262228 15203 263004
rect 15141 262216 15203 262228
rect 15259 263004 15321 263016
rect 15259 262228 15271 263004
rect 15305 262228 15321 263004
rect 15259 262216 15321 262228
rect 15351 263004 15413 263016
rect 15351 262228 15367 263004
rect 15401 262228 15413 263004
rect 15351 262216 15413 262228
rect 15469 263004 15531 263016
rect 15469 262228 15481 263004
rect 15515 262228 15531 263004
rect 15469 262216 15531 262228
rect 15561 263004 15623 263016
rect 15561 262228 15577 263004
rect 15611 262228 15623 263004
rect 15561 262216 15623 262228
rect 15679 263004 15741 263016
rect 15679 262228 15691 263004
rect 15725 262228 15741 263004
rect 15679 262216 15741 262228
rect 15771 263004 15833 263016
rect 15771 262228 15787 263004
rect 15821 262228 15833 263004
rect 15771 262216 15833 262228
rect 15889 263004 15951 263016
rect 15889 262228 15901 263004
rect 15935 262228 15951 263004
rect 15889 262216 15951 262228
rect 15981 263004 16043 263016
rect 15981 262228 15997 263004
rect 16031 262228 16043 263004
rect 15981 262216 16043 262228
rect 16099 263004 16161 263016
rect 16099 262228 16111 263004
rect 16145 262228 16161 263004
rect 16099 262216 16161 262228
rect 16191 263004 16253 263016
rect 16191 262228 16207 263004
rect 16241 262228 16253 263004
rect 16191 262216 16253 262228
rect 16309 263004 16371 263016
rect 16309 262228 16321 263004
rect 16355 262228 16371 263004
rect 16309 262216 16371 262228
rect 16401 263004 16463 263016
rect 16401 262228 16417 263004
rect 16451 262228 16463 263004
rect 16401 262216 16463 262228
rect 16519 263004 16581 263016
rect 16519 262228 16531 263004
rect 16565 262228 16581 263004
rect 16519 262216 16581 262228
rect 16611 263004 16673 263016
rect 16611 262228 16627 263004
rect 16661 262228 16673 263004
rect 16611 262216 16673 262228
rect 16729 263004 16791 263016
rect 16729 262228 16741 263004
rect 16775 262228 16791 263004
rect 16729 262216 16791 262228
rect 16821 263004 16883 263016
rect 16821 262228 16837 263004
rect 16871 262228 16883 263004
rect 16821 262216 16883 262228
rect 16939 263004 17001 263016
rect 16939 262228 16951 263004
rect 16985 262228 17001 263004
rect 16939 262216 17001 262228
rect 17031 263004 17093 263016
rect 17031 262228 17047 263004
rect 17081 262228 17093 263004
rect 17031 262216 17093 262228
rect 17149 263004 17211 263016
rect 17149 262228 17161 263004
rect 17195 262228 17211 263004
rect 17149 262216 17211 262228
rect 17241 263004 17303 263016
rect 17241 262228 17257 263004
rect 17291 262228 17303 263004
rect 17241 262216 17303 262228
rect 17359 263004 17421 263016
rect 17359 262228 17371 263004
rect 17405 262228 17421 263004
rect 17359 262216 17421 262228
rect 17451 263004 17513 263016
rect 17451 262228 17467 263004
rect 17501 262228 17513 263004
rect 17451 262216 17513 262228
rect 17569 263004 17631 263016
rect 17569 262228 17581 263004
rect 17615 262228 17631 263004
rect 17569 262216 17631 262228
rect 17661 263004 17723 263016
rect 17661 262228 17677 263004
rect 17711 262228 17723 263004
rect 17661 262216 17723 262228
rect 17779 263004 17841 263016
rect 17779 262228 17791 263004
rect 17825 262228 17841 263004
rect 17779 262216 17841 262228
rect 17871 263004 17933 263016
rect 17871 262228 17887 263004
rect 17921 262228 17933 263004
rect 17871 262216 17933 262228
rect 17989 263004 18051 263016
rect 17989 262228 18001 263004
rect 18035 262228 18051 263004
rect 17989 262216 18051 262228
rect 18081 263004 18143 263016
rect 18081 262228 18097 263004
rect 18131 262228 18143 263004
rect 18081 262216 18143 262228
rect 18199 263004 18261 263016
rect 18199 262228 18211 263004
rect 18245 262228 18261 263004
rect 18199 262216 18261 262228
rect 18291 263004 18353 263016
rect 18291 262228 18307 263004
rect 18341 262228 18353 263004
rect 18291 262216 18353 262228
rect 18409 263004 18471 263016
rect 18409 262228 18421 263004
rect 18455 262228 18471 263004
rect 18409 262216 18471 262228
rect 18501 263004 18563 263016
rect 18501 262228 18517 263004
rect 18551 262228 18563 263004
rect 18501 262216 18563 262228
rect 18619 263004 18681 263016
rect 18619 262228 18631 263004
rect 18665 262228 18681 263004
rect 18619 262216 18681 262228
rect 18711 263004 18773 263016
rect 18711 262228 18727 263004
rect 18761 262228 18773 263004
rect 18711 262216 18773 262228
rect 18829 263004 18891 263016
rect 18829 262228 18841 263004
rect 18875 262228 18891 263004
rect 18829 262216 18891 262228
rect 18921 263004 18983 263016
rect 18921 262228 18937 263004
rect 18971 262228 18983 263004
rect 18921 262216 18983 262228
rect 19039 263004 19101 263016
rect 19039 262228 19051 263004
rect 19085 262228 19101 263004
rect 19039 262216 19101 262228
rect 19131 263004 19193 263016
rect 19131 262228 19147 263004
rect 19181 262228 19193 263004
rect 19131 262216 19193 262228
rect 19249 263004 19311 263016
rect 19249 262228 19261 263004
rect 19295 262228 19311 263004
rect 19249 262216 19311 262228
rect 19341 263004 19403 263016
rect 19341 262228 19357 263004
rect 19391 262228 19403 263004
rect 19341 262216 19403 262228
rect 19459 263004 19521 263016
rect 19459 262228 19471 263004
rect 19505 262228 19521 263004
rect 19459 262216 19521 262228
rect 19551 263004 19613 263016
rect 19551 262228 19567 263004
rect 19601 262228 19613 263004
rect 19551 262216 19613 262228
rect 19669 263004 19731 263016
rect 19669 262228 19681 263004
rect 19715 262228 19731 263004
rect 19669 262216 19731 262228
rect 19761 263004 19823 263016
rect 19761 262228 19777 263004
rect 19811 262228 19823 263004
rect 19761 262216 19823 262228
rect 19879 263004 19941 263016
rect 19879 262228 19891 263004
rect 19925 262228 19941 263004
rect 19879 262216 19941 262228
rect 19971 263004 20033 263016
rect 19971 262228 19987 263004
rect 20021 262228 20033 263004
rect 19971 262216 20033 262228
rect 20089 263004 20151 263016
rect 20089 262228 20101 263004
rect 20135 262228 20151 263004
rect 20089 262216 20151 262228
rect 20181 263004 20243 263016
rect 20181 262228 20197 263004
rect 20231 262228 20243 263004
rect 20181 262216 20243 262228
rect 20299 263004 20361 263016
rect 20299 262228 20311 263004
rect 20345 262228 20361 263004
rect 20299 262216 20361 262228
rect 20391 263004 20453 263016
rect 20391 262228 20407 263004
rect 20441 262228 20453 263004
rect 20391 262216 20453 262228
rect 20509 263004 20571 263016
rect 20509 262228 20521 263004
rect 20555 262228 20571 263004
rect 20509 262216 20571 262228
rect 20601 263004 20663 263016
rect 20601 262228 20617 263004
rect 20651 262228 20663 263004
rect 20601 262216 20663 262228
rect 20719 263004 20781 263016
rect 20719 262228 20731 263004
rect 20765 262228 20781 263004
rect 20719 262216 20781 262228
rect 20811 263004 20873 263016
rect 20811 262228 20827 263004
rect 20861 262228 20873 263004
rect 20811 262216 20873 262228
rect 20929 263004 20991 263016
rect 20929 262228 20941 263004
rect 20975 262228 20991 263004
rect 20929 262216 20991 262228
rect 21021 263004 21083 263016
rect 21021 262228 21037 263004
rect 21071 262228 21083 263004
rect 21021 262216 21083 262228
rect 21139 263004 21201 263016
rect 21139 262228 21151 263004
rect 21185 262228 21201 263004
rect 21139 262216 21201 262228
rect 21231 263004 21293 263016
rect 21231 262228 21247 263004
rect 21281 262228 21293 263004
rect 21231 262216 21293 262228
rect 21349 263004 21411 263016
rect 21349 262228 21361 263004
rect 21395 262228 21411 263004
rect 21349 262216 21411 262228
rect 21441 263004 21503 263016
rect 21441 262228 21457 263004
rect 21491 262228 21503 263004
rect 21441 262216 21503 262228
rect 21559 263004 21621 263016
rect 21559 262228 21571 263004
rect 21605 262228 21621 263004
rect 21559 262216 21621 262228
rect 21651 263004 21713 263016
rect 21651 262228 21667 263004
rect 21701 262228 21713 263004
rect 21651 262216 21713 262228
rect 21769 263004 21831 263016
rect 21769 262228 21781 263004
rect 21815 262228 21831 263004
rect 21769 262216 21831 262228
rect 21861 263004 21923 263016
rect 21861 262228 21877 263004
rect 21911 262228 21923 263004
rect 21861 262216 21923 262228
rect 21979 263004 22041 263016
rect 21979 262228 21991 263004
rect 22025 262228 22041 263004
rect 21979 262216 22041 262228
rect 22071 263004 22133 263016
rect 22071 262228 22087 263004
rect 22121 262228 22133 263004
rect 22071 262216 22133 262228
rect 22189 263004 22251 263016
rect 22189 262228 22201 263004
rect 22235 262228 22251 263004
rect 22189 262216 22251 262228
rect 22281 263004 22343 263016
rect 22281 262228 22297 263004
rect 22331 262228 22343 263004
rect 22281 262216 22343 262228
rect 22399 263004 22461 263016
rect 22399 262228 22411 263004
rect 22445 262228 22461 263004
rect 22399 262216 22461 262228
rect 22491 263004 22553 263016
rect 22491 262228 22507 263004
rect 22541 262228 22553 263004
rect 22491 262216 22553 262228
rect 22609 263004 22671 263016
rect 22609 262228 22621 263004
rect 22655 262228 22671 263004
rect 22609 262216 22671 262228
rect 22701 263004 22763 263016
rect 22701 262228 22717 263004
rect 22751 262228 22763 263004
rect 22701 262216 22763 262228
rect 22819 263004 22881 263016
rect 22819 262228 22831 263004
rect 22865 262228 22881 263004
rect 22819 262216 22881 262228
rect 22911 263004 22973 263016
rect 22911 262228 22927 263004
rect 22961 262228 22973 263004
rect 22911 262216 22973 262228
rect 23029 263004 23091 263016
rect 23029 262228 23041 263004
rect 23075 262228 23091 263004
rect 23029 262216 23091 262228
rect 23121 263004 23183 263016
rect 23121 262228 23137 263004
rect 23171 262228 23183 263004
rect 23121 262216 23183 262228
rect 23239 263004 23301 263016
rect 23239 262228 23251 263004
rect 23285 262228 23301 263004
rect 23239 262216 23301 262228
rect 23331 263004 23393 263016
rect 23331 262228 23347 263004
rect 23381 262228 23393 263004
rect 23331 262216 23393 262228
rect 23449 263004 23511 263016
rect 23449 262228 23461 263004
rect 23495 262228 23511 263004
rect 23449 262216 23511 262228
rect 23541 263004 23603 263016
rect 23541 262228 23557 263004
rect 23591 262228 23603 263004
rect 23541 262216 23603 262228
rect 23659 263004 23721 263016
rect 23659 262228 23671 263004
rect 23705 262228 23721 263004
rect 23659 262216 23721 262228
rect 23751 263004 23813 263016
rect 23751 262228 23767 263004
rect 23801 262228 23813 263004
rect 23751 262216 23813 262228
rect 23869 263004 23931 263016
rect 23869 262228 23881 263004
rect 23915 262228 23931 263004
rect 23869 262216 23931 262228
rect 23961 263004 24023 263016
rect 23961 262228 23977 263004
rect 24011 262228 24023 263004
rect 23961 262216 24023 262228
rect 24079 263004 24141 263016
rect 24079 262228 24091 263004
rect 24125 262228 24141 263004
rect 24079 262216 24141 262228
rect 24171 263004 24233 263016
rect 24171 262228 24187 263004
rect 24221 262228 24233 263004
rect 24171 262216 24233 262228
rect 24289 263004 24351 263016
rect 24289 262228 24301 263004
rect 24335 262228 24351 263004
rect 24289 262216 24351 262228
rect 24381 263004 24443 263016
rect 24381 262228 24397 263004
rect 24431 262228 24443 263004
rect 24381 262216 24443 262228
rect 24499 263004 24561 263016
rect 24499 262228 24511 263004
rect 24545 262228 24561 263004
rect 24499 262216 24561 262228
rect 24591 263004 24653 263016
rect 24591 262228 24607 263004
rect 24641 262228 24653 263004
rect 24591 262216 24653 262228
rect 24709 263004 24771 263016
rect 24709 262228 24721 263004
rect 24755 262228 24771 263004
rect 24709 262216 24771 262228
rect 24801 263004 24863 263016
rect 24801 262228 24817 263004
rect 24851 262228 24863 263004
rect 24801 262216 24863 262228
rect 24919 263004 24981 263016
rect 24919 262228 24931 263004
rect 24965 262228 24981 263004
rect 24919 262216 24981 262228
rect 25011 263004 25073 263016
rect 25011 262228 25027 263004
rect 25061 262228 25073 263004
rect 25011 262216 25073 262228
rect 25129 263004 25191 263016
rect 25129 262228 25141 263004
rect 25175 262228 25191 263004
rect 25129 262216 25191 262228
rect 25221 263004 25283 263016
rect 25221 262228 25237 263004
rect 25271 262228 25283 263004
rect 25221 262216 25283 262228
rect 25339 263004 25401 263016
rect 25339 262228 25351 263004
rect 25385 262228 25401 263004
rect 25339 262216 25401 262228
rect 25431 263004 25493 263016
rect 25431 262228 25447 263004
rect 25481 262228 25493 263004
rect 25431 262216 25493 262228
rect 25549 263004 25611 263016
rect 25549 262228 25561 263004
rect 25595 262228 25611 263004
rect 25549 262216 25611 262228
rect 25641 263004 25703 263016
rect 25641 262228 25657 263004
rect 25691 262228 25703 263004
rect 25641 262216 25703 262228
rect 25759 263004 25821 263016
rect 25759 262228 25771 263004
rect 25805 262228 25821 263004
rect 25759 262216 25821 262228
rect 25851 263004 25913 263016
rect 25851 262228 25867 263004
rect 25901 262228 25913 263004
rect 25851 262216 25913 262228
rect 25969 263004 26031 263016
rect 25969 262228 25981 263004
rect 26015 262228 26031 263004
rect 25969 262216 26031 262228
rect 26061 263004 26123 263016
rect 26061 262228 26077 263004
rect 26111 262228 26123 263004
rect 26061 262216 26123 262228
rect 26179 263004 26241 263016
rect 26179 262228 26191 263004
rect 26225 262228 26241 263004
rect 26179 262216 26241 262228
rect 26271 263004 26333 263016
rect 26271 262228 26287 263004
rect 26321 262228 26333 263004
rect 26271 262216 26333 262228
rect 26389 263004 26451 263016
rect 26389 262228 26401 263004
rect 26435 262228 26451 263004
rect 26389 262216 26451 262228
rect 26481 263004 26543 263016
rect 26481 262228 26497 263004
rect 26531 262228 26543 263004
rect 26481 262216 26543 262228
rect 26599 263004 26661 263016
rect 26599 262228 26611 263004
rect 26645 262228 26661 263004
rect 26599 262216 26661 262228
rect 26691 263004 26753 263016
rect 26691 262228 26707 263004
rect 26741 262228 26753 263004
rect 26691 262216 26753 262228
rect 26809 263004 26871 263016
rect 26809 262228 26821 263004
rect 26855 262228 26871 263004
rect 26809 262216 26871 262228
rect 26901 263004 26963 263016
rect 26901 262228 26917 263004
rect 26951 262228 26963 263004
rect 26901 262216 26963 262228
rect 27019 263004 27081 263016
rect 27019 262228 27031 263004
rect 27065 262228 27081 263004
rect 27019 262216 27081 262228
rect 27111 263004 27173 263016
rect 27111 262228 27127 263004
rect 27161 262228 27173 263004
rect 27111 262216 27173 262228
rect 27229 263004 27291 263016
rect 27229 262228 27241 263004
rect 27275 262228 27291 263004
rect 27229 262216 27291 262228
rect 27321 263004 27383 263016
rect 27321 262228 27337 263004
rect 27371 262228 27383 263004
rect 27321 262216 27383 262228
<< pdiff >>
rect -4061 254489 -3999 254501
rect -4061 253713 -4049 254489
rect -4015 253713 -3999 254489
rect -4061 253701 -3999 253713
rect -3969 254489 -3907 254501
rect -3969 253713 -3953 254489
rect -3919 253713 -3907 254489
rect -3969 253701 -3907 253713
rect -3851 254489 -3789 254501
rect -3851 253713 -3839 254489
rect -3805 253713 -3789 254489
rect -3851 253701 -3789 253713
rect -3759 254489 -3697 254501
rect -3759 253713 -3743 254489
rect -3709 253713 -3697 254489
rect -3759 253701 -3697 253713
rect -3641 254489 -3579 254501
rect -3641 253713 -3629 254489
rect -3595 253713 -3579 254489
rect -3641 253701 -3579 253713
rect -3549 254489 -3487 254501
rect -3549 253713 -3533 254489
rect -3499 253713 -3487 254489
rect -3549 253701 -3487 253713
rect -3431 254489 -3369 254501
rect -3431 253713 -3419 254489
rect -3385 253713 -3369 254489
rect -3431 253701 -3369 253713
rect -3339 254489 -3277 254501
rect -3339 253713 -3323 254489
rect -3289 253713 -3277 254489
rect -3339 253701 -3277 253713
rect -3221 254489 -3159 254501
rect -3221 253713 -3209 254489
rect -3175 253713 -3159 254489
rect -3221 253701 -3159 253713
rect -3129 254489 -3067 254501
rect -3129 253713 -3113 254489
rect -3079 253713 -3067 254489
rect -3129 253701 -3067 253713
rect -3011 254489 -2949 254501
rect -3011 253713 -2999 254489
rect -2965 253713 -2949 254489
rect -3011 253701 -2949 253713
rect -2919 254489 -2857 254501
rect -2919 253713 -2903 254489
rect -2869 253713 -2857 254489
rect -2919 253701 -2857 253713
rect -2801 254489 -2739 254501
rect -2801 253713 -2789 254489
rect -2755 253713 -2739 254489
rect -2801 253701 -2739 253713
rect -2709 254489 -2647 254501
rect -2709 253713 -2693 254489
rect -2659 253713 -2647 254489
rect -2709 253701 -2647 253713
rect -2591 254489 -2529 254501
rect -2591 253713 -2579 254489
rect -2545 253713 -2529 254489
rect -2591 253701 -2529 253713
rect -2499 254489 -2437 254501
rect -2499 253713 -2483 254489
rect -2449 253713 -2437 254489
rect -2499 253701 -2437 253713
rect -2381 254489 -2319 254501
rect -2381 253713 -2369 254489
rect -2335 253713 -2319 254489
rect -2381 253701 -2319 253713
rect -2289 254489 -2227 254501
rect -2289 253713 -2273 254489
rect -2239 253713 -2227 254489
rect -2289 253701 -2227 253713
rect -2171 254489 -2109 254501
rect -2171 253713 -2159 254489
rect -2125 253713 -2109 254489
rect -2171 253701 -2109 253713
rect -2079 254489 -2017 254501
rect -2079 253713 -2063 254489
rect -2029 253713 -2017 254489
rect -2079 253701 -2017 253713
rect -1961 254489 -1899 254501
rect -1961 253713 -1949 254489
rect -1915 253713 -1899 254489
rect -1961 253701 -1899 253713
rect -1869 254489 -1807 254501
rect -1869 253713 -1853 254489
rect -1819 253713 -1807 254489
rect -1869 253701 -1807 253713
rect -1751 254489 -1689 254501
rect -1751 253713 -1739 254489
rect -1705 253713 -1689 254489
rect -1751 253701 -1689 253713
rect -1659 254489 -1597 254501
rect -1659 253713 -1643 254489
rect -1609 253713 -1597 254489
rect -1659 253701 -1597 253713
rect -1541 254489 -1479 254501
rect -1541 253713 -1529 254489
rect -1495 253713 -1479 254489
rect -1541 253701 -1479 253713
rect -1449 254489 -1387 254501
rect -1449 253713 -1433 254489
rect -1399 253713 -1387 254489
rect -1449 253701 -1387 253713
rect -1331 254489 -1269 254501
rect -1331 253713 -1319 254489
rect -1285 253713 -1269 254489
rect -1331 253701 -1269 253713
rect -1239 254489 -1177 254501
rect -1239 253713 -1223 254489
rect -1189 253713 -1177 254489
rect -1239 253701 -1177 253713
rect -1121 254489 -1059 254501
rect -1121 253713 -1109 254489
rect -1075 253713 -1059 254489
rect -1121 253701 -1059 253713
rect -1029 254489 -967 254501
rect -1029 253713 -1013 254489
rect -979 253713 -967 254489
rect -1029 253701 -967 253713
rect -911 254489 -849 254501
rect -911 253713 -899 254489
rect -865 253713 -849 254489
rect -911 253701 -849 253713
rect -819 254489 -757 254501
rect -819 253713 -803 254489
rect -769 253713 -757 254489
rect -819 253701 -757 253713
rect -701 254489 -639 254501
rect -701 253713 -689 254489
rect -655 253713 -639 254489
rect -701 253701 -639 253713
rect -609 254489 -547 254501
rect -609 253713 -593 254489
rect -559 253713 -547 254489
rect -609 253701 -547 253713
rect -491 254489 -429 254501
rect -491 253713 -479 254489
rect -445 253713 -429 254489
rect -491 253701 -429 253713
rect -399 254489 -337 254501
rect -399 253713 -383 254489
rect -349 253713 -337 254489
rect -399 253701 -337 253713
rect -281 254489 -219 254501
rect -281 253713 -269 254489
rect -235 253713 -219 254489
rect -281 253701 -219 253713
rect -189 254489 -127 254501
rect -189 253713 -173 254489
rect -139 253713 -127 254489
rect -189 253701 -127 253713
rect -71 254489 -9 254501
rect -71 253713 -59 254489
rect -25 253713 -9 254489
rect -71 253701 -9 253713
rect 21 254489 83 254501
rect 21 253713 37 254489
rect 71 253713 83 254489
rect 21 253701 83 253713
rect 139 254489 201 254501
rect 139 253713 151 254489
rect 185 253713 201 254489
rect 139 253701 201 253713
rect 231 254489 293 254501
rect 231 253713 247 254489
rect 281 253713 293 254489
rect 231 253701 293 253713
rect 349 254489 411 254501
rect 349 253713 361 254489
rect 395 253713 411 254489
rect 349 253701 411 253713
rect 441 254489 503 254501
rect 441 253713 457 254489
rect 491 253713 503 254489
rect 441 253701 503 253713
rect 559 254489 621 254501
rect 559 253713 571 254489
rect 605 253713 621 254489
rect 559 253701 621 253713
rect 651 254489 713 254501
rect 651 253713 667 254489
rect 701 253713 713 254489
rect 651 253701 713 253713
rect 769 254489 831 254501
rect 769 253713 781 254489
rect 815 253713 831 254489
rect 769 253701 831 253713
rect 861 254489 923 254501
rect 861 253713 877 254489
rect 911 253713 923 254489
rect 861 253701 923 253713
rect 979 254489 1041 254501
rect 979 253713 991 254489
rect 1025 253713 1041 254489
rect 979 253701 1041 253713
rect 1071 254489 1133 254501
rect 1071 253713 1087 254489
rect 1121 253713 1133 254489
rect 1071 253701 1133 253713
rect 1189 254489 1251 254501
rect 1189 253713 1201 254489
rect 1235 253713 1251 254489
rect 1189 253701 1251 253713
rect 1281 254489 1343 254501
rect 1281 253713 1297 254489
rect 1331 253713 1343 254489
rect 1281 253701 1343 253713
rect 1399 254489 1461 254501
rect 1399 253713 1411 254489
rect 1445 253713 1461 254489
rect 1399 253701 1461 253713
rect 1491 254489 1553 254501
rect 1491 253713 1507 254489
rect 1541 253713 1553 254489
rect 1491 253701 1553 253713
rect 1609 254489 1671 254501
rect 1609 253713 1621 254489
rect 1655 253713 1671 254489
rect 1609 253701 1671 253713
rect 1701 254489 1763 254501
rect 1701 253713 1717 254489
rect 1751 253713 1763 254489
rect 1701 253701 1763 253713
rect 1819 254489 1881 254501
rect 1819 253713 1831 254489
rect 1865 253713 1881 254489
rect 1819 253701 1881 253713
rect 1911 254489 1973 254501
rect 1911 253713 1927 254489
rect 1961 253713 1973 254489
rect 1911 253701 1973 253713
rect 2029 254489 2091 254501
rect 2029 253713 2041 254489
rect 2075 253713 2091 254489
rect 2029 253701 2091 253713
rect 2121 254489 2183 254501
rect 2121 253713 2137 254489
rect 2171 253713 2183 254489
rect 2121 253701 2183 253713
rect 2239 254489 2301 254501
rect 2239 253713 2251 254489
rect 2285 253713 2301 254489
rect 2239 253701 2301 253713
rect 2331 254489 2393 254501
rect 2331 253713 2347 254489
rect 2381 253713 2393 254489
rect 2331 253701 2393 253713
rect 2449 254489 2511 254501
rect 2449 253713 2461 254489
rect 2495 253713 2511 254489
rect 2449 253701 2511 253713
rect 2541 254489 2603 254501
rect 2541 253713 2557 254489
rect 2591 253713 2603 254489
rect 2541 253701 2603 253713
rect 2659 254489 2721 254501
rect 2659 253713 2671 254489
rect 2705 253713 2721 254489
rect 2659 253701 2721 253713
rect 2751 254489 2813 254501
rect 2751 253713 2767 254489
rect 2801 253713 2813 254489
rect 2751 253701 2813 253713
rect 2869 254489 2931 254501
rect 2869 253713 2881 254489
rect 2915 253713 2931 254489
rect 2869 253701 2931 253713
rect 2961 254489 3023 254501
rect 2961 253713 2977 254489
rect 3011 253713 3023 254489
rect 2961 253701 3023 253713
rect 3079 254489 3141 254501
rect 3079 253713 3091 254489
rect 3125 253713 3141 254489
rect 3079 253701 3141 253713
rect 3171 254489 3233 254501
rect 3171 253713 3187 254489
rect 3221 253713 3233 254489
rect 3171 253701 3233 253713
rect 3289 254489 3351 254501
rect 3289 253713 3301 254489
rect 3335 253713 3351 254489
rect 3289 253701 3351 253713
rect 3381 254489 3443 254501
rect 3381 253713 3397 254489
rect 3431 253713 3443 254489
rect 3381 253701 3443 253713
rect 3499 254489 3561 254501
rect 3499 253713 3511 254489
rect 3545 253713 3561 254489
rect 3499 253701 3561 253713
rect 3591 254489 3653 254501
rect 3591 253713 3607 254489
rect 3641 253713 3653 254489
rect 3591 253701 3653 253713
rect 3709 254489 3771 254501
rect 3709 253713 3721 254489
rect 3755 253713 3771 254489
rect 3709 253701 3771 253713
rect 3801 254489 3863 254501
rect 3801 253713 3817 254489
rect 3851 253713 3863 254489
rect 3801 253701 3863 253713
rect 3919 254489 3981 254501
rect 3919 253713 3931 254489
rect 3965 253713 3981 254489
rect 3919 253701 3981 253713
rect 4011 254489 4073 254501
rect 4011 253713 4027 254489
rect 4061 253713 4073 254489
rect 4011 253701 4073 253713
rect 4129 254489 4191 254501
rect 4129 253713 4141 254489
rect 4175 253713 4191 254489
rect 4129 253701 4191 253713
rect 4221 254489 4283 254501
rect 4221 253713 4237 254489
rect 4271 253713 4283 254489
rect 4221 253701 4283 253713
rect 4339 254489 4401 254501
rect 4339 253713 4351 254489
rect 4385 253713 4401 254489
rect 4339 253701 4401 253713
rect 4431 254489 4493 254501
rect 4431 253713 4447 254489
rect 4481 253713 4493 254489
rect 4431 253701 4493 253713
rect 4549 254489 4611 254501
rect 4549 253713 4561 254489
rect 4595 253713 4611 254489
rect 4549 253701 4611 253713
rect 4641 254489 4703 254501
rect 4641 253713 4657 254489
rect 4691 253713 4703 254489
rect 4641 253701 4703 253713
rect 4759 254489 4821 254501
rect 4759 253713 4771 254489
rect 4805 253713 4821 254489
rect 4759 253701 4821 253713
rect 4851 254489 4913 254501
rect 4851 253713 4867 254489
rect 4901 253713 4913 254489
rect 4851 253701 4913 253713
rect 4969 254489 5031 254501
rect 4969 253713 4981 254489
rect 5015 253713 5031 254489
rect 4969 253701 5031 253713
rect 5061 254489 5123 254501
rect 5061 253713 5077 254489
rect 5111 253713 5123 254489
rect 5061 253701 5123 253713
rect 5179 254489 5241 254501
rect 5179 253713 5191 254489
rect 5225 253713 5241 254489
rect 5179 253701 5241 253713
rect 5271 254489 5333 254501
rect 5271 253713 5287 254489
rect 5321 253713 5333 254489
rect 5271 253701 5333 253713
rect 5389 254489 5451 254501
rect 5389 253713 5401 254489
rect 5435 253713 5451 254489
rect 5389 253701 5451 253713
rect 5481 254489 5543 254501
rect 5481 253713 5497 254489
rect 5531 253713 5543 254489
rect 5481 253701 5543 253713
rect 5599 254489 5661 254501
rect 5599 253713 5611 254489
rect 5645 253713 5661 254489
rect 5599 253701 5661 253713
rect 5691 254489 5753 254501
rect 5691 253713 5707 254489
rect 5741 253713 5753 254489
rect 5691 253701 5753 253713
rect 5809 254489 5871 254501
rect 5809 253713 5821 254489
rect 5855 253713 5871 254489
rect 5809 253701 5871 253713
rect 5901 254489 5963 254501
rect 5901 253713 5917 254489
rect 5951 253713 5963 254489
rect 5901 253701 5963 253713
rect 6019 254489 6081 254501
rect 6019 253713 6031 254489
rect 6065 253713 6081 254489
rect 6019 253701 6081 253713
rect 6111 254489 6173 254501
rect 6111 253713 6127 254489
rect 6161 253713 6173 254489
rect 6111 253701 6173 253713
rect 6229 254489 6291 254501
rect 6229 253713 6241 254489
rect 6275 253713 6291 254489
rect 6229 253701 6291 253713
rect 6321 254489 6383 254501
rect 6321 253713 6337 254489
rect 6371 253713 6383 254489
rect 6321 253701 6383 253713
rect 6439 254489 6501 254501
rect 6439 253713 6451 254489
rect 6485 253713 6501 254489
rect 6439 253701 6501 253713
rect 6531 254489 6593 254501
rect 6531 253713 6547 254489
rect 6581 253713 6593 254489
rect 6531 253701 6593 253713
rect 6649 254489 6711 254501
rect 6649 253713 6661 254489
rect 6695 253713 6711 254489
rect 6649 253701 6711 253713
rect 6741 254489 6803 254501
rect 6741 253713 6757 254489
rect 6791 253713 6803 254489
rect 6741 253701 6803 253713
rect 6859 254489 6921 254501
rect 6859 253713 6871 254489
rect 6905 253713 6921 254489
rect 6859 253701 6921 253713
rect 6951 254489 7013 254501
rect 6951 253713 6967 254489
rect 7001 253713 7013 254489
rect 6951 253701 7013 253713
rect 7069 254489 7131 254501
rect 7069 253713 7081 254489
rect 7115 253713 7131 254489
rect 7069 253701 7131 253713
rect 7161 254489 7223 254501
rect 7161 253713 7177 254489
rect 7211 253713 7223 254489
rect 7161 253701 7223 253713
rect 7279 254489 7341 254501
rect 7279 253713 7291 254489
rect 7325 253713 7341 254489
rect 7279 253701 7341 253713
rect 7371 254489 7433 254501
rect 7371 253713 7387 254489
rect 7421 253713 7433 254489
rect 7371 253701 7433 253713
rect 7489 254489 7551 254501
rect 7489 253713 7501 254489
rect 7535 253713 7551 254489
rect 7489 253701 7551 253713
rect 7581 254489 7643 254501
rect 7581 253713 7597 254489
rect 7631 253713 7643 254489
rect 7581 253701 7643 253713
rect 7699 254489 7761 254501
rect 7699 253713 7711 254489
rect 7745 253713 7761 254489
rect 7699 253701 7761 253713
rect 7791 254489 7853 254501
rect 7791 253713 7807 254489
rect 7841 253713 7853 254489
rect 7791 253701 7853 253713
rect 7909 254489 7971 254501
rect 7909 253713 7921 254489
rect 7955 253713 7971 254489
rect 7909 253701 7971 253713
rect 8001 254489 8063 254501
rect 8001 253713 8017 254489
rect 8051 253713 8063 254489
rect 8001 253701 8063 253713
rect 8119 254489 8181 254501
rect 8119 253713 8131 254489
rect 8165 253713 8181 254489
rect 8119 253701 8181 253713
rect 8211 254489 8273 254501
rect 8211 253713 8227 254489
rect 8261 253713 8273 254489
rect 8211 253701 8273 253713
rect 8329 254489 8391 254501
rect 8329 253713 8341 254489
rect 8375 253713 8391 254489
rect 8329 253701 8391 253713
rect 8421 254489 8483 254501
rect 8421 253713 8437 254489
rect 8471 253713 8483 254489
rect 8421 253701 8483 253713
rect 8539 254489 8601 254501
rect 8539 253713 8551 254489
rect 8585 253713 8601 254489
rect 8539 253701 8601 253713
rect 8631 254489 8693 254501
rect 8631 253713 8647 254489
rect 8681 253713 8693 254489
rect 8631 253701 8693 253713
rect 8749 254489 8811 254501
rect 8749 253713 8761 254489
rect 8795 253713 8811 254489
rect 8749 253701 8811 253713
rect 8841 254489 8903 254501
rect 8841 253713 8857 254489
rect 8891 253713 8903 254489
rect 8841 253701 8903 253713
rect 8959 254489 9021 254501
rect 8959 253713 8971 254489
rect 9005 253713 9021 254489
rect 8959 253701 9021 253713
rect 9051 254489 9113 254501
rect 9051 253713 9067 254489
rect 9101 253713 9113 254489
rect 9051 253701 9113 253713
rect 9169 254489 9231 254501
rect 9169 253713 9181 254489
rect 9215 253713 9231 254489
rect 9169 253701 9231 253713
rect 9261 254489 9323 254501
rect 9261 253713 9277 254489
rect 9311 253713 9323 254489
rect 9261 253701 9323 253713
rect 9379 254489 9441 254501
rect 9379 253713 9391 254489
rect 9425 253713 9441 254489
rect 9379 253701 9441 253713
rect 9471 254489 9533 254501
rect 9471 253713 9487 254489
rect 9521 253713 9533 254489
rect 9471 253701 9533 253713
rect 9589 254489 9651 254501
rect 9589 253713 9601 254489
rect 9635 253713 9651 254489
rect 9589 253701 9651 253713
rect 9681 254489 9743 254501
rect 9681 253713 9697 254489
rect 9731 253713 9743 254489
rect 9681 253701 9743 253713
rect 9799 254489 9861 254501
rect 9799 253713 9811 254489
rect 9845 253713 9861 254489
rect 9799 253701 9861 253713
rect 9891 254489 9953 254501
rect 9891 253713 9907 254489
rect 9941 253713 9953 254489
rect 9891 253701 9953 253713
rect 10009 254489 10071 254501
rect 10009 253713 10021 254489
rect 10055 253713 10071 254489
rect 10009 253701 10071 253713
rect 10101 254489 10163 254501
rect 10101 253713 10117 254489
rect 10151 253713 10163 254489
rect 10101 253701 10163 253713
rect 10219 254489 10281 254501
rect 10219 253713 10231 254489
rect 10265 253713 10281 254489
rect 10219 253701 10281 253713
rect 10311 254489 10373 254501
rect 10311 253713 10327 254489
rect 10361 253713 10373 254489
rect 10311 253701 10373 253713
rect 10429 254489 10491 254501
rect 10429 253713 10441 254489
rect 10475 253713 10491 254489
rect 10429 253701 10491 253713
rect 10521 254489 10583 254501
rect 10521 253713 10537 254489
rect 10571 253713 10583 254489
rect 10521 253701 10583 253713
rect 10639 254489 10701 254501
rect 10639 253713 10651 254489
rect 10685 253713 10701 254489
rect 10639 253701 10701 253713
rect 10731 254489 10793 254501
rect 10731 253713 10747 254489
rect 10781 253713 10793 254489
rect 10731 253701 10793 253713
rect 10849 254489 10911 254501
rect 10849 253713 10861 254489
rect 10895 253713 10911 254489
rect 10849 253701 10911 253713
rect 10941 254489 11003 254501
rect 10941 253713 10957 254489
rect 10991 253713 11003 254489
rect 10941 253701 11003 253713
rect 11059 254489 11121 254501
rect 11059 253713 11071 254489
rect 11105 253713 11121 254489
rect 11059 253701 11121 253713
rect 11151 254489 11213 254501
rect 11151 253713 11167 254489
rect 11201 253713 11213 254489
rect 11151 253701 11213 253713
rect 11269 254489 11331 254501
rect 11269 253713 11281 254489
rect 11315 253713 11331 254489
rect 11269 253701 11331 253713
rect 11361 254489 11423 254501
rect 11361 253713 11377 254489
rect 11411 253713 11423 254489
rect 11361 253701 11423 253713
rect 11479 254489 11541 254501
rect 11479 253713 11491 254489
rect 11525 253713 11541 254489
rect 11479 253701 11541 253713
rect 11571 254489 11633 254501
rect 11571 253713 11587 254489
rect 11621 253713 11633 254489
rect 11571 253701 11633 253713
rect 11689 254489 11751 254501
rect 11689 253713 11701 254489
rect 11735 253713 11751 254489
rect 11689 253701 11751 253713
rect 11781 254489 11843 254501
rect 11781 253713 11797 254489
rect 11831 253713 11843 254489
rect 11781 253701 11843 253713
rect 11899 254489 11961 254501
rect 11899 253713 11911 254489
rect 11945 253713 11961 254489
rect 11899 253701 11961 253713
rect 11991 254489 12053 254501
rect 11991 253713 12007 254489
rect 12041 253713 12053 254489
rect 11991 253701 12053 253713
rect 12109 254489 12171 254501
rect 12109 253713 12121 254489
rect 12155 253713 12171 254489
rect 12109 253701 12171 253713
rect 12201 254489 12263 254501
rect 12201 253713 12217 254489
rect 12251 253713 12263 254489
rect 12201 253701 12263 253713
rect 12319 254489 12381 254501
rect 12319 253713 12331 254489
rect 12365 253713 12381 254489
rect 12319 253701 12381 253713
rect 12411 254489 12473 254501
rect 12411 253713 12427 254489
rect 12461 253713 12473 254489
rect 12411 253701 12473 253713
rect 12529 254489 12591 254501
rect 12529 253713 12541 254489
rect 12575 253713 12591 254489
rect 12529 253701 12591 253713
rect 12621 254489 12683 254501
rect 12621 253713 12637 254489
rect 12671 253713 12683 254489
rect 12621 253701 12683 253713
rect 12739 254489 12801 254501
rect 12739 253713 12751 254489
rect 12785 253713 12801 254489
rect 12739 253701 12801 253713
rect 12831 254489 12893 254501
rect 12831 253713 12847 254489
rect 12881 253713 12893 254489
rect 12831 253701 12893 253713
rect 12949 254489 13011 254501
rect 12949 253713 12961 254489
rect 12995 253713 13011 254489
rect 12949 253701 13011 253713
rect 13041 254489 13103 254501
rect 13041 253713 13057 254489
rect 13091 253713 13103 254489
rect 13041 253701 13103 253713
rect 13159 254489 13221 254501
rect 13159 253713 13171 254489
rect 13205 253713 13221 254489
rect 13159 253701 13221 253713
rect 13251 254489 13313 254501
rect 13251 253713 13267 254489
rect 13301 253713 13313 254489
rect 13251 253701 13313 253713
rect 13369 254489 13431 254501
rect 13369 253713 13381 254489
rect 13415 253713 13431 254489
rect 13369 253701 13431 253713
rect 13461 254489 13523 254501
rect 13461 253713 13477 254489
rect 13511 253713 13523 254489
rect 13461 253701 13523 253713
rect 13579 254489 13641 254501
rect 13579 253713 13591 254489
rect 13625 253713 13641 254489
rect 13579 253701 13641 253713
rect 13671 254489 13733 254501
rect 13671 253713 13687 254489
rect 13721 253713 13733 254489
rect 13671 253701 13733 253713
rect 13789 254489 13851 254501
rect 13789 253713 13801 254489
rect 13835 253713 13851 254489
rect 13789 253701 13851 253713
rect 13881 254489 13943 254501
rect 13881 253713 13897 254489
rect 13931 253713 13943 254489
rect 13881 253701 13943 253713
rect 13999 254489 14061 254501
rect 13999 253713 14011 254489
rect 14045 253713 14061 254489
rect 13999 253701 14061 253713
rect 14091 254489 14153 254501
rect 14091 253713 14107 254489
rect 14141 253713 14153 254489
rect 14091 253701 14153 253713
rect 14209 254489 14271 254501
rect 14209 253713 14221 254489
rect 14255 253713 14271 254489
rect 14209 253701 14271 253713
rect 14301 254489 14363 254501
rect 14301 253713 14317 254489
rect 14351 253713 14363 254489
rect 14301 253701 14363 253713
rect 14419 254489 14481 254501
rect 14419 253713 14431 254489
rect 14465 253713 14481 254489
rect 14419 253701 14481 253713
rect 14511 254489 14573 254501
rect 14511 253713 14527 254489
rect 14561 253713 14573 254489
rect 14511 253701 14573 253713
rect 14629 254489 14691 254501
rect 14629 253713 14641 254489
rect 14675 253713 14691 254489
rect 14629 253701 14691 253713
rect 14721 254489 14783 254501
rect 14721 253713 14737 254489
rect 14771 253713 14783 254489
rect 14721 253701 14783 253713
rect 14839 254489 14901 254501
rect 14839 253713 14851 254489
rect 14885 253713 14901 254489
rect 14839 253701 14901 253713
rect 14931 254489 14993 254501
rect 14931 253713 14947 254489
rect 14981 253713 14993 254489
rect 14931 253701 14993 253713
rect 15049 254489 15111 254501
rect 15049 253713 15061 254489
rect 15095 253713 15111 254489
rect 15049 253701 15111 253713
rect 15141 254489 15203 254501
rect 15141 253713 15157 254489
rect 15191 253713 15203 254489
rect 15141 253701 15203 253713
rect 15259 254489 15321 254501
rect 15259 253713 15271 254489
rect 15305 253713 15321 254489
rect 15259 253701 15321 253713
rect 15351 254489 15413 254501
rect 15351 253713 15367 254489
rect 15401 253713 15413 254489
rect 15351 253701 15413 253713
rect 15469 254489 15531 254501
rect 15469 253713 15481 254489
rect 15515 253713 15531 254489
rect 15469 253701 15531 253713
rect 15561 254489 15623 254501
rect 15561 253713 15577 254489
rect 15611 253713 15623 254489
rect 15561 253701 15623 253713
rect 15679 254489 15741 254501
rect 15679 253713 15691 254489
rect 15725 253713 15741 254489
rect 15679 253701 15741 253713
rect 15771 254489 15833 254501
rect 15771 253713 15787 254489
rect 15821 253713 15833 254489
rect 15771 253701 15833 253713
rect 15889 254489 15951 254501
rect 15889 253713 15901 254489
rect 15935 253713 15951 254489
rect 15889 253701 15951 253713
rect 15981 254489 16043 254501
rect 15981 253713 15997 254489
rect 16031 253713 16043 254489
rect 15981 253701 16043 253713
rect 16099 254489 16161 254501
rect 16099 253713 16111 254489
rect 16145 253713 16161 254489
rect 16099 253701 16161 253713
rect 16191 254489 16253 254501
rect 16191 253713 16207 254489
rect 16241 253713 16253 254489
rect 16191 253701 16253 253713
rect 16309 254489 16371 254501
rect 16309 253713 16321 254489
rect 16355 253713 16371 254489
rect 16309 253701 16371 253713
rect 16401 254489 16463 254501
rect 16401 253713 16417 254489
rect 16451 253713 16463 254489
rect 16401 253701 16463 253713
rect 16519 254489 16581 254501
rect 16519 253713 16531 254489
rect 16565 253713 16581 254489
rect 16519 253701 16581 253713
rect 16611 254489 16673 254501
rect 16611 253713 16627 254489
rect 16661 253713 16673 254489
rect 16611 253701 16673 253713
rect 16729 254489 16791 254501
rect 16729 253713 16741 254489
rect 16775 253713 16791 254489
rect 16729 253701 16791 253713
rect 16821 254489 16883 254501
rect 16821 253713 16837 254489
rect 16871 253713 16883 254489
rect 16821 253701 16883 253713
rect 16939 254489 17001 254501
rect 16939 253713 16951 254489
rect 16985 253713 17001 254489
rect 16939 253701 17001 253713
rect 17031 254489 17093 254501
rect 17031 253713 17047 254489
rect 17081 253713 17093 254489
rect 17031 253701 17093 253713
rect 17149 254489 17211 254501
rect 17149 253713 17161 254489
rect 17195 253713 17211 254489
rect 17149 253701 17211 253713
rect 17241 254489 17303 254501
rect 17241 253713 17257 254489
rect 17291 253713 17303 254489
rect 17241 253701 17303 253713
rect 17359 254489 17421 254501
rect 17359 253713 17371 254489
rect 17405 253713 17421 254489
rect 17359 253701 17421 253713
rect 17451 254489 17513 254501
rect 17451 253713 17467 254489
rect 17501 253713 17513 254489
rect 17451 253701 17513 253713
rect 17569 254489 17631 254501
rect 17569 253713 17581 254489
rect 17615 253713 17631 254489
rect 17569 253701 17631 253713
rect 17661 254489 17723 254501
rect 17661 253713 17677 254489
rect 17711 253713 17723 254489
rect 17661 253701 17723 253713
rect 17779 254489 17841 254501
rect 17779 253713 17791 254489
rect 17825 253713 17841 254489
rect 17779 253701 17841 253713
rect 17871 254489 17933 254501
rect 17871 253713 17887 254489
rect 17921 253713 17933 254489
rect 17871 253701 17933 253713
rect 17989 254489 18051 254501
rect 17989 253713 18001 254489
rect 18035 253713 18051 254489
rect 17989 253701 18051 253713
rect 18081 254489 18143 254501
rect 18081 253713 18097 254489
rect 18131 253713 18143 254489
rect 18081 253701 18143 253713
rect 18199 254489 18261 254501
rect 18199 253713 18211 254489
rect 18245 253713 18261 254489
rect 18199 253701 18261 253713
rect 18291 254489 18353 254501
rect 18291 253713 18307 254489
rect 18341 253713 18353 254489
rect 18291 253701 18353 253713
rect 18409 254489 18471 254501
rect 18409 253713 18421 254489
rect 18455 253713 18471 254489
rect 18409 253701 18471 253713
rect 18501 254489 18563 254501
rect 18501 253713 18517 254489
rect 18551 253713 18563 254489
rect 18501 253701 18563 253713
rect 18619 254489 18681 254501
rect 18619 253713 18631 254489
rect 18665 253713 18681 254489
rect 18619 253701 18681 253713
rect 18711 254489 18773 254501
rect 18711 253713 18727 254489
rect 18761 253713 18773 254489
rect 18711 253701 18773 253713
rect 18829 254489 18891 254501
rect 18829 253713 18841 254489
rect 18875 253713 18891 254489
rect 18829 253701 18891 253713
rect 18921 254489 18983 254501
rect 18921 253713 18937 254489
rect 18971 253713 18983 254489
rect 18921 253701 18983 253713
rect 19039 254489 19101 254501
rect 19039 253713 19051 254489
rect 19085 253713 19101 254489
rect 19039 253701 19101 253713
rect 19131 254489 19193 254501
rect 19131 253713 19147 254489
rect 19181 253713 19193 254489
rect 19131 253701 19193 253713
rect 19249 254489 19311 254501
rect 19249 253713 19261 254489
rect 19295 253713 19311 254489
rect 19249 253701 19311 253713
rect 19341 254489 19403 254501
rect 19341 253713 19357 254489
rect 19391 253713 19403 254489
rect 19341 253701 19403 253713
rect 19459 254489 19521 254501
rect 19459 253713 19471 254489
rect 19505 253713 19521 254489
rect 19459 253701 19521 253713
rect 19551 254489 19613 254501
rect 19551 253713 19567 254489
rect 19601 253713 19613 254489
rect 19551 253701 19613 253713
rect 19669 254489 19731 254501
rect 19669 253713 19681 254489
rect 19715 253713 19731 254489
rect 19669 253701 19731 253713
rect 19761 254489 19823 254501
rect 19761 253713 19777 254489
rect 19811 253713 19823 254489
rect 19761 253701 19823 253713
rect 19879 254489 19941 254501
rect 19879 253713 19891 254489
rect 19925 253713 19941 254489
rect 19879 253701 19941 253713
rect 19971 254489 20033 254501
rect 19971 253713 19987 254489
rect 20021 253713 20033 254489
rect 19971 253701 20033 253713
rect 20089 254489 20151 254501
rect 20089 253713 20101 254489
rect 20135 253713 20151 254489
rect 20089 253701 20151 253713
rect 20181 254489 20243 254501
rect 20181 253713 20197 254489
rect 20231 253713 20243 254489
rect 20181 253701 20243 253713
rect 20299 254489 20361 254501
rect 20299 253713 20311 254489
rect 20345 253713 20361 254489
rect 20299 253701 20361 253713
rect 20391 254489 20453 254501
rect 20391 253713 20407 254489
rect 20441 253713 20453 254489
rect 20391 253701 20453 253713
rect 20509 254489 20571 254501
rect 20509 253713 20521 254489
rect 20555 253713 20571 254489
rect 20509 253701 20571 253713
rect 20601 254489 20663 254501
rect 20601 253713 20617 254489
rect 20651 253713 20663 254489
rect 20601 253701 20663 253713
rect 20719 254489 20781 254501
rect 20719 253713 20731 254489
rect 20765 253713 20781 254489
rect 20719 253701 20781 253713
rect 20811 254489 20873 254501
rect 20811 253713 20827 254489
rect 20861 253713 20873 254489
rect 20811 253701 20873 253713
rect 20929 254489 20991 254501
rect 20929 253713 20941 254489
rect 20975 253713 20991 254489
rect 20929 253701 20991 253713
rect 21021 254489 21083 254501
rect 21021 253713 21037 254489
rect 21071 253713 21083 254489
rect 21021 253701 21083 253713
rect 21139 254489 21201 254501
rect 21139 253713 21151 254489
rect 21185 253713 21201 254489
rect 21139 253701 21201 253713
rect 21231 254489 21293 254501
rect 21231 253713 21247 254489
rect 21281 253713 21293 254489
rect 21231 253701 21293 253713
rect 21349 254489 21411 254501
rect 21349 253713 21361 254489
rect 21395 253713 21411 254489
rect 21349 253701 21411 253713
rect 21441 254489 21503 254501
rect 21441 253713 21457 254489
rect 21491 253713 21503 254489
rect 21441 253701 21503 253713
rect 21559 254489 21621 254501
rect 21559 253713 21571 254489
rect 21605 253713 21621 254489
rect 21559 253701 21621 253713
rect 21651 254489 21713 254501
rect 21651 253713 21667 254489
rect 21701 253713 21713 254489
rect 21651 253701 21713 253713
rect 21769 254489 21831 254501
rect 21769 253713 21781 254489
rect 21815 253713 21831 254489
rect 21769 253701 21831 253713
rect 21861 254489 21923 254501
rect 21861 253713 21877 254489
rect 21911 253713 21923 254489
rect 21861 253701 21923 253713
rect 21979 254489 22041 254501
rect 21979 253713 21991 254489
rect 22025 253713 22041 254489
rect 21979 253701 22041 253713
rect 22071 254489 22133 254501
rect 22071 253713 22087 254489
rect 22121 253713 22133 254489
rect 22071 253701 22133 253713
rect 22189 254489 22251 254501
rect 22189 253713 22201 254489
rect 22235 253713 22251 254489
rect 22189 253701 22251 253713
rect 22281 254489 22343 254501
rect 22281 253713 22297 254489
rect 22331 253713 22343 254489
rect 22281 253701 22343 253713
rect 22399 254489 22461 254501
rect 22399 253713 22411 254489
rect 22445 253713 22461 254489
rect 22399 253701 22461 253713
rect 22491 254489 22553 254501
rect 22491 253713 22507 254489
rect 22541 253713 22553 254489
rect 22491 253701 22553 253713
rect 22609 254489 22671 254501
rect 22609 253713 22621 254489
rect 22655 253713 22671 254489
rect 22609 253701 22671 253713
rect 22701 254489 22763 254501
rect 22701 253713 22717 254489
rect 22751 253713 22763 254489
rect 22701 253701 22763 253713
rect 22819 254489 22881 254501
rect 22819 253713 22831 254489
rect 22865 253713 22881 254489
rect 22819 253701 22881 253713
rect 22911 254489 22973 254501
rect 22911 253713 22927 254489
rect 22961 253713 22973 254489
rect 22911 253701 22973 253713
rect 23029 254489 23091 254501
rect 23029 253713 23041 254489
rect 23075 253713 23091 254489
rect 23029 253701 23091 253713
rect 23121 254489 23183 254501
rect 23121 253713 23137 254489
rect 23171 253713 23183 254489
rect 23121 253701 23183 253713
rect 23239 254489 23301 254501
rect 23239 253713 23251 254489
rect 23285 253713 23301 254489
rect 23239 253701 23301 253713
rect 23331 254489 23393 254501
rect 23331 253713 23347 254489
rect 23381 253713 23393 254489
rect 23331 253701 23393 253713
rect 23449 254489 23511 254501
rect 23449 253713 23461 254489
rect 23495 253713 23511 254489
rect 23449 253701 23511 253713
rect 23541 254489 23603 254501
rect 23541 253713 23557 254489
rect 23591 253713 23603 254489
rect 23541 253701 23603 253713
rect 23659 254489 23721 254501
rect 23659 253713 23671 254489
rect 23705 253713 23721 254489
rect 23659 253701 23721 253713
rect 23751 254489 23813 254501
rect 23751 253713 23767 254489
rect 23801 253713 23813 254489
rect 23751 253701 23813 253713
rect 23869 254489 23931 254501
rect 23869 253713 23881 254489
rect 23915 253713 23931 254489
rect 23869 253701 23931 253713
rect 23961 254489 24023 254501
rect 23961 253713 23977 254489
rect 24011 253713 24023 254489
rect 23961 253701 24023 253713
rect 24079 254489 24141 254501
rect 24079 253713 24091 254489
rect 24125 253713 24141 254489
rect 24079 253701 24141 253713
rect 24171 254489 24233 254501
rect 24171 253713 24187 254489
rect 24221 253713 24233 254489
rect 24171 253701 24233 253713
rect 24289 254489 24351 254501
rect 24289 253713 24301 254489
rect 24335 253713 24351 254489
rect 24289 253701 24351 253713
rect 24381 254489 24443 254501
rect 24381 253713 24397 254489
rect 24431 253713 24443 254489
rect 24381 253701 24443 253713
rect 24499 254489 24561 254501
rect 24499 253713 24511 254489
rect 24545 253713 24561 254489
rect 24499 253701 24561 253713
rect 24591 254489 24653 254501
rect 24591 253713 24607 254489
rect 24641 253713 24653 254489
rect 24591 253701 24653 253713
rect 24709 254489 24771 254501
rect 24709 253713 24721 254489
rect 24755 253713 24771 254489
rect 24709 253701 24771 253713
rect 24801 254489 24863 254501
rect 24801 253713 24817 254489
rect 24851 253713 24863 254489
rect 24801 253701 24863 253713
rect 24919 254489 24981 254501
rect 24919 253713 24931 254489
rect 24965 253713 24981 254489
rect 24919 253701 24981 253713
rect 25011 254489 25073 254501
rect 25011 253713 25027 254489
rect 25061 253713 25073 254489
rect 25011 253701 25073 253713
rect 25129 254489 25191 254501
rect 25129 253713 25141 254489
rect 25175 253713 25191 254489
rect 25129 253701 25191 253713
rect 25221 254489 25283 254501
rect 25221 253713 25237 254489
rect 25271 253713 25283 254489
rect 25221 253701 25283 253713
rect 25339 254489 25401 254501
rect 25339 253713 25351 254489
rect 25385 253713 25401 254489
rect 25339 253701 25401 253713
rect 25431 254489 25493 254501
rect 25431 253713 25447 254489
rect 25481 253713 25493 254489
rect 25431 253701 25493 253713
rect 25549 254489 25611 254501
rect 25549 253713 25561 254489
rect 25595 253713 25611 254489
rect 25549 253701 25611 253713
rect 25641 254489 25703 254501
rect 25641 253713 25657 254489
rect 25691 253713 25703 254489
rect 25641 253701 25703 253713
rect 25759 254489 25821 254501
rect 25759 253713 25771 254489
rect 25805 253713 25821 254489
rect 25759 253701 25821 253713
rect 25851 254489 25913 254501
rect 25851 253713 25867 254489
rect 25901 253713 25913 254489
rect 25851 253701 25913 253713
rect 25969 254489 26031 254501
rect 25969 253713 25981 254489
rect 26015 253713 26031 254489
rect 25969 253701 26031 253713
rect 26061 254489 26123 254501
rect 26061 253713 26077 254489
rect 26111 253713 26123 254489
rect 26061 253701 26123 253713
rect 26179 254489 26241 254501
rect 26179 253713 26191 254489
rect 26225 253713 26241 254489
rect 26179 253701 26241 253713
rect 26271 254489 26333 254501
rect 26271 253713 26287 254489
rect 26321 253713 26333 254489
rect 26271 253701 26333 253713
rect 26389 254489 26451 254501
rect 26389 253713 26401 254489
rect 26435 253713 26451 254489
rect 26389 253701 26451 253713
rect 26481 254489 26543 254501
rect 26481 253713 26497 254489
rect 26531 253713 26543 254489
rect 26481 253701 26543 253713
rect 26599 254489 26661 254501
rect 26599 253713 26611 254489
rect 26645 253713 26661 254489
rect 26599 253701 26661 253713
rect 26691 254489 26753 254501
rect 26691 253713 26707 254489
rect 26741 253713 26753 254489
rect 26691 253701 26753 253713
rect 26809 254489 26871 254501
rect 26809 253713 26821 254489
rect 26855 253713 26871 254489
rect 26809 253701 26871 253713
rect 26901 254489 26963 254501
rect 26901 253713 26917 254489
rect 26951 253713 26963 254489
rect 26901 253701 26963 253713
rect 27019 254489 27081 254501
rect 27019 253713 27031 254489
rect 27065 253713 27081 254489
rect 27019 253701 27081 253713
rect 27111 254489 27173 254501
rect 27111 253713 27127 254489
rect 27161 253713 27173 254489
rect 27111 253701 27173 253713
rect 27229 254489 27291 254501
rect 27229 253713 27241 254489
rect 27275 253713 27291 254489
rect 27229 253701 27291 253713
rect 27321 254489 27383 254501
rect 27321 253713 27337 254489
rect 27371 253713 27383 254489
rect 27321 253701 27383 253713
rect -4061 253453 -3999 253465
rect -4061 252677 -4049 253453
rect -4015 252677 -3999 253453
rect -4061 252665 -3999 252677
rect -3969 253453 -3907 253465
rect -3969 252677 -3953 253453
rect -3919 252677 -3907 253453
rect -3969 252665 -3907 252677
rect -3851 253453 -3789 253465
rect -3851 252677 -3839 253453
rect -3805 252677 -3789 253453
rect -3851 252665 -3789 252677
rect -3759 253453 -3697 253465
rect -3759 252677 -3743 253453
rect -3709 252677 -3697 253453
rect -3759 252665 -3697 252677
rect -3641 253453 -3579 253465
rect -3641 252677 -3629 253453
rect -3595 252677 -3579 253453
rect -3641 252665 -3579 252677
rect -3549 253453 -3487 253465
rect -3549 252677 -3533 253453
rect -3499 252677 -3487 253453
rect -3549 252665 -3487 252677
rect -3431 253453 -3369 253465
rect -3431 252677 -3419 253453
rect -3385 252677 -3369 253453
rect -3431 252665 -3369 252677
rect -3339 253453 -3277 253465
rect -3339 252677 -3323 253453
rect -3289 252677 -3277 253453
rect -3339 252665 -3277 252677
rect -3221 253453 -3159 253465
rect -3221 252677 -3209 253453
rect -3175 252677 -3159 253453
rect -3221 252665 -3159 252677
rect -3129 253453 -3067 253465
rect -3129 252677 -3113 253453
rect -3079 252677 -3067 253453
rect -3129 252665 -3067 252677
rect -3011 253453 -2949 253465
rect -3011 252677 -2999 253453
rect -2965 252677 -2949 253453
rect -3011 252665 -2949 252677
rect -2919 253453 -2857 253465
rect -2919 252677 -2903 253453
rect -2869 252677 -2857 253453
rect -2919 252665 -2857 252677
rect -2801 253453 -2739 253465
rect -2801 252677 -2789 253453
rect -2755 252677 -2739 253453
rect -2801 252665 -2739 252677
rect -2709 253453 -2647 253465
rect -2709 252677 -2693 253453
rect -2659 252677 -2647 253453
rect -2709 252665 -2647 252677
rect -2591 253453 -2529 253465
rect -2591 252677 -2579 253453
rect -2545 252677 -2529 253453
rect -2591 252665 -2529 252677
rect -2499 253453 -2437 253465
rect -2499 252677 -2483 253453
rect -2449 252677 -2437 253453
rect -2499 252665 -2437 252677
rect -2381 253453 -2319 253465
rect -2381 252677 -2369 253453
rect -2335 252677 -2319 253453
rect -2381 252665 -2319 252677
rect -2289 253453 -2227 253465
rect -2289 252677 -2273 253453
rect -2239 252677 -2227 253453
rect -2289 252665 -2227 252677
rect -2171 253453 -2109 253465
rect -2171 252677 -2159 253453
rect -2125 252677 -2109 253453
rect -2171 252665 -2109 252677
rect -2079 253453 -2017 253465
rect -2079 252677 -2063 253453
rect -2029 252677 -2017 253453
rect -2079 252665 -2017 252677
rect -1961 253453 -1899 253465
rect -1961 252677 -1949 253453
rect -1915 252677 -1899 253453
rect -1961 252665 -1899 252677
rect -1869 253453 -1807 253465
rect -1869 252677 -1853 253453
rect -1819 252677 -1807 253453
rect -1869 252665 -1807 252677
rect -1751 253453 -1689 253465
rect -1751 252677 -1739 253453
rect -1705 252677 -1689 253453
rect -1751 252665 -1689 252677
rect -1659 253453 -1597 253465
rect -1659 252677 -1643 253453
rect -1609 252677 -1597 253453
rect -1659 252665 -1597 252677
rect -1541 253453 -1479 253465
rect -1541 252677 -1529 253453
rect -1495 252677 -1479 253453
rect -1541 252665 -1479 252677
rect -1449 253453 -1387 253465
rect -1449 252677 -1433 253453
rect -1399 252677 -1387 253453
rect -1449 252665 -1387 252677
rect -1331 253453 -1269 253465
rect -1331 252677 -1319 253453
rect -1285 252677 -1269 253453
rect -1331 252665 -1269 252677
rect -1239 253453 -1177 253465
rect -1239 252677 -1223 253453
rect -1189 252677 -1177 253453
rect -1239 252665 -1177 252677
rect -1121 253453 -1059 253465
rect -1121 252677 -1109 253453
rect -1075 252677 -1059 253453
rect -1121 252665 -1059 252677
rect -1029 253453 -967 253465
rect -1029 252677 -1013 253453
rect -979 252677 -967 253453
rect -1029 252665 -967 252677
rect -911 253453 -849 253465
rect -911 252677 -899 253453
rect -865 252677 -849 253453
rect -911 252665 -849 252677
rect -819 253453 -757 253465
rect -819 252677 -803 253453
rect -769 252677 -757 253453
rect -819 252665 -757 252677
rect -701 253453 -639 253465
rect -701 252677 -689 253453
rect -655 252677 -639 253453
rect -701 252665 -639 252677
rect -609 253453 -547 253465
rect -609 252677 -593 253453
rect -559 252677 -547 253453
rect -609 252665 -547 252677
rect -491 253453 -429 253465
rect -491 252677 -479 253453
rect -445 252677 -429 253453
rect -491 252665 -429 252677
rect -399 253453 -337 253465
rect -399 252677 -383 253453
rect -349 252677 -337 253453
rect -399 252665 -337 252677
rect -281 253453 -219 253465
rect -281 252677 -269 253453
rect -235 252677 -219 253453
rect -281 252665 -219 252677
rect -189 253453 -127 253465
rect -189 252677 -173 253453
rect -139 252677 -127 253453
rect -189 252665 -127 252677
rect -71 253453 -9 253465
rect -71 252677 -59 253453
rect -25 252677 -9 253453
rect -71 252665 -9 252677
rect 21 253453 83 253465
rect 21 252677 37 253453
rect 71 252677 83 253453
rect 21 252665 83 252677
rect 139 253453 201 253465
rect 139 252677 151 253453
rect 185 252677 201 253453
rect 139 252665 201 252677
rect 231 253453 293 253465
rect 231 252677 247 253453
rect 281 252677 293 253453
rect 231 252665 293 252677
rect 349 253453 411 253465
rect 349 252677 361 253453
rect 395 252677 411 253453
rect 349 252665 411 252677
rect 441 253453 503 253465
rect 441 252677 457 253453
rect 491 252677 503 253453
rect 441 252665 503 252677
rect 559 253453 621 253465
rect 559 252677 571 253453
rect 605 252677 621 253453
rect 559 252665 621 252677
rect 651 253453 713 253465
rect 651 252677 667 253453
rect 701 252677 713 253453
rect 651 252665 713 252677
rect 769 253453 831 253465
rect 769 252677 781 253453
rect 815 252677 831 253453
rect 769 252665 831 252677
rect 861 253453 923 253465
rect 861 252677 877 253453
rect 911 252677 923 253453
rect 861 252665 923 252677
rect 979 253453 1041 253465
rect 979 252677 991 253453
rect 1025 252677 1041 253453
rect 979 252665 1041 252677
rect 1071 253453 1133 253465
rect 1071 252677 1087 253453
rect 1121 252677 1133 253453
rect 1071 252665 1133 252677
rect 1189 253453 1251 253465
rect 1189 252677 1201 253453
rect 1235 252677 1251 253453
rect 1189 252665 1251 252677
rect 1281 253453 1343 253465
rect 1281 252677 1297 253453
rect 1331 252677 1343 253453
rect 1281 252665 1343 252677
rect 1399 253453 1461 253465
rect 1399 252677 1411 253453
rect 1445 252677 1461 253453
rect 1399 252665 1461 252677
rect 1491 253453 1553 253465
rect 1491 252677 1507 253453
rect 1541 252677 1553 253453
rect 1491 252665 1553 252677
rect 1609 253453 1671 253465
rect 1609 252677 1621 253453
rect 1655 252677 1671 253453
rect 1609 252665 1671 252677
rect 1701 253453 1763 253465
rect 1701 252677 1717 253453
rect 1751 252677 1763 253453
rect 1701 252665 1763 252677
rect 1819 253453 1881 253465
rect 1819 252677 1831 253453
rect 1865 252677 1881 253453
rect 1819 252665 1881 252677
rect 1911 253453 1973 253465
rect 1911 252677 1927 253453
rect 1961 252677 1973 253453
rect 1911 252665 1973 252677
rect 2029 253453 2091 253465
rect 2029 252677 2041 253453
rect 2075 252677 2091 253453
rect 2029 252665 2091 252677
rect 2121 253453 2183 253465
rect 2121 252677 2137 253453
rect 2171 252677 2183 253453
rect 2121 252665 2183 252677
rect 2239 253453 2301 253465
rect 2239 252677 2251 253453
rect 2285 252677 2301 253453
rect 2239 252665 2301 252677
rect 2331 253453 2393 253465
rect 2331 252677 2347 253453
rect 2381 252677 2393 253453
rect 2331 252665 2393 252677
rect 2449 253453 2511 253465
rect 2449 252677 2461 253453
rect 2495 252677 2511 253453
rect 2449 252665 2511 252677
rect 2541 253453 2603 253465
rect 2541 252677 2557 253453
rect 2591 252677 2603 253453
rect 2541 252665 2603 252677
rect 2659 253453 2721 253465
rect 2659 252677 2671 253453
rect 2705 252677 2721 253453
rect 2659 252665 2721 252677
rect 2751 253453 2813 253465
rect 2751 252677 2767 253453
rect 2801 252677 2813 253453
rect 2751 252665 2813 252677
rect 2869 253453 2931 253465
rect 2869 252677 2881 253453
rect 2915 252677 2931 253453
rect 2869 252665 2931 252677
rect 2961 253453 3023 253465
rect 2961 252677 2977 253453
rect 3011 252677 3023 253453
rect 2961 252665 3023 252677
rect 3079 253453 3141 253465
rect 3079 252677 3091 253453
rect 3125 252677 3141 253453
rect 3079 252665 3141 252677
rect 3171 253453 3233 253465
rect 3171 252677 3187 253453
rect 3221 252677 3233 253453
rect 3171 252665 3233 252677
rect 3289 253453 3351 253465
rect 3289 252677 3301 253453
rect 3335 252677 3351 253453
rect 3289 252665 3351 252677
rect 3381 253453 3443 253465
rect 3381 252677 3397 253453
rect 3431 252677 3443 253453
rect 3381 252665 3443 252677
rect 3499 253453 3561 253465
rect 3499 252677 3511 253453
rect 3545 252677 3561 253453
rect 3499 252665 3561 252677
rect 3591 253453 3653 253465
rect 3591 252677 3607 253453
rect 3641 252677 3653 253453
rect 3591 252665 3653 252677
rect 3709 253453 3771 253465
rect 3709 252677 3721 253453
rect 3755 252677 3771 253453
rect 3709 252665 3771 252677
rect 3801 253453 3863 253465
rect 3801 252677 3817 253453
rect 3851 252677 3863 253453
rect 3801 252665 3863 252677
rect 3919 253453 3981 253465
rect 3919 252677 3931 253453
rect 3965 252677 3981 253453
rect 3919 252665 3981 252677
rect 4011 253453 4073 253465
rect 4011 252677 4027 253453
rect 4061 252677 4073 253453
rect 4011 252665 4073 252677
rect 4129 253453 4191 253465
rect 4129 252677 4141 253453
rect 4175 252677 4191 253453
rect 4129 252665 4191 252677
rect 4221 253453 4283 253465
rect 4221 252677 4237 253453
rect 4271 252677 4283 253453
rect 4221 252665 4283 252677
rect 4339 253453 4401 253465
rect 4339 252677 4351 253453
rect 4385 252677 4401 253453
rect 4339 252665 4401 252677
rect 4431 253453 4493 253465
rect 4431 252677 4447 253453
rect 4481 252677 4493 253453
rect 4431 252665 4493 252677
rect 4549 253453 4611 253465
rect 4549 252677 4561 253453
rect 4595 252677 4611 253453
rect 4549 252665 4611 252677
rect 4641 253453 4703 253465
rect 4641 252677 4657 253453
rect 4691 252677 4703 253453
rect 4641 252665 4703 252677
rect 4759 253453 4821 253465
rect 4759 252677 4771 253453
rect 4805 252677 4821 253453
rect 4759 252665 4821 252677
rect 4851 253453 4913 253465
rect 4851 252677 4867 253453
rect 4901 252677 4913 253453
rect 4851 252665 4913 252677
rect 4969 253453 5031 253465
rect 4969 252677 4981 253453
rect 5015 252677 5031 253453
rect 4969 252665 5031 252677
rect 5061 253453 5123 253465
rect 5061 252677 5077 253453
rect 5111 252677 5123 253453
rect 5061 252665 5123 252677
rect 5179 253453 5241 253465
rect 5179 252677 5191 253453
rect 5225 252677 5241 253453
rect 5179 252665 5241 252677
rect 5271 253453 5333 253465
rect 5271 252677 5287 253453
rect 5321 252677 5333 253453
rect 5271 252665 5333 252677
rect 5389 253453 5451 253465
rect 5389 252677 5401 253453
rect 5435 252677 5451 253453
rect 5389 252665 5451 252677
rect 5481 253453 5543 253465
rect 5481 252677 5497 253453
rect 5531 252677 5543 253453
rect 5481 252665 5543 252677
rect 5599 253453 5661 253465
rect 5599 252677 5611 253453
rect 5645 252677 5661 253453
rect 5599 252665 5661 252677
rect 5691 253453 5753 253465
rect 5691 252677 5707 253453
rect 5741 252677 5753 253453
rect 5691 252665 5753 252677
rect 5809 253453 5871 253465
rect 5809 252677 5821 253453
rect 5855 252677 5871 253453
rect 5809 252665 5871 252677
rect 5901 253453 5963 253465
rect 5901 252677 5917 253453
rect 5951 252677 5963 253453
rect 5901 252665 5963 252677
rect 6019 253453 6081 253465
rect 6019 252677 6031 253453
rect 6065 252677 6081 253453
rect 6019 252665 6081 252677
rect 6111 253453 6173 253465
rect 6111 252677 6127 253453
rect 6161 252677 6173 253453
rect 6111 252665 6173 252677
rect 6229 253453 6291 253465
rect 6229 252677 6241 253453
rect 6275 252677 6291 253453
rect 6229 252665 6291 252677
rect 6321 253453 6383 253465
rect 6321 252677 6337 253453
rect 6371 252677 6383 253453
rect 6321 252665 6383 252677
rect 6439 253453 6501 253465
rect 6439 252677 6451 253453
rect 6485 252677 6501 253453
rect 6439 252665 6501 252677
rect 6531 253453 6593 253465
rect 6531 252677 6547 253453
rect 6581 252677 6593 253453
rect 6531 252665 6593 252677
rect 6649 253453 6711 253465
rect 6649 252677 6661 253453
rect 6695 252677 6711 253453
rect 6649 252665 6711 252677
rect 6741 253453 6803 253465
rect 6741 252677 6757 253453
rect 6791 252677 6803 253453
rect 6741 252665 6803 252677
rect 6859 253453 6921 253465
rect 6859 252677 6871 253453
rect 6905 252677 6921 253453
rect 6859 252665 6921 252677
rect 6951 253453 7013 253465
rect 6951 252677 6967 253453
rect 7001 252677 7013 253453
rect 6951 252665 7013 252677
rect 7069 253453 7131 253465
rect 7069 252677 7081 253453
rect 7115 252677 7131 253453
rect 7069 252665 7131 252677
rect 7161 253453 7223 253465
rect 7161 252677 7177 253453
rect 7211 252677 7223 253453
rect 7161 252665 7223 252677
rect 7279 253453 7341 253465
rect 7279 252677 7291 253453
rect 7325 252677 7341 253453
rect 7279 252665 7341 252677
rect 7371 253453 7433 253465
rect 7371 252677 7387 253453
rect 7421 252677 7433 253453
rect 7371 252665 7433 252677
rect 7489 253453 7551 253465
rect 7489 252677 7501 253453
rect 7535 252677 7551 253453
rect 7489 252665 7551 252677
rect 7581 253453 7643 253465
rect 7581 252677 7597 253453
rect 7631 252677 7643 253453
rect 7581 252665 7643 252677
rect 7699 253453 7761 253465
rect 7699 252677 7711 253453
rect 7745 252677 7761 253453
rect 7699 252665 7761 252677
rect 7791 253453 7853 253465
rect 7791 252677 7807 253453
rect 7841 252677 7853 253453
rect 7791 252665 7853 252677
rect 7909 253453 7971 253465
rect 7909 252677 7921 253453
rect 7955 252677 7971 253453
rect 7909 252665 7971 252677
rect 8001 253453 8063 253465
rect 8001 252677 8017 253453
rect 8051 252677 8063 253453
rect 8001 252665 8063 252677
rect 8119 253453 8181 253465
rect 8119 252677 8131 253453
rect 8165 252677 8181 253453
rect 8119 252665 8181 252677
rect 8211 253453 8273 253465
rect 8211 252677 8227 253453
rect 8261 252677 8273 253453
rect 8211 252665 8273 252677
rect 8329 253453 8391 253465
rect 8329 252677 8341 253453
rect 8375 252677 8391 253453
rect 8329 252665 8391 252677
rect 8421 253453 8483 253465
rect 8421 252677 8437 253453
rect 8471 252677 8483 253453
rect 8421 252665 8483 252677
rect 8539 253453 8601 253465
rect 8539 252677 8551 253453
rect 8585 252677 8601 253453
rect 8539 252665 8601 252677
rect 8631 253453 8693 253465
rect 8631 252677 8647 253453
rect 8681 252677 8693 253453
rect 8631 252665 8693 252677
rect 8749 253453 8811 253465
rect 8749 252677 8761 253453
rect 8795 252677 8811 253453
rect 8749 252665 8811 252677
rect 8841 253453 8903 253465
rect 8841 252677 8857 253453
rect 8891 252677 8903 253453
rect 8841 252665 8903 252677
rect 8959 253453 9021 253465
rect 8959 252677 8971 253453
rect 9005 252677 9021 253453
rect 8959 252665 9021 252677
rect 9051 253453 9113 253465
rect 9051 252677 9067 253453
rect 9101 252677 9113 253453
rect 9051 252665 9113 252677
rect 9169 253453 9231 253465
rect 9169 252677 9181 253453
rect 9215 252677 9231 253453
rect 9169 252665 9231 252677
rect 9261 253453 9323 253465
rect 9261 252677 9277 253453
rect 9311 252677 9323 253453
rect 9261 252665 9323 252677
rect 9379 253453 9441 253465
rect 9379 252677 9391 253453
rect 9425 252677 9441 253453
rect 9379 252665 9441 252677
rect 9471 253453 9533 253465
rect 9471 252677 9487 253453
rect 9521 252677 9533 253453
rect 9471 252665 9533 252677
rect 9589 253453 9651 253465
rect 9589 252677 9601 253453
rect 9635 252677 9651 253453
rect 9589 252665 9651 252677
rect 9681 253453 9743 253465
rect 9681 252677 9697 253453
rect 9731 252677 9743 253453
rect 9681 252665 9743 252677
rect 9799 253453 9861 253465
rect 9799 252677 9811 253453
rect 9845 252677 9861 253453
rect 9799 252665 9861 252677
rect 9891 253453 9953 253465
rect 9891 252677 9907 253453
rect 9941 252677 9953 253453
rect 9891 252665 9953 252677
rect 10009 253453 10071 253465
rect 10009 252677 10021 253453
rect 10055 252677 10071 253453
rect 10009 252665 10071 252677
rect 10101 253453 10163 253465
rect 10101 252677 10117 253453
rect 10151 252677 10163 253453
rect 10101 252665 10163 252677
rect 10219 253453 10281 253465
rect 10219 252677 10231 253453
rect 10265 252677 10281 253453
rect 10219 252665 10281 252677
rect 10311 253453 10373 253465
rect 10311 252677 10327 253453
rect 10361 252677 10373 253453
rect 10311 252665 10373 252677
rect 10429 253453 10491 253465
rect 10429 252677 10441 253453
rect 10475 252677 10491 253453
rect 10429 252665 10491 252677
rect 10521 253453 10583 253465
rect 10521 252677 10537 253453
rect 10571 252677 10583 253453
rect 10521 252665 10583 252677
rect 10639 253453 10701 253465
rect 10639 252677 10651 253453
rect 10685 252677 10701 253453
rect 10639 252665 10701 252677
rect 10731 253453 10793 253465
rect 10731 252677 10747 253453
rect 10781 252677 10793 253453
rect 10731 252665 10793 252677
rect 10849 253453 10911 253465
rect 10849 252677 10861 253453
rect 10895 252677 10911 253453
rect 10849 252665 10911 252677
rect 10941 253453 11003 253465
rect 10941 252677 10957 253453
rect 10991 252677 11003 253453
rect 10941 252665 11003 252677
rect 11059 253453 11121 253465
rect 11059 252677 11071 253453
rect 11105 252677 11121 253453
rect 11059 252665 11121 252677
rect 11151 253453 11213 253465
rect 11151 252677 11167 253453
rect 11201 252677 11213 253453
rect 11151 252665 11213 252677
rect 11269 253453 11331 253465
rect 11269 252677 11281 253453
rect 11315 252677 11331 253453
rect 11269 252665 11331 252677
rect 11361 253453 11423 253465
rect 11361 252677 11377 253453
rect 11411 252677 11423 253453
rect 11361 252665 11423 252677
rect 11479 253453 11541 253465
rect 11479 252677 11491 253453
rect 11525 252677 11541 253453
rect 11479 252665 11541 252677
rect 11571 253453 11633 253465
rect 11571 252677 11587 253453
rect 11621 252677 11633 253453
rect 11571 252665 11633 252677
rect 11689 253453 11751 253465
rect 11689 252677 11701 253453
rect 11735 252677 11751 253453
rect 11689 252665 11751 252677
rect 11781 253453 11843 253465
rect 11781 252677 11797 253453
rect 11831 252677 11843 253453
rect 11781 252665 11843 252677
rect 11899 253453 11961 253465
rect 11899 252677 11911 253453
rect 11945 252677 11961 253453
rect 11899 252665 11961 252677
rect 11991 253453 12053 253465
rect 11991 252677 12007 253453
rect 12041 252677 12053 253453
rect 11991 252665 12053 252677
rect 12109 253453 12171 253465
rect 12109 252677 12121 253453
rect 12155 252677 12171 253453
rect 12109 252665 12171 252677
rect 12201 253453 12263 253465
rect 12201 252677 12217 253453
rect 12251 252677 12263 253453
rect 12201 252665 12263 252677
rect 12319 253453 12381 253465
rect 12319 252677 12331 253453
rect 12365 252677 12381 253453
rect 12319 252665 12381 252677
rect 12411 253453 12473 253465
rect 12411 252677 12427 253453
rect 12461 252677 12473 253453
rect 12411 252665 12473 252677
rect 12529 253453 12591 253465
rect 12529 252677 12541 253453
rect 12575 252677 12591 253453
rect 12529 252665 12591 252677
rect 12621 253453 12683 253465
rect 12621 252677 12637 253453
rect 12671 252677 12683 253453
rect 12621 252665 12683 252677
rect 12739 253453 12801 253465
rect 12739 252677 12751 253453
rect 12785 252677 12801 253453
rect 12739 252665 12801 252677
rect 12831 253453 12893 253465
rect 12831 252677 12847 253453
rect 12881 252677 12893 253453
rect 12831 252665 12893 252677
rect 12949 253453 13011 253465
rect 12949 252677 12961 253453
rect 12995 252677 13011 253453
rect 12949 252665 13011 252677
rect 13041 253453 13103 253465
rect 13041 252677 13057 253453
rect 13091 252677 13103 253453
rect 13041 252665 13103 252677
rect 13159 253453 13221 253465
rect 13159 252677 13171 253453
rect 13205 252677 13221 253453
rect 13159 252665 13221 252677
rect 13251 253453 13313 253465
rect 13251 252677 13267 253453
rect 13301 252677 13313 253453
rect 13251 252665 13313 252677
rect 13369 253453 13431 253465
rect 13369 252677 13381 253453
rect 13415 252677 13431 253453
rect 13369 252665 13431 252677
rect 13461 253453 13523 253465
rect 13461 252677 13477 253453
rect 13511 252677 13523 253453
rect 13461 252665 13523 252677
rect 13579 253453 13641 253465
rect 13579 252677 13591 253453
rect 13625 252677 13641 253453
rect 13579 252665 13641 252677
rect 13671 253453 13733 253465
rect 13671 252677 13687 253453
rect 13721 252677 13733 253453
rect 13671 252665 13733 252677
rect 13789 253453 13851 253465
rect 13789 252677 13801 253453
rect 13835 252677 13851 253453
rect 13789 252665 13851 252677
rect 13881 253453 13943 253465
rect 13881 252677 13897 253453
rect 13931 252677 13943 253453
rect 13881 252665 13943 252677
rect 13999 253453 14061 253465
rect 13999 252677 14011 253453
rect 14045 252677 14061 253453
rect 13999 252665 14061 252677
rect 14091 253453 14153 253465
rect 14091 252677 14107 253453
rect 14141 252677 14153 253453
rect 14091 252665 14153 252677
rect 14209 253453 14271 253465
rect 14209 252677 14221 253453
rect 14255 252677 14271 253453
rect 14209 252665 14271 252677
rect 14301 253453 14363 253465
rect 14301 252677 14317 253453
rect 14351 252677 14363 253453
rect 14301 252665 14363 252677
rect 14419 253453 14481 253465
rect 14419 252677 14431 253453
rect 14465 252677 14481 253453
rect 14419 252665 14481 252677
rect 14511 253453 14573 253465
rect 14511 252677 14527 253453
rect 14561 252677 14573 253453
rect 14511 252665 14573 252677
rect 14629 253453 14691 253465
rect 14629 252677 14641 253453
rect 14675 252677 14691 253453
rect 14629 252665 14691 252677
rect 14721 253453 14783 253465
rect 14721 252677 14737 253453
rect 14771 252677 14783 253453
rect 14721 252665 14783 252677
rect 14839 253453 14901 253465
rect 14839 252677 14851 253453
rect 14885 252677 14901 253453
rect 14839 252665 14901 252677
rect 14931 253453 14993 253465
rect 14931 252677 14947 253453
rect 14981 252677 14993 253453
rect 14931 252665 14993 252677
rect 15049 253453 15111 253465
rect 15049 252677 15061 253453
rect 15095 252677 15111 253453
rect 15049 252665 15111 252677
rect 15141 253453 15203 253465
rect 15141 252677 15157 253453
rect 15191 252677 15203 253453
rect 15141 252665 15203 252677
rect 15259 253453 15321 253465
rect 15259 252677 15271 253453
rect 15305 252677 15321 253453
rect 15259 252665 15321 252677
rect 15351 253453 15413 253465
rect 15351 252677 15367 253453
rect 15401 252677 15413 253453
rect 15351 252665 15413 252677
rect 15469 253453 15531 253465
rect 15469 252677 15481 253453
rect 15515 252677 15531 253453
rect 15469 252665 15531 252677
rect 15561 253453 15623 253465
rect 15561 252677 15577 253453
rect 15611 252677 15623 253453
rect 15561 252665 15623 252677
rect 15679 253453 15741 253465
rect 15679 252677 15691 253453
rect 15725 252677 15741 253453
rect 15679 252665 15741 252677
rect 15771 253453 15833 253465
rect 15771 252677 15787 253453
rect 15821 252677 15833 253453
rect 15771 252665 15833 252677
rect 15889 253453 15951 253465
rect 15889 252677 15901 253453
rect 15935 252677 15951 253453
rect 15889 252665 15951 252677
rect 15981 253453 16043 253465
rect 15981 252677 15997 253453
rect 16031 252677 16043 253453
rect 15981 252665 16043 252677
rect 16099 253453 16161 253465
rect 16099 252677 16111 253453
rect 16145 252677 16161 253453
rect 16099 252665 16161 252677
rect 16191 253453 16253 253465
rect 16191 252677 16207 253453
rect 16241 252677 16253 253453
rect 16191 252665 16253 252677
rect 16309 253453 16371 253465
rect 16309 252677 16321 253453
rect 16355 252677 16371 253453
rect 16309 252665 16371 252677
rect 16401 253453 16463 253465
rect 16401 252677 16417 253453
rect 16451 252677 16463 253453
rect 16401 252665 16463 252677
rect 16519 253453 16581 253465
rect 16519 252677 16531 253453
rect 16565 252677 16581 253453
rect 16519 252665 16581 252677
rect 16611 253453 16673 253465
rect 16611 252677 16627 253453
rect 16661 252677 16673 253453
rect 16611 252665 16673 252677
rect 16729 253453 16791 253465
rect 16729 252677 16741 253453
rect 16775 252677 16791 253453
rect 16729 252665 16791 252677
rect 16821 253453 16883 253465
rect 16821 252677 16837 253453
rect 16871 252677 16883 253453
rect 16821 252665 16883 252677
rect 16939 253453 17001 253465
rect 16939 252677 16951 253453
rect 16985 252677 17001 253453
rect 16939 252665 17001 252677
rect 17031 253453 17093 253465
rect 17031 252677 17047 253453
rect 17081 252677 17093 253453
rect 17031 252665 17093 252677
rect 17149 253453 17211 253465
rect 17149 252677 17161 253453
rect 17195 252677 17211 253453
rect 17149 252665 17211 252677
rect 17241 253453 17303 253465
rect 17241 252677 17257 253453
rect 17291 252677 17303 253453
rect 17241 252665 17303 252677
rect 17359 253453 17421 253465
rect 17359 252677 17371 253453
rect 17405 252677 17421 253453
rect 17359 252665 17421 252677
rect 17451 253453 17513 253465
rect 17451 252677 17467 253453
rect 17501 252677 17513 253453
rect 17451 252665 17513 252677
rect 17569 253453 17631 253465
rect 17569 252677 17581 253453
rect 17615 252677 17631 253453
rect 17569 252665 17631 252677
rect 17661 253453 17723 253465
rect 17661 252677 17677 253453
rect 17711 252677 17723 253453
rect 17661 252665 17723 252677
rect 17779 253453 17841 253465
rect 17779 252677 17791 253453
rect 17825 252677 17841 253453
rect 17779 252665 17841 252677
rect 17871 253453 17933 253465
rect 17871 252677 17887 253453
rect 17921 252677 17933 253453
rect 17871 252665 17933 252677
rect 17989 253453 18051 253465
rect 17989 252677 18001 253453
rect 18035 252677 18051 253453
rect 17989 252665 18051 252677
rect 18081 253453 18143 253465
rect 18081 252677 18097 253453
rect 18131 252677 18143 253453
rect 18081 252665 18143 252677
rect 18199 253453 18261 253465
rect 18199 252677 18211 253453
rect 18245 252677 18261 253453
rect 18199 252665 18261 252677
rect 18291 253453 18353 253465
rect 18291 252677 18307 253453
rect 18341 252677 18353 253453
rect 18291 252665 18353 252677
rect 18409 253453 18471 253465
rect 18409 252677 18421 253453
rect 18455 252677 18471 253453
rect 18409 252665 18471 252677
rect 18501 253453 18563 253465
rect 18501 252677 18517 253453
rect 18551 252677 18563 253453
rect 18501 252665 18563 252677
rect 18619 253453 18681 253465
rect 18619 252677 18631 253453
rect 18665 252677 18681 253453
rect 18619 252665 18681 252677
rect 18711 253453 18773 253465
rect 18711 252677 18727 253453
rect 18761 252677 18773 253453
rect 18711 252665 18773 252677
rect 18829 253453 18891 253465
rect 18829 252677 18841 253453
rect 18875 252677 18891 253453
rect 18829 252665 18891 252677
rect 18921 253453 18983 253465
rect 18921 252677 18937 253453
rect 18971 252677 18983 253453
rect 18921 252665 18983 252677
rect 19039 253453 19101 253465
rect 19039 252677 19051 253453
rect 19085 252677 19101 253453
rect 19039 252665 19101 252677
rect 19131 253453 19193 253465
rect 19131 252677 19147 253453
rect 19181 252677 19193 253453
rect 19131 252665 19193 252677
rect 19249 253453 19311 253465
rect 19249 252677 19261 253453
rect 19295 252677 19311 253453
rect 19249 252665 19311 252677
rect 19341 253453 19403 253465
rect 19341 252677 19357 253453
rect 19391 252677 19403 253453
rect 19341 252665 19403 252677
rect 19459 253453 19521 253465
rect 19459 252677 19471 253453
rect 19505 252677 19521 253453
rect 19459 252665 19521 252677
rect 19551 253453 19613 253465
rect 19551 252677 19567 253453
rect 19601 252677 19613 253453
rect 19551 252665 19613 252677
rect 19669 253453 19731 253465
rect 19669 252677 19681 253453
rect 19715 252677 19731 253453
rect 19669 252665 19731 252677
rect 19761 253453 19823 253465
rect 19761 252677 19777 253453
rect 19811 252677 19823 253453
rect 19761 252665 19823 252677
rect 19879 253453 19941 253465
rect 19879 252677 19891 253453
rect 19925 252677 19941 253453
rect 19879 252665 19941 252677
rect 19971 253453 20033 253465
rect 19971 252677 19987 253453
rect 20021 252677 20033 253453
rect 19971 252665 20033 252677
rect 20089 253453 20151 253465
rect 20089 252677 20101 253453
rect 20135 252677 20151 253453
rect 20089 252665 20151 252677
rect 20181 253453 20243 253465
rect 20181 252677 20197 253453
rect 20231 252677 20243 253453
rect 20181 252665 20243 252677
rect 20299 253453 20361 253465
rect 20299 252677 20311 253453
rect 20345 252677 20361 253453
rect 20299 252665 20361 252677
rect 20391 253453 20453 253465
rect 20391 252677 20407 253453
rect 20441 252677 20453 253453
rect 20391 252665 20453 252677
rect 20509 253453 20571 253465
rect 20509 252677 20521 253453
rect 20555 252677 20571 253453
rect 20509 252665 20571 252677
rect 20601 253453 20663 253465
rect 20601 252677 20617 253453
rect 20651 252677 20663 253453
rect 20601 252665 20663 252677
rect 20719 253453 20781 253465
rect 20719 252677 20731 253453
rect 20765 252677 20781 253453
rect 20719 252665 20781 252677
rect 20811 253453 20873 253465
rect 20811 252677 20827 253453
rect 20861 252677 20873 253453
rect 20811 252665 20873 252677
rect 20929 253453 20991 253465
rect 20929 252677 20941 253453
rect 20975 252677 20991 253453
rect 20929 252665 20991 252677
rect 21021 253453 21083 253465
rect 21021 252677 21037 253453
rect 21071 252677 21083 253453
rect 21021 252665 21083 252677
rect 21139 253453 21201 253465
rect 21139 252677 21151 253453
rect 21185 252677 21201 253453
rect 21139 252665 21201 252677
rect 21231 253453 21293 253465
rect 21231 252677 21247 253453
rect 21281 252677 21293 253453
rect 21231 252665 21293 252677
rect 21349 253453 21411 253465
rect 21349 252677 21361 253453
rect 21395 252677 21411 253453
rect 21349 252665 21411 252677
rect 21441 253453 21503 253465
rect 21441 252677 21457 253453
rect 21491 252677 21503 253453
rect 21441 252665 21503 252677
rect 21559 253453 21621 253465
rect 21559 252677 21571 253453
rect 21605 252677 21621 253453
rect 21559 252665 21621 252677
rect 21651 253453 21713 253465
rect 21651 252677 21667 253453
rect 21701 252677 21713 253453
rect 21651 252665 21713 252677
rect 21769 253453 21831 253465
rect 21769 252677 21781 253453
rect 21815 252677 21831 253453
rect 21769 252665 21831 252677
rect 21861 253453 21923 253465
rect 21861 252677 21877 253453
rect 21911 252677 21923 253453
rect 21861 252665 21923 252677
rect 21979 253453 22041 253465
rect 21979 252677 21991 253453
rect 22025 252677 22041 253453
rect 21979 252665 22041 252677
rect 22071 253453 22133 253465
rect 22071 252677 22087 253453
rect 22121 252677 22133 253453
rect 22071 252665 22133 252677
rect 22189 253453 22251 253465
rect 22189 252677 22201 253453
rect 22235 252677 22251 253453
rect 22189 252665 22251 252677
rect 22281 253453 22343 253465
rect 22281 252677 22297 253453
rect 22331 252677 22343 253453
rect 22281 252665 22343 252677
rect 22399 253453 22461 253465
rect 22399 252677 22411 253453
rect 22445 252677 22461 253453
rect 22399 252665 22461 252677
rect 22491 253453 22553 253465
rect 22491 252677 22507 253453
rect 22541 252677 22553 253453
rect 22491 252665 22553 252677
rect 22609 253453 22671 253465
rect 22609 252677 22621 253453
rect 22655 252677 22671 253453
rect 22609 252665 22671 252677
rect 22701 253453 22763 253465
rect 22701 252677 22717 253453
rect 22751 252677 22763 253453
rect 22701 252665 22763 252677
rect 22819 253453 22881 253465
rect 22819 252677 22831 253453
rect 22865 252677 22881 253453
rect 22819 252665 22881 252677
rect 22911 253453 22973 253465
rect 22911 252677 22927 253453
rect 22961 252677 22973 253453
rect 22911 252665 22973 252677
rect 23029 253453 23091 253465
rect 23029 252677 23041 253453
rect 23075 252677 23091 253453
rect 23029 252665 23091 252677
rect 23121 253453 23183 253465
rect 23121 252677 23137 253453
rect 23171 252677 23183 253453
rect 23121 252665 23183 252677
rect 23239 253453 23301 253465
rect 23239 252677 23251 253453
rect 23285 252677 23301 253453
rect 23239 252665 23301 252677
rect 23331 253453 23393 253465
rect 23331 252677 23347 253453
rect 23381 252677 23393 253453
rect 23331 252665 23393 252677
rect 23449 253453 23511 253465
rect 23449 252677 23461 253453
rect 23495 252677 23511 253453
rect 23449 252665 23511 252677
rect 23541 253453 23603 253465
rect 23541 252677 23557 253453
rect 23591 252677 23603 253453
rect 23541 252665 23603 252677
rect 23659 253453 23721 253465
rect 23659 252677 23671 253453
rect 23705 252677 23721 253453
rect 23659 252665 23721 252677
rect 23751 253453 23813 253465
rect 23751 252677 23767 253453
rect 23801 252677 23813 253453
rect 23751 252665 23813 252677
rect 23869 253453 23931 253465
rect 23869 252677 23881 253453
rect 23915 252677 23931 253453
rect 23869 252665 23931 252677
rect 23961 253453 24023 253465
rect 23961 252677 23977 253453
rect 24011 252677 24023 253453
rect 23961 252665 24023 252677
rect 24079 253453 24141 253465
rect 24079 252677 24091 253453
rect 24125 252677 24141 253453
rect 24079 252665 24141 252677
rect 24171 253453 24233 253465
rect 24171 252677 24187 253453
rect 24221 252677 24233 253453
rect 24171 252665 24233 252677
rect 24289 253453 24351 253465
rect 24289 252677 24301 253453
rect 24335 252677 24351 253453
rect 24289 252665 24351 252677
rect 24381 253453 24443 253465
rect 24381 252677 24397 253453
rect 24431 252677 24443 253453
rect 24381 252665 24443 252677
rect 24499 253453 24561 253465
rect 24499 252677 24511 253453
rect 24545 252677 24561 253453
rect 24499 252665 24561 252677
rect 24591 253453 24653 253465
rect 24591 252677 24607 253453
rect 24641 252677 24653 253453
rect 24591 252665 24653 252677
rect 24709 253453 24771 253465
rect 24709 252677 24721 253453
rect 24755 252677 24771 253453
rect 24709 252665 24771 252677
rect 24801 253453 24863 253465
rect 24801 252677 24817 253453
rect 24851 252677 24863 253453
rect 24801 252665 24863 252677
rect 24919 253453 24981 253465
rect 24919 252677 24931 253453
rect 24965 252677 24981 253453
rect 24919 252665 24981 252677
rect 25011 253453 25073 253465
rect 25011 252677 25027 253453
rect 25061 252677 25073 253453
rect 25011 252665 25073 252677
rect 25129 253453 25191 253465
rect 25129 252677 25141 253453
rect 25175 252677 25191 253453
rect 25129 252665 25191 252677
rect 25221 253453 25283 253465
rect 25221 252677 25237 253453
rect 25271 252677 25283 253453
rect 25221 252665 25283 252677
rect 25339 253453 25401 253465
rect 25339 252677 25351 253453
rect 25385 252677 25401 253453
rect 25339 252665 25401 252677
rect 25431 253453 25493 253465
rect 25431 252677 25447 253453
rect 25481 252677 25493 253453
rect 25431 252665 25493 252677
rect 25549 253453 25611 253465
rect 25549 252677 25561 253453
rect 25595 252677 25611 253453
rect 25549 252665 25611 252677
rect 25641 253453 25703 253465
rect 25641 252677 25657 253453
rect 25691 252677 25703 253453
rect 25641 252665 25703 252677
rect 25759 253453 25821 253465
rect 25759 252677 25771 253453
rect 25805 252677 25821 253453
rect 25759 252665 25821 252677
rect 25851 253453 25913 253465
rect 25851 252677 25867 253453
rect 25901 252677 25913 253453
rect 25851 252665 25913 252677
rect 25969 253453 26031 253465
rect 25969 252677 25981 253453
rect 26015 252677 26031 253453
rect 25969 252665 26031 252677
rect 26061 253453 26123 253465
rect 26061 252677 26077 253453
rect 26111 252677 26123 253453
rect 26061 252665 26123 252677
rect 26179 253453 26241 253465
rect 26179 252677 26191 253453
rect 26225 252677 26241 253453
rect 26179 252665 26241 252677
rect 26271 253453 26333 253465
rect 26271 252677 26287 253453
rect 26321 252677 26333 253453
rect 26271 252665 26333 252677
rect 26389 253453 26451 253465
rect 26389 252677 26401 253453
rect 26435 252677 26451 253453
rect 26389 252665 26451 252677
rect 26481 253453 26543 253465
rect 26481 252677 26497 253453
rect 26531 252677 26543 253453
rect 26481 252665 26543 252677
rect 26599 253453 26661 253465
rect 26599 252677 26611 253453
rect 26645 252677 26661 253453
rect 26599 252665 26661 252677
rect 26691 253453 26753 253465
rect 26691 252677 26707 253453
rect 26741 252677 26753 253453
rect 26691 252665 26753 252677
rect 26809 253453 26871 253465
rect 26809 252677 26821 253453
rect 26855 252677 26871 253453
rect 26809 252665 26871 252677
rect 26901 253453 26963 253465
rect 26901 252677 26917 253453
rect 26951 252677 26963 253453
rect 26901 252665 26963 252677
rect 27019 253453 27081 253465
rect 27019 252677 27031 253453
rect 27065 252677 27081 253453
rect 27019 252665 27081 252677
rect 27111 253453 27173 253465
rect 27111 252677 27127 253453
rect 27161 252677 27173 253453
rect 27111 252665 27173 252677
rect 27229 253453 27291 253465
rect 27229 252677 27241 253453
rect 27275 252677 27291 253453
rect 27229 252665 27291 252677
rect 27321 253453 27383 253465
rect 27321 252677 27337 253453
rect 27371 252677 27383 253453
rect 27321 252665 27383 252677
rect -4061 252417 -3999 252429
rect -4061 251641 -4049 252417
rect -4015 251641 -3999 252417
rect -4061 251629 -3999 251641
rect -3969 252417 -3907 252429
rect -3969 251641 -3953 252417
rect -3919 251641 -3907 252417
rect -3969 251629 -3907 251641
rect -3851 252417 -3789 252429
rect -3851 251641 -3839 252417
rect -3805 251641 -3789 252417
rect -3851 251629 -3789 251641
rect -3759 252417 -3697 252429
rect -3759 251641 -3743 252417
rect -3709 251641 -3697 252417
rect -3759 251629 -3697 251641
rect -3641 252417 -3579 252429
rect -3641 251641 -3629 252417
rect -3595 251641 -3579 252417
rect -3641 251629 -3579 251641
rect -3549 252417 -3487 252429
rect -3549 251641 -3533 252417
rect -3499 251641 -3487 252417
rect -3549 251629 -3487 251641
rect -3431 252417 -3369 252429
rect -3431 251641 -3419 252417
rect -3385 251641 -3369 252417
rect -3431 251629 -3369 251641
rect -3339 252417 -3277 252429
rect -3339 251641 -3323 252417
rect -3289 251641 -3277 252417
rect -3339 251629 -3277 251641
rect -3221 252417 -3159 252429
rect -3221 251641 -3209 252417
rect -3175 251641 -3159 252417
rect -3221 251629 -3159 251641
rect -3129 252417 -3067 252429
rect -3129 251641 -3113 252417
rect -3079 251641 -3067 252417
rect -3129 251629 -3067 251641
rect -3011 252417 -2949 252429
rect -3011 251641 -2999 252417
rect -2965 251641 -2949 252417
rect -3011 251629 -2949 251641
rect -2919 252417 -2857 252429
rect -2919 251641 -2903 252417
rect -2869 251641 -2857 252417
rect -2919 251629 -2857 251641
rect -2801 252417 -2739 252429
rect -2801 251641 -2789 252417
rect -2755 251641 -2739 252417
rect -2801 251629 -2739 251641
rect -2709 252417 -2647 252429
rect -2709 251641 -2693 252417
rect -2659 251641 -2647 252417
rect -2709 251629 -2647 251641
rect -2591 252417 -2529 252429
rect -2591 251641 -2579 252417
rect -2545 251641 -2529 252417
rect -2591 251629 -2529 251641
rect -2499 252417 -2437 252429
rect -2499 251641 -2483 252417
rect -2449 251641 -2437 252417
rect -2499 251629 -2437 251641
rect -2381 252417 -2319 252429
rect -2381 251641 -2369 252417
rect -2335 251641 -2319 252417
rect -2381 251629 -2319 251641
rect -2289 252417 -2227 252429
rect -2289 251641 -2273 252417
rect -2239 251641 -2227 252417
rect -2289 251629 -2227 251641
rect -2171 252417 -2109 252429
rect -2171 251641 -2159 252417
rect -2125 251641 -2109 252417
rect -2171 251629 -2109 251641
rect -2079 252417 -2017 252429
rect -2079 251641 -2063 252417
rect -2029 251641 -2017 252417
rect -2079 251629 -2017 251641
rect -1961 252417 -1899 252429
rect -1961 251641 -1949 252417
rect -1915 251641 -1899 252417
rect -1961 251629 -1899 251641
rect -1869 252417 -1807 252429
rect -1869 251641 -1853 252417
rect -1819 251641 -1807 252417
rect -1869 251629 -1807 251641
rect -1751 252417 -1689 252429
rect -1751 251641 -1739 252417
rect -1705 251641 -1689 252417
rect -1751 251629 -1689 251641
rect -1659 252417 -1597 252429
rect -1659 251641 -1643 252417
rect -1609 251641 -1597 252417
rect -1659 251629 -1597 251641
rect -1541 252417 -1479 252429
rect -1541 251641 -1529 252417
rect -1495 251641 -1479 252417
rect -1541 251629 -1479 251641
rect -1449 252417 -1387 252429
rect -1449 251641 -1433 252417
rect -1399 251641 -1387 252417
rect -1449 251629 -1387 251641
rect -1331 252417 -1269 252429
rect -1331 251641 -1319 252417
rect -1285 251641 -1269 252417
rect -1331 251629 -1269 251641
rect -1239 252417 -1177 252429
rect -1239 251641 -1223 252417
rect -1189 251641 -1177 252417
rect -1239 251629 -1177 251641
rect -1121 252417 -1059 252429
rect -1121 251641 -1109 252417
rect -1075 251641 -1059 252417
rect -1121 251629 -1059 251641
rect -1029 252417 -967 252429
rect -1029 251641 -1013 252417
rect -979 251641 -967 252417
rect -1029 251629 -967 251641
rect -911 252417 -849 252429
rect -911 251641 -899 252417
rect -865 251641 -849 252417
rect -911 251629 -849 251641
rect -819 252417 -757 252429
rect -819 251641 -803 252417
rect -769 251641 -757 252417
rect -819 251629 -757 251641
rect -701 252417 -639 252429
rect -701 251641 -689 252417
rect -655 251641 -639 252417
rect -701 251629 -639 251641
rect -609 252417 -547 252429
rect -609 251641 -593 252417
rect -559 251641 -547 252417
rect -609 251629 -547 251641
rect -491 252417 -429 252429
rect -491 251641 -479 252417
rect -445 251641 -429 252417
rect -491 251629 -429 251641
rect -399 252417 -337 252429
rect -399 251641 -383 252417
rect -349 251641 -337 252417
rect -399 251629 -337 251641
rect -281 252417 -219 252429
rect -281 251641 -269 252417
rect -235 251641 -219 252417
rect -281 251629 -219 251641
rect -189 252417 -127 252429
rect -189 251641 -173 252417
rect -139 251641 -127 252417
rect -189 251629 -127 251641
rect -71 252417 -9 252429
rect -71 251641 -59 252417
rect -25 251641 -9 252417
rect -71 251629 -9 251641
rect 21 252417 83 252429
rect 21 251641 37 252417
rect 71 251641 83 252417
rect 21 251629 83 251641
rect 139 252417 201 252429
rect 139 251641 151 252417
rect 185 251641 201 252417
rect 139 251629 201 251641
rect 231 252417 293 252429
rect 231 251641 247 252417
rect 281 251641 293 252417
rect 231 251629 293 251641
rect 349 252417 411 252429
rect 349 251641 361 252417
rect 395 251641 411 252417
rect 349 251629 411 251641
rect 441 252417 503 252429
rect 441 251641 457 252417
rect 491 251641 503 252417
rect 441 251629 503 251641
rect 559 252417 621 252429
rect 559 251641 571 252417
rect 605 251641 621 252417
rect 559 251629 621 251641
rect 651 252417 713 252429
rect 651 251641 667 252417
rect 701 251641 713 252417
rect 651 251629 713 251641
rect 769 252417 831 252429
rect 769 251641 781 252417
rect 815 251641 831 252417
rect 769 251629 831 251641
rect 861 252417 923 252429
rect 861 251641 877 252417
rect 911 251641 923 252417
rect 861 251629 923 251641
rect 979 252417 1041 252429
rect 979 251641 991 252417
rect 1025 251641 1041 252417
rect 979 251629 1041 251641
rect 1071 252417 1133 252429
rect 1071 251641 1087 252417
rect 1121 251641 1133 252417
rect 1071 251629 1133 251641
rect 1189 252417 1251 252429
rect 1189 251641 1201 252417
rect 1235 251641 1251 252417
rect 1189 251629 1251 251641
rect 1281 252417 1343 252429
rect 1281 251641 1297 252417
rect 1331 251641 1343 252417
rect 1281 251629 1343 251641
rect 1399 252417 1461 252429
rect 1399 251641 1411 252417
rect 1445 251641 1461 252417
rect 1399 251629 1461 251641
rect 1491 252417 1553 252429
rect 1491 251641 1507 252417
rect 1541 251641 1553 252417
rect 1491 251629 1553 251641
rect 1609 252417 1671 252429
rect 1609 251641 1621 252417
rect 1655 251641 1671 252417
rect 1609 251629 1671 251641
rect 1701 252417 1763 252429
rect 1701 251641 1717 252417
rect 1751 251641 1763 252417
rect 1701 251629 1763 251641
rect 1819 252417 1881 252429
rect 1819 251641 1831 252417
rect 1865 251641 1881 252417
rect 1819 251629 1881 251641
rect 1911 252417 1973 252429
rect 1911 251641 1927 252417
rect 1961 251641 1973 252417
rect 1911 251629 1973 251641
rect 2029 252417 2091 252429
rect 2029 251641 2041 252417
rect 2075 251641 2091 252417
rect 2029 251629 2091 251641
rect 2121 252417 2183 252429
rect 2121 251641 2137 252417
rect 2171 251641 2183 252417
rect 2121 251629 2183 251641
rect 2239 252417 2301 252429
rect 2239 251641 2251 252417
rect 2285 251641 2301 252417
rect 2239 251629 2301 251641
rect 2331 252417 2393 252429
rect 2331 251641 2347 252417
rect 2381 251641 2393 252417
rect 2331 251629 2393 251641
rect 2449 252417 2511 252429
rect 2449 251641 2461 252417
rect 2495 251641 2511 252417
rect 2449 251629 2511 251641
rect 2541 252417 2603 252429
rect 2541 251641 2557 252417
rect 2591 251641 2603 252417
rect 2541 251629 2603 251641
rect 2659 252417 2721 252429
rect 2659 251641 2671 252417
rect 2705 251641 2721 252417
rect 2659 251629 2721 251641
rect 2751 252417 2813 252429
rect 2751 251641 2767 252417
rect 2801 251641 2813 252417
rect 2751 251629 2813 251641
rect 2869 252417 2931 252429
rect 2869 251641 2881 252417
rect 2915 251641 2931 252417
rect 2869 251629 2931 251641
rect 2961 252417 3023 252429
rect 2961 251641 2977 252417
rect 3011 251641 3023 252417
rect 2961 251629 3023 251641
rect 3079 252417 3141 252429
rect 3079 251641 3091 252417
rect 3125 251641 3141 252417
rect 3079 251629 3141 251641
rect 3171 252417 3233 252429
rect 3171 251641 3187 252417
rect 3221 251641 3233 252417
rect 3171 251629 3233 251641
rect 3289 252417 3351 252429
rect 3289 251641 3301 252417
rect 3335 251641 3351 252417
rect 3289 251629 3351 251641
rect 3381 252417 3443 252429
rect 3381 251641 3397 252417
rect 3431 251641 3443 252417
rect 3381 251629 3443 251641
rect 3499 252417 3561 252429
rect 3499 251641 3511 252417
rect 3545 251641 3561 252417
rect 3499 251629 3561 251641
rect 3591 252417 3653 252429
rect 3591 251641 3607 252417
rect 3641 251641 3653 252417
rect 3591 251629 3653 251641
rect 3709 252417 3771 252429
rect 3709 251641 3721 252417
rect 3755 251641 3771 252417
rect 3709 251629 3771 251641
rect 3801 252417 3863 252429
rect 3801 251641 3817 252417
rect 3851 251641 3863 252417
rect 3801 251629 3863 251641
rect 3919 252417 3981 252429
rect 3919 251641 3931 252417
rect 3965 251641 3981 252417
rect 3919 251629 3981 251641
rect 4011 252417 4073 252429
rect 4011 251641 4027 252417
rect 4061 251641 4073 252417
rect 4011 251629 4073 251641
rect 4129 252417 4191 252429
rect 4129 251641 4141 252417
rect 4175 251641 4191 252417
rect 4129 251629 4191 251641
rect 4221 252417 4283 252429
rect 4221 251641 4237 252417
rect 4271 251641 4283 252417
rect 4221 251629 4283 251641
rect 4339 252417 4401 252429
rect 4339 251641 4351 252417
rect 4385 251641 4401 252417
rect 4339 251629 4401 251641
rect 4431 252417 4493 252429
rect 4431 251641 4447 252417
rect 4481 251641 4493 252417
rect 4431 251629 4493 251641
rect 4549 252417 4611 252429
rect 4549 251641 4561 252417
rect 4595 251641 4611 252417
rect 4549 251629 4611 251641
rect 4641 252417 4703 252429
rect 4641 251641 4657 252417
rect 4691 251641 4703 252417
rect 4641 251629 4703 251641
rect 4759 252417 4821 252429
rect 4759 251641 4771 252417
rect 4805 251641 4821 252417
rect 4759 251629 4821 251641
rect 4851 252417 4913 252429
rect 4851 251641 4867 252417
rect 4901 251641 4913 252417
rect 4851 251629 4913 251641
rect 4969 252417 5031 252429
rect 4969 251641 4981 252417
rect 5015 251641 5031 252417
rect 4969 251629 5031 251641
rect 5061 252417 5123 252429
rect 5061 251641 5077 252417
rect 5111 251641 5123 252417
rect 5061 251629 5123 251641
rect 5179 252417 5241 252429
rect 5179 251641 5191 252417
rect 5225 251641 5241 252417
rect 5179 251629 5241 251641
rect 5271 252417 5333 252429
rect 5271 251641 5287 252417
rect 5321 251641 5333 252417
rect 5271 251629 5333 251641
rect 5389 252417 5451 252429
rect 5389 251641 5401 252417
rect 5435 251641 5451 252417
rect 5389 251629 5451 251641
rect 5481 252417 5543 252429
rect 5481 251641 5497 252417
rect 5531 251641 5543 252417
rect 5481 251629 5543 251641
rect 5599 252417 5661 252429
rect 5599 251641 5611 252417
rect 5645 251641 5661 252417
rect 5599 251629 5661 251641
rect 5691 252417 5753 252429
rect 5691 251641 5707 252417
rect 5741 251641 5753 252417
rect 5691 251629 5753 251641
rect 5809 252417 5871 252429
rect 5809 251641 5821 252417
rect 5855 251641 5871 252417
rect 5809 251629 5871 251641
rect 5901 252417 5963 252429
rect 5901 251641 5917 252417
rect 5951 251641 5963 252417
rect 5901 251629 5963 251641
rect 6019 252417 6081 252429
rect 6019 251641 6031 252417
rect 6065 251641 6081 252417
rect 6019 251629 6081 251641
rect 6111 252417 6173 252429
rect 6111 251641 6127 252417
rect 6161 251641 6173 252417
rect 6111 251629 6173 251641
rect 6229 252417 6291 252429
rect 6229 251641 6241 252417
rect 6275 251641 6291 252417
rect 6229 251629 6291 251641
rect 6321 252417 6383 252429
rect 6321 251641 6337 252417
rect 6371 251641 6383 252417
rect 6321 251629 6383 251641
rect 6439 252417 6501 252429
rect 6439 251641 6451 252417
rect 6485 251641 6501 252417
rect 6439 251629 6501 251641
rect 6531 252417 6593 252429
rect 6531 251641 6547 252417
rect 6581 251641 6593 252417
rect 6531 251629 6593 251641
rect 6649 252417 6711 252429
rect 6649 251641 6661 252417
rect 6695 251641 6711 252417
rect 6649 251629 6711 251641
rect 6741 252417 6803 252429
rect 6741 251641 6757 252417
rect 6791 251641 6803 252417
rect 6741 251629 6803 251641
rect 6859 252417 6921 252429
rect 6859 251641 6871 252417
rect 6905 251641 6921 252417
rect 6859 251629 6921 251641
rect 6951 252417 7013 252429
rect 6951 251641 6967 252417
rect 7001 251641 7013 252417
rect 6951 251629 7013 251641
rect 7069 252417 7131 252429
rect 7069 251641 7081 252417
rect 7115 251641 7131 252417
rect 7069 251629 7131 251641
rect 7161 252417 7223 252429
rect 7161 251641 7177 252417
rect 7211 251641 7223 252417
rect 7161 251629 7223 251641
rect 7279 252417 7341 252429
rect 7279 251641 7291 252417
rect 7325 251641 7341 252417
rect 7279 251629 7341 251641
rect 7371 252417 7433 252429
rect 7371 251641 7387 252417
rect 7421 251641 7433 252417
rect 7371 251629 7433 251641
rect 7489 252417 7551 252429
rect 7489 251641 7501 252417
rect 7535 251641 7551 252417
rect 7489 251629 7551 251641
rect 7581 252417 7643 252429
rect 7581 251641 7597 252417
rect 7631 251641 7643 252417
rect 7581 251629 7643 251641
rect 7699 252417 7761 252429
rect 7699 251641 7711 252417
rect 7745 251641 7761 252417
rect 7699 251629 7761 251641
rect 7791 252417 7853 252429
rect 7791 251641 7807 252417
rect 7841 251641 7853 252417
rect 7791 251629 7853 251641
rect 7909 252417 7971 252429
rect 7909 251641 7921 252417
rect 7955 251641 7971 252417
rect 7909 251629 7971 251641
rect 8001 252417 8063 252429
rect 8001 251641 8017 252417
rect 8051 251641 8063 252417
rect 8001 251629 8063 251641
rect 8119 252417 8181 252429
rect 8119 251641 8131 252417
rect 8165 251641 8181 252417
rect 8119 251629 8181 251641
rect 8211 252417 8273 252429
rect 8211 251641 8227 252417
rect 8261 251641 8273 252417
rect 8211 251629 8273 251641
rect 8329 252417 8391 252429
rect 8329 251641 8341 252417
rect 8375 251641 8391 252417
rect 8329 251629 8391 251641
rect 8421 252417 8483 252429
rect 8421 251641 8437 252417
rect 8471 251641 8483 252417
rect 8421 251629 8483 251641
rect 8539 252417 8601 252429
rect 8539 251641 8551 252417
rect 8585 251641 8601 252417
rect 8539 251629 8601 251641
rect 8631 252417 8693 252429
rect 8631 251641 8647 252417
rect 8681 251641 8693 252417
rect 8631 251629 8693 251641
rect 8749 252417 8811 252429
rect 8749 251641 8761 252417
rect 8795 251641 8811 252417
rect 8749 251629 8811 251641
rect 8841 252417 8903 252429
rect 8841 251641 8857 252417
rect 8891 251641 8903 252417
rect 8841 251629 8903 251641
rect 8959 252417 9021 252429
rect 8959 251641 8971 252417
rect 9005 251641 9021 252417
rect 8959 251629 9021 251641
rect 9051 252417 9113 252429
rect 9051 251641 9067 252417
rect 9101 251641 9113 252417
rect 9051 251629 9113 251641
rect 9169 252417 9231 252429
rect 9169 251641 9181 252417
rect 9215 251641 9231 252417
rect 9169 251629 9231 251641
rect 9261 252417 9323 252429
rect 9261 251641 9277 252417
rect 9311 251641 9323 252417
rect 9261 251629 9323 251641
rect 9379 252417 9441 252429
rect 9379 251641 9391 252417
rect 9425 251641 9441 252417
rect 9379 251629 9441 251641
rect 9471 252417 9533 252429
rect 9471 251641 9487 252417
rect 9521 251641 9533 252417
rect 9471 251629 9533 251641
rect 9589 252417 9651 252429
rect 9589 251641 9601 252417
rect 9635 251641 9651 252417
rect 9589 251629 9651 251641
rect 9681 252417 9743 252429
rect 9681 251641 9697 252417
rect 9731 251641 9743 252417
rect 9681 251629 9743 251641
rect 9799 252417 9861 252429
rect 9799 251641 9811 252417
rect 9845 251641 9861 252417
rect 9799 251629 9861 251641
rect 9891 252417 9953 252429
rect 9891 251641 9907 252417
rect 9941 251641 9953 252417
rect 9891 251629 9953 251641
rect 10009 252417 10071 252429
rect 10009 251641 10021 252417
rect 10055 251641 10071 252417
rect 10009 251629 10071 251641
rect 10101 252417 10163 252429
rect 10101 251641 10117 252417
rect 10151 251641 10163 252417
rect 10101 251629 10163 251641
rect 10219 252417 10281 252429
rect 10219 251641 10231 252417
rect 10265 251641 10281 252417
rect 10219 251629 10281 251641
rect 10311 252417 10373 252429
rect 10311 251641 10327 252417
rect 10361 251641 10373 252417
rect 10311 251629 10373 251641
rect 10429 252417 10491 252429
rect 10429 251641 10441 252417
rect 10475 251641 10491 252417
rect 10429 251629 10491 251641
rect 10521 252417 10583 252429
rect 10521 251641 10537 252417
rect 10571 251641 10583 252417
rect 10521 251629 10583 251641
rect 10639 252417 10701 252429
rect 10639 251641 10651 252417
rect 10685 251641 10701 252417
rect 10639 251629 10701 251641
rect 10731 252417 10793 252429
rect 10731 251641 10747 252417
rect 10781 251641 10793 252417
rect 10731 251629 10793 251641
rect 10849 252417 10911 252429
rect 10849 251641 10861 252417
rect 10895 251641 10911 252417
rect 10849 251629 10911 251641
rect 10941 252417 11003 252429
rect 10941 251641 10957 252417
rect 10991 251641 11003 252417
rect 10941 251629 11003 251641
rect 11059 252417 11121 252429
rect 11059 251641 11071 252417
rect 11105 251641 11121 252417
rect 11059 251629 11121 251641
rect 11151 252417 11213 252429
rect 11151 251641 11167 252417
rect 11201 251641 11213 252417
rect 11151 251629 11213 251641
rect 11269 252417 11331 252429
rect 11269 251641 11281 252417
rect 11315 251641 11331 252417
rect 11269 251629 11331 251641
rect 11361 252417 11423 252429
rect 11361 251641 11377 252417
rect 11411 251641 11423 252417
rect 11361 251629 11423 251641
rect 11479 252417 11541 252429
rect 11479 251641 11491 252417
rect 11525 251641 11541 252417
rect 11479 251629 11541 251641
rect 11571 252417 11633 252429
rect 11571 251641 11587 252417
rect 11621 251641 11633 252417
rect 11571 251629 11633 251641
rect 11689 252417 11751 252429
rect 11689 251641 11701 252417
rect 11735 251641 11751 252417
rect 11689 251629 11751 251641
rect 11781 252417 11843 252429
rect 11781 251641 11797 252417
rect 11831 251641 11843 252417
rect 11781 251629 11843 251641
rect 11899 252417 11961 252429
rect 11899 251641 11911 252417
rect 11945 251641 11961 252417
rect 11899 251629 11961 251641
rect 11991 252417 12053 252429
rect 11991 251641 12007 252417
rect 12041 251641 12053 252417
rect 11991 251629 12053 251641
rect 12109 252417 12171 252429
rect 12109 251641 12121 252417
rect 12155 251641 12171 252417
rect 12109 251629 12171 251641
rect 12201 252417 12263 252429
rect 12201 251641 12217 252417
rect 12251 251641 12263 252417
rect 12201 251629 12263 251641
rect 12319 252417 12381 252429
rect 12319 251641 12331 252417
rect 12365 251641 12381 252417
rect 12319 251629 12381 251641
rect 12411 252417 12473 252429
rect 12411 251641 12427 252417
rect 12461 251641 12473 252417
rect 12411 251629 12473 251641
rect 12529 252417 12591 252429
rect 12529 251641 12541 252417
rect 12575 251641 12591 252417
rect 12529 251629 12591 251641
rect 12621 252417 12683 252429
rect 12621 251641 12637 252417
rect 12671 251641 12683 252417
rect 12621 251629 12683 251641
rect 12739 252417 12801 252429
rect 12739 251641 12751 252417
rect 12785 251641 12801 252417
rect 12739 251629 12801 251641
rect 12831 252417 12893 252429
rect 12831 251641 12847 252417
rect 12881 251641 12893 252417
rect 12831 251629 12893 251641
rect 12949 252417 13011 252429
rect 12949 251641 12961 252417
rect 12995 251641 13011 252417
rect 12949 251629 13011 251641
rect 13041 252417 13103 252429
rect 13041 251641 13057 252417
rect 13091 251641 13103 252417
rect 13041 251629 13103 251641
rect 13159 252417 13221 252429
rect 13159 251641 13171 252417
rect 13205 251641 13221 252417
rect 13159 251629 13221 251641
rect 13251 252417 13313 252429
rect 13251 251641 13267 252417
rect 13301 251641 13313 252417
rect 13251 251629 13313 251641
rect 13369 252417 13431 252429
rect 13369 251641 13381 252417
rect 13415 251641 13431 252417
rect 13369 251629 13431 251641
rect 13461 252417 13523 252429
rect 13461 251641 13477 252417
rect 13511 251641 13523 252417
rect 13461 251629 13523 251641
rect 13579 252417 13641 252429
rect 13579 251641 13591 252417
rect 13625 251641 13641 252417
rect 13579 251629 13641 251641
rect 13671 252417 13733 252429
rect 13671 251641 13687 252417
rect 13721 251641 13733 252417
rect 13671 251629 13733 251641
rect 13789 252417 13851 252429
rect 13789 251641 13801 252417
rect 13835 251641 13851 252417
rect 13789 251629 13851 251641
rect 13881 252417 13943 252429
rect 13881 251641 13897 252417
rect 13931 251641 13943 252417
rect 13881 251629 13943 251641
rect 13999 252417 14061 252429
rect 13999 251641 14011 252417
rect 14045 251641 14061 252417
rect 13999 251629 14061 251641
rect 14091 252417 14153 252429
rect 14091 251641 14107 252417
rect 14141 251641 14153 252417
rect 14091 251629 14153 251641
rect 14209 252417 14271 252429
rect 14209 251641 14221 252417
rect 14255 251641 14271 252417
rect 14209 251629 14271 251641
rect 14301 252417 14363 252429
rect 14301 251641 14317 252417
rect 14351 251641 14363 252417
rect 14301 251629 14363 251641
rect 14419 252417 14481 252429
rect 14419 251641 14431 252417
rect 14465 251641 14481 252417
rect 14419 251629 14481 251641
rect 14511 252417 14573 252429
rect 14511 251641 14527 252417
rect 14561 251641 14573 252417
rect 14511 251629 14573 251641
rect 14629 252417 14691 252429
rect 14629 251641 14641 252417
rect 14675 251641 14691 252417
rect 14629 251629 14691 251641
rect 14721 252417 14783 252429
rect 14721 251641 14737 252417
rect 14771 251641 14783 252417
rect 14721 251629 14783 251641
rect 14839 252417 14901 252429
rect 14839 251641 14851 252417
rect 14885 251641 14901 252417
rect 14839 251629 14901 251641
rect 14931 252417 14993 252429
rect 14931 251641 14947 252417
rect 14981 251641 14993 252417
rect 14931 251629 14993 251641
rect 15049 252417 15111 252429
rect 15049 251641 15061 252417
rect 15095 251641 15111 252417
rect 15049 251629 15111 251641
rect 15141 252417 15203 252429
rect 15141 251641 15157 252417
rect 15191 251641 15203 252417
rect 15141 251629 15203 251641
rect 15259 252417 15321 252429
rect 15259 251641 15271 252417
rect 15305 251641 15321 252417
rect 15259 251629 15321 251641
rect 15351 252417 15413 252429
rect 15351 251641 15367 252417
rect 15401 251641 15413 252417
rect 15351 251629 15413 251641
rect 15469 252417 15531 252429
rect 15469 251641 15481 252417
rect 15515 251641 15531 252417
rect 15469 251629 15531 251641
rect 15561 252417 15623 252429
rect 15561 251641 15577 252417
rect 15611 251641 15623 252417
rect 15561 251629 15623 251641
rect 15679 252417 15741 252429
rect 15679 251641 15691 252417
rect 15725 251641 15741 252417
rect 15679 251629 15741 251641
rect 15771 252417 15833 252429
rect 15771 251641 15787 252417
rect 15821 251641 15833 252417
rect 15771 251629 15833 251641
rect 15889 252417 15951 252429
rect 15889 251641 15901 252417
rect 15935 251641 15951 252417
rect 15889 251629 15951 251641
rect 15981 252417 16043 252429
rect 15981 251641 15997 252417
rect 16031 251641 16043 252417
rect 15981 251629 16043 251641
rect 16099 252417 16161 252429
rect 16099 251641 16111 252417
rect 16145 251641 16161 252417
rect 16099 251629 16161 251641
rect 16191 252417 16253 252429
rect 16191 251641 16207 252417
rect 16241 251641 16253 252417
rect 16191 251629 16253 251641
rect 16309 252417 16371 252429
rect 16309 251641 16321 252417
rect 16355 251641 16371 252417
rect 16309 251629 16371 251641
rect 16401 252417 16463 252429
rect 16401 251641 16417 252417
rect 16451 251641 16463 252417
rect 16401 251629 16463 251641
rect 16519 252417 16581 252429
rect 16519 251641 16531 252417
rect 16565 251641 16581 252417
rect 16519 251629 16581 251641
rect 16611 252417 16673 252429
rect 16611 251641 16627 252417
rect 16661 251641 16673 252417
rect 16611 251629 16673 251641
rect 16729 252417 16791 252429
rect 16729 251641 16741 252417
rect 16775 251641 16791 252417
rect 16729 251629 16791 251641
rect 16821 252417 16883 252429
rect 16821 251641 16837 252417
rect 16871 251641 16883 252417
rect 16821 251629 16883 251641
rect 16939 252417 17001 252429
rect 16939 251641 16951 252417
rect 16985 251641 17001 252417
rect 16939 251629 17001 251641
rect 17031 252417 17093 252429
rect 17031 251641 17047 252417
rect 17081 251641 17093 252417
rect 17031 251629 17093 251641
rect 17149 252417 17211 252429
rect 17149 251641 17161 252417
rect 17195 251641 17211 252417
rect 17149 251629 17211 251641
rect 17241 252417 17303 252429
rect 17241 251641 17257 252417
rect 17291 251641 17303 252417
rect 17241 251629 17303 251641
rect 17359 252417 17421 252429
rect 17359 251641 17371 252417
rect 17405 251641 17421 252417
rect 17359 251629 17421 251641
rect 17451 252417 17513 252429
rect 17451 251641 17467 252417
rect 17501 251641 17513 252417
rect 17451 251629 17513 251641
rect 17569 252417 17631 252429
rect 17569 251641 17581 252417
rect 17615 251641 17631 252417
rect 17569 251629 17631 251641
rect 17661 252417 17723 252429
rect 17661 251641 17677 252417
rect 17711 251641 17723 252417
rect 17661 251629 17723 251641
rect 17779 252417 17841 252429
rect 17779 251641 17791 252417
rect 17825 251641 17841 252417
rect 17779 251629 17841 251641
rect 17871 252417 17933 252429
rect 17871 251641 17887 252417
rect 17921 251641 17933 252417
rect 17871 251629 17933 251641
rect 17989 252417 18051 252429
rect 17989 251641 18001 252417
rect 18035 251641 18051 252417
rect 17989 251629 18051 251641
rect 18081 252417 18143 252429
rect 18081 251641 18097 252417
rect 18131 251641 18143 252417
rect 18081 251629 18143 251641
rect 18199 252417 18261 252429
rect 18199 251641 18211 252417
rect 18245 251641 18261 252417
rect 18199 251629 18261 251641
rect 18291 252417 18353 252429
rect 18291 251641 18307 252417
rect 18341 251641 18353 252417
rect 18291 251629 18353 251641
rect 18409 252417 18471 252429
rect 18409 251641 18421 252417
rect 18455 251641 18471 252417
rect 18409 251629 18471 251641
rect 18501 252417 18563 252429
rect 18501 251641 18517 252417
rect 18551 251641 18563 252417
rect 18501 251629 18563 251641
rect 18619 252417 18681 252429
rect 18619 251641 18631 252417
rect 18665 251641 18681 252417
rect 18619 251629 18681 251641
rect 18711 252417 18773 252429
rect 18711 251641 18727 252417
rect 18761 251641 18773 252417
rect 18711 251629 18773 251641
rect 18829 252417 18891 252429
rect 18829 251641 18841 252417
rect 18875 251641 18891 252417
rect 18829 251629 18891 251641
rect 18921 252417 18983 252429
rect 18921 251641 18937 252417
rect 18971 251641 18983 252417
rect 18921 251629 18983 251641
rect 19039 252417 19101 252429
rect 19039 251641 19051 252417
rect 19085 251641 19101 252417
rect 19039 251629 19101 251641
rect 19131 252417 19193 252429
rect 19131 251641 19147 252417
rect 19181 251641 19193 252417
rect 19131 251629 19193 251641
rect 19249 252417 19311 252429
rect 19249 251641 19261 252417
rect 19295 251641 19311 252417
rect 19249 251629 19311 251641
rect 19341 252417 19403 252429
rect 19341 251641 19357 252417
rect 19391 251641 19403 252417
rect 19341 251629 19403 251641
rect 19459 252417 19521 252429
rect 19459 251641 19471 252417
rect 19505 251641 19521 252417
rect 19459 251629 19521 251641
rect 19551 252417 19613 252429
rect 19551 251641 19567 252417
rect 19601 251641 19613 252417
rect 19551 251629 19613 251641
rect 19669 252417 19731 252429
rect 19669 251641 19681 252417
rect 19715 251641 19731 252417
rect 19669 251629 19731 251641
rect 19761 252417 19823 252429
rect 19761 251641 19777 252417
rect 19811 251641 19823 252417
rect 19761 251629 19823 251641
rect 19879 252417 19941 252429
rect 19879 251641 19891 252417
rect 19925 251641 19941 252417
rect 19879 251629 19941 251641
rect 19971 252417 20033 252429
rect 19971 251641 19987 252417
rect 20021 251641 20033 252417
rect 19971 251629 20033 251641
rect 20089 252417 20151 252429
rect 20089 251641 20101 252417
rect 20135 251641 20151 252417
rect 20089 251629 20151 251641
rect 20181 252417 20243 252429
rect 20181 251641 20197 252417
rect 20231 251641 20243 252417
rect 20181 251629 20243 251641
rect 20299 252417 20361 252429
rect 20299 251641 20311 252417
rect 20345 251641 20361 252417
rect 20299 251629 20361 251641
rect 20391 252417 20453 252429
rect 20391 251641 20407 252417
rect 20441 251641 20453 252417
rect 20391 251629 20453 251641
rect 20509 252417 20571 252429
rect 20509 251641 20521 252417
rect 20555 251641 20571 252417
rect 20509 251629 20571 251641
rect 20601 252417 20663 252429
rect 20601 251641 20617 252417
rect 20651 251641 20663 252417
rect 20601 251629 20663 251641
rect 20719 252417 20781 252429
rect 20719 251641 20731 252417
rect 20765 251641 20781 252417
rect 20719 251629 20781 251641
rect 20811 252417 20873 252429
rect 20811 251641 20827 252417
rect 20861 251641 20873 252417
rect 20811 251629 20873 251641
rect 20929 252417 20991 252429
rect 20929 251641 20941 252417
rect 20975 251641 20991 252417
rect 20929 251629 20991 251641
rect 21021 252417 21083 252429
rect 21021 251641 21037 252417
rect 21071 251641 21083 252417
rect 21021 251629 21083 251641
rect 21139 252417 21201 252429
rect 21139 251641 21151 252417
rect 21185 251641 21201 252417
rect 21139 251629 21201 251641
rect 21231 252417 21293 252429
rect 21231 251641 21247 252417
rect 21281 251641 21293 252417
rect 21231 251629 21293 251641
rect 21349 252417 21411 252429
rect 21349 251641 21361 252417
rect 21395 251641 21411 252417
rect 21349 251629 21411 251641
rect 21441 252417 21503 252429
rect 21441 251641 21457 252417
rect 21491 251641 21503 252417
rect 21441 251629 21503 251641
rect 21559 252417 21621 252429
rect 21559 251641 21571 252417
rect 21605 251641 21621 252417
rect 21559 251629 21621 251641
rect 21651 252417 21713 252429
rect 21651 251641 21667 252417
rect 21701 251641 21713 252417
rect 21651 251629 21713 251641
rect 21769 252417 21831 252429
rect 21769 251641 21781 252417
rect 21815 251641 21831 252417
rect 21769 251629 21831 251641
rect 21861 252417 21923 252429
rect 21861 251641 21877 252417
rect 21911 251641 21923 252417
rect 21861 251629 21923 251641
rect 21979 252417 22041 252429
rect 21979 251641 21991 252417
rect 22025 251641 22041 252417
rect 21979 251629 22041 251641
rect 22071 252417 22133 252429
rect 22071 251641 22087 252417
rect 22121 251641 22133 252417
rect 22071 251629 22133 251641
rect 22189 252417 22251 252429
rect 22189 251641 22201 252417
rect 22235 251641 22251 252417
rect 22189 251629 22251 251641
rect 22281 252417 22343 252429
rect 22281 251641 22297 252417
rect 22331 251641 22343 252417
rect 22281 251629 22343 251641
rect 22399 252417 22461 252429
rect 22399 251641 22411 252417
rect 22445 251641 22461 252417
rect 22399 251629 22461 251641
rect 22491 252417 22553 252429
rect 22491 251641 22507 252417
rect 22541 251641 22553 252417
rect 22491 251629 22553 251641
rect 22609 252417 22671 252429
rect 22609 251641 22621 252417
rect 22655 251641 22671 252417
rect 22609 251629 22671 251641
rect 22701 252417 22763 252429
rect 22701 251641 22717 252417
rect 22751 251641 22763 252417
rect 22701 251629 22763 251641
rect 22819 252417 22881 252429
rect 22819 251641 22831 252417
rect 22865 251641 22881 252417
rect 22819 251629 22881 251641
rect 22911 252417 22973 252429
rect 22911 251641 22927 252417
rect 22961 251641 22973 252417
rect 22911 251629 22973 251641
rect 23029 252417 23091 252429
rect 23029 251641 23041 252417
rect 23075 251641 23091 252417
rect 23029 251629 23091 251641
rect 23121 252417 23183 252429
rect 23121 251641 23137 252417
rect 23171 251641 23183 252417
rect 23121 251629 23183 251641
rect 23239 252417 23301 252429
rect 23239 251641 23251 252417
rect 23285 251641 23301 252417
rect 23239 251629 23301 251641
rect 23331 252417 23393 252429
rect 23331 251641 23347 252417
rect 23381 251641 23393 252417
rect 23331 251629 23393 251641
rect 23449 252417 23511 252429
rect 23449 251641 23461 252417
rect 23495 251641 23511 252417
rect 23449 251629 23511 251641
rect 23541 252417 23603 252429
rect 23541 251641 23557 252417
rect 23591 251641 23603 252417
rect 23541 251629 23603 251641
rect 23659 252417 23721 252429
rect 23659 251641 23671 252417
rect 23705 251641 23721 252417
rect 23659 251629 23721 251641
rect 23751 252417 23813 252429
rect 23751 251641 23767 252417
rect 23801 251641 23813 252417
rect 23751 251629 23813 251641
rect 23869 252417 23931 252429
rect 23869 251641 23881 252417
rect 23915 251641 23931 252417
rect 23869 251629 23931 251641
rect 23961 252417 24023 252429
rect 23961 251641 23977 252417
rect 24011 251641 24023 252417
rect 23961 251629 24023 251641
rect 24079 252417 24141 252429
rect 24079 251641 24091 252417
rect 24125 251641 24141 252417
rect 24079 251629 24141 251641
rect 24171 252417 24233 252429
rect 24171 251641 24187 252417
rect 24221 251641 24233 252417
rect 24171 251629 24233 251641
rect 24289 252417 24351 252429
rect 24289 251641 24301 252417
rect 24335 251641 24351 252417
rect 24289 251629 24351 251641
rect 24381 252417 24443 252429
rect 24381 251641 24397 252417
rect 24431 251641 24443 252417
rect 24381 251629 24443 251641
rect 24499 252417 24561 252429
rect 24499 251641 24511 252417
rect 24545 251641 24561 252417
rect 24499 251629 24561 251641
rect 24591 252417 24653 252429
rect 24591 251641 24607 252417
rect 24641 251641 24653 252417
rect 24591 251629 24653 251641
rect 24709 252417 24771 252429
rect 24709 251641 24721 252417
rect 24755 251641 24771 252417
rect 24709 251629 24771 251641
rect 24801 252417 24863 252429
rect 24801 251641 24817 252417
rect 24851 251641 24863 252417
rect 24801 251629 24863 251641
rect 24919 252417 24981 252429
rect 24919 251641 24931 252417
rect 24965 251641 24981 252417
rect 24919 251629 24981 251641
rect 25011 252417 25073 252429
rect 25011 251641 25027 252417
rect 25061 251641 25073 252417
rect 25011 251629 25073 251641
rect 25129 252417 25191 252429
rect 25129 251641 25141 252417
rect 25175 251641 25191 252417
rect 25129 251629 25191 251641
rect 25221 252417 25283 252429
rect 25221 251641 25237 252417
rect 25271 251641 25283 252417
rect 25221 251629 25283 251641
rect 25339 252417 25401 252429
rect 25339 251641 25351 252417
rect 25385 251641 25401 252417
rect 25339 251629 25401 251641
rect 25431 252417 25493 252429
rect 25431 251641 25447 252417
rect 25481 251641 25493 252417
rect 25431 251629 25493 251641
rect 25549 252417 25611 252429
rect 25549 251641 25561 252417
rect 25595 251641 25611 252417
rect 25549 251629 25611 251641
rect 25641 252417 25703 252429
rect 25641 251641 25657 252417
rect 25691 251641 25703 252417
rect 25641 251629 25703 251641
rect 25759 252417 25821 252429
rect 25759 251641 25771 252417
rect 25805 251641 25821 252417
rect 25759 251629 25821 251641
rect 25851 252417 25913 252429
rect 25851 251641 25867 252417
rect 25901 251641 25913 252417
rect 25851 251629 25913 251641
rect 25969 252417 26031 252429
rect 25969 251641 25981 252417
rect 26015 251641 26031 252417
rect 25969 251629 26031 251641
rect 26061 252417 26123 252429
rect 26061 251641 26077 252417
rect 26111 251641 26123 252417
rect 26061 251629 26123 251641
rect 26179 252417 26241 252429
rect 26179 251641 26191 252417
rect 26225 251641 26241 252417
rect 26179 251629 26241 251641
rect 26271 252417 26333 252429
rect 26271 251641 26287 252417
rect 26321 251641 26333 252417
rect 26271 251629 26333 251641
rect 26389 252417 26451 252429
rect 26389 251641 26401 252417
rect 26435 251641 26451 252417
rect 26389 251629 26451 251641
rect 26481 252417 26543 252429
rect 26481 251641 26497 252417
rect 26531 251641 26543 252417
rect 26481 251629 26543 251641
rect 26599 252417 26661 252429
rect 26599 251641 26611 252417
rect 26645 251641 26661 252417
rect 26599 251629 26661 251641
rect 26691 252417 26753 252429
rect 26691 251641 26707 252417
rect 26741 251641 26753 252417
rect 26691 251629 26753 251641
rect 26809 252417 26871 252429
rect 26809 251641 26821 252417
rect 26855 251641 26871 252417
rect 26809 251629 26871 251641
rect 26901 252417 26963 252429
rect 26901 251641 26917 252417
rect 26951 251641 26963 252417
rect 26901 251629 26963 251641
rect 27019 252417 27081 252429
rect 27019 251641 27031 252417
rect 27065 251641 27081 252417
rect 27019 251629 27081 251641
rect 27111 252417 27173 252429
rect 27111 251641 27127 252417
rect 27161 251641 27173 252417
rect 27111 251629 27173 251641
rect 27229 252417 27291 252429
rect 27229 251641 27241 252417
rect 27275 251641 27291 252417
rect 27229 251629 27291 251641
rect 27321 252417 27383 252429
rect 27321 251641 27337 252417
rect 27371 251641 27383 252417
rect 27321 251629 27383 251641
rect -4061 251381 -3999 251393
rect -4061 250605 -4049 251381
rect -4015 250605 -3999 251381
rect -4061 250593 -3999 250605
rect -3969 251381 -3907 251393
rect -3969 250605 -3953 251381
rect -3919 250605 -3907 251381
rect -3969 250593 -3907 250605
rect -3851 251381 -3789 251393
rect -3851 250605 -3839 251381
rect -3805 250605 -3789 251381
rect -3851 250593 -3789 250605
rect -3759 251381 -3697 251393
rect -3759 250605 -3743 251381
rect -3709 250605 -3697 251381
rect -3759 250593 -3697 250605
rect -3641 251381 -3579 251393
rect -3641 250605 -3629 251381
rect -3595 250605 -3579 251381
rect -3641 250593 -3579 250605
rect -3549 251381 -3487 251393
rect -3549 250605 -3533 251381
rect -3499 250605 -3487 251381
rect -3549 250593 -3487 250605
rect -3431 251381 -3369 251393
rect -3431 250605 -3419 251381
rect -3385 250605 -3369 251381
rect -3431 250593 -3369 250605
rect -3339 251381 -3277 251393
rect -3339 250605 -3323 251381
rect -3289 250605 -3277 251381
rect -3339 250593 -3277 250605
rect -3221 251381 -3159 251393
rect -3221 250605 -3209 251381
rect -3175 250605 -3159 251381
rect -3221 250593 -3159 250605
rect -3129 251381 -3067 251393
rect -3129 250605 -3113 251381
rect -3079 250605 -3067 251381
rect -3129 250593 -3067 250605
rect -3011 251381 -2949 251393
rect -3011 250605 -2999 251381
rect -2965 250605 -2949 251381
rect -3011 250593 -2949 250605
rect -2919 251381 -2857 251393
rect -2919 250605 -2903 251381
rect -2869 250605 -2857 251381
rect -2919 250593 -2857 250605
rect -2801 251381 -2739 251393
rect -2801 250605 -2789 251381
rect -2755 250605 -2739 251381
rect -2801 250593 -2739 250605
rect -2709 251381 -2647 251393
rect -2709 250605 -2693 251381
rect -2659 250605 -2647 251381
rect -2709 250593 -2647 250605
rect -2591 251381 -2529 251393
rect -2591 250605 -2579 251381
rect -2545 250605 -2529 251381
rect -2591 250593 -2529 250605
rect -2499 251381 -2437 251393
rect -2499 250605 -2483 251381
rect -2449 250605 -2437 251381
rect -2499 250593 -2437 250605
rect -2381 251381 -2319 251393
rect -2381 250605 -2369 251381
rect -2335 250605 -2319 251381
rect -2381 250593 -2319 250605
rect -2289 251381 -2227 251393
rect -2289 250605 -2273 251381
rect -2239 250605 -2227 251381
rect -2289 250593 -2227 250605
rect -2171 251381 -2109 251393
rect -2171 250605 -2159 251381
rect -2125 250605 -2109 251381
rect -2171 250593 -2109 250605
rect -2079 251381 -2017 251393
rect -2079 250605 -2063 251381
rect -2029 250605 -2017 251381
rect -2079 250593 -2017 250605
rect -1961 251381 -1899 251393
rect -1961 250605 -1949 251381
rect -1915 250605 -1899 251381
rect -1961 250593 -1899 250605
rect -1869 251381 -1807 251393
rect -1869 250605 -1853 251381
rect -1819 250605 -1807 251381
rect -1869 250593 -1807 250605
rect -1751 251381 -1689 251393
rect -1751 250605 -1739 251381
rect -1705 250605 -1689 251381
rect -1751 250593 -1689 250605
rect -1659 251381 -1597 251393
rect -1659 250605 -1643 251381
rect -1609 250605 -1597 251381
rect -1659 250593 -1597 250605
rect -1541 251381 -1479 251393
rect -1541 250605 -1529 251381
rect -1495 250605 -1479 251381
rect -1541 250593 -1479 250605
rect -1449 251381 -1387 251393
rect -1449 250605 -1433 251381
rect -1399 250605 -1387 251381
rect -1449 250593 -1387 250605
rect -1331 251381 -1269 251393
rect -1331 250605 -1319 251381
rect -1285 250605 -1269 251381
rect -1331 250593 -1269 250605
rect -1239 251381 -1177 251393
rect -1239 250605 -1223 251381
rect -1189 250605 -1177 251381
rect -1239 250593 -1177 250605
rect -1121 251381 -1059 251393
rect -1121 250605 -1109 251381
rect -1075 250605 -1059 251381
rect -1121 250593 -1059 250605
rect -1029 251381 -967 251393
rect -1029 250605 -1013 251381
rect -979 250605 -967 251381
rect -1029 250593 -967 250605
rect -911 251381 -849 251393
rect -911 250605 -899 251381
rect -865 250605 -849 251381
rect -911 250593 -849 250605
rect -819 251381 -757 251393
rect -819 250605 -803 251381
rect -769 250605 -757 251381
rect -819 250593 -757 250605
rect -701 251381 -639 251393
rect -701 250605 -689 251381
rect -655 250605 -639 251381
rect -701 250593 -639 250605
rect -609 251381 -547 251393
rect -609 250605 -593 251381
rect -559 250605 -547 251381
rect -609 250593 -547 250605
rect -491 251381 -429 251393
rect -491 250605 -479 251381
rect -445 250605 -429 251381
rect -491 250593 -429 250605
rect -399 251381 -337 251393
rect -399 250605 -383 251381
rect -349 250605 -337 251381
rect -399 250593 -337 250605
rect -281 251381 -219 251393
rect -281 250605 -269 251381
rect -235 250605 -219 251381
rect -281 250593 -219 250605
rect -189 251381 -127 251393
rect -189 250605 -173 251381
rect -139 250605 -127 251381
rect -189 250593 -127 250605
rect -71 251381 -9 251393
rect -71 250605 -59 251381
rect -25 250605 -9 251381
rect -71 250593 -9 250605
rect 21 251381 83 251393
rect 21 250605 37 251381
rect 71 250605 83 251381
rect 21 250593 83 250605
rect 139 251381 201 251393
rect 139 250605 151 251381
rect 185 250605 201 251381
rect 139 250593 201 250605
rect 231 251381 293 251393
rect 231 250605 247 251381
rect 281 250605 293 251381
rect 231 250593 293 250605
rect 349 251381 411 251393
rect 349 250605 361 251381
rect 395 250605 411 251381
rect 349 250593 411 250605
rect 441 251381 503 251393
rect 441 250605 457 251381
rect 491 250605 503 251381
rect 441 250593 503 250605
rect 559 251381 621 251393
rect 559 250605 571 251381
rect 605 250605 621 251381
rect 559 250593 621 250605
rect 651 251381 713 251393
rect 651 250605 667 251381
rect 701 250605 713 251381
rect 651 250593 713 250605
rect 769 251381 831 251393
rect 769 250605 781 251381
rect 815 250605 831 251381
rect 769 250593 831 250605
rect 861 251381 923 251393
rect 861 250605 877 251381
rect 911 250605 923 251381
rect 861 250593 923 250605
rect 979 251381 1041 251393
rect 979 250605 991 251381
rect 1025 250605 1041 251381
rect 979 250593 1041 250605
rect 1071 251381 1133 251393
rect 1071 250605 1087 251381
rect 1121 250605 1133 251381
rect 1071 250593 1133 250605
rect 1189 251381 1251 251393
rect 1189 250605 1201 251381
rect 1235 250605 1251 251381
rect 1189 250593 1251 250605
rect 1281 251381 1343 251393
rect 1281 250605 1297 251381
rect 1331 250605 1343 251381
rect 1281 250593 1343 250605
rect 1399 251381 1461 251393
rect 1399 250605 1411 251381
rect 1445 250605 1461 251381
rect 1399 250593 1461 250605
rect 1491 251381 1553 251393
rect 1491 250605 1507 251381
rect 1541 250605 1553 251381
rect 1491 250593 1553 250605
rect 1609 251381 1671 251393
rect 1609 250605 1621 251381
rect 1655 250605 1671 251381
rect 1609 250593 1671 250605
rect 1701 251381 1763 251393
rect 1701 250605 1717 251381
rect 1751 250605 1763 251381
rect 1701 250593 1763 250605
rect 1819 251381 1881 251393
rect 1819 250605 1831 251381
rect 1865 250605 1881 251381
rect 1819 250593 1881 250605
rect 1911 251381 1973 251393
rect 1911 250605 1927 251381
rect 1961 250605 1973 251381
rect 1911 250593 1973 250605
rect 2029 251381 2091 251393
rect 2029 250605 2041 251381
rect 2075 250605 2091 251381
rect 2029 250593 2091 250605
rect 2121 251381 2183 251393
rect 2121 250605 2137 251381
rect 2171 250605 2183 251381
rect 2121 250593 2183 250605
rect 2239 251381 2301 251393
rect 2239 250605 2251 251381
rect 2285 250605 2301 251381
rect 2239 250593 2301 250605
rect 2331 251381 2393 251393
rect 2331 250605 2347 251381
rect 2381 250605 2393 251381
rect 2331 250593 2393 250605
rect 2449 251381 2511 251393
rect 2449 250605 2461 251381
rect 2495 250605 2511 251381
rect 2449 250593 2511 250605
rect 2541 251381 2603 251393
rect 2541 250605 2557 251381
rect 2591 250605 2603 251381
rect 2541 250593 2603 250605
rect 2659 251381 2721 251393
rect 2659 250605 2671 251381
rect 2705 250605 2721 251381
rect 2659 250593 2721 250605
rect 2751 251381 2813 251393
rect 2751 250605 2767 251381
rect 2801 250605 2813 251381
rect 2751 250593 2813 250605
rect 2869 251381 2931 251393
rect 2869 250605 2881 251381
rect 2915 250605 2931 251381
rect 2869 250593 2931 250605
rect 2961 251381 3023 251393
rect 2961 250605 2977 251381
rect 3011 250605 3023 251381
rect 2961 250593 3023 250605
rect 3079 251381 3141 251393
rect 3079 250605 3091 251381
rect 3125 250605 3141 251381
rect 3079 250593 3141 250605
rect 3171 251381 3233 251393
rect 3171 250605 3187 251381
rect 3221 250605 3233 251381
rect 3171 250593 3233 250605
rect 3289 251381 3351 251393
rect 3289 250605 3301 251381
rect 3335 250605 3351 251381
rect 3289 250593 3351 250605
rect 3381 251381 3443 251393
rect 3381 250605 3397 251381
rect 3431 250605 3443 251381
rect 3381 250593 3443 250605
rect 3499 251381 3561 251393
rect 3499 250605 3511 251381
rect 3545 250605 3561 251381
rect 3499 250593 3561 250605
rect 3591 251381 3653 251393
rect 3591 250605 3607 251381
rect 3641 250605 3653 251381
rect 3591 250593 3653 250605
rect 3709 251381 3771 251393
rect 3709 250605 3721 251381
rect 3755 250605 3771 251381
rect 3709 250593 3771 250605
rect 3801 251381 3863 251393
rect 3801 250605 3817 251381
rect 3851 250605 3863 251381
rect 3801 250593 3863 250605
rect 3919 251381 3981 251393
rect 3919 250605 3931 251381
rect 3965 250605 3981 251381
rect 3919 250593 3981 250605
rect 4011 251381 4073 251393
rect 4011 250605 4027 251381
rect 4061 250605 4073 251381
rect 4011 250593 4073 250605
rect 4129 251381 4191 251393
rect 4129 250605 4141 251381
rect 4175 250605 4191 251381
rect 4129 250593 4191 250605
rect 4221 251381 4283 251393
rect 4221 250605 4237 251381
rect 4271 250605 4283 251381
rect 4221 250593 4283 250605
rect 4339 251381 4401 251393
rect 4339 250605 4351 251381
rect 4385 250605 4401 251381
rect 4339 250593 4401 250605
rect 4431 251381 4493 251393
rect 4431 250605 4447 251381
rect 4481 250605 4493 251381
rect 4431 250593 4493 250605
rect 4549 251381 4611 251393
rect 4549 250605 4561 251381
rect 4595 250605 4611 251381
rect 4549 250593 4611 250605
rect 4641 251381 4703 251393
rect 4641 250605 4657 251381
rect 4691 250605 4703 251381
rect 4641 250593 4703 250605
rect 4759 251381 4821 251393
rect 4759 250605 4771 251381
rect 4805 250605 4821 251381
rect 4759 250593 4821 250605
rect 4851 251381 4913 251393
rect 4851 250605 4867 251381
rect 4901 250605 4913 251381
rect 4851 250593 4913 250605
rect 4969 251381 5031 251393
rect 4969 250605 4981 251381
rect 5015 250605 5031 251381
rect 4969 250593 5031 250605
rect 5061 251381 5123 251393
rect 5061 250605 5077 251381
rect 5111 250605 5123 251381
rect 5061 250593 5123 250605
rect 5179 251381 5241 251393
rect 5179 250605 5191 251381
rect 5225 250605 5241 251381
rect 5179 250593 5241 250605
rect 5271 251381 5333 251393
rect 5271 250605 5287 251381
rect 5321 250605 5333 251381
rect 5271 250593 5333 250605
rect 5389 251381 5451 251393
rect 5389 250605 5401 251381
rect 5435 250605 5451 251381
rect 5389 250593 5451 250605
rect 5481 251381 5543 251393
rect 5481 250605 5497 251381
rect 5531 250605 5543 251381
rect 5481 250593 5543 250605
rect 5599 251381 5661 251393
rect 5599 250605 5611 251381
rect 5645 250605 5661 251381
rect 5599 250593 5661 250605
rect 5691 251381 5753 251393
rect 5691 250605 5707 251381
rect 5741 250605 5753 251381
rect 5691 250593 5753 250605
rect 5809 251381 5871 251393
rect 5809 250605 5821 251381
rect 5855 250605 5871 251381
rect 5809 250593 5871 250605
rect 5901 251381 5963 251393
rect 5901 250605 5917 251381
rect 5951 250605 5963 251381
rect 5901 250593 5963 250605
rect 6019 251381 6081 251393
rect 6019 250605 6031 251381
rect 6065 250605 6081 251381
rect 6019 250593 6081 250605
rect 6111 251381 6173 251393
rect 6111 250605 6127 251381
rect 6161 250605 6173 251381
rect 6111 250593 6173 250605
rect 6229 251381 6291 251393
rect 6229 250605 6241 251381
rect 6275 250605 6291 251381
rect 6229 250593 6291 250605
rect 6321 251381 6383 251393
rect 6321 250605 6337 251381
rect 6371 250605 6383 251381
rect 6321 250593 6383 250605
rect 6439 251381 6501 251393
rect 6439 250605 6451 251381
rect 6485 250605 6501 251381
rect 6439 250593 6501 250605
rect 6531 251381 6593 251393
rect 6531 250605 6547 251381
rect 6581 250605 6593 251381
rect 6531 250593 6593 250605
rect 6649 251381 6711 251393
rect 6649 250605 6661 251381
rect 6695 250605 6711 251381
rect 6649 250593 6711 250605
rect 6741 251381 6803 251393
rect 6741 250605 6757 251381
rect 6791 250605 6803 251381
rect 6741 250593 6803 250605
rect 6859 251381 6921 251393
rect 6859 250605 6871 251381
rect 6905 250605 6921 251381
rect 6859 250593 6921 250605
rect 6951 251381 7013 251393
rect 6951 250605 6967 251381
rect 7001 250605 7013 251381
rect 6951 250593 7013 250605
rect 7069 251381 7131 251393
rect 7069 250605 7081 251381
rect 7115 250605 7131 251381
rect 7069 250593 7131 250605
rect 7161 251381 7223 251393
rect 7161 250605 7177 251381
rect 7211 250605 7223 251381
rect 7161 250593 7223 250605
rect 7279 251381 7341 251393
rect 7279 250605 7291 251381
rect 7325 250605 7341 251381
rect 7279 250593 7341 250605
rect 7371 251381 7433 251393
rect 7371 250605 7387 251381
rect 7421 250605 7433 251381
rect 7371 250593 7433 250605
rect 7489 251381 7551 251393
rect 7489 250605 7501 251381
rect 7535 250605 7551 251381
rect 7489 250593 7551 250605
rect 7581 251381 7643 251393
rect 7581 250605 7597 251381
rect 7631 250605 7643 251381
rect 7581 250593 7643 250605
rect 7699 251381 7761 251393
rect 7699 250605 7711 251381
rect 7745 250605 7761 251381
rect 7699 250593 7761 250605
rect 7791 251381 7853 251393
rect 7791 250605 7807 251381
rect 7841 250605 7853 251381
rect 7791 250593 7853 250605
rect 7909 251381 7971 251393
rect 7909 250605 7921 251381
rect 7955 250605 7971 251381
rect 7909 250593 7971 250605
rect 8001 251381 8063 251393
rect 8001 250605 8017 251381
rect 8051 250605 8063 251381
rect 8001 250593 8063 250605
rect 8119 251381 8181 251393
rect 8119 250605 8131 251381
rect 8165 250605 8181 251381
rect 8119 250593 8181 250605
rect 8211 251381 8273 251393
rect 8211 250605 8227 251381
rect 8261 250605 8273 251381
rect 8211 250593 8273 250605
rect 8329 251381 8391 251393
rect 8329 250605 8341 251381
rect 8375 250605 8391 251381
rect 8329 250593 8391 250605
rect 8421 251381 8483 251393
rect 8421 250605 8437 251381
rect 8471 250605 8483 251381
rect 8421 250593 8483 250605
rect 8539 251381 8601 251393
rect 8539 250605 8551 251381
rect 8585 250605 8601 251381
rect 8539 250593 8601 250605
rect 8631 251381 8693 251393
rect 8631 250605 8647 251381
rect 8681 250605 8693 251381
rect 8631 250593 8693 250605
rect 8749 251381 8811 251393
rect 8749 250605 8761 251381
rect 8795 250605 8811 251381
rect 8749 250593 8811 250605
rect 8841 251381 8903 251393
rect 8841 250605 8857 251381
rect 8891 250605 8903 251381
rect 8841 250593 8903 250605
rect 8959 251381 9021 251393
rect 8959 250605 8971 251381
rect 9005 250605 9021 251381
rect 8959 250593 9021 250605
rect 9051 251381 9113 251393
rect 9051 250605 9067 251381
rect 9101 250605 9113 251381
rect 9051 250593 9113 250605
rect 9169 251381 9231 251393
rect 9169 250605 9181 251381
rect 9215 250605 9231 251381
rect 9169 250593 9231 250605
rect 9261 251381 9323 251393
rect 9261 250605 9277 251381
rect 9311 250605 9323 251381
rect 9261 250593 9323 250605
rect 9379 251381 9441 251393
rect 9379 250605 9391 251381
rect 9425 250605 9441 251381
rect 9379 250593 9441 250605
rect 9471 251381 9533 251393
rect 9471 250605 9487 251381
rect 9521 250605 9533 251381
rect 9471 250593 9533 250605
rect 9589 251381 9651 251393
rect 9589 250605 9601 251381
rect 9635 250605 9651 251381
rect 9589 250593 9651 250605
rect 9681 251381 9743 251393
rect 9681 250605 9697 251381
rect 9731 250605 9743 251381
rect 9681 250593 9743 250605
rect 9799 251381 9861 251393
rect 9799 250605 9811 251381
rect 9845 250605 9861 251381
rect 9799 250593 9861 250605
rect 9891 251381 9953 251393
rect 9891 250605 9907 251381
rect 9941 250605 9953 251381
rect 9891 250593 9953 250605
rect 10009 251381 10071 251393
rect 10009 250605 10021 251381
rect 10055 250605 10071 251381
rect 10009 250593 10071 250605
rect 10101 251381 10163 251393
rect 10101 250605 10117 251381
rect 10151 250605 10163 251381
rect 10101 250593 10163 250605
rect 10219 251381 10281 251393
rect 10219 250605 10231 251381
rect 10265 250605 10281 251381
rect 10219 250593 10281 250605
rect 10311 251381 10373 251393
rect 10311 250605 10327 251381
rect 10361 250605 10373 251381
rect 10311 250593 10373 250605
rect 10429 251381 10491 251393
rect 10429 250605 10441 251381
rect 10475 250605 10491 251381
rect 10429 250593 10491 250605
rect 10521 251381 10583 251393
rect 10521 250605 10537 251381
rect 10571 250605 10583 251381
rect 10521 250593 10583 250605
rect 10639 251381 10701 251393
rect 10639 250605 10651 251381
rect 10685 250605 10701 251381
rect 10639 250593 10701 250605
rect 10731 251381 10793 251393
rect 10731 250605 10747 251381
rect 10781 250605 10793 251381
rect 10731 250593 10793 250605
rect 10849 251381 10911 251393
rect 10849 250605 10861 251381
rect 10895 250605 10911 251381
rect 10849 250593 10911 250605
rect 10941 251381 11003 251393
rect 10941 250605 10957 251381
rect 10991 250605 11003 251381
rect 10941 250593 11003 250605
rect 11059 251381 11121 251393
rect 11059 250605 11071 251381
rect 11105 250605 11121 251381
rect 11059 250593 11121 250605
rect 11151 251381 11213 251393
rect 11151 250605 11167 251381
rect 11201 250605 11213 251381
rect 11151 250593 11213 250605
rect 11269 251381 11331 251393
rect 11269 250605 11281 251381
rect 11315 250605 11331 251381
rect 11269 250593 11331 250605
rect 11361 251381 11423 251393
rect 11361 250605 11377 251381
rect 11411 250605 11423 251381
rect 11361 250593 11423 250605
rect 11479 251381 11541 251393
rect 11479 250605 11491 251381
rect 11525 250605 11541 251381
rect 11479 250593 11541 250605
rect 11571 251381 11633 251393
rect 11571 250605 11587 251381
rect 11621 250605 11633 251381
rect 11571 250593 11633 250605
rect 11689 251381 11751 251393
rect 11689 250605 11701 251381
rect 11735 250605 11751 251381
rect 11689 250593 11751 250605
rect 11781 251381 11843 251393
rect 11781 250605 11797 251381
rect 11831 250605 11843 251381
rect 11781 250593 11843 250605
rect 11899 251381 11961 251393
rect 11899 250605 11911 251381
rect 11945 250605 11961 251381
rect 11899 250593 11961 250605
rect 11991 251381 12053 251393
rect 11991 250605 12007 251381
rect 12041 250605 12053 251381
rect 11991 250593 12053 250605
rect 12109 251381 12171 251393
rect 12109 250605 12121 251381
rect 12155 250605 12171 251381
rect 12109 250593 12171 250605
rect 12201 251381 12263 251393
rect 12201 250605 12217 251381
rect 12251 250605 12263 251381
rect 12201 250593 12263 250605
rect 12319 251381 12381 251393
rect 12319 250605 12331 251381
rect 12365 250605 12381 251381
rect 12319 250593 12381 250605
rect 12411 251381 12473 251393
rect 12411 250605 12427 251381
rect 12461 250605 12473 251381
rect 12411 250593 12473 250605
rect 12529 251381 12591 251393
rect 12529 250605 12541 251381
rect 12575 250605 12591 251381
rect 12529 250593 12591 250605
rect 12621 251381 12683 251393
rect 12621 250605 12637 251381
rect 12671 250605 12683 251381
rect 12621 250593 12683 250605
rect 12739 251381 12801 251393
rect 12739 250605 12751 251381
rect 12785 250605 12801 251381
rect 12739 250593 12801 250605
rect 12831 251381 12893 251393
rect 12831 250605 12847 251381
rect 12881 250605 12893 251381
rect 12831 250593 12893 250605
rect 12949 251381 13011 251393
rect 12949 250605 12961 251381
rect 12995 250605 13011 251381
rect 12949 250593 13011 250605
rect 13041 251381 13103 251393
rect 13041 250605 13057 251381
rect 13091 250605 13103 251381
rect 13041 250593 13103 250605
rect 13159 251381 13221 251393
rect 13159 250605 13171 251381
rect 13205 250605 13221 251381
rect 13159 250593 13221 250605
rect 13251 251381 13313 251393
rect 13251 250605 13267 251381
rect 13301 250605 13313 251381
rect 13251 250593 13313 250605
rect 13369 251381 13431 251393
rect 13369 250605 13381 251381
rect 13415 250605 13431 251381
rect 13369 250593 13431 250605
rect 13461 251381 13523 251393
rect 13461 250605 13477 251381
rect 13511 250605 13523 251381
rect 13461 250593 13523 250605
rect 13579 251381 13641 251393
rect 13579 250605 13591 251381
rect 13625 250605 13641 251381
rect 13579 250593 13641 250605
rect 13671 251381 13733 251393
rect 13671 250605 13687 251381
rect 13721 250605 13733 251381
rect 13671 250593 13733 250605
rect 13789 251381 13851 251393
rect 13789 250605 13801 251381
rect 13835 250605 13851 251381
rect 13789 250593 13851 250605
rect 13881 251381 13943 251393
rect 13881 250605 13897 251381
rect 13931 250605 13943 251381
rect 13881 250593 13943 250605
rect 13999 251381 14061 251393
rect 13999 250605 14011 251381
rect 14045 250605 14061 251381
rect 13999 250593 14061 250605
rect 14091 251381 14153 251393
rect 14091 250605 14107 251381
rect 14141 250605 14153 251381
rect 14091 250593 14153 250605
rect 14209 251381 14271 251393
rect 14209 250605 14221 251381
rect 14255 250605 14271 251381
rect 14209 250593 14271 250605
rect 14301 251381 14363 251393
rect 14301 250605 14317 251381
rect 14351 250605 14363 251381
rect 14301 250593 14363 250605
rect 14419 251381 14481 251393
rect 14419 250605 14431 251381
rect 14465 250605 14481 251381
rect 14419 250593 14481 250605
rect 14511 251381 14573 251393
rect 14511 250605 14527 251381
rect 14561 250605 14573 251381
rect 14511 250593 14573 250605
rect 14629 251381 14691 251393
rect 14629 250605 14641 251381
rect 14675 250605 14691 251381
rect 14629 250593 14691 250605
rect 14721 251381 14783 251393
rect 14721 250605 14737 251381
rect 14771 250605 14783 251381
rect 14721 250593 14783 250605
rect 14839 251381 14901 251393
rect 14839 250605 14851 251381
rect 14885 250605 14901 251381
rect 14839 250593 14901 250605
rect 14931 251381 14993 251393
rect 14931 250605 14947 251381
rect 14981 250605 14993 251381
rect 14931 250593 14993 250605
rect 15049 251381 15111 251393
rect 15049 250605 15061 251381
rect 15095 250605 15111 251381
rect 15049 250593 15111 250605
rect 15141 251381 15203 251393
rect 15141 250605 15157 251381
rect 15191 250605 15203 251381
rect 15141 250593 15203 250605
rect 15259 251381 15321 251393
rect 15259 250605 15271 251381
rect 15305 250605 15321 251381
rect 15259 250593 15321 250605
rect 15351 251381 15413 251393
rect 15351 250605 15367 251381
rect 15401 250605 15413 251381
rect 15351 250593 15413 250605
rect 15469 251381 15531 251393
rect 15469 250605 15481 251381
rect 15515 250605 15531 251381
rect 15469 250593 15531 250605
rect 15561 251381 15623 251393
rect 15561 250605 15577 251381
rect 15611 250605 15623 251381
rect 15561 250593 15623 250605
rect 15679 251381 15741 251393
rect 15679 250605 15691 251381
rect 15725 250605 15741 251381
rect 15679 250593 15741 250605
rect 15771 251381 15833 251393
rect 15771 250605 15787 251381
rect 15821 250605 15833 251381
rect 15771 250593 15833 250605
rect 15889 251381 15951 251393
rect 15889 250605 15901 251381
rect 15935 250605 15951 251381
rect 15889 250593 15951 250605
rect 15981 251381 16043 251393
rect 15981 250605 15997 251381
rect 16031 250605 16043 251381
rect 15981 250593 16043 250605
rect 16099 251381 16161 251393
rect 16099 250605 16111 251381
rect 16145 250605 16161 251381
rect 16099 250593 16161 250605
rect 16191 251381 16253 251393
rect 16191 250605 16207 251381
rect 16241 250605 16253 251381
rect 16191 250593 16253 250605
rect 16309 251381 16371 251393
rect 16309 250605 16321 251381
rect 16355 250605 16371 251381
rect 16309 250593 16371 250605
rect 16401 251381 16463 251393
rect 16401 250605 16417 251381
rect 16451 250605 16463 251381
rect 16401 250593 16463 250605
rect 16519 251381 16581 251393
rect 16519 250605 16531 251381
rect 16565 250605 16581 251381
rect 16519 250593 16581 250605
rect 16611 251381 16673 251393
rect 16611 250605 16627 251381
rect 16661 250605 16673 251381
rect 16611 250593 16673 250605
rect 16729 251381 16791 251393
rect 16729 250605 16741 251381
rect 16775 250605 16791 251381
rect 16729 250593 16791 250605
rect 16821 251381 16883 251393
rect 16821 250605 16837 251381
rect 16871 250605 16883 251381
rect 16821 250593 16883 250605
rect 16939 251381 17001 251393
rect 16939 250605 16951 251381
rect 16985 250605 17001 251381
rect 16939 250593 17001 250605
rect 17031 251381 17093 251393
rect 17031 250605 17047 251381
rect 17081 250605 17093 251381
rect 17031 250593 17093 250605
rect 17149 251381 17211 251393
rect 17149 250605 17161 251381
rect 17195 250605 17211 251381
rect 17149 250593 17211 250605
rect 17241 251381 17303 251393
rect 17241 250605 17257 251381
rect 17291 250605 17303 251381
rect 17241 250593 17303 250605
rect 17359 251381 17421 251393
rect 17359 250605 17371 251381
rect 17405 250605 17421 251381
rect 17359 250593 17421 250605
rect 17451 251381 17513 251393
rect 17451 250605 17467 251381
rect 17501 250605 17513 251381
rect 17451 250593 17513 250605
rect 17569 251381 17631 251393
rect 17569 250605 17581 251381
rect 17615 250605 17631 251381
rect 17569 250593 17631 250605
rect 17661 251381 17723 251393
rect 17661 250605 17677 251381
rect 17711 250605 17723 251381
rect 17661 250593 17723 250605
rect 17779 251381 17841 251393
rect 17779 250605 17791 251381
rect 17825 250605 17841 251381
rect 17779 250593 17841 250605
rect 17871 251381 17933 251393
rect 17871 250605 17887 251381
rect 17921 250605 17933 251381
rect 17871 250593 17933 250605
rect 17989 251381 18051 251393
rect 17989 250605 18001 251381
rect 18035 250605 18051 251381
rect 17989 250593 18051 250605
rect 18081 251381 18143 251393
rect 18081 250605 18097 251381
rect 18131 250605 18143 251381
rect 18081 250593 18143 250605
rect 18199 251381 18261 251393
rect 18199 250605 18211 251381
rect 18245 250605 18261 251381
rect 18199 250593 18261 250605
rect 18291 251381 18353 251393
rect 18291 250605 18307 251381
rect 18341 250605 18353 251381
rect 18291 250593 18353 250605
rect 18409 251381 18471 251393
rect 18409 250605 18421 251381
rect 18455 250605 18471 251381
rect 18409 250593 18471 250605
rect 18501 251381 18563 251393
rect 18501 250605 18517 251381
rect 18551 250605 18563 251381
rect 18501 250593 18563 250605
rect 18619 251381 18681 251393
rect 18619 250605 18631 251381
rect 18665 250605 18681 251381
rect 18619 250593 18681 250605
rect 18711 251381 18773 251393
rect 18711 250605 18727 251381
rect 18761 250605 18773 251381
rect 18711 250593 18773 250605
rect 18829 251381 18891 251393
rect 18829 250605 18841 251381
rect 18875 250605 18891 251381
rect 18829 250593 18891 250605
rect 18921 251381 18983 251393
rect 18921 250605 18937 251381
rect 18971 250605 18983 251381
rect 18921 250593 18983 250605
rect 19039 251381 19101 251393
rect 19039 250605 19051 251381
rect 19085 250605 19101 251381
rect 19039 250593 19101 250605
rect 19131 251381 19193 251393
rect 19131 250605 19147 251381
rect 19181 250605 19193 251381
rect 19131 250593 19193 250605
rect 19249 251381 19311 251393
rect 19249 250605 19261 251381
rect 19295 250605 19311 251381
rect 19249 250593 19311 250605
rect 19341 251381 19403 251393
rect 19341 250605 19357 251381
rect 19391 250605 19403 251381
rect 19341 250593 19403 250605
rect 19459 251381 19521 251393
rect 19459 250605 19471 251381
rect 19505 250605 19521 251381
rect 19459 250593 19521 250605
rect 19551 251381 19613 251393
rect 19551 250605 19567 251381
rect 19601 250605 19613 251381
rect 19551 250593 19613 250605
rect 19669 251381 19731 251393
rect 19669 250605 19681 251381
rect 19715 250605 19731 251381
rect 19669 250593 19731 250605
rect 19761 251381 19823 251393
rect 19761 250605 19777 251381
rect 19811 250605 19823 251381
rect 19761 250593 19823 250605
rect 19879 251381 19941 251393
rect 19879 250605 19891 251381
rect 19925 250605 19941 251381
rect 19879 250593 19941 250605
rect 19971 251381 20033 251393
rect 19971 250605 19987 251381
rect 20021 250605 20033 251381
rect 19971 250593 20033 250605
rect 20089 251381 20151 251393
rect 20089 250605 20101 251381
rect 20135 250605 20151 251381
rect 20089 250593 20151 250605
rect 20181 251381 20243 251393
rect 20181 250605 20197 251381
rect 20231 250605 20243 251381
rect 20181 250593 20243 250605
rect 20299 251381 20361 251393
rect 20299 250605 20311 251381
rect 20345 250605 20361 251381
rect 20299 250593 20361 250605
rect 20391 251381 20453 251393
rect 20391 250605 20407 251381
rect 20441 250605 20453 251381
rect 20391 250593 20453 250605
rect 20509 251381 20571 251393
rect 20509 250605 20521 251381
rect 20555 250605 20571 251381
rect 20509 250593 20571 250605
rect 20601 251381 20663 251393
rect 20601 250605 20617 251381
rect 20651 250605 20663 251381
rect 20601 250593 20663 250605
rect 20719 251381 20781 251393
rect 20719 250605 20731 251381
rect 20765 250605 20781 251381
rect 20719 250593 20781 250605
rect 20811 251381 20873 251393
rect 20811 250605 20827 251381
rect 20861 250605 20873 251381
rect 20811 250593 20873 250605
rect 20929 251381 20991 251393
rect 20929 250605 20941 251381
rect 20975 250605 20991 251381
rect 20929 250593 20991 250605
rect 21021 251381 21083 251393
rect 21021 250605 21037 251381
rect 21071 250605 21083 251381
rect 21021 250593 21083 250605
rect 21139 251381 21201 251393
rect 21139 250605 21151 251381
rect 21185 250605 21201 251381
rect 21139 250593 21201 250605
rect 21231 251381 21293 251393
rect 21231 250605 21247 251381
rect 21281 250605 21293 251381
rect 21231 250593 21293 250605
rect 21349 251381 21411 251393
rect 21349 250605 21361 251381
rect 21395 250605 21411 251381
rect 21349 250593 21411 250605
rect 21441 251381 21503 251393
rect 21441 250605 21457 251381
rect 21491 250605 21503 251381
rect 21441 250593 21503 250605
rect 21559 251381 21621 251393
rect 21559 250605 21571 251381
rect 21605 250605 21621 251381
rect 21559 250593 21621 250605
rect 21651 251381 21713 251393
rect 21651 250605 21667 251381
rect 21701 250605 21713 251381
rect 21651 250593 21713 250605
rect 21769 251381 21831 251393
rect 21769 250605 21781 251381
rect 21815 250605 21831 251381
rect 21769 250593 21831 250605
rect 21861 251381 21923 251393
rect 21861 250605 21877 251381
rect 21911 250605 21923 251381
rect 21861 250593 21923 250605
rect 21979 251381 22041 251393
rect 21979 250605 21991 251381
rect 22025 250605 22041 251381
rect 21979 250593 22041 250605
rect 22071 251381 22133 251393
rect 22071 250605 22087 251381
rect 22121 250605 22133 251381
rect 22071 250593 22133 250605
rect 22189 251381 22251 251393
rect 22189 250605 22201 251381
rect 22235 250605 22251 251381
rect 22189 250593 22251 250605
rect 22281 251381 22343 251393
rect 22281 250605 22297 251381
rect 22331 250605 22343 251381
rect 22281 250593 22343 250605
rect 22399 251381 22461 251393
rect 22399 250605 22411 251381
rect 22445 250605 22461 251381
rect 22399 250593 22461 250605
rect 22491 251381 22553 251393
rect 22491 250605 22507 251381
rect 22541 250605 22553 251381
rect 22491 250593 22553 250605
rect 22609 251381 22671 251393
rect 22609 250605 22621 251381
rect 22655 250605 22671 251381
rect 22609 250593 22671 250605
rect 22701 251381 22763 251393
rect 22701 250605 22717 251381
rect 22751 250605 22763 251381
rect 22701 250593 22763 250605
rect 22819 251381 22881 251393
rect 22819 250605 22831 251381
rect 22865 250605 22881 251381
rect 22819 250593 22881 250605
rect 22911 251381 22973 251393
rect 22911 250605 22927 251381
rect 22961 250605 22973 251381
rect 22911 250593 22973 250605
rect 23029 251381 23091 251393
rect 23029 250605 23041 251381
rect 23075 250605 23091 251381
rect 23029 250593 23091 250605
rect 23121 251381 23183 251393
rect 23121 250605 23137 251381
rect 23171 250605 23183 251381
rect 23121 250593 23183 250605
rect 23239 251381 23301 251393
rect 23239 250605 23251 251381
rect 23285 250605 23301 251381
rect 23239 250593 23301 250605
rect 23331 251381 23393 251393
rect 23331 250605 23347 251381
rect 23381 250605 23393 251381
rect 23331 250593 23393 250605
rect 23449 251381 23511 251393
rect 23449 250605 23461 251381
rect 23495 250605 23511 251381
rect 23449 250593 23511 250605
rect 23541 251381 23603 251393
rect 23541 250605 23557 251381
rect 23591 250605 23603 251381
rect 23541 250593 23603 250605
rect 23659 251381 23721 251393
rect 23659 250605 23671 251381
rect 23705 250605 23721 251381
rect 23659 250593 23721 250605
rect 23751 251381 23813 251393
rect 23751 250605 23767 251381
rect 23801 250605 23813 251381
rect 23751 250593 23813 250605
rect 23869 251381 23931 251393
rect 23869 250605 23881 251381
rect 23915 250605 23931 251381
rect 23869 250593 23931 250605
rect 23961 251381 24023 251393
rect 23961 250605 23977 251381
rect 24011 250605 24023 251381
rect 23961 250593 24023 250605
rect 24079 251381 24141 251393
rect 24079 250605 24091 251381
rect 24125 250605 24141 251381
rect 24079 250593 24141 250605
rect 24171 251381 24233 251393
rect 24171 250605 24187 251381
rect 24221 250605 24233 251381
rect 24171 250593 24233 250605
rect 24289 251381 24351 251393
rect 24289 250605 24301 251381
rect 24335 250605 24351 251381
rect 24289 250593 24351 250605
rect 24381 251381 24443 251393
rect 24381 250605 24397 251381
rect 24431 250605 24443 251381
rect 24381 250593 24443 250605
rect 24499 251381 24561 251393
rect 24499 250605 24511 251381
rect 24545 250605 24561 251381
rect 24499 250593 24561 250605
rect 24591 251381 24653 251393
rect 24591 250605 24607 251381
rect 24641 250605 24653 251381
rect 24591 250593 24653 250605
rect 24709 251381 24771 251393
rect 24709 250605 24721 251381
rect 24755 250605 24771 251381
rect 24709 250593 24771 250605
rect 24801 251381 24863 251393
rect 24801 250605 24817 251381
rect 24851 250605 24863 251381
rect 24801 250593 24863 250605
rect 24919 251381 24981 251393
rect 24919 250605 24931 251381
rect 24965 250605 24981 251381
rect 24919 250593 24981 250605
rect 25011 251381 25073 251393
rect 25011 250605 25027 251381
rect 25061 250605 25073 251381
rect 25011 250593 25073 250605
rect 25129 251381 25191 251393
rect 25129 250605 25141 251381
rect 25175 250605 25191 251381
rect 25129 250593 25191 250605
rect 25221 251381 25283 251393
rect 25221 250605 25237 251381
rect 25271 250605 25283 251381
rect 25221 250593 25283 250605
rect 25339 251381 25401 251393
rect 25339 250605 25351 251381
rect 25385 250605 25401 251381
rect 25339 250593 25401 250605
rect 25431 251381 25493 251393
rect 25431 250605 25447 251381
rect 25481 250605 25493 251381
rect 25431 250593 25493 250605
rect 25549 251381 25611 251393
rect 25549 250605 25561 251381
rect 25595 250605 25611 251381
rect 25549 250593 25611 250605
rect 25641 251381 25703 251393
rect 25641 250605 25657 251381
rect 25691 250605 25703 251381
rect 25641 250593 25703 250605
rect 25759 251381 25821 251393
rect 25759 250605 25771 251381
rect 25805 250605 25821 251381
rect 25759 250593 25821 250605
rect 25851 251381 25913 251393
rect 25851 250605 25867 251381
rect 25901 250605 25913 251381
rect 25851 250593 25913 250605
rect 25969 251381 26031 251393
rect 25969 250605 25981 251381
rect 26015 250605 26031 251381
rect 25969 250593 26031 250605
rect 26061 251381 26123 251393
rect 26061 250605 26077 251381
rect 26111 250605 26123 251381
rect 26061 250593 26123 250605
rect 26179 251381 26241 251393
rect 26179 250605 26191 251381
rect 26225 250605 26241 251381
rect 26179 250593 26241 250605
rect 26271 251381 26333 251393
rect 26271 250605 26287 251381
rect 26321 250605 26333 251381
rect 26271 250593 26333 250605
rect 26389 251381 26451 251393
rect 26389 250605 26401 251381
rect 26435 250605 26451 251381
rect 26389 250593 26451 250605
rect 26481 251381 26543 251393
rect 26481 250605 26497 251381
rect 26531 250605 26543 251381
rect 26481 250593 26543 250605
rect 26599 251381 26661 251393
rect 26599 250605 26611 251381
rect 26645 250605 26661 251381
rect 26599 250593 26661 250605
rect 26691 251381 26753 251393
rect 26691 250605 26707 251381
rect 26741 250605 26753 251381
rect 26691 250593 26753 250605
rect 26809 251381 26871 251393
rect 26809 250605 26821 251381
rect 26855 250605 26871 251381
rect 26809 250593 26871 250605
rect 26901 251381 26963 251393
rect 26901 250605 26917 251381
rect 26951 250605 26963 251381
rect 26901 250593 26963 250605
rect 27019 251381 27081 251393
rect 27019 250605 27031 251381
rect 27065 250605 27081 251381
rect 27019 250593 27081 250605
rect 27111 251381 27173 251393
rect 27111 250605 27127 251381
rect 27161 250605 27173 251381
rect 27111 250593 27173 250605
rect 27229 251381 27291 251393
rect 27229 250605 27241 251381
rect 27275 250605 27291 251381
rect 27229 250593 27291 250605
rect 27321 251381 27383 251393
rect 27321 250605 27337 251381
rect 27371 250605 27383 251381
rect 27321 250593 27383 250605
rect -4061 250345 -3999 250357
rect -4061 249569 -4049 250345
rect -4015 249569 -3999 250345
rect -4061 249557 -3999 249569
rect -3969 250345 -3907 250357
rect -3969 249569 -3953 250345
rect -3919 249569 -3907 250345
rect -3969 249557 -3907 249569
rect -3851 250345 -3789 250357
rect -3851 249569 -3839 250345
rect -3805 249569 -3789 250345
rect -3851 249557 -3789 249569
rect -3759 250345 -3697 250357
rect -3759 249569 -3743 250345
rect -3709 249569 -3697 250345
rect -3759 249557 -3697 249569
rect -3641 250345 -3579 250357
rect -3641 249569 -3629 250345
rect -3595 249569 -3579 250345
rect -3641 249557 -3579 249569
rect -3549 250345 -3487 250357
rect -3549 249569 -3533 250345
rect -3499 249569 -3487 250345
rect -3549 249557 -3487 249569
rect -3431 250345 -3369 250357
rect -3431 249569 -3419 250345
rect -3385 249569 -3369 250345
rect -3431 249557 -3369 249569
rect -3339 250345 -3277 250357
rect -3339 249569 -3323 250345
rect -3289 249569 -3277 250345
rect -3339 249557 -3277 249569
rect -3221 250345 -3159 250357
rect -3221 249569 -3209 250345
rect -3175 249569 -3159 250345
rect -3221 249557 -3159 249569
rect -3129 250345 -3067 250357
rect -3129 249569 -3113 250345
rect -3079 249569 -3067 250345
rect -3129 249557 -3067 249569
rect -3011 250345 -2949 250357
rect -3011 249569 -2999 250345
rect -2965 249569 -2949 250345
rect -3011 249557 -2949 249569
rect -2919 250345 -2857 250357
rect -2919 249569 -2903 250345
rect -2869 249569 -2857 250345
rect -2919 249557 -2857 249569
rect -2801 250345 -2739 250357
rect -2801 249569 -2789 250345
rect -2755 249569 -2739 250345
rect -2801 249557 -2739 249569
rect -2709 250345 -2647 250357
rect -2709 249569 -2693 250345
rect -2659 249569 -2647 250345
rect -2709 249557 -2647 249569
rect -2591 250345 -2529 250357
rect -2591 249569 -2579 250345
rect -2545 249569 -2529 250345
rect -2591 249557 -2529 249569
rect -2499 250345 -2437 250357
rect -2499 249569 -2483 250345
rect -2449 249569 -2437 250345
rect -2499 249557 -2437 249569
rect -2381 250345 -2319 250357
rect -2381 249569 -2369 250345
rect -2335 249569 -2319 250345
rect -2381 249557 -2319 249569
rect -2289 250345 -2227 250357
rect -2289 249569 -2273 250345
rect -2239 249569 -2227 250345
rect -2289 249557 -2227 249569
rect -2171 250345 -2109 250357
rect -2171 249569 -2159 250345
rect -2125 249569 -2109 250345
rect -2171 249557 -2109 249569
rect -2079 250345 -2017 250357
rect -2079 249569 -2063 250345
rect -2029 249569 -2017 250345
rect -2079 249557 -2017 249569
rect -1961 250345 -1899 250357
rect -1961 249569 -1949 250345
rect -1915 249569 -1899 250345
rect -1961 249557 -1899 249569
rect -1869 250345 -1807 250357
rect -1869 249569 -1853 250345
rect -1819 249569 -1807 250345
rect -1869 249557 -1807 249569
rect -1751 250345 -1689 250357
rect -1751 249569 -1739 250345
rect -1705 249569 -1689 250345
rect -1751 249557 -1689 249569
rect -1659 250345 -1597 250357
rect -1659 249569 -1643 250345
rect -1609 249569 -1597 250345
rect -1659 249557 -1597 249569
rect -1541 250345 -1479 250357
rect -1541 249569 -1529 250345
rect -1495 249569 -1479 250345
rect -1541 249557 -1479 249569
rect -1449 250345 -1387 250357
rect -1449 249569 -1433 250345
rect -1399 249569 -1387 250345
rect -1449 249557 -1387 249569
rect -1331 250345 -1269 250357
rect -1331 249569 -1319 250345
rect -1285 249569 -1269 250345
rect -1331 249557 -1269 249569
rect -1239 250345 -1177 250357
rect -1239 249569 -1223 250345
rect -1189 249569 -1177 250345
rect -1239 249557 -1177 249569
rect -1121 250345 -1059 250357
rect -1121 249569 -1109 250345
rect -1075 249569 -1059 250345
rect -1121 249557 -1059 249569
rect -1029 250345 -967 250357
rect -1029 249569 -1013 250345
rect -979 249569 -967 250345
rect -1029 249557 -967 249569
rect -911 250345 -849 250357
rect -911 249569 -899 250345
rect -865 249569 -849 250345
rect -911 249557 -849 249569
rect -819 250345 -757 250357
rect -819 249569 -803 250345
rect -769 249569 -757 250345
rect -819 249557 -757 249569
rect -701 250345 -639 250357
rect -701 249569 -689 250345
rect -655 249569 -639 250345
rect -701 249557 -639 249569
rect -609 250345 -547 250357
rect -609 249569 -593 250345
rect -559 249569 -547 250345
rect -609 249557 -547 249569
rect -491 250345 -429 250357
rect -491 249569 -479 250345
rect -445 249569 -429 250345
rect -491 249557 -429 249569
rect -399 250345 -337 250357
rect -399 249569 -383 250345
rect -349 249569 -337 250345
rect -399 249557 -337 249569
rect -281 250345 -219 250357
rect -281 249569 -269 250345
rect -235 249569 -219 250345
rect -281 249557 -219 249569
rect -189 250345 -127 250357
rect -189 249569 -173 250345
rect -139 249569 -127 250345
rect -189 249557 -127 249569
rect -71 250345 -9 250357
rect -71 249569 -59 250345
rect -25 249569 -9 250345
rect -71 249557 -9 249569
rect 21 250345 83 250357
rect 21 249569 37 250345
rect 71 249569 83 250345
rect 21 249557 83 249569
rect 139 250345 201 250357
rect 139 249569 151 250345
rect 185 249569 201 250345
rect 139 249557 201 249569
rect 231 250345 293 250357
rect 231 249569 247 250345
rect 281 249569 293 250345
rect 231 249557 293 249569
rect 349 250345 411 250357
rect 349 249569 361 250345
rect 395 249569 411 250345
rect 349 249557 411 249569
rect 441 250345 503 250357
rect 441 249569 457 250345
rect 491 249569 503 250345
rect 441 249557 503 249569
rect 559 250345 621 250357
rect 559 249569 571 250345
rect 605 249569 621 250345
rect 559 249557 621 249569
rect 651 250345 713 250357
rect 651 249569 667 250345
rect 701 249569 713 250345
rect 651 249557 713 249569
rect 769 250345 831 250357
rect 769 249569 781 250345
rect 815 249569 831 250345
rect 769 249557 831 249569
rect 861 250345 923 250357
rect 861 249569 877 250345
rect 911 249569 923 250345
rect 861 249557 923 249569
rect 979 250345 1041 250357
rect 979 249569 991 250345
rect 1025 249569 1041 250345
rect 979 249557 1041 249569
rect 1071 250345 1133 250357
rect 1071 249569 1087 250345
rect 1121 249569 1133 250345
rect 1071 249557 1133 249569
rect 1189 250345 1251 250357
rect 1189 249569 1201 250345
rect 1235 249569 1251 250345
rect 1189 249557 1251 249569
rect 1281 250345 1343 250357
rect 1281 249569 1297 250345
rect 1331 249569 1343 250345
rect 1281 249557 1343 249569
rect 1399 250345 1461 250357
rect 1399 249569 1411 250345
rect 1445 249569 1461 250345
rect 1399 249557 1461 249569
rect 1491 250345 1553 250357
rect 1491 249569 1507 250345
rect 1541 249569 1553 250345
rect 1491 249557 1553 249569
rect 1609 250345 1671 250357
rect 1609 249569 1621 250345
rect 1655 249569 1671 250345
rect 1609 249557 1671 249569
rect 1701 250345 1763 250357
rect 1701 249569 1717 250345
rect 1751 249569 1763 250345
rect 1701 249557 1763 249569
rect 1819 250345 1881 250357
rect 1819 249569 1831 250345
rect 1865 249569 1881 250345
rect 1819 249557 1881 249569
rect 1911 250345 1973 250357
rect 1911 249569 1927 250345
rect 1961 249569 1973 250345
rect 1911 249557 1973 249569
rect 2029 250345 2091 250357
rect 2029 249569 2041 250345
rect 2075 249569 2091 250345
rect 2029 249557 2091 249569
rect 2121 250345 2183 250357
rect 2121 249569 2137 250345
rect 2171 249569 2183 250345
rect 2121 249557 2183 249569
rect 2239 250345 2301 250357
rect 2239 249569 2251 250345
rect 2285 249569 2301 250345
rect 2239 249557 2301 249569
rect 2331 250345 2393 250357
rect 2331 249569 2347 250345
rect 2381 249569 2393 250345
rect 2331 249557 2393 249569
rect 2449 250345 2511 250357
rect 2449 249569 2461 250345
rect 2495 249569 2511 250345
rect 2449 249557 2511 249569
rect 2541 250345 2603 250357
rect 2541 249569 2557 250345
rect 2591 249569 2603 250345
rect 2541 249557 2603 249569
rect 2659 250345 2721 250357
rect 2659 249569 2671 250345
rect 2705 249569 2721 250345
rect 2659 249557 2721 249569
rect 2751 250345 2813 250357
rect 2751 249569 2767 250345
rect 2801 249569 2813 250345
rect 2751 249557 2813 249569
rect 2869 250345 2931 250357
rect 2869 249569 2881 250345
rect 2915 249569 2931 250345
rect 2869 249557 2931 249569
rect 2961 250345 3023 250357
rect 2961 249569 2977 250345
rect 3011 249569 3023 250345
rect 2961 249557 3023 249569
rect 3079 250345 3141 250357
rect 3079 249569 3091 250345
rect 3125 249569 3141 250345
rect 3079 249557 3141 249569
rect 3171 250345 3233 250357
rect 3171 249569 3187 250345
rect 3221 249569 3233 250345
rect 3171 249557 3233 249569
rect 3289 250345 3351 250357
rect 3289 249569 3301 250345
rect 3335 249569 3351 250345
rect 3289 249557 3351 249569
rect 3381 250345 3443 250357
rect 3381 249569 3397 250345
rect 3431 249569 3443 250345
rect 3381 249557 3443 249569
rect 3499 250345 3561 250357
rect 3499 249569 3511 250345
rect 3545 249569 3561 250345
rect 3499 249557 3561 249569
rect 3591 250345 3653 250357
rect 3591 249569 3607 250345
rect 3641 249569 3653 250345
rect 3591 249557 3653 249569
rect 3709 250345 3771 250357
rect 3709 249569 3721 250345
rect 3755 249569 3771 250345
rect 3709 249557 3771 249569
rect 3801 250345 3863 250357
rect 3801 249569 3817 250345
rect 3851 249569 3863 250345
rect 3801 249557 3863 249569
rect 3919 250345 3981 250357
rect 3919 249569 3931 250345
rect 3965 249569 3981 250345
rect 3919 249557 3981 249569
rect 4011 250345 4073 250357
rect 4011 249569 4027 250345
rect 4061 249569 4073 250345
rect 4011 249557 4073 249569
rect 4129 250345 4191 250357
rect 4129 249569 4141 250345
rect 4175 249569 4191 250345
rect 4129 249557 4191 249569
rect 4221 250345 4283 250357
rect 4221 249569 4237 250345
rect 4271 249569 4283 250345
rect 4221 249557 4283 249569
rect 4339 250345 4401 250357
rect 4339 249569 4351 250345
rect 4385 249569 4401 250345
rect 4339 249557 4401 249569
rect 4431 250345 4493 250357
rect 4431 249569 4447 250345
rect 4481 249569 4493 250345
rect 4431 249557 4493 249569
rect 4549 250345 4611 250357
rect 4549 249569 4561 250345
rect 4595 249569 4611 250345
rect 4549 249557 4611 249569
rect 4641 250345 4703 250357
rect 4641 249569 4657 250345
rect 4691 249569 4703 250345
rect 4641 249557 4703 249569
rect 4759 250345 4821 250357
rect 4759 249569 4771 250345
rect 4805 249569 4821 250345
rect 4759 249557 4821 249569
rect 4851 250345 4913 250357
rect 4851 249569 4867 250345
rect 4901 249569 4913 250345
rect 4851 249557 4913 249569
rect 4969 250345 5031 250357
rect 4969 249569 4981 250345
rect 5015 249569 5031 250345
rect 4969 249557 5031 249569
rect 5061 250345 5123 250357
rect 5061 249569 5077 250345
rect 5111 249569 5123 250345
rect 5061 249557 5123 249569
rect 5179 250345 5241 250357
rect 5179 249569 5191 250345
rect 5225 249569 5241 250345
rect 5179 249557 5241 249569
rect 5271 250345 5333 250357
rect 5271 249569 5287 250345
rect 5321 249569 5333 250345
rect 5271 249557 5333 249569
rect 5389 250345 5451 250357
rect 5389 249569 5401 250345
rect 5435 249569 5451 250345
rect 5389 249557 5451 249569
rect 5481 250345 5543 250357
rect 5481 249569 5497 250345
rect 5531 249569 5543 250345
rect 5481 249557 5543 249569
rect 5599 250345 5661 250357
rect 5599 249569 5611 250345
rect 5645 249569 5661 250345
rect 5599 249557 5661 249569
rect 5691 250345 5753 250357
rect 5691 249569 5707 250345
rect 5741 249569 5753 250345
rect 5691 249557 5753 249569
rect 5809 250345 5871 250357
rect 5809 249569 5821 250345
rect 5855 249569 5871 250345
rect 5809 249557 5871 249569
rect 5901 250345 5963 250357
rect 5901 249569 5917 250345
rect 5951 249569 5963 250345
rect 5901 249557 5963 249569
rect 6019 250345 6081 250357
rect 6019 249569 6031 250345
rect 6065 249569 6081 250345
rect 6019 249557 6081 249569
rect 6111 250345 6173 250357
rect 6111 249569 6127 250345
rect 6161 249569 6173 250345
rect 6111 249557 6173 249569
rect 6229 250345 6291 250357
rect 6229 249569 6241 250345
rect 6275 249569 6291 250345
rect 6229 249557 6291 249569
rect 6321 250345 6383 250357
rect 6321 249569 6337 250345
rect 6371 249569 6383 250345
rect 6321 249557 6383 249569
rect 6439 250345 6501 250357
rect 6439 249569 6451 250345
rect 6485 249569 6501 250345
rect 6439 249557 6501 249569
rect 6531 250345 6593 250357
rect 6531 249569 6547 250345
rect 6581 249569 6593 250345
rect 6531 249557 6593 249569
rect 6649 250345 6711 250357
rect 6649 249569 6661 250345
rect 6695 249569 6711 250345
rect 6649 249557 6711 249569
rect 6741 250345 6803 250357
rect 6741 249569 6757 250345
rect 6791 249569 6803 250345
rect 6741 249557 6803 249569
rect 6859 250345 6921 250357
rect 6859 249569 6871 250345
rect 6905 249569 6921 250345
rect 6859 249557 6921 249569
rect 6951 250345 7013 250357
rect 6951 249569 6967 250345
rect 7001 249569 7013 250345
rect 6951 249557 7013 249569
rect 7069 250345 7131 250357
rect 7069 249569 7081 250345
rect 7115 249569 7131 250345
rect 7069 249557 7131 249569
rect 7161 250345 7223 250357
rect 7161 249569 7177 250345
rect 7211 249569 7223 250345
rect 7161 249557 7223 249569
rect 7279 250345 7341 250357
rect 7279 249569 7291 250345
rect 7325 249569 7341 250345
rect 7279 249557 7341 249569
rect 7371 250345 7433 250357
rect 7371 249569 7387 250345
rect 7421 249569 7433 250345
rect 7371 249557 7433 249569
rect 7489 250345 7551 250357
rect 7489 249569 7501 250345
rect 7535 249569 7551 250345
rect 7489 249557 7551 249569
rect 7581 250345 7643 250357
rect 7581 249569 7597 250345
rect 7631 249569 7643 250345
rect 7581 249557 7643 249569
rect 7699 250345 7761 250357
rect 7699 249569 7711 250345
rect 7745 249569 7761 250345
rect 7699 249557 7761 249569
rect 7791 250345 7853 250357
rect 7791 249569 7807 250345
rect 7841 249569 7853 250345
rect 7791 249557 7853 249569
rect 7909 250345 7971 250357
rect 7909 249569 7921 250345
rect 7955 249569 7971 250345
rect 7909 249557 7971 249569
rect 8001 250345 8063 250357
rect 8001 249569 8017 250345
rect 8051 249569 8063 250345
rect 8001 249557 8063 249569
rect 8119 250345 8181 250357
rect 8119 249569 8131 250345
rect 8165 249569 8181 250345
rect 8119 249557 8181 249569
rect 8211 250345 8273 250357
rect 8211 249569 8227 250345
rect 8261 249569 8273 250345
rect 8211 249557 8273 249569
rect 8329 250345 8391 250357
rect 8329 249569 8341 250345
rect 8375 249569 8391 250345
rect 8329 249557 8391 249569
rect 8421 250345 8483 250357
rect 8421 249569 8437 250345
rect 8471 249569 8483 250345
rect 8421 249557 8483 249569
rect 8539 250345 8601 250357
rect 8539 249569 8551 250345
rect 8585 249569 8601 250345
rect 8539 249557 8601 249569
rect 8631 250345 8693 250357
rect 8631 249569 8647 250345
rect 8681 249569 8693 250345
rect 8631 249557 8693 249569
rect 8749 250345 8811 250357
rect 8749 249569 8761 250345
rect 8795 249569 8811 250345
rect 8749 249557 8811 249569
rect 8841 250345 8903 250357
rect 8841 249569 8857 250345
rect 8891 249569 8903 250345
rect 8841 249557 8903 249569
rect 8959 250345 9021 250357
rect 8959 249569 8971 250345
rect 9005 249569 9021 250345
rect 8959 249557 9021 249569
rect 9051 250345 9113 250357
rect 9051 249569 9067 250345
rect 9101 249569 9113 250345
rect 9051 249557 9113 249569
rect 9169 250345 9231 250357
rect 9169 249569 9181 250345
rect 9215 249569 9231 250345
rect 9169 249557 9231 249569
rect 9261 250345 9323 250357
rect 9261 249569 9277 250345
rect 9311 249569 9323 250345
rect 9261 249557 9323 249569
rect 9379 250345 9441 250357
rect 9379 249569 9391 250345
rect 9425 249569 9441 250345
rect 9379 249557 9441 249569
rect 9471 250345 9533 250357
rect 9471 249569 9487 250345
rect 9521 249569 9533 250345
rect 9471 249557 9533 249569
rect 9589 250345 9651 250357
rect 9589 249569 9601 250345
rect 9635 249569 9651 250345
rect 9589 249557 9651 249569
rect 9681 250345 9743 250357
rect 9681 249569 9697 250345
rect 9731 249569 9743 250345
rect 9681 249557 9743 249569
rect 9799 250345 9861 250357
rect 9799 249569 9811 250345
rect 9845 249569 9861 250345
rect 9799 249557 9861 249569
rect 9891 250345 9953 250357
rect 9891 249569 9907 250345
rect 9941 249569 9953 250345
rect 9891 249557 9953 249569
rect 10009 250345 10071 250357
rect 10009 249569 10021 250345
rect 10055 249569 10071 250345
rect 10009 249557 10071 249569
rect 10101 250345 10163 250357
rect 10101 249569 10117 250345
rect 10151 249569 10163 250345
rect 10101 249557 10163 249569
rect 10219 250345 10281 250357
rect 10219 249569 10231 250345
rect 10265 249569 10281 250345
rect 10219 249557 10281 249569
rect 10311 250345 10373 250357
rect 10311 249569 10327 250345
rect 10361 249569 10373 250345
rect 10311 249557 10373 249569
rect 10429 250345 10491 250357
rect 10429 249569 10441 250345
rect 10475 249569 10491 250345
rect 10429 249557 10491 249569
rect 10521 250345 10583 250357
rect 10521 249569 10537 250345
rect 10571 249569 10583 250345
rect 10521 249557 10583 249569
rect 10639 250345 10701 250357
rect 10639 249569 10651 250345
rect 10685 249569 10701 250345
rect 10639 249557 10701 249569
rect 10731 250345 10793 250357
rect 10731 249569 10747 250345
rect 10781 249569 10793 250345
rect 10731 249557 10793 249569
rect 10849 250345 10911 250357
rect 10849 249569 10861 250345
rect 10895 249569 10911 250345
rect 10849 249557 10911 249569
rect 10941 250345 11003 250357
rect 10941 249569 10957 250345
rect 10991 249569 11003 250345
rect 10941 249557 11003 249569
rect 11059 250345 11121 250357
rect 11059 249569 11071 250345
rect 11105 249569 11121 250345
rect 11059 249557 11121 249569
rect 11151 250345 11213 250357
rect 11151 249569 11167 250345
rect 11201 249569 11213 250345
rect 11151 249557 11213 249569
rect 11269 250345 11331 250357
rect 11269 249569 11281 250345
rect 11315 249569 11331 250345
rect 11269 249557 11331 249569
rect 11361 250345 11423 250357
rect 11361 249569 11377 250345
rect 11411 249569 11423 250345
rect 11361 249557 11423 249569
rect 11479 250345 11541 250357
rect 11479 249569 11491 250345
rect 11525 249569 11541 250345
rect 11479 249557 11541 249569
rect 11571 250345 11633 250357
rect 11571 249569 11587 250345
rect 11621 249569 11633 250345
rect 11571 249557 11633 249569
rect 11689 250345 11751 250357
rect 11689 249569 11701 250345
rect 11735 249569 11751 250345
rect 11689 249557 11751 249569
rect 11781 250345 11843 250357
rect 11781 249569 11797 250345
rect 11831 249569 11843 250345
rect 11781 249557 11843 249569
rect 11899 250345 11961 250357
rect 11899 249569 11911 250345
rect 11945 249569 11961 250345
rect 11899 249557 11961 249569
rect 11991 250345 12053 250357
rect 11991 249569 12007 250345
rect 12041 249569 12053 250345
rect 11991 249557 12053 249569
rect 12109 250345 12171 250357
rect 12109 249569 12121 250345
rect 12155 249569 12171 250345
rect 12109 249557 12171 249569
rect 12201 250345 12263 250357
rect 12201 249569 12217 250345
rect 12251 249569 12263 250345
rect 12201 249557 12263 249569
rect 12319 250345 12381 250357
rect 12319 249569 12331 250345
rect 12365 249569 12381 250345
rect 12319 249557 12381 249569
rect 12411 250345 12473 250357
rect 12411 249569 12427 250345
rect 12461 249569 12473 250345
rect 12411 249557 12473 249569
rect 12529 250345 12591 250357
rect 12529 249569 12541 250345
rect 12575 249569 12591 250345
rect 12529 249557 12591 249569
rect 12621 250345 12683 250357
rect 12621 249569 12637 250345
rect 12671 249569 12683 250345
rect 12621 249557 12683 249569
rect 12739 250345 12801 250357
rect 12739 249569 12751 250345
rect 12785 249569 12801 250345
rect 12739 249557 12801 249569
rect 12831 250345 12893 250357
rect 12831 249569 12847 250345
rect 12881 249569 12893 250345
rect 12831 249557 12893 249569
rect 12949 250345 13011 250357
rect 12949 249569 12961 250345
rect 12995 249569 13011 250345
rect 12949 249557 13011 249569
rect 13041 250345 13103 250357
rect 13041 249569 13057 250345
rect 13091 249569 13103 250345
rect 13041 249557 13103 249569
rect 13159 250345 13221 250357
rect 13159 249569 13171 250345
rect 13205 249569 13221 250345
rect 13159 249557 13221 249569
rect 13251 250345 13313 250357
rect 13251 249569 13267 250345
rect 13301 249569 13313 250345
rect 13251 249557 13313 249569
rect 13369 250345 13431 250357
rect 13369 249569 13381 250345
rect 13415 249569 13431 250345
rect 13369 249557 13431 249569
rect 13461 250345 13523 250357
rect 13461 249569 13477 250345
rect 13511 249569 13523 250345
rect 13461 249557 13523 249569
rect 13579 250345 13641 250357
rect 13579 249569 13591 250345
rect 13625 249569 13641 250345
rect 13579 249557 13641 249569
rect 13671 250345 13733 250357
rect 13671 249569 13687 250345
rect 13721 249569 13733 250345
rect 13671 249557 13733 249569
rect 13789 250345 13851 250357
rect 13789 249569 13801 250345
rect 13835 249569 13851 250345
rect 13789 249557 13851 249569
rect 13881 250345 13943 250357
rect 13881 249569 13897 250345
rect 13931 249569 13943 250345
rect 13881 249557 13943 249569
rect 13999 250345 14061 250357
rect 13999 249569 14011 250345
rect 14045 249569 14061 250345
rect 13999 249557 14061 249569
rect 14091 250345 14153 250357
rect 14091 249569 14107 250345
rect 14141 249569 14153 250345
rect 14091 249557 14153 249569
rect 14209 250345 14271 250357
rect 14209 249569 14221 250345
rect 14255 249569 14271 250345
rect 14209 249557 14271 249569
rect 14301 250345 14363 250357
rect 14301 249569 14317 250345
rect 14351 249569 14363 250345
rect 14301 249557 14363 249569
rect 14419 250345 14481 250357
rect 14419 249569 14431 250345
rect 14465 249569 14481 250345
rect 14419 249557 14481 249569
rect 14511 250345 14573 250357
rect 14511 249569 14527 250345
rect 14561 249569 14573 250345
rect 14511 249557 14573 249569
rect 14629 250345 14691 250357
rect 14629 249569 14641 250345
rect 14675 249569 14691 250345
rect 14629 249557 14691 249569
rect 14721 250345 14783 250357
rect 14721 249569 14737 250345
rect 14771 249569 14783 250345
rect 14721 249557 14783 249569
rect 14839 250345 14901 250357
rect 14839 249569 14851 250345
rect 14885 249569 14901 250345
rect 14839 249557 14901 249569
rect 14931 250345 14993 250357
rect 14931 249569 14947 250345
rect 14981 249569 14993 250345
rect 14931 249557 14993 249569
rect 15049 250345 15111 250357
rect 15049 249569 15061 250345
rect 15095 249569 15111 250345
rect 15049 249557 15111 249569
rect 15141 250345 15203 250357
rect 15141 249569 15157 250345
rect 15191 249569 15203 250345
rect 15141 249557 15203 249569
rect 15259 250345 15321 250357
rect 15259 249569 15271 250345
rect 15305 249569 15321 250345
rect 15259 249557 15321 249569
rect 15351 250345 15413 250357
rect 15351 249569 15367 250345
rect 15401 249569 15413 250345
rect 15351 249557 15413 249569
rect 15469 250345 15531 250357
rect 15469 249569 15481 250345
rect 15515 249569 15531 250345
rect 15469 249557 15531 249569
rect 15561 250345 15623 250357
rect 15561 249569 15577 250345
rect 15611 249569 15623 250345
rect 15561 249557 15623 249569
rect 15679 250345 15741 250357
rect 15679 249569 15691 250345
rect 15725 249569 15741 250345
rect 15679 249557 15741 249569
rect 15771 250345 15833 250357
rect 15771 249569 15787 250345
rect 15821 249569 15833 250345
rect 15771 249557 15833 249569
rect 15889 250345 15951 250357
rect 15889 249569 15901 250345
rect 15935 249569 15951 250345
rect 15889 249557 15951 249569
rect 15981 250345 16043 250357
rect 15981 249569 15997 250345
rect 16031 249569 16043 250345
rect 15981 249557 16043 249569
rect 16099 250345 16161 250357
rect 16099 249569 16111 250345
rect 16145 249569 16161 250345
rect 16099 249557 16161 249569
rect 16191 250345 16253 250357
rect 16191 249569 16207 250345
rect 16241 249569 16253 250345
rect 16191 249557 16253 249569
rect 16309 250345 16371 250357
rect 16309 249569 16321 250345
rect 16355 249569 16371 250345
rect 16309 249557 16371 249569
rect 16401 250345 16463 250357
rect 16401 249569 16417 250345
rect 16451 249569 16463 250345
rect 16401 249557 16463 249569
rect 16519 250345 16581 250357
rect 16519 249569 16531 250345
rect 16565 249569 16581 250345
rect 16519 249557 16581 249569
rect 16611 250345 16673 250357
rect 16611 249569 16627 250345
rect 16661 249569 16673 250345
rect 16611 249557 16673 249569
rect 16729 250345 16791 250357
rect 16729 249569 16741 250345
rect 16775 249569 16791 250345
rect 16729 249557 16791 249569
rect 16821 250345 16883 250357
rect 16821 249569 16837 250345
rect 16871 249569 16883 250345
rect 16821 249557 16883 249569
rect 16939 250345 17001 250357
rect 16939 249569 16951 250345
rect 16985 249569 17001 250345
rect 16939 249557 17001 249569
rect 17031 250345 17093 250357
rect 17031 249569 17047 250345
rect 17081 249569 17093 250345
rect 17031 249557 17093 249569
rect 17149 250345 17211 250357
rect 17149 249569 17161 250345
rect 17195 249569 17211 250345
rect 17149 249557 17211 249569
rect 17241 250345 17303 250357
rect 17241 249569 17257 250345
rect 17291 249569 17303 250345
rect 17241 249557 17303 249569
rect 17359 250345 17421 250357
rect 17359 249569 17371 250345
rect 17405 249569 17421 250345
rect 17359 249557 17421 249569
rect 17451 250345 17513 250357
rect 17451 249569 17467 250345
rect 17501 249569 17513 250345
rect 17451 249557 17513 249569
rect 17569 250345 17631 250357
rect 17569 249569 17581 250345
rect 17615 249569 17631 250345
rect 17569 249557 17631 249569
rect 17661 250345 17723 250357
rect 17661 249569 17677 250345
rect 17711 249569 17723 250345
rect 17661 249557 17723 249569
rect 17779 250345 17841 250357
rect 17779 249569 17791 250345
rect 17825 249569 17841 250345
rect 17779 249557 17841 249569
rect 17871 250345 17933 250357
rect 17871 249569 17887 250345
rect 17921 249569 17933 250345
rect 17871 249557 17933 249569
rect 17989 250345 18051 250357
rect 17989 249569 18001 250345
rect 18035 249569 18051 250345
rect 17989 249557 18051 249569
rect 18081 250345 18143 250357
rect 18081 249569 18097 250345
rect 18131 249569 18143 250345
rect 18081 249557 18143 249569
rect 18199 250345 18261 250357
rect 18199 249569 18211 250345
rect 18245 249569 18261 250345
rect 18199 249557 18261 249569
rect 18291 250345 18353 250357
rect 18291 249569 18307 250345
rect 18341 249569 18353 250345
rect 18291 249557 18353 249569
rect 18409 250345 18471 250357
rect 18409 249569 18421 250345
rect 18455 249569 18471 250345
rect 18409 249557 18471 249569
rect 18501 250345 18563 250357
rect 18501 249569 18517 250345
rect 18551 249569 18563 250345
rect 18501 249557 18563 249569
rect 18619 250345 18681 250357
rect 18619 249569 18631 250345
rect 18665 249569 18681 250345
rect 18619 249557 18681 249569
rect 18711 250345 18773 250357
rect 18711 249569 18727 250345
rect 18761 249569 18773 250345
rect 18711 249557 18773 249569
rect 18829 250345 18891 250357
rect 18829 249569 18841 250345
rect 18875 249569 18891 250345
rect 18829 249557 18891 249569
rect 18921 250345 18983 250357
rect 18921 249569 18937 250345
rect 18971 249569 18983 250345
rect 18921 249557 18983 249569
rect 19039 250345 19101 250357
rect 19039 249569 19051 250345
rect 19085 249569 19101 250345
rect 19039 249557 19101 249569
rect 19131 250345 19193 250357
rect 19131 249569 19147 250345
rect 19181 249569 19193 250345
rect 19131 249557 19193 249569
rect 19249 250345 19311 250357
rect 19249 249569 19261 250345
rect 19295 249569 19311 250345
rect 19249 249557 19311 249569
rect 19341 250345 19403 250357
rect 19341 249569 19357 250345
rect 19391 249569 19403 250345
rect 19341 249557 19403 249569
rect 19459 250345 19521 250357
rect 19459 249569 19471 250345
rect 19505 249569 19521 250345
rect 19459 249557 19521 249569
rect 19551 250345 19613 250357
rect 19551 249569 19567 250345
rect 19601 249569 19613 250345
rect 19551 249557 19613 249569
rect 19669 250345 19731 250357
rect 19669 249569 19681 250345
rect 19715 249569 19731 250345
rect 19669 249557 19731 249569
rect 19761 250345 19823 250357
rect 19761 249569 19777 250345
rect 19811 249569 19823 250345
rect 19761 249557 19823 249569
rect 19879 250345 19941 250357
rect 19879 249569 19891 250345
rect 19925 249569 19941 250345
rect 19879 249557 19941 249569
rect 19971 250345 20033 250357
rect 19971 249569 19987 250345
rect 20021 249569 20033 250345
rect 19971 249557 20033 249569
rect 20089 250345 20151 250357
rect 20089 249569 20101 250345
rect 20135 249569 20151 250345
rect 20089 249557 20151 249569
rect 20181 250345 20243 250357
rect 20181 249569 20197 250345
rect 20231 249569 20243 250345
rect 20181 249557 20243 249569
rect 20299 250345 20361 250357
rect 20299 249569 20311 250345
rect 20345 249569 20361 250345
rect 20299 249557 20361 249569
rect 20391 250345 20453 250357
rect 20391 249569 20407 250345
rect 20441 249569 20453 250345
rect 20391 249557 20453 249569
rect 20509 250345 20571 250357
rect 20509 249569 20521 250345
rect 20555 249569 20571 250345
rect 20509 249557 20571 249569
rect 20601 250345 20663 250357
rect 20601 249569 20617 250345
rect 20651 249569 20663 250345
rect 20601 249557 20663 249569
rect 20719 250345 20781 250357
rect 20719 249569 20731 250345
rect 20765 249569 20781 250345
rect 20719 249557 20781 249569
rect 20811 250345 20873 250357
rect 20811 249569 20827 250345
rect 20861 249569 20873 250345
rect 20811 249557 20873 249569
rect 20929 250345 20991 250357
rect 20929 249569 20941 250345
rect 20975 249569 20991 250345
rect 20929 249557 20991 249569
rect 21021 250345 21083 250357
rect 21021 249569 21037 250345
rect 21071 249569 21083 250345
rect 21021 249557 21083 249569
rect 21139 250345 21201 250357
rect 21139 249569 21151 250345
rect 21185 249569 21201 250345
rect 21139 249557 21201 249569
rect 21231 250345 21293 250357
rect 21231 249569 21247 250345
rect 21281 249569 21293 250345
rect 21231 249557 21293 249569
rect 21349 250345 21411 250357
rect 21349 249569 21361 250345
rect 21395 249569 21411 250345
rect 21349 249557 21411 249569
rect 21441 250345 21503 250357
rect 21441 249569 21457 250345
rect 21491 249569 21503 250345
rect 21441 249557 21503 249569
rect 21559 250345 21621 250357
rect 21559 249569 21571 250345
rect 21605 249569 21621 250345
rect 21559 249557 21621 249569
rect 21651 250345 21713 250357
rect 21651 249569 21667 250345
rect 21701 249569 21713 250345
rect 21651 249557 21713 249569
rect 21769 250345 21831 250357
rect 21769 249569 21781 250345
rect 21815 249569 21831 250345
rect 21769 249557 21831 249569
rect 21861 250345 21923 250357
rect 21861 249569 21877 250345
rect 21911 249569 21923 250345
rect 21861 249557 21923 249569
rect 21979 250345 22041 250357
rect 21979 249569 21991 250345
rect 22025 249569 22041 250345
rect 21979 249557 22041 249569
rect 22071 250345 22133 250357
rect 22071 249569 22087 250345
rect 22121 249569 22133 250345
rect 22071 249557 22133 249569
rect 22189 250345 22251 250357
rect 22189 249569 22201 250345
rect 22235 249569 22251 250345
rect 22189 249557 22251 249569
rect 22281 250345 22343 250357
rect 22281 249569 22297 250345
rect 22331 249569 22343 250345
rect 22281 249557 22343 249569
rect 22399 250345 22461 250357
rect 22399 249569 22411 250345
rect 22445 249569 22461 250345
rect 22399 249557 22461 249569
rect 22491 250345 22553 250357
rect 22491 249569 22507 250345
rect 22541 249569 22553 250345
rect 22491 249557 22553 249569
rect 22609 250345 22671 250357
rect 22609 249569 22621 250345
rect 22655 249569 22671 250345
rect 22609 249557 22671 249569
rect 22701 250345 22763 250357
rect 22701 249569 22717 250345
rect 22751 249569 22763 250345
rect 22701 249557 22763 249569
rect 22819 250345 22881 250357
rect 22819 249569 22831 250345
rect 22865 249569 22881 250345
rect 22819 249557 22881 249569
rect 22911 250345 22973 250357
rect 22911 249569 22927 250345
rect 22961 249569 22973 250345
rect 22911 249557 22973 249569
rect 23029 250345 23091 250357
rect 23029 249569 23041 250345
rect 23075 249569 23091 250345
rect 23029 249557 23091 249569
rect 23121 250345 23183 250357
rect 23121 249569 23137 250345
rect 23171 249569 23183 250345
rect 23121 249557 23183 249569
rect 23239 250345 23301 250357
rect 23239 249569 23251 250345
rect 23285 249569 23301 250345
rect 23239 249557 23301 249569
rect 23331 250345 23393 250357
rect 23331 249569 23347 250345
rect 23381 249569 23393 250345
rect 23331 249557 23393 249569
rect 23449 250345 23511 250357
rect 23449 249569 23461 250345
rect 23495 249569 23511 250345
rect 23449 249557 23511 249569
rect 23541 250345 23603 250357
rect 23541 249569 23557 250345
rect 23591 249569 23603 250345
rect 23541 249557 23603 249569
rect 23659 250345 23721 250357
rect 23659 249569 23671 250345
rect 23705 249569 23721 250345
rect 23659 249557 23721 249569
rect 23751 250345 23813 250357
rect 23751 249569 23767 250345
rect 23801 249569 23813 250345
rect 23751 249557 23813 249569
rect 23869 250345 23931 250357
rect 23869 249569 23881 250345
rect 23915 249569 23931 250345
rect 23869 249557 23931 249569
rect 23961 250345 24023 250357
rect 23961 249569 23977 250345
rect 24011 249569 24023 250345
rect 23961 249557 24023 249569
rect 24079 250345 24141 250357
rect 24079 249569 24091 250345
rect 24125 249569 24141 250345
rect 24079 249557 24141 249569
rect 24171 250345 24233 250357
rect 24171 249569 24187 250345
rect 24221 249569 24233 250345
rect 24171 249557 24233 249569
rect 24289 250345 24351 250357
rect 24289 249569 24301 250345
rect 24335 249569 24351 250345
rect 24289 249557 24351 249569
rect 24381 250345 24443 250357
rect 24381 249569 24397 250345
rect 24431 249569 24443 250345
rect 24381 249557 24443 249569
rect 24499 250345 24561 250357
rect 24499 249569 24511 250345
rect 24545 249569 24561 250345
rect 24499 249557 24561 249569
rect 24591 250345 24653 250357
rect 24591 249569 24607 250345
rect 24641 249569 24653 250345
rect 24591 249557 24653 249569
rect 24709 250345 24771 250357
rect 24709 249569 24721 250345
rect 24755 249569 24771 250345
rect 24709 249557 24771 249569
rect 24801 250345 24863 250357
rect 24801 249569 24817 250345
rect 24851 249569 24863 250345
rect 24801 249557 24863 249569
rect 24919 250345 24981 250357
rect 24919 249569 24931 250345
rect 24965 249569 24981 250345
rect 24919 249557 24981 249569
rect 25011 250345 25073 250357
rect 25011 249569 25027 250345
rect 25061 249569 25073 250345
rect 25011 249557 25073 249569
rect 25129 250345 25191 250357
rect 25129 249569 25141 250345
rect 25175 249569 25191 250345
rect 25129 249557 25191 249569
rect 25221 250345 25283 250357
rect 25221 249569 25237 250345
rect 25271 249569 25283 250345
rect 25221 249557 25283 249569
rect 25339 250345 25401 250357
rect 25339 249569 25351 250345
rect 25385 249569 25401 250345
rect 25339 249557 25401 249569
rect 25431 250345 25493 250357
rect 25431 249569 25447 250345
rect 25481 249569 25493 250345
rect 25431 249557 25493 249569
rect 25549 250345 25611 250357
rect 25549 249569 25561 250345
rect 25595 249569 25611 250345
rect 25549 249557 25611 249569
rect 25641 250345 25703 250357
rect 25641 249569 25657 250345
rect 25691 249569 25703 250345
rect 25641 249557 25703 249569
rect 25759 250345 25821 250357
rect 25759 249569 25771 250345
rect 25805 249569 25821 250345
rect 25759 249557 25821 249569
rect 25851 250345 25913 250357
rect 25851 249569 25867 250345
rect 25901 249569 25913 250345
rect 25851 249557 25913 249569
rect 25969 250345 26031 250357
rect 25969 249569 25981 250345
rect 26015 249569 26031 250345
rect 25969 249557 26031 249569
rect 26061 250345 26123 250357
rect 26061 249569 26077 250345
rect 26111 249569 26123 250345
rect 26061 249557 26123 249569
rect 26179 250345 26241 250357
rect 26179 249569 26191 250345
rect 26225 249569 26241 250345
rect 26179 249557 26241 249569
rect 26271 250345 26333 250357
rect 26271 249569 26287 250345
rect 26321 249569 26333 250345
rect 26271 249557 26333 249569
rect 26389 250345 26451 250357
rect 26389 249569 26401 250345
rect 26435 249569 26451 250345
rect 26389 249557 26451 249569
rect 26481 250345 26543 250357
rect 26481 249569 26497 250345
rect 26531 249569 26543 250345
rect 26481 249557 26543 249569
rect 26599 250345 26661 250357
rect 26599 249569 26611 250345
rect 26645 249569 26661 250345
rect 26599 249557 26661 249569
rect 26691 250345 26753 250357
rect 26691 249569 26707 250345
rect 26741 249569 26753 250345
rect 26691 249557 26753 249569
rect 26809 250345 26871 250357
rect 26809 249569 26821 250345
rect 26855 249569 26871 250345
rect 26809 249557 26871 249569
rect 26901 250345 26963 250357
rect 26901 249569 26917 250345
rect 26951 249569 26963 250345
rect 26901 249557 26963 249569
rect 27019 250345 27081 250357
rect 27019 249569 27031 250345
rect 27065 249569 27081 250345
rect 27019 249557 27081 249569
rect 27111 250345 27173 250357
rect 27111 249569 27127 250345
rect 27161 249569 27173 250345
rect 27111 249557 27173 249569
rect 27229 250345 27291 250357
rect 27229 249569 27241 250345
rect 27275 249569 27291 250345
rect 27229 249557 27291 249569
rect 27321 250345 27383 250357
rect 27321 249569 27337 250345
rect 27371 249569 27383 250345
rect 27321 249557 27383 249569
rect -4061 249180 -3999 249192
rect -4061 248404 -4049 249180
rect -4015 248404 -3999 249180
rect -4061 248392 -3999 248404
rect -3969 249180 -3907 249192
rect -3969 248404 -3953 249180
rect -3919 248404 -3907 249180
rect -3969 248392 -3907 248404
rect -3851 249180 -3789 249192
rect -3851 248404 -3839 249180
rect -3805 248404 -3789 249180
rect -3851 248392 -3789 248404
rect -3759 249180 -3697 249192
rect -3759 248404 -3743 249180
rect -3709 248404 -3697 249180
rect -3759 248392 -3697 248404
rect -3641 249180 -3579 249192
rect -3641 248404 -3629 249180
rect -3595 248404 -3579 249180
rect -3641 248392 -3579 248404
rect -3549 249180 -3487 249192
rect -3549 248404 -3533 249180
rect -3499 248404 -3487 249180
rect -3549 248392 -3487 248404
rect -3431 249180 -3369 249192
rect -3431 248404 -3419 249180
rect -3385 248404 -3369 249180
rect -3431 248392 -3369 248404
rect -3339 249180 -3277 249192
rect -3339 248404 -3323 249180
rect -3289 248404 -3277 249180
rect -3339 248392 -3277 248404
rect -3221 249180 -3159 249192
rect -3221 248404 -3209 249180
rect -3175 248404 -3159 249180
rect -3221 248392 -3159 248404
rect -3129 249180 -3067 249192
rect -3129 248404 -3113 249180
rect -3079 248404 -3067 249180
rect -3129 248392 -3067 248404
rect -3011 249180 -2949 249192
rect -3011 248404 -2999 249180
rect -2965 248404 -2949 249180
rect -3011 248392 -2949 248404
rect -2919 249180 -2857 249192
rect -2919 248404 -2903 249180
rect -2869 248404 -2857 249180
rect -2919 248392 -2857 248404
rect -2801 249180 -2739 249192
rect -2801 248404 -2789 249180
rect -2755 248404 -2739 249180
rect -2801 248392 -2739 248404
rect -2709 249180 -2647 249192
rect -2709 248404 -2693 249180
rect -2659 248404 -2647 249180
rect -2709 248392 -2647 248404
rect -2591 249180 -2529 249192
rect -2591 248404 -2579 249180
rect -2545 248404 -2529 249180
rect -2591 248392 -2529 248404
rect -2499 249180 -2437 249192
rect -2499 248404 -2483 249180
rect -2449 248404 -2437 249180
rect -2499 248392 -2437 248404
rect -2381 249180 -2319 249192
rect -2381 248404 -2369 249180
rect -2335 248404 -2319 249180
rect -2381 248392 -2319 248404
rect -2289 249180 -2227 249192
rect -2289 248404 -2273 249180
rect -2239 248404 -2227 249180
rect -2289 248392 -2227 248404
rect -2171 249180 -2109 249192
rect -2171 248404 -2159 249180
rect -2125 248404 -2109 249180
rect -2171 248392 -2109 248404
rect -2079 249180 -2017 249192
rect -2079 248404 -2063 249180
rect -2029 248404 -2017 249180
rect -2079 248392 -2017 248404
rect -1961 249180 -1899 249192
rect -1961 248404 -1949 249180
rect -1915 248404 -1899 249180
rect -1961 248392 -1899 248404
rect -1869 249180 -1807 249192
rect -1869 248404 -1853 249180
rect -1819 248404 -1807 249180
rect -1869 248392 -1807 248404
rect -1751 249180 -1689 249192
rect -1751 248404 -1739 249180
rect -1705 248404 -1689 249180
rect -1751 248392 -1689 248404
rect -1659 249180 -1597 249192
rect -1659 248404 -1643 249180
rect -1609 248404 -1597 249180
rect -1659 248392 -1597 248404
rect -1541 249180 -1479 249192
rect -1541 248404 -1529 249180
rect -1495 248404 -1479 249180
rect -1541 248392 -1479 248404
rect -1449 249180 -1387 249192
rect -1449 248404 -1433 249180
rect -1399 248404 -1387 249180
rect -1449 248392 -1387 248404
rect -1331 249180 -1269 249192
rect -1331 248404 -1319 249180
rect -1285 248404 -1269 249180
rect -1331 248392 -1269 248404
rect -1239 249180 -1177 249192
rect -1239 248404 -1223 249180
rect -1189 248404 -1177 249180
rect -1239 248392 -1177 248404
rect -1121 249180 -1059 249192
rect -1121 248404 -1109 249180
rect -1075 248404 -1059 249180
rect -1121 248392 -1059 248404
rect -1029 249180 -967 249192
rect -1029 248404 -1013 249180
rect -979 248404 -967 249180
rect -1029 248392 -967 248404
rect -911 249180 -849 249192
rect -911 248404 -899 249180
rect -865 248404 -849 249180
rect -911 248392 -849 248404
rect -819 249180 -757 249192
rect -819 248404 -803 249180
rect -769 248404 -757 249180
rect -819 248392 -757 248404
rect -701 249180 -639 249192
rect -701 248404 -689 249180
rect -655 248404 -639 249180
rect -701 248392 -639 248404
rect -609 249180 -547 249192
rect -609 248404 -593 249180
rect -559 248404 -547 249180
rect -609 248392 -547 248404
rect -491 249180 -429 249192
rect -491 248404 -479 249180
rect -445 248404 -429 249180
rect -491 248392 -429 248404
rect -399 249180 -337 249192
rect -399 248404 -383 249180
rect -349 248404 -337 249180
rect -399 248392 -337 248404
rect -281 249180 -219 249192
rect -281 248404 -269 249180
rect -235 248404 -219 249180
rect -281 248392 -219 248404
rect -189 249180 -127 249192
rect -189 248404 -173 249180
rect -139 248404 -127 249180
rect -189 248392 -127 248404
rect -71 249180 -9 249192
rect -71 248404 -59 249180
rect -25 248404 -9 249180
rect -71 248392 -9 248404
rect 21 249180 83 249192
rect 21 248404 37 249180
rect 71 248404 83 249180
rect 21 248392 83 248404
rect 139 249180 201 249192
rect 139 248404 151 249180
rect 185 248404 201 249180
rect 139 248392 201 248404
rect 231 249180 293 249192
rect 231 248404 247 249180
rect 281 248404 293 249180
rect 231 248392 293 248404
rect 349 249180 411 249192
rect 349 248404 361 249180
rect 395 248404 411 249180
rect 349 248392 411 248404
rect 441 249180 503 249192
rect 441 248404 457 249180
rect 491 248404 503 249180
rect 441 248392 503 248404
rect 559 249180 621 249192
rect 559 248404 571 249180
rect 605 248404 621 249180
rect 559 248392 621 248404
rect 651 249180 713 249192
rect 651 248404 667 249180
rect 701 248404 713 249180
rect 651 248392 713 248404
rect 769 249180 831 249192
rect 769 248404 781 249180
rect 815 248404 831 249180
rect 769 248392 831 248404
rect 861 249180 923 249192
rect 861 248404 877 249180
rect 911 248404 923 249180
rect 861 248392 923 248404
rect 979 249180 1041 249192
rect 979 248404 991 249180
rect 1025 248404 1041 249180
rect 979 248392 1041 248404
rect 1071 249180 1133 249192
rect 1071 248404 1087 249180
rect 1121 248404 1133 249180
rect 1071 248392 1133 248404
rect 1189 249180 1251 249192
rect 1189 248404 1201 249180
rect 1235 248404 1251 249180
rect 1189 248392 1251 248404
rect 1281 249180 1343 249192
rect 1281 248404 1297 249180
rect 1331 248404 1343 249180
rect 1281 248392 1343 248404
rect 1399 249180 1461 249192
rect 1399 248404 1411 249180
rect 1445 248404 1461 249180
rect 1399 248392 1461 248404
rect 1491 249180 1553 249192
rect 1491 248404 1507 249180
rect 1541 248404 1553 249180
rect 1491 248392 1553 248404
rect 1609 249180 1671 249192
rect 1609 248404 1621 249180
rect 1655 248404 1671 249180
rect 1609 248392 1671 248404
rect 1701 249180 1763 249192
rect 1701 248404 1717 249180
rect 1751 248404 1763 249180
rect 1701 248392 1763 248404
rect 1819 249180 1881 249192
rect 1819 248404 1831 249180
rect 1865 248404 1881 249180
rect 1819 248392 1881 248404
rect 1911 249180 1973 249192
rect 1911 248404 1927 249180
rect 1961 248404 1973 249180
rect 1911 248392 1973 248404
rect 2029 249180 2091 249192
rect 2029 248404 2041 249180
rect 2075 248404 2091 249180
rect 2029 248392 2091 248404
rect 2121 249180 2183 249192
rect 2121 248404 2137 249180
rect 2171 248404 2183 249180
rect 2121 248392 2183 248404
rect 2239 249180 2301 249192
rect 2239 248404 2251 249180
rect 2285 248404 2301 249180
rect 2239 248392 2301 248404
rect 2331 249180 2393 249192
rect 2331 248404 2347 249180
rect 2381 248404 2393 249180
rect 2331 248392 2393 248404
rect 2449 249180 2511 249192
rect 2449 248404 2461 249180
rect 2495 248404 2511 249180
rect 2449 248392 2511 248404
rect 2541 249180 2603 249192
rect 2541 248404 2557 249180
rect 2591 248404 2603 249180
rect 2541 248392 2603 248404
rect 2659 249180 2721 249192
rect 2659 248404 2671 249180
rect 2705 248404 2721 249180
rect 2659 248392 2721 248404
rect 2751 249180 2813 249192
rect 2751 248404 2767 249180
rect 2801 248404 2813 249180
rect 2751 248392 2813 248404
rect 2869 249180 2931 249192
rect 2869 248404 2881 249180
rect 2915 248404 2931 249180
rect 2869 248392 2931 248404
rect 2961 249180 3023 249192
rect 2961 248404 2977 249180
rect 3011 248404 3023 249180
rect 2961 248392 3023 248404
rect 3079 249180 3141 249192
rect 3079 248404 3091 249180
rect 3125 248404 3141 249180
rect 3079 248392 3141 248404
rect 3171 249180 3233 249192
rect 3171 248404 3187 249180
rect 3221 248404 3233 249180
rect 3171 248392 3233 248404
rect 3289 249180 3351 249192
rect 3289 248404 3301 249180
rect 3335 248404 3351 249180
rect 3289 248392 3351 248404
rect 3381 249180 3443 249192
rect 3381 248404 3397 249180
rect 3431 248404 3443 249180
rect 3381 248392 3443 248404
rect 3499 249180 3561 249192
rect 3499 248404 3511 249180
rect 3545 248404 3561 249180
rect 3499 248392 3561 248404
rect 3591 249180 3653 249192
rect 3591 248404 3607 249180
rect 3641 248404 3653 249180
rect 3591 248392 3653 248404
rect 3709 249180 3771 249192
rect 3709 248404 3721 249180
rect 3755 248404 3771 249180
rect 3709 248392 3771 248404
rect 3801 249180 3863 249192
rect 3801 248404 3817 249180
rect 3851 248404 3863 249180
rect 3801 248392 3863 248404
rect 3919 249180 3981 249192
rect 3919 248404 3931 249180
rect 3965 248404 3981 249180
rect 3919 248392 3981 248404
rect 4011 249180 4073 249192
rect 4011 248404 4027 249180
rect 4061 248404 4073 249180
rect 4011 248392 4073 248404
rect 4129 249180 4191 249192
rect 4129 248404 4141 249180
rect 4175 248404 4191 249180
rect 4129 248392 4191 248404
rect 4221 249180 4283 249192
rect 4221 248404 4237 249180
rect 4271 248404 4283 249180
rect 4221 248392 4283 248404
rect 4339 249180 4401 249192
rect 4339 248404 4351 249180
rect 4385 248404 4401 249180
rect 4339 248392 4401 248404
rect 4431 249180 4493 249192
rect 4431 248404 4447 249180
rect 4481 248404 4493 249180
rect 4431 248392 4493 248404
rect 4549 249180 4611 249192
rect 4549 248404 4561 249180
rect 4595 248404 4611 249180
rect 4549 248392 4611 248404
rect 4641 249180 4703 249192
rect 4641 248404 4657 249180
rect 4691 248404 4703 249180
rect 4641 248392 4703 248404
rect 4759 249180 4821 249192
rect 4759 248404 4771 249180
rect 4805 248404 4821 249180
rect 4759 248392 4821 248404
rect 4851 249180 4913 249192
rect 4851 248404 4867 249180
rect 4901 248404 4913 249180
rect 4851 248392 4913 248404
rect 4969 249180 5031 249192
rect 4969 248404 4981 249180
rect 5015 248404 5031 249180
rect 4969 248392 5031 248404
rect 5061 249180 5123 249192
rect 5061 248404 5077 249180
rect 5111 248404 5123 249180
rect 5061 248392 5123 248404
rect 5179 249180 5241 249192
rect 5179 248404 5191 249180
rect 5225 248404 5241 249180
rect 5179 248392 5241 248404
rect 5271 249180 5333 249192
rect 5271 248404 5287 249180
rect 5321 248404 5333 249180
rect 5271 248392 5333 248404
rect 5389 249180 5451 249192
rect 5389 248404 5401 249180
rect 5435 248404 5451 249180
rect 5389 248392 5451 248404
rect 5481 249180 5543 249192
rect 5481 248404 5497 249180
rect 5531 248404 5543 249180
rect 5481 248392 5543 248404
rect 5599 249180 5661 249192
rect 5599 248404 5611 249180
rect 5645 248404 5661 249180
rect 5599 248392 5661 248404
rect 5691 249180 5753 249192
rect 5691 248404 5707 249180
rect 5741 248404 5753 249180
rect 5691 248392 5753 248404
rect 5809 249180 5871 249192
rect 5809 248404 5821 249180
rect 5855 248404 5871 249180
rect 5809 248392 5871 248404
rect 5901 249180 5963 249192
rect 5901 248404 5917 249180
rect 5951 248404 5963 249180
rect 5901 248392 5963 248404
rect 6019 249180 6081 249192
rect 6019 248404 6031 249180
rect 6065 248404 6081 249180
rect 6019 248392 6081 248404
rect 6111 249180 6173 249192
rect 6111 248404 6127 249180
rect 6161 248404 6173 249180
rect 6111 248392 6173 248404
rect 6229 249180 6291 249192
rect 6229 248404 6241 249180
rect 6275 248404 6291 249180
rect 6229 248392 6291 248404
rect 6321 249180 6383 249192
rect 6321 248404 6337 249180
rect 6371 248404 6383 249180
rect 6321 248392 6383 248404
rect 6439 249180 6501 249192
rect 6439 248404 6451 249180
rect 6485 248404 6501 249180
rect 6439 248392 6501 248404
rect 6531 249180 6593 249192
rect 6531 248404 6547 249180
rect 6581 248404 6593 249180
rect 6531 248392 6593 248404
rect 6649 249180 6711 249192
rect 6649 248404 6661 249180
rect 6695 248404 6711 249180
rect 6649 248392 6711 248404
rect 6741 249180 6803 249192
rect 6741 248404 6757 249180
rect 6791 248404 6803 249180
rect 6741 248392 6803 248404
rect 6859 249180 6921 249192
rect 6859 248404 6871 249180
rect 6905 248404 6921 249180
rect 6859 248392 6921 248404
rect 6951 249180 7013 249192
rect 6951 248404 6967 249180
rect 7001 248404 7013 249180
rect 6951 248392 7013 248404
rect 7069 249180 7131 249192
rect 7069 248404 7081 249180
rect 7115 248404 7131 249180
rect 7069 248392 7131 248404
rect 7161 249180 7223 249192
rect 7161 248404 7177 249180
rect 7211 248404 7223 249180
rect 7161 248392 7223 248404
rect 7279 249180 7341 249192
rect 7279 248404 7291 249180
rect 7325 248404 7341 249180
rect 7279 248392 7341 248404
rect 7371 249180 7433 249192
rect 7371 248404 7387 249180
rect 7421 248404 7433 249180
rect 7371 248392 7433 248404
rect 7489 249180 7551 249192
rect 7489 248404 7501 249180
rect 7535 248404 7551 249180
rect 7489 248392 7551 248404
rect 7581 249180 7643 249192
rect 7581 248404 7597 249180
rect 7631 248404 7643 249180
rect 7581 248392 7643 248404
rect 7699 249180 7761 249192
rect 7699 248404 7711 249180
rect 7745 248404 7761 249180
rect 7699 248392 7761 248404
rect 7791 249180 7853 249192
rect 7791 248404 7807 249180
rect 7841 248404 7853 249180
rect 7791 248392 7853 248404
rect 7909 249180 7971 249192
rect 7909 248404 7921 249180
rect 7955 248404 7971 249180
rect 7909 248392 7971 248404
rect 8001 249180 8063 249192
rect 8001 248404 8017 249180
rect 8051 248404 8063 249180
rect 8001 248392 8063 248404
rect 8119 249180 8181 249192
rect 8119 248404 8131 249180
rect 8165 248404 8181 249180
rect 8119 248392 8181 248404
rect 8211 249180 8273 249192
rect 8211 248404 8227 249180
rect 8261 248404 8273 249180
rect 8211 248392 8273 248404
rect 8329 249180 8391 249192
rect 8329 248404 8341 249180
rect 8375 248404 8391 249180
rect 8329 248392 8391 248404
rect 8421 249180 8483 249192
rect 8421 248404 8437 249180
rect 8471 248404 8483 249180
rect 8421 248392 8483 248404
rect 8539 249180 8601 249192
rect 8539 248404 8551 249180
rect 8585 248404 8601 249180
rect 8539 248392 8601 248404
rect 8631 249180 8693 249192
rect 8631 248404 8647 249180
rect 8681 248404 8693 249180
rect 8631 248392 8693 248404
rect 8749 249180 8811 249192
rect 8749 248404 8761 249180
rect 8795 248404 8811 249180
rect 8749 248392 8811 248404
rect 8841 249180 8903 249192
rect 8841 248404 8857 249180
rect 8891 248404 8903 249180
rect 8841 248392 8903 248404
rect 8959 249180 9021 249192
rect 8959 248404 8971 249180
rect 9005 248404 9021 249180
rect 8959 248392 9021 248404
rect 9051 249180 9113 249192
rect 9051 248404 9067 249180
rect 9101 248404 9113 249180
rect 9051 248392 9113 248404
rect 9169 249180 9231 249192
rect 9169 248404 9181 249180
rect 9215 248404 9231 249180
rect 9169 248392 9231 248404
rect 9261 249180 9323 249192
rect 9261 248404 9277 249180
rect 9311 248404 9323 249180
rect 9261 248392 9323 248404
rect 9379 249180 9441 249192
rect 9379 248404 9391 249180
rect 9425 248404 9441 249180
rect 9379 248392 9441 248404
rect 9471 249180 9533 249192
rect 9471 248404 9487 249180
rect 9521 248404 9533 249180
rect 9471 248392 9533 248404
rect 9589 249180 9651 249192
rect 9589 248404 9601 249180
rect 9635 248404 9651 249180
rect 9589 248392 9651 248404
rect 9681 249180 9743 249192
rect 9681 248404 9697 249180
rect 9731 248404 9743 249180
rect 9681 248392 9743 248404
rect 9799 249180 9861 249192
rect 9799 248404 9811 249180
rect 9845 248404 9861 249180
rect 9799 248392 9861 248404
rect 9891 249180 9953 249192
rect 9891 248404 9907 249180
rect 9941 248404 9953 249180
rect 9891 248392 9953 248404
rect 10009 249180 10071 249192
rect 10009 248404 10021 249180
rect 10055 248404 10071 249180
rect 10009 248392 10071 248404
rect 10101 249180 10163 249192
rect 10101 248404 10117 249180
rect 10151 248404 10163 249180
rect 10101 248392 10163 248404
rect 10219 249180 10281 249192
rect 10219 248404 10231 249180
rect 10265 248404 10281 249180
rect 10219 248392 10281 248404
rect 10311 249180 10373 249192
rect 10311 248404 10327 249180
rect 10361 248404 10373 249180
rect 10311 248392 10373 248404
rect 10429 249180 10491 249192
rect 10429 248404 10441 249180
rect 10475 248404 10491 249180
rect 10429 248392 10491 248404
rect 10521 249180 10583 249192
rect 10521 248404 10537 249180
rect 10571 248404 10583 249180
rect 10521 248392 10583 248404
rect 10639 249180 10701 249192
rect 10639 248404 10651 249180
rect 10685 248404 10701 249180
rect 10639 248392 10701 248404
rect 10731 249180 10793 249192
rect 10731 248404 10747 249180
rect 10781 248404 10793 249180
rect 10731 248392 10793 248404
rect 10849 249180 10911 249192
rect 10849 248404 10861 249180
rect 10895 248404 10911 249180
rect 10849 248392 10911 248404
rect 10941 249180 11003 249192
rect 10941 248404 10957 249180
rect 10991 248404 11003 249180
rect 10941 248392 11003 248404
rect 11059 249180 11121 249192
rect 11059 248404 11071 249180
rect 11105 248404 11121 249180
rect 11059 248392 11121 248404
rect 11151 249180 11213 249192
rect 11151 248404 11167 249180
rect 11201 248404 11213 249180
rect 11151 248392 11213 248404
rect 11269 249180 11331 249192
rect 11269 248404 11281 249180
rect 11315 248404 11331 249180
rect 11269 248392 11331 248404
rect 11361 249180 11423 249192
rect 11361 248404 11377 249180
rect 11411 248404 11423 249180
rect 11361 248392 11423 248404
rect 11479 249180 11541 249192
rect 11479 248404 11491 249180
rect 11525 248404 11541 249180
rect 11479 248392 11541 248404
rect 11571 249180 11633 249192
rect 11571 248404 11587 249180
rect 11621 248404 11633 249180
rect 11571 248392 11633 248404
rect 11689 249180 11751 249192
rect 11689 248404 11701 249180
rect 11735 248404 11751 249180
rect 11689 248392 11751 248404
rect 11781 249180 11843 249192
rect 11781 248404 11797 249180
rect 11831 248404 11843 249180
rect 11781 248392 11843 248404
rect 11899 249180 11961 249192
rect 11899 248404 11911 249180
rect 11945 248404 11961 249180
rect 11899 248392 11961 248404
rect 11991 249180 12053 249192
rect 11991 248404 12007 249180
rect 12041 248404 12053 249180
rect 11991 248392 12053 248404
rect 12109 249180 12171 249192
rect 12109 248404 12121 249180
rect 12155 248404 12171 249180
rect 12109 248392 12171 248404
rect 12201 249180 12263 249192
rect 12201 248404 12217 249180
rect 12251 248404 12263 249180
rect 12201 248392 12263 248404
rect 12319 249180 12381 249192
rect 12319 248404 12331 249180
rect 12365 248404 12381 249180
rect 12319 248392 12381 248404
rect 12411 249180 12473 249192
rect 12411 248404 12427 249180
rect 12461 248404 12473 249180
rect 12411 248392 12473 248404
rect 12529 249180 12591 249192
rect 12529 248404 12541 249180
rect 12575 248404 12591 249180
rect 12529 248392 12591 248404
rect 12621 249180 12683 249192
rect 12621 248404 12637 249180
rect 12671 248404 12683 249180
rect 12621 248392 12683 248404
rect 12739 249180 12801 249192
rect 12739 248404 12751 249180
rect 12785 248404 12801 249180
rect 12739 248392 12801 248404
rect 12831 249180 12893 249192
rect 12831 248404 12847 249180
rect 12881 248404 12893 249180
rect 12831 248392 12893 248404
rect 12949 249180 13011 249192
rect 12949 248404 12961 249180
rect 12995 248404 13011 249180
rect 12949 248392 13011 248404
rect 13041 249180 13103 249192
rect 13041 248404 13057 249180
rect 13091 248404 13103 249180
rect 13041 248392 13103 248404
rect 13159 249180 13221 249192
rect 13159 248404 13171 249180
rect 13205 248404 13221 249180
rect 13159 248392 13221 248404
rect 13251 249180 13313 249192
rect 13251 248404 13267 249180
rect 13301 248404 13313 249180
rect 13251 248392 13313 248404
rect 13369 249180 13431 249192
rect 13369 248404 13381 249180
rect 13415 248404 13431 249180
rect 13369 248392 13431 248404
rect 13461 249180 13523 249192
rect 13461 248404 13477 249180
rect 13511 248404 13523 249180
rect 13461 248392 13523 248404
rect 13579 249180 13641 249192
rect 13579 248404 13591 249180
rect 13625 248404 13641 249180
rect 13579 248392 13641 248404
rect 13671 249180 13733 249192
rect 13671 248404 13687 249180
rect 13721 248404 13733 249180
rect 13671 248392 13733 248404
rect 13789 249180 13851 249192
rect 13789 248404 13801 249180
rect 13835 248404 13851 249180
rect 13789 248392 13851 248404
rect 13881 249180 13943 249192
rect 13881 248404 13897 249180
rect 13931 248404 13943 249180
rect 13881 248392 13943 248404
rect 13999 249180 14061 249192
rect 13999 248404 14011 249180
rect 14045 248404 14061 249180
rect 13999 248392 14061 248404
rect 14091 249180 14153 249192
rect 14091 248404 14107 249180
rect 14141 248404 14153 249180
rect 14091 248392 14153 248404
rect 14209 249180 14271 249192
rect 14209 248404 14221 249180
rect 14255 248404 14271 249180
rect 14209 248392 14271 248404
rect 14301 249180 14363 249192
rect 14301 248404 14317 249180
rect 14351 248404 14363 249180
rect 14301 248392 14363 248404
rect 14419 249180 14481 249192
rect 14419 248404 14431 249180
rect 14465 248404 14481 249180
rect 14419 248392 14481 248404
rect 14511 249180 14573 249192
rect 14511 248404 14527 249180
rect 14561 248404 14573 249180
rect 14511 248392 14573 248404
rect 14629 249180 14691 249192
rect 14629 248404 14641 249180
rect 14675 248404 14691 249180
rect 14629 248392 14691 248404
rect 14721 249180 14783 249192
rect 14721 248404 14737 249180
rect 14771 248404 14783 249180
rect 14721 248392 14783 248404
rect 14839 249180 14901 249192
rect 14839 248404 14851 249180
rect 14885 248404 14901 249180
rect 14839 248392 14901 248404
rect 14931 249180 14993 249192
rect 14931 248404 14947 249180
rect 14981 248404 14993 249180
rect 14931 248392 14993 248404
rect 15049 249180 15111 249192
rect 15049 248404 15061 249180
rect 15095 248404 15111 249180
rect 15049 248392 15111 248404
rect 15141 249180 15203 249192
rect 15141 248404 15157 249180
rect 15191 248404 15203 249180
rect 15141 248392 15203 248404
rect 15259 249180 15321 249192
rect 15259 248404 15271 249180
rect 15305 248404 15321 249180
rect 15259 248392 15321 248404
rect 15351 249180 15413 249192
rect 15351 248404 15367 249180
rect 15401 248404 15413 249180
rect 15351 248392 15413 248404
rect 15469 249180 15531 249192
rect 15469 248404 15481 249180
rect 15515 248404 15531 249180
rect 15469 248392 15531 248404
rect 15561 249180 15623 249192
rect 15561 248404 15577 249180
rect 15611 248404 15623 249180
rect 15561 248392 15623 248404
rect 15679 249180 15741 249192
rect 15679 248404 15691 249180
rect 15725 248404 15741 249180
rect 15679 248392 15741 248404
rect 15771 249180 15833 249192
rect 15771 248404 15787 249180
rect 15821 248404 15833 249180
rect 15771 248392 15833 248404
rect 15889 249180 15951 249192
rect 15889 248404 15901 249180
rect 15935 248404 15951 249180
rect 15889 248392 15951 248404
rect 15981 249180 16043 249192
rect 15981 248404 15997 249180
rect 16031 248404 16043 249180
rect 15981 248392 16043 248404
rect 16099 249180 16161 249192
rect 16099 248404 16111 249180
rect 16145 248404 16161 249180
rect 16099 248392 16161 248404
rect 16191 249180 16253 249192
rect 16191 248404 16207 249180
rect 16241 248404 16253 249180
rect 16191 248392 16253 248404
rect 16309 249180 16371 249192
rect 16309 248404 16321 249180
rect 16355 248404 16371 249180
rect 16309 248392 16371 248404
rect 16401 249180 16463 249192
rect 16401 248404 16417 249180
rect 16451 248404 16463 249180
rect 16401 248392 16463 248404
rect 16519 249180 16581 249192
rect 16519 248404 16531 249180
rect 16565 248404 16581 249180
rect 16519 248392 16581 248404
rect 16611 249180 16673 249192
rect 16611 248404 16627 249180
rect 16661 248404 16673 249180
rect 16611 248392 16673 248404
rect 16729 249180 16791 249192
rect 16729 248404 16741 249180
rect 16775 248404 16791 249180
rect 16729 248392 16791 248404
rect 16821 249180 16883 249192
rect 16821 248404 16837 249180
rect 16871 248404 16883 249180
rect 16821 248392 16883 248404
rect 16939 249180 17001 249192
rect 16939 248404 16951 249180
rect 16985 248404 17001 249180
rect 16939 248392 17001 248404
rect 17031 249180 17093 249192
rect 17031 248404 17047 249180
rect 17081 248404 17093 249180
rect 17031 248392 17093 248404
rect 17149 249180 17211 249192
rect 17149 248404 17161 249180
rect 17195 248404 17211 249180
rect 17149 248392 17211 248404
rect 17241 249180 17303 249192
rect 17241 248404 17257 249180
rect 17291 248404 17303 249180
rect 17241 248392 17303 248404
rect 17359 249180 17421 249192
rect 17359 248404 17371 249180
rect 17405 248404 17421 249180
rect 17359 248392 17421 248404
rect 17451 249180 17513 249192
rect 17451 248404 17467 249180
rect 17501 248404 17513 249180
rect 17451 248392 17513 248404
rect 17569 249180 17631 249192
rect 17569 248404 17581 249180
rect 17615 248404 17631 249180
rect 17569 248392 17631 248404
rect 17661 249180 17723 249192
rect 17661 248404 17677 249180
rect 17711 248404 17723 249180
rect 17661 248392 17723 248404
rect 17779 249180 17841 249192
rect 17779 248404 17791 249180
rect 17825 248404 17841 249180
rect 17779 248392 17841 248404
rect 17871 249180 17933 249192
rect 17871 248404 17887 249180
rect 17921 248404 17933 249180
rect 17871 248392 17933 248404
rect 17989 249180 18051 249192
rect 17989 248404 18001 249180
rect 18035 248404 18051 249180
rect 17989 248392 18051 248404
rect 18081 249180 18143 249192
rect 18081 248404 18097 249180
rect 18131 248404 18143 249180
rect 18081 248392 18143 248404
rect 18199 249180 18261 249192
rect 18199 248404 18211 249180
rect 18245 248404 18261 249180
rect 18199 248392 18261 248404
rect 18291 249180 18353 249192
rect 18291 248404 18307 249180
rect 18341 248404 18353 249180
rect 18291 248392 18353 248404
rect 18409 249180 18471 249192
rect 18409 248404 18421 249180
rect 18455 248404 18471 249180
rect 18409 248392 18471 248404
rect 18501 249180 18563 249192
rect 18501 248404 18517 249180
rect 18551 248404 18563 249180
rect 18501 248392 18563 248404
rect 18619 249180 18681 249192
rect 18619 248404 18631 249180
rect 18665 248404 18681 249180
rect 18619 248392 18681 248404
rect 18711 249180 18773 249192
rect 18711 248404 18727 249180
rect 18761 248404 18773 249180
rect 18711 248392 18773 248404
rect 18829 249180 18891 249192
rect 18829 248404 18841 249180
rect 18875 248404 18891 249180
rect 18829 248392 18891 248404
rect 18921 249180 18983 249192
rect 18921 248404 18937 249180
rect 18971 248404 18983 249180
rect 18921 248392 18983 248404
rect 19039 249180 19101 249192
rect 19039 248404 19051 249180
rect 19085 248404 19101 249180
rect 19039 248392 19101 248404
rect 19131 249180 19193 249192
rect 19131 248404 19147 249180
rect 19181 248404 19193 249180
rect 19131 248392 19193 248404
rect 19249 249180 19311 249192
rect 19249 248404 19261 249180
rect 19295 248404 19311 249180
rect 19249 248392 19311 248404
rect 19341 249180 19403 249192
rect 19341 248404 19357 249180
rect 19391 248404 19403 249180
rect 19341 248392 19403 248404
rect 19459 249180 19521 249192
rect 19459 248404 19471 249180
rect 19505 248404 19521 249180
rect 19459 248392 19521 248404
rect 19551 249180 19613 249192
rect 19551 248404 19567 249180
rect 19601 248404 19613 249180
rect 19551 248392 19613 248404
rect 19669 249180 19731 249192
rect 19669 248404 19681 249180
rect 19715 248404 19731 249180
rect 19669 248392 19731 248404
rect 19761 249180 19823 249192
rect 19761 248404 19777 249180
rect 19811 248404 19823 249180
rect 19761 248392 19823 248404
rect 19879 249180 19941 249192
rect 19879 248404 19891 249180
rect 19925 248404 19941 249180
rect 19879 248392 19941 248404
rect 19971 249180 20033 249192
rect 19971 248404 19987 249180
rect 20021 248404 20033 249180
rect 19971 248392 20033 248404
rect 20089 249180 20151 249192
rect 20089 248404 20101 249180
rect 20135 248404 20151 249180
rect 20089 248392 20151 248404
rect 20181 249180 20243 249192
rect 20181 248404 20197 249180
rect 20231 248404 20243 249180
rect 20181 248392 20243 248404
rect 20299 249180 20361 249192
rect 20299 248404 20311 249180
rect 20345 248404 20361 249180
rect 20299 248392 20361 248404
rect 20391 249180 20453 249192
rect 20391 248404 20407 249180
rect 20441 248404 20453 249180
rect 20391 248392 20453 248404
rect 20509 249180 20571 249192
rect 20509 248404 20521 249180
rect 20555 248404 20571 249180
rect 20509 248392 20571 248404
rect 20601 249180 20663 249192
rect 20601 248404 20617 249180
rect 20651 248404 20663 249180
rect 20601 248392 20663 248404
rect 20719 249180 20781 249192
rect 20719 248404 20731 249180
rect 20765 248404 20781 249180
rect 20719 248392 20781 248404
rect 20811 249180 20873 249192
rect 20811 248404 20827 249180
rect 20861 248404 20873 249180
rect 20811 248392 20873 248404
rect 20929 249180 20991 249192
rect 20929 248404 20941 249180
rect 20975 248404 20991 249180
rect 20929 248392 20991 248404
rect 21021 249180 21083 249192
rect 21021 248404 21037 249180
rect 21071 248404 21083 249180
rect 21021 248392 21083 248404
rect 21139 249180 21201 249192
rect 21139 248404 21151 249180
rect 21185 248404 21201 249180
rect 21139 248392 21201 248404
rect 21231 249180 21293 249192
rect 21231 248404 21247 249180
rect 21281 248404 21293 249180
rect 21231 248392 21293 248404
rect 21349 249180 21411 249192
rect 21349 248404 21361 249180
rect 21395 248404 21411 249180
rect 21349 248392 21411 248404
rect 21441 249180 21503 249192
rect 21441 248404 21457 249180
rect 21491 248404 21503 249180
rect 21441 248392 21503 248404
rect 21559 249180 21621 249192
rect 21559 248404 21571 249180
rect 21605 248404 21621 249180
rect 21559 248392 21621 248404
rect 21651 249180 21713 249192
rect 21651 248404 21667 249180
rect 21701 248404 21713 249180
rect 21651 248392 21713 248404
rect 21769 249180 21831 249192
rect 21769 248404 21781 249180
rect 21815 248404 21831 249180
rect 21769 248392 21831 248404
rect 21861 249180 21923 249192
rect 21861 248404 21877 249180
rect 21911 248404 21923 249180
rect 21861 248392 21923 248404
rect 21979 249180 22041 249192
rect 21979 248404 21991 249180
rect 22025 248404 22041 249180
rect 21979 248392 22041 248404
rect 22071 249180 22133 249192
rect 22071 248404 22087 249180
rect 22121 248404 22133 249180
rect 22071 248392 22133 248404
rect 22189 249180 22251 249192
rect 22189 248404 22201 249180
rect 22235 248404 22251 249180
rect 22189 248392 22251 248404
rect 22281 249180 22343 249192
rect 22281 248404 22297 249180
rect 22331 248404 22343 249180
rect 22281 248392 22343 248404
rect 22399 249180 22461 249192
rect 22399 248404 22411 249180
rect 22445 248404 22461 249180
rect 22399 248392 22461 248404
rect 22491 249180 22553 249192
rect 22491 248404 22507 249180
rect 22541 248404 22553 249180
rect 22491 248392 22553 248404
rect 22609 249180 22671 249192
rect 22609 248404 22621 249180
rect 22655 248404 22671 249180
rect 22609 248392 22671 248404
rect 22701 249180 22763 249192
rect 22701 248404 22717 249180
rect 22751 248404 22763 249180
rect 22701 248392 22763 248404
rect 22819 249180 22881 249192
rect 22819 248404 22831 249180
rect 22865 248404 22881 249180
rect 22819 248392 22881 248404
rect 22911 249180 22973 249192
rect 22911 248404 22927 249180
rect 22961 248404 22973 249180
rect 22911 248392 22973 248404
rect 23029 249180 23091 249192
rect 23029 248404 23041 249180
rect 23075 248404 23091 249180
rect 23029 248392 23091 248404
rect 23121 249180 23183 249192
rect 23121 248404 23137 249180
rect 23171 248404 23183 249180
rect 23121 248392 23183 248404
rect 23239 249180 23301 249192
rect 23239 248404 23251 249180
rect 23285 248404 23301 249180
rect 23239 248392 23301 248404
rect 23331 249180 23393 249192
rect 23331 248404 23347 249180
rect 23381 248404 23393 249180
rect 23331 248392 23393 248404
rect 23449 249180 23511 249192
rect 23449 248404 23461 249180
rect 23495 248404 23511 249180
rect 23449 248392 23511 248404
rect 23541 249180 23603 249192
rect 23541 248404 23557 249180
rect 23591 248404 23603 249180
rect 23541 248392 23603 248404
rect 23659 249180 23721 249192
rect 23659 248404 23671 249180
rect 23705 248404 23721 249180
rect 23659 248392 23721 248404
rect 23751 249180 23813 249192
rect 23751 248404 23767 249180
rect 23801 248404 23813 249180
rect 23751 248392 23813 248404
rect 23869 249180 23931 249192
rect 23869 248404 23881 249180
rect 23915 248404 23931 249180
rect 23869 248392 23931 248404
rect 23961 249180 24023 249192
rect 23961 248404 23977 249180
rect 24011 248404 24023 249180
rect 23961 248392 24023 248404
rect 24079 249180 24141 249192
rect 24079 248404 24091 249180
rect 24125 248404 24141 249180
rect 24079 248392 24141 248404
rect 24171 249180 24233 249192
rect 24171 248404 24187 249180
rect 24221 248404 24233 249180
rect 24171 248392 24233 248404
rect 24289 249180 24351 249192
rect 24289 248404 24301 249180
rect 24335 248404 24351 249180
rect 24289 248392 24351 248404
rect 24381 249180 24443 249192
rect 24381 248404 24397 249180
rect 24431 248404 24443 249180
rect 24381 248392 24443 248404
rect 24499 249180 24561 249192
rect 24499 248404 24511 249180
rect 24545 248404 24561 249180
rect 24499 248392 24561 248404
rect 24591 249180 24653 249192
rect 24591 248404 24607 249180
rect 24641 248404 24653 249180
rect 24591 248392 24653 248404
rect 24709 249180 24771 249192
rect 24709 248404 24721 249180
rect 24755 248404 24771 249180
rect 24709 248392 24771 248404
rect 24801 249180 24863 249192
rect 24801 248404 24817 249180
rect 24851 248404 24863 249180
rect 24801 248392 24863 248404
rect 24919 249180 24981 249192
rect 24919 248404 24931 249180
rect 24965 248404 24981 249180
rect 24919 248392 24981 248404
rect 25011 249180 25073 249192
rect 25011 248404 25027 249180
rect 25061 248404 25073 249180
rect 25011 248392 25073 248404
rect 25129 249180 25191 249192
rect 25129 248404 25141 249180
rect 25175 248404 25191 249180
rect 25129 248392 25191 248404
rect 25221 249180 25283 249192
rect 25221 248404 25237 249180
rect 25271 248404 25283 249180
rect 25221 248392 25283 248404
rect 25339 249180 25401 249192
rect 25339 248404 25351 249180
rect 25385 248404 25401 249180
rect 25339 248392 25401 248404
rect 25431 249180 25493 249192
rect 25431 248404 25447 249180
rect 25481 248404 25493 249180
rect 25431 248392 25493 248404
rect 25549 249180 25611 249192
rect 25549 248404 25561 249180
rect 25595 248404 25611 249180
rect 25549 248392 25611 248404
rect 25641 249180 25703 249192
rect 25641 248404 25657 249180
rect 25691 248404 25703 249180
rect 25641 248392 25703 248404
rect 25759 249180 25821 249192
rect 25759 248404 25771 249180
rect 25805 248404 25821 249180
rect 25759 248392 25821 248404
rect 25851 249180 25913 249192
rect 25851 248404 25867 249180
rect 25901 248404 25913 249180
rect 25851 248392 25913 248404
rect 25969 249180 26031 249192
rect 25969 248404 25981 249180
rect 26015 248404 26031 249180
rect 25969 248392 26031 248404
rect 26061 249180 26123 249192
rect 26061 248404 26077 249180
rect 26111 248404 26123 249180
rect 26061 248392 26123 248404
rect 26179 249180 26241 249192
rect 26179 248404 26191 249180
rect 26225 248404 26241 249180
rect 26179 248392 26241 248404
rect 26271 249180 26333 249192
rect 26271 248404 26287 249180
rect 26321 248404 26333 249180
rect 26271 248392 26333 248404
rect 26389 249180 26451 249192
rect 26389 248404 26401 249180
rect 26435 248404 26451 249180
rect 26389 248392 26451 248404
rect 26481 249180 26543 249192
rect 26481 248404 26497 249180
rect 26531 248404 26543 249180
rect 26481 248392 26543 248404
rect 26599 249180 26661 249192
rect 26599 248404 26611 249180
rect 26645 248404 26661 249180
rect 26599 248392 26661 248404
rect 26691 249180 26753 249192
rect 26691 248404 26707 249180
rect 26741 248404 26753 249180
rect 26691 248392 26753 248404
rect 26809 249180 26871 249192
rect 26809 248404 26821 249180
rect 26855 248404 26871 249180
rect 26809 248392 26871 248404
rect 26901 249180 26963 249192
rect 26901 248404 26917 249180
rect 26951 248404 26963 249180
rect 26901 248392 26963 248404
rect 27019 249180 27081 249192
rect 27019 248404 27031 249180
rect 27065 248404 27081 249180
rect 27019 248392 27081 248404
rect 27111 249180 27173 249192
rect 27111 248404 27127 249180
rect 27161 248404 27173 249180
rect 27111 248392 27173 248404
rect 27229 249180 27291 249192
rect 27229 248404 27241 249180
rect 27275 248404 27291 249180
rect 27229 248392 27291 248404
rect 27321 249180 27383 249192
rect 27321 248404 27337 249180
rect 27371 248404 27383 249180
rect 27321 248392 27383 248404
rect -4061 248144 -3999 248156
rect -4061 247368 -4049 248144
rect -4015 247368 -3999 248144
rect -4061 247356 -3999 247368
rect -3969 248144 -3907 248156
rect -3969 247368 -3953 248144
rect -3919 247368 -3907 248144
rect -3969 247356 -3907 247368
rect -3851 248144 -3789 248156
rect -3851 247368 -3839 248144
rect -3805 247368 -3789 248144
rect -3851 247356 -3789 247368
rect -3759 248144 -3697 248156
rect -3759 247368 -3743 248144
rect -3709 247368 -3697 248144
rect -3759 247356 -3697 247368
rect -3641 248144 -3579 248156
rect -3641 247368 -3629 248144
rect -3595 247368 -3579 248144
rect -3641 247356 -3579 247368
rect -3549 248144 -3487 248156
rect -3549 247368 -3533 248144
rect -3499 247368 -3487 248144
rect -3549 247356 -3487 247368
rect -3431 248144 -3369 248156
rect -3431 247368 -3419 248144
rect -3385 247368 -3369 248144
rect -3431 247356 -3369 247368
rect -3339 248144 -3277 248156
rect -3339 247368 -3323 248144
rect -3289 247368 -3277 248144
rect -3339 247356 -3277 247368
rect -3221 248144 -3159 248156
rect -3221 247368 -3209 248144
rect -3175 247368 -3159 248144
rect -3221 247356 -3159 247368
rect -3129 248144 -3067 248156
rect -3129 247368 -3113 248144
rect -3079 247368 -3067 248144
rect -3129 247356 -3067 247368
rect -3011 248144 -2949 248156
rect -3011 247368 -2999 248144
rect -2965 247368 -2949 248144
rect -3011 247356 -2949 247368
rect -2919 248144 -2857 248156
rect -2919 247368 -2903 248144
rect -2869 247368 -2857 248144
rect -2919 247356 -2857 247368
rect -2801 248144 -2739 248156
rect -2801 247368 -2789 248144
rect -2755 247368 -2739 248144
rect -2801 247356 -2739 247368
rect -2709 248144 -2647 248156
rect -2709 247368 -2693 248144
rect -2659 247368 -2647 248144
rect -2709 247356 -2647 247368
rect -2591 248144 -2529 248156
rect -2591 247368 -2579 248144
rect -2545 247368 -2529 248144
rect -2591 247356 -2529 247368
rect -2499 248144 -2437 248156
rect -2499 247368 -2483 248144
rect -2449 247368 -2437 248144
rect -2499 247356 -2437 247368
rect -2381 248144 -2319 248156
rect -2381 247368 -2369 248144
rect -2335 247368 -2319 248144
rect -2381 247356 -2319 247368
rect -2289 248144 -2227 248156
rect -2289 247368 -2273 248144
rect -2239 247368 -2227 248144
rect -2289 247356 -2227 247368
rect -2171 248144 -2109 248156
rect -2171 247368 -2159 248144
rect -2125 247368 -2109 248144
rect -2171 247356 -2109 247368
rect -2079 248144 -2017 248156
rect -2079 247368 -2063 248144
rect -2029 247368 -2017 248144
rect -2079 247356 -2017 247368
rect -1961 248144 -1899 248156
rect -1961 247368 -1949 248144
rect -1915 247368 -1899 248144
rect -1961 247356 -1899 247368
rect -1869 248144 -1807 248156
rect -1869 247368 -1853 248144
rect -1819 247368 -1807 248144
rect -1869 247356 -1807 247368
rect -1751 248144 -1689 248156
rect -1751 247368 -1739 248144
rect -1705 247368 -1689 248144
rect -1751 247356 -1689 247368
rect -1659 248144 -1597 248156
rect -1659 247368 -1643 248144
rect -1609 247368 -1597 248144
rect -1659 247356 -1597 247368
rect -1541 248144 -1479 248156
rect -1541 247368 -1529 248144
rect -1495 247368 -1479 248144
rect -1541 247356 -1479 247368
rect -1449 248144 -1387 248156
rect -1449 247368 -1433 248144
rect -1399 247368 -1387 248144
rect -1449 247356 -1387 247368
rect -1331 248144 -1269 248156
rect -1331 247368 -1319 248144
rect -1285 247368 -1269 248144
rect -1331 247356 -1269 247368
rect -1239 248144 -1177 248156
rect -1239 247368 -1223 248144
rect -1189 247368 -1177 248144
rect -1239 247356 -1177 247368
rect -1121 248144 -1059 248156
rect -1121 247368 -1109 248144
rect -1075 247368 -1059 248144
rect -1121 247356 -1059 247368
rect -1029 248144 -967 248156
rect -1029 247368 -1013 248144
rect -979 247368 -967 248144
rect -1029 247356 -967 247368
rect -911 248144 -849 248156
rect -911 247368 -899 248144
rect -865 247368 -849 248144
rect -911 247356 -849 247368
rect -819 248144 -757 248156
rect -819 247368 -803 248144
rect -769 247368 -757 248144
rect -819 247356 -757 247368
rect -701 248144 -639 248156
rect -701 247368 -689 248144
rect -655 247368 -639 248144
rect -701 247356 -639 247368
rect -609 248144 -547 248156
rect -609 247368 -593 248144
rect -559 247368 -547 248144
rect -609 247356 -547 247368
rect -491 248144 -429 248156
rect -491 247368 -479 248144
rect -445 247368 -429 248144
rect -491 247356 -429 247368
rect -399 248144 -337 248156
rect -399 247368 -383 248144
rect -349 247368 -337 248144
rect -399 247356 -337 247368
rect -281 248144 -219 248156
rect -281 247368 -269 248144
rect -235 247368 -219 248144
rect -281 247356 -219 247368
rect -189 248144 -127 248156
rect -189 247368 -173 248144
rect -139 247368 -127 248144
rect -189 247356 -127 247368
rect -71 248144 -9 248156
rect -71 247368 -59 248144
rect -25 247368 -9 248144
rect -71 247356 -9 247368
rect 21 248144 83 248156
rect 21 247368 37 248144
rect 71 247368 83 248144
rect 21 247356 83 247368
rect 139 248144 201 248156
rect 139 247368 151 248144
rect 185 247368 201 248144
rect 139 247356 201 247368
rect 231 248144 293 248156
rect 231 247368 247 248144
rect 281 247368 293 248144
rect 231 247356 293 247368
rect 349 248144 411 248156
rect 349 247368 361 248144
rect 395 247368 411 248144
rect 349 247356 411 247368
rect 441 248144 503 248156
rect 441 247368 457 248144
rect 491 247368 503 248144
rect 441 247356 503 247368
rect 559 248144 621 248156
rect 559 247368 571 248144
rect 605 247368 621 248144
rect 559 247356 621 247368
rect 651 248144 713 248156
rect 651 247368 667 248144
rect 701 247368 713 248144
rect 651 247356 713 247368
rect 769 248144 831 248156
rect 769 247368 781 248144
rect 815 247368 831 248144
rect 769 247356 831 247368
rect 861 248144 923 248156
rect 861 247368 877 248144
rect 911 247368 923 248144
rect 861 247356 923 247368
rect 979 248144 1041 248156
rect 979 247368 991 248144
rect 1025 247368 1041 248144
rect 979 247356 1041 247368
rect 1071 248144 1133 248156
rect 1071 247368 1087 248144
rect 1121 247368 1133 248144
rect 1071 247356 1133 247368
rect 1189 248144 1251 248156
rect 1189 247368 1201 248144
rect 1235 247368 1251 248144
rect 1189 247356 1251 247368
rect 1281 248144 1343 248156
rect 1281 247368 1297 248144
rect 1331 247368 1343 248144
rect 1281 247356 1343 247368
rect 1399 248144 1461 248156
rect 1399 247368 1411 248144
rect 1445 247368 1461 248144
rect 1399 247356 1461 247368
rect 1491 248144 1553 248156
rect 1491 247368 1507 248144
rect 1541 247368 1553 248144
rect 1491 247356 1553 247368
rect 1609 248144 1671 248156
rect 1609 247368 1621 248144
rect 1655 247368 1671 248144
rect 1609 247356 1671 247368
rect 1701 248144 1763 248156
rect 1701 247368 1717 248144
rect 1751 247368 1763 248144
rect 1701 247356 1763 247368
rect 1819 248144 1881 248156
rect 1819 247368 1831 248144
rect 1865 247368 1881 248144
rect 1819 247356 1881 247368
rect 1911 248144 1973 248156
rect 1911 247368 1927 248144
rect 1961 247368 1973 248144
rect 1911 247356 1973 247368
rect 2029 248144 2091 248156
rect 2029 247368 2041 248144
rect 2075 247368 2091 248144
rect 2029 247356 2091 247368
rect 2121 248144 2183 248156
rect 2121 247368 2137 248144
rect 2171 247368 2183 248144
rect 2121 247356 2183 247368
rect 2239 248144 2301 248156
rect 2239 247368 2251 248144
rect 2285 247368 2301 248144
rect 2239 247356 2301 247368
rect 2331 248144 2393 248156
rect 2331 247368 2347 248144
rect 2381 247368 2393 248144
rect 2331 247356 2393 247368
rect 2449 248144 2511 248156
rect 2449 247368 2461 248144
rect 2495 247368 2511 248144
rect 2449 247356 2511 247368
rect 2541 248144 2603 248156
rect 2541 247368 2557 248144
rect 2591 247368 2603 248144
rect 2541 247356 2603 247368
rect 2659 248144 2721 248156
rect 2659 247368 2671 248144
rect 2705 247368 2721 248144
rect 2659 247356 2721 247368
rect 2751 248144 2813 248156
rect 2751 247368 2767 248144
rect 2801 247368 2813 248144
rect 2751 247356 2813 247368
rect 2869 248144 2931 248156
rect 2869 247368 2881 248144
rect 2915 247368 2931 248144
rect 2869 247356 2931 247368
rect 2961 248144 3023 248156
rect 2961 247368 2977 248144
rect 3011 247368 3023 248144
rect 2961 247356 3023 247368
rect 3079 248144 3141 248156
rect 3079 247368 3091 248144
rect 3125 247368 3141 248144
rect 3079 247356 3141 247368
rect 3171 248144 3233 248156
rect 3171 247368 3187 248144
rect 3221 247368 3233 248144
rect 3171 247356 3233 247368
rect 3289 248144 3351 248156
rect 3289 247368 3301 248144
rect 3335 247368 3351 248144
rect 3289 247356 3351 247368
rect 3381 248144 3443 248156
rect 3381 247368 3397 248144
rect 3431 247368 3443 248144
rect 3381 247356 3443 247368
rect 3499 248144 3561 248156
rect 3499 247368 3511 248144
rect 3545 247368 3561 248144
rect 3499 247356 3561 247368
rect 3591 248144 3653 248156
rect 3591 247368 3607 248144
rect 3641 247368 3653 248144
rect 3591 247356 3653 247368
rect 3709 248144 3771 248156
rect 3709 247368 3721 248144
rect 3755 247368 3771 248144
rect 3709 247356 3771 247368
rect 3801 248144 3863 248156
rect 3801 247368 3817 248144
rect 3851 247368 3863 248144
rect 3801 247356 3863 247368
rect 3919 248144 3981 248156
rect 3919 247368 3931 248144
rect 3965 247368 3981 248144
rect 3919 247356 3981 247368
rect 4011 248144 4073 248156
rect 4011 247368 4027 248144
rect 4061 247368 4073 248144
rect 4011 247356 4073 247368
rect 4129 248144 4191 248156
rect 4129 247368 4141 248144
rect 4175 247368 4191 248144
rect 4129 247356 4191 247368
rect 4221 248144 4283 248156
rect 4221 247368 4237 248144
rect 4271 247368 4283 248144
rect 4221 247356 4283 247368
rect 4339 248144 4401 248156
rect 4339 247368 4351 248144
rect 4385 247368 4401 248144
rect 4339 247356 4401 247368
rect 4431 248144 4493 248156
rect 4431 247368 4447 248144
rect 4481 247368 4493 248144
rect 4431 247356 4493 247368
rect 4549 248144 4611 248156
rect 4549 247368 4561 248144
rect 4595 247368 4611 248144
rect 4549 247356 4611 247368
rect 4641 248144 4703 248156
rect 4641 247368 4657 248144
rect 4691 247368 4703 248144
rect 4641 247356 4703 247368
rect 4759 248144 4821 248156
rect 4759 247368 4771 248144
rect 4805 247368 4821 248144
rect 4759 247356 4821 247368
rect 4851 248144 4913 248156
rect 4851 247368 4867 248144
rect 4901 247368 4913 248144
rect 4851 247356 4913 247368
rect 4969 248144 5031 248156
rect 4969 247368 4981 248144
rect 5015 247368 5031 248144
rect 4969 247356 5031 247368
rect 5061 248144 5123 248156
rect 5061 247368 5077 248144
rect 5111 247368 5123 248144
rect 5061 247356 5123 247368
rect 5179 248144 5241 248156
rect 5179 247368 5191 248144
rect 5225 247368 5241 248144
rect 5179 247356 5241 247368
rect 5271 248144 5333 248156
rect 5271 247368 5287 248144
rect 5321 247368 5333 248144
rect 5271 247356 5333 247368
rect 5389 248144 5451 248156
rect 5389 247368 5401 248144
rect 5435 247368 5451 248144
rect 5389 247356 5451 247368
rect 5481 248144 5543 248156
rect 5481 247368 5497 248144
rect 5531 247368 5543 248144
rect 5481 247356 5543 247368
rect 5599 248144 5661 248156
rect 5599 247368 5611 248144
rect 5645 247368 5661 248144
rect 5599 247356 5661 247368
rect 5691 248144 5753 248156
rect 5691 247368 5707 248144
rect 5741 247368 5753 248144
rect 5691 247356 5753 247368
rect 5809 248144 5871 248156
rect 5809 247368 5821 248144
rect 5855 247368 5871 248144
rect 5809 247356 5871 247368
rect 5901 248144 5963 248156
rect 5901 247368 5917 248144
rect 5951 247368 5963 248144
rect 5901 247356 5963 247368
rect 6019 248144 6081 248156
rect 6019 247368 6031 248144
rect 6065 247368 6081 248144
rect 6019 247356 6081 247368
rect 6111 248144 6173 248156
rect 6111 247368 6127 248144
rect 6161 247368 6173 248144
rect 6111 247356 6173 247368
rect 6229 248144 6291 248156
rect 6229 247368 6241 248144
rect 6275 247368 6291 248144
rect 6229 247356 6291 247368
rect 6321 248144 6383 248156
rect 6321 247368 6337 248144
rect 6371 247368 6383 248144
rect 6321 247356 6383 247368
rect 6439 248144 6501 248156
rect 6439 247368 6451 248144
rect 6485 247368 6501 248144
rect 6439 247356 6501 247368
rect 6531 248144 6593 248156
rect 6531 247368 6547 248144
rect 6581 247368 6593 248144
rect 6531 247356 6593 247368
rect 6649 248144 6711 248156
rect 6649 247368 6661 248144
rect 6695 247368 6711 248144
rect 6649 247356 6711 247368
rect 6741 248144 6803 248156
rect 6741 247368 6757 248144
rect 6791 247368 6803 248144
rect 6741 247356 6803 247368
rect 6859 248144 6921 248156
rect 6859 247368 6871 248144
rect 6905 247368 6921 248144
rect 6859 247356 6921 247368
rect 6951 248144 7013 248156
rect 6951 247368 6967 248144
rect 7001 247368 7013 248144
rect 6951 247356 7013 247368
rect 7069 248144 7131 248156
rect 7069 247368 7081 248144
rect 7115 247368 7131 248144
rect 7069 247356 7131 247368
rect 7161 248144 7223 248156
rect 7161 247368 7177 248144
rect 7211 247368 7223 248144
rect 7161 247356 7223 247368
rect 7279 248144 7341 248156
rect 7279 247368 7291 248144
rect 7325 247368 7341 248144
rect 7279 247356 7341 247368
rect 7371 248144 7433 248156
rect 7371 247368 7387 248144
rect 7421 247368 7433 248144
rect 7371 247356 7433 247368
rect 7489 248144 7551 248156
rect 7489 247368 7501 248144
rect 7535 247368 7551 248144
rect 7489 247356 7551 247368
rect 7581 248144 7643 248156
rect 7581 247368 7597 248144
rect 7631 247368 7643 248144
rect 7581 247356 7643 247368
rect 7699 248144 7761 248156
rect 7699 247368 7711 248144
rect 7745 247368 7761 248144
rect 7699 247356 7761 247368
rect 7791 248144 7853 248156
rect 7791 247368 7807 248144
rect 7841 247368 7853 248144
rect 7791 247356 7853 247368
rect 7909 248144 7971 248156
rect 7909 247368 7921 248144
rect 7955 247368 7971 248144
rect 7909 247356 7971 247368
rect 8001 248144 8063 248156
rect 8001 247368 8017 248144
rect 8051 247368 8063 248144
rect 8001 247356 8063 247368
rect 8119 248144 8181 248156
rect 8119 247368 8131 248144
rect 8165 247368 8181 248144
rect 8119 247356 8181 247368
rect 8211 248144 8273 248156
rect 8211 247368 8227 248144
rect 8261 247368 8273 248144
rect 8211 247356 8273 247368
rect 8329 248144 8391 248156
rect 8329 247368 8341 248144
rect 8375 247368 8391 248144
rect 8329 247356 8391 247368
rect 8421 248144 8483 248156
rect 8421 247368 8437 248144
rect 8471 247368 8483 248144
rect 8421 247356 8483 247368
rect 8539 248144 8601 248156
rect 8539 247368 8551 248144
rect 8585 247368 8601 248144
rect 8539 247356 8601 247368
rect 8631 248144 8693 248156
rect 8631 247368 8647 248144
rect 8681 247368 8693 248144
rect 8631 247356 8693 247368
rect 8749 248144 8811 248156
rect 8749 247368 8761 248144
rect 8795 247368 8811 248144
rect 8749 247356 8811 247368
rect 8841 248144 8903 248156
rect 8841 247368 8857 248144
rect 8891 247368 8903 248144
rect 8841 247356 8903 247368
rect 8959 248144 9021 248156
rect 8959 247368 8971 248144
rect 9005 247368 9021 248144
rect 8959 247356 9021 247368
rect 9051 248144 9113 248156
rect 9051 247368 9067 248144
rect 9101 247368 9113 248144
rect 9051 247356 9113 247368
rect 9169 248144 9231 248156
rect 9169 247368 9181 248144
rect 9215 247368 9231 248144
rect 9169 247356 9231 247368
rect 9261 248144 9323 248156
rect 9261 247368 9277 248144
rect 9311 247368 9323 248144
rect 9261 247356 9323 247368
rect 9379 248144 9441 248156
rect 9379 247368 9391 248144
rect 9425 247368 9441 248144
rect 9379 247356 9441 247368
rect 9471 248144 9533 248156
rect 9471 247368 9487 248144
rect 9521 247368 9533 248144
rect 9471 247356 9533 247368
rect 9589 248144 9651 248156
rect 9589 247368 9601 248144
rect 9635 247368 9651 248144
rect 9589 247356 9651 247368
rect 9681 248144 9743 248156
rect 9681 247368 9697 248144
rect 9731 247368 9743 248144
rect 9681 247356 9743 247368
rect 9799 248144 9861 248156
rect 9799 247368 9811 248144
rect 9845 247368 9861 248144
rect 9799 247356 9861 247368
rect 9891 248144 9953 248156
rect 9891 247368 9907 248144
rect 9941 247368 9953 248144
rect 9891 247356 9953 247368
rect 10009 248144 10071 248156
rect 10009 247368 10021 248144
rect 10055 247368 10071 248144
rect 10009 247356 10071 247368
rect 10101 248144 10163 248156
rect 10101 247368 10117 248144
rect 10151 247368 10163 248144
rect 10101 247356 10163 247368
rect 10219 248144 10281 248156
rect 10219 247368 10231 248144
rect 10265 247368 10281 248144
rect 10219 247356 10281 247368
rect 10311 248144 10373 248156
rect 10311 247368 10327 248144
rect 10361 247368 10373 248144
rect 10311 247356 10373 247368
rect 10429 248144 10491 248156
rect 10429 247368 10441 248144
rect 10475 247368 10491 248144
rect 10429 247356 10491 247368
rect 10521 248144 10583 248156
rect 10521 247368 10537 248144
rect 10571 247368 10583 248144
rect 10521 247356 10583 247368
rect 10639 248144 10701 248156
rect 10639 247368 10651 248144
rect 10685 247368 10701 248144
rect 10639 247356 10701 247368
rect 10731 248144 10793 248156
rect 10731 247368 10747 248144
rect 10781 247368 10793 248144
rect 10731 247356 10793 247368
rect 10849 248144 10911 248156
rect 10849 247368 10861 248144
rect 10895 247368 10911 248144
rect 10849 247356 10911 247368
rect 10941 248144 11003 248156
rect 10941 247368 10957 248144
rect 10991 247368 11003 248144
rect 10941 247356 11003 247368
rect 11059 248144 11121 248156
rect 11059 247368 11071 248144
rect 11105 247368 11121 248144
rect 11059 247356 11121 247368
rect 11151 248144 11213 248156
rect 11151 247368 11167 248144
rect 11201 247368 11213 248144
rect 11151 247356 11213 247368
rect 11269 248144 11331 248156
rect 11269 247368 11281 248144
rect 11315 247368 11331 248144
rect 11269 247356 11331 247368
rect 11361 248144 11423 248156
rect 11361 247368 11377 248144
rect 11411 247368 11423 248144
rect 11361 247356 11423 247368
rect 11479 248144 11541 248156
rect 11479 247368 11491 248144
rect 11525 247368 11541 248144
rect 11479 247356 11541 247368
rect 11571 248144 11633 248156
rect 11571 247368 11587 248144
rect 11621 247368 11633 248144
rect 11571 247356 11633 247368
rect 11689 248144 11751 248156
rect 11689 247368 11701 248144
rect 11735 247368 11751 248144
rect 11689 247356 11751 247368
rect 11781 248144 11843 248156
rect 11781 247368 11797 248144
rect 11831 247368 11843 248144
rect 11781 247356 11843 247368
rect 11899 248144 11961 248156
rect 11899 247368 11911 248144
rect 11945 247368 11961 248144
rect 11899 247356 11961 247368
rect 11991 248144 12053 248156
rect 11991 247368 12007 248144
rect 12041 247368 12053 248144
rect 11991 247356 12053 247368
rect 12109 248144 12171 248156
rect 12109 247368 12121 248144
rect 12155 247368 12171 248144
rect 12109 247356 12171 247368
rect 12201 248144 12263 248156
rect 12201 247368 12217 248144
rect 12251 247368 12263 248144
rect 12201 247356 12263 247368
rect 12319 248144 12381 248156
rect 12319 247368 12331 248144
rect 12365 247368 12381 248144
rect 12319 247356 12381 247368
rect 12411 248144 12473 248156
rect 12411 247368 12427 248144
rect 12461 247368 12473 248144
rect 12411 247356 12473 247368
rect 12529 248144 12591 248156
rect 12529 247368 12541 248144
rect 12575 247368 12591 248144
rect 12529 247356 12591 247368
rect 12621 248144 12683 248156
rect 12621 247368 12637 248144
rect 12671 247368 12683 248144
rect 12621 247356 12683 247368
rect 12739 248144 12801 248156
rect 12739 247368 12751 248144
rect 12785 247368 12801 248144
rect 12739 247356 12801 247368
rect 12831 248144 12893 248156
rect 12831 247368 12847 248144
rect 12881 247368 12893 248144
rect 12831 247356 12893 247368
rect 12949 248144 13011 248156
rect 12949 247368 12961 248144
rect 12995 247368 13011 248144
rect 12949 247356 13011 247368
rect 13041 248144 13103 248156
rect 13041 247368 13057 248144
rect 13091 247368 13103 248144
rect 13041 247356 13103 247368
rect 13159 248144 13221 248156
rect 13159 247368 13171 248144
rect 13205 247368 13221 248144
rect 13159 247356 13221 247368
rect 13251 248144 13313 248156
rect 13251 247368 13267 248144
rect 13301 247368 13313 248144
rect 13251 247356 13313 247368
rect 13369 248144 13431 248156
rect 13369 247368 13381 248144
rect 13415 247368 13431 248144
rect 13369 247356 13431 247368
rect 13461 248144 13523 248156
rect 13461 247368 13477 248144
rect 13511 247368 13523 248144
rect 13461 247356 13523 247368
rect 13579 248144 13641 248156
rect 13579 247368 13591 248144
rect 13625 247368 13641 248144
rect 13579 247356 13641 247368
rect 13671 248144 13733 248156
rect 13671 247368 13687 248144
rect 13721 247368 13733 248144
rect 13671 247356 13733 247368
rect 13789 248144 13851 248156
rect 13789 247368 13801 248144
rect 13835 247368 13851 248144
rect 13789 247356 13851 247368
rect 13881 248144 13943 248156
rect 13881 247368 13897 248144
rect 13931 247368 13943 248144
rect 13881 247356 13943 247368
rect 13999 248144 14061 248156
rect 13999 247368 14011 248144
rect 14045 247368 14061 248144
rect 13999 247356 14061 247368
rect 14091 248144 14153 248156
rect 14091 247368 14107 248144
rect 14141 247368 14153 248144
rect 14091 247356 14153 247368
rect 14209 248144 14271 248156
rect 14209 247368 14221 248144
rect 14255 247368 14271 248144
rect 14209 247356 14271 247368
rect 14301 248144 14363 248156
rect 14301 247368 14317 248144
rect 14351 247368 14363 248144
rect 14301 247356 14363 247368
rect 14419 248144 14481 248156
rect 14419 247368 14431 248144
rect 14465 247368 14481 248144
rect 14419 247356 14481 247368
rect 14511 248144 14573 248156
rect 14511 247368 14527 248144
rect 14561 247368 14573 248144
rect 14511 247356 14573 247368
rect 14629 248144 14691 248156
rect 14629 247368 14641 248144
rect 14675 247368 14691 248144
rect 14629 247356 14691 247368
rect 14721 248144 14783 248156
rect 14721 247368 14737 248144
rect 14771 247368 14783 248144
rect 14721 247356 14783 247368
rect 14839 248144 14901 248156
rect 14839 247368 14851 248144
rect 14885 247368 14901 248144
rect 14839 247356 14901 247368
rect 14931 248144 14993 248156
rect 14931 247368 14947 248144
rect 14981 247368 14993 248144
rect 14931 247356 14993 247368
rect 15049 248144 15111 248156
rect 15049 247368 15061 248144
rect 15095 247368 15111 248144
rect 15049 247356 15111 247368
rect 15141 248144 15203 248156
rect 15141 247368 15157 248144
rect 15191 247368 15203 248144
rect 15141 247356 15203 247368
rect 15259 248144 15321 248156
rect 15259 247368 15271 248144
rect 15305 247368 15321 248144
rect 15259 247356 15321 247368
rect 15351 248144 15413 248156
rect 15351 247368 15367 248144
rect 15401 247368 15413 248144
rect 15351 247356 15413 247368
rect 15469 248144 15531 248156
rect 15469 247368 15481 248144
rect 15515 247368 15531 248144
rect 15469 247356 15531 247368
rect 15561 248144 15623 248156
rect 15561 247368 15577 248144
rect 15611 247368 15623 248144
rect 15561 247356 15623 247368
rect 15679 248144 15741 248156
rect 15679 247368 15691 248144
rect 15725 247368 15741 248144
rect 15679 247356 15741 247368
rect 15771 248144 15833 248156
rect 15771 247368 15787 248144
rect 15821 247368 15833 248144
rect 15771 247356 15833 247368
rect 15889 248144 15951 248156
rect 15889 247368 15901 248144
rect 15935 247368 15951 248144
rect 15889 247356 15951 247368
rect 15981 248144 16043 248156
rect 15981 247368 15997 248144
rect 16031 247368 16043 248144
rect 15981 247356 16043 247368
rect 16099 248144 16161 248156
rect 16099 247368 16111 248144
rect 16145 247368 16161 248144
rect 16099 247356 16161 247368
rect 16191 248144 16253 248156
rect 16191 247368 16207 248144
rect 16241 247368 16253 248144
rect 16191 247356 16253 247368
rect 16309 248144 16371 248156
rect 16309 247368 16321 248144
rect 16355 247368 16371 248144
rect 16309 247356 16371 247368
rect 16401 248144 16463 248156
rect 16401 247368 16417 248144
rect 16451 247368 16463 248144
rect 16401 247356 16463 247368
rect 16519 248144 16581 248156
rect 16519 247368 16531 248144
rect 16565 247368 16581 248144
rect 16519 247356 16581 247368
rect 16611 248144 16673 248156
rect 16611 247368 16627 248144
rect 16661 247368 16673 248144
rect 16611 247356 16673 247368
rect 16729 248144 16791 248156
rect 16729 247368 16741 248144
rect 16775 247368 16791 248144
rect 16729 247356 16791 247368
rect 16821 248144 16883 248156
rect 16821 247368 16837 248144
rect 16871 247368 16883 248144
rect 16821 247356 16883 247368
rect 16939 248144 17001 248156
rect 16939 247368 16951 248144
rect 16985 247368 17001 248144
rect 16939 247356 17001 247368
rect 17031 248144 17093 248156
rect 17031 247368 17047 248144
rect 17081 247368 17093 248144
rect 17031 247356 17093 247368
rect 17149 248144 17211 248156
rect 17149 247368 17161 248144
rect 17195 247368 17211 248144
rect 17149 247356 17211 247368
rect 17241 248144 17303 248156
rect 17241 247368 17257 248144
rect 17291 247368 17303 248144
rect 17241 247356 17303 247368
rect 17359 248144 17421 248156
rect 17359 247368 17371 248144
rect 17405 247368 17421 248144
rect 17359 247356 17421 247368
rect 17451 248144 17513 248156
rect 17451 247368 17467 248144
rect 17501 247368 17513 248144
rect 17451 247356 17513 247368
rect 17569 248144 17631 248156
rect 17569 247368 17581 248144
rect 17615 247368 17631 248144
rect 17569 247356 17631 247368
rect 17661 248144 17723 248156
rect 17661 247368 17677 248144
rect 17711 247368 17723 248144
rect 17661 247356 17723 247368
rect 17779 248144 17841 248156
rect 17779 247368 17791 248144
rect 17825 247368 17841 248144
rect 17779 247356 17841 247368
rect 17871 248144 17933 248156
rect 17871 247368 17887 248144
rect 17921 247368 17933 248144
rect 17871 247356 17933 247368
rect 17989 248144 18051 248156
rect 17989 247368 18001 248144
rect 18035 247368 18051 248144
rect 17989 247356 18051 247368
rect 18081 248144 18143 248156
rect 18081 247368 18097 248144
rect 18131 247368 18143 248144
rect 18081 247356 18143 247368
rect 18199 248144 18261 248156
rect 18199 247368 18211 248144
rect 18245 247368 18261 248144
rect 18199 247356 18261 247368
rect 18291 248144 18353 248156
rect 18291 247368 18307 248144
rect 18341 247368 18353 248144
rect 18291 247356 18353 247368
rect 18409 248144 18471 248156
rect 18409 247368 18421 248144
rect 18455 247368 18471 248144
rect 18409 247356 18471 247368
rect 18501 248144 18563 248156
rect 18501 247368 18517 248144
rect 18551 247368 18563 248144
rect 18501 247356 18563 247368
rect 18619 248144 18681 248156
rect 18619 247368 18631 248144
rect 18665 247368 18681 248144
rect 18619 247356 18681 247368
rect 18711 248144 18773 248156
rect 18711 247368 18727 248144
rect 18761 247368 18773 248144
rect 18711 247356 18773 247368
rect 18829 248144 18891 248156
rect 18829 247368 18841 248144
rect 18875 247368 18891 248144
rect 18829 247356 18891 247368
rect 18921 248144 18983 248156
rect 18921 247368 18937 248144
rect 18971 247368 18983 248144
rect 18921 247356 18983 247368
rect 19039 248144 19101 248156
rect 19039 247368 19051 248144
rect 19085 247368 19101 248144
rect 19039 247356 19101 247368
rect 19131 248144 19193 248156
rect 19131 247368 19147 248144
rect 19181 247368 19193 248144
rect 19131 247356 19193 247368
rect 19249 248144 19311 248156
rect 19249 247368 19261 248144
rect 19295 247368 19311 248144
rect 19249 247356 19311 247368
rect 19341 248144 19403 248156
rect 19341 247368 19357 248144
rect 19391 247368 19403 248144
rect 19341 247356 19403 247368
rect 19459 248144 19521 248156
rect 19459 247368 19471 248144
rect 19505 247368 19521 248144
rect 19459 247356 19521 247368
rect 19551 248144 19613 248156
rect 19551 247368 19567 248144
rect 19601 247368 19613 248144
rect 19551 247356 19613 247368
rect 19669 248144 19731 248156
rect 19669 247368 19681 248144
rect 19715 247368 19731 248144
rect 19669 247356 19731 247368
rect 19761 248144 19823 248156
rect 19761 247368 19777 248144
rect 19811 247368 19823 248144
rect 19761 247356 19823 247368
rect 19879 248144 19941 248156
rect 19879 247368 19891 248144
rect 19925 247368 19941 248144
rect 19879 247356 19941 247368
rect 19971 248144 20033 248156
rect 19971 247368 19987 248144
rect 20021 247368 20033 248144
rect 19971 247356 20033 247368
rect 20089 248144 20151 248156
rect 20089 247368 20101 248144
rect 20135 247368 20151 248144
rect 20089 247356 20151 247368
rect 20181 248144 20243 248156
rect 20181 247368 20197 248144
rect 20231 247368 20243 248144
rect 20181 247356 20243 247368
rect 20299 248144 20361 248156
rect 20299 247368 20311 248144
rect 20345 247368 20361 248144
rect 20299 247356 20361 247368
rect 20391 248144 20453 248156
rect 20391 247368 20407 248144
rect 20441 247368 20453 248144
rect 20391 247356 20453 247368
rect 20509 248144 20571 248156
rect 20509 247368 20521 248144
rect 20555 247368 20571 248144
rect 20509 247356 20571 247368
rect 20601 248144 20663 248156
rect 20601 247368 20617 248144
rect 20651 247368 20663 248144
rect 20601 247356 20663 247368
rect 20719 248144 20781 248156
rect 20719 247368 20731 248144
rect 20765 247368 20781 248144
rect 20719 247356 20781 247368
rect 20811 248144 20873 248156
rect 20811 247368 20827 248144
rect 20861 247368 20873 248144
rect 20811 247356 20873 247368
rect 20929 248144 20991 248156
rect 20929 247368 20941 248144
rect 20975 247368 20991 248144
rect 20929 247356 20991 247368
rect 21021 248144 21083 248156
rect 21021 247368 21037 248144
rect 21071 247368 21083 248144
rect 21021 247356 21083 247368
rect 21139 248144 21201 248156
rect 21139 247368 21151 248144
rect 21185 247368 21201 248144
rect 21139 247356 21201 247368
rect 21231 248144 21293 248156
rect 21231 247368 21247 248144
rect 21281 247368 21293 248144
rect 21231 247356 21293 247368
rect 21349 248144 21411 248156
rect 21349 247368 21361 248144
rect 21395 247368 21411 248144
rect 21349 247356 21411 247368
rect 21441 248144 21503 248156
rect 21441 247368 21457 248144
rect 21491 247368 21503 248144
rect 21441 247356 21503 247368
rect 21559 248144 21621 248156
rect 21559 247368 21571 248144
rect 21605 247368 21621 248144
rect 21559 247356 21621 247368
rect 21651 248144 21713 248156
rect 21651 247368 21667 248144
rect 21701 247368 21713 248144
rect 21651 247356 21713 247368
rect 21769 248144 21831 248156
rect 21769 247368 21781 248144
rect 21815 247368 21831 248144
rect 21769 247356 21831 247368
rect 21861 248144 21923 248156
rect 21861 247368 21877 248144
rect 21911 247368 21923 248144
rect 21861 247356 21923 247368
rect 21979 248144 22041 248156
rect 21979 247368 21991 248144
rect 22025 247368 22041 248144
rect 21979 247356 22041 247368
rect 22071 248144 22133 248156
rect 22071 247368 22087 248144
rect 22121 247368 22133 248144
rect 22071 247356 22133 247368
rect 22189 248144 22251 248156
rect 22189 247368 22201 248144
rect 22235 247368 22251 248144
rect 22189 247356 22251 247368
rect 22281 248144 22343 248156
rect 22281 247368 22297 248144
rect 22331 247368 22343 248144
rect 22281 247356 22343 247368
rect 22399 248144 22461 248156
rect 22399 247368 22411 248144
rect 22445 247368 22461 248144
rect 22399 247356 22461 247368
rect 22491 248144 22553 248156
rect 22491 247368 22507 248144
rect 22541 247368 22553 248144
rect 22491 247356 22553 247368
rect 22609 248144 22671 248156
rect 22609 247368 22621 248144
rect 22655 247368 22671 248144
rect 22609 247356 22671 247368
rect 22701 248144 22763 248156
rect 22701 247368 22717 248144
rect 22751 247368 22763 248144
rect 22701 247356 22763 247368
rect 22819 248144 22881 248156
rect 22819 247368 22831 248144
rect 22865 247368 22881 248144
rect 22819 247356 22881 247368
rect 22911 248144 22973 248156
rect 22911 247368 22927 248144
rect 22961 247368 22973 248144
rect 22911 247356 22973 247368
rect 23029 248144 23091 248156
rect 23029 247368 23041 248144
rect 23075 247368 23091 248144
rect 23029 247356 23091 247368
rect 23121 248144 23183 248156
rect 23121 247368 23137 248144
rect 23171 247368 23183 248144
rect 23121 247356 23183 247368
rect 23239 248144 23301 248156
rect 23239 247368 23251 248144
rect 23285 247368 23301 248144
rect 23239 247356 23301 247368
rect 23331 248144 23393 248156
rect 23331 247368 23347 248144
rect 23381 247368 23393 248144
rect 23331 247356 23393 247368
rect 23449 248144 23511 248156
rect 23449 247368 23461 248144
rect 23495 247368 23511 248144
rect 23449 247356 23511 247368
rect 23541 248144 23603 248156
rect 23541 247368 23557 248144
rect 23591 247368 23603 248144
rect 23541 247356 23603 247368
rect 23659 248144 23721 248156
rect 23659 247368 23671 248144
rect 23705 247368 23721 248144
rect 23659 247356 23721 247368
rect 23751 248144 23813 248156
rect 23751 247368 23767 248144
rect 23801 247368 23813 248144
rect 23751 247356 23813 247368
rect 23869 248144 23931 248156
rect 23869 247368 23881 248144
rect 23915 247368 23931 248144
rect 23869 247356 23931 247368
rect 23961 248144 24023 248156
rect 23961 247368 23977 248144
rect 24011 247368 24023 248144
rect 23961 247356 24023 247368
rect 24079 248144 24141 248156
rect 24079 247368 24091 248144
rect 24125 247368 24141 248144
rect 24079 247356 24141 247368
rect 24171 248144 24233 248156
rect 24171 247368 24187 248144
rect 24221 247368 24233 248144
rect 24171 247356 24233 247368
rect 24289 248144 24351 248156
rect 24289 247368 24301 248144
rect 24335 247368 24351 248144
rect 24289 247356 24351 247368
rect 24381 248144 24443 248156
rect 24381 247368 24397 248144
rect 24431 247368 24443 248144
rect 24381 247356 24443 247368
rect 24499 248144 24561 248156
rect 24499 247368 24511 248144
rect 24545 247368 24561 248144
rect 24499 247356 24561 247368
rect 24591 248144 24653 248156
rect 24591 247368 24607 248144
rect 24641 247368 24653 248144
rect 24591 247356 24653 247368
rect 24709 248144 24771 248156
rect 24709 247368 24721 248144
rect 24755 247368 24771 248144
rect 24709 247356 24771 247368
rect 24801 248144 24863 248156
rect 24801 247368 24817 248144
rect 24851 247368 24863 248144
rect 24801 247356 24863 247368
rect 24919 248144 24981 248156
rect 24919 247368 24931 248144
rect 24965 247368 24981 248144
rect 24919 247356 24981 247368
rect 25011 248144 25073 248156
rect 25011 247368 25027 248144
rect 25061 247368 25073 248144
rect 25011 247356 25073 247368
rect 25129 248144 25191 248156
rect 25129 247368 25141 248144
rect 25175 247368 25191 248144
rect 25129 247356 25191 247368
rect 25221 248144 25283 248156
rect 25221 247368 25237 248144
rect 25271 247368 25283 248144
rect 25221 247356 25283 247368
rect 25339 248144 25401 248156
rect 25339 247368 25351 248144
rect 25385 247368 25401 248144
rect 25339 247356 25401 247368
rect 25431 248144 25493 248156
rect 25431 247368 25447 248144
rect 25481 247368 25493 248144
rect 25431 247356 25493 247368
rect 25549 248144 25611 248156
rect 25549 247368 25561 248144
rect 25595 247368 25611 248144
rect 25549 247356 25611 247368
rect 25641 248144 25703 248156
rect 25641 247368 25657 248144
rect 25691 247368 25703 248144
rect 25641 247356 25703 247368
rect 25759 248144 25821 248156
rect 25759 247368 25771 248144
rect 25805 247368 25821 248144
rect 25759 247356 25821 247368
rect 25851 248144 25913 248156
rect 25851 247368 25867 248144
rect 25901 247368 25913 248144
rect 25851 247356 25913 247368
rect 25969 248144 26031 248156
rect 25969 247368 25981 248144
rect 26015 247368 26031 248144
rect 25969 247356 26031 247368
rect 26061 248144 26123 248156
rect 26061 247368 26077 248144
rect 26111 247368 26123 248144
rect 26061 247356 26123 247368
rect 26179 248144 26241 248156
rect 26179 247368 26191 248144
rect 26225 247368 26241 248144
rect 26179 247356 26241 247368
rect 26271 248144 26333 248156
rect 26271 247368 26287 248144
rect 26321 247368 26333 248144
rect 26271 247356 26333 247368
rect 26389 248144 26451 248156
rect 26389 247368 26401 248144
rect 26435 247368 26451 248144
rect 26389 247356 26451 247368
rect 26481 248144 26543 248156
rect 26481 247368 26497 248144
rect 26531 247368 26543 248144
rect 26481 247356 26543 247368
rect 26599 248144 26661 248156
rect 26599 247368 26611 248144
rect 26645 247368 26661 248144
rect 26599 247356 26661 247368
rect 26691 248144 26753 248156
rect 26691 247368 26707 248144
rect 26741 247368 26753 248144
rect 26691 247356 26753 247368
rect 26809 248144 26871 248156
rect 26809 247368 26821 248144
rect 26855 247368 26871 248144
rect 26809 247356 26871 247368
rect 26901 248144 26963 248156
rect 26901 247368 26917 248144
rect 26951 247368 26963 248144
rect 26901 247356 26963 247368
rect 27019 248144 27081 248156
rect 27019 247368 27031 248144
rect 27065 247368 27081 248144
rect 27019 247356 27081 247368
rect 27111 248144 27173 248156
rect 27111 247368 27127 248144
rect 27161 247368 27173 248144
rect 27111 247356 27173 247368
rect 27229 248144 27291 248156
rect 27229 247368 27241 248144
rect 27275 247368 27291 248144
rect 27229 247356 27291 247368
rect 27321 248144 27383 248156
rect 27321 247368 27337 248144
rect 27371 247368 27383 248144
rect 27321 247356 27383 247368
rect -4061 247108 -3999 247120
rect -4061 246332 -4049 247108
rect -4015 246332 -3999 247108
rect -4061 246320 -3999 246332
rect -3969 247108 -3907 247120
rect -3969 246332 -3953 247108
rect -3919 246332 -3907 247108
rect -3969 246320 -3907 246332
rect -3851 247108 -3789 247120
rect -3851 246332 -3839 247108
rect -3805 246332 -3789 247108
rect -3851 246320 -3789 246332
rect -3759 247108 -3697 247120
rect -3759 246332 -3743 247108
rect -3709 246332 -3697 247108
rect -3759 246320 -3697 246332
rect -3641 247108 -3579 247120
rect -3641 246332 -3629 247108
rect -3595 246332 -3579 247108
rect -3641 246320 -3579 246332
rect -3549 247108 -3487 247120
rect -3549 246332 -3533 247108
rect -3499 246332 -3487 247108
rect -3549 246320 -3487 246332
rect -3431 247108 -3369 247120
rect -3431 246332 -3419 247108
rect -3385 246332 -3369 247108
rect -3431 246320 -3369 246332
rect -3339 247108 -3277 247120
rect -3339 246332 -3323 247108
rect -3289 246332 -3277 247108
rect -3339 246320 -3277 246332
rect -3221 247108 -3159 247120
rect -3221 246332 -3209 247108
rect -3175 246332 -3159 247108
rect -3221 246320 -3159 246332
rect -3129 247108 -3067 247120
rect -3129 246332 -3113 247108
rect -3079 246332 -3067 247108
rect -3129 246320 -3067 246332
rect -3011 247108 -2949 247120
rect -3011 246332 -2999 247108
rect -2965 246332 -2949 247108
rect -3011 246320 -2949 246332
rect -2919 247108 -2857 247120
rect -2919 246332 -2903 247108
rect -2869 246332 -2857 247108
rect -2919 246320 -2857 246332
rect -2801 247108 -2739 247120
rect -2801 246332 -2789 247108
rect -2755 246332 -2739 247108
rect -2801 246320 -2739 246332
rect -2709 247108 -2647 247120
rect -2709 246332 -2693 247108
rect -2659 246332 -2647 247108
rect -2709 246320 -2647 246332
rect -2591 247108 -2529 247120
rect -2591 246332 -2579 247108
rect -2545 246332 -2529 247108
rect -2591 246320 -2529 246332
rect -2499 247108 -2437 247120
rect -2499 246332 -2483 247108
rect -2449 246332 -2437 247108
rect -2499 246320 -2437 246332
rect -2381 247108 -2319 247120
rect -2381 246332 -2369 247108
rect -2335 246332 -2319 247108
rect -2381 246320 -2319 246332
rect -2289 247108 -2227 247120
rect -2289 246332 -2273 247108
rect -2239 246332 -2227 247108
rect -2289 246320 -2227 246332
rect -2171 247108 -2109 247120
rect -2171 246332 -2159 247108
rect -2125 246332 -2109 247108
rect -2171 246320 -2109 246332
rect -2079 247108 -2017 247120
rect -2079 246332 -2063 247108
rect -2029 246332 -2017 247108
rect -2079 246320 -2017 246332
rect -1961 247108 -1899 247120
rect -1961 246332 -1949 247108
rect -1915 246332 -1899 247108
rect -1961 246320 -1899 246332
rect -1869 247108 -1807 247120
rect -1869 246332 -1853 247108
rect -1819 246332 -1807 247108
rect -1869 246320 -1807 246332
rect -1751 247108 -1689 247120
rect -1751 246332 -1739 247108
rect -1705 246332 -1689 247108
rect -1751 246320 -1689 246332
rect -1659 247108 -1597 247120
rect -1659 246332 -1643 247108
rect -1609 246332 -1597 247108
rect -1659 246320 -1597 246332
rect -1541 247108 -1479 247120
rect -1541 246332 -1529 247108
rect -1495 246332 -1479 247108
rect -1541 246320 -1479 246332
rect -1449 247108 -1387 247120
rect -1449 246332 -1433 247108
rect -1399 246332 -1387 247108
rect -1449 246320 -1387 246332
rect -1331 247108 -1269 247120
rect -1331 246332 -1319 247108
rect -1285 246332 -1269 247108
rect -1331 246320 -1269 246332
rect -1239 247108 -1177 247120
rect -1239 246332 -1223 247108
rect -1189 246332 -1177 247108
rect -1239 246320 -1177 246332
rect -1121 247108 -1059 247120
rect -1121 246332 -1109 247108
rect -1075 246332 -1059 247108
rect -1121 246320 -1059 246332
rect -1029 247108 -967 247120
rect -1029 246332 -1013 247108
rect -979 246332 -967 247108
rect -1029 246320 -967 246332
rect -911 247108 -849 247120
rect -911 246332 -899 247108
rect -865 246332 -849 247108
rect -911 246320 -849 246332
rect -819 247108 -757 247120
rect -819 246332 -803 247108
rect -769 246332 -757 247108
rect -819 246320 -757 246332
rect -701 247108 -639 247120
rect -701 246332 -689 247108
rect -655 246332 -639 247108
rect -701 246320 -639 246332
rect -609 247108 -547 247120
rect -609 246332 -593 247108
rect -559 246332 -547 247108
rect -609 246320 -547 246332
rect -491 247108 -429 247120
rect -491 246332 -479 247108
rect -445 246332 -429 247108
rect -491 246320 -429 246332
rect -399 247108 -337 247120
rect -399 246332 -383 247108
rect -349 246332 -337 247108
rect -399 246320 -337 246332
rect -281 247108 -219 247120
rect -281 246332 -269 247108
rect -235 246332 -219 247108
rect -281 246320 -219 246332
rect -189 247108 -127 247120
rect -189 246332 -173 247108
rect -139 246332 -127 247108
rect -189 246320 -127 246332
rect -71 247108 -9 247120
rect -71 246332 -59 247108
rect -25 246332 -9 247108
rect -71 246320 -9 246332
rect 21 247108 83 247120
rect 21 246332 37 247108
rect 71 246332 83 247108
rect 21 246320 83 246332
rect 139 247108 201 247120
rect 139 246332 151 247108
rect 185 246332 201 247108
rect 139 246320 201 246332
rect 231 247108 293 247120
rect 231 246332 247 247108
rect 281 246332 293 247108
rect 231 246320 293 246332
rect 349 247108 411 247120
rect 349 246332 361 247108
rect 395 246332 411 247108
rect 349 246320 411 246332
rect 441 247108 503 247120
rect 441 246332 457 247108
rect 491 246332 503 247108
rect 441 246320 503 246332
rect 559 247108 621 247120
rect 559 246332 571 247108
rect 605 246332 621 247108
rect 559 246320 621 246332
rect 651 247108 713 247120
rect 651 246332 667 247108
rect 701 246332 713 247108
rect 651 246320 713 246332
rect 769 247108 831 247120
rect 769 246332 781 247108
rect 815 246332 831 247108
rect 769 246320 831 246332
rect 861 247108 923 247120
rect 861 246332 877 247108
rect 911 246332 923 247108
rect 861 246320 923 246332
rect 979 247108 1041 247120
rect 979 246332 991 247108
rect 1025 246332 1041 247108
rect 979 246320 1041 246332
rect 1071 247108 1133 247120
rect 1071 246332 1087 247108
rect 1121 246332 1133 247108
rect 1071 246320 1133 246332
rect 1189 247108 1251 247120
rect 1189 246332 1201 247108
rect 1235 246332 1251 247108
rect 1189 246320 1251 246332
rect 1281 247108 1343 247120
rect 1281 246332 1297 247108
rect 1331 246332 1343 247108
rect 1281 246320 1343 246332
rect 1399 247108 1461 247120
rect 1399 246332 1411 247108
rect 1445 246332 1461 247108
rect 1399 246320 1461 246332
rect 1491 247108 1553 247120
rect 1491 246332 1507 247108
rect 1541 246332 1553 247108
rect 1491 246320 1553 246332
rect 1609 247108 1671 247120
rect 1609 246332 1621 247108
rect 1655 246332 1671 247108
rect 1609 246320 1671 246332
rect 1701 247108 1763 247120
rect 1701 246332 1717 247108
rect 1751 246332 1763 247108
rect 1701 246320 1763 246332
rect 1819 247108 1881 247120
rect 1819 246332 1831 247108
rect 1865 246332 1881 247108
rect 1819 246320 1881 246332
rect 1911 247108 1973 247120
rect 1911 246332 1927 247108
rect 1961 246332 1973 247108
rect 1911 246320 1973 246332
rect 2029 247108 2091 247120
rect 2029 246332 2041 247108
rect 2075 246332 2091 247108
rect 2029 246320 2091 246332
rect 2121 247108 2183 247120
rect 2121 246332 2137 247108
rect 2171 246332 2183 247108
rect 2121 246320 2183 246332
rect 2239 247108 2301 247120
rect 2239 246332 2251 247108
rect 2285 246332 2301 247108
rect 2239 246320 2301 246332
rect 2331 247108 2393 247120
rect 2331 246332 2347 247108
rect 2381 246332 2393 247108
rect 2331 246320 2393 246332
rect 2449 247108 2511 247120
rect 2449 246332 2461 247108
rect 2495 246332 2511 247108
rect 2449 246320 2511 246332
rect 2541 247108 2603 247120
rect 2541 246332 2557 247108
rect 2591 246332 2603 247108
rect 2541 246320 2603 246332
rect 2659 247108 2721 247120
rect 2659 246332 2671 247108
rect 2705 246332 2721 247108
rect 2659 246320 2721 246332
rect 2751 247108 2813 247120
rect 2751 246332 2767 247108
rect 2801 246332 2813 247108
rect 2751 246320 2813 246332
rect 2869 247108 2931 247120
rect 2869 246332 2881 247108
rect 2915 246332 2931 247108
rect 2869 246320 2931 246332
rect 2961 247108 3023 247120
rect 2961 246332 2977 247108
rect 3011 246332 3023 247108
rect 2961 246320 3023 246332
rect 3079 247108 3141 247120
rect 3079 246332 3091 247108
rect 3125 246332 3141 247108
rect 3079 246320 3141 246332
rect 3171 247108 3233 247120
rect 3171 246332 3187 247108
rect 3221 246332 3233 247108
rect 3171 246320 3233 246332
rect 3289 247108 3351 247120
rect 3289 246332 3301 247108
rect 3335 246332 3351 247108
rect 3289 246320 3351 246332
rect 3381 247108 3443 247120
rect 3381 246332 3397 247108
rect 3431 246332 3443 247108
rect 3381 246320 3443 246332
rect 3499 247108 3561 247120
rect 3499 246332 3511 247108
rect 3545 246332 3561 247108
rect 3499 246320 3561 246332
rect 3591 247108 3653 247120
rect 3591 246332 3607 247108
rect 3641 246332 3653 247108
rect 3591 246320 3653 246332
rect 3709 247108 3771 247120
rect 3709 246332 3721 247108
rect 3755 246332 3771 247108
rect 3709 246320 3771 246332
rect 3801 247108 3863 247120
rect 3801 246332 3817 247108
rect 3851 246332 3863 247108
rect 3801 246320 3863 246332
rect 3919 247108 3981 247120
rect 3919 246332 3931 247108
rect 3965 246332 3981 247108
rect 3919 246320 3981 246332
rect 4011 247108 4073 247120
rect 4011 246332 4027 247108
rect 4061 246332 4073 247108
rect 4011 246320 4073 246332
rect 4129 247108 4191 247120
rect 4129 246332 4141 247108
rect 4175 246332 4191 247108
rect 4129 246320 4191 246332
rect 4221 247108 4283 247120
rect 4221 246332 4237 247108
rect 4271 246332 4283 247108
rect 4221 246320 4283 246332
rect 4339 247108 4401 247120
rect 4339 246332 4351 247108
rect 4385 246332 4401 247108
rect 4339 246320 4401 246332
rect 4431 247108 4493 247120
rect 4431 246332 4447 247108
rect 4481 246332 4493 247108
rect 4431 246320 4493 246332
rect 4549 247108 4611 247120
rect 4549 246332 4561 247108
rect 4595 246332 4611 247108
rect 4549 246320 4611 246332
rect 4641 247108 4703 247120
rect 4641 246332 4657 247108
rect 4691 246332 4703 247108
rect 4641 246320 4703 246332
rect 4759 247108 4821 247120
rect 4759 246332 4771 247108
rect 4805 246332 4821 247108
rect 4759 246320 4821 246332
rect 4851 247108 4913 247120
rect 4851 246332 4867 247108
rect 4901 246332 4913 247108
rect 4851 246320 4913 246332
rect 4969 247108 5031 247120
rect 4969 246332 4981 247108
rect 5015 246332 5031 247108
rect 4969 246320 5031 246332
rect 5061 247108 5123 247120
rect 5061 246332 5077 247108
rect 5111 246332 5123 247108
rect 5061 246320 5123 246332
rect 5179 247108 5241 247120
rect 5179 246332 5191 247108
rect 5225 246332 5241 247108
rect 5179 246320 5241 246332
rect 5271 247108 5333 247120
rect 5271 246332 5287 247108
rect 5321 246332 5333 247108
rect 5271 246320 5333 246332
rect 5389 247108 5451 247120
rect 5389 246332 5401 247108
rect 5435 246332 5451 247108
rect 5389 246320 5451 246332
rect 5481 247108 5543 247120
rect 5481 246332 5497 247108
rect 5531 246332 5543 247108
rect 5481 246320 5543 246332
rect 5599 247108 5661 247120
rect 5599 246332 5611 247108
rect 5645 246332 5661 247108
rect 5599 246320 5661 246332
rect 5691 247108 5753 247120
rect 5691 246332 5707 247108
rect 5741 246332 5753 247108
rect 5691 246320 5753 246332
rect 5809 247108 5871 247120
rect 5809 246332 5821 247108
rect 5855 246332 5871 247108
rect 5809 246320 5871 246332
rect 5901 247108 5963 247120
rect 5901 246332 5917 247108
rect 5951 246332 5963 247108
rect 5901 246320 5963 246332
rect 6019 247108 6081 247120
rect 6019 246332 6031 247108
rect 6065 246332 6081 247108
rect 6019 246320 6081 246332
rect 6111 247108 6173 247120
rect 6111 246332 6127 247108
rect 6161 246332 6173 247108
rect 6111 246320 6173 246332
rect 6229 247108 6291 247120
rect 6229 246332 6241 247108
rect 6275 246332 6291 247108
rect 6229 246320 6291 246332
rect 6321 247108 6383 247120
rect 6321 246332 6337 247108
rect 6371 246332 6383 247108
rect 6321 246320 6383 246332
rect 6439 247108 6501 247120
rect 6439 246332 6451 247108
rect 6485 246332 6501 247108
rect 6439 246320 6501 246332
rect 6531 247108 6593 247120
rect 6531 246332 6547 247108
rect 6581 246332 6593 247108
rect 6531 246320 6593 246332
rect 6649 247108 6711 247120
rect 6649 246332 6661 247108
rect 6695 246332 6711 247108
rect 6649 246320 6711 246332
rect 6741 247108 6803 247120
rect 6741 246332 6757 247108
rect 6791 246332 6803 247108
rect 6741 246320 6803 246332
rect 6859 247108 6921 247120
rect 6859 246332 6871 247108
rect 6905 246332 6921 247108
rect 6859 246320 6921 246332
rect 6951 247108 7013 247120
rect 6951 246332 6967 247108
rect 7001 246332 7013 247108
rect 6951 246320 7013 246332
rect 7069 247108 7131 247120
rect 7069 246332 7081 247108
rect 7115 246332 7131 247108
rect 7069 246320 7131 246332
rect 7161 247108 7223 247120
rect 7161 246332 7177 247108
rect 7211 246332 7223 247108
rect 7161 246320 7223 246332
rect 7279 247108 7341 247120
rect 7279 246332 7291 247108
rect 7325 246332 7341 247108
rect 7279 246320 7341 246332
rect 7371 247108 7433 247120
rect 7371 246332 7387 247108
rect 7421 246332 7433 247108
rect 7371 246320 7433 246332
rect 7489 247108 7551 247120
rect 7489 246332 7501 247108
rect 7535 246332 7551 247108
rect 7489 246320 7551 246332
rect 7581 247108 7643 247120
rect 7581 246332 7597 247108
rect 7631 246332 7643 247108
rect 7581 246320 7643 246332
rect 7699 247108 7761 247120
rect 7699 246332 7711 247108
rect 7745 246332 7761 247108
rect 7699 246320 7761 246332
rect 7791 247108 7853 247120
rect 7791 246332 7807 247108
rect 7841 246332 7853 247108
rect 7791 246320 7853 246332
rect 7909 247108 7971 247120
rect 7909 246332 7921 247108
rect 7955 246332 7971 247108
rect 7909 246320 7971 246332
rect 8001 247108 8063 247120
rect 8001 246332 8017 247108
rect 8051 246332 8063 247108
rect 8001 246320 8063 246332
rect 8119 247108 8181 247120
rect 8119 246332 8131 247108
rect 8165 246332 8181 247108
rect 8119 246320 8181 246332
rect 8211 247108 8273 247120
rect 8211 246332 8227 247108
rect 8261 246332 8273 247108
rect 8211 246320 8273 246332
rect 8329 247108 8391 247120
rect 8329 246332 8341 247108
rect 8375 246332 8391 247108
rect 8329 246320 8391 246332
rect 8421 247108 8483 247120
rect 8421 246332 8437 247108
rect 8471 246332 8483 247108
rect 8421 246320 8483 246332
rect 8539 247108 8601 247120
rect 8539 246332 8551 247108
rect 8585 246332 8601 247108
rect 8539 246320 8601 246332
rect 8631 247108 8693 247120
rect 8631 246332 8647 247108
rect 8681 246332 8693 247108
rect 8631 246320 8693 246332
rect 8749 247108 8811 247120
rect 8749 246332 8761 247108
rect 8795 246332 8811 247108
rect 8749 246320 8811 246332
rect 8841 247108 8903 247120
rect 8841 246332 8857 247108
rect 8891 246332 8903 247108
rect 8841 246320 8903 246332
rect 8959 247108 9021 247120
rect 8959 246332 8971 247108
rect 9005 246332 9021 247108
rect 8959 246320 9021 246332
rect 9051 247108 9113 247120
rect 9051 246332 9067 247108
rect 9101 246332 9113 247108
rect 9051 246320 9113 246332
rect 9169 247108 9231 247120
rect 9169 246332 9181 247108
rect 9215 246332 9231 247108
rect 9169 246320 9231 246332
rect 9261 247108 9323 247120
rect 9261 246332 9277 247108
rect 9311 246332 9323 247108
rect 9261 246320 9323 246332
rect 9379 247108 9441 247120
rect 9379 246332 9391 247108
rect 9425 246332 9441 247108
rect 9379 246320 9441 246332
rect 9471 247108 9533 247120
rect 9471 246332 9487 247108
rect 9521 246332 9533 247108
rect 9471 246320 9533 246332
rect 9589 247108 9651 247120
rect 9589 246332 9601 247108
rect 9635 246332 9651 247108
rect 9589 246320 9651 246332
rect 9681 247108 9743 247120
rect 9681 246332 9697 247108
rect 9731 246332 9743 247108
rect 9681 246320 9743 246332
rect 9799 247108 9861 247120
rect 9799 246332 9811 247108
rect 9845 246332 9861 247108
rect 9799 246320 9861 246332
rect 9891 247108 9953 247120
rect 9891 246332 9907 247108
rect 9941 246332 9953 247108
rect 9891 246320 9953 246332
rect 10009 247108 10071 247120
rect 10009 246332 10021 247108
rect 10055 246332 10071 247108
rect 10009 246320 10071 246332
rect 10101 247108 10163 247120
rect 10101 246332 10117 247108
rect 10151 246332 10163 247108
rect 10101 246320 10163 246332
rect 10219 247108 10281 247120
rect 10219 246332 10231 247108
rect 10265 246332 10281 247108
rect 10219 246320 10281 246332
rect 10311 247108 10373 247120
rect 10311 246332 10327 247108
rect 10361 246332 10373 247108
rect 10311 246320 10373 246332
rect 10429 247108 10491 247120
rect 10429 246332 10441 247108
rect 10475 246332 10491 247108
rect 10429 246320 10491 246332
rect 10521 247108 10583 247120
rect 10521 246332 10537 247108
rect 10571 246332 10583 247108
rect 10521 246320 10583 246332
rect 10639 247108 10701 247120
rect 10639 246332 10651 247108
rect 10685 246332 10701 247108
rect 10639 246320 10701 246332
rect 10731 247108 10793 247120
rect 10731 246332 10747 247108
rect 10781 246332 10793 247108
rect 10731 246320 10793 246332
rect 10849 247108 10911 247120
rect 10849 246332 10861 247108
rect 10895 246332 10911 247108
rect 10849 246320 10911 246332
rect 10941 247108 11003 247120
rect 10941 246332 10957 247108
rect 10991 246332 11003 247108
rect 10941 246320 11003 246332
rect 11059 247108 11121 247120
rect 11059 246332 11071 247108
rect 11105 246332 11121 247108
rect 11059 246320 11121 246332
rect 11151 247108 11213 247120
rect 11151 246332 11167 247108
rect 11201 246332 11213 247108
rect 11151 246320 11213 246332
rect 11269 247108 11331 247120
rect 11269 246332 11281 247108
rect 11315 246332 11331 247108
rect 11269 246320 11331 246332
rect 11361 247108 11423 247120
rect 11361 246332 11377 247108
rect 11411 246332 11423 247108
rect 11361 246320 11423 246332
rect 11479 247108 11541 247120
rect 11479 246332 11491 247108
rect 11525 246332 11541 247108
rect 11479 246320 11541 246332
rect 11571 247108 11633 247120
rect 11571 246332 11587 247108
rect 11621 246332 11633 247108
rect 11571 246320 11633 246332
rect 11689 247108 11751 247120
rect 11689 246332 11701 247108
rect 11735 246332 11751 247108
rect 11689 246320 11751 246332
rect 11781 247108 11843 247120
rect 11781 246332 11797 247108
rect 11831 246332 11843 247108
rect 11781 246320 11843 246332
rect 11899 247108 11961 247120
rect 11899 246332 11911 247108
rect 11945 246332 11961 247108
rect 11899 246320 11961 246332
rect 11991 247108 12053 247120
rect 11991 246332 12007 247108
rect 12041 246332 12053 247108
rect 11991 246320 12053 246332
rect 12109 247108 12171 247120
rect 12109 246332 12121 247108
rect 12155 246332 12171 247108
rect 12109 246320 12171 246332
rect 12201 247108 12263 247120
rect 12201 246332 12217 247108
rect 12251 246332 12263 247108
rect 12201 246320 12263 246332
rect 12319 247108 12381 247120
rect 12319 246332 12331 247108
rect 12365 246332 12381 247108
rect 12319 246320 12381 246332
rect 12411 247108 12473 247120
rect 12411 246332 12427 247108
rect 12461 246332 12473 247108
rect 12411 246320 12473 246332
rect 12529 247108 12591 247120
rect 12529 246332 12541 247108
rect 12575 246332 12591 247108
rect 12529 246320 12591 246332
rect 12621 247108 12683 247120
rect 12621 246332 12637 247108
rect 12671 246332 12683 247108
rect 12621 246320 12683 246332
rect 12739 247108 12801 247120
rect 12739 246332 12751 247108
rect 12785 246332 12801 247108
rect 12739 246320 12801 246332
rect 12831 247108 12893 247120
rect 12831 246332 12847 247108
rect 12881 246332 12893 247108
rect 12831 246320 12893 246332
rect 12949 247108 13011 247120
rect 12949 246332 12961 247108
rect 12995 246332 13011 247108
rect 12949 246320 13011 246332
rect 13041 247108 13103 247120
rect 13041 246332 13057 247108
rect 13091 246332 13103 247108
rect 13041 246320 13103 246332
rect 13159 247108 13221 247120
rect 13159 246332 13171 247108
rect 13205 246332 13221 247108
rect 13159 246320 13221 246332
rect 13251 247108 13313 247120
rect 13251 246332 13267 247108
rect 13301 246332 13313 247108
rect 13251 246320 13313 246332
rect 13369 247108 13431 247120
rect 13369 246332 13381 247108
rect 13415 246332 13431 247108
rect 13369 246320 13431 246332
rect 13461 247108 13523 247120
rect 13461 246332 13477 247108
rect 13511 246332 13523 247108
rect 13461 246320 13523 246332
rect 13579 247108 13641 247120
rect 13579 246332 13591 247108
rect 13625 246332 13641 247108
rect 13579 246320 13641 246332
rect 13671 247108 13733 247120
rect 13671 246332 13687 247108
rect 13721 246332 13733 247108
rect 13671 246320 13733 246332
rect 13789 247108 13851 247120
rect 13789 246332 13801 247108
rect 13835 246332 13851 247108
rect 13789 246320 13851 246332
rect 13881 247108 13943 247120
rect 13881 246332 13897 247108
rect 13931 246332 13943 247108
rect 13881 246320 13943 246332
rect 13999 247108 14061 247120
rect 13999 246332 14011 247108
rect 14045 246332 14061 247108
rect 13999 246320 14061 246332
rect 14091 247108 14153 247120
rect 14091 246332 14107 247108
rect 14141 246332 14153 247108
rect 14091 246320 14153 246332
rect 14209 247108 14271 247120
rect 14209 246332 14221 247108
rect 14255 246332 14271 247108
rect 14209 246320 14271 246332
rect 14301 247108 14363 247120
rect 14301 246332 14317 247108
rect 14351 246332 14363 247108
rect 14301 246320 14363 246332
rect 14419 247108 14481 247120
rect 14419 246332 14431 247108
rect 14465 246332 14481 247108
rect 14419 246320 14481 246332
rect 14511 247108 14573 247120
rect 14511 246332 14527 247108
rect 14561 246332 14573 247108
rect 14511 246320 14573 246332
rect 14629 247108 14691 247120
rect 14629 246332 14641 247108
rect 14675 246332 14691 247108
rect 14629 246320 14691 246332
rect 14721 247108 14783 247120
rect 14721 246332 14737 247108
rect 14771 246332 14783 247108
rect 14721 246320 14783 246332
rect 14839 247108 14901 247120
rect 14839 246332 14851 247108
rect 14885 246332 14901 247108
rect 14839 246320 14901 246332
rect 14931 247108 14993 247120
rect 14931 246332 14947 247108
rect 14981 246332 14993 247108
rect 14931 246320 14993 246332
rect 15049 247108 15111 247120
rect 15049 246332 15061 247108
rect 15095 246332 15111 247108
rect 15049 246320 15111 246332
rect 15141 247108 15203 247120
rect 15141 246332 15157 247108
rect 15191 246332 15203 247108
rect 15141 246320 15203 246332
rect 15259 247108 15321 247120
rect 15259 246332 15271 247108
rect 15305 246332 15321 247108
rect 15259 246320 15321 246332
rect 15351 247108 15413 247120
rect 15351 246332 15367 247108
rect 15401 246332 15413 247108
rect 15351 246320 15413 246332
rect 15469 247108 15531 247120
rect 15469 246332 15481 247108
rect 15515 246332 15531 247108
rect 15469 246320 15531 246332
rect 15561 247108 15623 247120
rect 15561 246332 15577 247108
rect 15611 246332 15623 247108
rect 15561 246320 15623 246332
rect 15679 247108 15741 247120
rect 15679 246332 15691 247108
rect 15725 246332 15741 247108
rect 15679 246320 15741 246332
rect 15771 247108 15833 247120
rect 15771 246332 15787 247108
rect 15821 246332 15833 247108
rect 15771 246320 15833 246332
rect 15889 247108 15951 247120
rect 15889 246332 15901 247108
rect 15935 246332 15951 247108
rect 15889 246320 15951 246332
rect 15981 247108 16043 247120
rect 15981 246332 15997 247108
rect 16031 246332 16043 247108
rect 15981 246320 16043 246332
rect 16099 247108 16161 247120
rect 16099 246332 16111 247108
rect 16145 246332 16161 247108
rect 16099 246320 16161 246332
rect 16191 247108 16253 247120
rect 16191 246332 16207 247108
rect 16241 246332 16253 247108
rect 16191 246320 16253 246332
rect 16309 247108 16371 247120
rect 16309 246332 16321 247108
rect 16355 246332 16371 247108
rect 16309 246320 16371 246332
rect 16401 247108 16463 247120
rect 16401 246332 16417 247108
rect 16451 246332 16463 247108
rect 16401 246320 16463 246332
rect 16519 247108 16581 247120
rect 16519 246332 16531 247108
rect 16565 246332 16581 247108
rect 16519 246320 16581 246332
rect 16611 247108 16673 247120
rect 16611 246332 16627 247108
rect 16661 246332 16673 247108
rect 16611 246320 16673 246332
rect 16729 247108 16791 247120
rect 16729 246332 16741 247108
rect 16775 246332 16791 247108
rect 16729 246320 16791 246332
rect 16821 247108 16883 247120
rect 16821 246332 16837 247108
rect 16871 246332 16883 247108
rect 16821 246320 16883 246332
rect 16939 247108 17001 247120
rect 16939 246332 16951 247108
rect 16985 246332 17001 247108
rect 16939 246320 17001 246332
rect 17031 247108 17093 247120
rect 17031 246332 17047 247108
rect 17081 246332 17093 247108
rect 17031 246320 17093 246332
rect 17149 247108 17211 247120
rect 17149 246332 17161 247108
rect 17195 246332 17211 247108
rect 17149 246320 17211 246332
rect 17241 247108 17303 247120
rect 17241 246332 17257 247108
rect 17291 246332 17303 247108
rect 17241 246320 17303 246332
rect 17359 247108 17421 247120
rect 17359 246332 17371 247108
rect 17405 246332 17421 247108
rect 17359 246320 17421 246332
rect 17451 247108 17513 247120
rect 17451 246332 17467 247108
rect 17501 246332 17513 247108
rect 17451 246320 17513 246332
rect 17569 247108 17631 247120
rect 17569 246332 17581 247108
rect 17615 246332 17631 247108
rect 17569 246320 17631 246332
rect 17661 247108 17723 247120
rect 17661 246332 17677 247108
rect 17711 246332 17723 247108
rect 17661 246320 17723 246332
rect 17779 247108 17841 247120
rect 17779 246332 17791 247108
rect 17825 246332 17841 247108
rect 17779 246320 17841 246332
rect 17871 247108 17933 247120
rect 17871 246332 17887 247108
rect 17921 246332 17933 247108
rect 17871 246320 17933 246332
rect 17989 247108 18051 247120
rect 17989 246332 18001 247108
rect 18035 246332 18051 247108
rect 17989 246320 18051 246332
rect 18081 247108 18143 247120
rect 18081 246332 18097 247108
rect 18131 246332 18143 247108
rect 18081 246320 18143 246332
rect 18199 247108 18261 247120
rect 18199 246332 18211 247108
rect 18245 246332 18261 247108
rect 18199 246320 18261 246332
rect 18291 247108 18353 247120
rect 18291 246332 18307 247108
rect 18341 246332 18353 247108
rect 18291 246320 18353 246332
rect 18409 247108 18471 247120
rect 18409 246332 18421 247108
rect 18455 246332 18471 247108
rect 18409 246320 18471 246332
rect 18501 247108 18563 247120
rect 18501 246332 18517 247108
rect 18551 246332 18563 247108
rect 18501 246320 18563 246332
rect 18619 247108 18681 247120
rect 18619 246332 18631 247108
rect 18665 246332 18681 247108
rect 18619 246320 18681 246332
rect 18711 247108 18773 247120
rect 18711 246332 18727 247108
rect 18761 246332 18773 247108
rect 18711 246320 18773 246332
rect 18829 247108 18891 247120
rect 18829 246332 18841 247108
rect 18875 246332 18891 247108
rect 18829 246320 18891 246332
rect 18921 247108 18983 247120
rect 18921 246332 18937 247108
rect 18971 246332 18983 247108
rect 18921 246320 18983 246332
rect 19039 247108 19101 247120
rect 19039 246332 19051 247108
rect 19085 246332 19101 247108
rect 19039 246320 19101 246332
rect 19131 247108 19193 247120
rect 19131 246332 19147 247108
rect 19181 246332 19193 247108
rect 19131 246320 19193 246332
rect 19249 247108 19311 247120
rect 19249 246332 19261 247108
rect 19295 246332 19311 247108
rect 19249 246320 19311 246332
rect 19341 247108 19403 247120
rect 19341 246332 19357 247108
rect 19391 246332 19403 247108
rect 19341 246320 19403 246332
rect 19459 247108 19521 247120
rect 19459 246332 19471 247108
rect 19505 246332 19521 247108
rect 19459 246320 19521 246332
rect 19551 247108 19613 247120
rect 19551 246332 19567 247108
rect 19601 246332 19613 247108
rect 19551 246320 19613 246332
rect 19669 247108 19731 247120
rect 19669 246332 19681 247108
rect 19715 246332 19731 247108
rect 19669 246320 19731 246332
rect 19761 247108 19823 247120
rect 19761 246332 19777 247108
rect 19811 246332 19823 247108
rect 19761 246320 19823 246332
rect 19879 247108 19941 247120
rect 19879 246332 19891 247108
rect 19925 246332 19941 247108
rect 19879 246320 19941 246332
rect 19971 247108 20033 247120
rect 19971 246332 19987 247108
rect 20021 246332 20033 247108
rect 19971 246320 20033 246332
rect 20089 247108 20151 247120
rect 20089 246332 20101 247108
rect 20135 246332 20151 247108
rect 20089 246320 20151 246332
rect 20181 247108 20243 247120
rect 20181 246332 20197 247108
rect 20231 246332 20243 247108
rect 20181 246320 20243 246332
rect 20299 247108 20361 247120
rect 20299 246332 20311 247108
rect 20345 246332 20361 247108
rect 20299 246320 20361 246332
rect 20391 247108 20453 247120
rect 20391 246332 20407 247108
rect 20441 246332 20453 247108
rect 20391 246320 20453 246332
rect 20509 247108 20571 247120
rect 20509 246332 20521 247108
rect 20555 246332 20571 247108
rect 20509 246320 20571 246332
rect 20601 247108 20663 247120
rect 20601 246332 20617 247108
rect 20651 246332 20663 247108
rect 20601 246320 20663 246332
rect 20719 247108 20781 247120
rect 20719 246332 20731 247108
rect 20765 246332 20781 247108
rect 20719 246320 20781 246332
rect 20811 247108 20873 247120
rect 20811 246332 20827 247108
rect 20861 246332 20873 247108
rect 20811 246320 20873 246332
rect 20929 247108 20991 247120
rect 20929 246332 20941 247108
rect 20975 246332 20991 247108
rect 20929 246320 20991 246332
rect 21021 247108 21083 247120
rect 21021 246332 21037 247108
rect 21071 246332 21083 247108
rect 21021 246320 21083 246332
rect 21139 247108 21201 247120
rect 21139 246332 21151 247108
rect 21185 246332 21201 247108
rect 21139 246320 21201 246332
rect 21231 247108 21293 247120
rect 21231 246332 21247 247108
rect 21281 246332 21293 247108
rect 21231 246320 21293 246332
rect 21349 247108 21411 247120
rect 21349 246332 21361 247108
rect 21395 246332 21411 247108
rect 21349 246320 21411 246332
rect 21441 247108 21503 247120
rect 21441 246332 21457 247108
rect 21491 246332 21503 247108
rect 21441 246320 21503 246332
rect 21559 247108 21621 247120
rect 21559 246332 21571 247108
rect 21605 246332 21621 247108
rect 21559 246320 21621 246332
rect 21651 247108 21713 247120
rect 21651 246332 21667 247108
rect 21701 246332 21713 247108
rect 21651 246320 21713 246332
rect 21769 247108 21831 247120
rect 21769 246332 21781 247108
rect 21815 246332 21831 247108
rect 21769 246320 21831 246332
rect 21861 247108 21923 247120
rect 21861 246332 21877 247108
rect 21911 246332 21923 247108
rect 21861 246320 21923 246332
rect 21979 247108 22041 247120
rect 21979 246332 21991 247108
rect 22025 246332 22041 247108
rect 21979 246320 22041 246332
rect 22071 247108 22133 247120
rect 22071 246332 22087 247108
rect 22121 246332 22133 247108
rect 22071 246320 22133 246332
rect 22189 247108 22251 247120
rect 22189 246332 22201 247108
rect 22235 246332 22251 247108
rect 22189 246320 22251 246332
rect 22281 247108 22343 247120
rect 22281 246332 22297 247108
rect 22331 246332 22343 247108
rect 22281 246320 22343 246332
rect 22399 247108 22461 247120
rect 22399 246332 22411 247108
rect 22445 246332 22461 247108
rect 22399 246320 22461 246332
rect 22491 247108 22553 247120
rect 22491 246332 22507 247108
rect 22541 246332 22553 247108
rect 22491 246320 22553 246332
rect 22609 247108 22671 247120
rect 22609 246332 22621 247108
rect 22655 246332 22671 247108
rect 22609 246320 22671 246332
rect 22701 247108 22763 247120
rect 22701 246332 22717 247108
rect 22751 246332 22763 247108
rect 22701 246320 22763 246332
rect 22819 247108 22881 247120
rect 22819 246332 22831 247108
rect 22865 246332 22881 247108
rect 22819 246320 22881 246332
rect 22911 247108 22973 247120
rect 22911 246332 22927 247108
rect 22961 246332 22973 247108
rect 22911 246320 22973 246332
rect 23029 247108 23091 247120
rect 23029 246332 23041 247108
rect 23075 246332 23091 247108
rect 23029 246320 23091 246332
rect 23121 247108 23183 247120
rect 23121 246332 23137 247108
rect 23171 246332 23183 247108
rect 23121 246320 23183 246332
rect 23239 247108 23301 247120
rect 23239 246332 23251 247108
rect 23285 246332 23301 247108
rect 23239 246320 23301 246332
rect 23331 247108 23393 247120
rect 23331 246332 23347 247108
rect 23381 246332 23393 247108
rect 23331 246320 23393 246332
rect 23449 247108 23511 247120
rect 23449 246332 23461 247108
rect 23495 246332 23511 247108
rect 23449 246320 23511 246332
rect 23541 247108 23603 247120
rect 23541 246332 23557 247108
rect 23591 246332 23603 247108
rect 23541 246320 23603 246332
rect 23659 247108 23721 247120
rect 23659 246332 23671 247108
rect 23705 246332 23721 247108
rect 23659 246320 23721 246332
rect 23751 247108 23813 247120
rect 23751 246332 23767 247108
rect 23801 246332 23813 247108
rect 23751 246320 23813 246332
rect 23869 247108 23931 247120
rect 23869 246332 23881 247108
rect 23915 246332 23931 247108
rect 23869 246320 23931 246332
rect 23961 247108 24023 247120
rect 23961 246332 23977 247108
rect 24011 246332 24023 247108
rect 23961 246320 24023 246332
rect 24079 247108 24141 247120
rect 24079 246332 24091 247108
rect 24125 246332 24141 247108
rect 24079 246320 24141 246332
rect 24171 247108 24233 247120
rect 24171 246332 24187 247108
rect 24221 246332 24233 247108
rect 24171 246320 24233 246332
rect 24289 247108 24351 247120
rect 24289 246332 24301 247108
rect 24335 246332 24351 247108
rect 24289 246320 24351 246332
rect 24381 247108 24443 247120
rect 24381 246332 24397 247108
rect 24431 246332 24443 247108
rect 24381 246320 24443 246332
rect 24499 247108 24561 247120
rect 24499 246332 24511 247108
rect 24545 246332 24561 247108
rect 24499 246320 24561 246332
rect 24591 247108 24653 247120
rect 24591 246332 24607 247108
rect 24641 246332 24653 247108
rect 24591 246320 24653 246332
rect 24709 247108 24771 247120
rect 24709 246332 24721 247108
rect 24755 246332 24771 247108
rect 24709 246320 24771 246332
rect 24801 247108 24863 247120
rect 24801 246332 24817 247108
rect 24851 246332 24863 247108
rect 24801 246320 24863 246332
rect 24919 247108 24981 247120
rect 24919 246332 24931 247108
rect 24965 246332 24981 247108
rect 24919 246320 24981 246332
rect 25011 247108 25073 247120
rect 25011 246332 25027 247108
rect 25061 246332 25073 247108
rect 25011 246320 25073 246332
rect 25129 247108 25191 247120
rect 25129 246332 25141 247108
rect 25175 246332 25191 247108
rect 25129 246320 25191 246332
rect 25221 247108 25283 247120
rect 25221 246332 25237 247108
rect 25271 246332 25283 247108
rect 25221 246320 25283 246332
rect 25339 247108 25401 247120
rect 25339 246332 25351 247108
rect 25385 246332 25401 247108
rect 25339 246320 25401 246332
rect 25431 247108 25493 247120
rect 25431 246332 25447 247108
rect 25481 246332 25493 247108
rect 25431 246320 25493 246332
rect 25549 247108 25611 247120
rect 25549 246332 25561 247108
rect 25595 246332 25611 247108
rect 25549 246320 25611 246332
rect 25641 247108 25703 247120
rect 25641 246332 25657 247108
rect 25691 246332 25703 247108
rect 25641 246320 25703 246332
rect 25759 247108 25821 247120
rect 25759 246332 25771 247108
rect 25805 246332 25821 247108
rect 25759 246320 25821 246332
rect 25851 247108 25913 247120
rect 25851 246332 25867 247108
rect 25901 246332 25913 247108
rect 25851 246320 25913 246332
rect 25969 247108 26031 247120
rect 25969 246332 25981 247108
rect 26015 246332 26031 247108
rect 25969 246320 26031 246332
rect 26061 247108 26123 247120
rect 26061 246332 26077 247108
rect 26111 246332 26123 247108
rect 26061 246320 26123 246332
rect 26179 247108 26241 247120
rect 26179 246332 26191 247108
rect 26225 246332 26241 247108
rect 26179 246320 26241 246332
rect 26271 247108 26333 247120
rect 26271 246332 26287 247108
rect 26321 246332 26333 247108
rect 26271 246320 26333 246332
rect 26389 247108 26451 247120
rect 26389 246332 26401 247108
rect 26435 246332 26451 247108
rect 26389 246320 26451 246332
rect 26481 247108 26543 247120
rect 26481 246332 26497 247108
rect 26531 246332 26543 247108
rect 26481 246320 26543 246332
rect 26599 247108 26661 247120
rect 26599 246332 26611 247108
rect 26645 246332 26661 247108
rect 26599 246320 26661 246332
rect 26691 247108 26753 247120
rect 26691 246332 26707 247108
rect 26741 246332 26753 247108
rect 26691 246320 26753 246332
rect 26809 247108 26871 247120
rect 26809 246332 26821 247108
rect 26855 246332 26871 247108
rect 26809 246320 26871 246332
rect 26901 247108 26963 247120
rect 26901 246332 26917 247108
rect 26951 246332 26963 247108
rect 26901 246320 26963 246332
rect 27019 247108 27081 247120
rect 27019 246332 27031 247108
rect 27065 246332 27081 247108
rect 27019 246320 27081 246332
rect 27111 247108 27173 247120
rect 27111 246332 27127 247108
rect 27161 246332 27173 247108
rect 27111 246320 27173 246332
rect 27229 247108 27291 247120
rect 27229 246332 27241 247108
rect 27275 246332 27291 247108
rect 27229 246320 27291 246332
rect 27321 247108 27383 247120
rect 27321 246332 27337 247108
rect 27371 246332 27383 247108
rect 27321 246320 27383 246332
rect -4061 246072 -3999 246084
rect -4061 245296 -4049 246072
rect -4015 245296 -3999 246072
rect -4061 245284 -3999 245296
rect -3969 246072 -3907 246084
rect -3969 245296 -3953 246072
rect -3919 245296 -3907 246072
rect -3969 245284 -3907 245296
rect -3851 246072 -3789 246084
rect -3851 245296 -3839 246072
rect -3805 245296 -3789 246072
rect -3851 245284 -3789 245296
rect -3759 246072 -3697 246084
rect -3759 245296 -3743 246072
rect -3709 245296 -3697 246072
rect -3759 245284 -3697 245296
rect -3641 246072 -3579 246084
rect -3641 245296 -3629 246072
rect -3595 245296 -3579 246072
rect -3641 245284 -3579 245296
rect -3549 246072 -3487 246084
rect -3549 245296 -3533 246072
rect -3499 245296 -3487 246072
rect -3549 245284 -3487 245296
rect -3431 246072 -3369 246084
rect -3431 245296 -3419 246072
rect -3385 245296 -3369 246072
rect -3431 245284 -3369 245296
rect -3339 246072 -3277 246084
rect -3339 245296 -3323 246072
rect -3289 245296 -3277 246072
rect -3339 245284 -3277 245296
rect -3221 246072 -3159 246084
rect -3221 245296 -3209 246072
rect -3175 245296 -3159 246072
rect -3221 245284 -3159 245296
rect -3129 246072 -3067 246084
rect -3129 245296 -3113 246072
rect -3079 245296 -3067 246072
rect -3129 245284 -3067 245296
rect -3011 246072 -2949 246084
rect -3011 245296 -2999 246072
rect -2965 245296 -2949 246072
rect -3011 245284 -2949 245296
rect -2919 246072 -2857 246084
rect -2919 245296 -2903 246072
rect -2869 245296 -2857 246072
rect -2919 245284 -2857 245296
rect -2801 246072 -2739 246084
rect -2801 245296 -2789 246072
rect -2755 245296 -2739 246072
rect -2801 245284 -2739 245296
rect -2709 246072 -2647 246084
rect -2709 245296 -2693 246072
rect -2659 245296 -2647 246072
rect -2709 245284 -2647 245296
rect -2591 246072 -2529 246084
rect -2591 245296 -2579 246072
rect -2545 245296 -2529 246072
rect -2591 245284 -2529 245296
rect -2499 246072 -2437 246084
rect -2499 245296 -2483 246072
rect -2449 245296 -2437 246072
rect -2499 245284 -2437 245296
rect -2381 246072 -2319 246084
rect -2381 245296 -2369 246072
rect -2335 245296 -2319 246072
rect -2381 245284 -2319 245296
rect -2289 246072 -2227 246084
rect -2289 245296 -2273 246072
rect -2239 245296 -2227 246072
rect -2289 245284 -2227 245296
rect -2171 246072 -2109 246084
rect -2171 245296 -2159 246072
rect -2125 245296 -2109 246072
rect -2171 245284 -2109 245296
rect -2079 246072 -2017 246084
rect -2079 245296 -2063 246072
rect -2029 245296 -2017 246072
rect -2079 245284 -2017 245296
rect -1961 246072 -1899 246084
rect -1961 245296 -1949 246072
rect -1915 245296 -1899 246072
rect -1961 245284 -1899 245296
rect -1869 246072 -1807 246084
rect -1869 245296 -1853 246072
rect -1819 245296 -1807 246072
rect -1869 245284 -1807 245296
rect -1751 246072 -1689 246084
rect -1751 245296 -1739 246072
rect -1705 245296 -1689 246072
rect -1751 245284 -1689 245296
rect -1659 246072 -1597 246084
rect -1659 245296 -1643 246072
rect -1609 245296 -1597 246072
rect -1659 245284 -1597 245296
rect -1541 246072 -1479 246084
rect -1541 245296 -1529 246072
rect -1495 245296 -1479 246072
rect -1541 245284 -1479 245296
rect -1449 246072 -1387 246084
rect -1449 245296 -1433 246072
rect -1399 245296 -1387 246072
rect -1449 245284 -1387 245296
rect -1331 246072 -1269 246084
rect -1331 245296 -1319 246072
rect -1285 245296 -1269 246072
rect -1331 245284 -1269 245296
rect -1239 246072 -1177 246084
rect -1239 245296 -1223 246072
rect -1189 245296 -1177 246072
rect -1239 245284 -1177 245296
rect -1121 246072 -1059 246084
rect -1121 245296 -1109 246072
rect -1075 245296 -1059 246072
rect -1121 245284 -1059 245296
rect -1029 246072 -967 246084
rect -1029 245296 -1013 246072
rect -979 245296 -967 246072
rect -1029 245284 -967 245296
rect -911 246072 -849 246084
rect -911 245296 -899 246072
rect -865 245296 -849 246072
rect -911 245284 -849 245296
rect -819 246072 -757 246084
rect -819 245296 -803 246072
rect -769 245296 -757 246072
rect -819 245284 -757 245296
rect -701 246072 -639 246084
rect -701 245296 -689 246072
rect -655 245296 -639 246072
rect -701 245284 -639 245296
rect -609 246072 -547 246084
rect -609 245296 -593 246072
rect -559 245296 -547 246072
rect -609 245284 -547 245296
rect -491 246072 -429 246084
rect -491 245296 -479 246072
rect -445 245296 -429 246072
rect -491 245284 -429 245296
rect -399 246072 -337 246084
rect -399 245296 -383 246072
rect -349 245296 -337 246072
rect -399 245284 -337 245296
rect -281 246072 -219 246084
rect -281 245296 -269 246072
rect -235 245296 -219 246072
rect -281 245284 -219 245296
rect -189 246072 -127 246084
rect -189 245296 -173 246072
rect -139 245296 -127 246072
rect -189 245284 -127 245296
rect -71 246072 -9 246084
rect -71 245296 -59 246072
rect -25 245296 -9 246072
rect -71 245284 -9 245296
rect 21 246072 83 246084
rect 21 245296 37 246072
rect 71 245296 83 246072
rect 21 245284 83 245296
rect 139 246072 201 246084
rect 139 245296 151 246072
rect 185 245296 201 246072
rect 139 245284 201 245296
rect 231 246072 293 246084
rect 231 245296 247 246072
rect 281 245296 293 246072
rect 231 245284 293 245296
rect 349 246072 411 246084
rect 349 245296 361 246072
rect 395 245296 411 246072
rect 349 245284 411 245296
rect 441 246072 503 246084
rect 441 245296 457 246072
rect 491 245296 503 246072
rect 441 245284 503 245296
rect 559 246072 621 246084
rect 559 245296 571 246072
rect 605 245296 621 246072
rect 559 245284 621 245296
rect 651 246072 713 246084
rect 651 245296 667 246072
rect 701 245296 713 246072
rect 651 245284 713 245296
rect 769 246072 831 246084
rect 769 245296 781 246072
rect 815 245296 831 246072
rect 769 245284 831 245296
rect 861 246072 923 246084
rect 861 245296 877 246072
rect 911 245296 923 246072
rect 861 245284 923 245296
rect 979 246072 1041 246084
rect 979 245296 991 246072
rect 1025 245296 1041 246072
rect 979 245284 1041 245296
rect 1071 246072 1133 246084
rect 1071 245296 1087 246072
rect 1121 245296 1133 246072
rect 1071 245284 1133 245296
rect 1189 246072 1251 246084
rect 1189 245296 1201 246072
rect 1235 245296 1251 246072
rect 1189 245284 1251 245296
rect 1281 246072 1343 246084
rect 1281 245296 1297 246072
rect 1331 245296 1343 246072
rect 1281 245284 1343 245296
rect 1399 246072 1461 246084
rect 1399 245296 1411 246072
rect 1445 245296 1461 246072
rect 1399 245284 1461 245296
rect 1491 246072 1553 246084
rect 1491 245296 1507 246072
rect 1541 245296 1553 246072
rect 1491 245284 1553 245296
rect 1609 246072 1671 246084
rect 1609 245296 1621 246072
rect 1655 245296 1671 246072
rect 1609 245284 1671 245296
rect 1701 246072 1763 246084
rect 1701 245296 1717 246072
rect 1751 245296 1763 246072
rect 1701 245284 1763 245296
rect 1819 246072 1881 246084
rect 1819 245296 1831 246072
rect 1865 245296 1881 246072
rect 1819 245284 1881 245296
rect 1911 246072 1973 246084
rect 1911 245296 1927 246072
rect 1961 245296 1973 246072
rect 1911 245284 1973 245296
rect 2029 246072 2091 246084
rect 2029 245296 2041 246072
rect 2075 245296 2091 246072
rect 2029 245284 2091 245296
rect 2121 246072 2183 246084
rect 2121 245296 2137 246072
rect 2171 245296 2183 246072
rect 2121 245284 2183 245296
rect 2239 246072 2301 246084
rect 2239 245296 2251 246072
rect 2285 245296 2301 246072
rect 2239 245284 2301 245296
rect 2331 246072 2393 246084
rect 2331 245296 2347 246072
rect 2381 245296 2393 246072
rect 2331 245284 2393 245296
rect 2449 246072 2511 246084
rect 2449 245296 2461 246072
rect 2495 245296 2511 246072
rect 2449 245284 2511 245296
rect 2541 246072 2603 246084
rect 2541 245296 2557 246072
rect 2591 245296 2603 246072
rect 2541 245284 2603 245296
rect 2659 246072 2721 246084
rect 2659 245296 2671 246072
rect 2705 245296 2721 246072
rect 2659 245284 2721 245296
rect 2751 246072 2813 246084
rect 2751 245296 2767 246072
rect 2801 245296 2813 246072
rect 2751 245284 2813 245296
rect 2869 246072 2931 246084
rect 2869 245296 2881 246072
rect 2915 245296 2931 246072
rect 2869 245284 2931 245296
rect 2961 246072 3023 246084
rect 2961 245296 2977 246072
rect 3011 245296 3023 246072
rect 2961 245284 3023 245296
rect 3079 246072 3141 246084
rect 3079 245296 3091 246072
rect 3125 245296 3141 246072
rect 3079 245284 3141 245296
rect 3171 246072 3233 246084
rect 3171 245296 3187 246072
rect 3221 245296 3233 246072
rect 3171 245284 3233 245296
rect 3289 246072 3351 246084
rect 3289 245296 3301 246072
rect 3335 245296 3351 246072
rect 3289 245284 3351 245296
rect 3381 246072 3443 246084
rect 3381 245296 3397 246072
rect 3431 245296 3443 246072
rect 3381 245284 3443 245296
rect 3499 246072 3561 246084
rect 3499 245296 3511 246072
rect 3545 245296 3561 246072
rect 3499 245284 3561 245296
rect 3591 246072 3653 246084
rect 3591 245296 3607 246072
rect 3641 245296 3653 246072
rect 3591 245284 3653 245296
rect 3709 246072 3771 246084
rect 3709 245296 3721 246072
rect 3755 245296 3771 246072
rect 3709 245284 3771 245296
rect 3801 246072 3863 246084
rect 3801 245296 3817 246072
rect 3851 245296 3863 246072
rect 3801 245284 3863 245296
rect 3919 246072 3981 246084
rect 3919 245296 3931 246072
rect 3965 245296 3981 246072
rect 3919 245284 3981 245296
rect 4011 246072 4073 246084
rect 4011 245296 4027 246072
rect 4061 245296 4073 246072
rect 4011 245284 4073 245296
rect 4129 246072 4191 246084
rect 4129 245296 4141 246072
rect 4175 245296 4191 246072
rect 4129 245284 4191 245296
rect 4221 246072 4283 246084
rect 4221 245296 4237 246072
rect 4271 245296 4283 246072
rect 4221 245284 4283 245296
rect 4339 246072 4401 246084
rect 4339 245296 4351 246072
rect 4385 245296 4401 246072
rect 4339 245284 4401 245296
rect 4431 246072 4493 246084
rect 4431 245296 4447 246072
rect 4481 245296 4493 246072
rect 4431 245284 4493 245296
rect 4549 246072 4611 246084
rect 4549 245296 4561 246072
rect 4595 245296 4611 246072
rect 4549 245284 4611 245296
rect 4641 246072 4703 246084
rect 4641 245296 4657 246072
rect 4691 245296 4703 246072
rect 4641 245284 4703 245296
rect 4759 246072 4821 246084
rect 4759 245296 4771 246072
rect 4805 245296 4821 246072
rect 4759 245284 4821 245296
rect 4851 246072 4913 246084
rect 4851 245296 4867 246072
rect 4901 245296 4913 246072
rect 4851 245284 4913 245296
rect 4969 246072 5031 246084
rect 4969 245296 4981 246072
rect 5015 245296 5031 246072
rect 4969 245284 5031 245296
rect 5061 246072 5123 246084
rect 5061 245296 5077 246072
rect 5111 245296 5123 246072
rect 5061 245284 5123 245296
rect 5179 246072 5241 246084
rect 5179 245296 5191 246072
rect 5225 245296 5241 246072
rect 5179 245284 5241 245296
rect 5271 246072 5333 246084
rect 5271 245296 5287 246072
rect 5321 245296 5333 246072
rect 5271 245284 5333 245296
rect 5389 246072 5451 246084
rect 5389 245296 5401 246072
rect 5435 245296 5451 246072
rect 5389 245284 5451 245296
rect 5481 246072 5543 246084
rect 5481 245296 5497 246072
rect 5531 245296 5543 246072
rect 5481 245284 5543 245296
rect 5599 246072 5661 246084
rect 5599 245296 5611 246072
rect 5645 245296 5661 246072
rect 5599 245284 5661 245296
rect 5691 246072 5753 246084
rect 5691 245296 5707 246072
rect 5741 245296 5753 246072
rect 5691 245284 5753 245296
rect 5809 246072 5871 246084
rect 5809 245296 5821 246072
rect 5855 245296 5871 246072
rect 5809 245284 5871 245296
rect 5901 246072 5963 246084
rect 5901 245296 5917 246072
rect 5951 245296 5963 246072
rect 5901 245284 5963 245296
rect 6019 246072 6081 246084
rect 6019 245296 6031 246072
rect 6065 245296 6081 246072
rect 6019 245284 6081 245296
rect 6111 246072 6173 246084
rect 6111 245296 6127 246072
rect 6161 245296 6173 246072
rect 6111 245284 6173 245296
rect 6229 246072 6291 246084
rect 6229 245296 6241 246072
rect 6275 245296 6291 246072
rect 6229 245284 6291 245296
rect 6321 246072 6383 246084
rect 6321 245296 6337 246072
rect 6371 245296 6383 246072
rect 6321 245284 6383 245296
rect 6439 246072 6501 246084
rect 6439 245296 6451 246072
rect 6485 245296 6501 246072
rect 6439 245284 6501 245296
rect 6531 246072 6593 246084
rect 6531 245296 6547 246072
rect 6581 245296 6593 246072
rect 6531 245284 6593 245296
rect 6649 246072 6711 246084
rect 6649 245296 6661 246072
rect 6695 245296 6711 246072
rect 6649 245284 6711 245296
rect 6741 246072 6803 246084
rect 6741 245296 6757 246072
rect 6791 245296 6803 246072
rect 6741 245284 6803 245296
rect 6859 246072 6921 246084
rect 6859 245296 6871 246072
rect 6905 245296 6921 246072
rect 6859 245284 6921 245296
rect 6951 246072 7013 246084
rect 6951 245296 6967 246072
rect 7001 245296 7013 246072
rect 6951 245284 7013 245296
rect 7069 246072 7131 246084
rect 7069 245296 7081 246072
rect 7115 245296 7131 246072
rect 7069 245284 7131 245296
rect 7161 246072 7223 246084
rect 7161 245296 7177 246072
rect 7211 245296 7223 246072
rect 7161 245284 7223 245296
rect 7279 246072 7341 246084
rect 7279 245296 7291 246072
rect 7325 245296 7341 246072
rect 7279 245284 7341 245296
rect 7371 246072 7433 246084
rect 7371 245296 7387 246072
rect 7421 245296 7433 246072
rect 7371 245284 7433 245296
rect 7489 246072 7551 246084
rect 7489 245296 7501 246072
rect 7535 245296 7551 246072
rect 7489 245284 7551 245296
rect 7581 246072 7643 246084
rect 7581 245296 7597 246072
rect 7631 245296 7643 246072
rect 7581 245284 7643 245296
rect 7699 246072 7761 246084
rect 7699 245296 7711 246072
rect 7745 245296 7761 246072
rect 7699 245284 7761 245296
rect 7791 246072 7853 246084
rect 7791 245296 7807 246072
rect 7841 245296 7853 246072
rect 7791 245284 7853 245296
rect 7909 246072 7971 246084
rect 7909 245296 7921 246072
rect 7955 245296 7971 246072
rect 7909 245284 7971 245296
rect 8001 246072 8063 246084
rect 8001 245296 8017 246072
rect 8051 245296 8063 246072
rect 8001 245284 8063 245296
rect 8119 246072 8181 246084
rect 8119 245296 8131 246072
rect 8165 245296 8181 246072
rect 8119 245284 8181 245296
rect 8211 246072 8273 246084
rect 8211 245296 8227 246072
rect 8261 245296 8273 246072
rect 8211 245284 8273 245296
rect 8329 246072 8391 246084
rect 8329 245296 8341 246072
rect 8375 245296 8391 246072
rect 8329 245284 8391 245296
rect 8421 246072 8483 246084
rect 8421 245296 8437 246072
rect 8471 245296 8483 246072
rect 8421 245284 8483 245296
rect 8539 246072 8601 246084
rect 8539 245296 8551 246072
rect 8585 245296 8601 246072
rect 8539 245284 8601 245296
rect 8631 246072 8693 246084
rect 8631 245296 8647 246072
rect 8681 245296 8693 246072
rect 8631 245284 8693 245296
rect 8749 246072 8811 246084
rect 8749 245296 8761 246072
rect 8795 245296 8811 246072
rect 8749 245284 8811 245296
rect 8841 246072 8903 246084
rect 8841 245296 8857 246072
rect 8891 245296 8903 246072
rect 8841 245284 8903 245296
rect 8959 246072 9021 246084
rect 8959 245296 8971 246072
rect 9005 245296 9021 246072
rect 8959 245284 9021 245296
rect 9051 246072 9113 246084
rect 9051 245296 9067 246072
rect 9101 245296 9113 246072
rect 9051 245284 9113 245296
rect 9169 246072 9231 246084
rect 9169 245296 9181 246072
rect 9215 245296 9231 246072
rect 9169 245284 9231 245296
rect 9261 246072 9323 246084
rect 9261 245296 9277 246072
rect 9311 245296 9323 246072
rect 9261 245284 9323 245296
rect 9379 246072 9441 246084
rect 9379 245296 9391 246072
rect 9425 245296 9441 246072
rect 9379 245284 9441 245296
rect 9471 246072 9533 246084
rect 9471 245296 9487 246072
rect 9521 245296 9533 246072
rect 9471 245284 9533 245296
rect 9589 246072 9651 246084
rect 9589 245296 9601 246072
rect 9635 245296 9651 246072
rect 9589 245284 9651 245296
rect 9681 246072 9743 246084
rect 9681 245296 9697 246072
rect 9731 245296 9743 246072
rect 9681 245284 9743 245296
rect 9799 246072 9861 246084
rect 9799 245296 9811 246072
rect 9845 245296 9861 246072
rect 9799 245284 9861 245296
rect 9891 246072 9953 246084
rect 9891 245296 9907 246072
rect 9941 245296 9953 246072
rect 9891 245284 9953 245296
rect 10009 246072 10071 246084
rect 10009 245296 10021 246072
rect 10055 245296 10071 246072
rect 10009 245284 10071 245296
rect 10101 246072 10163 246084
rect 10101 245296 10117 246072
rect 10151 245296 10163 246072
rect 10101 245284 10163 245296
rect 10219 246072 10281 246084
rect 10219 245296 10231 246072
rect 10265 245296 10281 246072
rect 10219 245284 10281 245296
rect 10311 246072 10373 246084
rect 10311 245296 10327 246072
rect 10361 245296 10373 246072
rect 10311 245284 10373 245296
rect 10429 246072 10491 246084
rect 10429 245296 10441 246072
rect 10475 245296 10491 246072
rect 10429 245284 10491 245296
rect 10521 246072 10583 246084
rect 10521 245296 10537 246072
rect 10571 245296 10583 246072
rect 10521 245284 10583 245296
rect 10639 246072 10701 246084
rect 10639 245296 10651 246072
rect 10685 245296 10701 246072
rect 10639 245284 10701 245296
rect 10731 246072 10793 246084
rect 10731 245296 10747 246072
rect 10781 245296 10793 246072
rect 10731 245284 10793 245296
rect 10849 246072 10911 246084
rect 10849 245296 10861 246072
rect 10895 245296 10911 246072
rect 10849 245284 10911 245296
rect 10941 246072 11003 246084
rect 10941 245296 10957 246072
rect 10991 245296 11003 246072
rect 10941 245284 11003 245296
rect 11059 246072 11121 246084
rect 11059 245296 11071 246072
rect 11105 245296 11121 246072
rect 11059 245284 11121 245296
rect 11151 246072 11213 246084
rect 11151 245296 11167 246072
rect 11201 245296 11213 246072
rect 11151 245284 11213 245296
rect 11269 246072 11331 246084
rect 11269 245296 11281 246072
rect 11315 245296 11331 246072
rect 11269 245284 11331 245296
rect 11361 246072 11423 246084
rect 11361 245296 11377 246072
rect 11411 245296 11423 246072
rect 11361 245284 11423 245296
rect 11479 246072 11541 246084
rect 11479 245296 11491 246072
rect 11525 245296 11541 246072
rect 11479 245284 11541 245296
rect 11571 246072 11633 246084
rect 11571 245296 11587 246072
rect 11621 245296 11633 246072
rect 11571 245284 11633 245296
rect 11689 246072 11751 246084
rect 11689 245296 11701 246072
rect 11735 245296 11751 246072
rect 11689 245284 11751 245296
rect 11781 246072 11843 246084
rect 11781 245296 11797 246072
rect 11831 245296 11843 246072
rect 11781 245284 11843 245296
rect 11899 246072 11961 246084
rect 11899 245296 11911 246072
rect 11945 245296 11961 246072
rect 11899 245284 11961 245296
rect 11991 246072 12053 246084
rect 11991 245296 12007 246072
rect 12041 245296 12053 246072
rect 11991 245284 12053 245296
rect 12109 246072 12171 246084
rect 12109 245296 12121 246072
rect 12155 245296 12171 246072
rect 12109 245284 12171 245296
rect 12201 246072 12263 246084
rect 12201 245296 12217 246072
rect 12251 245296 12263 246072
rect 12201 245284 12263 245296
rect 12319 246072 12381 246084
rect 12319 245296 12331 246072
rect 12365 245296 12381 246072
rect 12319 245284 12381 245296
rect 12411 246072 12473 246084
rect 12411 245296 12427 246072
rect 12461 245296 12473 246072
rect 12411 245284 12473 245296
rect 12529 246072 12591 246084
rect 12529 245296 12541 246072
rect 12575 245296 12591 246072
rect 12529 245284 12591 245296
rect 12621 246072 12683 246084
rect 12621 245296 12637 246072
rect 12671 245296 12683 246072
rect 12621 245284 12683 245296
rect 12739 246072 12801 246084
rect 12739 245296 12751 246072
rect 12785 245296 12801 246072
rect 12739 245284 12801 245296
rect 12831 246072 12893 246084
rect 12831 245296 12847 246072
rect 12881 245296 12893 246072
rect 12831 245284 12893 245296
rect 12949 246072 13011 246084
rect 12949 245296 12961 246072
rect 12995 245296 13011 246072
rect 12949 245284 13011 245296
rect 13041 246072 13103 246084
rect 13041 245296 13057 246072
rect 13091 245296 13103 246072
rect 13041 245284 13103 245296
rect 13159 246072 13221 246084
rect 13159 245296 13171 246072
rect 13205 245296 13221 246072
rect 13159 245284 13221 245296
rect 13251 246072 13313 246084
rect 13251 245296 13267 246072
rect 13301 245296 13313 246072
rect 13251 245284 13313 245296
rect 13369 246072 13431 246084
rect 13369 245296 13381 246072
rect 13415 245296 13431 246072
rect 13369 245284 13431 245296
rect 13461 246072 13523 246084
rect 13461 245296 13477 246072
rect 13511 245296 13523 246072
rect 13461 245284 13523 245296
rect 13579 246072 13641 246084
rect 13579 245296 13591 246072
rect 13625 245296 13641 246072
rect 13579 245284 13641 245296
rect 13671 246072 13733 246084
rect 13671 245296 13687 246072
rect 13721 245296 13733 246072
rect 13671 245284 13733 245296
rect 13789 246072 13851 246084
rect 13789 245296 13801 246072
rect 13835 245296 13851 246072
rect 13789 245284 13851 245296
rect 13881 246072 13943 246084
rect 13881 245296 13897 246072
rect 13931 245296 13943 246072
rect 13881 245284 13943 245296
rect 13999 246072 14061 246084
rect 13999 245296 14011 246072
rect 14045 245296 14061 246072
rect 13999 245284 14061 245296
rect 14091 246072 14153 246084
rect 14091 245296 14107 246072
rect 14141 245296 14153 246072
rect 14091 245284 14153 245296
rect 14209 246072 14271 246084
rect 14209 245296 14221 246072
rect 14255 245296 14271 246072
rect 14209 245284 14271 245296
rect 14301 246072 14363 246084
rect 14301 245296 14317 246072
rect 14351 245296 14363 246072
rect 14301 245284 14363 245296
rect 14419 246072 14481 246084
rect 14419 245296 14431 246072
rect 14465 245296 14481 246072
rect 14419 245284 14481 245296
rect 14511 246072 14573 246084
rect 14511 245296 14527 246072
rect 14561 245296 14573 246072
rect 14511 245284 14573 245296
rect 14629 246072 14691 246084
rect 14629 245296 14641 246072
rect 14675 245296 14691 246072
rect 14629 245284 14691 245296
rect 14721 246072 14783 246084
rect 14721 245296 14737 246072
rect 14771 245296 14783 246072
rect 14721 245284 14783 245296
rect 14839 246072 14901 246084
rect 14839 245296 14851 246072
rect 14885 245296 14901 246072
rect 14839 245284 14901 245296
rect 14931 246072 14993 246084
rect 14931 245296 14947 246072
rect 14981 245296 14993 246072
rect 14931 245284 14993 245296
rect 15049 246072 15111 246084
rect 15049 245296 15061 246072
rect 15095 245296 15111 246072
rect 15049 245284 15111 245296
rect 15141 246072 15203 246084
rect 15141 245296 15157 246072
rect 15191 245296 15203 246072
rect 15141 245284 15203 245296
rect 15259 246072 15321 246084
rect 15259 245296 15271 246072
rect 15305 245296 15321 246072
rect 15259 245284 15321 245296
rect 15351 246072 15413 246084
rect 15351 245296 15367 246072
rect 15401 245296 15413 246072
rect 15351 245284 15413 245296
rect 15469 246072 15531 246084
rect 15469 245296 15481 246072
rect 15515 245296 15531 246072
rect 15469 245284 15531 245296
rect 15561 246072 15623 246084
rect 15561 245296 15577 246072
rect 15611 245296 15623 246072
rect 15561 245284 15623 245296
rect 15679 246072 15741 246084
rect 15679 245296 15691 246072
rect 15725 245296 15741 246072
rect 15679 245284 15741 245296
rect 15771 246072 15833 246084
rect 15771 245296 15787 246072
rect 15821 245296 15833 246072
rect 15771 245284 15833 245296
rect 15889 246072 15951 246084
rect 15889 245296 15901 246072
rect 15935 245296 15951 246072
rect 15889 245284 15951 245296
rect 15981 246072 16043 246084
rect 15981 245296 15997 246072
rect 16031 245296 16043 246072
rect 15981 245284 16043 245296
rect 16099 246072 16161 246084
rect 16099 245296 16111 246072
rect 16145 245296 16161 246072
rect 16099 245284 16161 245296
rect 16191 246072 16253 246084
rect 16191 245296 16207 246072
rect 16241 245296 16253 246072
rect 16191 245284 16253 245296
rect 16309 246072 16371 246084
rect 16309 245296 16321 246072
rect 16355 245296 16371 246072
rect 16309 245284 16371 245296
rect 16401 246072 16463 246084
rect 16401 245296 16417 246072
rect 16451 245296 16463 246072
rect 16401 245284 16463 245296
rect 16519 246072 16581 246084
rect 16519 245296 16531 246072
rect 16565 245296 16581 246072
rect 16519 245284 16581 245296
rect 16611 246072 16673 246084
rect 16611 245296 16627 246072
rect 16661 245296 16673 246072
rect 16611 245284 16673 245296
rect 16729 246072 16791 246084
rect 16729 245296 16741 246072
rect 16775 245296 16791 246072
rect 16729 245284 16791 245296
rect 16821 246072 16883 246084
rect 16821 245296 16837 246072
rect 16871 245296 16883 246072
rect 16821 245284 16883 245296
rect 16939 246072 17001 246084
rect 16939 245296 16951 246072
rect 16985 245296 17001 246072
rect 16939 245284 17001 245296
rect 17031 246072 17093 246084
rect 17031 245296 17047 246072
rect 17081 245296 17093 246072
rect 17031 245284 17093 245296
rect 17149 246072 17211 246084
rect 17149 245296 17161 246072
rect 17195 245296 17211 246072
rect 17149 245284 17211 245296
rect 17241 246072 17303 246084
rect 17241 245296 17257 246072
rect 17291 245296 17303 246072
rect 17241 245284 17303 245296
rect 17359 246072 17421 246084
rect 17359 245296 17371 246072
rect 17405 245296 17421 246072
rect 17359 245284 17421 245296
rect 17451 246072 17513 246084
rect 17451 245296 17467 246072
rect 17501 245296 17513 246072
rect 17451 245284 17513 245296
rect 17569 246072 17631 246084
rect 17569 245296 17581 246072
rect 17615 245296 17631 246072
rect 17569 245284 17631 245296
rect 17661 246072 17723 246084
rect 17661 245296 17677 246072
rect 17711 245296 17723 246072
rect 17661 245284 17723 245296
rect 17779 246072 17841 246084
rect 17779 245296 17791 246072
rect 17825 245296 17841 246072
rect 17779 245284 17841 245296
rect 17871 246072 17933 246084
rect 17871 245296 17887 246072
rect 17921 245296 17933 246072
rect 17871 245284 17933 245296
rect 17989 246072 18051 246084
rect 17989 245296 18001 246072
rect 18035 245296 18051 246072
rect 17989 245284 18051 245296
rect 18081 246072 18143 246084
rect 18081 245296 18097 246072
rect 18131 245296 18143 246072
rect 18081 245284 18143 245296
rect 18199 246072 18261 246084
rect 18199 245296 18211 246072
rect 18245 245296 18261 246072
rect 18199 245284 18261 245296
rect 18291 246072 18353 246084
rect 18291 245296 18307 246072
rect 18341 245296 18353 246072
rect 18291 245284 18353 245296
rect 18409 246072 18471 246084
rect 18409 245296 18421 246072
rect 18455 245296 18471 246072
rect 18409 245284 18471 245296
rect 18501 246072 18563 246084
rect 18501 245296 18517 246072
rect 18551 245296 18563 246072
rect 18501 245284 18563 245296
rect 18619 246072 18681 246084
rect 18619 245296 18631 246072
rect 18665 245296 18681 246072
rect 18619 245284 18681 245296
rect 18711 246072 18773 246084
rect 18711 245296 18727 246072
rect 18761 245296 18773 246072
rect 18711 245284 18773 245296
rect 18829 246072 18891 246084
rect 18829 245296 18841 246072
rect 18875 245296 18891 246072
rect 18829 245284 18891 245296
rect 18921 246072 18983 246084
rect 18921 245296 18937 246072
rect 18971 245296 18983 246072
rect 18921 245284 18983 245296
rect 19039 246072 19101 246084
rect 19039 245296 19051 246072
rect 19085 245296 19101 246072
rect 19039 245284 19101 245296
rect 19131 246072 19193 246084
rect 19131 245296 19147 246072
rect 19181 245296 19193 246072
rect 19131 245284 19193 245296
rect 19249 246072 19311 246084
rect 19249 245296 19261 246072
rect 19295 245296 19311 246072
rect 19249 245284 19311 245296
rect 19341 246072 19403 246084
rect 19341 245296 19357 246072
rect 19391 245296 19403 246072
rect 19341 245284 19403 245296
rect 19459 246072 19521 246084
rect 19459 245296 19471 246072
rect 19505 245296 19521 246072
rect 19459 245284 19521 245296
rect 19551 246072 19613 246084
rect 19551 245296 19567 246072
rect 19601 245296 19613 246072
rect 19551 245284 19613 245296
rect 19669 246072 19731 246084
rect 19669 245296 19681 246072
rect 19715 245296 19731 246072
rect 19669 245284 19731 245296
rect 19761 246072 19823 246084
rect 19761 245296 19777 246072
rect 19811 245296 19823 246072
rect 19761 245284 19823 245296
rect 19879 246072 19941 246084
rect 19879 245296 19891 246072
rect 19925 245296 19941 246072
rect 19879 245284 19941 245296
rect 19971 246072 20033 246084
rect 19971 245296 19987 246072
rect 20021 245296 20033 246072
rect 19971 245284 20033 245296
rect 20089 246072 20151 246084
rect 20089 245296 20101 246072
rect 20135 245296 20151 246072
rect 20089 245284 20151 245296
rect 20181 246072 20243 246084
rect 20181 245296 20197 246072
rect 20231 245296 20243 246072
rect 20181 245284 20243 245296
rect 20299 246072 20361 246084
rect 20299 245296 20311 246072
rect 20345 245296 20361 246072
rect 20299 245284 20361 245296
rect 20391 246072 20453 246084
rect 20391 245296 20407 246072
rect 20441 245296 20453 246072
rect 20391 245284 20453 245296
rect 20509 246072 20571 246084
rect 20509 245296 20521 246072
rect 20555 245296 20571 246072
rect 20509 245284 20571 245296
rect 20601 246072 20663 246084
rect 20601 245296 20617 246072
rect 20651 245296 20663 246072
rect 20601 245284 20663 245296
rect 20719 246072 20781 246084
rect 20719 245296 20731 246072
rect 20765 245296 20781 246072
rect 20719 245284 20781 245296
rect 20811 246072 20873 246084
rect 20811 245296 20827 246072
rect 20861 245296 20873 246072
rect 20811 245284 20873 245296
rect 20929 246072 20991 246084
rect 20929 245296 20941 246072
rect 20975 245296 20991 246072
rect 20929 245284 20991 245296
rect 21021 246072 21083 246084
rect 21021 245296 21037 246072
rect 21071 245296 21083 246072
rect 21021 245284 21083 245296
rect 21139 246072 21201 246084
rect 21139 245296 21151 246072
rect 21185 245296 21201 246072
rect 21139 245284 21201 245296
rect 21231 246072 21293 246084
rect 21231 245296 21247 246072
rect 21281 245296 21293 246072
rect 21231 245284 21293 245296
rect 21349 246072 21411 246084
rect 21349 245296 21361 246072
rect 21395 245296 21411 246072
rect 21349 245284 21411 245296
rect 21441 246072 21503 246084
rect 21441 245296 21457 246072
rect 21491 245296 21503 246072
rect 21441 245284 21503 245296
rect 21559 246072 21621 246084
rect 21559 245296 21571 246072
rect 21605 245296 21621 246072
rect 21559 245284 21621 245296
rect 21651 246072 21713 246084
rect 21651 245296 21667 246072
rect 21701 245296 21713 246072
rect 21651 245284 21713 245296
rect 21769 246072 21831 246084
rect 21769 245296 21781 246072
rect 21815 245296 21831 246072
rect 21769 245284 21831 245296
rect 21861 246072 21923 246084
rect 21861 245296 21877 246072
rect 21911 245296 21923 246072
rect 21861 245284 21923 245296
rect 21979 246072 22041 246084
rect 21979 245296 21991 246072
rect 22025 245296 22041 246072
rect 21979 245284 22041 245296
rect 22071 246072 22133 246084
rect 22071 245296 22087 246072
rect 22121 245296 22133 246072
rect 22071 245284 22133 245296
rect 22189 246072 22251 246084
rect 22189 245296 22201 246072
rect 22235 245296 22251 246072
rect 22189 245284 22251 245296
rect 22281 246072 22343 246084
rect 22281 245296 22297 246072
rect 22331 245296 22343 246072
rect 22281 245284 22343 245296
rect 22399 246072 22461 246084
rect 22399 245296 22411 246072
rect 22445 245296 22461 246072
rect 22399 245284 22461 245296
rect 22491 246072 22553 246084
rect 22491 245296 22507 246072
rect 22541 245296 22553 246072
rect 22491 245284 22553 245296
rect 22609 246072 22671 246084
rect 22609 245296 22621 246072
rect 22655 245296 22671 246072
rect 22609 245284 22671 245296
rect 22701 246072 22763 246084
rect 22701 245296 22717 246072
rect 22751 245296 22763 246072
rect 22701 245284 22763 245296
rect 22819 246072 22881 246084
rect 22819 245296 22831 246072
rect 22865 245296 22881 246072
rect 22819 245284 22881 245296
rect 22911 246072 22973 246084
rect 22911 245296 22927 246072
rect 22961 245296 22973 246072
rect 22911 245284 22973 245296
rect 23029 246072 23091 246084
rect 23029 245296 23041 246072
rect 23075 245296 23091 246072
rect 23029 245284 23091 245296
rect 23121 246072 23183 246084
rect 23121 245296 23137 246072
rect 23171 245296 23183 246072
rect 23121 245284 23183 245296
rect 23239 246072 23301 246084
rect 23239 245296 23251 246072
rect 23285 245296 23301 246072
rect 23239 245284 23301 245296
rect 23331 246072 23393 246084
rect 23331 245296 23347 246072
rect 23381 245296 23393 246072
rect 23331 245284 23393 245296
rect 23449 246072 23511 246084
rect 23449 245296 23461 246072
rect 23495 245296 23511 246072
rect 23449 245284 23511 245296
rect 23541 246072 23603 246084
rect 23541 245296 23557 246072
rect 23591 245296 23603 246072
rect 23541 245284 23603 245296
rect 23659 246072 23721 246084
rect 23659 245296 23671 246072
rect 23705 245296 23721 246072
rect 23659 245284 23721 245296
rect 23751 246072 23813 246084
rect 23751 245296 23767 246072
rect 23801 245296 23813 246072
rect 23751 245284 23813 245296
rect 23869 246072 23931 246084
rect 23869 245296 23881 246072
rect 23915 245296 23931 246072
rect 23869 245284 23931 245296
rect 23961 246072 24023 246084
rect 23961 245296 23977 246072
rect 24011 245296 24023 246072
rect 23961 245284 24023 245296
rect 24079 246072 24141 246084
rect 24079 245296 24091 246072
rect 24125 245296 24141 246072
rect 24079 245284 24141 245296
rect 24171 246072 24233 246084
rect 24171 245296 24187 246072
rect 24221 245296 24233 246072
rect 24171 245284 24233 245296
rect 24289 246072 24351 246084
rect 24289 245296 24301 246072
rect 24335 245296 24351 246072
rect 24289 245284 24351 245296
rect 24381 246072 24443 246084
rect 24381 245296 24397 246072
rect 24431 245296 24443 246072
rect 24381 245284 24443 245296
rect 24499 246072 24561 246084
rect 24499 245296 24511 246072
rect 24545 245296 24561 246072
rect 24499 245284 24561 245296
rect 24591 246072 24653 246084
rect 24591 245296 24607 246072
rect 24641 245296 24653 246072
rect 24591 245284 24653 245296
rect 24709 246072 24771 246084
rect 24709 245296 24721 246072
rect 24755 245296 24771 246072
rect 24709 245284 24771 245296
rect 24801 246072 24863 246084
rect 24801 245296 24817 246072
rect 24851 245296 24863 246072
rect 24801 245284 24863 245296
rect 24919 246072 24981 246084
rect 24919 245296 24931 246072
rect 24965 245296 24981 246072
rect 24919 245284 24981 245296
rect 25011 246072 25073 246084
rect 25011 245296 25027 246072
rect 25061 245296 25073 246072
rect 25011 245284 25073 245296
rect 25129 246072 25191 246084
rect 25129 245296 25141 246072
rect 25175 245296 25191 246072
rect 25129 245284 25191 245296
rect 25221 246072 25283 246084
rect 25221 245296 25237 246072
rect 25271 245296 25283 246072
rect 25221 245284 25283 245296
rect 25339 246072 25401 246084
rect 25339 245296 25351 246072
rect 25385 245296 25401 246072
rect 25339 245284 25401 245296
rect 25431 246072 25493 246084
rect 25431 245296 25447 246072
rect 25481 245296 25493 246072
rect 25431 245284 25493 245296
rect 25549 246072 25611 246084
rect 25549 245296 25561 246072
rect 25595 245296 25611 246072
rect 25549 245284 25611 245296
rect 25641 246072 25703 246084
rect 25641 245296 25657 246072
rect 25691 245296 25703 246072
rect 25641 245284 25703 245296
rect 25759 246072 25821 246084
rect 25759 245296 25771 246072
rect 25805 245296 25821 246072
rect 25759 245284 25821 245296
rect 25851 246072 25913 246084
rect 25851 245296 25867 246072
rect 25901 245296 25913 246072
rect 25851 245284 25913 245296
rect 25969 246072 26031 246084
rect 25969 245296 25981 246072
rect 26015 245296 26031 246072
rect 25969 245284 26031 245296
rect 26061 246072 26123 246084
rect 26061 245296 26077 246072
rect 26111 245296 26123 246072
rect 26061 245284 26123 245296
rect 26179 246072 26241 246084
rect 26179 245296 26191 246072
rect 26225 245296 26241 246072
rect 26179 245284 26241 245296
rect 26271 246072 26333 246084
rect 26271 245296 26287 246072
rect 26321 245296 26333 246072
rect 26271 245284 26333 245296
rect 26389 246072 26451 246084
rect 26389 245296 26401 246072
rect 26435 245296 26451 246072
rect 26389 245284 26451 245296
rect 26481 246072 26543 246084
rect 26481 245296 26497 246072
rect 26531 245296 26543 246072
rect 26481 245284 26543 245296
rect 26599 246072 26661 246084
rect 26599 245296 26611 246072
rect 26645 245296 26661 246072
rect 26599 245284 26661 245296
rect 26691 246072 26753 246084
rect 26691 245296 26707 246072
rect 26741 245296 26753 246072
rect 26691 245284 26753 245296
rect 26809 246072 26871 246084
rect 26809 245296 26821 246072
rect 26855 245296 26871 246072
rect 26809 245284 26871 245296
rect 26901 246072 26963 246084
rect 26901 245296 26917 246072
rect 26951 245296 26963 246072
rect 26901 245284 26963 245296
rect 27019 246072 27081 246084
rect 27019 245296 27031 246072
rect 27065 245296 27081 246072
rect 27019 245284 27081 245296
rect 27111 246072 27173 246084
rect 27111 245296 27127 246072
rect 27161 245296 27173 246072
rect 27111 245284 27173 245296
rect 27229 246072 27291 246084
rect 27229 245296 27241 246072
rect 27275 245296 27291 246072
rect 27229 245284 27291 245296
rect 27321 246072 27383 246084
rect 27321 245296 27337 246072
rect 27371 245296 27383 246072
rect 27321 245284 27383 245296
rect -4061 245036 -3999 245048
rect -4061 244260 -4049 245036
rect -4015 244260 -3999 245036
rect -4061 244248 -3999 244260
rect -3969 245036 -3907 245048
rect -3969 244260 -3953 245036
rect -3919 244260 -3907 245036
rect -3969 244248 -3907 244260
rect -3851 245036 -3789 245048
rect -3851 244260 -3839 245036
rect -3805 244260 -3789 245036
rect -3851 244248 -3789 244260
rect -3759 245036 -3697 245048
rect -3759 244260 -3743 245036
rect -3709 244260 -3697 245036
rect -3759 244248 -3697 244260
rect -3641 245036 -3579 245048
rect -3641 244260 -3629 245036
rect -3595 244260 -3579 245036
rect -3641 244248 -3579 244260
rect -3549 245036 -3487 245048
rect -3549 244260 -3533 245036
rect -3499 244260 -3487 245036
rect -3549 244248 -3487 244260
rect -3431 245036 -3369 245048
rect -3431 244260 -3419 245036
rect -3385 244260 -3369 245036
rect -3431 244248 -3369 244260
rect -3339 245036 -3277 245048
rect -3339 244260 -3323 245036
rect -3289 244260 -3277 245036
rect -3339 244248 -3277 244260
rect -3221 245036 -3159 245048
rect -3221 244260 -3209 245036
rect -3175 244260 -3159 245036
rect -3221 244248 -3159 244260
rect -3129 245036 -3067 245048
rect -3129 244260 -3113 245036
rect -3079 244260 -3067 245036
rect -3129 244248 -3067 244260
rect -3011 245036 -2949 245048
rect -3011 244260 -2999 245036
rect -2965 244260 -2949 245036
rect -3011 244248 -2949 244260
rect -2919 245036 -2857 245048
rect -2919 244260 -2903 245036
rect -2869 244260 -2857 245036
rect -2919 244248 -2857 244260
rect -2801 245036 -2739 245048
rect -2801 244260 -2789 245036
rect -2755 244260 -2739 245036
rect -2801 244248 -2739 244260
rect -2709 245036 -2647 245048
rect -2709 244260 -2693 245036
rect -2659 244260 -2647 245036
rect -2709 244248 -2647 244260
rect -2591 245036 -2529 245048
rect -2591 244260 -2579 245036
rect -2545 244260 -2529 245036
rect -2591 244248 -2529 244260
rect -2499 245036 -2437 245048
rect -2499 244260 -2483 245036
rect -2449 244260 -2437 245036
rect -2499 244248 -2437 244260
rect -2381 245036 -2319 245048
rect -2381 244260 -2369 245036
rect -2335 244260 -2319 245036
rect -2381 244248 -2319 244260
rect -2289 245036 -2227 245048
rect -2289 244260 -2273 245036
rect -2239 244260 -2227 245036
rect -2289 244248 -2227 244260
rect -2171 245036 -2109 245048
rect -2171 244260 -2159 245036
rect -2125 244260 -2109 245036
rect -2171 244248 -2109 244260
rect -2079 245036 -2017 245048
rect -2079 244260 -2063 245036
rect -2029 244260 -2017 245036
rect -2079 244248 -2017 244260
rect -1961 245036 -1899 245048
rect -1961 244260 -1949 245036
rect -1915 244260 -1899 245036
rect -1961 244248 -1899 244260
rect -1869 245036 -1807 245048
rect -1869 244260 -1853 245036
rect -1819 244260 -1807 245036
rect -1869 244248 -1807 244260
rect -1751 245036 -1689 245048
rect -1751 244260 -1739 245036
rect -1705 244260 -1689 245036
rect -1751 244248 -1689 244260
rect -1659 245036 -1597 245048
rect -1659 244260 -1643 245036
rect -1609 244260 -1597 245036
rect -1659 244248 -1597 244260
rect -1541 245036 -1479 245048
rect -1541 244260 -1529 245036
rect -1495 244260 -1479 245036
rect -1541 244248 -1479 244260
rect -1449 245036 -1387 245048
rect -1449 244260 -1433 245036
rect -1399 244260 -1387 245036
rect -1449 244248 -1387 244260
rect -1331 245036 -1269 245048
rect -1331 244260 -1319 245036
rect -1285 244260 -1269 245036
rect -1331 244248 -1269 244260
rect -1239 245036 -1177 245048
rect -1239 244260 -1223 245036
rect -1189 244260 -1177 245036
rect -1239 244248 -1177 244260
rect -1121 245036 -1059 245048
rect -1121 244260 -1109 245036
rect -1075 244260 -1059 245036
rect -1121 244248 -1059 244260
rect -1029 245036 -967 245048
rect -1029 244260 -1013 245036
rect -979 244260 -967 245036
rect -1029 244248 -967 244260
rect -911 245036 -849 245048
rect -911 244260 -899 245036
rect -865 244260 -849 245036
rect -911 244248 -849 244260
rect -819 245036 -757 245048
rect -819 244260 -803 245036
rect -769 244260 -757 245036
rect -819 244248 -757 244260
rect -701 245036 -639 245048
rect -701 244260 -689 245036
rect -655 244260 -639 245036
rect -701 244248 -639 244260
rect -609 245036 -547 245048
rect -609 244260 -593 245036
rect -559 244260 -547 245036
rect -609 244248 -547 244260
rect -491 245036 -429 245048
rect -491 244260 -479 245036
rect -445 244260 -429 245036
rect -491 244248 -429 244260
rect -399 245036 -337 245048
rect -399 244260 -383 245036
rect -349 244260 -337 245036
rect -399 244248 -337 244260
rect -281 245036 -219 245048
rect -281 244260 -269 245036
rect -235 244260 -219 245036
rect -281 244248 -219 244260
rect -189 245036 -127 245048
rect -189 244260 -173 245036
rect -139 244260 -127 245036
rect -189 244248 -127 244260
rect -71 245036 -9 245048
rect -71 244260 -59 245036
rect -25 244260 -9 245036
rect -71 244248 -9 244260
rect 21 245036 83 245048
rect 21 244260 37 245036
rect 71 244260 83 245036
rect 21 244248 83 244260
rect 139 245036 201 245048
rect 139 244260 151 245036
rect 185 244260 201 245036
rect 139 244248 201 244260
rect 231 245036 293 245048
rect 231 244260 247 245036
rect 281 244260 293 245036
rect 231 244248 293 244260
rect 349 245036 411 245048
rect 349 244260 361 245036
rect 395 244260 411 245036
rect 349 244248 411 244260
rect 441 245036 503 245048
rect 441 244260 457 245036
rect 491 244260 503 245036
rect 441 244248 503 244260
rect 559 245036 621 245048
rect 559 244260 571 245036
rect 605 244260 621 245036
rect 559 244248 621 244260
rect 651 245036 713 245048
rect 651 244260 667 245036
rect 701 244260 713 245036
rect 651 244248 713 244260
rect 769 245036 831 245048
rect 769 244260 781 245036
rect 815 244260 831 245036
rect 769 244248 831 244260
rect 861 245036 923 245048
rect 861 244260 877 245036
rect 911 244260 923 245036
rect 861 244248 923 244260
rect 979 245036 1041 245048
rect 979 244260 991 245036
rect 1025 244260 1041 245036
rect 979 244248 1041 244260
rect 1071 245036 1133 245048
rect 1071 244260 1087 245036
rect 1121 244260 1133 245036
rect 1071 244248 1133 244260
rect 1189 245036 1251 245048
rect 1189 244260 1201 245036
rect 1235 244260 1251 245036
rect 1189 244248 1251 244260
rect 1281 245036 1343 245048
rect 1281 244260 1297 245036
rect 1331 244260 1343 245036
rect 1281 244248 1343 244260
rect 1399 245036 1461 245048
rect 1399 244260 1411 245036
rect 1445 244260 1461 245036
rect 1399 244248 1461 244260
rect 1491 245036 1553 245048
rect 1491 244260 1507 245036
rect 1541 244260 1553 245036
rect 1491 244248 1553 244260
rect 1609 245036 1671 245048
rect 1609 244260 1621 245036
rect 1655 244260 1671 245036
rect 1609 244248 1671 244260
rect 1701 245036 1763 245048
rect 1701 244260 1717 245036
rect 1751 244260 1763 245036
rect 1701 244248 1763 244260
rect 1819 245036 1881 245048
rect 1819 244260 1831 245036
rect 1865 244260 1881 245036
rect 1819 244248 1881 244260
rect 1911 245036 1973 245048
rect 1911 244260 1927 245036
rect 1961 244260 1973 245036
rect 1911 244248 1973 244260
rect 2029 245036 2091 245048
rect 2029 244260 2041 245036
rect 2075 244260 2091 245036
rect 2029 244248 2091 244260
rect 2121 245036 2183 245048
rect 2121 244260 2137 245036
rect 2171 244260 2183 245036
rect 2121 244248 2183 244260
rect 2239 245036 2301 245048
rect 2239 244260 2251 245036
rect 2285 244260 2301 245036
rect 2239 244248 2301 244260
rect 2331 245036 2393 245048
rect 2331 244260 2347 245036
rect 2381 244260 2393 245036
rect 2331 244248 2393 244260
rect 2449 245036 2511 245048
rect 2449 244260 2461 245036
rect 2495 244260 2511 245036
rect 2449 244248 2511 244260
rect 2541 245036 2603 245048
rect 2541 244260 2557 245036
rect 2591 244260 2603 245036
rect 2541 244248 2603 244260
rect 2659 245036 2721 245048
rect 2659 244260 2671 245036
rect 2705 244260 2721 245036
rect 2659 244248 2721 244260
rect 2751 245036 2813 245048
rect 2751 244260 2767 245036
rect 2801 244260 2813 245036
rect 2751 244248 2813 244260
rect 2869 245036 2931 245048
rect 2869 244260 2881 245036
rect 2915 244260 2931 245036
rect 2869 244248 2931 244260
rect 2961 245036 3023 245048
rect 2961 244260 2977 245036
rect 3011 244260 3023 245036
rect 2961 244248 3023 244260
rect 3079 245036 3141 245048
rect 3079 244260 3091 245036
rect 3125 244260 3141 245036
rect 3079 244248 3141 244260
rect 3171 245036 3233 245048
rect 3171 244260 3187 245036
rect 3221 244260 3233 245036
rect 3171 244248 3233 244260
rect 3289 245036 3351 245048
rect 3289 244260 3301 245036
rect 3335 244260 3351 245036
rect 3289 244248 3351 244260
rect 3381 245036 3443 245048
rect 3381 244260 3397 245036
rect 3431 244260 3443 245036
rect 3381 244248 3443 244260
rect 3499 245036 3561 245048
rect 3499 244260 3511 245036
rect 3545 244260 3561 245036
rect 3499 244248 3561 244260
rect 3591 245036 3653 245048
rect 3591 244260 3607 245036
rect 3641 244260 3653 245036
rect 3591 244248 3653 244260
rect 3709 245036 3771 245048
rect 3709 244260 3721 245036
rect 3755 244260 3771 245036
rect 3709 244248 3771 244260
rect 3801 245036 3863 245048
rect 3801 244260 3817 245036
rect 3851 244260 3863 245036
rect 3801 244248 3863 244260
rect 3919 245036 3981 245048
rect 3919 244260 3931 245036
rect 3965 244260 3981 245036
rect 3919 244248 3981 244260
rect 4011 245036 4073 245048
rect 4011 244260 4027 245036
rect 4061 244260 4073 245036
rect 4011 244248 4073 244260
rect 4129 245036 4191 245048
rect 4129 244260 4141 245036
rect 4175 244260 4191 245036
rect 4129 244248 4191 244260
rect 4221 245036 4283 245048
rect 4221 244260 4237 245036
rect 4271 244260 4283 245036
rect 4221 244248 4283 244260
rect 4339 245036 4401 245048
rect 4339 244260 4351 245036
rect 4385 244260 4401 245036
rect 4339 244248 4401 244260
rect 4431 245036 4493 245048
rect 4431 244260 4447 245036
rect 4481 244260 4493 245036
rect 4431 244248 4493 244260
rect 4549 245036 4611 245048
rect 4549 244260 4561 245036
rect 4595 244260 4611 245036
rect 4549 244248 4611 244260
rect 4641 245036 4703 245048
rect 4641 244260 4657 245036
rect 4691 244260 4703 245036
rect 4641 244248 4703 244260
rect 4759 245036 4821 245048
rect 4759 244260 4771 245036
rect 4805 244260 4821 245036
rect 4759 244248 4821 244260
rect 4851 245036 4913 245048
rect 4851 244260 4867 245036
rect 4901 244260 4913 245036
rect 4851 244248 4913 244260
rect 4969 245036 5031 245048
rect 4969 244260 4981 245036
rect 5015 244260 5031 245036
rect 4969 244248 5031 244260
rect 5061 245036 5123 245048
rect 5061 244260 5077 245036
rect 5111 244260 5123 245036
rect 5061 244248 5123 244260
rect 5179 245036 5241 245048
rect 5179 244260 5191 245036
rect 5225 244260 5241 245036
rect 5179 244248 5241 244260
rect 5271 245036 5333 245048
rect 5271 244260 5287 245036
rect 5321 244260 5333 245036
rect 5271 244248 5333 244260
rect 5389 245036 5451 245048
rect 5389 244260 5401 245036
rect 5435 244260 5451 245036
rect 5389 244248 5451 244260
rect 5481 245036 5543 245048
rect 5481 244260 5497 245036
rect 5531 244260 5543 245036
rect 5481 244248 5543 244260
rect 5599 245036 5661 245048
rect 5599 244260 5611 245036
rect 5645 244260 5661 245036
rect 5599 244248 5661 244260
rect 5691 245036 5753 245048
rect 5691 244260 5707 245036
rect 5741 244260 5753 245036
rect 5691 244248 5753 244260
rect 5809 245036 5871 245048
rect 5809 244260 5821 245036
rect 5855 244260 5871 245036
rect 5809 244248 5871 244260
rect 5901 245036 5963 245048
rect 5901 244260 5917 245036
rect 5951 244260 5963 245036
rect 5901 244248 5963 244260
rect 6019 245036 6081 245048
rect 6019 244260 6031 245036
rect 6065 244260 6081 245036
rect 6019 244248 6081 244260
rect 6111 245036 6173 245048
rect 6111 244260 6127 245036
rect 6161 244260 6173 245036
rect 6111 244248 6173 244260
rect 6229 245036 6291 245048
rect 6229 244260 6241 245036
rect 6275 244260 6291 245036
rect 6229 244248 6291 244260
rect 6321 245036 6383 245048
rect 6321 244260 6337 245036
rect 6371 244260 6383 245036
rect 6321 244248 6383 244260
rect 6439 245036 6501 245048
rect 6439 244260 6451 245036
rect 6485 244260 6501 245036
rect 6439 244248 6501 244260
rect 6531 245036 6593 245048
rect 6531 244260 6547 245036
rect 6581 244260 6593 245036
rect 6531 244248 6593 244260
rect 6649 245036 6711 245048
rect 6649 244260 6661 245036
rect 6695 244260 6711 245036
rect 6649 244248 6711 244260
rect 6741 245036 6803 245048
rect 6741 244260 6757 245036
rect 6791 244260 6803 245036
rect 6741 244248 6803 244260
rect 6859 245036 6921 245048
rect 6859 244260 6871 245036
rect 6905 244260 6921 245036
rect 6859 244248 6921 244260
rect 6951 245036 7013 245048
rect 6951 244260 6967 245036
rect 7001 244260 7013 245036
rect 6951 244248 7013 244260
rect 7069 245036 7131 245048
rect 7069 244260 7081 245036
rect 7115 244260 7131 245036
rect 7069 244248 7131 244260
rect 7161 245036 7223 245048
rect 7161 244260 7177 245036
rect 7211 244260 7223 245036
rect 7161 244248 7223 244260
rect 7279 245036 7341 245048
rect 7279 244260 7291 245036
rect 7325 244260 7341 245036
rect 7279 244248 7341 244260
rect 7371 245036 7433 245048
rect 7371 244260 7387 245036
rect 7421 244260 7433 245036
rect 7371 244248 7433 244260
rect 7489 245036 7551 245048
rect 7489 244260 7501 245036
rect 7535 244260 7551 245036
rect 7489 244248 7551 244260
rect 7581 245036 7643 245048
rect 7581 244260 7597 245036
rect 7631 244260 7643 245036
rect 7581 244248 7643 244260
rect 7699 245036 7761 245048
rect 7699 244260 7711 245036
rect 7745 244260 7761 245036
rect 7699 244248 7761 244260
rect 7791 245036 7853 245048
rect 7791 244260 7807 245036
rect 7841 244260 7853 245036
rect 7791 244248 7853 244260
rect 7909 245036 7971 245048
rect 7909 244260 7921 245036
rect 7955 244260 7971 245036
rect 7909 244248 7971 244260
rect 8001 245036 8063 245048
rect 8001 244260 8017 245036
rect 8051 244260 8063 245036
rect 8001 244248 8063 244260
rect 8119 245036 8181 245048
rect 8119 244260 8131 245036
rect 8165 244260 8181 245036
rect 8119 244248 8181 244260
rect 8211 245036 8273 245048
rect 8211 244260 8227 245036
rect 8261 244260 8273 245036
rect 8211 244248 8273 244260
rect 8329 245036 8391 245048
rect 8329 244260 8341 245036
rect 8375 244260 8391 245036
rect 8329 244248 8391 244260
rect 8421 245036 8483 245048
rect 8421 244260 8437 245036
rect 8471 244260 8483 245036
rect 8421 244248 8483 244260
rect 8539 245036 8601 245048
rect 8539 244260 8551 245036
rect 8585 244260 8601 245036
rect 8539 244248 8601 244260
rect 8631 245036 8693 245048
rect 8631 244260 8647 245036
rect 8681 244260 8693 245036
rect 8631 244248 8693 244260
rect 8749 245036 8811 245048
rect 8749 244260 8761 245036
rect 8795 244260 8811 245036
rect 8749 244248 8811 244260
rect 8841 245036 8903 245048
rect 8841 244260 8857 245036
rect 8891 244260 8903 245036
rect 8841 244248 8903 244260
rect 8959 245036 9021 245048
rect 8959 244260 8971 245036
rect 9005 244260 9021 245036
rect 8959 244248 9021 244260
rect 9051 245036 9113 245048
rect 9051 244260 9067 245036
rect 9101 244260 9113 245036
rect 9051 244248 9113 244260
rect 9169 245036 9231 245048
rect 9169 244260 9181 245036
rect 9215 244260 9231 245036
rect 9169 244248 9231 244260
rect 9261 245036 9323 245048
rect 9261 244260 9277 245036
rect 9311 244260 9323 245036
rect 9261 244248 9323 244260
rect 9379 245036 9441 245048
rect 9379 244260 9391 245036
rect 9425 244260 9441 245036
rect 9379 244248 9441 244260
rect 9471 245036 9533 245048
rect 9471 244260 9487 245036
rect 9521 244260 9533 245036
rect 9471 244248 9533 244260
rect 9589 245036 9651 245048
rect 9589 244260 9601 245036
rect 9635 244260 9651 245036
rect 9589 244248 9651 244260
rect 9681 245036 9743 245048
rect 9681 244260 9697 245036
rect 9731 244260 9743 245036
rect 9681 244248 9743 244260
rect 9799 245036 9861 245048
rect 9799 244260 9811 245036
rect 9845 244260 9861 245036
rect 9799 244248 9861 244260
rect 9891 245036 9953 245048
rect 9891 244260 9907 245036
rect 9941 244260 9953 245036
rect 9891 244248 9953 244260
rect 10009 245036 10071 245048
rect 10009 244260 10021 245036
rect 10055 244260 10071 245036
rect 10009 244248 10071 244260
rect 10101 245036 10163 245048
rect 10101 244260 10117 245036
rect 10151 244260 10163 245036
rect 10101 244248 10163 244260
rect 10219 245036 10281 245048
rect 10219 244260 10231 245036
rect 10265 244260 10281 245036
rect 10219 244248 10281 244260
rect 10311 245036 10373 245048
rect 10311 244260 10327 245036
rect 10361 244260 10373 245036
rect 10311 244248 10373 244260
rect 10429 245036 10491 245048
rect 10429 244260 10441 245036
rect 10475 244260 10491 245036
rect 10429 244248 10491 244260
rect 10521 245036 10583 245048
rect 10521 244260 10537 245036
rect 10571 244260 10583 245036
rect 10521 244248 10583 244260
rect 10639 245036 10701 245048
rect 10639 244260 10651 245036
rect 10685 244260 10701 245036
rect 10639 244248 10701 244260
rect 10731 245036 10793 245048
rect 10731 244260 10747 245036
rect 10781 244260 10793 245036
rect 10731 244248 10793 244260
rect 10849 245036 10911 245048
rect 10849 244260 10861 245036
rect 10895 244260 10911 245036
rect 10849 244248 10911 244260
rect 10941 245036 11003 245048
rect 10941 244260 10957 245036
rect 10991 244260 11003 245036
rect 10941 244248 11003 244260
rect 11059 245036 11121 245048
rect 11059 244260 11071 245036
rect 11105 244260 11121 245036
rect 11059 244248 11121 244260
rect 11151 245036 11213 245048
rect 11151 244260 11167 245036
rect 11201 244260 11213 245036
rect 11151 244248 11213 244260
rect 11269 245036 11331 245048
rect 11269 244260 11281 245036
rect 11315 244260 11331 245036
rect 11269 244248 11331 244260
rect 11361 245036 11423 245048
rect 11361 244260 11377 245036
rect 11411 244260 11423 245036
rect 11361 244248 11423 244260
rect 11479 245036 11541 245048
rect 11479 244260 11491 245036
rect 11525 244260 11541 245036
rect 11479 244248 11541 244260
rect 11571 245036 11633 245048
rect 11571 244260 11587 245036
rect 11621 244260 11633 245036
rect 11571 244248 11633 244260
rect 11689 245036 11751 245048
rect 11689 244260 11701 245036
rect 11735 244260 11751 245036
rect 11689 244248 11751 244260
rect 11781 245036 11843 245048
rect 11781 244260 11797 245036
rect 11831 244260 11843 245036
rect 11781 244248 11843 244260
rect 11899 245036 11961 245048
rect 11899 244260 11911 245036
rect 11945 244260 11961 245036
rect 11899 244248 11961 244260
rect 11991 245036 12053 245048
rect 11991 244260 12007 245036
rect 12041 244260 12053 245036
rect 11991 244248 12053 244260
rect 12109 245036 12171 245048
rect 12109 244260 12121 245036
rect 12155 244260 12171 245036
rect 12109 244248 12171 244260
rect 12201 245036 12263 245048
rect 12201 244260 12217 245036
rect 12251 244260 12263 245036
rect 12201 244248 12263 244260
rect 12319 245036 12381 245048
rect 12319 244260 12331 245036
rect 12365 244260 12381 245036
rect 12319 244248 12381 244260
rect 12411 245036 12473 245048
rect 12411 244260 12427 245036
rect 12461 244260 12473 245036
rect 12411 244248 12473 244260
rect 12529 245036 12591 245048
rect 12529 244260 12541 245036
rect 12575 244260 12591 245036
rect 12529 244248 12591 244260
rect 12621 245036 12683 245048
rect 12621 244260 12637 245036
rect 12671 244260 12683 245036
rect 12621 244248 12683 244260
rect 12739 245036 12801 245048
rect 12739 244260 12751 245036
rect 12785 244260 12801 245036
rect 12739 244248 12801 244260
rect 12831 245036 12893 245048
rect 12831 244260 12847 245036
rect 12881 244260 12893 245036
rect 12831 244248 12893 244260
rect 12949 245036 13011 245048
rect 12949 244260 12961 245036
rect 12995 244260 13011 245036
rect 12949 244248 13011 244260
rect 13041 245036 13103 245048
rect 13041 244260 13057 245036
rect 13091 244260 13103 245036
rect 13041 244248 13103 244260
rect 13159 245036 13221 245048
rect 13159 244260 13171 245036
rect 13205 244260 13221 245036
rect 13159 244248 13221 244260
rect 13251 245036 13313 245048
rect 13251 244260 13267 245036
rect 13301 244260 13313 245036
rect 13251 244248 13313 244260
rect 13369 245036 13431 245048
rect 13369 244260 13381 245036
rect 13415 244260 13431 245036
rect 13369 244248 13431 244260
rect 13461 245036 13523 245048
rect 13461 244260 13477 245036
rect 13511 244260 13523 245036
rect 13461 244248 13523 244260
rect 13579 245036 13641 245048
rect 13579 244260 13591 245036
rect 13625 244260 13641 245036
rect 13579 244248 13641 244260
rect 13671 245036 13733 245048
rect 13671 244260 13687 245036
rect 13721 244260 13733 245036
rect 13671 244248 13733 244260
rect 13789 245036 13851 245048
rect 13789 244260 13801 245036
rect 13835 244260 13851 245036
rect 13789 244248 13851 244260
rect 13881 245036 13943 245048
rect 13881 244260 13897 245036
rect 13931 244260 13943 245036
rect 13881 244248 13943 244260
rect 13999 245036 14061 245048
rect 13999 244260 14011 245036
rect 14045 244260 14061 245036
rect 13999 244248 14061 244260
rect 14091 245036 14153 245048
rect 14091 244260 14107 245036
rect 14141 244260 14153 245036
rect 14091 244248 14153 244260
rect 14209 245036 14271 245048
rect 14209 244260 14221 245036
rect 14255 244260 14271 245036
rect 14209 244248 14271 244260
rect 14301 245036 14363 245048
rect 14301 244260 14317 245036
rect 14351 244260 14363 245036
rect 14301 244248 14363 244260
rect 14419 245036 14481 245048
rect 14419 244260 14431 245036
rect 14465 244260 14481 245036
rect 14419 244248 14481 244260
rect 14511 245036 14573 245048
rect 14511 244260 14527 245036
rect 14561 244260 14573 245036
rect 14511 244248 14573 244260
rect 14629 245036 14691 245048
rect 14629 244260 14641 245036
rect 14675 244260 14691 245036
rect 14629 244248 14691 244260
rect 14721 245036 14783 245048
rect 14721 244260 14737 245036
rect 14771 244260 14783 245036
rect 14721 244248 14783 244260
rect 14839 245036 14901 245048
rect 14839 244260 14851 245036
rect 14885 244260 14901 245036
rect 14839 244248 14901 244260
rect 14931 245036 14993 245048
rect 14931 244260 14947 245036
rect 14981 244260 14993 245036
rect 14931 244248 14993 244260
rect 15049 245036 15111 245048
rect 15049 244260 15061 245036
rect 15095 244260 15111 245036
rect 15049 244248 15111 244260
rect 15141 245036 15203 245048
rect 15141 244260 15157 245036
rect 15191 244260 15203 245036
rect 15141 244248 15203 244260
rect 15259 245036 15321 245048
rect 15259 244260 15271 245036
rect 15305 244260 15321 245036
rect 15259 244248 15321 244260
rect 15351 245036 15413 245048
rect 15351 244260 15367 245036
rect 15401 244260 15413 245036
rect 15351 244248 15413 244260
rect 15469 245036 15531 245048
rect 15469 244260 15481 245036
rect 15515 244260 15531 245036
rect 15469 244248 15531 244260
rect 15561 245036 15623 245048
rect 15561 244260 15577 245036
rect 15611 244260 15623 245036
rect 15561 244248 15623 244260
rect 15679 245036 15741 245048
rect 15679 244260 15691 245036
rect 15725 244260 15741 245036
rect 15679 244248 15741 244260
rect 15771 245036 15833 245048
rect 15771 244260 15787 245036
rect 15821 244260 15833 245036
rect 15771 244248 15833 244260
rect 15889 245036 15951 245048
rect 15889 244260 15901 245036
rect 15935 244260 15951 245036
rect 15889 244248 15951 244260
rect 15981 245036 16043 245048
rect 15981 244260 15997 245036
rect 16031 244260 16043 245036
rect 15981 244248 16043 244260
rect 16099 245036 16161 245048
rect 16099 244260 16111 245036
rect 16145 244260 16161 245036
rect 16099 244248 16161 244260
rect 16191 245036 16253 245048
rect 16191 244260 16207 245036
rect 16241 244260 16253 245036
rect 16191 244248 16253 244260
rect 16309 245036 16371 245048
rect 16309 244260 16321 245036
rect 16355 244260 16371 245036
rect 16309 244248 16371 244260
rect 16401 245036 16463 245048
rect 16401 244260 16417 245036
rect 16451 244260 16463 245036
rect 16401 244248 16463 244260
rect 16519 245036 16581 245048
rect 16519 244260 16531 245036
rect 16565 244260 16581 245036
rect 16519 244248 16581 244260
rect 16611 245036 16673 245048
rect 16611 244260 16627 245036
rect 16661 244260 16673 245036
rect 16611 244248 16673 244260
rect 16729 245036 16791 245048
rect 16729 244260 16741 245036
rect 16775 244260 16791 245036
rect 16729 244248 16791 244260
rect 16821 245036 16883 245048
rect 16821 244260 16837 245036
rect 16871 244260 16883 245036
rect 16821 244248 16883 244260
rect 16939 245036 17001 245048
rect 16939 244260 16951 245036
rect 16985 244260 17001 245036
rect 16939 244248 17001 244260
rect 17031 245036 17093 245048
rect 17031 244260 17047 245036
rect 17081 244260 17093 245036
rect 17031 244248 17093 244260
rect 17149 245036 17211 245048
rect 17149 244260 17161 245036
rect 17195 244260 17211 245036
rect 17149 244248 17211 244260
rect 17241 245036 17303 245048
rect 17241 244260 17257 245036
rect 17291 244260 17303 245036
rect 17241 244248 17303 244260
rect 17359 245036 17421 245048
rect 17359 244260 17371 245036
rect 17405 244260 17421 245036
rect 17359 244248 17421 244260
rect 17451 245036 17513 245048
rect 17451 244260 17467 245036
rect 17501 244260 17513 245036
rect 17451 244248 17513 244260
rect 17569 245036 17631 245048
rect 17569 244260 17581 245036
rect 17615 244260 17631 245036
rect 17569 244248 17631 244260
rect 17661 245036 17723 245048
rect 17661 244260 17677 245036
rect 17711 244260 17723 245036
rect 17661 244248 17723 244260
rect 17779 245036 17841 245048
rect 17779 244260 17791 245036
rect 17825 244260 17841 245036
rect 17779 244248 17841 244260
rect 17871 245036 17933 245048
rect 17871 244260 17887 245036
rect 17921 244260 17933 245036
rect 17871 244248 17933 244260
rect 17989 245036 18051 245048
rect 17989 244260 18001 245036
rect 18035 244260 18051 245036
rect 17989 244248 18051 244260
rect 18081 245036 18143 245048
rect 18081 244260 18097 245036
rect 18131 244260 18143 245036
rect 18081 244248 18143 244260
rect 18199 245036 18261 245048
rect 18199 244260 18211 245036
rect 18245 244260 18261 245036
rect 18199 244248 18261 244260
rect 18291 245036 18353 245048
rect 18291 244260 18307 245036
rect 18341 244260 18353 245036
rect 18291 244248 18353 244260
rect 18409 245036 18471 245048
rect 18409 244260 18421 245036
rect 18455 244260 18471 245036
rect 18409 244248 18471 244260
rect 18501 245036 18563 245048
rect 18501 244260 18517 245036
rect 18551 244260 18563 245036
rect 18501 244248 18563 244260
rect 18619 245036 18681 245048
rect 18619 244260 18631 245036
rect 18665 244260 18681 245036
rect 18619 244248 18681 244260
rect 18711 245036 18773 245048
rect 18711 244260 18727 245036
rect 18761 244260 18773 245036
rect 18711 244248 18773 244260
rect 18829 245036 18891 245048
rect 18829 244260 18841 245036
rect 18875 244260 18891 245036
rect 18829 244248 18891 244260
rect 18921 245036 18983 245048
rect 18921 244260 18937 245036
rect 18971 244260 18983 245036
rect 18921 244248 18983 244260
rect 19039 245036 19101 245048
rect 19039 244260 19051 245036
rect 19085 244260 19101 245036
rect 19039 244248 19101 244260
rect 19131 245036 19193 245048
rect 19131 244260 19147 245036
rect 19181 244260 19193 245036
rect 19131 244248 19193 244260
rect 19249 245036 19311 245048
rect 19249 244260 19261 245036
rect 19295 244260 19311 245036
rect 19249 244248 19311 244260
rect 19341 245036 19403 245048
rect 19341 244260 19357 245036
rect 19391 244260 19403 245036
rect 19341 244248 19403 244260
rect 19459 245036 19521 245048
rect 19459 244260 19471 245036
rect 19505 244260 19521 245036
rect 19459 244248 19521 244260
rect 19551 245036 19613 245048
rect 19551 244260 19567 245036
rect 19601 244260 19613 245036
rect 19551 244248 19613 244260
rect 19669 245036 19731 245048
rect 19669 244260 19681 245036
rect 19715 244260 19731 245036
rect 19669 244248 19731 244260
rect 19761 245036 19823 245048
rect 19761 244260 19777 245036
rect 19811 244260 19823 245036
rect 19761 244248 19823 244260
rect 19879 245036 19941 245048
rect 19879 244260 19891 245036
rect 19925 244260 19941 245036
rect 19879 244248 19941 244260
rect 19971 245036 20033 245048
rect 19971 244260 19987 245036
rect 20021 244260 20033 245036
rect 19971 244248 20033 244260
rect 20089 245036 20151 245048
rect 20089 244260 20101 245036
rect 20135 244260 20151 245036
rect 20089 244248 20151 244260
rect 20181 245036 20243 245048
rect 20181 244260 20197 245036
rect 20231 244260 20243 245036
rect 20181 244248 20243 244260
rect 20299 245036 20361 245048
rect 20299 244260 20311 245036
rect 20345 244260 20361 245036
rect 20299 244248 20361 244260
rect 20391 245036 20453 245048
rect 20391 244260 20407 245036
rect 20441 244260 20453 245036
rect 20391 244248 20453 244260
rect 20509 245036 20571 245048
rect 20509 244260 20521 245036
rect 20555 244260 20571 245036
rect 20509 244248 20571 244260
rect 20601 245036 20663 245048
rect 20601 244260 20617 245036
rect 20651 244260 20663 245036
rect 20601 244248 20663 244260
rect 20719 245036 20781 245048
rect 20719 244260 20731 245036
rect 20765 244260 20781 245036
rect 20719 244248 20781 244260
rect 20811 245036 20873 245048
rect 20811 244260 20827 245036
rect 20861 244260 20873 245036
rect 20811 244248 20873 244260
rect 20929 245036 20991 245048
rect 20929 244260 20941 245036
rect 20975 244260 20991 245036
rect 20929 244248 20991 244260
rect 21021 245036 21083 245048
rect 21021 244260 21037 245036
rect 21071 244260 21083 245036
rect 21021 244248 21083 244260
rect 21139 245036 21201 245048
rect 21139 244260 21151 245036
rect 21185 244260 21201 245036
rect 21139 244248 21201 244260
rect 21231 245036 21293 245048
rect 21231 244260 21247 245036
rect 21281 244260 21293 245036
rect 21231 244248 21293 244260
rect 21349 245036 21411 245048
rect 21349 244260 21361 245036
rect 21395 244260 21411 245036
rect 21349 244248 21411 244260
rect 21441 245036 21503 245048
rect 21441 244260 21457 245036
rect 21491 244260 21503 245036
rect 21441 244248 21503 244260
rect 21559 245036 21621 245048
rect 21559 244260 21571 245036
rect 21605 244260 21621 245036
rect 21559 244248 21621 244260
rect 21651 245036 21713 245048
rect 21651 244260 21667 245036
rect 21701 244260 21713 245036
rect 21651 244248 21713 244260
rect 21769 245036 21831 245048
rect 21769 244260 21781 245036
rect 21815 244260 21831 245036
rect 21769 244248 21831 244260
rect 21861 245036 21923 245048
rect 21861 244260 21877 245036
rect 21911 244260 21923 245036
rect 21861 244248 21923 244260
rect 21979 245036 22041 245048
rect 21979 244260 21991 245036
rect 22025 244260 22041 245036
rect 21979 244248 22041 244260
rect 22071 245036 22133 245048
rect 22071 244260 22087 245036
rect 22121 244260 22133 245036
rect 22071 244248 22133 244260
rect 22189 245036 22251 245048
rect 22189 244260 22201 245036
rect 22235 244260 22251 245036
rect 22189 244248 22251 244260
rect 22281 245036 22343 245048
rect 22281 244260 22297 245036
rect 22331 244260 22343 245036
rect 22281 244248 22343 244260
rect 22399 245036 22461 245048
rect 22399 244260 22411 245036
rect 22445 244260 22461 245036
rect 22399 244248 22461 244260
rect 22491 245036 22553 245048
rect 22491 244260 22507 245036
rect 22541 244260 22553 245036
rect 22491 244248 22553 244260
rect 22609 245036 22671 245048
rect 22609 244260 22621 245036
rect 22655 244260 22671 245036
rect 22609 244248 22671 244260
rect 22701 245036 22763 245048
rect 22701 244260 22717 245036
rect 22751 244260 22763 245036
rect 22701 244248 22763 244260
rect 22819 245036 22881 245048
rect 22819 244260 22831 245036
rect 22865 244260 22881 245036
rect 22819 244248 22881 244260
rect 22911 245036 22973 245048
rect 22911 244260 22927 245036
rect 22961 244260 22973 245036
rect 22911 244248 22973 244260
rect 23029 245036 23091 245048
rect 23029 244260 23041 245036
rect 23075 244260 23091 245036
rect 23029 244248 23091 244260
rect 23121 245036 23183 245048
rect 23121 244260 23137 245036
rect 23171 244260 23183 245036
rect 23121 244248 23183 244260
rect 23239 245036 23301 245048
rect 23239 244260 23251 245036
rect 23285 244260 23301 245036
rect 23239 244248 23301 244260
rect 23331 245036 23393 245048
rect 23331 244260 23347 245036
rect 23381 244260 23393 245036
rect 23331 244248 23393 244260
rect 23449 245036 23511 245048
rect 23449 244260 23461 245036
rect 23495 244260 23511 245036
rect 23449 244248 23511 244260
rect 23541 245036 23603 245048
rect 23541 244260 23557 245036
rect 23591 244260 23603 245036
rect 23541 244248 23603 244260
rect 23659 245036 23721 245048
rect 23659 244260 23671 245036
rect 23705 244260 23721 245036
rect 23659 244248 23721 244260
rect 23751 245036 23813 245048
rect 23751 244260 23767 245036
rect 23801 244260 23813 245036
rect 23751 244248 23813 244260
rect 23869 245036 23931 245048
rect 23869 244260 23881 245036
rect 23915 244260 23931 245036
rect 23869 244248 23931 244260
rect 23961 245036 24023 245048
rect 23961 244260 23977 245036
rect 24011 244260 24023 245036
rect 23961 244248 24023 244260
rect 24079 245036 24141 245048
rect 24079 244260 24091 245036
rect 24125 244260 24141 245036
rect 24079 244248 24141 244260
rect 24171 245036 24233 245048
rect 24171 244260 24187 245036
rect 24221 244260 24233 245036
rect 24171 244248 24233 244260
rect 24289 245036 24351 245048
rect 24289 244260 24301 245036
rect 24335 244260 24351 245036
rect 24289 244248 24351 244260
rect 24381 245036 24443 245048
rect 24381 244260 24397 245036
rect 24431 244260 24443 245036
rect 24381 244248 24443 244260
rect 24499 245036 24561 245048
rect 24499 244260 24511 245036
rect 24545 244260 24561 245036
rect 24499 244248 24561 244260
rect 24591 245036 24653 245048
rect 24591 244260 24607 245036
rect 24641 244260 24653 245036
rect 24591 244248 24653 244260
rect 24709 245036 24771 245048
rect 24709 244260 24721 245036
rect 24755 244260 24771 245036
rect 24709 244248 24771 244260
rect 24801 245036 24863 245048
rect 24801 244260 24817 245036
rect 24851 244260 24863 245036
rect 24801 244248 24863 244260
rect 24919 245036 24981 245048
rect 24919 244260 24931 245036
rect 24965 244260 24981 245036
rect 24919 244248 24981 244260
rect 25011 245036 25073 245048
rect 25011 244260 25027 245036
rect 25061 244260 25073 245036
rect 25011 244248 25073 244260
rect 25129 245036 25191 245048
rect 25129 244260 25141 245036
rect 25175 244260 25191 245036
rect 25129 244248 25191 244260
rect 25221 245036 25283 245048
rect 25221 244260 25237 245036
rect 25271 244260 25283 245036
rect 25221 244248 25283 244260
rect 25339 245036 25401 245048
rect 25339 244260 25351 245036
rect 25385 244260 25401 245036
rect 25339 244248 25401 244260
rect 25431 245036 25493 245048
rect 25431 244260 25447 245036
rect 25481 244260 25493 245036
rect 25431 244248 25493 244260
rect 25549 245036 25611 245048
rect 25549 244260 25561 245036
rect 25595 244260 25611 245036
rect 25549 244248 25611 244260
rect 25641 245036 25703 245048
rect 25641 244260 25657 245036
rect 25691 244260 25703 245036
rect 25641 244248 25703 244260
rect 25759 245036 25821 245048
rect 25759 244260 25771 245036
rect 25805 244260 25821 245036
rect 25759 244248 25821 244260
rect 25851 245036 25913 245048
rect 25851 244260 25867 245036
rect 25901 244260 25913 245036
rect 25851 244248 25913 244260
rect 25969 245036 26031 245048
rect 25969 244260 25981 245036
rect 26015 244260 26031 245036
rect 25969 244248 26031 244260
rect 26061 245036 26123 245048
rect 26061 244260 26077 245036
rect 26111 244260 26123 245036
rect 26061 244248 26123 244260
rect 26179 245036 26241 245048
rect 26179 244260 26191 245036
rect 26225 244260 26241 245036
rect 26179 244248 26241 244260
rect 26271 245036 26333 245048
rect 26271 244260 26287 245036
rect 26321 244260 26333 245036
rect 26271 244248 26333 244260
rect 26389 245036 26451 245048
rect 26389 244260 26401 245036
rect 26435 244260 26451 245036
rect 26389 244248 26451 244260
rect 26481 245036 26543 245048
rect 26481 244260 26497 245036
rect 26531 244260 26543 245036
rect 26481 244248 26543 244260
rect 26599 245036 26661 245048
rect 26599 244260 26611 245036
rect 26645 244260 26661 245036
rect 26599 244248 26661 244260
rect 26691 245036 26753 245048
rect 26691 244260 26707 245036
rect 26741 244260 26753 245036
rect 26691 244248 26753 244260
rect 26809 245036 26871 245048
rect 26809 244260 26821 245036
rect 26855 244260 26871 245036
rect 26809 244248 26871 244260
rect 26901 245036 26963 245048
rect 26901 244260 26917 245036
rect 26951 244260 26963 245036
rect 26901 244248 26963 244260
rect 27019 245036 27081 245048
rect 27019 244260 27031 245036
rect 27065 244260 27081 245036
rect 27019 244248 27081 244260
rect 27111 245036 27173 245048
rect 27111 244260 27127 245036
rect 27161 244260 27173 245036
rect 27111 244248 27173 244260
rect 27229 245036 27291 245048
rect 27229 244260 27241 245036
rect 27275 244260 27291 245036
rect 27229 244248 27291 244260
rect 27321 245036 27383 245048
rect 27321 244260 27337 245036
rect 27371 244260 27383 245036
rect 27321 244248 27383 244260
<< ndiffc >>
rect -4049 263250 -4015 264026
rect -3953 263250 -3919 264026
rect -3839 263250 -3805 264026
rect -3743 263250 -3709 264026
rect -3629 263250 -3595 264026
rect -3533 263250 -3499 264026
rect -3419 263250 -3385 264026
rect -3323 263250 -3289 264026
rect -3209 263250 -3175 264026
rect -3113 263250 -3079 264026
rect -2999 263250 -2965 264026
rect -2903 263250 -2869 264026
rect -2789 263250 -2755 264026
rect -2693 263250 -2659 264026
rect -2579 263250 -2545 264026
rect -2483 263250 -2449 264026
rect -2369 263250 -2335 264026
rect -2273 263250 -2239 264026
rect -2159 263250 -2125 264026
rect -2063 263250 -2029 264026
rect -1949 263250 -1915 264026
rect -1853 263250 -1819 264026
rect -1739 263250 -1705 264026
rect -1643 263250 -1609 264026
rect -1529 263250 -1495 264026
rect -1433 263250 -1399 264026
rect -1319 263250 -1285 264026
rect -1223 263250 -1189 264026
rect -1109 263250 -1075 264026
rect -1013 263250 -979 264026
rect -899 263250 -865 264026
rect -803 263250 -769 264026
rect -689 263250 -655 264026
rect -593 263250 -559 264026
rect -479 263250 -445 264026
rect -383 263250 -349 264026
rect -269 263250 -235 264026
rect -173 263250 -139 264026
rect -59 263250 -25 264026
rect 37 263250 71 264026
rect 151 263250 185 264026
rect 247 263250 281 264026
rect 361 263250 395 264026
rect 457 263250 491 264026
rect 571 263250 605 264026
rect 667 263250 701 264026
rect 781 263250 815 264026
rect 877 263250 911 264026
rect 991 263250 1025 264026
rect 1087 263250 1121 264026
rect 1201 263250 1235 264026
rect 1297 263250 1331 264026
rect 1411 263250 1445 264026
rect 1507 263250 1541 264026
rect 1621 263250 1655 264026
rect 1717 263250 1751 264026
rect 1831 263250 1865 264026
rect 1927 263250 1961 264026
rect 2041 263250 2075 264026
rect 2137 263250 2171 264026
rect 2251 263250 2285 264026
rect 2347 263250 2381 264026
rect 2461 263250 2495 264026
rect 2557 263250 2591 264026
rect 2671 263250 2705 264026
rect 2767 263250 2801 264026
rect 2881 263250 2915 264026
rect 2977 263250 3011 264026
rect 3091 263250 3125 264026
rect 3187 263250 3221 264026
rect 3301 263250 3335 264026
rect 3397 263250 3431 264026
rect 3511 263250 3545 264026
rect 3607 263250 3641 264026
rect 3721 263250 3755 264026
rect 3817 263250 3851 264026
rect 3931 263250 3965 264026
rect 4027 263250 4061 264026
rect 4141 263250 4175 264026
rect 4237 263250 4271 264026
rect 4351 263250 4385 264026
rect 4447 263250 4481 264026
rect 4561 263250 4595 264026
rect 4657 263250 4691 264026
rect 4771 263250 4805 264026
rect 4867 263250 4901 264026
rect 4981 263250 5015 264026
rect 5077 263250 5111 264026
rect 5191 263250 5225 264026
rect 5287 263250 5321 264026
rect 5401 263250 5435 264026
rect 5497 263250 5531 264026
rect 5611 263250 5645 264026
rect 5707 263250 5741 264026
rect 5821 263250 5855 264026
rect 5917 263250 5951 264026
rect 6031 263250 6065 264026
rect 6127 263250 6161 264026
rect 6241 263250 6275 264026
rect 6337 263250 6371 264026
rect 6451 263250 6485 264026
rect 6547 263250 6581 264026
rect 6661 263250 6695 264026
rect 6757 263250 6791 264026
rect 6871 263250 6905 264026
rect 6967 263250 7001 264026
rect 7081 263250 7115 264026
rect 7177 263250 7211 264026
rect 7291 263250 7325 264026
rect 7387 263250 7421 264026
rect 7501 263250 7535 264026
rect 7597 263250 7631 264026
rect 7711 263250 7745 264026
rect 7807 263250 7841 264026
rect 7921 263250 7955 264026
rect 8017 263250 8051 264026
rect 8131 263250 8165 264026
rect 8227 263250 8261 264026
rect 8341 263250 8375 264026
rect 8437 263250 8471 264026
rect 8551 263250 8585 264026
rect 8647 263250 8681 264026
rect 8761 263250 8795 264026
rect 8857 263250 8891 264026
rect 8971 263250 9005 264026
rect 9067 263250 9101 264026
rect 9181 263250 9215 264026
rect 9277 263250 9311 264026
rect 9391 263250 9425 264026
rect 9487 263250 9521 264026
rect 9601 263250 9635 264026
rect 9697 263250 9731 264026
rect 9811 263250 9845 264026
rect 9907 263250 9941 264026
rect 10021 263250 10055 264026
rect 10117 263250 10151 264026
rect 10231 263250 10265 264026
rect 10327 263250 10361 264026
rect 10441 263250 10475 264026
rect 10537 263250 10571 264026
rect 10651 263250 10685 264026
rect 10747 263250 10781 264026
rect 10861 263250 10895 264026
rect 10957 263250 10991 264026
rect 11071 263250 11105 264026
rect 11167 263250 11201 264026
rect 11281 263250 11315 264026
rect 11377 263250 11411 264026
rect 11491 263250 11525 264026
rect 11587 263250 11621 264026
rect 11701 263250 11735 264026
rect 11797 263250 11831 264026
rect 11911 263250 11945 264026
rect 12007 263250 12041 264026
rect 12121 263250 12155 264026
rect 12217 263250 12251 264026
rect 12331 263250 12365 264026
rect 12427 263250 12461 264026
rect 12541 263250 12575 264026
rect 12637 263250 12671 264026
rect 12751 263250 12785 264026
rect 12847 263250 12881 264026
rect 12961 263250 12995 264026
rect 13057 263250 13091 264026
rect 13171 263250 13205 264026
rect 13267 263250 13301 264026
rect 13381 263250 13415 264026
rect 13477 263250 13511 264026
rect 13591 263250 13625 264026
rect 13687 263250 13721 264026
rect 13801 263250 13835 264026
rect 13897 263250 13931 264026
rect 14011 263250 14045 264026
rect 14107 263250 14141 264026
rect 14221 263250 14255 264026
rect 14317 263250 14351 264026
rect 14431 263250 14465 264026
rect 14527 263250 14561 264026
rect 14641 263250 14675 264026
rect 14737 263250 14771 264026
rect 14851 263250 14885 264026
rect 14947 263250 14981 264026
rect 15061 263250 15095 264026
rect 15157 263250 15191 264026
rect 15271 263250 15305 264026
rect 15367 263250 15401 264026
rect 15481 263250 15515 264026
rect 15577 263250 15611 264026
rect 15691 263250 15725 264026
rect 15787 263250 15821 264026
rect 15901 263250 15935 264026
rect 15997 263250 16031 264026
rect 16111 263250 16145 264026
rect 16207 263250 16241 264026
rect 16321 263250 16355 264026
rect 16417 263250 16451 264026
rect 16531 263250 16565 264026
rect 16627 263250 16661 264026
rect 16741 263250 16775 264026
rect 16837 263250 16871 264026
rect 16951 263250 16985 264026
rect 17047 263250 17081 264026
rect 17161 263250 17195 264026
rect 17257 263250 17291 264026
rect 17371 263250 17405 264026
rect 17467 263250 17501 264026
rect 17581 263250 17615 264026
rect 17677 263250 17711 264026
rect 17791 263250 17825 264026
rect 17887 263250 17921 264026
rect 18001 263250 18035 264026
rect 18097 263250 18131 264026
rect 18211 263250 18245 264026
rect 18307 263250 18341 264026
rect 18421 263250 18455 264026
rect 18517 263250 18551 264026
rect 18631 263250 18665 264026
rect 18727 263250 18761 264026
rect 18841 263250 18875 264026
rect 18937 263250 18971 264026
rect 19051 263250 19085 264026
rect 19147 263250 19181 264026
rect 19261 263250 19295 264026
rect 19357 263250 19391 264026
rect 19471 263250 19505 264026
rect 19567 263250 19601 264026
rect 19681 263250 19715 264026
rect 19777 263250 19811 264026
rect 19891 263250 19925 264026
rect 19987 263250 20021 264026
rect 20101 263250 20135 264026
rect 20197 263250 20231 264026
rect 20311 263250 20345 264026
rect 20407 263250 20441 264026
rect 20521 263250 20555 264026
rect 20617 263250 20651 264026
rect 20731 263250 20765 264026
rect 20827 263250 20861 264026
rect 20941 263250 20975 264026
rect 21037 263250 21071 264026
rect 21151 263250 21185 264026
rect 21247 263250 21281 264026
rect 21361 263250 21395 264026
rect 21457 263250 21491 264026
rect 21571 263250 21605 264026
rect 21667 263250 21701 264026
rect 21781 263250 21815 264026
rect 21877 263250 21911 264026
rect 21991 263250 22025 264026
rect 22087 263250 22121 264026
rect 22201 263250 22235 264026
rect 22297 263250 22331 264026
rect 22411 263250 22445 264026
rect 22507 263250 22541 264026
rect 22621 263250 22655 264026
rect 22717 263250 22751 264026
rect 22831 263250 22865 264026
rect 22927 263250 22961 264026
rect 23041 263250 23075 264026
rect 23137 263250 23171 264026
rect 23251 263250 23285 264026
rect 23347 263250 23381 264026
rect 23461 263250 23495 264026
rect 23557 263250 23591 264026
rect 23671 263250 23705 264026
rect 23767 263250 23801 264026
rect 23881 263250 23915 264026
rect 23977 263250 24011 264026
rect 24091 263250 24125 264026
rect 24187 263250 24221 264026
rect 24301 263250 24335 264026
rect 24397 263250 24431 264026
rect 24511 263250 24545 264026
rect 24607 263250 24641 264026
rect 24721 263250 24755 264026
rect 24817 263250 24851 264026
rect 24931 263250 24965 264026
rect 25027 263250 25061 264026
rect 25141 263250 25175 264026
rect 25237 263250 25271 264026
rect 25351 263250 25385 264026
rect 25447 263250 25481 264026
rect 25561 263250 25595 264026
rect 25657 263250 25691 264026
rect 25771 263250 25805 264026
rect 25867 263250 25901 264026
rect 25981 263250 26015 264026
rect 26077 263250 26111 264026
rect 26191 263250 26225 264026
rect 26287 263250 26321 264026
rect 26401 263250 26435 264026
rect 26497 263250 26531 264026
rect 26611 263250 26645 264026
rect 26707 263250 26741 264026
rect 26821 263250 26855 264026
rect 26917 263250 26951 264026
rect 27031 263250 27065 264026
rect 27127 263250 27161 264026
rect 27241 263250 27275 264026
rect 27337 263250 27371 264026
rect -4049 262228 -4015 263004
rect -3953 262228 -3919 263004
rect -3839 262228 -3805 263004
rect -3743 262228 -3709 263004
rect -3629 262228 -3595 263004
rect -3533 262228 -3499 263004
rect -3419 262228 -3385 263004
rect -3323 262228 -3289 263004
rect -3209 262228 -3175 263004
rect -3113 262228 -3079 263004
rect -2999 262228 -2965 263004
rect -2903 262228 -2869 263004
rect -2789 262228 -2755 263004
rect -2693 262228 -2659 263004
rect -2579 262228 -2545 263004
rect -2483 262228 -2449 263004
rect -2369 262228 -2335 263004
rect -2273 262228 -2239 263004
rect -2159 262228 -2125 263004
rect -2063 262228 -2029 263004
rect -1949 262228 -1915 263004
rect -1853 262228 -1819 263004
rect -1739 262228 -1705 263004
rect -1643 262228 -1609 263004
rect -1529 262228 -1495 263004
rect -1433 262228 -1399 263004
rect -1319 262228 -1285 263004
rect -1223 262228 -1189 263004
rect -1109 262228 -1075 263004
rect -1013 262228 -979 263004
rect -899 262228 -865 263004
rect -803 262228 -769 263004
rect -689 262228 -655 263004
rect -593 262228 -559 263004
rect -479 262228 -445 263004
rect -383 262228 -349 263004
rect -269 262228 -235 263004
rect -173 262228 -139 263004
rect -59 262228 -25 263004
rect 37 262228 71 263004
rect 151 262228 185 263004
rect 247 262228 281 263004
rect 361 262228 395 263004
rect 457 262228 491 263004
rect 571 262228 605 263004
rect 667 262228 701 263004
rect 781 262228 815 263004
rect 877 262228 911 263004
rect 991 262228 1025 263004
rect 1087 262228 1121 263004
rect 1201 262228 1235 263004
rect 1297 262228 1331 263004
rect 1411 262228 1445 263004
rect 1507 262228 1541 263004
rect 1621 262228 1655 263004
rect 1717 262228 1751 263004
rect 1831 262228 1865 263004
rect 1927 262228 1961 263004
rect 2041 262228 2075 263004
rect 2137 262228 2171 263004
rect 2251 262228 2285 263004
rect 2347 262228 2381 263004
rect 2461 262228 2495 263004
rect 2557 262228 2591 263004
rect 2671 262228 2705 263004
rect 2767 262228 2801 263004
rect 2881 262228 2915 263004
rect 2977 262228 3011 263004
rect 3091 262228 3125 263004
rect 3187 262228 3221 263004
rect 3301 262228 3335 263004
rect 3397 262228 3431 263004
rect 3511 262228 3545 263004
rect 3607 262228 3641 263004
rect 3721 262228 3755 263004
rect 3817 262228 3851 263004
rect 3931 262228 3965 263004
rect 4027 262228 4061 263004
rect 4141 262228 4175 263004
rect 4237 262228 4271 263004
rect 4351 262228 4385 263004
rect 4447 262228 4481 263004
rect 4561 262228 4595 263004
rect 4657 262228 4691 263004
rect 4771 262228 4805 263004
rect 4867 262228 4901 263004
rect 4981 262228 5015 263004
rect 5077 262228 5111 263004
rect 5191 262228 5225 263004
rect 5287 262228 5321 263004
rect 5401 262228 5435 263004
rect 5497 262228 5531 263004
rect 5611 262228 5645 263004
rect 5707 262228 5741 263004
rect 5821 262228 5855 263004
rect 5917 262228 5951 263004
rect 6031 262228 6065 263004
rect 6127 262228 6161 263004
rect 6241 262228 6275 263004
rect 6337 262228 6371 263004
rect 6451 262228 6485 263004
rect 6547 262228 6581 263004
rect 6661 262228 6695 263004
rect 6757 262228 6791 263004
rect 6871 262228 6905 263004
rect 6967 262228 7001 263004
rect 7081 262228 7115 263004
rect 7177 262228 7211 263004
rect 7291 262228 7325 263004
rect 7387 262228 7421 263004
rect 7501 262228 7535 263004
rect 7597 262228 7631 263004
rect 7711 262228 7745 263004
rect 7807 262228 7841 263004
rect 7921 262228 7955 263004
rect 8017 262228 8051 263004
rect 8131 262228 8165 263004
rect 8227 262228 8261 263004
rect 8341 262228 8375 263004
rect 8437 262228 8471 263004
rect 8551 262228 8585 263004
rect 8647 262228 8681 263004
rect 8761 262228 8795 263004
rect 8857 262228 8891 263004
rect 8971 262228 9005 263004
rect 9067 262228 9101 263004
rect 9181 262228 9215 263004
rect 9277 262228 9311 263004
rect 9391 262228 9425 263004
rect 9487 262228 9521 263004
rect 9601 262228 9635 263004
rect 9697 262228 9731 263004
rect 9811 262228 9845 263004
rect 9907 262228 9941 263004
rect 10021 262228 10055 263004
rect 10117 262228 10151 263004
rect 10231 262228 10265 263004
rect 10327 262228 10361 263004
rect 10441 262228 10475 263004
rect 10537 262228 10571 263004
rect 10651 262228 10685 263004
rect 10747 262228 10781 263004
rect 10861 262228 10895 263004
rect 10957 262228 10991 263004
rect 11071 262228 11105 263004
rect 11167 262228 11201 263004
rect 11281 262228 11315 263004
rect 11377 262228 11411 263004
rect 11491 262228 11525 263004
rect 11587 262228 11621 263004
rect 11701 262228 11735 263004
rect 11797 262228 11831 263004
rect 11911 262228 11945 263004
rect 12007 262228 12041 263004
rect 12121 262228 12155 263004
rect 12217 262228 12251 263004
rect 12331 262228 12365 263004
rect 12427 262228 12461 263004
rect 12541 262228 12575 263004
rect 12637 262228 12671 263004
rect 12751 262228 12785 263004
rect 12847 262228 12881 263004
rect 12961 262228 12995 263004
rect 13057 262228 13091 263004
rect 13171 262228 13205 263004
rect 13267 262228 13301 263004
rect 13381 262228 13415 263004
rect 13477 262228 13511 263004
rect 13591 262228 13625 263004
rect 13687 262228 13721 263004
rect 13801 262228 13835 263004
rect 13897 262228 13931 263004
rect 14011 262228 14045 263004
rect 14107 262228 14141 263004
rect 14221 262228 14255 263004
rect 14317 262228 14351 263004
rect 14431 262228 14465 263004
rect 14527 262228 14561 263004
rect 14641 262228 14675 263004
rect 14737 262228 14771 263004
rect 14851 262228 14885 263004
rect 14947 262228 14981 263004
rect 15061 262228 15095 263004
rect 15157 262228 15191 263004
rect 15271 262228 15305 263004
rect 15367 262228 15401 263004
rect 15481 262228 15515 263004
rect 15577 262228 15611 263004
rect 15691 262228 15725 263004
rect 15787 262228 15821 263004
rect 15901 262228 15935 263004
rect 15997 262228 16031 263004
rect 16111 262228 16145 263004
rect 16207 262228 16241 263004
rect 16321 262228 16355 263004
rect 16417 262228 16451 263004
rect 16531 262228 16565 263004
rect 16627 262228 16661 263004
rect 16741 262228 16775 263004
rect 16837 262228 16871 263004
rect 16951 262228 16985 263004
rect 17047 262228 17081 263004
rect 17161 262228 17195 263004
rect 17257 262228 17291 263004
rect 17371 262228 17405 263004
rect 17467 262228 17501 263004
rect 17581 262228 17615 263004
rect 17677 262228 17711 263004
rect 17791 262228 17825 263004
rect 17887 262228 17921 263004
rect 18001 262228 18035 263004
rect 18097 262228 18131 263004
rect 18211 262228 18245 263004
rect 18307 262228 18341 263004
rect 18421 262228 18455 263004
rect 18517 262228 18551 263004
rect 18631 262228 18665 263004
rect 18727 262228 18761 263004
rect 18841 262228 18875 263004
rect 18937 262228 18971 263004
rect 19051 262228 19085 263004
rect 19147 262228 19181 263004
rect 19261 262228 19295 263004
rect 19357 262228 19391 263004
rect 19471 262228 19505 263004
rect 19567 262228 19601 263004
rect 19681 262228 19715 263004
rect 19777 262228 19811 263004
rect 19891 262228 19925 263004
rect 19987 262228 20021 263004
rect 20101 262228 20135 263004
rect 20197 262228 20231 263004
rect 20311 262228 20345 263004
rect 20407 262228 20441 263004
rect 20521 262228 20555 263004
rect 20617 262228 20651 263004
rect 20731 262228 20765 263004
rect 20827 262228 20861 263004
rect 20941 262228 20975 263004
rect 21037 262228 21071 263004
rect 21151 262228 21185 263004
rect 21247 262228 21281 263004
rect 21361 262228 21395 263004
rect 21457 262228 21491 263004
rect 21571 262228 21605 263004
rect 21667 262228 21701 263004
rect 21781 262228 21815 263004
rect 21877 262228 21911 263004
rect 21991 262228 22025 263004
rect 22087 262228 22121 263004
rect 22201 262228 22235 263004
rect 22297 262228 22331 263004
rect 22411 262228 22445 263004
rect 22507 262228 22541 263004
rect 22621 262228 22655 263004
rect 22717 262228 22751 263004
rect 22831 262228 22865 263004
rect 22927 262228 22961 263004
rect 23041 262228 23075 263004
rect 23137 262228 23171 263004
rect 23251 262228 23285 263004
rect 23347 262228 23381 263004
rect 23461 262228 23495 263004
rect 23557 262228 23591 263004
rect 23671 262228 23705 263004
rect 23767 262228 23801 263004
rect 23881 262228 23915 263004
rect 23977 262228 24011 263004
rect 24091 262228 24125 263004
rect 24187 262228 24221 263004
rect 24301 262228 24335 263004
rect 24397 262228 24431 263004
rect 24511 262228 24545 263004
rect 24607 262228 24641 263004
rect 24721 262228 24755 263004
rect 24817 262228 24851 263004
rect 24931 262228 24965 263004
rect 25027 262228 25061 263004
rect 25141 262228 25175 263004
rect 25237 262228 25271 263004
rect 25351 262228 25385 263004
rect 25447 262228 25481 263004
rect 25561 262228 25595 263004
rect 25657 262228 25691 263004
rect 25771 262228 25805 263004
rect 25867 262228 25901 263004
rect 25981 262228 26015 263004
rect 26077 262228 26111 263004
rect 26191 262228 26225 263004
rect 26287 262228 26321 263004
rect 26401 262228 26435 263004
rect 26497 262228 26531 263004
rect 26611 262228 26645 263004
rect 26707 262228 26741 263004
rect 26821 262228 26855 263004
rect 26917 262228 26951 263004
rect 27031 262228 27065 263004
rect 27127 262228 27161 263004
rect 27241 262228 27275 263004
rect 27337 262228 27371 263004
<< pdiffc >>
rect -4049 253713 -4015 254489
rect -3953 253713 -3919 254489
rect -3839 253713 -3805 254489
rect -3743 253713 -3709 254489
rect -3629 253713 -3595 254489
rect -3533 253713 -3499 254489
rect -3419 253713 -3385 254489
rect -3323 253713 -3289 254489
rect -3209 253713 -3175 254489
rect -3113 253713 -3079 254489
rect -2999 253713 -2965 254489
rect -2903 253713 -2869 254489
rect -2789 253713 -2755 254489
rect -2693 253713 -2659 254489
rect -2579 253713 -2545 254489
rect -2483 253713 -2449 254489
rect -2369 253713 -2335 254489
rect -2273 253713 -2239 254489
rect -2159 253713 -2125 254489
rect -2063 253713 -2029 254489
rect -1949 253713 -1915 254489
rect -1853 253713 -1819 254489
rect -1739 253713 -1705 254489
rect -1643 253713 -1609 254489
rect -1529 253713 -1495 254489
rect -1433 253713 -1399 254489
rect -1319 253713 -1285 254489
rect -1223 253713 -1189 254489
rect -1109 253713 -1075 254489
rect -1013 253713 -979 254489
rect -899 253713 -865 254489
rect -803 253713 -769 254489
rect -689 253713 -655 254489
rect -593 253713 -559 254489
rect -479 253713 -445 254489
rect -383 253713 -349 254489
rect -269 253713 -235 254489
rect -173 253713 -139 254489
rect -59 253713 -25 254489
rect 37 253713 71 254489
rect 151 253713 185 254489
rect 247 253713 281 254489
rect 361 253713 395 254489
rect 457 253713 491 254489
rect 571 253713 605 254489
rect 667 253713 701 254489
rect 781 253713 815 254489
rect 877 253713 911 254489
rect 991 253713 1025 254489
rect 1087 253713 1121 254489
rect 1201 253713 1235 254489
rect 1297 253713 1331 254489
rect 1411 253713 1445 254489
rect 1507 253713 1541 254489
rect 1621 253713 1655 254489
rect 1717 253713 1751 254489
rect 1831 253713 1865 254489
rect 1927 253713 1961 254489
rect 2041 253713 2075 254489
rect 2137 253713 2171 254489
rect 2251 253713 2285 254489
rect 2347 253713 2381 254489
rect 2461 253713 2495 254489
rect 2557 253713 2591 254489
rect 2671 253713 2705 254489
rect 2767 253713 2801 254489
rect 2881 253713 2915 254489
rect 2977 253713 3011 254489
rect 3091 253713 3125 254489
rect 3187 253713 3221 254489
rect 3301 253713 3335 254489
rect 3397 253713 3431 254489
rect 3511 253713 3545 254489
rect 3607 253713 3641 254489
rect 3721 253713 3755 254489
rect 3817 253713 3851 254489
rect 3931 253713 3965 254489
rect 4027 253713 4061 254489
rect 4141 253713 4175 254489
rect 4237 253713 4271 254489
rect 4351 253713 4385 254489
rect 4447 253713 4481 254489
rect 4561 253713 4595 254489
rect 4657 253713 4691 254489
rect 4771 253713 4805 254489
rect 4867 253713 4901 254489
rect 4981 253713 5015 254489
rect 5077 253713 5111 254489
rect 5191 253713 5225 254489
rect 5287 253713 5321 254489
rect 5401 253713 5435 254489
rect 5497 253713 5531 254489
rect 5611 253713 5645 254489
rect 5707 253713 5741 254489
rect 5821 253713 5855 254489
rect 5917 253713 5951 254489
rect 6031 253713 6065 254489
rect 6127 253713 6161 254489
rect 6241 253713 6275 254489
rect 6337 253713 6371 254489
rect 6451 253713 6485 254489
rect 6547 253713 6581 254489
rect 6661 253713 6695 254489
rect 6757 253713 6791 254489
rect 6871 253713 6905 254489
rect 6967 253713 7001 254489
rect 7081 253713 7115 254489
rect 7177 253713 7211 254489
rect 7291 253713 7325 254489
rect 7387 253713 7421 254489
rect 7501 253713 7535 254489
rect 7597 253713 7631 254489
rect 7711 253713 7745 254489
rect 7807 253713 7841 254489
rect 7921 253713 7955 254489
rect 8017 253713 8051 254489
rect 8131 253713 8165 254489
rect 8227 253713 8261 254489
rect 8341 253713 8375 254489
rect 8437 253713 8471 254489
rect 8551 253713 8585 254489
rect 8647 253713 8681 254489
rect 8761 253713 8795 254489
rect 8857 253713 8891 254489
rect 8971 253713 9005 254489
rect 9067 253713 9101 254489
rect 9181 253713 9215 254489
rect 9277 253713 9311 254489
rect 9391 253713 9425 254489
rect 9487 253713 9521 254489
rect 9601 253713 9635 254489
rect 9697 253713 9731 254489
rect 9811 253713 9845 254489
rect 9907 253713 9941 254489
rect 10021 253713 10055 254489
rect 10117 253713 10151 254489
rect 10231 253713 10265 254489
rect 10327 253713 10361 254489
rect 10441 253713 10475 254489
rect 10537 253713 10571 254489
rect 10651 253713 10685 254489
rect 10747 253713 10781 254489
rect 10861 253713 10895 254489
rect 10957 253713 10991 254489
rect 11071 253713 11105 254489
rect 11167 253713 11201 254489
rect 11281 253713 11315 254489
rect 11377 253713 11411 254489
rect 11491 253713 11525 254489
rect 11587 253713 11621 254489
rect 11701 253713 11735 254489
rect 11797 253713 11831 254489
rect 11911 253713 11945 254489
rect 12007 253713 12041 254489
rect 12121 253713 12155 254489
rect 12217 253713 12251 254489
rect 12331 253713 12365 254489
rect 12427 253713 12461 254489
rect 12541 253713 12575 254489
rect 12637 253713 12671 254489
rect 12751 253713 12785 254489
rect 12847 253713 12881 254489
rect 12961 253713 12995 254489
rect 13057 253713 13091 254489
rect 13171 253713 13205 254489
rect 13267 253713 13301 254489
rect 13381 253713 13415 254489
rect 13477 253713 13511 254489
rect 13591 253713 13625 254489
rect 13687 253713 13721 254489
rect 13801 253713 13835 254489
rect 13897 253713 13931 254489
rect 14011 253713 14045 254489
rect 14107 253713 14141 254489
rect 14221 253713 14255 254489
rect 14317 253713 14351 254489
rect 14431 253713 14465 254489
rect 14527 253713 14561 254489
rect 14641 253713 14675 254489
rect 14737 253713 14771 254489
rect 14851 253713 14885 254489
rect 14947 253713 14981 254489
rect 15061 253713 15095 254489
rect 15157 253713 15191 254489
rect 15271 253713 15305 254489
rect 15367 253713 15401 254489
rect 15481 253713 15515 254489
rect 15577 253713 15611 254489
rect 15691 253713 15725 254489
rect 15787 253713 15821 254489
rect 15901 253713 15935 254489
rect 15997 253713 16031 254489
rect 16111 253713 16145 254489
rect 16207 253713 16241 254489
rect 16321 253713 16355 254489
rect 16417 253713 16451 254489
rect 16531 253713 16565 254489
rect 16627 253713 16661 254489
rect 16741 253713 16775 254489
rect 16837 253713 16871 254489
rect 16951 253713 16985 254489
rect 17047 253713 17081 254489
rect 17161 253713 17195 254489
rect 17257 253713 17291 254489
rect 17371 253713 17405 254489
rect 17467 253713 17501 254489
rect 17581 253713 17615 254489
rect 17677 253713 17711 254489
rect 17791 253713 17825 254489
rect 17887 253713 17921 254489
rect 18001 253713 18035 254489
rect 18097 253713 18131 254489
rect 18211 253713 18245 254489
rect 18307 253713 18341 254489
rect 18421 253713 18455 254489
rect 18517 253713 18551 254489
rect 18631 253713 18665 254489
rect 18727 253713 18761 254489
rect 18841 253713 18875 254489
rect 18937 253713 18971 254489
rect 19051 253713 19085 254489
rect 19147 253713 19181 254489
rect 19261 253713 19295 254489
rect 19357 253713 19391 254489
rect 19471 253713 19505 254489
rect 19567 253713 19601 254489
rect 19681 253713 19715 254489
rect 19777 253713 19811 254489
rect 19891 253713 19925 254489
rect 19987 253713 20021 254489
rect 20101 253713 20135 254489
rect 20197 253713 20231 254489
rect 20311 253713 20345 254489
rect 20407 253713 20441 254489
rect 20521 253713 20555 254489
rect 20617 253713 20651 254489
rect 20731 253713 20765 254489
rect 20827 253713 20861 254489
rect 20941 253713 20975 254489
rect 21037 253713 21071 254489
rect 21151 253713 21185 254489
rect 21247 253713 21281 254489
rect 21361 253713 21395 254489
rect 21457 253713 21491 254489
rect 21571 253713 21605 254489
rect 21667 253713 21701 254489
rect 21781 253713 21815 254489
rect 21877 253713 21911 254489
rect 21991 253713 22025 254489
rect 22087 253713 22121 254489
rect 22201 253713 22235 254489
rect 22297 253713 22331 254489
rect 22411 253713 22445 254489
rect 22507 253713 22541 254489
rect 22621 253713 22655 254489
rect 22717 253713 22751 254489
rect 22831 253713 22865 254489
rect 22927 253713 22961 254489
rect 23041 253713 23075 254489
rect 23137 253713 23171 254489
rect 23251 253713 23285 254489
rect 23347 253713 23381 254489
rect 23461 253713 23495 254489
rect 23557 253713 23591 254489
rect 23671 253713 23705 254489
rect 23767 253713 23801 254489
rect 23881 253713 23915 254489
rect 23977 253713 24011 254489
rect 24091 253713 24125 254489
rect 24187 253713 24221 254489
rect 24301 253713 24335 254489
rect 24397 253713 24431 254489
rect 24511 253713 24545 254489
rect 24607 253713 24641 254489
rect 24721 253713 24755 254489
rect 24817 253713 24851 254489
rect 24931 253713 24965 254489
rect 25027 253713 25061 254489
rect 25141 253713 25175 254489
rect 25237 253713 25271 254489
rect 25351 253713 25385 254489
rect 25447 253713 25481 254489
rect 25561 253713 25595 254489
rect 25657 253713 25691 254489
rect 25771 253713 25805 254489
rect 25867 253713 25901 254489
rect 25981 253713 26015 254489
rect 26077 253713 26111 254489
rect 26191 253713 26225 254489
rect 26287 253713 26321 254489
rect 26401 253713 26435 254489
rect 26497 253713 26531 254489
rect 26611 253713 26645 254489
rect 26707 253713 26741 254489
rect 26821 253713 26855 254489
rect 26917 253713 26951 254489
rect 27031 253713 27065 254489
rect 27127 253713 27161 254489
rect 27241 253713 27275 254489
rect 27337 253713 27371 254489
rect -4049 252677 -4015 253453
rect -3953 252677 -3919 253453
rect -3839 252677 -3805 253453
rect -3743 252677 -3709 253453
rect -3629 252677 -3595 253453
rect -3533 252677 -3499 253453
rect -3419 252677 -3385 253453
rect -3323 252677 -3289 253453
rect -3209 252677 -3175 253453
rect -3113 252677 -3079 253453
rect -2999 252677 -2965 253453
rect -2903 252677 -2869 253453
rect -2789 252677 -2755 253453
rect -2693 252677 -2659 253453
rect -2579 252677 -2545 253453
rect -2483 252677 -2449 253453
rect -2369 252677 -2335 253453
rect -2273 252677 -2239 253453
rect -2159 252677 -2125 253453
rect -2063 252677 -2029 253453
rect -1949 252677 -1915 253453
rect -1853 252677 -1819 253453
rect -1739 252677 -1705 253453
rect -1643 252677 -1609 253453
rect -1529 252677 -1495 253453
rect -1433 252677 -1399 253453
rect -1319 252677 -1285 253453
rect -1223 252677 -1189 253453
rect -1109 252677 -1075 253453
rect -1013 252677 -979 253453
rect -899 252677 -865 253453
rect -803 252677 -769 253453
rect -689 252677 -655 253453
rect -593 252677 -559 253453
rect -479 252677 -445 253453
rect -383 252677 -349 253453
rect -269 252677 -235 253453
rect -173 252677 -139 253453
rect -59 252677 -25 253453
rect 37 252677 71 253453
rect 151 252677 185 253453
rect 247 252677 281 253453
rect 361 252677 395 253453
rect 457 252677 491 253453
rect 571 252677 605 253453
rect 667 252677 701 253453
rect 781 252677 815 253453
rect 877 252677 911 253453
rect 991 252677 1025 253453
rect 1087 252677 1121 253453
rect 1201 252677 1235 253453
rect 1297 252677 1331 253453
rect 1411 252677 1445 253453
rect 1507 252677 1541 253453
rect 1621 252677 1655 253453
rect 1717 252677 1751 253453
rect 1831 252677 1865 253453
rect 1927 252677 1961 253453
rect 2041 252677 2075 253453
rect 2137 252677 2171 253453
rect 2251 252677 2285 253453
rect 2347 252677 2381 253453
rect 2461 252677 2495 253453
rect 2557 252677 2591 253453
rect 2671 252677 2705 253453
rect 2767 252677 2801 253453
rect 2881 252677 2915 253453
rect 2977 252677 3011 253453
rect 3091 252677 3125 253453
rect 3187 252677 3221 253453
rect 3301 252677 3335 253453
rect 3397 252677 3431 253453
rect 3511 252677 3545 253453
rect 3607 252677 3641 253453
rect 3721 252677 3755 253453
rect 3817 252677 3851 253453
rect 3931 252677 3965 253453
rect 4027 252677 4061 253453
rect 4141 252677 4175 253453
rect 4237 252677 4271 253453
rect 4351 252677 4385 253453
rect 4447 252677 4481 253453
rect 4561 252677 4595 253453
rect 4657 252677 4691 253453
rect 4771 252677 4805 253453
rect 4867 252677 4901 253453
rect 4981 252677 5015 253453
rect 5077 252677 5111 253453
rect 5191 252677 5225 253453
rect 5287 252677 5321 253453
rect 5401 252677 5435 253453
rect 5497 252677 5531 253453
rect 5611 252677 5645 253453
rect 5707 252677 5741 253453
rect 5821 252677 5855 253453
rect 5917 252677 5951 253453
rect 6031 252677 6065 253453
rect 6127 252677 6161 253453
rect 6241 252677 6275 253453
rect 6337 252677 6371 253453
rect 6451 252677 6485 253453
rect 6547 252677 6581 253453
rect 6661 252677 6695 253453
rect 6757 252677 6791 253453
rect 6871 252677 6905 253453
rect 6967 252677 7001 253453
rect 7081 252677 7115 253453
rect 7177 252677 7211 253453
rect 7291 252677 7325 253453
rect 7387 252677 7421 253453
rect 7501 252677 7535 253453
rect 7597 252677 7631 253453
rect 7711 252677 7745 253453
rect 7807 252677 7841 253453
rect 7921 252677 7955 253453
rect 8017 252677 8051 253453
rect 8131 252677 8165 253453
rect 8227 252677 8261 253453
rect 8341 252677 8375 253453
rect 8437 252677 8471 253453
rect 8551 252677 8585 253453
rect 8647 252677 8681 253453
rect 8761 252677 8795 253453
rect 8857 252677 8891 253453
rect 8971 252677 9005 253453
rect 9067 252677 9101 253453
rect 9181 252677 9215 253453
rect 9277 252677 9311 253453
rect 9391 252677 9425 253453
rect 9487 252677 9521 253453
rect 9601 252677 9635 253453
rect 9697 252677 9731 253453
rect 9811 252677 9845 253453
rect 9907 252677 9941 253453
rect 10021 252677 10055 253453
rect 10117 252677 10151 253453
rect 10231 252677 10265 253453
rect 10327 252677 10361 253453
rect 10441 252677 10475 253453
rect 10537 252677 10571 253453
rect 10651 252677 10685 253453
rect 10747 252677 10781 253453
rect 10861 252677 10895 253453
rect 10957 252677 10991 253453
rect 11071 252677 11105 253453
rect 11167 252677 11201 253453
rect 11281 252677 11315 253453
rect 11377 252677 11411 253453
rect 11491 252677 11525 253453
rect 11587 252677 11621 253453
rect 11701 252677 11735 253453
rect 11797 252677 11831 253453
rect 11911 252677 11945 253453
rect 12007 252677 12041 253453
rect 12121 252677 12155 253453
rect 12217 252677 12251 253453
rect 12331 252677 12365 253453
rect 12427 252677 12461 253453
rect 12541 252677 12575 253453
rect 12637 252677 12671 253453
rect 12751 252677 12785 253453
rect 12847 252677 12881 253453
rect 12961 252677 12995 253453
rect 13057 252677 13091 253453
rect 13171 252677 13205 253453
rect 13267 252677 13301 253453
rect 13381 252677 13415 253453
rect 13477 252677 13511 253453
rect 13591 252677 13625 253453
rect 13687 252677 13721 253453
rect 13801 252677 13835 253453
rect 13897 252677 13931 253453
rect 14011 252677 14045 253453
rect 14107 252677 14141 253453
rect 14221 252677 14255 253453
rect 14317 252677 14351 253453
rect 14431 252677 14465 253453
rect 14527 252677 14561 253453
rect 14641 252677 14675 253453
rect 14737 252677 14771 253453
rect 14851 252677 14885 253453
rect 14947 252677 14981 253453
rect 15061 252677 15095 253453
rect 15157 252677 15191 253453
rect 15271 252677 15305 253453
rect 15367 252677 15401 253453
rect 15481 252677 15515 253453
rect 15577 252677 15611 253453
rect 15691 252677 15725 253453
rect 15787 252677 15821 253453
rect 15901 252677 15935 253453
rect 15997 252677 16031 253453
rect 16111 252677 16145 253453
rect 16207 252677 16241 253453
rect 16321 252677 16355 253453
rect 16417 252677 16451 253453
rect 16531 252677 16565 253453
rect 16627 252677 16661 253453
rect 16741 252677 16775 253453
rect 16837 252677 16871 253453
rect 16951 252677 16985 253453
rect 17047 252677 17081 253453
rect 17161 252677 17195 253453
rect 17257 252677 17291 253453
rect 17371 252677 17405 253453
rect 17467 252677 17501 253453
rect 17581 252677 17615 253453
rect 17677 252677 17711 253453
rect 17791 252677 17825 253453
rect 17887 252677 17921 253453
rect 18001 252677 18035 253453
rect 18097 252677 18131 253453
rect 18211 252677 18245 253453
rect 18307 252677 18341 253453
rect 18421 252677 18455 253453
rect 18517 252677 18551 253453
rect 18631 252677 18665 253453
rect 18727 252677 18761 253453
rect 18841 252677 18875 253453
rect 18937 252677 18971 253453
rect 19051 252677 19085 253453
rect 19147 252677 19181 253453
rect 19261 252677 19295 253453
rect 19357 252677 19391 253453
rect 19471 252677 19505 253453
rect 19567 252677 19601 253453
rect 19681 252677 19715 253453
rect 19777 252677 19811 253453
rect 19891 252677 19925 253453
rect 19987 252677 20021 253453
rect 20101 252677 20135 253453
rect 20197 252677 20231 253453
rect 20311 252677 20345 253453
rect 20407 252677 20441 253453
rect 20521 252677 20555 253453
rect 20617 252677 20651 253453
rect 20731 252677 20765 253453
rect 20827 252677 20861 253453
rect 20941 252677 20975 253453
rect 21037 252677 21071 253453
rect 21151 252677 21185 253453
rect 21247 252677 21281 253453
rect 21361 252677 21395 253453
rect 21457 252677 21491 253453
rect 21571 252677 21605 253453
rect 21667 252677 21701 253453
rect 21781 252677 21815 253453
rect 21877 252677 21911 253453
rect 21991 252677 22025 253453
rect 22087 252677 22121 253453
rect 22201 252677 22235 253453
rect 22297 252677 22331 253453
rect 22411 252677 22445 253453
rect 22507 252677 22541 253453
rect 22621 252677 22655 253453
rect 22717 252677 22751 253453
rect 22831 252677 22865 253453
rect 22927 252677 22961 253453
rect 23041 252677 23075 253453
rect 23137 252677 23171 253453
rect 23251 252677 23285 253453
rect 23347 252677 23381 253453
rect 23461 252677 23495 253453
rect 23557 252677 23591 253453
rect 23671 252677 23705 253453
rect 23767 252677 23801 253453
rect 23881 252677 23915 253453
rect 23977 252677 24011 253453
rect 24091 252677 24125 253453
rect 24187 252677 24221 253453
rect 24301 252677 24335 253453
rect 24397 252677 24431 253453
rect 24511 252677 24545 253453
rect 24607 252677 24641 253453
rect 24721 252677 24755 253453
rect 24817 252677 24851 253453
rect 24931 252677 24965 253453
rect 25027 252677 25061 253453
rect 25141 252677 25175 253453
rect 25237 252677 25271 253453
rect 25351 252677 25385 253453
rect 25447 252677 25481 253453
rect 25561 252677 25595 253453
rect 25657 252677 25691 253453
rect 25771 252677 25805 253453
rect 25867 252677 25901 253453
rect 25981 252677 26015 253453
rect 26077 252677 26111 253453
rect 26191 252677 26225 253453
rect 26287 252677 26321 253453
rect 26401 252677 26435 253453
rect 26497 252677 26531 253453
rect 26611 252677 26645 253453
rect 26707 252677 26741 253453
rect 26821 252677 26855 253453
rect 26917 252677 26951 253453
rect 27031 252677 27065 253453
rect 27127 252677 27161 253453
rect 27241 252677 27275 253453
rect 27337 252677 27371 253453
rect -4049 251641 -4015 252417
rect -3953 251641 -3919 252417
rect -3839 251641 -3805 252417
rect -3743 251641 -3709 252417
rect -3629 251641 -3595 252417
rect -3533 251641 -3499 252417
rect -3419 251641 -3385 252417
rect -3323 251641 -3289 252417
rect -3209 251641 -3175 252417
rect -3113 251641 -3079 252417
rect -2999 251641 -2965 252417
rect -2903 251641 -2869 252417
rect -2789 251641 -2755 252417
rect -2693 251641 -2659 252417
rect -2579 251641 -2545 252417
rect -2483 251641 -2449 252417
rect -2369 251641 -2335 252417
rect -2273 251641 -2239 252417
rect -2159 251641 -2125 252417
rect -2063 251641 -2029 252417
rect -1949 251641 -1915 252417
rect -1853 251641 -1819 252417
rect -1739 251641 -1705 252417
rect -1643 251641 -1609 252417
rect -1529 251641 -1495 252417
rect -1433 251641 -1399 252417
rect -1319 251641 -1285 252417
rect -1223 251641 -1189 252417
rect -1109 251641 -1075 252417
rect -1013 251641 -979 252417
rect -899 251641 -865 252417
rect -803 251641 -769 252417
rect -689 251641 -655 252417
rect -593 251641 -559 252417
rect -479 251641 -445 252417
rect -383 251641 -349 252417
rect -269 251641 -235 252417
rect -173 251641 -139 252417
rect -59 251641 -25 252417
rect 37 251641 71 252417
rect 151 251641 185 252417
rect 247 251641 281 252417
rect 361 251641 395 252417
rect 457 251641 491 252417
rect 571 251641 605 252417
rect 667 251641 701 252417
rect 781 251641 815 252417
rect 877 251641 911 252417
rect 991 251641 1025 252417
rect 1087 251641 1121 252417
rect 1201 251641 1235 252417
rect 1297 251641 1331 252417
rect 1411 251641 1445 252417
rect 1507 251641 1541 252417
rect 1621 251641 1655 252417
rect 1717 251641 1751 252417
rect 1831 251641 1865 252417
rect 1927 251641 1961 252417
rect 2041 251641 2075 252417
rect 2137 251641 2171 252417
rect 2251 251641 2285 252417
rect 2347 251641 2381 252417
rect 2461 251641 2495 252417
rect 2557 251641 2591 252417
rect 2671 251641 2705 252417
rect 2767 251641 2801 252417
rect 2881 251641 2915 252417
rect 2977 251641 3011 252417
rect 3091 251641 3125 252417
rect 3187 251641 3221 252417
rect 3301 251641 3335 252417
rect 3397 251641 3431 252417
rect 3511 251641 3545 252417
rect 3607 251641 3641 252417
rect 3721 251641 3755 252417
rect 3817 251641 3851 252417
rect 3931 251641 3965 252417
rect 4027 251641 4061 252417
rect 4141 251641 4175 252417
rect 4237 251641 4271 252417
rect 4351 251641 4385 252417
rect 4447 251641 4481 252417
rect 4561 251641 4595 252417
rect 4657 251641 4691 252417
rect 4771 251641 4805 252417
rect 4867 251641 4901 252417
rect 4981 251641 5015 252417
rect 5077 251641 5111 252417
rect 5191 251641 5225 252417
rect 5287 251641 5321 252417
rect 5401 251641 5435 252417
rect 5497 251641 5531 252417
rect 5611 251641 5645 252417
rect 5707 251641 5741 252417
rect 5821 251641 5855 252417
rect 5917 251641 5951 252417
rect 6031 251641 6065 252417
rect 6127 251641 6161 252417
rect 6241 251641 6275 252417
rect 6337 251641 6371 252417
rect 6451 251641 6485 252417
rect 6547 251641 6581 252417
rect 6661 251641 6695 252417
rect 6757 251641 6791 252417
rect 6871 251641 6905 252417
rect 6967 251641 7001 252417
rect 7081 251641 7115 252417
rect 7177 251641 7211 252417
rect 7291 251641 7325 252417
rect 7387 251641 7421 252417
rect 7501 251641 7535 252417
rect 7597 251641 7631 252417
rect 7711 251641 7745 252417
rect 7807 251641 7841 252417
rect 7921 251641 7955 252417
rect 8017 251641 8051 252417
rect 8131 251641 8165 252417
rect 8227 251641 8261 252417
rect 8341 251641 8375 252417
rect 8437 251641 8471 252417
rect 8551 251641 8585 252417
rect 8647 251641 8681 252417
rect 8761 251641 8795 252417
rect 8857 251641 8891 252417
rect 8971 251641 9005 252417
rect 9067 251641 9101 252417
rect 9181 251641 9215 252417
rect 9277 251641 9311 252417
rect 9391 251641 9425 252417
rect 9487 251641 9521 252417
rect 9601 251641 9635 252417
rect 9697 251641 9731 252417
rect 9811 251641 9845 252417
rect 9907 251641 9941 252417
rect 10021 251641 10055 252417
rect 10117 251641 10151 252417
rect 10231 251641 10265 252417
rect 10327 251641 10361 252417
rect 10441 251641 10475 252417
rect 10537 251641 10571 252417
rect 10651 251641 10685 252417
rect 10747 251641 10781 252417
rect 10861 251641 10895 252417
rect 10957 251641 10991 252417
rect 11071 251641 11105 252417
rect 11167 251641 11201 252417
rect 11281 251641 11315 252417
rect 11377 251641 11411 252417
rect 11491 251641 11525 252417
rect 11587 251641 11621 252417
rect 11701 251641 11735 252417
rect 11797 251641 11831 252417
rect 11911 251641 11945 252417
rect 12007 251641 12041 252417
rect 12121 251641 12155 252417
rect 12217 251641 12251 252417
rect 12331 251641 12365 252417
rect 12427 251641 12461 252417
rect 12541 251641 12575 252417
rect 12637 251641 12671 252417
rect 12751 251641 12785 252417
rect 12847 251641 12881 252417
rect 12961 251641 12995 252417
rect 13057 251641 13091 252417
rect 13171 251641 13205 252417
rect 13267 251641 13301 252417
rect 13381 251641 13415 252417
rect 13477 251641 13511 252417
rect 13591 251641 13625 252417
rect 13687 251641 13721 252417
rect 13801 251641 13835 252417
rect 13897 251641 13931 252417
rect 14011 251641 14045 252417
rect 14107 251641 14141 252417
rect 14221 251641 14255 252417
rect 14317 251641 14351 252417
rect 14431 251641 14465 252417
rect 14527 251641 14561 252417
rect 14641 251641 14675 252417
rect 14737 251641 14771 252417
rect 14851 251641 14885 252417
rect 14947 251641 14981 252417
rect 15061 251641 15095 252417
rect 15157 251641 15191 252417
rect 15271 251641 15305 252417
rect 15367 251641 15401 252417
rect 15481 251641 15515 252417
rect 15577 251641 15611 252417
rect 15691 251641 15725 252417
rect 15787 251641 15821 252417
rect 15901 251641 15935 252417
rect 15997 251641 16031 252417
rect 16111 251641 16145 252417
rect 16207 251641 16241 252417
rect 16321 251641 16355 252417
rect 16417 251641 16451 252417
rect 16531 251641 16565 252417
rect 16627 251641 16661 252417
rect 16741 251641 16775 252417
rect 16837 251641 16871 252417
rect 16951 251641 16985 252417
rect 17047 251641 17081 252417
rect 17161 251641 17195 252417
rect 17257 251641 17291 252417
rect 17371 251641 17405 252417
rect 17467 251641 17501 252417
rect 17581 251641 17615 252417
rect 17677 251641 17711 252417
rect 17791 251641 17825 252417
rect 17887 251641 17921 252417
rect 18001 251641 18035 252417
rect 18097 251641 18131 252417
rect 18211 251641 18245 252417
rect 18307 251641 18341 252417
rect 18421 251641 18455 252417
rect 18517 251641 18551 252417
rect 18631 251641 18665 252417
rect 18727 251641 18761 252417
rect 18841 251641 18875 252417
rect 18937 251641 18971 252417
rect 19051 251641 19085 252417
rect 19147 251641 19181 252417
rect 19261 251641 19295 252417
rect 19357 251641 19391 252417
rect 19471 251641 19505 252417
rect 19567 251641 19601 252417
rect 19681 251641 19715 252417
rect 19777 251641 19811 252417
rect 19891 251641 19925 252417
rect 19987 251641 20021 252417
rect 20101 251641 20135 252417
rect 20197 251641 20231 252417
rect 20311 251641 20345 252417
rect 20407 251641 20441 252417
rect 20521 251641 20555 252417
rect 20617 251641 20651 252417
rect 20731 251641 20765 252417
rect 20827 251641 20861 252417
rect 20941 251641 20975 252417
rect 21037 251641 21071 252417
rect 21151 251641 21185 252417
rect 21247 251641 21281 252417
rect 21361 251641 21395 252417
rect 21457 251641 21491 252417
rect 21571 251641 21605 252417
rect 21667 251641 21701 252417
rect 21781 251641 21815 252417
rect 21877 251641 21911 252417
rect 21991 251641 22025 252417
rect 22087 251641 22121 252417
rect 22201 251641 22235 252417
rect 22297 251641 22331 252417
rect 22411 251641 22445 252417
rect 22507 251641 22541 252417
rect 22621 251641 22655 252417
rect 22717 251641 22751 252417
rect 22831 251641 22865 252417
rect 22927 251641 22961 252417
rect 23041 251641 23075 252417
rect 23137 251641 23171 252417
rect 23251 251641 23285 252417
rect 23347 251641 23381 252417
rect 23461 251641 23495 252417
rect 23557 251641 23591 252417
rect 23671 251641 23705 252417
rect 23767 251641 23801 252417
rect 23881 251641 23915 252417
rect 23977 251641 24011 252417
rect 24091 251641 24125 252417
rect 24187 251641 24221 252417
rect 24301 251641 24335 252417
rect 24397 251641 24431 252417
rect 24511 251641 24545 252417
rect 24607 251641 24641 252417
rect 24721 251641 24755 252417
rect 24817 251641 24851 252417
rect 24931 251641 24965 252417
rect 25027 251641 25061 252417
rect 25141 251641 25175 252417
rect 25237 251641 25271 252417
rect 25351 251641 25385 252417
rect 25447 251641 25481 252417
rect 25561 251641 25595 252417
rect 25657 251641 25691 252417
rect 25771 251641 25805 252417
rect 25867 251641 25901 252417
rect 25981 251641 26015 252417
rect 26077 251641 26111 252417
rect 26191 251641 26225 252417
rect 26287 251641 26321 252417
rect 26401 251641 26435 252417
rect 26497 251641 26531 252417
rect 26611 251641 26645 252417
rect 26707 251641 26741 252417
rect 26821 251641 26855 252417
rect 26917 251641 26951 252417
rect 27031 251641 27065 252417
rect 27127 251641 27161 252417
rect 27241 251641 27275 252417
rect 27337 251641 27371 252417
rect -4049 250605 -4015 251381
rect -3953 250605 -3919 251381
rect -3839 250605 -3805 251381
rect -3743 250605 -3709 251381
rect -3629 250605 -3595 251381
rect -3533 250605 -3499 251381
rect -3419 250605 -3385 251381
rect -3323 250605 -3289 251381
rect -3209 250605 -3175 251381
rect -3113 250605 -3079 251381
rect -2999 250605 -2965 251381
rect -2903 250605 -2869 251381
rect -2789 250605 -2755 251381
rect -2693 250605 -2659 251381
rect -2579 250605 -2545 251381
rect -2483 250605 -2449 251381
rect -2369 250605 -2335 251381
rect -2273 250605 -2239 251381
rect -2159 250605 -2125 251381
rect -2063 250605 -2029 251381
rect -1949 250605 -1915 251381
rect -1853 250605 -1819 251381
rect -1739 250605 -1705 251381
rect -1643 250605 -1609 251381
rect -1529 250605 -1495 251381
rect -1433 250605 -1399 251381
rect -1319 250605 -1285 251381
rect -1223 250605 -1189 251381
rect -1109 250605 -1075 251381
rect -1013 250605 -979 251381
rect -899 250605 -865 251381
rect -803 250605 -769 251381
rect -689 250605 -655 251381
rect -593 250605 -559 251381
rect -479 250605 -445 251381
rect -383 250605 -349 251381
rect -269 250605 -235 251381
rect -173 250605 -139 251381
rect -59 250605 -25 251381
rect 37 250605 71 251381
rect 151 250605 185 251381
rect 247 250605 281 251381
rect 361 250605 395 251381
rect 457 250605 491 251381
rect 571 250605 605 251381
rect 667 250605 701 251381
rect 781 250605 815 251381
rect 877 250605 911 251381
rect 991 250605 1025 251381
rect 1087 250605 1121 251381
rect 1201 250605 1235 251381
rect 1297 250605 1331 251381
rect 1411 250605 1445 251381
rect 1507 250605 1541 251381
rect 1621 250605 1655 251381
rect 1717 250605 1751 251381
rect 1831 250605 1865 251381
rect 1927 250605 1961 251381
rect 2041 250605 2075 251381
rect 2137 250605 2171 251381
rect 2251 250605 2285 251381
rect 2347 250605 2381 251381
rect 2461 250605 2495 251381
rect 2557 250605 2591 251381
rect 2671 250605 2705 251381
rect 2767 250605 2801 251381
rect 2881 250605 2915 251381
rect 2977 250605 3011 251381
rect 3091 250605 3125 251381
rect 3187 250605 3221 251381
rect 3301 250605 3335 251381
rect 3397 250605 3431 251381
rect 3511 250605 3545 251381
rect 3607 250605 3641 251381
rect 3721 250605 3755 251381
rect 3817 250605 3851 251381
rect 3931 250605 3965 251381
rect 4027 250605 4061 251381
rect 4141 250605 4175 251381
rect 4237 250605 4271 251381
rect 4351 250605 4385 251381
rect 4447 250605 4481 251381
rect 4561 250605 4595 251381
rect 4657 250605 4691 251381
rect 4771 250605 4805 251381
rect 4867 250605 4901 251381
rect 4981 250605 5015 251381
rect 5077 250605 5111 251381
rect 5191 250605 5225 251381
rect 5287 250605 5321 251381
rect 5401 250605 5435 251381
rect 5497 250605 5531 251381
rect 5611 250605 5645 251381
rect 5707 250605 5741 251381
rect 5821 250605 5855 251381
rect 5917 250605 5951 251381
rect 6031 250605 6065 251381
rect 6127 250605 6161 251381
rect 6241 250605 6275 251381
rect 6337 250605 6371 251381
rect 6451 250605 6485 251381
rect 6547 250605 6581 251381
rect 6661 250605 6695 251381
rect 6757 250605 6791 251381
rect 6871 250605 6905 251381
rect 6967 250605 7001 251381
rect 7081 250605 7115 251381
rect 7177 250605 7211 251381
rect 7291 250605 7325 251381
rect 7387 250605 7421 251381
rect 7501 250605 7535 251381
rect 7597 250605 7631 251381
rect 7711 250605 7745 251381
rect 7807 250605 7841 251381
rect 7921 250605 7955 251381
rect 8017 250605 8051 251381
rect 8131 250605 8165 251381
rect 8227 250605 8261 251381
rect 8341 250605 8375 251381
rect 8437 250605 8471 251381
rect 8551 250605 8585 251381
rect 8647 250605 8681 251381
rect 8761 250605 8795 251381
rect 8857 250605 8891 251381
rect 8971 250605 9005 251381
rect 9067 250605 9101 251381
rect 9181 250605 9215 251381
rect 9277 250605 9311 251381
rect 9391 250605 9425 251381
rect 9487 250605 9521 251381
rect 9601 250605 9635 251381
rect 9697 250605 9731 251381
rect 9811 250605 9845 251381
rect 9907 250605 9941 251381
rect 10021 250605 10055 251381
rect 10117 250605 10151 251381
rect 10231 250605 10265 251381
rect 10327 250605 10361 251381
rect 10441 250605 10475 251381
rect 10537 250605 10571 251381
rect 10651 250605 10685 251381
rect 10747 250605 10781 251381
rect 10861 250605 10895 251381
rect 10957 250605 10991 251381
rect 11071 250605 11105 251381
rect 11167 250605 11201 251381
rect 11281 250605 11315 251381
rect 11377 250605 11411 251381
rect 11491 250605 11525 251381
rect 11587 250605 11621 251381
rect 11701 250605 11735 251381
rect 11797 250605 11831 251381
rect 11911 250605 11945 251381
rect 12007 250605 12041 251381
rect 12121 250605 12155 251381
rect 12217 250605 12251 251381
rect 12331 250605 12365 251381
rect 12427 250605 12461 251381
rect 12541 250605 12575 251381
rect 12637 250605 12671 251381
rect 12751 250605 12785 251381
rect 12847 250605 12881 251381
rect 12961 250605 12995 251381
rect 13057 250605 13091 251381
rect 13171 250605 13205 251381
rect 13267 250605 13301 251381
rect 13381 250605 13415 251381
rect 13477 250605 13511 251381
rect 13591 250605 13625 251381
rect 13687 250605 13721 251381
rect 13801 250605 13835 251381
rect 13897 250605 13931 251381
rect 14011 250605 14045 251381
rect 14107 250605 14141 251381
rect 14221 250605 14255 251381
rect 14317 250605 14351 251381
rect 14431 250605 14465 251381
rect 14527 250605 14561 251381
rect 14641 250605 14675 251381
rect 14737 250605 14771 251381
rect 14851 250605 14885 251381
rect 14947 250605 14981 251381
rect 15061 250605 15095 251381
rect 15157 250605 15191 251381
rect 15271 250605 15305 251381
rect 15367 250605 15401 251381
rect 15481 250605 15515 251381
rect 15577 250605 15611 251381
rect 15691 250605 15725 251381
rect 15787 250605 15821 251381
rect 15901 250605 15935 251381
rect 15997 250605 16031 251381
rect 16111 250605 16145 251381
rect 16207 250605 16241 251381
rect 16321 250605 16355 251381
rect 16417 250605 16451 251381
rect 16531 250605 16565 251381
rect 16627 250605 16661 251381
rect 16741 250605 16775 251381
rect 16837 250605 16871 251381
rect 16951 250605 16985 251381
rect 17047 250605 17081 251381
rect 17161 250605 17195 251381
rect 17257 250605 17291 251381
rect 17371 250605 17405 251381
rect 17467 250605 17501 251381
rect 17581 250605 17615 251381
rect 17677 250605 17711 251381
rect 17791 250605 17825 251381
rect 17887 250605 17921 251381
rect 18001 250605 18035 251381
rect 18097 250605 18131 251381
rect 18211 250605 18245 251381
rect 18307 250605 18341 251381
rect 18421 250605 18455 251381
rect 18517 250605 18551 251381
rect 18631 250605 18665 251381
rect 18727 250605 18761 251381
rect 18841 250605 18875 251381
rect 18937 250605 18971 251381
rect 19051 250605 19085 251381
rect 19147 250605 19181 251381
rect 19261 250605 19295 251381
rect 19357 250605 19391 251381
rect 19471 250605 19505 251381
rect 19567 250605 19601 251381
rect 19681 250605 19715 251381
rect 19777 250605 19811 251381
rect 19891 250605 19925 251381
rect 19987 250605 20021 251381
rect 20101 250605 20135 251381
rect 20197 250605 20231 251381
rect 20311 250605 20345 251381
rect 20407 250605 20441 251381
rect 20521 250605 20555 251381
rect 20617 250605 20651 251381
rect 20731 250605 20765 251381
rect 20827 250605 20861 251381
rect 20941 250605 20975 251381
rect 21037 250605 21071 251381
rect 21151 250605 21185 251381
rect 21247 250605 21281 251381
rect 21361 250605 21395 251381
rect 21457 250605 21491 251381
rect 21571 250605 21605 251381
rect 21667 250605 21701 251381
rect 21781 250605 21815 251381
rect 21877 250605 21911 251381
rect 21991 250605 22025 251381
rect 22087 250605 22121 251381
rect 22201 250605 22235 251381
rect 22297 250605 22331 251381
rect 22411 250605 22445 251381
rect 22507 250605 22541 251381
rect 22621 250605 22655 251381
rect 22717 250605 22751 251381
rect 22831 250605 22865 251381
rect 22927 250605 22961 251381
rect 23041 250605 23075 251381
rect 23137 250605 23171 251381
rect 23251 250605 23285 251381
rect 23347 250605 23381 251381
rect 23461 250605 23495 251381
rect 23557 250605 23591 251381
rect 23671 250605 23705 251381
rect 23767 250605 23801 251381
rect 23881 250605 23915 251381
rect 23977 250605 24011 251381
rect 24091 250605 24125 251381
rect 24187 250605 24221 251381
rect 24301 250605 24335 251381
rect 24397 250605 24431 251381
rect 24511 250605 24545 251381
rect 24607 250605 24641 251381
rect 24721 250605 24755 251381
rect 24817 250605 24851 251381
rect 24931 250605 24965 251381
rect 25027 250605 25061 251381
rect 25141 250605 25175 251381
rect 25237 250605 25271 251381
rect 25351 250605 25385 251381
rect 25447 250605 25481 251381
rect 25561 250605 25595 251381
rect 25657 250605 25691 251381
rect 25771 250605 25805 251381
rect 25867 250605 25901 251381
rect 25981 250605 26015 251381
rect 26077 250605 26111 251381
rect 26191 250605 26225 251381
rect 26287 250605 26321 251381
rect 26401 250605 26435 251381
rect 26497 250605 26531 251381
rect 26611 250605 26645 251381
rect 26707 250605 26741 251381
rect 26821 250605 26855 251381
rect 26917 250605 26951 251381
rect 27031 250605 27065 251381
rect 27127 250605 27161 251381
rect 27241 250605 27275 251381
rect 27337 250605 27371 251381
rect -4049 249569 -4015 250345
rect -3953 249569 -3919 250345
rect -3839 249569 -3805 250345
rect -3743 249569 -3709 250345
rect -3629 249569 -3595 250345
rect -3533 249569 -3499 250345
rect -3419 249569 -3385 250345
rect -3323 249569 -3289 250345
rect -3209 249569 -3175 250345
rect -3113 249569 -3079 250345
rect -2999 249569 -2965 250345
rect -2903 249569 -2869 250345
rect -2789 249569 -2755 250345
rect -2693 249569 -2659 250345
rect -2579 249569 -2545 250345
rect -2483 249569 -2449 250345
rect -2369 249569 -2335 250345
rect -2273 249569 -2239 250345
rect -2159 249569 -2125 250345
rect -2063 249569 -2029 250345
rect -1949 249569 -1915 250345
rect -1853 249569 -1819 250345
rect -1739 249569 -1705 250345
rect -1643 249569 -1609 250345
rect -1529 249569 -1495 250345
rect -1433 249569 -1399 250345
rect -1319 249569 -1285 250345
rect -1223 249569 -1189 250345
rect -1109 249569 -1075 250345
rect -1013 249569 -979 250345
rect -899 249569 -865 250345
rect -803 249569 -769 250345
rect -689 249569 -655 250345
rect -593 249569 -559 250345
rect -479 249569 -445 250345
rect -383 249569 -349 250345
rect -269 249569 -235 250345
rect -173 249569 -139 250345
rect -59 249569 -25 250345
rect 37 249569 71 250345
rect 151 249569 185 250345
rect 247 249569 281 250345
rect 361 249569 395 250345
rect 457 249569 491 250345
rect 571 249569 605 250345
rect 667 249569 701 250345
rect 781 249569 815 250345
rect 877 249569 911 250345
rect 991 249569 1025 250345
rect 1087 249569 1121 250345
rect 1201 249569 1235 250345
rect 1297 249569 1331 250345
rect 1411 249569 1445 250345
rect 1507 249569 1541 250345
rect 1621 249569 1655 250345
rect 1717 249569 1751 250345
rect 1831 249569 1865 250345
rect 1927 249569 1961 250345
rect 2041 249569 2075 250345
rect 2137 249569 2171 250345
rect 2251 249569 2285 250345
rect 2347 249569 2381 250345
rect 2461 249569 2495 250345
rect 2557 249569 2591 250345
rect 2671 249569 2705 250345
rect 2767 249569 2801 250345
rect 2881 249569 2915 250345
rect 2977 249569 3011 250345
rect 3091 249569 3125 250345
rect 3187 249569 3221 250345
rect 3301 249569 3335 250345
rect 3397 249569 3431 250345
rect 3511 249569 3545 250345
rect 3607 249569 3641 250345
rect 3721 249569 3755 250345
rect 3817 249569 3851 250345
rect 3931 249569 3965 250345
rect 4027 249569 4061 250345
rect 4141 249569 4175 250345
rect 4237 249569 4271 250345
rect 4351 249569 4385 250345
rect 4447 249569 4481 250345
rect 4561 249569 4595 250345
rect 4657 249569 4691 250345
rect 4771 249569 4805 250345
rect 4867 249569 4901 250345
rect 4981 249569 5015 250345
rect 5077 249569 5111 250345
rect 5191 249569 5225 250345
rect 5287 249569 5321 250345
rect 5401 249569 5435 250345
rect 5497 249569 5531 250345
rect 5611 249569 5645 250345
rect 5707 249569 5741 250345
rect 5821 249569 5855 250345
rect 5917 249569 5951 250345
rect 6031 249569 6065 250345
rect 6127 249569 6161 250345
rect 6241 249569 6275 250345
rect 6337 249569 6371 250345
rect 6451 249569 6485 250345
rect 6547 249569 6581 250345
rect 6661 249569 6695 250345
rect 6757 249569 6791 250345
rect 6871 249569 6905 250345
rect 6967 249569 7001 250345
rect 7081 249569 7115 250345
rect 7177 249569 7211 250345
rect 7291 249569 7325 250345
rect 7387 249569 7421 250345
rect 7501 249569 7535 250345
rect 7597 249569 7631 250345
rect 7711 249569 7745 250345
rect 7807 249569 7841 250345
rect 7921 249569 7955 250345
rect 8017 249569 8051 250345
rect 8131 249569 8165 250345
rect 8227 249569 8261 250345
rect 8341 249569 8375 250345
rect 8437 249569 8471 250345
rect 8551 249569 8585 250345
rect 8647 249569 8681 250345
rect 8761 249569 8795 250345
rect 8857 249569 8891 250345
rect 8971 249569 9005 250345
rect 9067 249569 9101 250345
rect 9181 249569 9215 250345
rect 9277 249569 9311 250345
rect 9391 249569 9425 250345
rect 9487 249569 9521 250345
rect 9601 249569 9635 250345
rect 9697 249569 9731 250345
rect 9811 249569 9845 250345
rect 9907 249569 9941 250345
rect 10021 249569 10055 250345
rect 10117 249569 10151 250345
rect 10231 249569 10265 250345
rect 10327 249569 10361 250345
rect 10441 249569 10475 250345
rect 10537 249569 10571 250345
rect 10651 249569 10685 250345
rect 10747 249569 10781 250345
rect 10861 249569 10895 250345
rect 10957 249569 10991 250345
rect 11071 249569 11105 250345
rect 11167 249569 11201 250345
rect 11281 249569 11315 250345
rect 11377 249569 11411 250345
rect 11491 249569 11525 250345
rect 11587 249569 11621 250345
rect 11701 249569 11735 250345
rect 11797 249569 11831 250345
rect 11911 249569 11945 250345
rect 12007 249569 12041 250345
rect 12121 249569 12155 250345
rect 12217 249569 12251 250345
rect 12331 249569 12365 250345
rect 12427 249569 12461 250345
rect 12541 249569 12575 250345
rect 12637 249569 12671 250345
rect 12751 249569 12785 250345
rect 12847 249569 12881 250345
rect 12961 249569 12995 250345
rect 13057 249569 13091 250345
rect 13171 249569 13205 250345
rect 13267 249569 13301 250345
rect 13381 249569 13415 250345
rect 13477 249569 13511 250345
rect 13591 249569 13625 250345
rect 13687 249569 13721 250345
rect 13801 249569 13835 250345
rect 13897 249569 13931 250345
rect 14011 249569 14045 250345
rect 14107 249569 14141 250345
rect 14221 249569 14255 250345
rect 14317 249569 14351 250345
rect 14431 249569 14465 250345
rect 14527 249569 14561 250345
rect 14641 249569 14675 250345
rect 14737 249569 14771 250345
rect 14851 249569 14885 250345
rect 14947 249569 14981 250345
rect 15061 249569 15095 250345
rect 15157 249569 15191 250345
rect 15271 249569 15305 250345
rect 15367 249569 15401 250345
rect 15481 249569 15515 250345
rect 15577 249569 15611 250345
rect 15691 249569 15725 250345
rect 15787 249569 15821 250345
rect 15901 249569 15935 250345
rect 15997 249569 16031 250345
rect 16111 249569 16145 250345
rect 16207 249569 16241 250345
rect 16321 249569 16355 250345
rect 16417 249569 16451 250345
rect 16531 249569 16565 250345
rect 16627 249569 16661 250345
rect 16741 249569 16775 250345
rect 16837 249569 16871 250345
rect 16951 249569 16985 250345
rect 17047 249569 17081 250345
rect 17161 249569 17195 250345
rect 17257 249569 17291 250345
rect 17371 249569 17405 250345
rect 17467 249569 17501 250345
rect 17581 249569 17615 250345
rect 17677 249569 17711 250345
rect 17791 249569 17825 250345
rect 17887 249569 17921 250345
rect 18001 249569 18035 250345
rect 18097 249569 18131 250345
rect 18211 249569 18245 250345
rect 18307 249569 18341 250345
rect 18421 249569 18455 250345
rect 18517 249569 18551 250345
rect 18631 249569 18665 250345
rect 18727 249569 18761 250345
rect 18841 249569 18875 250345
rect 18937 249569 18971 250345
rect 19051 249569 19085 250345
rect 19147 249569 19181 250345
rect 19261 249569 19295 250345
rect 19357 249569 19391 250345
rect 19471 249569 19505 250345
rect 19567 249569 19601 250345
rect 19681 249569 19715 250345
rect 19777 249569 19811 250345
rect 19891 249569 19925 250345
rect 19987 249569 20021 250345
rect 20101 249569 20135 250345
rect 20197 249569 20231 250345
rect 20311 249569 20345 250345
rect 20407 249569 20441 250345
rect 20521 249569 20555 250345
rect 20617 249569 20651 250345
rect 20731 249569 20765 250345
rect 20827 249569 20861 250345
rect 20941 249569 20975 250345
rect 21037 249569 21071 250345
rect 21151 249569 21185 250345
rect 21247 249569 21281 250345
rect 21361 249569 21395 250345
rect 21457 249569 21491 250345
rect 21571 249569 21605 250345
rect 21667 249569 21701 250345
rect 21781 249569 21815 250345
rect 21877 249569 21911 250345
rect 21991 249569 22025 250345
rect 22087 249569 22121 250345
rect 22201 249569 22235 250345
rect 22297 249569 22331 250345
rect 22411 249569 22445 250345
rect 22507 249569 22541 250345
rect 22621 249569 22655 250345
rect 22717 249569 22751 250345
rect 22831 249569 22865 250345
rect 22927 249569 22961 250345
rect 23041 249569 23075 250345
rect 23137 249569 23171 250345
rect 23251 249569 23285 250345
rect 23347 249569 23381 250345
rect 23461 249569 23495 250345
rect 23557 249569 23591 250345
rect 23671 249569 23705 250345
rect 23767 249569 23801 250345
rect 23881 249569 23915 250345
rect 23977 249569 24011 250345
rect 24091 249569 24125 250345
rect 24187 249569 24221 250345
rect 24301 249569 24335 250345
rect 24397 249569 24431 250345
rect 24511 249569 24545 250345
rect 24607 249569 24641 250345
rect 24721 249569 24755 250345
rect 24817 249569 24851 250345
rect 24931 249569 24965 250345
rect 25027 249569 25061 250345
rect 25141 249569 25175 250345
rect 25237 249569 25271 250345
rect 25351 249569 25385 250345
rect 25447 249569 25481 250345
rect 25561 249569 25595 250345
rect 25657 249569 25691 250345
rect 25771 249569 25805 250345
rect 25867 249569 25901 250345
rect 25981 249569 26015 250345
rect 26077 249569 26111 250345
rect 26191 249569 26225 250345
rect 26287 249569 26321 250345
rect 26401 249569 26435 250345
rect 26497 249569 26531 250345
rect 26611 249569 26645 250345
rect 26707 249569 26741 250345
rect 26821 249569 26855 250345
rect 26917 249569 26951 250345
rect 27031 249569 27065 250345
rect 27127 249569 27161 250345
rect 27241 249569 27275 250345
rect 27337 249569 27371 250345
rect -4049 248404 -4015 249180
rect -3953 248404 -3919 249180
rect -3839 248404 -3805 249180
rect -3743 248404 -3709 249180
rect -3629 248404 -3595 249180
rect -3533 248404 -3499 249180
rect -3419 248404 -3385 249180
rect -3323 248404 -3289 249180
rect -3209 248404 -3175 249180
rect -3113 248404 -3079 249180
rect -2999 248404 -2965 249180
rect -2903 248404 -2869 249180
rect -2789 248404 -2755 249180
rect -2693 248404 -2659 249180
rect -2579 248404 -2545 249180
rect -2483 248404 -2449 249180
rect -2369 248404 -2335 249180
rect -2273 248404 -2239 249180
rect -2159 248404 -2125 249180
rect -2063 248404 -2029 249180
rect -1949 248404 -1915 249180
rect -1853 248404 -1819 249180
rect -1739 248404 -1705 249180
rect -1643 248404 -1609 249180
rect -1529 248404 -1495 249180
rect -1433 248404 -1399 249180
rect -1319 248404 -1285 249180
rect -1223 248404 -1189 249180
rect -1109 248404 -1075 249180
rect -1013 248404 -979 249180
rect -899 248404 -865 249180
rect -803 248404 -769 249180
rect -689 248404 -655 249180
rect -593 248404 -559 249180
rect -479 248404 -445 249180
rect -383 248404 -349 249180
rect -269 248404 -235 249180
rect -173 248404 -139 249180
rect -59 248404 -25 249180
rect 37 248404 71 249180
rect 151 248404 185 249180
rect 247 248404 281 249180
rect 361 248404 395 249180
rect 457 248404 491 249180
rect 571 248404 605 249180
rect 667 248404 701 249180
rect 781 248404 815 249180
rect 877 248404 911 249180
rect 991 248404 1025 249180
rect 1087 248404 1121 249180
rect 1201 248404 1235 249180
rect 1297 248404 1331 249180
rect 1411 248404 1445 249180
rect 1507 248404 1541 249180
rect 1621 248404 1655 249180
rect 1717 248404 1751 249180
rect 1831 248404 1865 249180
rect 1927 248404 1961 249180
rect 2041 248404 2075 249180
rect 2137 248404 2171 249180
rect 2251 248404 2285 249180
rect 2347 248404 2381 249180
rect 2461 248404 2495 249180
rect 2557 248404 2591 249180
rect 2671 248404 2705 249180
rect 2767 248404 2801 249180
rect 2881 248404 2915 249180
rect 2977 248404 3011 249180
rect 3091 248404 3125 249180
rect 3187 248404 3221 249180
rect 3301 248404 3335 249180
rect 3397 248404 3431 249180
rect 3511 248404 3545 249180
rect 3607 248404 3641 249180
rect 3721 248404 3755 249180
rect 3817 248404 3851 249180
rect 3931 248404 3965 249180
rect 4027 248404 4061 249180
rect 4141 248404 4175 249180
rect 4237 248404 4271 249180
rect 4351 248404 4385 249180
rect 4447 248404 4481 249180
rect 4561 248404 4595 249180
rect 4657 248404 4691 249180
rect 4771 248404 4805 249180
rect 4867 248404 4901 249180
rect 4981 248404 5015 249180
rect 5077 248404 5111 249180
rect 5191 248404 5225 249180
rect 5287 248404 5321 249180
rect 5401 248404 5435 249180
rect 5497 248404 5531 249180
rect 5611 248404 5645 249180
rect 5707 248404 5741 249180
rect 5821 248404 5855 249180
rect 5917 248404 5951 249180
rect 6031 248404 6065 249180
rect 6127 248404 6161 249180
rect 6241 248404 6275 249180
rect 6337 248404 6371 249180
rect 6451 248404 6485 249180
rect 6547 248404 6581 249180
rect 6661 248404 6695 249180
rect 6757 248404 6791 249180
rect 6871 248404 6905 249180
rect 6967 248404 7001 249180
rect 7081 248404 7115 249180
rect 7177 248404 7211 249180
rect 7291 248404 7325 249180
rect 7387 248404 7421 249180
rect 7501 248404 7535 249180
rect 7597 248404 7631 249180
rect 7711 248404 7745 249180
rect 7807 248404 7841 249180
rect 7921 248404 7955 249180
rect 8017 248404 8051 249180
rect 8131 248404 8165 249180
rect 8227 248404 8261 249180
rect 8341 248404 8375 249180
rect 8437 248404 8471 249180
rect 8551 248404 8585 249180
rect 8647 248404 8681 249180
rect 8761 248404 8795 249180
rect 8857 248404 8891 249180
rect 8971 248404 9005 249180
rect 9067 248404 9101 249180
rect 9181 248404 9215 249180
rect 9277 248404 9311 249180
rect 9391 248404 9425 249180
rect 9487 248404 9521 249180
rect 9601 248404 9635 249180
rect 9697 248404 9731 249180
rect 9811 248404 9845 249180
rect 9907 248404 9941 249180
rect 10021 248404 10055 249180
rect 10117 248404 10151 249180
rect 10231 248404 10265 249180
rect 10327 248404 10361 249180
rect 10441 248404 10475 249180
rect 10537 248404 10571 249180
rect 10651 248404 10685 249180
rect 10747 248404 10781 249180
rect 10861 248404 10895 249180
rect 10957 248404 10991 249180
rect 11071 248404 11105 249180
rect 11167 248404 11201 249180
rect 11281 248404 11315 249180
rect 11377 248404 11411 249180
rect 11491 248404 11525 249180
rect 11587 248404 11621 249180
rect 11701 248404 11735 249180
rect 11797 248404 11831 249180
rect 11911 248404 11945 249180
rect 12007 248404 12041 249180
rect 12121 248404 12155 249180
rect 12217 248404 12251 249180
rect 12331 248404 12365 249180
rect 12427 248404 12461 249180
rect 12541 248404 12575 249180
rect 12637 248404 12671 249180
rect 12751 248404 12785 249180
rect 12847 248404 12881 249180
rect 12961 248404 12995 249180
rect 13057 248404 13091 249180
rect 13171 248404 13205 249180
rect 13267 248404 13301 249180
rect 13381 248404 13415 249180
rect 13477 248404 13511 249180
rect 13591 248404 13625 249180
rect 13687 248404 13721 249180
rect 13801 248404 13835 249180
rect 13897 248404 13931 249180
rect 14011 248404 14045 249180
rect 14107 248404 14141 249180
rect 14221 248404 14255 249180
rect 14317 248404 14351 249180
rect 14431 248404 14465 249180
rect 14527 248404 14561 249180
rect 14641 248404 14675 249180
rect 14737 248404 14771 249180
rect 14851 248404 14885 249180
rect 14947 248404 14981 249180
rect 15061 248404 15095 249180
rect 15157 248404 15191 249180
rect 15271 248404 15305 249180
rect 15367 248404 15401 249180
rect 15481 248404 15515 249180
rect 15577 248404 15611 249180
rect 15691 248404 15725 249180
rect 15787 248404 15821 249180
rect 15901 248404 15935 249180
rect 15997 248404 16031 249180
rect 16111 248404 16145 249180
rect 16207 248404 16241 249180
rect 16321 248404 16355 249180
rect 16417 248404 16451 249180
rect 16531 248404 16565 249180
rect 16627 248404 16661 249180
rect 16741 248404 16775 249180
rect 16837 248404 16871 249180
rect 16951 248404 16985 249180
rect 17047 248404 17081 249180
rect 17161 248404 17195 249180
rect 17257 248404 17291 249180
rect 17371 248404 17405 249180
rect 17467 248404 17501 249180
rect 17581 248404 17615 249180
rect 17677 248404 17711 249180
rect 17791 248404 17825 249180
rect 17887 248404 17921 249180
rect 18001 248404 18035 249180
rect 18097 248404 18131 249180
rect 18211 248404 18245 249180
rect 18307 248404 18341 249180
rect 18421 248404 18455 249180
rect 18517 248404 18551 249180
rect 18631 248404 18665 249180
rect 18727 248404 18761 249180
rect 18841 248404 18875 249180
rect 18937 248404 18971 249180
rect 19051 248404 19085 249180
rect 19147 248404 19181 249180
rect 19261 248404 19295 249180
rect 19357 248404 19391 249180
rect 19471 248404 19505 249180
rect 19567 248404 19601 249180
rect 19681 248404 19715 249180
rect 19777 248404 19811 249180
rect 19891 248404 19925 249180
rect 19987 248404 20021 249180
rect 20101 248404 20135 249180
rect 20197 248404 20231 249180
rect 20311 248404 20345 249180
rect 20407 248404 20441 249180
rect 20521 248404 20555 249180
rect 20617 248404 20651 249180
rect 20731 248404 20765 249180
rect 20827 248404 20861 249180
rect 20941 248404 20975 249180
rect 21037 248404 21071 249180
rect 21151 248404 21185 249180
rect 21247 248404 21281 249180
rect 21361 248404 21395 249180
rect 21457 248404 21491 249180
rect 21571 248404 21605 249180
rect 21667 248404 21701 249180
rect 21781 248404 21815 249180
rect 21877 248404 21911 249180
rect 21991 248404 22025 249180
rect 22087 248404 22121 249180
rect 22201 248404 22235 249180
rect 22297 248404 22331 249180
rect 22411 248404 22445 249180
rect 22507 248404 22541 249180
rect 22621 248404 22655 249180
rect 22717 248404 22751 249180
rect 22831 248404 22865 249180
rect 22927 248404 22961 249180
rect 23041 248404 23075 249180
rect 23137 248404 23171 249180
rect 23251 248404 23285 249180
rect 23347 248404 23381 249180
rect 23461 248404 23495 249180
rect 23557 248404 23591 249180
rect 23671 248404 23705 249180
rect 23767 248404 23801 249180
rect 23881 248404 23915 249180
rect 23977 248404 24011 249180
rect 24091 248404 24125 249180
rect 24187 248404 24221 249180
rect 24301 248404 24335 249180
rect 24397 248404 24431 249180
rect 24511 248404 24545 249180
rect 24607 248404 24641 249180
rect 24721 248404 24755 249180
rect 24817 248404 24851 249180
rect 24931 248404 24965 249180
rect 25027 248404 25061 249180
rect 25141 248404 25175 249180
rect 25237 248404 25271 249180
rect 25351 248404 25385 249180
rect 25447 248404 25481 249180
rect 25561 248404 25595 249180
rect 25657 248404 25691 249180
rect 25771 248404 25805 249180
rect 25867 248404 25901 249180
rect 25981 248404 26015 249180
rect 26077 248404 26111 249180
rect 26191 248404 26225 249180
rect 26287 248404 26321 249180
rect 26401 248404 26435 249180
rect 26497 248404 26531 249180
rect 26611 248404 26645 249180
rect 26707 248404 26741 249180
rect 26821 248404 26855 249180
rect 26917 248404 26951 249180
rect 27031 248404 27065 249180
rect 27127 248404 27161 249180
rect 27241 248404 27275 249180
rect 27337 248404 27371 249180
rect -4049 247368 -4015 248144
rect -3953 247368 -3919 248144
rect -3839 247368 -3805 248144
rect -3743 247368 -3709 248144
rect -3629 247368 -3595 248144
rect -3533 247368 -3499 248144
rect -3419 247368 -3385 248144
rect -3323 247368 -3289 248144
rect -3209 247368 -3175 248144
rect -3113 247368 -3079 248144
rect -2999 247368 -2965 248144
rect -2903 247368 -2869 248144
rect -2789 247368 -2755 248144
rect -2693 247368 -2659 248144
rect -2579 247368 -2545 248144
rect -2483 247368 -2449 248144
rect -2369 247368 -2335 248144
rect -2273 247368 -2239 248144
rect -2159 247368 -2125 248144
rect -2063 247368 -2029 248144
rect -1949 247368 -1915 248144
rect -1853 247368 -1819 248144
rect -1739 247368 -1705 248144
rect -1643 247368 -1609 248144
rect -1529 247368 -1495 248144
rect -1433 247368 -1399 248144
rect -1319 247368 -1285 248144
rect -1223 247368 -1189 248144
rect -1109 247368 -1075 248144
rect -1013 247368 -979 248144
rect -899 247368 -865 248144
rect -803 247368 -769 248144
rect -689 247368 -655 248144
rect -593 247368 -559 248144
rect -479 247368 -445 248144
rect -383 247368 -349 248144
rect -269 247368 -235 248144
rect -173 247368 -139 248144
rect -59 247368 -25 248144
rect 37 247368 71 248144
rect 151 247368 185 248144
rect 247 247368 281 248144
rect 361 247368 395 248144
rect 457 247368 491 248144
rect 571 247368 605 248144
rect 667 247368 701 248144
rect 781 247368 815 248144
rect 877 247368 911 248144
rect 991 247368 1025 248144
rect 1087 247368 1121 248144
rect 1201 247368 1235 248144
rect 1297 247368 1331 248144
rect 1411 247368 1445 248144
rect 1507 247368 1541 248144
rect 1621 247368 1655 248144
rect 1717 247368 1751 248144
rect 1831 247368 1865 248144
rect 1927 247368 1961 248144
rect 2041 247368 2075 248144
rect 2137 247368 2171 248144
rect 2251 247368 2285 248144
rect 2347 247368 2381 248144
rect 2461 247368 2495 248144
rect 2557 247368 2591 248144
rect 2671 247368 2705 248144
rect 2767 247368 2801 248144
rect 2881 247368 2915 248144
rect 2977 247368 3011 248144
rect 3091 247368 3125 248144
rect 3187 247368 3221 248144
rect 3301 247368 3335 248144
rect 3397 247368 3431 248144
rect 3511 247368 3545 248144
rect 3607 247368 3641 248144
rect 3721 247368 3755 248144
rect 3817 247368 3851 248144
rect 3931 247368 3965 248144
rect 4027 247368 4061 248144
rect 4141 247368 4175 248144
rect 4237 247368 4271 248144
rect 4351 247368 4385 248144
rect 4447 247368 4481 248144
rect 4561 247368 4595 248144
rect 4657 247368 4691 248144
rect 4771 247368 4805 248144
rect 4867 247368 4901 248144
rect 4981 247368 5015 248144
rect 5077 247368 5111 248144
rect 5191 247368 5225 248144
rect 5287 247368 5321 248144
rect 5401 247368 5435 248144
rect 5497 247368 5531 248144
rect 5611 247368 5645 248144
rect 5707 247368 5741 248144
rect 5821 247368 5855 248144
rect 5917 247368 5951 248144
rect 6031 247368 6065 248144
rect 6127 247368 6161 248144
rect 6241 247368 6275 248144
rect 6337 247368 6371 248144
rect 6451 247368 6485 248144
rect 6547 247368 6581 248144
rect 6661 247368 6695 248144
rect 6757 247368 6791 248144
rect 6871 247368 6905 248144
rect 6967 247368 7001 248144
rect 7081 247368 7115 248144
rect 7177 247368 7211 248144
rect 7291 247368 7325 248144
rect 7387 247368 7421 248144
rect 7501 247368 7535 248144
rect 7597 247368 7631 248144
rect 7711 247368 7745 248144
rect 7807 247368 7841 248144
rect 7921 247368 7955 248144
rect 8017 247368 8051 248144
rect 8131 247368 8165 248144
rect 8227 247368 8261 248144
rect 8341 247368 8375 248144
rect 8437 247368 8471 248144
rect 8551 247368 8585 248144
rect 8647 247368 8681 248144
rect 8761 247368 8795 248144
rect 8857 247368 8891 248144
rect 8971 247368 9005 248144
rect 9067 247368 9101 248144
rect 9181 247368 9215 248144
rect 9277 247368 9311 248144
rect 9391 247368 9425 248144
rect 9487 247368 9521 248144
rect 9601 247368 9635 248144
rect 9697 247368 9731 248144
rect 9811 247368 9845 248144
rect 9907 247368 9941 248144
rect 10021 247368 10055 248144
rect 10117 247368 10151 248144
rect 10231 247368 10265 248144
rect 10327 247368 10361 248144
rect 10441 247368 10475 248144
rect 10537 247368 10571 248144
rect 10651 247368 10685 248144
rect 10747 247368 10781 248144
rect 10861 247368 10895 248144
rect 10957 247368 10991 248144
rect 11071 247368 11105 248144
rect 11167 247368 11201 248144
rect 11281 247368 11315 248144
rect 11377 247368 11411 248144
rect 11491 247368 11525 248144
rect 11587 247368 11621 248144
rect 11701 247368 11735 248144
rect 11797 247368 11831 248144
rect 11911 247368 11945 248144
rect 12007 247368 12041 248144
rect 12121 247368 12155 248144
rect 12217 247368 12251 248144
rect 12331 247368 12365 248144
rect 12427 247368 12461 248144
rect 12541 247368 12575 248144
rect 12637 247368 12671 248144
rect 12751 247368 12785 248144
rect 12847 247368 12881 248144
rect 12961 247368 12995 248144
rect 13057 247368 13091 248144
rect 13171 247368 13205 248144
rect 13267 247368 13301 248144
rect 13381 247368 13415 248144
rect 13477 247368 13511 248144
rect 13591 247368 13625 248144
rect 13687 247368 13721 248144
rect 13801 247368 13835 248144
rect 13897 247368 13931 248144
rect 14011 247368 14045 248144
rect 14107 247368 14141 248144
rect 14221 247368 14255 248144
rect 14317 247368 14351 248144
rect 14431 247368 14465 248144
rect 14527 247368 14561 248144
rect 14641 247368 14675 248144
rect 14737 247368 14771 248144
rect 14851 247368 14885 248144
rect 14947 247368 14981 248144
rect 15061 247368 15095 248144
rect 15157 247368 15191 248144
rect 15271 247368 15305 248144
rect 15367 247368 15401 248144
rect 15481 247368 15515 248144
rect 15577 247368 15611 248144
rect 15691 247368 15725 248144
rect 15787 247368 15821 248144
rect 15901 247368 15935 248144
rect 15997 247368 16031 248144
rect 16111 247368 16145 248144
rect 16207 247368 16241 248144
rect 16321 247368 16355 248144
rect 16417 247368 16451 248144
rect 16531 247368 16565 248144
rect 16627 247368 16661 248144
rect 16741 247368 16775 248144
rect 16837 247368 16871 248144
rect 16951 247368 16985 248144
rect 17047 247368 17081 248144
rect 17161 247368 17195 248144
rect 17257 247368 17291 248144
rect 17371 247368 17405 248144
rect 17467 247368 17501 248144
rect 17581 247368 17615 248144
rect 17677 247368 17711 248144
rect 17791 247368 17825 248144
rect 17887 247368 17921 248144
rect 18001 247368 18035 248144
rect 18097 247368 18131 248144
rect 18211 247368 18245 248144
rect 18307 247368 18341 248144
rect 18421 247368 18455 248144
rect 18517 247368 18551 248144
rect 18631 247368 18665 248144
rect 18727 247368 18761 248144
rect 18841 247368 18875 248144
rect 18937 247368 18971 248144
rect 19051 247368 19085 248144
rect 19147 247368 19181 248144
rect 19261 247368 19295 248144
rect 19357 247368 19391 248144
rect 19471 247368 19505 248144
rect 19567 247368 19601 248144
rect 19681 247368 19715 248144
rect 19777 247368 19811 248144
rect 19891 247368 19925 248144
rect 19987 247368 20021 248144
rect 20101 247368 20135 248144
rect 20197 247368 20231 248144
rect 20311 247368 20345 248144
rect 20407 247368 20441 248144
rect 20521 247368 20555 248144
rect 20617 247368 20651 248144
rect 20731 247368 20765 248144
rect 20827 247368 20861 248144
rect 20941 247368 20975 248144
rect 21037 247368 21071 248144
rect 21151 247368 21185 248144
rect 21247 247368 21281 248144
rect 21361 247368 21395 248144
rect 21457 247368 21491 248144
rect 21571 247368 21605 248144
rect 21667 247368 21701 248144
rect 21781 247368 21815 248144
rect 21877 247368 21911 248144
rect 21991 247368 22025 248144
rect 22087 247368 22121 248144
rect 22201 247368 22235 248144
rect 22297 247368 22331 248144
rect 22411 247368 22445 248144
rect 22507 247368 22541 248144
rect 22621 247368 22655 248144
rect 22717 247368 22751 248144
rect 22831 247368 22865 248144
rect 22927 247368 22961 248144
rect 23041 247368 23075 248144
rect 23137 247368 23171 248144
rect 23251 247368 23285 248144
rect 23347 247368 23381 248144
rect 23461 247368 23495 248144
rect 23557 247368 23591 248144
rect 23671 247368 23705 248144
rect 23767 247368 23801 248144
rect 23881 247368 23915 248144
rect 23977 247368 24011 248144
rect 24091 247368 24125 248144
rect 24187 247368 24221 248144
rect 24301 247368 24335 248144
rect 24397 247368 24431 248144
rect 24511 247368 24545 248144
rect 24607 247368 24641 248144
rect 24721 247368 24755 248144
rect 24817 247368 24851 248144
rect 24931 247368 24965 248144
rect 25027 247368 25061 248144
rect 25141 247368 25175 248144
rect 25237 247368 25271 248144
rect 25351 247368 25385 248144
rect 25447 247368 25481 248144
rect 25561 247368 25595 248144
rect 25657 247368 25691 248144
rect 25771 247368 25805 248144
rect 25867 247368 25901 248144
rect 25981 247368 26015 248144
rect 26077 247368 26111 248144
rect 26191 247368 26225 248144
rect 26287 247368 26321 248144
rect 26401 247368 26435 248144
rect 26497 247368 26531 248144
rect 26611 247368 26645 248144
rect 26707 247368 26741 248144
rect 26821 247368 26855 248144
rect 26917 247368 26951 248144
rect 27031 247368 27065 248144
rect 27127 247368 27161 248144
rect 27241 247368 27275 248144
rect 27337 247368 27371 248144
rect -4049 246332 -4015 247108
rect -3953 246332 -3919 247108
rect -3839 246332 -3805 247108
rect -3743 246332 -3709 247108
rect -3629 246332 -3595 247108
rect -3533 246332 -3499 247108
rect -3419 246332 -3385 247108
rect -3323 246332 -3289 247108
rect -3209 246332 -3175 247108
rect -3113 246332 -3079 247108
rect -2999 246332 -2965 247108
rect -2903 246332 -2869 247108
rect -2789 246332 -2755 247108
rect -2693 246332 -2659 247108
rect -2579 246332 -2545 247108
rect -2483 246332 -2449 247108
rect -2369 246332 -2335 247108
rect -2273 246332 -2239 247108
rect -2159 246332 -2125 247108
rect -2063 246332 -2029 247108
rect -1949 246332 -1915 247108
rect -1853 246332 -1819 247108
rect -1739 246332 -1705 247108
rect -1643 246332 -1609 247108
rect -1529 246332 -1495 247108
rect -1433 246332 -1399 247108
rect -1319 246332 -1285 247108
rect -1223 246332 -1189 247108
rect -1109 246332 -1075 247108
rect -1013 246332 -979 247108
rect -899 246332 -865 247108
rect -803 246332 -769 247108
rect -689 246332 -655 247108
rect -593 246332 -559 247108
rect -479 246332 -445 247108
rect -383 246332 -349 247108
rect -269 246332 -235 247108
rect -173 246332 -139 247108
rect -59 246332 -25 247108
rect 37 246332 71 247108
rect 151 246332 185 247108
rect 247 246332 281 247108
rect 361 246332 395 247108
rect 457 246332 491 247108
rect 571 246332 605 247108
rect 667 246332 701 247108
rect 781 246332 815 247108
rect 877 246332 911 247108
rect 991 246332 1025 247108
rect 1087 246332 1121 247108
rect 1201 246332 1235 247108
rect 1297 246332 1331 247108
rect 1411 246332 1445 247108
rect 1507 246332 1541 247108
rect 1621 246332 1655 247108
rect 1717 246332 1751 247108
rect 1831 246332 1865 247108
rect 1927 246332 1961 247108
rect 2041 246332 2075 247108
rect 2137 246332 2171 247108
rect 2251 246332 2285 247108
rect 2347 246332 2381 247108
rect 2461 246332 2495 247108
rect 2557 246332 2591 247108
rect 2671 246332 2705 247108
rect 2767 246332 2801 247108
rect 2881 246332 2915 247108
rect 2977 246332 3011 247108
rect 3091 246332 3125 247108
rect 3187 246332 3221 247108
rect 3301 246332 3335 247108
rect 3397 246332 3431 247108
rect 3511 246332 3545 247108
rect 3607 246332 3641 247108
rect 3721 246332 3755 247108
rect 3817 246332 3851 247108
rect 3931 246332 3965 247108
rect 4027 246332 4061 247108
rect 4141 246332 4175 247108
rect 4237 246332 4271 247108
rect 4351 246332 4385 247108
rect 4447 246332 4481 247108
rect 4561 246332 4595 247108
rect 4657 246332 4691 247108
rect 4771 246332 4805 247108
rect 4867 246332 4901 247108
rect 4981 246332 5015 247108
rect 5077 246332 5111 247108
rect 5191 246332 5225 247108
rect 5287 246332 5321 247108
rect 5401 246332 5435 247108
rect 5497 246332 5531 247108
rect 5611 246332 5645 247108
rect 5707 246332 5741 247108
rect 5821 246332 5855 247108
rect 5917 246332 5951 247108
rect 6031 246332 6065 247108
rect 6127 246332 6161 247108
rect 6241 246332 6275 247108
rect 6337 246332 6371 247108
rect 6451 246332 6485 247108
rect 6547 246332 6581 247108
rect 6661 246332 6695 247108
rect 6757 246332 6791 247108
rect 6871 246332 6905 247108
rect 6967 246332 7001 247108
rect 7081 246332 7115 247108
rect 7177 246332 7211 247108
rect 7291 246332 7325 247108
rect 7387 246332 7421 247108
rect 7501 246332 7535 247108
rect 7597 246332 7631 247108
rect 7711 246332 7745 247108
rect 7807 246332 7841 247108
rect 7921 246332 7955 247108
rect 8017 246332 8051 247108
rect 8131 246332 8165 247108
rect 8227 246332 8261 247108
rect 8341 246332 8375 247108
rect 8437 246332 8471 247108
rect 8551 246332 8585 247108
rect 8647 246332 8681 247108
rect 8761 246332 8795 247108
rect 8857 246332 8891 247108
rect 8971 246332 9005 247108
rect 9067 246332 9101 247108
rect 9181 246332 9215 247108
rect 9277 246332 9311 247108
rect 9391 246332 9425 247108
rect 9487 246332 9521 247108
rect 9601 246332 9635 247108
rect 9697 246332 9731 247108
rect 9811 246332 9845 247108
rect 9907 246332 9941 247108
rect 10021 246332 10055 247108
rect 10117 246332 10151 247108
rect 10231 246332 10265 247108
rect 10327 246332 10361 247108
rect 10441 246332 10475 247108
rect 10537 246332 10571 247108
rect 10651 246332 10685 247108
rect 10747 246332 10781 247108
rect 10861 246332 10895 247108
rect 10957 246332 10991 247108
rect 11071 246332 11105 247108
rect 11167 246332 11201 247108
rect 11281 246332 11315 247108
rect 11377 246332 11411 247108
rect 11491 246332 11525 247108
rect 11587 246332 11621 247108
rect 11701 246332 11735 247108
rect 11797 246332 11831 247108
rect 11911 246332 11945 247108
rect 12007 246332 12041 247108
rect 12121 246332 12155 247108
rect 12217 246332 12251 247108
rect 12331 246332 12365 247108
rect 12427 246332 12461 247108
rect 12541 246332 12575 247108
rect 12637 246332 12671 247108
rect 12751 246332 12785 247108
rect 12847 246332 12881 247108
rect 12961 246332 12995 247108
rect 13057 246332 13091 247108
rect 13171 246332 13205 247108
rect 13267 246332 13301 247108
rect 13381 246332 13415 247108
rect 13477 246332 13511 247108
rect 13591 246332 13625 247108
rect 13687 246332 13721 247108
rect 13801 246332 13835 247108
rect 13897 246332 13931 247108
rect 14011 246332 14045 247108
rect 14107 246332 14141 247108
rect 14221 246332 14255 247108
rect 14317 246332 14351 247108
rect 14431 246332 14465 247108
rect 14527 246332 14561 247108
rect 14641 246332 14675 247108
rect 14737 246332 14771 247108
rect 14851 246332 14885 247108
rect 14947 246332 14981 247108
rect 15061 246332 15095 247108
rect 15157 246332 15191 247108
rect 15271 246332 15305 247108
rect 15367 246332 15401 247108
rect 15481 246332 15515 247108
rect 15577 246332 15611 247108
rect 15691 246332 15725 247108
rect 15787 246332 15821 247108
rect 15901 246332 15935 247108
rect 15997 246332 16031 247108
rect 16111 246332 16145 247108
rect 16207 246332 16241 247108
rect 16321 246332 16355 247108
rect 16417 246332 16451 247108
rect 16531 246332 16565 247108
rect 16627 246332 16661 247108
rect 16741 246332 16775 247108
rect 16837 246332 16871 247108
rect 16951 246332 16985 247108
rect 17047 246332 17081 247108
rect 17161 246332 17195 247108
rect 17257 246332 17291 247108
rect 17371 246332 17405 247108
rect 17467 246332 17501 247108
rect 17581 246332 17615 247108
rect 17677 246332 17711 247108
rect 17791 246332 17825 247108
rect 17887 246332 17921 247108
rect 18001 246332 18035 247108
rect 18097 246332 18131 247108
rect 18211 246332 18245 247108
rect 18307 246332 18341 247108
rect 18421 246332 18455 247108
rect 18517 246332 18551 247108
rect 18631 246332 18665 247108
rect 18727 246332 18761 247108
rect 18841 246332 18875 247108
rect 18937 246332 18971 247108
rect 19051 246332 19085 247108
rect 19147 246332 19181 247108
rect 19261 246332 19295 247108
rect 19357 246332 19391 247108
rect 19471 246332 19505 247108
rect 19567 246332 19601 247108
rect 19681 246332 19715 247108
rect 19777 246332 19811 247108
rect 19891 246332 19925 247108
rect 19987 246332 20021 247108
rect 20101 246332 20135 247108
rect 20197 246332 20231 247108
rect 20311 246332 20345 247108
rect 20407 246332 20441 247108
rect 20521 246332 20555 247108
rect 20617 246332 20651 247108
rect 20731 246332 20765 247108
rect 20827 246332 20861 247108
rect 20941 246332 20975 247108
rect 21037 246332 21071 247108
rect 21151 246332 21185 247108
rect 21247 246332 21281 247108
rect 21361 246332 21395 247108
rect 21457 246332 21491 247108
rect 21571 246332 21605 247108
rect 21667 246332 21701 247108
rect 21781 246332 21815 247108
rect 21877 246332 21911 247108
rect 21991 246332 22025 247108
rect 22087 246332 22121 247108
rect 22201 246332 22235 247108
rect 22297 246332 22331 247108
rect 22411 246332 22445 247108
rect 22507 246332 22541 247108
rect 22621 246332 22655 247108
rect 22717 246332 22751 247108
rect 22831 246332 22865 247108
rect 22927 246332 22961 247108
rect 23041 246332 23075 247108
rect 23137 246332 23171 247108
rect 23251 246332 23285 247108
rect 23347 246332 23381 247108
rect 23461 246332 23495 247108
rect 23557 246332 23591 247108
rect 23671 246332 23705 247108
rect 23767 246332 23801 247108
rect 23881 246332 23915 247108
rect 23977 246332 24011 247108
rect 24091 246332 24125 247108
rect 24187 246332 24221 247108
rect 24301 246332 24335 247108
rect 24397 246332 24431 247108
rect 24511 246332 24545 247108
rect 24607 246332 24641 247108
rect 24721 246332 24755 247108
rect 24817 246332 24851 247108
rect 24931 246332 24965 247108
rect 25027 246332 25061 247108
rect 25141 246332 25175 247108
rect 25237 246332 25271 247108
rect 25351 246332 25385 247108
rect 25447 246332 25481 247108
rect 25561 246332 25595 247108
rect 25657 246332 25691 247108
rect 25771 246332 25805 247108
rect 25867 246332 25901 247108
rect 25981 246332 26015 247108
rect 26077 246332 26111 247108
rect 26191 246332 26225 247108
rect 26287 246332 26321 247108
rect 26401 246332 26435 247108
rect 26497 246332 26531 247108
rect 26611 246332 26645 247108
rect 26707 246332 26741 247108
rect 26821 246332 26855 247108
rect 26917 246332 26951 247108
rect 27031 246332 27065 247108
rect 27127 246332 27161 247108
rect 27241 246332 27275 247108
rect 27337 246332 27371 247108
rect -4049 245296 -4015 246072
rect -3953 245296 -3919 246072
rect -3839 245296 -3805 246072
rect -3743 245296 -3709 246072
rect -3629 245296 -3595 246072
rect -3533 245296 -3499 246072
rect -3419 245296 -3385 246072
rect -3323 245296 -3289 246072
rect -3209 245296 -3175 246072
rect -3113 245296 -3079 246072
rect -2999 245296 -2965 246072
rect -2903 245296 -2869 246072
rect -2789 245296 -2755 246072
rect -2693 245296 -2659 246072
rect -2579 245296 -2545 246072
rect -2483 245296 -2449 246072
rect -2369 245296 -2335 246072
rect -2273 245296 -2239 246072
rect -2159 245296 -2125 246072
rect -2063 245296 -2029 246072
rect -1949 245296 -1915 246072
rect -1853 245296 -1819 246072
rect -1739 245296 -1705 246072
rect -1643 245296 -1609 246072
rect -1529 245296 -1495 246072
rect -1433 245296 -1399 246072
rect -1319 245296 -1285 246072
rect -1223 245296 -1189 246072
rect -1109 245296 -1075 246072
rect -1013 245296 -979 246072
rect -899 245296 -865 246072
rect -803 245296 -769 246072
rect -689 245296 -655 246072
rect -593 245296 -559 246072
rect -479 245296 -445 246072
rect -383 245296 -349 246072
rect -269 245296 -235 246072
rect -173 245296 -139 246072
rect -59 245296 -25 246072
rect 37 245296 71 246072
rect 151 245296 185 246072
rect 247 245296 281 246072
rect 361 245296 395 246072
rect 457 245296 491 246072
rect 571 245296 605 246072
rect 667 245296 701 246072
rect 781 245296 815 246072
rect 877 245296 911 246072
rect 991 245296 1025 246072
rect 1087 245296 1121 246072
rect 1201 245296 1235 246072
rect 1297 245296 1331 246072
rect 1411 245296 1445 246072
rect 1507 245296 1541 246072
rect 1621 245296 1655 246072
rect 1717 245296 1751 246072
rect 1831 245296 1865 246072
rect 1927 245296 1961 246072
rect 2041 245296 2075 246072
rect 2137 245296 2171 246072
rect 2251 245296 2285 246072
rect 2347 245296 2381 246072
rect 2461 245296 2495 246072
rect 2557 245296 2591 246072
rect 2671 245296 2705 246072
rect 2767 245296 2801 246072
rect 2881 245296 2915 246072
rect 2977 245296 3011 246072
rect 3091 245296 3125 246072
rect 3187 245296 3221 246072
rect 3301 245296 3335 246072
rect 3397 245296 3431 246072
rect 3511 245296 3545 246072
rect 3607 245296 3641 246072
rect 3721 245296 3755 246072
rect 3817 245296 3851 246072
rect 3931 245296 3965 246072
rect 4027 245296 4061 246072
rect 4141 245296 4175 246072
rect 4237 245296 4271 246072
rect 4351 245296 4385 246072
rect 4447 245296 4481 246072
rect 4561 245296 4595 246072
rect 4657 245296 4691 246072
rect 4771 245296 4805 246072
rect 4867 245296 4901 246072
rect 4981 245296 5015 246072
rect 5077 245296 5111 246072
rect 5191 245296 5225 246072
rect 5287 245296 5321 246072
rect 5401 245296 5435 246072
rect 5497 245296 5531 246072
rect 5611 245296 5645 246072
rect 5707 245296 5741 246072
rect 5821 245296 5855 246072
rect 5917 245296 5951 246072
rect 6031 245296 6065 246072
rect 6127 245296 6161 246072
rect 6241 245296 6275 246072
rect 6337 245296 6371 246072
rect 6451 245296 6485 246072
rect 6547 245296 6581 246072
rect 6661 245296 6695 246072
rect 6757 245296 6791 246072
rect 6871 245296 6905 246072
rect 6967 245296 7001 246072
rect 7081 245296 7115 246072
rect 7177 245296 7211 246072
rect 7291 245296 7325 246072
rect 7387 245296 7421 246072
rect 7501 245296 7535 246072
rect 7597 245296 7631 246072
rect 7711 245296 7745 246072
rect 7807 245296 7841 246072
rect 7921 245296 7955 246072
rect 8017 245296 8051 246072
rect 8131 245296 8165 246072
rect 8227 245296 8261 246072
rect 8341 245296 8375 246072
rect 8437 245296 8471 246072
rect 8551 245296 8585 246072
rect 8647 245296 8681 246072
rect 8761 245296 8795 246072
rect 8857 245296 8891 246072
rect 8971 245296 9005 246072
rect 9067 245296 9101 246072
rect 9181 245296 9215 246072
rect 9277 245296 9311 246072
rect 9391 245296 9425 246072
rect 9487 245296 9521 246072
rect 9601 245296 9635 246072
rect 9697 245296 9731 246072
rect 9811 245296 9845 246072
rect 9907 245296 9941 246072
rect 10021 245296 10055 246072
rect 10117 245296 10151 246072
rect 10231 245296 10265 246072
rect 10327 245296 10361 246072
rect 10441 245296 10475 246072
rect 10537 245296 10571 246072
rect 10651 245296 10685 246072
rect 10747 245296 10781 246072
rect 10861 245296 10895 246072
rect 10957 245296 10991 246072
rect 11071 245296 11105 246072
rect 11167 245296 11201 246072
rect 11281 245296 11315 246072
rect 11377 245296 11411 246072
rect 11491 245296 11525 246072
rect 11587 245296 11621 246072
rect 11701 245296 11735 246072
rect 11797 245296 11831 246072
rect 11911 245296 11945 246072
rect 12007 245296 12041 246072
rect 12121 245296 12155 246072
rect 12217 245296 12251 246072
rect 12331 245296 12365 246072
rect 12427 245296 12461 246072
rect 12541 245296 12575 246072
rect 12637 245296 12671 246072
rect 12751 245296 12785 246072
rect 12847 245296 12881 246072
rect 12961 245296 12995 246072
rect 13057 245296 13091 246072
rect 13171 245296 13205 246072
rect 13267 245296 13301 246072
rect 13381 245296 13415 246072
rect 13477 245296 13511 246072
rect 13591 245296 13625 246072
rect 13687 245296 13721 246072
rect 13801 245296 13835 246072
rect 13897 245296 13931 246072
rect 14011 245296 14045 246072
rect 14107 245296 14141 246072
rect 14221 245296 14255 246072
rect 14317 245296 14351 246072
rect 14431 245296 14465 246072
rect 14527 245296 14561 246072
rect 14641 245296 14675 246072
rect 14737 245296 14771 246072
rect 14851 245296 14885 246072
rect 14947 245296 14981 246072
rect 15061 245296 15095 246072
rect 15157 245296 15191 246072
rect 15271 245296 15305 246072
rect 15367 245296 15401 246072
rect 15481 245296 15515 246072
rect 15577 245296 15611 246072
rect 15691 245296 15725 246072
rect 15787 245296 15821 246072
rect 15901 245296 15935 246072
rect 15997 245296 16031 246072
rect 16111 245296 16145 246072
rect 16207 245296 16241 246072
rect 16321 245296 16355 246072
rect 16417 245296 16451 246072
rect 16531 245296 16565 246072
rect 16627 245296 16661 246072
rect 16741 245296 16775 246072
rect 16837 245296 16871 246072
rect 16951 245296 16985 246072
rect 17047 245296 17081 246072
rect 17161 245296 17195 246072
rect 17257 245296 17291 246072
rect 17371 245296 17405 246072
rect 17467 245296 17501 246072
rect 17581 245296 17615 246072
rect 17677 245296 17711 246072
rect 17791 245296 17825 246072
rect 17887 245296 17921 246072
rect 18001 245296 18035 246072
rect 18097 245296 18131 246072
rect 18211 245296 18245 246072
rect 18307 245296 18341 246072
rect 18421 245296 18455 246072
rect 18517 245296 18551 246072
rect 18631 245296 18665 246072
rect 18727 245296 18761 246072
rect 18841 245296 18875 246072
rect 18937 245296 18971 246072
rect 19051 245296 19085 246072
rect 19147 245296 19181 246072
rect 19261 245296 19295 246072
rect 19357 245296 19391 246072
rect 19471 245296 19505 246072
rect 19567 245296 19601 246072
rect 19681 245296 19715 246072
rect 19777 245296 19811 246072
rect 19891 245296 19925 246072
rect 19987 245296 20021 246072
rect 20101 245296 20135 246072
rect 20197 245296 20231 246072
rect 20311 245296 20345 246072
rect 20407 245296 20441 246072
rect 20521 245296 20555 246072
rect 20617 245296 20651 246072
rect 20731 245296 20765 246072
rect 20827 245296 20861 246072
rect 20941 245296 20975 246072
rect 21037 245296 21071 246072
rect 21151 245296 21185 246072
rect 21247 245296 21281 246072
rect 21361 245296 21395 246072
rect 21457 245296 21491 246072
rect 21571 245296 21605 246072
rect 21667 245296 21701 246072
rect 21781 245296 21815 246072
rect 21877 245296 21911 246072
rect 21991 245296 22025 246072
rect 22087 245296 22121 246072
rect 22201 245296 22235 246072
rect 22297 245296 22331 246072
rect 22411 245296 22445 246072
rect 22507 245296 22541 246072
rect 22621 245296 22655 246072
rect 22717 245296 22751 246072
rect 22831 245296 22865 246072
rect 22927 245296 22961 246072
rect 23041 245296 23075 246072
rect 23137 245296 23171 246072
rect 23251 245296 23285 246072
rect 23347 245296 23381 246072
rect 23461 245296 23495 246072
rect 23557 245296 23591 246072
rect 23671 245296 23705 246072
rect 23767 245296 23801 246072
rect 23881 245296 23915 246072
rect 23977 245296 24011 246072
rect 24091 245296 24125 246072
rect 24187 245296 24221 246072
rect 24301 245296 24335 246072
rect 24397 245296 24431 246072
rect 24511 245296 24545 246072
rect 24607 245296 24641 246072
rect 24721 245296 24755 246072
rect 24817 245296 24851 246072
rect 24931 245296 24965 246072
rect 25027 245296 25061 246072
rect 25141 245296 25175 246072
rect 25237 245296 25271 246072
rect 25351 245296 25385 246072
rect 25447 245296 25481 246072
rect 25561 245296 25595 246072
rect 25657 245296 25691 246072
rect 25771 245296 25805 246072
rect 25867 245296 25901 246072
rect 25981 245296 26015 246072
rect 26077 245296 26111 246072
rect 26191 245296 26225 246072
rect 26287 245296 26321 246072
rect 26401 245296 26435 246072
rect 26497 245296 26531 246072
rect 26611 245296 26645 246072
rect 26707 245296 26741 246072
rect 26821 245296 26855 246072
rect 26917 245296 26951 246072
rect 27031 245296 27065 246072
rect 27127 245296 27161 246072
rect 27241 245296 27275 246072
rect 27337 245296 27371 246072
rect -4049 244260 -4015 245036
rect -3953 244260 -3919 245036
rect -3839 244260 -3805 245036
rect -3743 244260 -3709 245036
rect -3629 244260 -3595 245036
rect -3533 244260 -3499 245036
rect -3419 244260 -3385 245036
rect -3323 244260 -3289 245036
rect -3209 244260 -3175 245036
rect -3113 244260 -3079 245036
rect -2999 244260 -2965 245036
rect -2903 244260 -2869 245036
rect -2789 244260 -2755 245036
rect -2693 244260 -2659 245036
rect -2579 244260 -2545 245036
rect -2483 244260 -2449 245036
rect -2369 244260 -2335 245036
rect -2273 244260 -2239 245036
rect -2159 244260 -2125 245036
rect -2063 244260 -2029 245036
rect -1949 244260 -1915 245036
rect -1853 244260 -1819 245036
rect -1739 244260 -1705 245036
rect -1643 244260 -1609 245036
rect -1529 244260 -1495 245036
rect -1433 244260 -1399 245036
rect -1319 244260 -1285 245036
rect -1223 244260 -1189 245036
rect -1109 244260 -1075 245036
rect -1013 244260 -979 245036
rect -899 244260 -865 245036
rect -803 244260 -769 245036
rect -689 244260 -655 245036
rect -593 244260 -559 245036
rect -479 244260 -445 245036
rect -383 244260 -349 245036
rect -269 244260 -235 245036
rect -173 244260 -139 245036
rect -59 244260 -25 245036
rect 37 244260 71 245036
rect 151 244260 185 245036
rect 247 244260 281 245036
rect 361 244260 395 245036
rect 457 244260 491 245036
rect 571 244260 605 245036
rect 667 244260 701 245036
rect 781 244260 815 245036
rect 877 244260 911 245036
rect 991 244260 1025 245036
rect 1087 244260 1121 245036
rect 1201 244260 1235 245036
rect 1297 244260 1331 245036
rect 1411 244260 1445 245036
rect 1507 244260 1541 245036
rect 1621 244260 1655 245036
rect 1717 244260 1751 245036
rect 1831 244260 1865 245036
rect 1927 244260 1961 245036
rect 2041 244260 2075 245036
rect 2137 244260 2171 245036
rect 2251 244260 2285 245036
rect 2347 244260 2381 245036
rect 2461 244260 2495 245036
rect 2557 244260 2591 245036
rect 2671 244260 2705 245036
rect 2767 244260 2801 245036
rect 2881 244260 2915 245036
rect 2977 244260 3011 245036
rect 3091 244260 3125 245036
rect 3187 244260 3221 245036
rect 3301 244260 3335 245036
rect 3397 244260 3431 245036
rect 3511 244260 3545 245036
rect 3607 244260 3641 245036
rect 3721 244260 3755 245036
rect 3817 244260 3851 245036
rect 3931 244260 3965 245036
rect 4027 244260 4061 245036
rect 4141 244260 4175 245036
rect 4237 244260 4271 245036
rect 4351 244260 4385 245036
rect 4447 244260 4481 245036
rect 4561 244260 4595 245036
rect 4657 244260 4691 245036
rect 4771 244260 4805 245036
rect 4867 244260 4901 245036
rect 4981 244260 5015 245036
rect 5077 244260 5111 245036
rect 5191 244260 5225 245036
rect 5287 244260 5321 245036
rect 5401 244260 5435 245036
rect 5497 244260 5531 245036
rect 5611 244260 5645 245036
rect 5707 244260 5741 245036
rect 5821 244260 5855 245036
rect 5917 244260 5951 245036
rect 6031 244260 6065 245036
rect 6127 244260 6161 245036
rect 6241 244260 6275 245036
rect 6337 244260 6371 245036
rect 6451 244260 6485 245036
rect 6547 244260 6581 245036
rect 6661 244260 6695 245036
rect 6757 244260 6791 245036
rect 6871 244260 6905 245036
rect 6967 244260 7001 245036
rect 7081 244260 7115 245036
rect 7177 244260 7211 245036
rect 7291 244260 7325 245036
rect 7387 244260 7421 245036
rect 7501 244260 7535 245036
rect 7597 244260 7631 245036
rect 7711 244260 7745 245036
rect 7807 244260 7841 245036
rect 7921 244260 7955 245036
rect 8017 244260 8051 245036
rect 8131 244260 8165 245036
rect 8227 244260 8261 245036
rect 8341 244260 8375 245036
rect 8437 244260 8471 245036
rect 8551 244260 8585 245036
rect 8647 244260 8681 245036
rect 8761 244260 8795 245036
rect 8857 244260 8891 245036
rect 8971 244260 9005 245036
rect 9067 244260 9101 245036
rect 9181 244260 9215 245036
rect 9277 244260 9311 245036
rect 9391 244260 9425 245036
rect 9487 244260 9521 245036
rect 9601 244260 9635 245036
rect 9697 244260 9731 245036
rect 9811 244260 9845 245036
rect 9907 244260 9941 245036
rect 10021 244260 10055 245036
rect 10117 244260 10151 245036
rect 10231 244260 10265 245036
rect 10327 244260 10361 245036
rect 10441 244260 10475 245036
rect 10537 244260 10571 245036
rect 10651 244260 10685 245036
rect 10747 244260 10781 245036
rect 10861 244260 10895 245036
rect 10957 244260 10991 245036
rect 11071 244260 11105 245036
rect 11167 244260 11201 245036
rect 11281 244260 11315 245036
rect 11377 244260 11411 245036
rect 11491 244260 11525 245036
rect 11587 244260 11621 245036
rect 11701 244260 11735 245036
rect 11797 244260 11831 245036
rect 11911 244260 11945 245036
rect 12007 244260 12041 245036
rect 12121 244260 12155 245036
rect 12217 244260 12251 245036
rect 12331 244260 12365 245036
rect 12427 244260 12461 245036
rect 12541 244260 12575 245036
rect 12637 244260 12671 245036
rect 12751 244260 12785 245036
rect 12847 244260 12881 245036
rect 12961 244260 12995 245036
rect 13057 244260 13091 245036
rect 13171 244260 13205 245036
rect 13267 244260 13301 245036
rect 13381 244260 13415 245036
rect 13477 244260 13511 245036
rect 13591 244260 13625 245036
rect 13687 244260 13721 245036
rect 13801 244260 13835 245036
rect 13897 244260 13931 245036
rect 14011 244260 14045 245036
rect 14107 244260 14141 245036
rect 14221 244260 14255 245036
rect 14317 244260 14351 245036
rect 14431 244260 14465 245036
rect 14527 244260 14561 245036
rect 14641 244260 14675 245036
rect 14737 244260 14771 245036
rect 14851 244260 14885 245036
rect 14947 244260 14981 245036
rect 15061 244260 15095 245036
rect 15157 244260 15191 245036
rect 15271 244260 15305 245036
rect 15367 244260 15401 245036
rect 15481 244260 15515 245036
rect 15577 244260 15611 245036
rect 15691 244260 15725 245036
rect 15787 244260 15821 245036
rect 15901 244260 15935 245036
rect 15997 244260 16031 245036
rect 16111 244260 16145 245036
rect 16207 244260 16241 245036
rect 16321 244260 16355 245036
rect 16417 244260 16451 245036
rect 16531 244260 16565 245036
rect 16627 244260 16661 245036
rect 16741 244260 16775 245036
rect 16837 244260 16871 245036
rect 16951 244260 16985 245036
rect 17047 244260 17081 245036
rect 17161 244260 17195 245036
rect 17257 244260 17291 245036
rect 17371 244260 17405 245036
rect 17467 244260 17501 245036
rect 17581 244260 17615 245036
rect 17677 244260 17711 245036
rect 17791 244260 17825 245036
rect 17887 244260 17921 245036
rect 18001 244260 18035 245036
rect 18097 244260 18131 245036
rect 18211 244260 18245 245036
rect 18307 244260 18341 245036
rect 18421 244260 18455 245036
rect 18517 244260 18551 245036
rect 18631 244260 18665 245036
rect 18727 244260 18761 245036
rect 18841 244260 18875 245036
rect 18937 244260 18971 245036
rect 19051 244260 19085 245036
rect 19147 244260 19181 245036
rect 19261 244260 19295 245036
rect 19357 244260 19391 245036
rect 19471 244260 19505 245036
rect 19567 244260 19601 245036
rect 19681 244260 19715 245036
rect 19777 244260 19811 245036
rect 19891 244260 19925 245036
rect 19987 244260 20021 245036
rect 20101 244260 20135 245036
rect 20197 244260 20231 245036
rect 20311 244260 20345 245036
rect 20407 244260 20441 245036
rect 20521 244260 20555 245036
rect 20617 244260 20651 245036
rect 20731 244260 20765 245036
rect 20827 244260 20861 245036
rect 20941 244260 20975 245036
rect 21037 244260 21071 245036
rect 21151 244260 21185 245036
rect 21247 244260 21281 245036
rect 21361 244260 21395 245036
rect 21457 244260 21491 245036
rect 21571 244260 21605 245036
rect 21667 244260 21701 245036
rect 21781 244260 21815 245036
rect 21877 244260 21911 245036
rect 21991 244260 22025 245036
rect 22087 244260 22121 245036
rect 22201 244260 22235 245036
rect 22297 244260 22331 245036
rect 22411 244260 22445 245036
rect 22507 244260 22541 245036
rect 22621 244260 22655 245036
rect 22717 244260 22751 245036
rect 22831 244260 22865 245036
rect 22927 244260 22961 245036
rect 23041 244260 23075 245036
rect 23137 244260 23171 245036
rect 23251 244260 23285 245036
rect 23347 244260 23381 245036
rect 23461 244260 23495 245036
rect 23557 244260 23591 245036
rect 23671 244260 23705 245036
rect 23767 244260 23801 245036
rect 23881 244260 23915 245036
rect 23977 244260 24011 245036
rect 24091 244260 24125 245036
rect 24187 244260 24221 245036
rect 24301 244260 24335 245036
rect 24397 244260 24431 245036
rect 24511 244260 24545 245036
rect 24607 244260 24641 245036
rect 24721 244260 24755 245036
rect 24817 244260 24851 245036
rect 24931 244260 24965 245036
rect 25027 244260 25061 245036
rect 25141 244260 25175 245036
rect 25237 244260 25271 245036
rect 25351 244260 25385 245036
rect 25447 244260 25481 245036
rect 25561 244260 25595 245036
rect 25657 244260 25691 245036
rect 25771 244260 25805 245036
rect 25867 244260 25901 245036
rect 25981 244260 26015 245036
rect 26077 244260 26111 245036
rect 26191 244260 26225 245036
rect 26287 244260 26321 245036
rect 26401 244260 26435 245036
rect 26497 244260 26531 245036
rect 26611 244260 26645 245036
rect 26707 244260 26741 245036
rect 26821 244260 26855 245036
rect 26917 244260 26951 245036
rect 27031 244260 27065 245036
rect 27127 244260 27161 245036
rect 27241 244260 27275 245036
rect 27337 244260 27371 245036
<< psubdiff >>
rect -4163 264178 -4067 264212
rect 27389 264178 27485 264212
rect -4163 264116 -4129 264178
rect 27451 264116 27485 264178
rect -4163 262076 -4129 262138
rect 27451 262076 27485 262138
rect -4163 262042 -4067 262076
rect 27389 262042 27485 262076
<< nsubdiff >>
rect -4163 254650 -4067 254684
rect 27389 254650 27485 254684
rect -4163 254588 -4129 254650
rect 27451 254588 27485 254650
rect -4163 249408 -4129 249470
rect 27451 249408 27485 249470
rect -4163 249341 -4067 249408
rect 27389 249375 27485 249408
rect 27389 249341 27485 249374
rect -4163 249279 -4129 249341
rect 27451 249279 27485 249341
rect -4163 244099 -4129 244161
rect 27451 244099 27485 244161
rect -4163 244065 -4067 244099
rect 27389 244065 27485 244099
<< psubdiffcont >>
rect -4067 264178 27389 264212
rect -4163 262138 -4129 264116
rect 27451 262138 27485 264116
rect -4067 262042 27389 262076
<< nsubdiffcont >>
rect -4067 254650 27389 254684
rect -4163 249470 -4129 254588
rect 27451 249470 27485 254588
rect -4067 249375 27389 249408
rect -4067 249374 27485 249375
rect -4067 249341 27389 249374
rect -4163 244161 -4129 249279
rect 27451 244161 27485 249279
rect -4067 244065 27389 244099
<< poly >>
rect -4017 264110 -3888 264126
rect -4017 264076 -4001 264110
rect -3905 264076 -3888 264110
rect -4017 264060 -3888 264076
rect -3597 264110 -3468 264126
rect -3597 264076 -3581 264110
rect -3485 264076 -3468 264110
rect -3999 264038 -3969 264060
rect -3789 264038 -3759 264064
rect -3597 264060 -3468 264076
rect -3177 264110 -3048 264126
rect -3177 264076 -3161 264110
rect -3065 264076 -3048 264110
rect -3579 264038 -3549 264060
rect -3369 264038 -3339 264064
rect -3177 264060 -3048 264076
rect -2757 264110 -2628 264126
rect -2757 264076 -2741 264110
rect -2645 264076 -2628 264110
rect -3159 264038 -3129 264060
rect -2949 264038 -2919 264064
rect -2757 264060 -2628 264076
rect -2337 264110 -2208 264126
rect -2337 264076 -2321 264110
rect -2225 264076 -2208 264110
rect -2739 264038 -2709 264060
rect -2529 264038 -2499 264064
rect -2337 264060 -2208 264076
rect -1917 264110 -1788 264126
rect -1917 264076 -1901 264110
rect -1805 264076 -1788 264110
rect -2319 264038 -2289 264060
rect -2109 264038 -2079 264064
rect -1917 264060 -1788 264076
rect -1497 264110 -1368 264126
rect -1497 264076 -1481 264110
rect -1385 264076 -1368 264110
rect -1899 264038 -1869 264060
rect -1689 264038 -1659 264064
rect -1497 264060 -1368 264076
rect -1077 264110 -948 264126
rect -1077 264076 -1061 264110
rect -965 264076 -948 264110
rect -1479 264038 -1449 264060
rect -1269 264038 -1239 264064
rect -1077 264060 -948 264076
rect -657 264110 -528 264126
rect -657 264076 -641 264110
rect -545 264076 -528 264110
rect -1059 264038 -1029 264060
rect -849 264038 -819 264064
rect -657 264060 -528 264076
rect -237 264110 -108 264126
rect -237 264076 -221 264110
rect -125 264076 -108 264110
rect -639 264038 -609 264060
rect -429 264038 -399 264064
rect -237 264060 -108 264076
rect 183 264110 312 264126
rect 183 264076 199 264110
rect 295 264076 312 264110
rect -219 264038 -189 264060
rect -9 264038 21 264064
rect 183 264060 312 264076
rect 603 264110 732 264126
rect 603 264076 619 264110
rect 715 264076 732 264110
rect 201 264038 231 264060
rect 411 264038 441 264064
rect 603 264060 732 264076
rect 1023 264110 1152 264126
rect 1023 264076 1039 264110
rect 1135 264076 1152 264110
rect 621 264038 651 264060
rect 831 264038 861 264064
rect 1023 264060 1152 264076
rect 1443 264110 1572 264126
rect 1443 264076 1459 264110
rect 1555 264076 1572 264110
rect 1041 264038 1071 264060
rect 1251 264038 1281 264064
rect 1443 264060 1572 264076
rect 1863 264110 1992 264126
rect 1863 264076 1879 264110
rect 1975 264076 1992 264110
rect 1461 264038 1491 264060
rect 1671 264038 1701 264064
rect 1863 264060 1992 264076
rect 2283 264110 2412 264126
rect 2283 264076 2299 264110
rect 2395 264076 2412 264110
rect 1881 264038 1911 264060
rect 2091 264038 2121 264064
rect 2283 264060 2412 264076
rect 2703 264110 2832 264126
rect 2703 264076 2719 264110
rect 2815 264076 2832 264110
rect 2301 264038 2331 264060
rect 2511 264038 2541 264064
rect 2703 264060 2832 264076
rect 3123 264110 3252 264126
rect 3123 264076 3139 264110
rect 3235 264076 3252 264110
rect 2721 264038 2751 264060
rect 2931 264038 2961 264064
rect 3123 264060 3252 264076
rect 3543 264110 3672 264126
rect 3543 264076 3559 264110
rect 3655 264076 3672 264110
rect 3141 264038 3171 264060
rect 3351 264038 3381 264064
rect 3543 264060 3672 264076
rect 3963 264110 4092 264126
rect 3963 264076 3979 264110
rect 4075 264076 4092 264110
rect 3561 264038 3591 264060
rect 3771 264038 3801 264064
rect 3963 264060 4092 264076
rect 4383 264110 4512 264126
rect 4383 264076 4399 264110
rect 4495 264076 4512 264110
rect 3981 264038 4011 264060
rect 4191 264038 4221 264064
rect 4383 264060 4512 264076
rect 4803 264110 4932 264126
rect 4803 264076 4819 264110
rect 4915 264076 4932 264110
rect 4401 264038 4431 264060
rect 4611 264038 4641 264064
rect 4803 264060 4932 264076
rect 5223 264110 5352 264126
rect 5223 264076 5239 264110
rect 5335 264076 5352 264110
rect 4821 264038 4851 264060
rect 5031 264038 5061 264064
rect 5223 264060 5352 264076
rect 5643 264110 5772 264126
rect 5643 264076 5659 264110
rect 5755 264076 5772 264110
rect 5241 264038 5271 264060
rect 5451 264038 5481 264064
rect 5643 264060 5772 264076
rect 6063 264110 6192 264126
rect 6063 264076 6079 264110
rect 6175 264076 6192 264110
rect 5661 264038 5691 264060
rect 5871 264038 5901 264064
rect 6063 264060 6192 264076
rect 6483 264110 6612 264126
rect 6483 264076 6499 264110
rect 6595 264076 6612 264110
rect 6081 264038 6111 264060
rect 6291 264038 6321 264064
rect 6483 264060 6612 264076
rect 6903 264110 7032 264126
rect 6903 264076 6919 264110
rect 7015 264076 7032 264110
rect 6501 264038 6531 264060
rect 6711 264038 6741 264064
rect 6903 264060 7032 264076
rect 7323 264110 7452 264126
rect 7323 264076 7339 264110
rect 7435 264076 7452 264110
rect 6921 264038 6951 264060
rect 7131 264038 7161 264064
rect 7323 264060 7452 264076
rect 7743 264110 7872 264126
rect 7743 264076 7759 264110
rect 7855 264076 7872 264110
rect 7341 264038 7371 264060
rect 7551 264038 7581 264064
rect 7743 264060 7872 264076
rect 8163 264110 8292 264126
rect 8163 264076 8179 264110
rect 8275 264076 8292 264110
rect 7761 264038 7791 264060
rect 7971 264038 8001 264064
rect 8163 264060 8292 264076
rect 8583 264110 8712 264126
rect 8583 264076 8599 264110
rect 8695 264076 8712 264110
rect 8181 264038 8211 264060
rect 8391 264038 8421 264064
rect 8583 264060 8712 264076
rect 9003 264110 9132 264126
rect 9003 264076 9019 264110
rect 9115 264076 9132 264110
rect 8601 264038 8631 264060
rect 8811 264038 8841 264064
rect 9003 264060 9132 264076
rect 9423 264110 9552 264126
rect 9423 264076 9439 264110
rect 9535 264076 9552 264110
rect 9021 264038 9051 264060
rect 9231 264038 9261 264064
rect 9423 264060 9552 264076
rect 9843 264110 9972 264126
rect 9843 264076 9859 264110
rect 9955 264076 9972 264110
rect 9441 264038 9471 264060
rect 9651 264038 9681 264064
rect 9843 264060 9972 264076
rect 10263 264110 10392 264126
rect 10263 264076 10279 264110
rect 10375 264076 10392 264110
rect 9861 264038 9891 264060
rect 10071 264038 10101 264064
rect 10263 264060 10392 264076
rect 10683 264110 10812 264126
rect 10683 264076 10699 264110
rect 10795 264076 10812 264110
rect 10281 264038 10311 264060
rect 10491 264038 10521 264064
rect 10683 264060 10812 264076
rect 11103 264110 11232 264126
rect 11103 264076 11119 264110
rect 11215 264076 11232 264110
rect 10701 264038 10731 264060
rect 10911 264038 10941 264064
rect 11103 264060 11232 264076
rect 11523 264110 11652 264126
rect 11523 264076 11539 264110
rect 11635 264076 11652 264110
rect 11121 264038 11151 264060
rect 11331 264038 11361 264064
rect 11523 264060 11652 264076
rect 11943 264110 12072 264126
rect 11943 264076 11959 264110
rect 12055 264076 12072 264110
rect 11541 264038 11571 264060
rect 11751 264038 11781 264064
rect 11943 264060 12072 264076
rect 12363 264110 12492 264126
rect 12363 264076 12379 264110
rect 12475 264076 12492 264110
rect 11961 264038 11991 264060
rect 12171 264038 12201 264064
rect 12363 264060 12492 264076
rect 12783 264110 12912 264126
rect 12783 264076 12799 264110
rect 12895 264076 12912 264110
rect 12381 264038 12411 264060
rect 12591 264038 12621 264064
rect 12783 264060 12912 264076
rect 13203 264110 13332 264126
rect 13203 264076 13219 264110
rect 13315 264076 13332 264110
rect 12801 264038 12831 264060
rect 13011 264038 13041 264064
rect 13203 264060 13332 264076
rect 13623 264110 13752 264126
rect 13623 264076 13639 264110
rect 13735 264076 13752 264110
rect 13221 264038 13251 264060
rect 13431 264038 13461 264064
rect 13623 264060 13752 264076
rect 14043 264110 14172 264126
rect 14043 264076 14059 264110
rect 14155 264076 14172 264110
rect 13641 264038 13671 264060
rect 13851 264038 13881 264064
rect 14043 264060 14172 264076
rect 14463 264110 14592 264126
rect 14463 264076 14479 264110
rect 14575 264076 14592 264110
rect 14061 264038 14091 264060
rect 14271 264038 14301 264064
rect 14463 264060 14592 264076
rect 14883 264110 15012 264126
rect 14883 264076 14899 264110
rect 14995 264076 15012 264110
rect 14481 264038 14511 264060
rect 14691 264038 14721 264064
rect 14883 264060 15012 264076
rect 15303 264110 15432 264126
rect 15303 264076 15319 264110
rect 15415 264076 15432 264110
rect 14901 264038 14931 264060
rect 15111 264038 15141 264064
rect 15303 264060 15432 264076
rect 15723 264110 15852 264126
rect 15723 264076 15739 264110
rect 15835 264076 15852 264110
rect 15321 264038 15351 264060
rect 15531 264038 15561 264064
rect 15723 264060 15852 264076
rect 16143 264110 16272 264126
rect 16143 264076 16159 264110
rect 16255 264076 16272 264110
rect 15741 264038 15771 264060
rect 15951 264038 15981 264064
rect 16143 264060 16272 264076
rect 16563 264110 16692 264126
rect 16563 264076 16579 264110
rect 16675 264076 16692 264110
rect 16161 264038 16191 264060
rect 16371 264038 16401 264064
rect 16563 264060 16692 264076
rect 16983 264110 17112 264126
rect 16983 264076 16999 264110
rect 17095 264076 17112 264110
rect 16581 264038 16611 264060
rect 16791 264038 16821 264064
rect 16983 264060 17112 264076
rect 17403 264110 17532 264126
rect 17403 264076 17419 264110
rect 17515 264076 17532 264110
rect 17001 264038 17031 264060
rect 17211 264038 17241 264064
rect 17403 264060 17532 264076
rect 17823 264110 17952 264126
rect 17823 264076 17839 264110
rect 17935 264076 17952 264110
rect 17421 264038 17451 264060
rect 17631 264038 17661 264064
rect 17823 264060 17952 264076
rect 18243 264110 18372 264126
rect 18243 264076 18259 264110
rect 18355 264076 18372 264110
rect 17841 264038 17871 264060
rect 18051 264038 18081 264064
rect 18243 264060 18372 264076
rect 18663 264110 18792 264126
rect 18663 264076 18679 264110
rect 18775 264076 18792 264110
rect 18261 264038 18291 264060
rect 18471 264038 18501 264064
rect 18663 264060 18792 264076
rect 19083 264110 19212 264126
rect 19083 264076 19099 264110
rect 19195 264076 19212 264110
rect 18681 264038 18711 264060
rect 18891 264038 18921 264064
rect 19083 264060 19212 264076
rect 19503 264110 19632 264126
rect 19503 264076 19519 264110
rect 19615 264076 19632 264110
rect 19101 264038 19131 264060
rect 19311 264038 19341 264064
rect 19503 264060 19632 264076
rect 19923 264110 20052 264126
rect 19923 264076 19939 264110
rect 20035 264076 20052 264110
rect 19521 264038 19551 264060
rect 19731 264038 19761 264064
rect 19923 264060 20052 264076
rect 20343 264110 20472 264126
rect 20343 264076 20359 264110
rect 20455 264076 20472 264110
rect 19941 264038 19971 264060
rect 20151 264038 20181 264064
rect 20343 264060 20472 264076
rect 20763 264110 20892 264126
rect 20763 264076 20779 264110
rect 20875 264076 20892 264110
rect 20361 264038 20391 264060
rect 20571 264038 20601 264064
rect 20763 264060 20892 264076
rect 21183 264110 21312 264126
rect 21183 264076 21199 264110
rect 21295 264076 21312 264110
rect 20781 264038 20811 264060
rect 20991 264038 21021 264064
rect 21183 264060 21312 264076
rect 21603 264110 21732 264126
rect 21603 264076 21619 264110
rect 21715 264076 21732 264110
rect 21201 264038 21231 264060
rect 21411 264038 21441 264064
rect 21603 264060 21732 264076
rect 22023 264110 22152 264126
rect 22023 264076 22039 264110
rect 22135 264076 22152 264110
rect 21621 264038 21651 264060
rect 21831 264038 21861 264064
rect 22023 264060 22152 264076
rect 22443 264110 22572 264126
rect 22443 264076 22459 264110
rect 22555 264076 22572 264110
rect 22041 264038 22071 264060
rect 22251 264038 22281 264064
rect 22443 264060 22572 264076
rect 22863 264110 22992 264126
rect 22863 264076 22879 264110
rect 22975 264076 22992 264110
rect 22461 264038 22491 264060
rect 22671 264038 22701 264064
rect 22863 264060 22992 264076
rect 23283 264110 23412 264126
rect 23283 264076 23299 264110
rect 23395 264076 23412 264110
rect 22881 264038 22911 264060
rect 23091 264038 23121 264064
rect 23283 264060 23412 264076
rect 23703 264110 23832 264126
rect 23703 264076 23719 264110
rect 23815 264076 23832 264110
rect 23301 264038 23331 264060
rect 23511 264038 23541 264064
rect 23703 264060 23832 264076
rect 24123 264110 24252 264126
rect 24123 264076 24139 264110
rect 24235 264076 24252 264110
rect 23721 264038 23751 264060
rect 23931 264038 23961 264064
rect 24123 264060 24252 264076
rect 24543 264110 24672 264126
rect 24543 264076 24559 264110
rect 24655 264076 24672 264110
rect 24141 264038 24171 264060
rect 24351 264038 24381 264064
rect 24543 264060 24672 264076
rect 24963 264110 25092 264126
rect 24963 264076 24979 264110
rect 25075 264076 25092 264110
rect 24561 264038 24591 264060
rect 24771 264038 24801 264064
rect 24963 264060 25092 264076
rect 25383 264110 25512 264126
rect 25383 264076 25399 264110
rect 25495 264076 25512 264110
rect 24981 264038 25011 264060
rect 25191 264038 25221 264064
rect 25383 264060 25512 264076
rect 25803 264110 25932 264126
rect 25803 264076 25819 264110
rect 25915 264076 25932 264110
rect 25401 264038 25431 264060
rect 25611 264038 25641 264064
rect 25803 264060 25932 264076
rect 26223 264110 26352 264126
rect 26223 264076 26239 264110
rect 26335 264076 26352 264110
rect 25821 264038 25851 264060
rect 26031 264038 26061 264064
rect 26223 264060 26352 264076
rect 26643 264110 26772 264126
rect 26643 264076 26659 264110
rect 26755 264076 26772 264110
rect 26241 264038 26271 264060
rect 26451 264038 26481 264064
rect 26643 264060 26772 264076
rect 27063 264110 27192 264126
rect 27063 264076 27079 264110
rect 27175 264076 27192 264110
rect 26661 264038 26691 264060
rect 26871 264038 26901 264064
rect 27063 264060 27192 264076
rect 27081 264038 27111 264060
rect 27291 264038 27321 264064
rect -3999 263210 -3969 263238
rect -3789 263214 -3759 263238
rect -3807 263198 -3741 263214
rect -3579 263210 -3549 263238
rect -3369 263214 -3339 263238
rect -3807 263164 -3791 263198
rect -3757 263164 -3741 263198
rect -3807 263090 -3741 263164
rect -3807 263056 -3791 263090
rect -3757 263056 -3741 263090
rect -3999 263016 -3969 263044
rect -3807 263040 -3741 263056
rect -3387 263198 -3321 263214
rect -3159 263210 -3129 263238
rect -2949 263214 -2919 263238
rect -3387 263164 -3371 263198
rect -3337 263164 -3321 263198
rect -3387 263090 -3321 263164
rect -3387 263056 -3371 263090
rect -3337 263056 -3321 263090
rect -3789 263016 -3759 263040
rect -3579 263016 -3549 263044
rect -3387 263040 -3321 263056
rect -2967 263198 -2901 263214
rect -2739 263210 -2709 263238
rect -2529 263214 -2499 263238
rect -2967 263164 -2951 263198
rect -2917 263164 -2901 263198
rect -2967 263090 -2901 263164
rect -2967 263056 -2951 263090
rect -2917 263056 -2901 263090
rect -3369 263016 -3339 263040
rect -3159 263016 -3129 263044
rect -2967 263040 -2901 263056
rect -2547 263198 -2481 263214
rect -2319 263210 -2289 263238
rect -2109 263214 -2079 263238
rect -2547 263164 -2531 263198
rect -2497 263164 -2481 263198
rect -2547 263090 -2481 263164
rect -2547 263056 -2531 263090
rect -2497 263056 -2481 263090
rect -2949 263016 -2919 263040
rect -2739 263016 -2709 263044
rect -2547 263040 -2481 263056
rect -2127 263198 -2061 263214
rect -1899 263210 -1869 263238
rect -1689 263214 -1659 263238
rect -2127 263164 -2111 263198
rect -2077 263164 -2061 263198
rect -2127 263090 -2061 263164
rect -2127 263056 -2111 263090
rect -2077 263056 -2061 263090
rect -2529 263016 -2499 263040
rect -2319 263016 -2289 263044
rect -2127 263040 -2061 263056
rect -1707 263198 -1641 263214
rect -1479 263210 -1449 263238
rect -1269 263214 -1239 263238
rect -1707 263164 -1691 263198
rect -1657 263164 -1641 263198
rect -1707 263090 -1641 263164
rect -1707 263056 -1691 263090
rect -1657 263056 -1641 263090
rect -2109 263016 -2079 263040
rect -1899 263016 -1869 263044
rect -1707 263040 -1641 263056
rect -1287 263198 -1221 263214
rect -1059 263210 -1029 263238
rect -849 263214 -819 263238
rect -1287 263164 -1271 263198
rect -1237 263164 -1221 263198
rect -1287 263090 -1221 263164
rect -1287 263056 -1271 263090
rect -1237 263056 -1221 263090
rect -1689 263016 -1659 263040
rect -1479 263016 -1449 263044
rect -1287 263040 -1221 263056
rect -867 263198 -801 263214
rect -639 263210 -609 263238
rect -429 263214 -399 263238
rect -867 263164 -851 263198
rect -817 263164 -801 263198
rect -867 263090 -801 263164
rect -867 263056 -851 263090
rect -817 263056 -801 263090
rect -1269 263016 -1239 263040
rect -1059 263016 -1029 263044
rect -867 263040 -801 263056
rect -447 263198 -381 263214
rect -219 263210 -189 263238
rect -9 263214 21 263238
rect -447 263164 -431 263198
rect -397 263164 -381 263198
rect -447 263090 -381 263164
rect -447 263056 -431 263090
rect -397 263056 -381 263090
rect -849 263016 -819 263040
rect -639 263016 -609 263044
rect -447 263040 -381 263056
rect -27 263198 39 263214
rect 201 263210 231 263238
rect 411 263214 441 263238
rect -27 263164 -11 263198
rect 23 263164 39 263198
rect -27 263090 39 263164
rect -27 263056 -11 263090
rect 23 263056 39 263090
rect -429 263016 -399 263040
rect -219 263016 -189 263044
rect -27 263040 39 263056
rect 393 263198 459 263214
rect 621 263210 651 263238
rect 831 263214 861 263238
rect 393 263164 409 263198
rect 443 263164 459 263198
rect 393 263090 459 263164
rect 393 263056 409 263090
rect 443 263056 459 263090
rect -9 263016 21 263040
rect 201 263016 231 263044
rect 393 263040 459 263056
rect 813 263198 879 263214
rect 1041 263210 1071 263238
rect 1251 263214 1281 263238
rect 813 263164 829 263198
rect 863 263164 879 263198
rect 813 263090 879 263164
rect 813 263056 829 263090
rect 863 263056 879 263090
rect 411 263016 441 263040
rect 621 263016 651 263044
rect 813 263040 879 263056
rect 1233 263198 1299 263214
rect 1461 263210 1491 263238
rect 1671 263214 1701 263238
rect 1233 263164 1249 263198
rect 1283 263164 1299 263198
rect 1233 263090 1299 263164
rect 1233 263056 1249 263090
rect 1283 263056 1299 263090
rect 831 263016 861 263040
rect 1041 263016 1071 263044
rect 1233 263040 1299 263056
rect 1653 263198 1719 263214
rect 1881 263210 1911 263238
rect 2091 263214 2121 263238
rect 1653 263164 1669 263198
rect 1703 263164 1719 263198
rect 1653 263090 1719 263164
rect 1653 263056 1669 263090
rect 1703 263056 1719 263090
rect 1251 263016 1281 263040
rect 1461 263016 1491 263044
rect 1653 263040 1719 263056
rect 2073 263198 2139 263214
rect 2301 263210 2331 263238
rect 2511 263214 2541 263238
rect 2073 263164 2089 263198
rect 2123 263164 2139 263198
rect 2073 263090 2139 263164
rect 2073 263056 2089 263090
rect 2123 263056 2139 263090
rect 1671 263016 1701 263040
rect 1881 263016 1911 263044
rect 2073 263040 2139 263056
rect 2493 263198 2559 263214
rect 2721 263210 2751 263238
rect 2931 263214 2961 263238
rect 2493 263164 2509 263198
rect 2543 263164 2559 263198
rect 2493 263090 2559 263164
rect 2493 263056 2509 263090
rect 2543 263056 2559 263090
rect 2091 263016 2121 263040
rect 2301 263016 2331 263044
rect 2493 263040 2559 263056
rect 2913 263198 2979 263214
rect 3141 263210 3171 263238
rect 3351 263214 3381 263238
rect 2913 263164 2929 263198
rect 2963 263164 2979 263198
rect 2913 263090 2979 263164
rect 2913 263056 2929 263090
rect 2963 263056 2979 263090
rect 2511 263016 2541 263040
rect 2721 263016 2751 263044
rect 2913 263040 2979 263056
rect 3333 263198 3399 263214
rect 3561 263210 3591 263238
rect 3771 263214 3801 263238
rect 3333 263164 3349 263198
rect 3383 263164 3399 263198
rect 3333 263090 3399 263164
rect 3333 263056 3349 263090
rect 3383 263056 3399 263090
rect 2931 263016 2961 263040
rect 3141 263016 3171 263044
rect 3333 263040 3399 263056
rect 3753 263198 3819 263214
rect 3981 263210 4011 263238
rect 4191 263214 4221 263238
rect 3753 263164 3769 263198
rect 3803 263164 3819 263198
rect 3753 263090 3819 263164
rect 3753 263056 3769 263090
rect 3803 263056 3819 263090
rect 3351 263016 3381 263040
rect 3561 263016 3591 263044
rect 3753 263040 3819 263056
rect 4173 263198 4239 263214
rect 4401 263210 4431 263238
rect 4611 263214 4641 263238
rect 4173 263164 4189 263198
rect 4223 263164 4239 263198
rect 4173 263090 4239 263164
rect 4173 263056 4189 263090
rect 4223 263056 4239 263090
rect 3771 263016 3801 263040
rect 3981 263016 4011 263044
rect 4173 263040 4239 263056
rect 4593 263198 4659 263214
rect 4821 263210 4851 263238
rect 5031 263214 5061 263238
rect 4593 263164 4609 263198
rect 4643 263164 4659 263198
rect 4593 263090 4659 263164
rect 4593 263056 4609 263090
rect 4643 263056 4659 263090
rect 4191 263016 4221 263040
rect 4401 263016 4431 263044
rect 4593 263040 4659 263056
rect 5013 263198 5079 263214
rect 5241 263210 5271 263238
rect 5451 263214 5481 263238
rect 5013 263164 5029 263198
rect 5063 263164 5079 263198
rect 5013 263090 5079 263164
rect 5013 263056 5029 263090
rect 5063 263056 5079 263090
rect 4611 263016 4641 263040
rect 4821 263016 4851 263044
rect 5013 263040 5079 263056
rect 5433 263198 5499 263214
rect 5661 263210 5691 263238
rect 5871 263214 5901 263238
rect 5433 263164 5449 263198
rect 5483 263164 5499 263198
rect 5433 263090 5499 263164
rect 5433 263056 5449 263090
rect 5483 263056 5499 263090
rect 5031 263016 5061 263040
rect 5241 263016 5271 263044
rect 5433 263040 5499 263056
rect 5853 263198 5919 263214
rect 6081 263210 6111 263238
rect 6291 263214 6321 263238
rect 5853 263164 5869 263198
rect 5903 263164 5919 263198
rect 5853 263090 5919 263164
rect 5853 263056 5869 263090
rect 5903 263056 5919 263090
rect 5451 263016 5481 263040
rect 5661 263016 5691 263044
rect 5853 263040 5919 263056
rect 6273 263198 6339 263214
rect 6501 263210 6531 263238
rect 6711 263214 6741 263238
rect 6273 263164 6289 263198
rect 6323 263164 6339 263198
rect 6273 263090 6339 263164
rect 6273 263056 6289 263090
rect 6323 263056 6339 263090
rect 5871 263016 5901 263040
rect 6081 263016 6111 263044
rect 6273 263040 6339 263056
rect 6693 263198 6759 263214
rect 6921 263210 6951 263238
rect 7131 263214 7161 263238
rect 6693 263164 6709 263198
rect 6743 263164 6759 263198
rect 6693 263090 6759 263164
rect 6693 263056 6709 263090
rect 6743 263056 6759 263090
rect 6291 263016 6321 263040
rect 6501 263016 6531 263044
rect 6693 263040 6759 263056
rect 7113 263198 7179 263214
rect 7341 263210 7371 263238
rect 7551 263214 7581 263238
rect 7113 263164 7129 263198
rect 7163 263164 7179 263198
rect 7113 263090 7179 263164
rect 7113 263056 7129 263090
rect 7163 263056 7179 263090
rect 6711 263016 6741 263040
rect 6921 263016 6951 263044
rect 7113 263040 7179 263056
rect 7533 263198 7599 263214
rect 7761 263210 7791 263238
rect 7971 263214 8001 263238
rect 7533 263164 7549 263198
rect 7583 263164 7599 263198
rect 7533 263090 7599 263164
rect 7533 263056 7549 263090
rect 7583 263056 7599 263090
rect 7131 263016 7161 263040
rect 7341 263016 7371 263044
rect 7533 263040 7599 263056
rect 7953 263198 8019 263214
rect 8181 263210 8211 263238
rect 8391 263214 8421 263238
rect 7953 263164 7969 263198
rect 8003 263164 8019 263198
rect 7953 263090 8019 263164
rect 7953 263056 7969 263090
rect 8003 263056 8019 263090
rect 7551 263016 7581 263040
rect 7761 263016 7791 263044
rect 7953 263040 8019 263056
rect 8373 263198 8439 263214
rect 8601 263210 8631 263238
rect 8811 263214 8841 263238
rect 8373 263164 8389 263198
rect 8423 263164 8439 263198
rect 8373 263090 8439 263164
rect 8373 263056 8389 263090
rect 8423 263056 8439 263090
rect 7971 263016 8001 263040
rect 8181 263016 8211 263044
rect 8373 263040 8439 263056
rect 8793 263198 8859 263214
rect 9021 263210 9051 263238
rect 9231 263214 9261 263238
rect 8793 263164 8809 263198
rect 8843 263164 8859 263198
rect 8793 263090 8859 263164
rect 8793 263056 8809 263090
rect 8843 263056 8859 263090
rect 8391 263016 8421 263040
rect 8601 263016 8631 263044
rect 8793 263040 8859 263056
rect 9213 263198 9279 263214
rect 9441 263210 9471 263238
rect 9651 263214 9681 263238
rect 9213 263164 9229 263198
rect 9263 263164 9279 263198
rect 9213 263090 9279 263164
rect 9213 263056 9229 263090
rect 9263 263056 9279 263090
rect 8811 263016 8841 263040
rect 9021 263016 9051 263044
rect 9213 263040 9279 263056
rect 9633 263198 9699 263214
rect 9861 263210 9891 263238
rect 10071 263214 10101 263238
rect 9633 263164 9649 263198
rect 9683 263164 9699 263198
rect 9633 263090 9699 263164
rect 9633 263056 9649 263090
rect 9683 263056 9699 263090
rect 9231 263016 9261 263040
rect 9441 263016 9471 263044
rect 9633 263040 9699 263056
rect 10053 263198 10119 263214
rect 10281 263210 10311 263238
rect 10491 263214 10521 263238
rect 10053 263164 10069 263198
rect 10103 263164 10119 263198
rect 10053 263090 10119 263164
rect 10053 263056 10069 263090
rect 10103 263056 10119 263090
rect 9651 263016 9681 263040
rect 9861 263016 9891 263044
rect 10053 263040 10119 263056
rect 10473 263198 10539 263214
rect 10701 263210 10731 263238
rect 10911 263214 10941 263238
rect 10473 263164 10489 263198
rect 10523 263164 10539 263198
rect 10473 263090 10539 263164
rect 10473 263056 10489 263090
rect 10523 263056 10539 263090
rect 10071 263016 10101 263040
rect 10281 263016 10311 263044
rect 10473 263040 10539 263056
rect 10893 263198 10959 263214
rect 11121 263210 11151 263238
rect 11331 263214 11361 263238
rect 10893 263164 10909 263198
rect 10943 263164 10959 263198
rect 10893 263090 10959 263164
rect 10893 263056 10909 263090
rect 10943 263056 10959 263090
rect 10491 263016 10521 263040
rect 10701 263016 10731 263044
rect 10893 263040 10959 263056
rect 11313 263198 11379 263214
rect 11541 263210 11571 263238
rect 11751 263214 11781 263238
rect 11313 263164 11329 263198
rect 11363 263164 11379 263198
rect 11313 263090 11379 263164
rect 11313 263056 11329 263090
rect 11363 263056 11379 263090
rect 10911 263016 10941 263040
rect 11121 263016 11151 263044
rect 11313 263040 11379 263056
rect 11733 263198 11799 263214
rect 11961 263210 11991 263238
rect 12171 263214 12201 263238
rect 11733 263164 11749 263198
rect 11783 263164 11799 263198
rect 11733 263090 11799 263164
rect 11733 263056 11749 263090
rect 11783 263056 11799 263090
rect 11331 263016 11361 263040
rect 11541 263016 11571 263044
rect 11733 263040 11799 263056
rect 12153 263198 12219 263214
rect 12381 263210 12411 263238
rect 12591 263214 12621 263238
rect 12153 263164 12169 263198
rect 12203 263164 12219 263198
rect 12153 263090 12219 263164
rect 12153 263056 12169 263090
rect 12203 263056 12219 263090
rect 11751 263016 11781 263040
rect 11961 263016 11991 263044
rect 12153 263040 12219 263056
rect 12573 263198 12639 263214
rect 12801 263210 12831 263238
rect 13011 263214 13041 263238
rect 12573 263164 12589 263198
rect 12623 263164 12639 263198
rect 12573 263090 12639 263164
rect 12573 263056 12589 263090
rect 12623 263056 12639 263090
rect 12171 263016 12201 263040
rect 12381 263016 12411 263044
rect 12573 263040 12639 263056
rect 12993 263198 13059 263214
rect 13221 263210 13251 263238
rect 13431 263214 13461 263238
rect 12993 263164 13009 263198
rect 13043 263164 13059 263198
rect 12993 263090 13059 263164
rect 12993 263056 13009 263090
rect 13043 263056 13059 263090
rect 12591 263016 12621 263040
rect 12801 263016 12831 263044
rect 12993 263040 13059 263056
rect 13413 263198 13479 263214
rect 13641 263210 13671 263238
rect 13851 263214 13881 263238
rect 13413 263164 13429 263198
rect 13463 263164 13479 263198
rect 13413 263090 13479 263164
rect 13413 263056 13429 263090
rect 13463 263056 13479 263090
rect 13011 263016 13041 263040
rect 13221 263016 13251 263044
rect 13413 263040 13479 263056
rect 13833 263198 13899 263214
rect 14061 263210 14091 263238
rect 14271 263214 14301 263238
rect 13833 263164 13849 263198
rect 13883 263164 13899 263198
rect 13833 263090 13899 263164
rect 13833 263056 13849 263090
rect 13883 263056 13899 263090
rect 13431 263016 13461 263040
rect 13641 263016 13671 263044
rect 13833 263040 13899 263056
rect 14253 263198 14319 263214
rect 14481 263210 14511 263238
rect 14691 263214 14721 263238
rect 14253 263164 14269 263198
rect 14303 263164 14319 263198
rect 14253 263090 14319 263164
rect 14253 263056 14269 263090
rect 14303 263056 14319 263090
rect 13851 263016 13881 263040
rect 14061 263016 14091 263044
rect 14253 263040 14319 263056
rect 14673 263198 14739 263214
rect 14901 263210 14931 263238
rect 15111 263214 15141 263238
rect 14673 263164 14689 263198
rect 14723 263164 14739 263198
rect 14673 263090 14739 263164
rect 14673 263056 14689 263090
rect 14723 263056 14739 263090
rect 14271 263016 14301 263040
rect 14481 263016 14511 263044
rect 14673 263040 14739 263056
rect 15093 263198 15159 263214
rect 15321 263210 15351 263238
rect 15531 263214 15561 263238
rect 15093 263164 15109 263198
rect 15143 263164 15159 263198
rect 15093 263090 15159 263164
rect 15093 263056 15109 263090
rect 15143 263056 15159 263090
rect 14691 263016 14721 263040
rect 14901 263016 14931 263044
rect 15093 263040 15159 263056
rect 15513 263198 15579 263214
rect 15741 263210 15771 263238
rect 15951 263214 15981 263238
rect 15513 263164 15529 263198
rect 15563 263164 15579 263198
rect 15513 263090 15579 263164
rect 15513 263056 15529 263090
rect 15563 263056 15579 263090
rect 15111 263016 15141 263040
rect 15321 263016 15351 263044
rect 15513 263040 15579 263056
rect 15933 263198 15999 263214
rect 16161 263210 16191 263238
rect 16371 263214 16401 263238
rect 15933 263164 15949 263198
rect 15983 263164 15999 263198
rect 15933 263090 15999 263164
rect 15933 263056 15949 263090
rect 15983 263056 15999 263090
rect 15531 263016 15561 263040
rect 15741 263016 15771 263044
rect 15933 263040 15999 263056
rect 16353 263198 16419 263214
rect 16581 263210 16611 263238
rect 16791 263214 16821 263238
rect 16353 263164 16369 263198
rect 16403 263164 16419 263198
rect 16353 263090 16419 263164
rect 16353 263056 16369 263090
rect 16403 263056 16419 263090
rect 15951 263016 15981 263040
rect 16161 263016 16191 263044
rect 16353 263040 16419 263056
rect 16773 263198 16839 263214
rect 17001 263210 17031 263238
rect 17211 263214 17241 263238
rect 16773 263164 16789 263198
rect 16823 263164 16839 263198
rect 16773 263090 16839 263164
rect 16773 263056 16789 263090
rect 16823 263056 16839 263090
rect 16371 263016 16401 263040
rect 16581 263016 16611 263044
rect 16773 263040 16839 263056
rect 17193 263198 17259 263214
rect 17421 263210 17451 263238
rect 17631 263214 17661 263238
rect 17193 263164 17209 263198
rect 17243 263164 17259 263198
rect 17193 263090 17259 263164
rect 17193 263056 17209 263090
rect 17243 263056 17259 263090
rect 16791 263016 16821 263040
rect 17001 263016 17031 263044
rect 17193 263040 17259 263056
rect 17613 263198 17679 263214
rect 17841 263210 17871 263238
rect 18051 263214 18081 263238
rect 17613 263164 17629 263198
rect 17663 263164 17679 263198
rect 17613 263090 17679 263164
rect 17613 263056 17629 263090
rect 17663 263056 17679 263090
rect 17211 263016 17241 263040
rect 17421 263016 17451 263044
rect 17613 263040 17679 263056
rect 18033 263198 18099 263214
rect 18261 263210 18291 263238
rect 18471 263214 18501 263238
rect 18033 263164 18049 263198
rect 18083 263164 18099 263198
rect 18033 263090 18099 263164
rect 18033 263056 18049 263090
rect 18083 263056 18099 263090
rect 17631 263016 17661 263040
rect 17841 263016 17871 263044
rect 18033 263040 18099 263056
rect 18453 263198 18519 263214
rect 18681 263210 18711 263238
rect 18891 263214 18921 263238
rect 18453 263164 18469 263198
rect 18503 263164 18519 263198
rect 18453 263090 18519 263164
rect 18453 263056 18469 263090
rect 18503 263056 18519 263090
rect 18051 263016 18081 263040
rect 18261 263016 18291 263044
rect 18453 263040 18519 263056
rect 18873 263198 18939 263214
rect 19101 263210 19131 263238
rect 19311 263214 19341 263238
rect 18873 263164 18889 263198
rect 18923 263164 18939 263198
rect 18873 263090 18939 263164
rect 18873 263056 18889 263090
rect 18923 263056 18939 263090
rect 18471 263016 18501 263040
rect 18681 263016 18711 263044
rect 18873 263040 18939 263056
rect 19293 263198 19359 263214
rect 19521 263210 19551 263238
rect 19731 263214 19761 263238
rect 19293 263164 19309 263198
rect 19343 263164 19359 263198
rect 19293 263090 19359 263164
rect 19293 263056 19309 263090
rect 19343 263056 19359 263090
rect 18891 263016 18921 263040
rect 19101 263016 19131 263044
rect 19293 263040 19359 263056
rect 19713 263198 19779 263214
rect 19941 263210 19971 263238
rect 20151 263214 20181 263238
rect 19713 263164 19729 263198
rect 19763 263164 19779 263198
rect 19713 263090 19779 263164
rect 19713 263056 19729 263090
rect 19763 263056 19779 263090
rect 19311 263016 19341 263040
rect 19521 263016 19551 263044
rect 19713 263040 19779 263056
rect 20133 263198 20199 263214
rect 20361 263210 20391 263238
rect 20571 263214 20601 263238
rect 20133 263164 20149 263198
rect 20183 263164 20199 263198
rect 20133 263090 20199 263164
rect 20133 263056 20149 263090
rect 20183 263056 20199 263090
rect 19731 263016 19761 263040
rect 19941 263016 19971 263044
rect 20133 263040 20199 263056
rect 20553 263198 20619 263214
rect 20781 263210 20811 263238
rect 20991 263214 21021 263238
rect 20553 263164 20569 263198
rect 20603 263164 20619 263198
rect 20553 263090 20619 263164
rect 20553 263056 20569 263090
rect 20603 263056 20619 263090
rect 20151 263016 20181 263040
rect 20361 263016 20391 263044
rect 20553 263040 20619 263056
rect 20973 263198 21039 263214
rect 21201 263210 21231 263238
rect 21411 263214 21441 263238
rect 20973 263164 20989 263198
rect 21023 263164 21039 263198
rect 20973 263090 21039 263164
rect 20973 263056 20989 263090
rect 21023 263056 21039 263090
rect 20571 263016 20601 263040
rect 20781 263016 20811 263044
rect 20973 263040 21039 263056
rect 21393 263198 21459 263214
rect 21621 263210 21651 263238
rect 21831 263214 21861 263238
rect 21393 263164 21409 263198
rect 21443 263164 21459 263198
rect 21393 263090 21459 263164
rect 21393 263056 21409 263090
rect 21443 263056 21459 263090
rect 20991 263016 21021 263040
rect 21201 263016 21231 263044
rect 21393 263040 21459 263056
rect 21813 263198 21879 263214
rect 22041 263210 22071 263238
rect 22251 263214 22281 263238
rect 21813 263164 21829 263198
rect 21863 263164 21879 263198
rect 21813 263090 21879 263164
rect 21813 263056 21829 263090
rect 21863 263056 21879 263090
rect 21411 263016 21441 263040
rect 21621 263016 21651 263044
rect 21813 263040 21879 263056
rect 22233 263198 22299 263214
rect 22461 263210 22491 263238
rect 22671 263214 22701 263238
rect 22233 263164 22249 263198
rect 22283 263164 22299 263198
rect 22233 263090 22299 263164
rect 22233 263056 22249 263090
rect 22283 263056 22299 263090
rect 21831 263016 21861 263040
rect 22041 263016 22071 263044
rect 22233 263040 22299 263056
rect 22653 263198 22719 263214
rect 22881 263210 22911 263238
rect 23091 263214 23121 263238
rect 22653 263164 22669 263198
rect 22703 263164 22719 263198
rect 22653 263090 22719 263164
rect 22653 263056 22669 263090
rect 22703 263056 22719 263090
rect 22251 263016 22281 263040
rect 22461 263016 22491 263044
rect 22653 263040 22719 263056
rect 23073 263198 23139 263214
rect 23301 263210 23331 263238
rect 23511 263214 23541 263238
rect 23073 263164 23089 263198
rect 23123 263164 23139 263198
rect 23073 263090 23139 263164
rect 23073 263056 23089 263090
rect 23123 263056 23139 263090
rect 22671 263016 22701 263040
rect 22881 263016 22911 263044
rect 23073 263040 23139 263056
rect 23493 263198 23559 263214
rect 23721 263210 23751 263238
rect 23931 263214 23961 263238
rect 23493 263164 23509 263198
rect 23543 263164 23559 263198
rect 23493 263090 23559 263164
rect 23493 263056 23509 263090
rect 23543 263056 23559 263090
rect 23091 263016 23121 263040
rect 23301 263016 23331 263044
rect 23493 263040 23559 263056
rect 23913 263198 23979 263214
rect 24141 263210 24171 263238
rect 24351 263214 24381 263238
rect 23913 263164 23929 263198
rect 23963 263164 23979 263198
rect 23913 263090 23979 263164
rect 23913 263056 23929 263090
rect 23963 263056 23979 263090
rect 23511 263016 23541 263040
rect 23721 263016 23751 263044
rect 23913 263040 23979 263056
rect 24333 263198 24399 263214
rect 24561 263210 24591 263238
rect 24771 263214 24801 263238
rect 24333 263164 24349 263198
rect 24383 263164 24399 263198
rect 24333 263090 24399 263164
rect 24333 263056 24349 263090
rect 24383 263056 24399 263090
rect 23931 263016 23961 263040
rect 24141 263016 24171 263044
rect 24333 263040 24399 263056
rect 24753 263198 24819 263214
rect 24981 263210 25011 263238
rect 25191 263214 25221 263238
rect 24753 263164 24769 263198
rect 24803 263164 24819 263198
rect 24753 263090 24819 263164
rect 24753 263056 24769 263090
rect 24803 263056 24819 263090
rect 24351 263016 24381 263040
rect 24561 263016 24591 263044
rect 24753 263040 24819 263056
rect 25173 263198 25239 263214
rect 25401 263210 25431 263238
rect 25611 263214 25641 263238
rect 25173 263164 25189 263198
rect 25223 263164 25239 263198
rect 25173 263090 25239 263164
rect 25173 263056 25189 263090
rect 25223 263056 25239 263090
rect 24771 263016 24801 263040
rect 24981 263016 25011 263044
rect 25173 263040 25239 263056
rect 25593 263198 25659 263214
rect 25821 263210 25851 263238
rect 26031 263214 26061 263238
rect 25593 263164 25609 263198
rect 25643 263164 25659 263198
rect 25593 263090 25659 263164
rect 25593 263056 25609 263090
rect 25643 263056 25659 263090
rect 25191 263016 25221 263040
rect 25401 263016 25431 263044
rect 25593 263040 25659 263056
rect 26013 263198 26079 263214
rect 26241 263210 26271 263238
rect 26451 263214 26481 263238
rect 26013 263164 26029 263198
rect 26063 263164 26079 263198
rect 26013 263090 26079 263164
rect 26013 263056 26029 263090
rect 26063 263056 26079 263090
rect 25611 263016 25641 263040
rect 25821 263016 25851 263044
rect 26013 263040 26079 263056
rect 26433 263198 26499 263214
rect 26661 263210 26691 263238
rect 26871 263214 26901 263238
rect 26433 263164 26449 263198
rect 26483 263164 26499 263198
rect 26433 263090 26499 263164
rect 26433 263056 26449 263090
rect 26483 263056 26499 263090
rect 26031 263016 26061 263040
rect 26241 263016 26271 263044
rect 26433 263040 26499 263056
rect 26853 263198 26919 263214
rect 27081 263210 27111 263238
rect 27291 263214 27321 263238
rect 26853 263164 26869 263198
rect 26903 263164 26919 263198
rect 26853 263090 26919 263164
rect 26853 263056 26869 263090
rect 26903 263056 26919 263090
rect 26451 263016 26481 263040
rect 26661 263016 26691 263044
rect 26853 263040 26919 263056
rect 27273 263198 27339 263214
rect 27273 263164 27289 263198
rect 27323 263164 27339 263198
rect 27273 263090 27339 263164
rect 27273 263056 27289 263090
rect 27323 263056 27339 263090
rect 26871 263016 26901 263040
rect 27081 263016 27111 263044
rect 27273 263040 27339 263056
rect 27291 263016 27321 263040
rect -3999 262194 -3969 262216
rect -4017 262178 -3888 262194
rect -3789 262190 -3759 262216
rect -3579 262194 -3549 262216
rect -4017 262144 -4001 262178
rect -3905 262144 -3888 262178
rect -4017 262128 -3888 262144
rect -3597 262178 -3468 262194
rect -3369 262190 -3339 262216
rect -3159 262194 -3129 262216
rect -3597 262144 -3581 262178
rect -3485 262144 -3468 262178
rect -3597 262128 -3468 262144
rect -3177 262178 -3048 262194
rect -2949 262190 -2919 262216
rect -2739 262194 -2709 262216
rect -3177 262144 -3161 262178
rect -3065 262144 -3048 262178
rect -3177 262128 -3048 262144
rect -2757 262178 -2628 262194
rect -2529 262190 -2499 262216
rect -2319 262194 -2289 262216
rect -2757 262144 -2741 262178
rect -2645 262144 -2628 262178
rect -2757 262128 -2628 262144
rect -2337 262178 -2208 262194
rect -2109 262190 -2079 262216
rect -1899 262194 -1869 262216
rect -2337 262144 -2321 262178
rect -2225 262144 -2208 262178
rect -2337 262128 -2208 262144
rect -1917 262178 -1788 262194
rect -1689 262190 -1659 262216
rect -1479 262194 -1449 262216
rect -1917 262144 -1901 262178
rect -1805 262144 -1788 262178
rect -1917 262128 -1788 262144
rect -1497 262178 -1368 262194
rect -1269 262190 -1239 262216
rect -1059 262194 -1029 262216
rect -1497 262144 -1481 262178
rect -1385 262144 -1368 262178
rect -1497 262128 -1368 262144
rect -1077 262178 -948 262194
rect -849 262190 -819 262216
rect -639 262194 -609 262216
rect -1077 262144 -1061 262178
rect -965 262144 -948 262178
rect -1077 262128 -948 262144
rect -657 262178 -528 262194
rect -429 262190 -399 262216
rect -219 262194 -189 262216
rect -657 262144 -641 262178
rect -545 262144 -528 262178
rect -657 262128 -528 262144
rect -237 262178 -108 262194
rect -9 262190 21 262216
rect 201 262194 231 262216
rect -237 262144 -221 262178
rect -125 262144 -108 262178
rect -237 262128 -108 262144
rect 183 262178 312 262194
rect 411 262190 441 262216
rect 621 262194 651 262216
rect 183 262144 199 262178
rect 295 262144 312 262178
rect 183 262128 312 262144
rect 603 262178 732 262194
rect 831 262190 861 262216
rect 1041 262194 1071 262216
rect 603 262144 619 262178
rect 715 262144 732 262178
rect 603 262128 732 262144
rect 1023 262178 1152 262194
rect 1251 262190 1281 262216
rect 1461 262194 1491 262216
rect 1023 262144 1039 262178
rect 1135 262144 1152 262178
rect 1023 262128 1152 262144
rect 1443 262178 1572 262194
rect 1671 262190 1701 262216
rect 1881 262194 1911 262216
rect 1443 262144 1459 262178
rect 1555 262144 1572 262178
rect 1443 262128 1572 262144
rect 1863 262178 1992 262194
rect 2091 262190 2121 262216
rect 2301 262194 2331 262216
rect 1863 262144 1879 262178
rect 1975 262144 1992 262178
rect 1863 262128 1992 262144
rect 2283 262178 2412 262194
rect 2511 262190 2541 262216
rect 2721 262194 2751 262216
rect 2283 262144 2299 262178
rect 2395 262144 2412 262178
rect 2283 262128 2412 262144
rect 2703 262178 2832 262194
rect 2931 262190 2961 262216
rect 3141 262194 3171 262216
rect 2703 262144 2719 262178
rect 2815 262144 2832 262178
rect 2703 262128 2832 262144
rect 3123 262178 3252 262194
rect 3351 262190 3381 262216
rect 3561 262194 3591 262216
rect 3123 262144 3139 262178
rect 3235 262144 3252 262178
rect 3123 262128 3252 262144
rect 3543 262178 3672 262194
rect 3771 262190 3801 262216
rect 3981 262194 4011 262216
rect 3543 262144 3559 262178
rect 3655 262144 3672 262178
rect 3543 262128 3672 262144
rect 3963 262178 4092 262194
rect 4191 262190 4221 262216
rect 4401 262194 4431 262216
rect 3963 262144 3979 262178
rect 4075 262144 4092 262178
rect 3963 262128 4092 262144
rect 4383 262178 4512 262194
rect 4611 262190 4641 262216
rect 4821 262194 4851 262216
rect 4383 262144 4399 262178
rect 4495 262144 4512 262178
rect 4383 262128 4512 262144
rect 4803 262178 4932 262194
rect 5031 262190 5061 262216
rect 5241 262194 5271 262216
rect 4803 262144 4819 262178
rect 4915 262144 4932 262178
rect 4803 262128 4932 262144
rect 5223 262178 5352 262194
rect 5451 262190 5481 262216
rect 5661 262194 5691 262216
rect 5223 262144 5239 262178
rect 5335 262144 5352 262178
rect 5223 262128 5352 262144
rect 5643 262178 5772 262194
rect 5871 262190 5901 262216
rect 6081 262194 6111 262216
rect 5643 262144 5659 262178
rect 5755 262144 5772 262178
rect 5643 262128 5772 262144
rect 6063 262178 6192 262194
rect 6291 262190 6321 262216
rect 6501 262194 6531 262216
rect 6063 262144 6079 262178
rect 6175 262144 6192 262178
rect 6063 262128 6192 262144
rect 6483 262178 6612 262194
rect 6711 262190 6741 262216
rect 6921 262194 6951 262216
rect 6483 262144 6499 262178
rect 6595 262144 6612 262178
rect 6483 262128 6612 262144
rect 6903 262178 7032 262194
rect 7131 262190 7161 262216
rect 7341 262194 7371 262216
rect 6903 262144 6919 262178
rect 7015 262144 7032 262178
rect 6903 262128 7032 262144
rect 7323 262178 7452 262194
rect 7551 262190 7581 262216
rect 7761 262194 7791 262216
rect 7323 262144 7339 262178
rect 7435 262144 7452 262178
rect 7323 262128 7452 262144
rect 7743 262178 7872 262194
rect 7971 262190 8001 262216
rect 8181 262194 8211 262216
rect 7743 262144 7759 262178
rect 7855 262144 7872 262178
rect 7743 262128 7872 262144
rect 8163 262178 8292 262194
rect 8391 262190 8421 262216
rect 8601 262194 8631 262216
rect 8163 262144 8179 262178
rect 8275 262144 8292 262178
rect 8163 262128 8292 262144
rect 8583 262178 8712 262194
rect 8811 262190 8841 262216
rect 9021 262194 9051 262216
rect 8583 262144 8599 262178
rect 8695 262144 8712 262178
rect 8583 262128 8712 262144
rect 9003 262178 9132 262194
rect 9231 262190 9261 262216
rect 9441 262194 9471 262216
rect 9003 262144 9019 262178
rect 9115 262144 9132 262178
rect 9003 262128 9132 262144
rect 9423 262178 9552 262194
rect 9651 262190 9681 262216
rect 9861 262194 9891 262216
rect 9423 262144 9439 262178
rect 9535 262144 9552 262178
rect 9423 262128 9552 262144
rect 9843 262178 9972 262194
rect 10071 262190 10101 262216
rect 10281 262194 10311 262216
rect 9843 262144 9859 262178
rect 9955 262144 9972 262178
rect 9843 262128 9972 262144
rect 10263 262178 10392 262194
rect 10491 262190 10521 262216
rect 10701 262194 10731 262216
rect 10263 262144 10279 262178
rect 10375 262144 10392 262178
rect 10263 262128 10392 262144
rect 10683 262178 10812 262194
rect 10911 262190 10941 262216
rect 11121 262194 11151 262216
rect 10683 262144 10699 262178
rect 10795 262144 10812 262178
rect 10683 262128 10812 262144
rect 11103 262178 11232 262194
rect 11331 262190 11361 262216
rect 11541 262194 11571 262216
rect 11103 262144 11119 262178
rect 11215 262144 11232 262178
rect 11103 262128 11232 262144
rect 11523 262178 11652 262194
rect 11751 262190 11781 262216
rect 11961 262194 11991 262216
rect 11523 262144 11539 262178
rect 11635 262144 11652 262178
rect 11523 262128 11652 262144
rect 11943 262178 12072 262194
rect 12171 262190 12201 262216
rect 12381 262194 12411 262216
rect 11943 262144 11959 262178
rect 12055 262144 12072 262178
rect 11943 262128 12072 262144
rect 12363 262178 12492 262194
rect 12591 262190 12621 262216
rect 12801 262194 12831 262216
rect 12363 262144 12379 262178
rect 12475 262144 12492 262178
rect 12363 262128 12492 262144
rect 12783 262178 12912 262194
rect 13011 262190 13041 262216
rect 13221 262194 13251 262216
rect 12783 262144 12799 262178
rect 12895 262144 12912 262178
rect 12783 262128 12912 262144
rect 13203 262178 13332 262194
rect 13431 262190 13461 262216
rect 13641 262194 13671 262216
rect 13203 262144 13219 262178
rect 13315 262144 13332 262178
rect 13203 262128 13332 262144
rect 13623 262178 13752 262194
rect 13851 262190 13881 262216
rect 14061 262194 14091 262216
rect 13623 262144 13639 262178
rect 13735 262144 13752 262178
rect 13623 262128 13752 262144
rect 14043 262178 14172 262194
rect 14271 262190 14301 262216
rect 14481 262194 14511 262216
rect 14043 262144 14059 262178
rect 14155 262144 14172 262178
rect 14043 262128 14172 262144
rect 14463 262178 14592 262194
rect 14691 262190 14721 262216
rect 14901 262194 14931 262216
rect 14463 262144 14479 262178
rect 14575 262144 14592 262178
rect 14463 262128 14592 262144
rect 14883 262178 15012 262194
rect 15111 262190 15141 262216
rect 15321 262194 15351 262216
rect 14883 262144 14899 262178
rect 14995 262144 15012 262178
rect 14883 262128 15012 262144
rect 15303 262178 15432 262194
rect 15531 262190 15561 262216
rect 15741 262194 15771 262216
rect 15303 262144 15319 262178
rect 15415 262144 15432 262178
rect 15303 262128 15432 262144
rect 15723 262178 15852 262194
rect 15951 262190 15981 262216
rect 16161 262194 16191 262216
rect 15723 262144 15739 262178
rect 15835 262144 15852 262178
rect 15723 262128 15852 262144
rect 16143 262178 16272 262194
rect 16371 262190 16401 262216
rect 16581 262194 16611 262216
rect 16143 262144 16159 262178
rect 16255 262144 16272 262178
rect 16143 262128 16272 262144
rect 16563 262178 16692 262194
rect 16791 262190 16821 262216
rect 17001 262194 17031 262216
rect 16563 262144 16579 262178
rect 16675 262144 16692 262178
rect 16563 262128 16692 262144
rect 16983 262178 17112 262194
rect 17211 262190 17241 262216
rect 17421 262194 17451 262216
rect 16983 262144 16999 262178
rect 17095 262144 17112 262178
rect 16983 262128 17112 262144
rect 17403 262178 17532 262194
rect 17631 262190 17661 262216
rect 17841 262194 17871 262216
rect 17403 262144 17419 262178
rect 17515 262144 17532 262178
rect 17403 262128 17532 262144
rect 17823 262178 17952 262194
rect 18051 262190 18081 262216
rect 18261 262194 18291 262216
rect 17823 262144 17839 262178
rect 17935 262144 17952 262178
rect 17823 262128 17952 262144
rect 18243 262178 18372 262194
rect 18471 262190 18501 262216
rect 18681 262194 18711 262216
rect 18243 262144 18259 262178
rect 18355 262144 18372 262178
rect 18243 262128 18372 262144
rect 18663 262178 18792 262194
rect 18891 262190 18921 262216
rect 19101 262194 19131 262216
rect 18663 262144 18679 262178
rect 18775 262144 18792 262178
rect 18663 262128 18792 262144
rect 19083 262178 19212 262194
rect 19311 262190 19341 262216
rect 19521 262194 19551 262216
rect 19083 262144 19099 262178
rect 19195 262144 19212 262178
rect 19083 262128 19212 262144
rect 19503 262178 19632 262194
rect 19731 262190 19761 262216
rect 19941 262194 19971 262216
rect 19503 262144 19519 262178
rect 19615 262144 19632 262178
rect 19503 262128 19632 262144
rect 19923 262178 20052 262194
rect 20151 262190 20181 262216
rect 20361 262194 20391 262216
rect 19923 262144 19939 262178
rect 20035 262144 20052 262178
rect 19923 262128 20052 262144
rect 20343 262178 20472 262194
rect 20571 262190 20601 262216
rect 20781 262194 20811 262216
rect 20343 262144 20359 262178
rect 20455 262144 20472 262178
rect 20343 262128 20472 262144
rect 20763 262178 20892 262194
rect 20991 262190 21021 262216
rect 21201 262194 21231 262216
rect 20763 262144 20779 262178
rect 20875 262144 20892 262178
rect 20763 262128 20892 262144
rect 21183 262178 21312 262194
rect 21411 262190 21441 262216
rect 21621 262194 21651 262216
rect 21183 262144 21199 262178
rect 21295 262144 21312 262178
rect 21183 262128 21312 262144
rect 21603 262178 21732 262194
rect 21831 262190 21861 262216
rect 22041 262194 22071 262216
rect 21603 262144 21619 262178
rect 21715 262144 21732 262178
rect 21603 262128 21732 262144
rect 22023 262178 22152 262194
rect 22251 262190 22281 262216
rect 22461 262194 22491 262216
rect 22023 262144 22039 262178
rect 22135 262144 22152 262178
rect 22023 262128 22152 262144
rect 22443 262178 22572 262194
rect 22671 262190 22701 262216
rect 22881 262194 22911 262216
rect 22443 262144 22459 262178
rect 22555 262144 22572 262178
rect 22443 262128 22572 262144
rect 22863 262178 22992 262194
rect 23091 262190 23121 262216
rect 23301 262194 23331 262216
rect 22863 262144 22879 262178
rect 22975 262144 22992 262178
rect 22863 262128 22992 262144
rect 23283 262178 23412 262194
rect 23511 262190 23541 262216
rect 23721 262194 23751 262216
rect 23283 262144 23299 262178
rect 23395 262144 23412 262178
rect 23283 262128 23412 262144
rect 23703 262178 23832 262194
rect 23931 262190 23961 262216
rect 24141 262194 24171 262216
rect 23703 262144 23719 262178
rect 23815 262144 23832 262178
rect 23703 262128 23832 262144
rect 24123 262178 24252 262194
rect 24351 262190 24381 262216
rect 24561 262194 24591 262216
rect 24123 262144 24139 262178
rect 24235 262144 24252 262178
rect 24123 262128 24252 262144
rect 24543 262178 24672 262194
rect 24771 262190 24801 262216
rect 24981 262194 25011 262216
rect 24543 262144 24559 262178
rect 24655 262144 24672 262178
rect 24543 262128 24672 262144
rect 24963 262178 25092 262194
rect 25191 262190 25221 262216
rect 25401 262194 25431 262216
rect 24963 262144 24979 262178
rect 25075 262144 25092 262178
rect 24963 262128 25092 262144
rect 25383 262178 25512 262194
rect 25611 262190 25641 262216
rect 25821 262194 25851 262216
rect 25383 262144 25399 262178
rect 25495 262144 25512 262178
rect 25383 262128 25512 262144
rect 25803 262178 25932 262194
rect 26031 262190 26061 262216
rect 26241 262194 26271 262216
rect 25803 262144 25819 262178
rect 25915 262144 25932 262178
rect 25803 262128 25932 262144
rect 26223 262178 26352 262194
rect 26451 262190 26481 262216
rect 26661 262194 26691 262216
rect 26223 262144 26239 262178
rect 26335 262144 26352 262178
rect 26223 262128 26352 262144
rect 26643 262178 26772 262194
rect 26871 262190 26901 262216
rect 27081 262194 27111 262216
rect 26643 262144 26659 262178
rect 26755 262144 26772 262178
rect 26643 262128 26772 262144
rect 27063 262178 27192 262194
rect 27291 262190 27321 262216
rect 27063 262144 27079 262178
rect 27175 262144 27192 262178
rect 27063 262128 27192 262144
rect -4017 254582 -3888 254598
rect -4017 254548 -4001 254582
rect -3905 254548 -3888 254582
rect -4017 254532 -3888 254548
rect -3597 254582 -3468 254598
rect -3597 254548 -3581 254582
rect -3485 254548 -3468 254582
rect -3597 254532 -3468 254548
rect -3177 254582 -3048 254598
rect -3177 254548 -3161 254582
rect -3065 254548 -3048 254582
rect -3177 254532 -3048 254548
rect -2757 254582 -2628 254598
rect -2757 254548 -2741 254582
rect -2645 254548 -2628 254582
rect -2757 254532 -2628 254548
rect -2337 254582 -2208 254598
rect -2337 254548 -2321 254582
rect -2225 254548 -2208 254582
rect -2337 254532 -2208 254548
rect -1917 254582 -1788 254598
rect -1917 254548 -1901 254582
rect -1805 254548 -1788 254582
rect -1917 254532 -1788 254548
rect -1497 254582 -1368 254598
rect -1497 254548 -1481 254582
rect -1385 254548 -1368 254582
rect -1497 254532 -1368 254548
rect -1077 254582 -948 254598
rect -1077 254548 -1061 254582
rect -965 254548 -948 254582
rect -1077 254532 -948 254548
rect -657 254582 -528 254598
rect -657 254548 -641 254582
rect -545 254548 -528 254582
rect -657 254532 -528 254548
rect -237 254582 -108 254598
rect -237 254548 -221 254582
rect -125 254548 -108 254582
rect -237 254532 -108 254548
rect 183 254582 312 254598
rect 183 254548 199 254582
rect 295 254548 312 254582
rect 183 254532 312 254548
rect 603 254582 732 254598
rect 603 254548 619 254582
rect 715 254548 732 254582
rect 603 254532 732 254548
rect 1023 254582 1152 254598
rect 1023 254548 1039 254582
rect 1135 254548 1152 254582
rect 1023 254532 1152 254548
rect 1443 254582 1572 254598
rect 1443 254548 1459 254582
rect 1555 254548 1572 254582
rect 1443 254532 1572 254548
rect 1863 254582 1992 254598
rect 1863 254548 1879 254582
rect 1975 254548 1992 254582
rect 1863 254532 1992 254548
rect 2283 254582 2412 254598
rect 2283 254548 2299 254582
rect 2395 254548 2412 254582
rect 2283 254532 2412 254548
rect 2703 254582 2832 254598
rect 2703 254548 2719 254582
rect 2815 254548 2832 254582
rect 2703 254532 2832 254548
rect 3123 254582 3252 254598
rect 3123 254548 3139 254582
rect 3235 254548 3252 254582
rect 3123 254532 3252 254548
rect 3543 254582 3672 254598
rect 3543 254548 3559 254582
rect 3655 254548 3672 254582
rect 3543 254532 3672 254548
rect 3963 254582 4092 254598
rect 3963 254548 3979 254582
rect 4075 254548 4092 254582
rect 3963 254532 4092 254548
rect 4383 254582 4512 254598
rect 4383 254548 4399 254582
rect 4495 254548 4512 254582
rect 4383 254532 4512 254548
rect 4803 254582 4932 254598
rect 4803 254548 4819 254582
rect 4915 254548 4932 254582
rect 4803 254532 4932 254548
rect 5223 254582 5352 254598
rect 5223 254548 5239 254582
rect 5335 254548 5352 254582
rect 5223 254532 5352 254548
rect 5643 254582 5772 254598
rect 5643 254548 5659 254582
rect 5755 254548 5772 254582
rect 5643 254532 5772 254548
rect 6063 254582 6192 254598
rect 6063 254548 6079 254582
rect 6175 254548 6192 254582
rect 6063 254532 6192 254548
rect 6483 254582 6612 254598
rect 6483 254548 6499 254582
rect 6595 254548 6612 254582
rect 6483 254532 6612 254548
rect 6903 254582 7032 254598
rect 6903 254548 6919 254582
rect 7015 254548 7032 254582
rect 6903 254532 7032 254548
rect 7323 254582 7452 254598
rect 7323 254548 7339 254582
rect 7435 254548 7452 254582
rect 7323 254532 7452 254548
rect 7743 254582 7872 254598
rect 7743 254548 7759 254582
rect 7855 254548 7872 254582
rect 7743 254532 7872 254548
rect 8163 254582 8292 254598
rect 8163 254548 8179 254582
rect 8275 254548 8292 254582
rect 8163 254532 8292 254548
rect 8583 254582 8712 254598
rect 8583 254548 8599 254582
rect 8695 254548 8712 254582
rect 8583 254532 8712 254548
rect 9003 254582 9132 254598
rect 9003 254548 9019 254582
rect 9115 254548 9132 254582
rect 9003 254532 9132 254548
rect 9423 254582 9552 254598
rect 9423 254548 9439 254582
rect 9535 254548 9552 254582
rect 9423 254532 9552 254548
rect 9843 254582 9972 254598
rect 9843 254548 9859 254582
rect 9955 254548 9972 254582
rect 9843 254532 9972 254548
rect 10263 254582 10392 254598
rect 10263 254548 10279 254582
rect 10375 254548 10392 254582
rect 10263 254532 10392 254548
rect 10683 254582 10812 254598
rect 10683 254548 10699 254582
rect 10795 254548 10812 254582
rect 10683 254532 10812 254548
rect 11103 254582 11232 254598
rect 11103 254548 11119 254582
rect 11215 254548 11232 254582
rect 11103 254532 11232 254548
rect 11523 254582 11652 254598
rect 11523 254548 11539 254582
rect 11635 254548 11652 254582
rect 11523 254532 11652 254548
rect 11943 254582 12072 254598
rect 11943 254548 11959 254582
rect 12055 254548 12072 254582
rect 11943 254532 12072 254548
rect 12363 254582 12492 254598
rect 12363 254548 12379 254582
rect 12475 254548 12492 254582
rect 12363 254532 12492 254548
rect 12783 254582 12912 254598
rect 12783 254548 12799 254582
rect 12895 254548 12912 254582
rect 12783 254532 12912 254548
rect 13203 254582 13332 254598
rect 13203 254548 13219 254582
rect 13315 254548 13332 254582
rect 13203 254532 13332 254548
rect 13623 254582 13752 254598
rect 13623 254548 13639 254582
rect 13735 254548 13752 254582
rect 13623 254532 13752 254548
rect 14043 254582 14172 254598
rect 14043 254548 14059 254582
rect 14155 254548 14172 254582
rect 14043 254532 14172 254548
rect 14463 254582 14592 254598
rect 14463 254548 14479 254582
rect 14575 254548 14592 254582
rect 14463 254532 14592 254548
rect 14883 254582 15012 254598
rect 14883 254548 14899 254582
rect 14995 254548 15012 254582
rect 14883 254532 15012 254548
rect 15303 254582 15432 254598
rect 15303 254548 15319 254582
rect 15415 254548 15432 254582
rect 15303 254532 15432 254548
rect 15723 254582 15852 254598
rect 15723 254548 15739 254582
rect 15835 254548 15852 254582
rect 15723 254532 15852 254548
rect 16143 254582 16272 254598
rect 16143 254548 16159 254582
rect 16255 254548 16272 254582
rect 16143 254532 16272 254548
rect 16563 254582 16692 254598
rect 16563 254548 16579 254582
rect 16675 254548 16692 254582
rect 16563 254532 16692 254548
rect 16983 254582 17112 254598
rect 16983 254548 16999 254582
rect 17095 254548 17112 254582
rect 16983 254532 17112 254548
rect 17403 254582 17532 254598
rect 17403 254548 17419 254582
rect 17515 254548 17532 254582
rect 17403 254532 17532 254548
rect 17823 254582 17952 254598
rect 17823 254548 17839 254582
rect 17935 254548 17952 254582
rect 17823 254532 17952 254548
rect 18243 254582 18372 254598
rect 18243 254548 18259 254582
rect 18355 254548 18372 254582
rect 18243 254532 18372 254548
rect 18663 254582 18792 254598
rect 18663 254548 18679 254582
rect 18775 254548 18792 254582
rect 18663 254532 18792 254548
rect 19083 254582 19212 254598
rect 19083 254548 19099 254582
rect 19195 254548 19212 254582
rect 19083 254532 19212 254548
rect 19503 254582 19632 254598
rect 19503 254548 19519 254582
rect 19615 254548 19632 254582
rect 19503 254532 19632 254548
rect 19923 254582 20052 254598
rect 19923 254548 19939 254582
rect 20035 254548 20052 254582
rect 19923 254532 20052 254548
rect 20343 254582 20472 254598
rect 20343 254548 20359 254582
rect 20455 254548 20472 254582
rect 20343 254532 20472 254548
rect 20763 254582 20892 254598
rect 20763 254548 20779 254582
rect 20875 254548 20892 254582
rect 20763 254532 20892 254548
rect 21183 254582 21312 254598
rect 21183 254548 21199 254582
rect 21295 254548 21312 254582
rect 21183 254532 21312 254548
rect 21603 254582 21732 254598
rect 21603 254548 21619 254582
rect 21715 254548 21732 254582
rect 21603 254532 21732 254548
rect 22023 254582 22152 254598
rect 22023 254548 22039 254582
rect 22135 254548 22152 254582
rect 22023 254532 22152 254548
rect 22443 254582 22572 254598
rect 22443 254548 22459 254582
rect 22555 254548 22572 254582
rect 22443 254532 22572 254548
rect 22863 254582 22992 254598
rect 22863 254548 22879 254582
rect 22975 254548 22992 254582
rect 22863 254532 22992 254548
rect 23283 254582 23412 254598
rect 23283 254548 23299 254582
rect 23395 254548 23412 254582
rect 23283 254532 23412 254548
rect 23703 254582 23832 254598
rect 23703 254548 23719 254582
rect 23815 254548 23832 254582
rect 23703 254532 23832 254548
rect 24123 254582 24252 254598
rect 24123 254548 24139 254582
rect 24235 254548 24252 254582
rect 24123 254532 24252 254548
rect 24543 254582 24672 254598
rect 24543 254548 24559 254582
rect 24655 254548 24672 254582
rect 24543 254532 24672 254548
rect 24963 254582 25092 254598
rect 24963 254548 24979 254582
rect 25075 254548 25092 254582
rect 24963 254532 25092 254548
rect 25383 254582 25512 254598
rect 25383 254548 25399 254582
rect 25495 254548 25512 254582
rect 25383 254532 25512 254548
rect 25803 254582 25932 254598
rect 25803 254548 25819 254582
rect 25915 254548 25932 254582
rect 25803 254532 25932 254548
rect 26223 254582 26352 254598
rect 26223 254548 26239 254582
rect 26335 254548 26352 254582
rect 26223 254532 26352 254548
rect 26643 254582 26772 254598
rect 26643 254548 26659 254582
rect 26755 254548 26772 254582
rect 26643 254532 26772 254548
rect 27063 254582 27192 254598
rect 27063 254548 27079 254582
rect 27175 254548 27192 254582
rect 27063 254532 27192 254548
rect -3999 254501 -3969 254532
rect -3789 254501 -3759 254527
rect -3579 254501 -3549 254532
rect -3369 254501 -3339 254527
rect -3159 254501 -3129 254532
rect -2949 254501 -2919 254527
rect -2739 254501 -2709 254532
rect -2529 254501 -2499 254527
rect -2319 254501 -2289 254532
rect -2109 254501 -2079 254527
rect -1899 254501 -1869 254532
rect -1689 254501 -1659 254527
rect -1479 254501 -1449 254532
rect -1269 254501 -1239 254527
rect -1059 254501 -1029 254532
rect -849 254501 -819 254527
rect -639 254501 -609 254532
rect -429 254501 -399 254527
rect -219 254501 -189 254532
rect -9 254501 21 254527
rect 201 254501 231 254532
rect 411 254501 441 254527
rect 621 254501 651 254532
rect 831 254501 861 254527
rect 1041 254501 1071 254532
rect 1251 254501 1281 254527
rect 1461 254501 1491 254532
rect 1671 254501 1701 254527
rect 1881 254501 1911 254532
rect 2091 254501 2121 254527
rect 2301 254501 2331 254532
rect 2511 254501 2541 254527
rect 2721 254501 2751 254532
rect 2931 254501 2961 254527
rect 3141 254501 3171 254532
rect 3351 254501 3381 254527
rect 3561 254501 3591 254532
rect 3771 254501 3801 254527
rect 3981 254501 4011 254532
rect 4191 254501 4221 254527
rect 4401 254501 4431 254532
rect 4611 254501 4641 254527
rect 4821 254501 4851 254532
rect 5031 254501 5061 254527
rect 5241 254501 5271 254532
rect 5451 254501 5481 254527
rect 5661 254501 5691 254532
rect 5871 254501 5901 254527
rect 6081 254501 6111 254532
rect 6291 254501 6321 254527
rect 6501 254501 6531 254532
rect 6711 254501 6741 254527
rect 6921 254501 6951 254532
rect 7131 254501 7161 254527
rect 7341 254501 7371 254532
rect 7551 254501 7581 254527
rect 7761 254501 7791 254532
rect 7971 254501 8001 254527
rect 8181 254501 8211 254532
rect 8391 254501 8421 254527
rect 8601 254501 8631 254532
rect 8811 254501 8841 254527
rect 9021 254501 9051 254532
rect 9231 254501 9261 254527
rect 9441 254501 9471 254532
rect 9651 254501 9681 254527
rect 9861 254501 9891 254532
rect 10071 254501 10101 254527
rect 10281 254501 10311 254532
rect 10491 254501 10521 254527
rect 10701 254501 10731 254532
rect 10911 254501 10941 254527
rect 11121 254501 11151 254532
rect 11331 254501 11361 254527
rect 11541 254501 11571 254532
rect 11751 254501 11781 254527
rect 11961 254501 11991 254532
rect 12171 254501 12201 254527
rect 12381 254501 12411 254532
rect 12591 254501 12621 254527
rect 12801 254501 12831 254532
rect 13011 254501 13041 254527
rect 13221 254501 13251 254532
rect 13431 254501 13461 254527
rect 13641 254501 13671 254532
rect 13851 254501 13881 254527
rect 14061 254501 14091 254532
rect 14271 254501 14301 254527
rect 14481 254501 14511 254532
rect 14691 254501 14721 254527
rect 14901 254501 14931 254532
rect 15111 254501 15141 254527
rect 15321 254501 15351 254532
rect 15531 254501 15561 254527
rect 15741 254501 15771 254532
rect 15951 254501 15981 254527
rect 16161 254501 16191 254532
rect 16371 254501 16401 254527
rect 16581 254501 16611 254532
rect 16791 254501 16821 254527
rect 17001 254501 17031 254532
rect 17211 254501 17241 254527
rect 17421 254501 17451 254532
rect 17631 254501 17661 254527
rect 17841 254501 17871 254532
rect 18051 254501 18081 254527
rect 18261 254501 18291 254532
rect 18471 254501 18501 254527
rect 18681 254501 18711 254532
rect 18891 254501 18921 254527
rect 19101 254501 19131 254532
rect 19311 254501 19341 254527
rect 19521 254501 19551 254532
rect 19731 254501 19761 254527
rect 19941 254501 19971 254532
rect 20151 254501 20181 254527
rect 20361 254501 20391 254532
rect 20571 254501 20601 254527
rect 20781 254501 20811 254532
rect 20991 254501 21021 254527
rect 21201 254501 21231 254532
rect 21411 254501 21441 254527
rect 21621 254501 21651 254532
rect 21831 254501 21861 254527
rect 22041 254501 22071 254532
rect 22251 254501 22281 254527
rect 22461 254501 22491 254532
rect 22671 254501 22701 254527
rect 22881 254501 22911 254532
rect 23091 254501 23121 254527
rect 23301 254501 23331 254532
rect 23511 254501 23541 254527
rect 23721 254501 23751 254532
rect 23931 254501 23961 254527
rect 24141 254501 24171 254532
rect 24351 254501 24381 254527
rect 24561 254501 24591 254532
rect 24771 254501 24801 254527
rect 24981 254501 25011 254532
rect 25191 254501 25221 254527
rect 25401 254501 25431 254532
rect 25611 254501 25641 254527
rect 25821 254501 25851 254532
rect 26031 254501 26061 254527
rect 26241 254501 26271 254532
rect 26451 254501 26481 254527
rect 26661 254501 26691 254532
rect 26871 254501 26901 254527
rect 27081 254501 27111 254532
rect 27291 254501 27321 254527
rect -3999 253675 -3969 253701
rect -3789 253670 -3759 253701
rect -3579 253675 -3549 253701
rect -3369 253670 -3339 253701
rect -3159 253675 -3129 253701
rect -2949 253670 -2919 253701
rect -2739 253675 -2709 253701
rect -2529 253670 -2499 253701
rect -2319 253675 -2289 253701
rect -2109 253670 -2079 253701
rect -1899 253675 -1869 253701
rect -1689 253670 -1659 253701
rect -1479 253675 -1449 253701
rect -1269 253670 -1239 253701
rect -1059 253675 -1029 253701
rect -849 253670 -819 253701
rect -639 253675 -609 253701
rect -429 253670 -399 253701
rect -219 253675 -189 253701
rect -9 253670 21 253701
rect 201 253675 231 253701
rect 411 253670 441 253701
rect 621 253675 651 253701
rect 831 253670 861 253701
rect 1041 253675 1071 253701
rect 1251 253670 1281 253701
rect 1461 253675 1491 253701
rect 1671 253670 1701 253701
rect 1881 253675 1911 253701
rect 2091 253670 2121 253701
rect 2301 253675 2331 253701
rect 2511 253670 2541 253701
rect 2721 253675 2751 253701
rect 2931 253670 2961 253701
rect 3141 253675 3171 253701
rect 3351 253670 3381 253701
rect 3561 253675 3591 253701
rect 3771 253670 3801 253701
rect 3981 253675 4011 253701
rect 4191 253670 4221 253701
rect 4401 253675 4431 253701
rect 4611 253670 4641 253701
rect 4821 253675 4851 253701
rect 5031 253670 5061 253701
rect 5241 253675 5271 253701
rect 5451 253670 5481 253701
rect 5661 253675 5691 253701
rect 5871 253670 5901 253701
rect 6081 253675 6111 253701
rect 6291 253670 6321 253701
rect 6501 253675 6531 253701
rect 6711 253670 6741 253701
rect 6921 253675 6951 253701
rect 7131 253670 7161 253701
rect 7341 253675 7371 253701
rect 7551 253670 7581 253701
rect 7761 253675 7791 253701
rect 7971 253670 8001 253701
rect 8181 253675 8211 253701
rect 8391 253670 8421 253701
rect 8601 253675 8631 253701
rect 8811 253670 8841 253701
rect 9021 253675 9051 253701
rect 9231 253670 9261 253701
rect 9441 253675 9471 253701
rect 9651 253670 9681 253701
rect 9861 253675 9891 253701
rect 10071 253670 10101 253701
rect 10281 253675 10311 253701
rect 10491 253670 10521 253701
rect 10701 253675 10731 253701
rect 10911 253670 10941 253701
rect 11121 253675 11151 253701
rect 11331 253670 11361 253701
rect 11541 253675 11571 253701
rect 11751 253670 11781 253701
rect 11961 253675 11991 253701
rect 12171 253670 12201 253701
rect 12381 253675 12411 253701
rect 12591 253670 12621 253701
rect 12801 253675 12831 253701
rect 13011 253670 13041 253701
rect 13221 253675 13251 253701
rect 13431 253670 13461 253701
rect 13641 253675 13671 253701
rect 13851 253670 13881 253701
rect 14061 253675 14091 253701
rect 14271 253670 14301 253701
rect 14481 253675 14511 253701
rect 14691 253670 14721 253701
rect 14901 253675 14931 253701
rect 15111 253670 15141 253701
rect 15321 253675 15351 253701
rect 15531 253670 15561 253701
rect 15741 253675 15771 253701
rect 15951 253670 15981 253701
rect 16161 253675 16191 253701
rect 16371 253670 16401 253701
rect 16581 253675 16611 253701
rect 16791 253670 16821 253701
rect 17001 253675 17031 253701
rect 17211 253670 17241 253701
rect 17421 253675 17451 253701
rect 17631 253670 17661 253701
rect 17841 253675 17871 253701
rect 18051 253670 18081 253701
rect 18261 253675 18291 253701
rect 18471 253670 18501 253701
rect 18681 253675 18711 253701
rect 18891 253670 18921 253701
rect 19101 253675 19131 253701
rect 19311 253670 19341 253701
rect 19521 253675 19551 253701
rect 19731 253670 19761 253701
rect 19941 253675 19971 253701
rect 20151 253670 20181 253701
rect 20361 253675 20391 253701
rect 20571 253670 20601 253701
rect 20781 253675 20811 253701
rect 20991 253670 21021 253701
rect 21201 253675 21231 253701
rect 21411 253670 21441 253701
rect 21621 253675 21651 253701
rect 21831 253670 21861 253701
rect 22041 253675 22071 253701
rect 22251 253670 22281 253701
rect 22461 253675 22491 253701
rect 22671 253670 22701 253701
rect 22881 253675 22911 253701
rect 23091 253670 23121 253701
rect 23301 253675 23331 253701
rect 23511 253670 23541 253701
rect 23721 253675 23751 253701
rect 23931 253670 23961 253701
rect 24141 253675 24171 253701
rect 24351 253670 24381 253701
rect 24561 253675 24591 253701
rect 24771 253670 24801 253701
rect 24981 253675 25011 253701
rect 25191 253670 25221 253701
rect 25401 253675 25431 253701
rect 25611 253670 25641 253701
rect 25821 253675 25851 253701
rect 26031 253670 26061 253701
rect 26241 253675 26271 253701
rect 26451 253670 26481 253701
rect 26661 253675 26691 253701
rect 26871 253670 26901 253701
rect 27081 253675 27111 253701
rect 27291 253670 27321 253701
rect -3807 253654 -3741 253670
rect -3807 253512 -3791 253654
rect -3757 253512 -3741 253654
rect -3807 253496 -3741 253512
rect -3387 253654 -3321 253670
rect -3387 253512 -3371 253654
rect -3337 253512 -3321 253654
rect -3387 253496 -3321 253512
rect -2967 253654 -2901 253670
rect -2967 253512 -2951 253654
rect -2917 253512 -2901 253654
rect -2967 253496 -2901 253512
rect -2547 253654 -2481 253670
rect -2547 253512 -2531 253654
rect -2497 253512 -2481 253654
rect -2547 253496 -2481 253512
rect -2127 253654 -2061 253670
rect -2127 253512 -2111 253654
rect -2077 253512 -2061 253654
rect -2127 253496 -2061 253512
rect -1707 253654 -1641 253670
rect -1707 253512 -1691 253654
rect -1657 253512 -1641 253654
rect -1707 253496 -1641 253512
rect -1287 253654 -1221 253670
rect -1287 253512 -1271 253654
rect -1237 253512 -1221 253654
rect -1287 253496 -1221 253512
rect -867 253654 -801 253670
rect -867 253512 -851 253654
rect -817 253512 -801 253654
rect -867 253496 -801 253512
rect -447 253654 -381 253670
rect -447 253512 -431 253654
rect -397 253512 -381 253654
rect -447 253496 -381 253512
rect -27 253654 39 253670
rect -27 253512 -11 253654
rect 23 253512 39 253654
rect -27 253496 39 253512
rect 393 253654 459 253670
rect 393 253512 409 253654
rect 443 253512 459 253654
rect 393 253496 459 253512
rect 813 253654 879 253670
rect 813 253512 829 253654
rect 863 253512 879 253654
rect 813 253496 879 253512
rect 1233 253654 1299 253670
rect 1233 253512 1249 253654
rect 1283 253512 1299 253654
rect 1233 253496 1299 253512
rect 1653 253654 1719 253670
rect 1653 253512 1669 253654
rect 1703 253512 1719 253654
rect 1653 253496 1719 253512
rect 2073 253654 2139 253670
rect 2073 253512 2089 253654
rect 2123 253512 2139 253654
rect 2073 253496 2139 253512
rect 2493 253654 2559 253670
rect 2493 253512 2509 253654
rect 2543 253512 2559 253654
rect 2493 253496 2559 253512
rect 2913 253654 2979 253670
rect 2913 253512 2929 253654
rect 2963 253512 2979 253654
rect 2913 253496 2979 253512
rect 3333 253654 3399 253670
rect 3333 253512 3349 253654
rect 3383 253512 3399 253654
rect 3333 253496 3399 253512
rect 3753 253654 3819 253670
rect 3753 253512 3769 253654
rect 3803 253512 3819 253654
rect 3753 253496 3819 253512
rect 4173 253654 4239 253670
rect 4173 253512 4189 253654
rect 4223 253512 4239 253654
rect 4173 253496 4239 253512
rect 4593 253654 4659 253670
rect 4593 253512 4609 253654
rect 4643 253512 4659 253654
rect 4593 253496 4659 253512
rect 5013 253654 5079 253670
rect 5013 253512 5029 253654
rect 5063 253512 5079 253654
rect 5013 253496 5079 253512
rect 5433 253654 5499 253670
rect 5433 253512 5449 253654
rect 5483 253512 5499 253654
rect 5433 253496 5499 253512
rect 5853 253654 5919 253670
rect 5853 253512 5869 253654
rect 5903 253512 5919 253654
rect 5853 253496 5919 253512
rect 6273 253654 6339 253670
rect 6273 253512 6289 253654
rect 6323 253512 6339 253654
rect 6273 253496 6339 253512
rect 6693 253654 6759 253670
rect 6693 253512 6709 253654
rect 6743 253512 6759 253654
rect 6693 253496 6759 253512
rect 7113 253654 7179 253670
rect 7113 253512 7129 253654
rect 7163 253512 7179 253654
rect 7113 253496 7179 253512
rect 7533 253654 7599 253670
rect 7533 253512 7549 253654
rect 7583 253512 7599 253654
rect 7533 253496 7599 253512
rect 7953 253654 8019 253670
rect 7953 253512 7969 253654
rect 8003 253512 8019 253654
rect 7953 253496 8019 253512
rect 8373 253654 8439 253670
rect 8373 253512 8389 253654
rect 8423 253512 8439 253654
rect 8373 253496 8439 253512
rect 8793 253654 8859 253670
rect 8793 253512 8809 253654
rect 8843 253512 8859 253654
rect 8793 253496 8859 253512
rect 9213 253654 9279 253670
rect 9213 253512 9229 253654
rect 9263 253512 9279 253654
rect 9213 253496 9279 253512
rect 9633 253654 9699 253670
rect 9633 253512 9649 253654
rect 9683 253512 9699 253654
rect 9633 253496 9699 253512
rect 10053 253654 10119 253670
rect 10053 253512 10069 253654
rect 10103 253512 10119 253654
rect 10053 253496 10119 253512
rect 10473 253654 10539 253670
rect 10473 253512 10489 253654
rect 10523 253512 10539 253654
rect 10473 253496 10539 253512
rect 10893 253654 10959 253670
rect 10893 253512 10909 253654
rect 10943 253512 10959 253654
rect 10893 253496 10959 253512
rect 11313 253654 11379 253670
rect 11313 253512 11329 253654
rect 11363 253512 11379 253654
rect 11313 253496 11379 253512
rect 11733 253654 11799 253670
rect 11733 253512 11749 253654
rect 11783 253512 11799 253654
rect 11733 253496 11799 253512
rect 12153 253654 12219 253670
rect 12153 253512 12169 253654
rect 12203 253512 12219 253654
rect 12153 253496 12219 253512
rect 12573 253654 12639 253670
rect 12573 253512 12589 253654
rect 12623 253512 12639 253654
rect 12573 253496 12639 253512
rect 12993 253654 13059 253670
rect 12993 253512 13009 253654
rect 13043 253512 13059 253654
rect 12993 253496 13059 253512
rect 13413 253654 13479 253670
rect 13413 253512 13429 253654
rect 13463 253512 13479 253654
rect 13413 253496 13479 253512
rect 13833 253654 13899 253670
rect 13833 253512 13849 253654
rect 13883 253512 13899 253654
rect 13833 253496 13899 253512
rect 14253 253654 14319 253670
rect 14253 253512 14269 253654
rect 14303 253512 14319 253654
rect 14253 253496 14319 253512
rect 14673 253654 14739 253670
rect 14673 253512 14689 253654
rect 14723 253512 14739 253654
rect 14673 253496 14739 253512
rect 15093 253654 15159 253670
rect 15093 253512 15109 253654
rect 15143 253512 15159 253654
rect 15093 253496 15159 253512
rect 15513 253654 15579 253670
rect 15513 253512 15529 253654
rect 15563 253512 15579 253654
rect 15513 253496 15579 253512
rect 15933 253654 15999 253670
rect 15933 253512 15949 253654
rect 15983 253512 15999 253654
rect 15933 253496 15999 253512
rect 16353 253654 16419 253670
rect 16353 253512 16369 253654
rect 16403 253512 16419 253654
rect 16353 253496 16419 253512
rect 16773 253654 16839 253670
rect 16773 253512 16789 253654
rect 16823 253512 16839 253654
rect 16773 253496 16839 253512
rect 17193 253654 17259 253670
rect 17193 253512 17209 253654
rect 17243 253512 17259 253654
rect 17193 253496 17259 253512
rect 17613 253654 17679 253670
rect 17613 253512 17629 253654
rect 17663 253512 17679 253654
rect 17613 253496 17679 253512
rect 18033 253654 18099 253670
rect 18033 253512 18049 253654
rect 18083 253512 18099 253654
rect 18033 253496 18099 253512
rect 18453 253654 18519 253670
rect 18453 253512 18469 253654
rect 18503 253512 18519 253654
rect 18453 253496 18519 253512
rect 18873 253654 18939 253670
rect 18873 253512 18889 253654
rect 18923 253512 18939 253654
rect 18873 253496 18939 253512
rect 19293 253654 19359 253670
rect 19293 253512 19309 253654
rect 19343 253512 19359 253654
rect 19293 253496 19359 253512
rect 19713 253654 19779 253670
rect 19713 253512 19729 253654
rect 19763 253512 19779 253654
rect 19713 253496 19779 253512
rect 20133 253654 20199 253670
rect 20133 253512 20149 253654
rect 20183 253512 20199 253654
rect 20133 253496 20199 253512
rect 20553 253654 20619 253670
rect 20553 253512 20569 253654
rect 20603 253512 20619 253654
rect 20553 253496 20619 253512
rect 20973 253654 21039 253670
rect 20973 253512 20989 253654
rect 21023 253512 21039 253654
rect 20973 253496 21039 253512
rect 21393 253654 21459 253670
rect 21393 253512 21409 253654
rect 21443 253512 21459 253654
rect 21393 253496 21459 253512
rect 21813 253654 21879 253670
rect 21813 253512 21829 253654
rect 21863 253512 21879 253654
rect 21813 253496 21879 253512
rect 22233 253654 22299 253670
rect 22233 253512 22249 253654
rect 22283 253512 22299 253654
rect 22233 253496 22299 253512
rect 22653 253654 22719 253670
rect 22653 253512 22669 253654
rect 22703 253512 22719 253654
rect 22653 253496 22719 253512
rect 23073 253654 23139 253670
rect 23073 253512 23089 253654
rect 23123 253512 23139 253654
rect 23073 253496 23139 253512
rect 23493 253654 23559 253670
rect 23493 253512 23509 253654
rect 23543 253512 23559 253654
rect 23493 253496 23559 253512
rect 23913 253654 23979 253670
rect 23913 253512 23929 253654
rect 23963 253512 23979 253654
rect 23913 253496 23979 253512
rect 24333 253654 24399 253670
rect 24333 253512 24349 253654
rect 24383 253512 24399 253654
rect 24333 253496 24399 253512
rect 24753 253654 24819 253670
rect 24753 253512 24769 253654
rect 24803 253512 24819 253654
rect 24753 253496 24819 253512
rect 25173 253654 25239 253670
rect 25173 253512 25189 253654
rect 25223 253512 25239 253654
rect 25173 253496 25239 253512
rect 25593 253654 25659 253670
rect 25593 253512 25609 253654
rect 25643 253512 25659 253654
rect 25593 253496 25659 253512
rect 26013 253654 26079 253670
rect 26013 253512 26029 253654
rect 26063 253512 26079 253654
rect 26013 253496 26079 253512
rect 26433 253654 26499 253670
rect 26433 253512 26449 253654
rect 26483 253512 26499 253654
rect 26433 253496 26499 253512
rect 26853 253654 26919 253670
rect 26853 253512 26869 253654
rect 26903 253512 26919 253654
rect 26853 253496 26919 253512
rect 27273 253654 27339 253670
rect 27273 253512 27289 253654
rect 27323 253512 27339 253654
rect 27273 253496 27339 253512
rect -3999 253465 -3969 253491
rect -3789 253465 -3759 253496
rect -3579 253465 -3549 253491
rect -3369 253465 -3339 253496
rect -3159 253465 -3129 253491
rect -2949 253465 -2919 253496
rect -2739 253465 -2709 253491
rect -2529 253465 -2499 253496
rect -2319 253465 -2289 253491
rect -2109 253465 -2079 253496
rect -1899 253465 -1869 253491
rect -1689 253465 -1659 253496
rect -1479 253465 -1449 253491
rect -1269 253465 -1239 253496
rect -1059 253465 -1029 253491
rect -849 253465 -819 253496
rect -639 253465 -609 253491
rect -429 253465 -399 253496
rect -219 253465 -189 253491
rect -9 253465 21 253496
rect 201 253465 231 253491
rect 411 253465 441 253496
rect 621 253465 651 253491
rect 831 253465 861 253496
rect 1041 253465 1071 253491
rect 1251 253465 1281 253496
rect 1461 253465 1491 253491
rect 1671 253465 1701 253496
rect 1881 253465 1911 253491
rect 2091 253465 2121 253496
rect 2301 253465 2331 253491
rect 2511 253465 2541 253496
rect 2721 253465 2751 253491
rect 2931 253465 2961 253496
rect 3141 253465 3171 253491
rect 3351 253465 3381 253496
rect 3561 253465 3591 253491
rect 3771 253465 3801 253496
rect 3981 253465 4011 253491
rect 4191 253465 4221 253496
rect 4401 253465 4431 253491
rect 4611 253465 4641 253496
rect 4821 253465 4851 253491
rect 5031 253465 5061 253496
rect 5241 253465 5271 253491
rect 5451 253465 5481 253496
rect 5661 253465 5691 253491
rect 5871 253465 5901 253496
rect 6081 253465 6111 253491
rect 6291 253465 6321 253496
rect 6501 253465 6531 253491
rect 6711 253465 6741 253496
rect 6921 253465 6951 253491
rect 7131 253465 7161 253496
rect 7341 253465 7371 253491
rect 7551 253465 7581 253496
rect 7761 253465 7791 253491
rect 7971 253465 8001 253496
rect 8181 253465 8211 253491
rect 8391 253465 8421 253496
rect 8601 253465 8631 253491
rect 8811 253465 8841 253496
rect 9021 253465 9051 253491
rect 9231 253465 9261 253496
rect 9441 253465 9471 253491
rect 9651 253465 9681 253496
rect 9861 253465 9891 253491
rect 10071 253465 10101 253496
rect 10281 253465 10311 253491
rect 10491 253465 10521 253496
rect 10701 253465 10731 253491
rect 10911 253465 10941 253496
rect 11121 253465 11151 253491
rect 11331 253465 11361 253496
rect 11541 253465 11571 253491
rect 11751 253465 11781 253496
rect 11961 253465 11991 253491
rect 12171 253465 12201 253496
rect 12381 253465 12411 253491
rect 12591 253465 12621 253496
rect 12801 253465 12831 253491
rect 13011 253465 13041 253496
rect 13221 253465 13251 253491
rect 13431 253465 13461 253496
rect 13641 253465 13671 253491
rect 13851 253465 13881 253496
rect 14061 253465 14091 253491
rect 14271 253465 14301 253496
rect 14481 253465 14511 253491
rect 14691 253465 14721 253496
rect 14901 253465 14931 253491
rect 15111 253465 15141 253496
rect 15321 253465 15351 253491
rect 15531 253465 15561 253496
rect 15741 253465 15771 253491
rect 15951 253465 15981 253496
rect 16161 253465 16191 253491
rect 16371 253465 16401 253496
rect 16581 253465 16611 253491
rect 16791 253465 16821 253496
rect 17001 253465 17031 253491
rect 17211 253465 17241 253496
rect 17421 253465 17451 253491
rect 17631 253465 17661 253496
rect 17841 253465 17871 253491
rect 18051 253465 18081 253496
rect 18261 253465 18291 253491
rect 18471 253465 18501 253496
rect 18681 253465 18711 253491
rect 18891 253465 18921 253496
rect 19101 253465 19131 253491
rect 19311 253465 19341 253496
rect 19521 253465 19551 253491
rect 19731 253465 19761 253496
rect 19941 253465 19971 253491
rect 20151 253465 20181 253496
rect 20361 253465 20391 253491
rect 20571 253465 20601 253496
rect 20781 253465 20811 253491
rect 20991 253465 21021 253496
rect 21201 253465 21231 253491
rect 21411 253465 21441 253496
rect 21621 253465 21651 253491
rect 21831 253465 21861 253496
rect 22041 253465 22071 253491
rect 22251 253465 22281 253496
rect 22461 253465 22491 253491
rect 22671 253465 22701 253496
rect 22881 253465 22911 253491
rect 23091 253465 23121 253496
rect 23301 253465 23331 253491
rect 23511 253465 23541 253496
rect 23721 253465 23751 253491
rect 23931 253465 23961 253496
rect 24141 253465 24171 253491
rect 24351 253465 24381 253496
rect 24561 253465 24591 253491
rect 24771 253465 24801 253496
rect 24981 253465 25011 253491
rect 25191 253465 25221 253496
rect 25401 253465 25431 253491
rect 25611 253465 25641 253496
rect 25821 253465 25851 253491
rect 26031 253465 26061 253496
rect 26241 253465 26271 253491
rect 26451 253465 26481 253496
rect 26661 253465 26691 253491
rect 26871 253465 26901 253496
rect 27081 253465 27111 253491
rect 27291 253465 27321 253496
rect -3999 252634 -3969 252665
rect -3789 252639 -3759 252665
rect -3579 252634 -3549 252665
rect -3369 252639 -3339 252665
rect -3159 252634 -3129 252665
rect -2949 252639 -2919 252665
rect -2739 252634 -2709 252665
rect -2529 252639 -2499 252665
rect -2319 252634 -2289 252665
rect -2109 252639 -2079 252665
rect -1899 252634 -1869 252665
rect -1689 252639 -1659 252665
rect -1479 252634 -1449 252665
rect -1269 252639 -1239 252665
rect -1059 252634 -1029 252665
rect -849 252639 -819 252665
rect -639 252634 -609 252665
rect -429 252639 -399 252665
rect -219 252634 -189 252665
rect -9 252639 21 252665
rect 201 252634 231 252665
rect 411 252639 441 252665
rect 621 252634 651 252665
rect 831 252639 861 252665
rect 1041 252634 1071 252665
rect 1251 252639 1281 252665
rect 1461 252634 1491 252665
rect 1671 252639 1701 252665
rect 1881 252634 1911 252665
rect 2091 252639 2121 252665
rect 2301 252634 2331 252665
rect 2511 252639 2541 252665
rect 2721 252634 2751 252665
rect 2931 252639 2961 252665
rect 3141 252634 3171 252665
rect 3351 252639 3381 252665
rect 3561 252634 3591 252665
rect 3771 252639 3801 252665
rect 3981 252634 4011 252665
rect 4191 252639 4221 252665
rect 4401 252634 4431 252665
rect 4611 252639 4641 252665
rect 4821 252634 4851 252665
rect 5031 252639 5061 252665
rect 5241 252634 5271 252665
rect 5451 252639 5481 252665
rect 5661 252634 5691 252665
rect 5871 252639 5901 252665
rect 6081 252634 6111 252665
rect 6291 252639 6321 252665
rect 6501 252634 6531 252665
rect 6711 252639 6741 252665
rect 6921 252634 6951 252665
rect 7131 252639 7161 252665
rect 7341 252634 7371 252665
rect 7551 252639 7581 252665
rect 7761 252634 7791 252665
rect 7971 252639 8001 252665
rect 8181 252634 8211 252665
rect 8391 252639 8421 252665
rect 8601 252634 8631 252665
rect 8811 252639 8841 252665
rect 9021 252634 9051 252665
rect 9231 252639 9261 252665
rect 9441 252634 9471 252665
rect 9651 252639 9681 252665
rect 9861 252634 9891 252665
rect 10071 252639 10101 252665
rect 10281 252634 10311 252665
rect 10491 252639 10521 252665
rect 10701 252634 10731 252665
rect 10911 252639 10941 252665
rect 11121 252634 11151 252665
rect 11331 252639 11361 252665
rect 11541 252634 11571 252665
rect 11751 252639 11781 252665
rect 11961 252634 11991 252665
rect 12171 252639 12201 252665
rect 12381 252634 12411 252665
rect 12591 252639 12621 252665
rect 12801 252634 12831 252665
rect 13011 252639 13041 252665
rect 13221 252634 13251 252665
rect 13431 252639 13461 252665
rect 13641 252634 13671 252665
rect 13851 252639 13881 252665
rect 14061 252634 14091 252665
rect 14271 252639 14301 252665
rect 14481 252634 14511 252665
rect 14691 252639 14721 252665
rect 14901 252634 14931 252665
rect 15111 252639 15141 252665
rect 15321 252634 15351 252665
rect 15531 252639 15561 252665
rect 15741 252634 15771 252665
rect 15951 252639 15981 252665
rect 16161 252634 16191 252665
rect 16371 252639 16401 252665
rect 16581 252634 16611 252665
rect 16791 252639 16821 252665
rect 17001 252634 17031 252665
rect 17211 252639 17241 252665
rect 17421 252634 17451 252665
rect 17631 252639 17661 252665
rect 17841 252634 17871 252665
rect 18051 252639 18081 252665
rect 18261 252634 18291 252665
rect 18471 252639 18501 252665
rect 18681 252634 18711 252665
rect 18891 252639 18921 252665
rect 19101 252634 19131 252665
rect 19311 252639 19341 252665
rect 19521 252634 19551 252665
rect 19731 252639 19761 252665
rect 19941 252634 19971 252665
rect 20151 252639 20181 252665
rect 20361 252634 20391 252665
rect 20571 252639 20601 252665
rect 20781 252634 20811 252665
rect 20991 252639 21021 252665
rect 21201 252634 21231 252665
rect 21411 252639 21441 252665
rect 21621 252634 21651 252665
rect 21831 252639 21861 252665
rect 22041 252634 22071 252665
rect 22251 252639 22281 252665
rect 22461 252634 22491 252665
rect 22671 252639 22701 252665
rect 22881 252634 22911 252665
rect 23091 252639 23121 252665
rect 23301 252634 23331 252665
rect 23511 252639 23541 252665
rect 23721 252634 23751 252665
rect 23931 252639 23961 252665
rect 24141 252634 24171 252665
rect 24351 252639 24381 252665
rect 24561 252634 24591 252665
rect 24771 252639 24801 252665
rect 24981 252634 25011 252665
rect 25191 252639 25221 252665
rect 25401 252634 25431 252665
rect 25611 252639 25641 252665
rect 25821 252634 25851 252665
rect 26031 252639 26061 252665
rect 26241 252634 26271 252665
rect 26451 252639 26481 252665
rect 26661 252634 26691 252665
rect 26871 252639 26901 252665
rect 27081 252634 27111 252665
rect 27291 252639 27321 252665
rect -4017 252618 -3951 252634
rect -4017 252476 -4001 252618
rect -3967 252476 -3951 252618
rect -4017 252460 -3951 252476
rect -3597 252618 -3531 252634
rect -3597 252476 -3581 252618
rect -3547 252476 -3531 252618
rect -3597 252460 -3531 252476
rect -3177 252618 -3111 252634
rect -3177 252476 -3161 252618
rect -3127 252476 -3111 252618
rect -3177 252460 -3111 252476
rect -2757 252618 -2691 252634
rect -2757 252476 -2741 252618
rect -2707 252476 -2691 252618
rect -2757 252460 -2691 252476
rect -2337 252618 -2271 252634
rect -2337 252476 -2321 252618
rect -2287 252476 -2271 252618
rect -2337 252460 -2271 252476
rect -1917 252618 -1851 252634
rect -1917 252476 -1901 252618
rect -1867 252476 -1851 252618
rect -1917 252460 -1851 252476
rect -1497 252618 -1431 252634
rect -1497 252476 -1481 252618
rect -1447 252476 -1431 252618
rect -1497 252460 -1431 252476
rect -1077 252618 -1011 252634
rect -1077 252476 -1061 252618
rect -1027 252476 -1011 252618
rect -1077 252460 -1011 252476
rect -657 252618 -591 252634
rect -657 252476 -641 252618
rect -607 252476 -591 252618
rect -657 252460 -591 252476
rect -237 252618 -171 252634
rect -237 252476 -221 252618
rect -187 252476 -171 252618
rect -237 252460 -171 252476
rect 183 252618 249 252634
rect 183 252476 199 252618
rect 233 252476 249 252618
rect 183 252460 249 252476
rect 603 252618 669 252634
rect 603 252476 619 252618
rect 653 252476 669 252618
rect 603 252460 669 252476
rect 1023 252618 1089 252634
rect 1023 252476 1039 252618
rect 1073 252476 1089 252618
rect 1023 252460 1089 252476
rect 1443 252618 1509 252634
rect 1443 252476 1459 252618
rect 1493 252476 1509 252618
rect 1443 252460 1509 252476
rect 1863 252618 1929 252634
rect 1863 252476 1879 252618
rect 1913 252476 1929 252618
rect 1863 252460 1929 252476
rect 2283 252618 2349 252634
rect 2283 252476 2299 252618
rect 2333 252476 2349 252618
rect 2283 252460 2349 252476
rect 2703 252618 2769 252634
rect 2703 252476 2719 252618
rect 2753 252476 2769 252618
rect 2703 252460 2769 252476
rect 3123 252618 3189 252634
rect 3123 252476 3139 252618
rect 3173 252476 3189 252618
rect 3123 252460 3189 252476
rect 3543 252618 3609 252634
rect 3543 252476 3559 252618
rect 3593 252476 3609 252618
rect 3543 252460 3609 252476
rect 3963 252618 4029 252634
rect 3963 252476 3979 252618
rect 4013 252476 4029 252618
rect 3963 252460 4029 252476
rect 4383 252618 4449 252634
rect 4383 252476 4399 252618
rect 4433 252476 4449 252618
rect 4383 252460 4449 252476
rect 4803 252618 4869 252634
rect 4803 252476 4819 252618
rect 4853 252476 4869 252618
rect 4803 252460 4869 252476
rect 5223 252618 5289 252634
rect 5223 252476 5239 252618
rect 5273 252476 5289 252618
rect 5223 252460 5289 252476
rect 5643 252618 5709 252634
rect 5643 252476 5659 252618
rect 5693 252476 5709 252618
rect 5643 252460 5709 252476
rect 6063 252618 6129 252634
rect 6063 252476 6079 252618
rect 6113 252476 6129 252618
rect 6063 252460 6129 252476
rect 6483 252618 6549 252634
rect 6483 252476 6499 252618
rect 6533 252476 6549 252618
rect 6483 252460 6549 252476
rect 6903 252618 6969 252634
rect 6903 252476 6919 252618
rect 6953 252476 6969 252618
rect 6903 252460 6969 252476
rect 7323 252618 7389 252634
rect 7323 252476 7339 252618
rect 7373 252476 7389 252618
rect 7323 252460 7389 252476
rect 7743 252618 7809 252634
rect 7743 252476 7759 252618
rect 7793 252476 7809 252618
rect 7743 252460 7809 252476
rect 8163 252618 8229 252634
rect 8163 252476 8179 252618
rect 8213 252476 8229 252618
rect 8163 252460 8229 252476
rect 8583 252618 8649 252634
rect 8583 252476 8599 252618
rect 8633 252476 8649 252618
rect 8583 252460 8649 252476
rect 9003 252618 9069 252634
rect 9003 252476 9019 252618
rect 9053 252476 9069 252618
rect 9003 252460 9069 252476
rect 9423 252618 9489 252634
rect 9423 252476 9439 252618
rect 9473 252476 9489 252618
rect 9423 252460 9489 252476
rect 9843 252618 9909 252634
rect 9843 252476 9859 252618
rect 9893 252476 9909 252618
rect 9843 252460 9909 252476
rect 10263 252618 10329 252634
rect 10263 252476 10279 252618
rect 10313 252476 10329 252618
rect 10263 252460 10329 252476
rect 10683 252618 10749 252634
rect 10683 252476 10699 252618
rect 10733 252476 10749 252618
rect 10683 252460 10749 252476
rect 11103 252618 11169 252634
rect 11103 252476 11119 252618
rect 11153 252476 11169 252618
rect 11103 252460 11169 252476
rect 11523 252618 11589 252634
rect 11523 252476 11539 252618
rect 11573 252476 11589 252618
rect 11523 252460 11589 252476
rect 11943 252618 12009 252634
rect 11943 252476 11959 252618
rect 11993 252476 12009 252618
rect 11943 252460 12009 252476
rect 12363 252618 12429 252634
rect 12363 252476 12379 252618
rect 12413 252476 12429 252618
rect 12363 252460 12429 252476
rect 12783 252618 12849 252634
rect 12783 252476 12799 252618
rect 12833 252476 12849 252618
rect 12783 252460 12849 252476
rect 13203 252618 13269 252634
rect 13203 252476 13219 252618
rect 13253 252476 13269 252618
rect 13203 252460 13269 252476
rect 13623 252618 13689 252634
rect 13623 252476 13639 252618
rect 13673 252476 13689 252618
rect 13623 252460 13689 252476
rect 14043 252618 14109 252634
rect 14043 252476 14059 252618
rect 14093 252476 14109 252618
rect 14043 252460 14109 252476
rect 14463 252618 14529 252634
rect 14463 252476 14479 252618
rect 14513 252476 14529 252618
rect 14463 252460 14529 252476
rect 14883 252618 14949 252634
rect 14883 252476 14899 252618
rect 14933 252476 14949 252618
rect 14883 252460 14949 252476
rect 15303 252618 15369 252634
rect 15303 252476 15319 252618
rect 15353 252476 15369 252618
rect 15303 252460 15369 252476
rect 15723 252618 15789 252634
rect 15723 252476 15739 252618
rect 15773 252476 15789 252618
rect 15723 252460 15789 252476
rect 16143 252618 16209 252634
rect 16143 252476 16159 252618
rect 16193 252476 16209 252618
rect 16143 252460 16209 252476
rect 16563 252618 16629 252634
rect 16563 252476 16579 252618
rect 16613 252476 16629 252618
rect 16563 252460 16629 252476
rect 16983 252618 17049 252634
rect 16983 252476 16999 252618
rect 17033 252476 17049 252618
rect 16983 252460 17049 252476
rect 17403 252618 17469 252634
rect 17403 252476 17419 252618
rect 17453 252476 17469 252618
rect 17403 252460 17469 252476
rect 17823 252618 17889 252634
rect 17823 252476 17839 252618
rect 17873 252476 17889 252618
rect 17823 252460 17889 252476
rect 18243 252618 18309 252634
rect 18243 252476 18259 252618
rect 18293 252476 18309 252618
rect 18243 252460 18309 252476
rect 18663 252618 18729 252634
rect 18663 252476 18679 252618
rect 18713 252476 18729 252618
rect 18663 252460 18729 252476
rect 19083 252618 19149 252634
rect 19083 252476 19099 252618
rect 19133 252476 19149 252618
rect 19083 252460 19149 252476
rect 19503 252618 19569 252634
rect 19503 252476 19519 252618
rect 19553 252476 19569 252618
rect 19503 252460 19569 252476
rect 19923 252618 19989 252634
rect 19923 252476 19939 252618
rect 19973 252476 19989 252618
rect 19923 252460 19989 252476
rect 20343 252618 20409 252634
rect 20343 252476 20359 252618
rect 20393 252476 20409 252618
rect 20343 252460 20409 252476
rect 20763 252618 20829 252634
rect 20763 252476 20779 252618
rect 20813 252476 20829 252618
rect 20763 252460 20829 252476
rect 21183 252618 21249 252634
rect 21183 252476 21199 252618
rect 21233 252476 21249 252618
rect 21183 252460 21249 252476
rect 21603 252618 21669 252634
rect 21603 252476 21619 252618
rect 21653 252476 21669 252618
rect 21603 252460 21669 252476
rect 22023 252618 22089 252634
rect 22023 252476 22039 252618
rect 22073 252476 22089 252618
rect 22023 252460 22089 252476
rect 22443 252618 22509 252634
rect 22443 252476 22459 252618
rect 22493 252476 22509 252618
rect 22443 252460 22509 252476
rect 22863 252618 22929 252634
rect 22863 252476 22879 252618
rect 22913 252476 22929 252618
rect 22863 252460 22929 252476
rect 23283 252618 23349 252634
rect 23283 252476 23299 252618
rect 23333 252476 23349 252618
rect 23283 252460 23349 252476
rect 23703 252618 23769 252634
rect 23703 252476 23719 252618
rect 23753 252476 23769 252618
rect 23703 252460 23769 252476
rect 24123 252618 24189 252634
rect 24123 252476 24139 252618
rect 24173 252476 24189 252618
rect 24123 252460 24189 252476
rect 24543 252618 24609 252634
rect 24543 252476 24559 252618
rect 24593 252476 24609 252618
rect 24543 252460 24609 252476
rect 24963 252618 25029 252634
rect 24963 252476 24979 252618
rect 25013 252476 25029 252618
rect 24963 252460 25029 252476
rect 25383 252618 25449 252634
rect 25383 252476 25399 252618
rect 25433 252476 25449 252618
rect 25383 252460 25449 252476
rect 25803 252618 25869 252634
rect 25803 252476 25819 252618
rect 25853 252476 25869 252618
rect 25803 252460 25869 252476
rect 26223 252618 26289 252634
rect 26223 252476 26239 252618
rect 26273 252476 26289 252618
rect 26223 252460 26289 252476
rect 26643 252618 26709 252634
rect 26643 252476 26659 252618
rect 26693 252476 26709 252618
rect 26643 252460 26709 252476
rect 27063 252618 27129 252634
rect 27063 252476 27079 252618
rect 27113 252476 27129 252618
rect 27063 252460 27129 252476
rect -3999 252429 -3969 252460
rect -3789 252429 -3759 252455
rect -3579 252429 -3549 252460
rect -3369 252429 -3339 252455
rect -3159 252429 -3129 252460
rect -2949 252429 -2919 252455
rect -2739 252429 -2709 252460
rect -2529 252429 -2499 252455
rect -2319 252429 -2289 252460
rect -2109 252429 -2079 252455
rect -1899 252429 -1869 252460
rect -1689 252429 -1659 252455
rect -1479 252429 -1449 252460
rect -1269 252429 -1239 252455
rect -1059 252429 -1029 252460
rect -849 252429 -819 252455
rect -639 252429 -609 252460
rect -429 252429 -399 252455
rect -219 252429 -189 252460
rect -9 252429 21 252455
rect 201 252429 231 252460
rect 411 252429 441 252455
rect 621 252429 651 252460
rect 831 252429 861 252455
rect 1041 252429 1071 252460
rect 1251 252429 1281 252455
rect 1461 252429 1491 252460
rect 1671 252429 1701 252455
rect 1881 252429 1911 252460
rect 2091 252429 2121 252455
rect 2301 252429 2331 252460
rect 2511 252429 2541 252455
rect 2721 252429 2751 252460
rect 2931 252429 2961 252455
rect 3141 252429 3171 252460
rect 3351 252429 3381 252455
rect 3561 252429 3591 252460
rect 3771 252429 3801 252455
rect 3981 252429 4011 252460
rect 4191 252429 4221 252455
rect 4401 252429 4431 252460
rect 4611 252429 4641 252455
rect 4821 252429 4851 252460
rect 5031 252429 5061 252455
rect 5241 252429 5271 252460
rect 5451 252429 5481 252455
rect 5661 252429 5691 252460
rect 5871 252429 5901 252455
rect 6081 252429 6111 252460
rect 6291 252429 6321 252455
rect 6501 252429 6531 252460
rect 6711 252429 6741 252455
rect 6921 252429 6951 252460
rect 7131 252429 7161 252455
rect 7341 252429 7371 252460
rect 7551 252429 7581 252455
rect 7761 252429 7791 252460
rect 7971 252429 8001 252455
rect 8181 252429 8211 252460
rect 8391 252429 8421 252455
rect 8601 252429 8631 252460
rect 8811 252429 8841 252455
rect 9021 252429 9051 252460
rect 9231 252429 9261 252455
rect 9441 252429 9471 252460
rect 9651 252429 9681 252455
rect 9861 252429 9891 252460
rect 10071 252429 10101 252455
rect 10281 252429 10311 252460
rect 10491 252429 10521 252455
rect 10701 252429 10731 252460
rect 10911 252429 10941 252455
rect 11121 252429 11151 252460
rect 11331 252429 11361 252455
rect 11541 252429 11571 252460
rect 11751 252429 11781 252455
rect 11961 252429 11991 252460
rect 12171 252429 12201 252455
rect 12381 252429 12411 252460
rect 12591 252429 12621 252455
rect 12801 252429 12831 252460
rect 13011 252429 13041 252455
rect 13221 252429 13251 252460
rect 13431 252429 13461 252455
rect 13641 252429 13671 252460
rect 13851 252429 13881 252455
rect 14061 252429 14091 252460
rect 14271 252429 14301 252455
rect 14481 252429 14511 252460
rect 14691 252429 14721 252455
rect 14901 252429 14931 252460
rect 15111 252429 15141 252455
rect 15321 252429 15351 252460
rect 15531 252429 15561 252455
rect 15741 252429 15771 252460
rect 15951 252429 15981 252455
rect 16161 252429 16191 252460
rect 16371 252429 16401 252455
rect 16581 252429 16611 252460
rect 16791 252429 16821 252455
rect 17001 252429 17031 252460
rect 17211 252429 17241 252455
rect 17421 252429 17451 252460
rect 17631 252429 17661 252455
rect 17841 252429 17871 252460
rect 18051 252429 18081 252455
rect 18261 252429 18291 252460
rect 18471 252429 18501 252455
rect 18681 252429 18711 252460
rect 18891 252429 18921 252455
rect 19101 252429 19131 252460
rect 19311 252429 19341 252455
rect 19521 252429 19551 252460
rect 19731 252429 19761 252455
rect 19941 252429 19971 252460
rect 20151 252429 20181 252455
rect 20361 252429 20391 252460
rect 20571 252429 20601 252455
rect 20781 252429 20811 252460
rect 20991 252429 21021 252455
rect 21201 252429 21231 252460
rect 21411 252429 21441 252455
rect 21621 252429 21651 252460
rect 21831 252429 21861 252455
rect 22041 252429 22071 252460
rect 22251 252429 22281 252455
rect 22461 252429 22491 252460
rect 22671 252429 22701 252455
rect 22881 252429 22911 252460
rect 23091 252429 23121 252455
rect 23301 252429 23331 252460
rect 23511 252429 23541 252455
rect 23721 252429 23751 252460
rect 23931 252429 23961 252455
rect 24141 252429 24171 252460
rect 24351 252429 24381 252455
rect 24561 252429 24591 252460
rect 24771 252429 24801 252455
rect 24981 252429 25011 252460
rect 25191 252429 25221 252455
rect 25401 252429 25431 252460
rect 25611 252429 25641 252455
rect 25821 252429 25851 252460
rect 26031 252429 26061 252455
rect 26241 252429 26271 252460
rect 26451 252429 26481 252455
rect 26661 252429 26691 252460
rect 26871 252429 26901 252455
rect 27081 252429 27111 252460
rect 27291 252429 27321 252455
rect -3999 251603 -3969 251629
rect -3789 251598 -3759 251629
rect -3579 251603 -3549 251629
rect -3369 251598 -3339 251629
rect -3159 251603 -3129 251629
rect -2949 251598 -2919 251629
rect -2739 251603 -2709 251629
rect -2529 251598 -2499 251629
rect -2319 251603 -2289 251629
rect -2109 251598 -2079 251629
rect -1899 251603 -1869 251629
rect -1689 251598 -1659 251629
rect -1479 251603 -1449 251629
rect -1269 251598 -1239 251629
rect -1059 251603 -1029 251629
rect -849 251598 -819 251629
rect -639 251603 -609 251629
rect -429 251598 -399 251629
rect -219 251603 -189 251629
rect -9 251598 21 251629
rect 201 251603 231 251629
rect 411 251598 441 251629
rect 621 251603 651 251629
rect 831 251598 861 251629
rect 1041 251603 1071 251629
rect 1251 251598 1281 251629
rect 1461 251603 1491 251629
rect 1671 251598 1701 251629
rect 1881 251603 1911 251629
rect 2091 251598 2121 251629
rect 2301 251603 2331 251629
rect 2511 251598 2541 251629
rect 2721 251603 2751 251629
rect 2931 251598 2961 251629
rect 3141 251603 3171 251629
rect 3351 251598 3381 251629
rect 3561 251603 3591 251629
rect 3771 251598 3801 251629
rect 3981 251603 4011 251629
rect 4191 251598 4221 251629
rect 4401 251603 4431 251629
rect 4611 251598 4641 251629
rect 4821 251603 4851 251629
rect 5031 251598 5061 251629
rect 5241 251603 5271 251629
rect 5451 251598 5481 251629
rect 5661 251603 5691 251629
rect 5871 251598 5901 251629
rect 6081 251603 6111 251629
rect 6291 251598 6321 251629
rect 6501 251603 6531 251629
rect 6711 251598 6741 251629
rect 6921 251603 6951 251629
rect 7131 251598 7161 251629
rect 7341 251603 7371 251629
rect 7551 251598 7581 251629
rect 7761 251603 7791 251629
rect 7971 251598 8001 251629
rect 8181 251603 8211 251629
rect 8391 251598 8421 251629
rect 8601 251603 8631 251629
rect 8811 251598 8841 251629
rect 9021 251603 9051 251629
rect 9231 251598 9261 251629
rect 9441 251603 9471 251629
rect 9651 251598 9681 251629
rect 9861 251603 9891 251629
rect 10071 251598 10101 251629
rect 10281 251603 10311 251629
rect 10491 251598 10521 251629
rect 10701 251603 10731 251629
rect 10911 251598 10941 251629
rect 11121 251603 11151 251629
rect 11331 251598 11361 251629
rect 11541 251603 11571 251629
rect 11751 251598 11781 251629
rect 11961 251603 11991 251629
rect 12171 251598 12201 251629
rect 12381 251603 12411 251629
rect 12591 251598 12621 251629
rect 12801 251603 12831 251629
rect 13011 251598 13041 251629
rect 13221 251603 13251 251629
rect 13431 251598 13461 251629
rect 13641 251603 13671 251629
rect 13851 251598 13881 251629
rect 14061 251603 14091 251629
rect 14271 251598 14301 251629
rect 14481 251603 14511 251629
rect 14691 251598 14721 251629
rect 14901 251603 14931 251629
rect 15111 251598 15141 251629
rect 15321 251603 15351 251629
rect 15531 251598 15561 251629
rect 15741 251603 15771 251629
rect 15951 251598 15981 251629
rect 16161 251603 16191 251629
rect 16371 251598 16401 251629
rect 16581 251603 16611 251629
rect 16791 251598 16821 251629
rect 17001 251603 17031 251629
rect 17211 251598 17241 251629
rect 17421 251603 17451 251629
rect 17631 251598 17661 251629
rect 17841 251603 17871 251629
rect 18051 251598 18081 251629
rect 18261 251603 18291 251629
rect 18471 251598 18501 251629
rect 18681 251603 18711 251629
rect 18891 251598 18921 251629
rect 19101 251603 19131 251629
rect 19311 251598 19341 251629
rect 19521 251603 19551 251629
rect 19731 251598 19761 251629
rect 19941 251603 19971 251629
rect 20151 251598 20181 251629
rect 20361 251603 20391 251629
rect 20571 251598 20601 251629
rect 20781 251603 20811 251629
rect 20991 251598 21021 251629
rect 21201 251603 21231 251629
rect 21411 251598 21441 251629
rect 21621 251603 21651 251629
rect 21831 251598 21861 251629
rect 22041 251603 22071 251629
rect 22251 251598 22281 251629
rect 22461 251603 22491 251629
rect 22671 251598 22701 251629
rect 22881 251603 22911 251629
rect 23091 251598 23121 251629
rect 23301 251603 23331 251629
rect 23511 251598 23541 251629
rect 23721 251603 23751 251629
rect 23931 251598 23961 251629
rect 24141 251603 24171 251629
rect 24351 251598 24381 251629
rect 24561 251603 24591 251629
rect 24771 251598 24801 251629
rect 24981 251603 25011 251629
rect 25191 251598 25221 251629
rect 25401 251603 25431 251629
rect 25611 251598 25641 251629
rect 25821 251603 25851 251629
rect 26031 251598 26061 251629
rect 26241 251603 26271 251629
rect 26451 251598 26481 251629
rect 26661 251603 26691 251629
rect 26871 251598 26901 251629
rect 27081 251603 27111 251629
rect 27291 251598 27321 251629
rect -3807 251582 -3741 251598
rect -3807 251440 -3791 251582
rect -3757 251440 -3741 251582
rect -3807 251424 -3741 251440
rect -3387 251582 -3321 251598
rect -3387 251440 -3371 251582
rect -3337 251440 -3321 251582
rect -3387 251424 -3321 251440
rect -2967 251582 -2901 251598
rect -2967 251440 -2951 251582
rect -2917 251440 -2901 251582
rect -2967 251424 -2901 251440
rect -2547 251582 -2481 251598
rect -2547 251440 -2531 251582
rect -2497 251440 -2481 251582
rect -2547 251424 -2481 251440
rect -2127 251582 -2061 251598
rect -2127 251440 -2111 251582
rect -2077 251440 -2061 251582
rect -2127 251424 -2061 251440
rect -1707 251582 -1641 251598
rect -1707 251440 -1691 251582
rect -1657 251440 -1641 251582
rect -1707 251424 -1641 251440
rect -1287 251582 -1221 251598
rect -1287 251440 -1271 251582
rect -1237 251440 -1221 251582
rect -1287 251424 -1221 251440
rect -867 251582 -801 251598
rect -867 251440 -851 251582
rect -817 251440 -801 251582
rect -867 251424 -801 251440
rect -447 251582 -381 251598
rect -447 251440 -431 251582
rect -397 251440 -381 251582
rect -447 251424 -381 251440
rect -27 251582 39 251598
rect -27 251440 -11 251582
rect 23 251440 39 251582
rect -27 251424 39 251440
rect 393 251582 459 251598
rect 393 251440 409 251582
rect 443 251440 459 251582
rect 393 251424 459 251440
rect 813 251582 879 251598
rect 813 251440 829 251582
rect 863 251440 879 251582
rect 813 251424 879 251440
rect 1233 251582 1299 251598
rect 1233 251440 1249 251582
rect 1283 251440 1299 251582
rect 1233 251424 1299 251440
rect 1653 251582 1719 251598
rect 1653 251440 1669 251582
rect 1703 251440 1719 251582
rect 1653 251424 1719 251440
rect 2073 251582 2139 251598
rect 2073 251440 2089 251582
rect 2123 251440 2139 251582
rect 2073 251424 2139 251440
rect 2493 251582 2559 251598
rect 2493 251440 2509 251582
rect 2543 251440 2559 251582
rect 2493 251424 2559 251440
rect 2913 251582 2979 251598
rect 2913 251440 2929 251582
rect 2963 251440 2979 251582
rect 2913 251424 2979 251440
rect 3333 251582 3399 251598
rect 3333 251440 3349 251582
rect 3383 251440 3399 251582
rect 3333 251424 3399 251440
rect 3753 251582 3819 251598
rect 3753 251440 3769 251582
rect 3803 251440 3819 251582
rect 3753 251424 3819 251440
rect 4173 251582 4239 251598
rect 4173 251440 4189 251582
rect 4223 251440 4239 251582
rect 4173 251424 4239 251440
rect 4593 251582 4659 251598
rect 4593 251440 4609 251582
rect 4643 251440 4659 251582
rect 4593 251424 4659 251440
rect 5013 251582 5079 251598
rect 5013 251440 5029 251582
rect 5063 251440 5079 251582
rect 5013 251424 5079 251440
rect 5433 251582 5499 251598
rect 5433 251440 5449 251582
rect 5483 251440 5499 251582
rect 5433 251424 5499 251440
rect 5853 251582 5919 251598
rect 5853 251440 5869 251582
rect 5903 251440 5919 251582
rect 5853 251424 5919 251440
rect 6273 251582 6339 251598
rect 6273 251440 6289 251582
rect 6323 251440 6339 251582
rect 6273 251424 6339 251440
rect 6693 251582 6759 251598
rect 6693 251440 6709 251582
rect 6743 251440 6759 251582
rect 6693 251424 6759 251440
rect 7113 251582 7179 251598
rect 7113 251440 7129 251582
rect 7163 251440 7179 251582
rect 7113 251424 7179 251440
rect 7533 251582 7599 251598
rect 7533 251440 7549 251582
rect 7583 251440 7599 251582
rect 7533 251424 7599 251440
rect 7953 251582 8019 251598
rect 7953 251440 7969 251582
rect 8003 251440 8019 251582
rect 7953 251424 8019 251440
rect 8373 251582 8439 251598
rect 8373 251440 8389 251582
rect 8423 251440 8439 251582
rect 8373 251424 8439 251440
rect 8793 251582 8859 251598
rect 8793 251440 8809 251582
rect 8843 251440 8859 251582
rect 8793 251424 8859 251440
rect 9213 251582 9279 251598
rect 9213 251440 9229 251582
rect 9263 251440 9279 251582
rect 9213 251424 9279 251440
rect 9633 251582 9699 251598
rect 9633 251440 9649 251582
rect 9683 251440 9699 251582
rect 9633 251424 9699 251440
rect 10053 251582 10119 251598
rect 10053 251440 10069 251582
rect 10103 251440 10119 251582
rect 10053 251424 10119 251440
rect 10473 251582 10539 251598
rect 10473 251440 10489 251582
rect 10523 251440 10539 251582
rect 10473 251424 10539 251440
rect 10893 251582 10959 251598
rect 10893 251440 10909 251582
rect 10943 251440 10959 251582
rect 10893 251424 10959 251440
rect 11313 251582 11379 251598
rect 11313 251440 11329 251582
rect 11363 251440 11379 251582
rect 11313 251424 11379 251440
rect 11733 251582 11799 251598
rect 11733 251440 11749 251582
rect 11783 251440 11799 251582
rect 11733 251424 11799 251440
rect 12153 251582 12219 251598
rect 12153 251440 12169 251582
rect 12203 251440 12219 251582
rect 12153 251424 12219 251440
rect 12573 251582 12639 251598
rect 12573 251440 12589 251582
rect 12623 251440 12639 251582
rect 12573 251424 12639 251440
rect 12993 251582 13059 251598
rect 12993 251440 13009 251582
rect 13043 251440 13059 251582
rect 12993 251424 13059 251440
rect 13413 251582 13479 251598
rect 13413 251440 13429 251582
rect 13463 251440 13479 251582
rect 13413 251424 13479 251440
rect 13833 251582 13899 251598
rect 13833 251440 13849 251582
rect 13883 251440 13899 251582
rect 13833 251424 13899 251440
rect 14253 251582 14319 251598
rect 14253 251440 14269 251582
rect 14303 251440 14319 251582
rect 14253 251424 14319 251440
rect 14673 251582 14739 251598
rect 14673 251440 14689 251582
rect 14723 251440 14739 251582
rect 14673 251424 14739 251440
rect 15093 251582 15159 251598
rect 15093 251440 15109 251582
rect 15143 251440 15159 251582
rect 15093 251424 15159 251440
rect 15513 251582 15579 251598
rect 15513 251440 15529 251582
rect 15563 251440 15579 251582
rect 15513 251424 15579 251440
rect 15933 251582 15999 251598
rect 15933 251440 15949 251582
rect 15983 251440 15999 251582
rect 15933 251424 15999 251440
rect 16353 251582 16419 251598
rect 16353 251440 16369 251582
rect 16403 251440 16419 251582
rect 16353 251424 16419 251440
rect 16773 251582 16839 251598
rect 16773 251440 16789 251582
rect 16823 251440 16839 251582
rect 16773 251424 16839 251440
rect 17193 251582 17259 251598
rect 17193 251440 17209 251582
rect 17243 251440 17259 251582
rect 17193 251424 17259 251440
rect 17613 251582 17679 251598
rect 17613 251440 17629 251582
rect 17663 251440 17679 251582
rect 17613 251424 17679 251440
rect 18033 251582 18099 251598
rect 18033 251440 18049 251582
rect 18083 251440 18099 251582
rect 18033 251424 18099 251440
rect 18453 251582 18519 251598
rect 18453 251440 18469 251582
rect 18503 251440 18519 251582
rect 18453 251424 18519 251440
rect 18873 251582 18939 251598
rect 18873 251440 18889 251582
rect 18923 251440 18939 251582
rect 18873 251424 18939 251440
rect 19293 251582 19359 251598
rect 19293 251440 19309 251582
rect 19343 251440 19359 251582
rect 19293 251424 19359 251440
rect 19713 251582 19779 251598
rect 19713 251440 19729 251582
rect 19763 251440 19779 251582
rect 19713 251424 19779 251440
rect 20133 251582 20199 251598
rect 20133 251440 20149 251582
rect 20183 251440 20199 251582
rect 20133 251424 20199 251440
rect 20553 251582 20619 251598
rect 20553 251440 20569 251582
rect 20603 251440 20619 251582
rect 20553 251424 20619 251440
rect 20973 251582 21039 251598
rect 20973 251440 20989 251582
rect 21023 251440 21039 251582
rect 20973 251424 21039 251440
rect 21393 251582 21459 251598
rect 21393 251440 21409 251582
rect 21443 251440 21459 251582
rect 21393 251424 21459 251440
rect 21813 251582 21879 251598
rect 21813 251440 21829 251582
rect 21863 251440 21879 251582
rect 21813 251424 21879 251440
rect 22233 251582 22299 251598
rect 22233 251440 22249 251582
rect 22283 251440 22299 251582
rect 22233 251424 22299 251440
rect 22653 251582 22719 251598
rect 22653 251440 22669 251582
rect 22703 251440 22719 251582
rect 22653 251424 22719 251440
rect 23073 251582 23139 251598
rect 23073 251440 23089 251582
rect 23123 251440 23139 251582
rect 23073 251424 23139 251440
rect 23493 251582 23559 251598
rect 23493 251440 23509 251582
rect 23543 251440 23559 251582
rect 23493 251424 23559 251440
rect 23913 251582 23979 251598
rect 23913 251440 23929 251582
rect 23963 251440 23979 251582
rect 23913 251424 23979 251440
rect 24333 251582 24399 251598
rect 24333 251440 24349 251582
rect 24383 251440 24399 251582
rect 24333 251424 24399 251440
rect 24753 251582 24819 251598
rect 24753 251440 24769 251582
rect 24803 251440 24819 251582
rect 24753 251424 24819 251440
rect 25173 251582 25239 251598
rect 25173 251440 25189 251582
rect 25223 251440 25239 251582
rect 25173 251424 25239 251440
rect 25593 251582 25659 251598
rect 25593 251440 25609 251582
rect 25643 251440 25659 251582
rect 25593 251424 25659 251440
rect 26013 251582 26079 251598
rect 26013 251440 26029 251582
rect 26063 251440 26079 251582
rect 26013 251424 26079 251440
rect 26433 251582 26499 251598
rect 26433 251440 26449 251582
rect 26483 251440 26499 251582
rect 26433 251424 26499 251440
rect 26853 251582 26919 251598
rect 26853 251440 26869 251582
rect 26903 251440 26919 251582
rect 26853 251424 26919 251440
rect 27273 251582 27339 251598
rect 27273 251440 27289 251582
rect 27323 251440 27339 251582
rect 27273 251424 27339 251440
rect -3999 251393 -3969 251419
rect -3789 251393 -3759 251424
rect -3579 251393 -3549 251419
rect -3369 251393 -3339 251424
rect -3159 251393 -3129 251419
rect -2949 251393 -2919 251424
rect -2739 251393 -2709 251419
rect -2529 251393 -2499 251424
rect -2319 251393 -2289 251419
rect -2109 251393 -2079 251424
rect -1899 251393 -1869 251419
rect -1689 251393 -1659 251424
rect -1479 251393 -1449 251419
rect -1269 251393 -1239 251424
rect -1059 251393 -1029 251419
rect -849 251393 -819 251424
rect -639 251393 -609 251419
rect -429 251393 -399 251424
rect -219 251393 -189 251419
rect -9 251393 21 251424
rect 201 251393 231 251419
rect 411 251393 441 251424
rect 621 251393 651 251419
rect 831 251393 861 251424
rect 1041 251393 1071 251419
rect 1251 251393 1281 251424
rect 1461 251393 1491 251419
rect 1671 251393 1701 251424
rect 1881 251393 1911 251419
rect 2091 251393 2121 251424
rect 2301 251393 2331 251419
rect 2511 251393 2541 251424
rect 2721 251393 2751 251419
rect 2931 251393 2961 251424
rect 3141 251393 3171 251419
rect 3351 251393 3381 251424
rect 3561 251393 3591 251419
rect 3771 251393 3801 251424
rect 3981 251393 4011 251419
rect 4191 251393 4221 251424
rect 4401 251393 4431 251419
rect 4611 251393 4641 251424
rect 4821 251393 4851 251419
rect 5031 251393 5061 251424
rect 5241 251393 5271 251419
rect 5451 251393 5481 251424
rect 5661 251393 5691 251419
rect 5871 251393 5901 251424
rect 6081 251393 6111 251419
rect 6291 251393 6321 251424
rect 6501 251393 6531 251419
rect 6711 251393 6741 251424
rect 6921 251393 6951 251419
rect 7131 251393 7161 251424
rect 7341 251393 7371 251419
rect 7551 251393 7581 251424
rect 7761 251393 7791 251419
rect 7971 251393 8001 251424
rect 8181 251393 8211 251419
rect 8391 251393 8421 251424
rect 8601 251393 8631 251419
rect 8811 251393 8841 251424
rect 9021 251393 9051 251419
rect 9231 251393 9261 251424
rect 9441 251393 9471 251419
rect 9651 251393 9681 251424
rect 9861 251393 9891 251419
rect 10071 251393 10101 251424
rect 10281 251393 10311 251419
rect 10491 251393 10521 251424
rect 10701 251393 10731 251419
rect 10911 251393 10941 251424
rect 11121 251393 11151 251419
rect 11331 251393 11361 251424
rect 11541 251393 11571 251419
rect 11751 251393 11781 251424
rect 11961 251393 11991 251419
rect 12171 251393 12201 251424
rect 12381 251393 12411 251419
rect 12591 251393 12621 251424
rect 12801 251393 12831 251419
rect 13011 251393 13041 251424
rect 13221 251393 13251 251419
rect 13431 251393 13461 251424
rect 13641 251393 13671 251419
rect 13851 251393 13881 251424
rect 14061 251393 14091 251419
rect 14271 251393 14301 251424
rect 14481 251393 14511 251419
rect 14691 251393 14721 251424
rect 14901 251393 14931 251419
rect 15111 251393 15141 251424
rect 15321 251393 15351 251419
rect 15531 251393 15561 251424
rect 15741 251393 15771 251419
rect 15951 251393 15981 251424
rect 16161 251393 16191 251419
rect 16371 251393 16401 251424
rect 16581 251393 16611 251419
rect 16791 251393 16821 251424
rect 17001 251393 17031 251419
rect 17211 251393 17241 251424
rect 17421 251393 17451 251419
rect 17631 251393 17661 251424
rect 17841 251393 17871 251419
rect 18051 251393 18081 251424
rect 18261 251393 18291 251419
rect 18471 251393 18501 251424
rect 18681 251393 18711 251419
rect 18891 251393 18921 251424
rect 19101 251393 19131 251419
rect 19311 251393 19341 251424
rect 19521 251393 19551 251419
rect 19731 251393 19761 251424
rect 19941 251393 19971 251419
rect 20151 251393 20181 251424
rect 20361 251393 20391 251419
rect 20571 251393 20601 251424
rect 20781 251393 20811 251419
rect 20991 251393 21021 251424
rect 21201 251393 21231 251419
rect 21411 251393 21441 251424
rect 21621 251393 21651 251419
rect 21831 251393 21861 251424
rect 22041 251393 22071 251419
rect 22251 251393 22281 251424
rect 22461 251393 22491 251419
rect 22671 251393 22701 251424
rect 22881 251393 22911 251419
rect 23091 251393 23121 251424
rect 23301 251393 23331 251419
rect 23511 251393 23541 251424
rect 23721 251393 23751 251419
rect 23931 251393 23961 251424
rect 24141 251393 24171 251419
rect 24351 251393 24381 251424
rect 24561 251393 24591 251419
rect 24771 251393 24801 251424
rect 24981 251393 25011 251419
rect 25191 251393 25221 251424
rect 25401 251393 25431 251419
rect 25611 251393 25641 251424
rect 25821 251393 25851 251419
rect 26031 251393 26061 251424
rect 26241 251393 26271 251419
rect 26451 251393 26481 251424
rect 26661 251393 26691 251419
rect 26871 251393 26901 251424
rect 27081 251393 27111 251419
rect 27291 251393 27321 251424
rect -3999 250562 -3969 250593
rect -3789 250567 -3759 250593
rect -3579 250562 -3549 250593
rect -3369 250567 -3339 250593
rect -3159 250562 -3129 250593
rect -2949 250567 -2919 250593
rect -2739 250562 -2709 250593
rect -2529 250567 -2499 250593
rect -2319 250562 -2289 250593
rect -2109 250567 -2079 250593
rect -1899 250562 -1869 250593
rect -1689 250567 -1659 250593
rect -1479 250562 -1449 250593
rect -1269 250567 -1239 250593
rect -1059 250562 -1029 250593
rect -849 250567 -819 250593
rect -639 250562 -609 250593
rect -429 250567 -399 250593
rect -219 250562 -189 250593
rect -9 250567 21 250593
rect 201 250562 231 250593
rect 411 250567 441 250593
rect 621 250562 651 250593
rect 831 250567 861 250593
rect 1041 250562 1071 250593
rect 1251 250567 1281 250593
rect 1461 250562 1491 250593
rect 1671 250567 1701 250593
rect 1881 250562 1911 250593
rect 2091 250567 2121 250593
rect 2301 250562 2331 250593
rect 2511 250567 2541 250593
rect 2721 250562 2751 250593
rect 2931 250567 2961 250593
rect 3141 250562 3171 250593
rect 3351 250567 3381 250593
rect 3561 250562 3591 250593
rect 3771 250567 3801 250593
rect 3981 250562 4011 250593
rect 4191 250567 4221 250593
rect 4401 250562 4431 250593
rect 4611 250567 4641 250593
rect 4821 250562 4851 250593
rect 5031 250567 5061 250593
rect 5241 250562 5271 250593
rect 5451 250567 5481 250593
rect 5661 250562 5691 250593
rect 5871 250567 5901 250593
rect 6081 250562 6111 250593
rect 6291 250567 6321 250593
rect 6501 250562 6531 250593
rect 6711 250567 6741 250593
rect 6921 250562 6951 250593
rect 7131 250567 7161 250593
rect 7341 250562 7371 250593
rect 7551 250567 7581 250593
rect 7761 250562 7791 250593
rect 7971 250567 8001 250593
rect 8181 250562 8211 250593
rect 8391 250567 8421 250593
rect 8601 250562 8631 250593
rect 8811 250567 8841 250593
rect 9021 250562 9051 250593
rect 9231 250567 9261 250593
rect 9441 250562 9471 250593
rect 9651 250567 9681 250593
rect 9861 250562 9891 250593
rect 10071 250567 10101 250593
rect 10281 250562 10311 250593
rect 10491 250567 10521 250593
rect 10701 250562 10731 250593
rect 10911 250567 10941 250593
rect 11121 250562 11151 250593
rect 11331 250567 11361 250593
rect 11541 250562 11571 250593
rect 11751 250567 11781 250593
rect 11961 250562 11991 250593
rect 12171 250567 12201 250593
rect 12381 250562 12411 250593
rect 12591 250567 12621 250593
rect 12801 250562 12831 250593
rect 13011 250567 13041 250593
rect 13221 250562 13251 250593
rect 13431 250567 13461 250593
rect 13641 250562 13671 250593
rect 13851 250567 13881 250593
rect 14061 250562 14091 250593
rect 14271 250567 14301 250593
rect 14481 250562 14511 250593
rect 14691 250567 14721 250593
rect 14901 250562 14931 250593
rect 15111 250567 15141 250593
rect 15321 250562 15351 250593
rect 15531 250567 15561 250593
rect 15741 250562 15771 250593
rect 15951 250567 15981 250593
rect 16161 250562 16191 250593
rect 16371 250567 16401 250593
rect 16581 250562 16611 250593
rect 16791 250567 16821 250593
rect 17001 250562 17031 250593
rect 17211 250567 17241 250593
rect 17421 250562 17451 250593
rect 17631 250567 17661 250593
rect 17841 250562 17871 250593
rect 18051 250567 18081 250593
rect 18261 250562 18291 250593
rect 18471 250567 18501 250593
rect 18681 250562 18711 250593
rect 18891 250567 18921 250593
rect 19101 250562 19131 250593
rect 19311 250567 19341 250593
rect 19521 250562 19551 250593
rect 19731 250567 19761 250593
rect 19941 250562 19971 250593
rect 20151 250567 20181 250593
rect 20361 250562 20391 250593
rect 20571 250567 20601 250593
rect 20781 250562 20811 250593
rect 20991 250567 21021 250593
rect 21201 250562 21231 250593
rect 21411 250567 21441 250593
rect 21621 250562 21651 250593
rect 21831 250567 21861 250593
rect 22041 250562 22071 250593
rect 22251 250567 22281 250593
rect 22461 250562 22491 250593
rect 22671 250567 22701 250593
rect 22881 250562 22911 250593
rect 23091 250567 23121 250593
rect 23301 250562 23331 250593
rect 23511 250567 23541 250593
rect 23721 250562 23751 250593
rect 23931 250567 23961 250593
rect 24141 250562 24171 250593
rect 24351 250567 24381 250593
rect 24561 250562 24591 250593
rect 24771 250567 24801 250593
rect 24981 250562 25011 250593
rect 25191 250567 25221 250593
rect 25401 250562 25431 250593
rect 25611 250567 25641 250593
rect 25821 250562 25851 250593
rect 26031 250567 26061 250593
rect 26241 250562 26271 250593
rect 26451 250567 26481 250593
rect 26661 250562 26691 250593
rect 26871 250567 26901 250593
rect 27081 250562 27111 250593
rect 27291 250567 27321 250593
rect -4017 250546 -3951 250562
rect -4017 250404 -4001 250546
rect -3967 250404 -3951 250546
rect -4017 250388 -3951 250404
rect -3597 250546 -3531 250562
rect -3597 250404 -3581 250546
rect -3547 250404 -3531 250546
rect -3597 250388 -3531 250404
rect -3177 250546 -3111 250562
rect -3177 250404 -3161 250546
rect -3127 250404 -3111 250546
rect -3177 250388 -3111 250404
rect -2757 250546 -2691 250562
rect -2757 250404 -2741 250546
rect -2707 250404 -2691 250546
rect -2757 250388 -2691 250404
rect -2337 250546 -2271 250562
rect -2337 250404 -2321 250546
rect -2287 250404 -2271 250546
rect -2337 250388 -2271 250404
rect -1917 250546 -1851 250562
rect -1917 250404 -1901 250546
rect -1867 250404 -1851 250546
rect -1917 250388 -1851 250404
rect -1497 250546 -1431 250562
rect -1497 250404 -1481 250546
rect -1447 250404 -1431 250546
rect -1497 250388 -1431 250404
rect -1077 250546 -1011 250562
rect -1077 250404 -1061 250546
rect -1027 250404 -1011 250546
rect -1077 250388 -1011 250404
rect -657 250546 -591 250562
rect -657 250404 -641 250546
rect -607 250404 -591 250546
rect -657 250388 -591 250404
rect -237 250546 -171 250562
rect -237 250404 -221 250546
rect -187 250404 -171 250546
rect -237 250388 -171 250404
rect 183 250546 249 250562
rect 183 250404 199 250546
rect 233 250404 249 250546
rect 183 250388 249 250404
rect 603 250546 669 250562
rect 603 250404 619 250546
rect 653 250404 669 250546
rect 603 250388 669 250404
rect 1023 250546 1089 250562
rect 1023 250404 1039 250546
rect 1073 250404 1089 250546
rect 1023 250388 1089 250404
rect 1443 250546 1509 250562
rect 1443 250404 1459 250546
rect 1493 250404 1509 250546
rect 1443 250388 1509 250404
rect 1863 250546 1929 250562
rect 1863 250404 1879 250546
rect 1913 250404 1929 250546
rect 1863 250388 1929 250404
rect 2283 250546 2349 250562
rect 2283 250404 2299 250546
rect 2333 250404 2349 250546
rect 2283 250388 2349 250404
rect 2703 250546 2769 250562
rect 2703 250404 2719 250546
rect 2753 250404 2769 250546
rect 2703 250388 2769 250404
rect 3123 250546 3189 250562
rect 3123 250404 3139 250546
rect 3173 250404 3189 250546
rect 3123 250388 3189 250404
rect 3543 250546 3609 250562
rect 3543 250404 3559 250546
rect 3593 250404 3609 250546
rect 3543 250388 3609 250404
rect 3963 250546 4029 250562
rect 3963 250404 3979 250546
rect 4013 250404 4029 250546
rect 3963 250388 4029 250404
rect 4383 250546 4449 250562
rect 4383 250404 4399 250546
rect 4433 250404 4449 250546
rect 4383 250388 4449 250404
rect 4803 250546 4869 250562
rect 4803 250404 4819 250546
rect 4853 250404 4869 250546
rect 4803 250388 4869 250404
rect 5223 250546 5289 250562
rect 5223 250404 5239 250546
rect 5273 250404 5289 250546
rect 5223 250388 5289 250404
rect 5643 250546 5709 250562
rect 5643 250404 5659 250546
rect 5693 250404 5709 250546
rect 5643 250388 5709 250404
rect 6063 250546 6129 250562
rect 6063 250404 6079 250546
rect 6113 250404 6129 250546
rect 6063 250388 6129 250404
rect 6483 250546 6549 250562
rect 6483 250404 6499 250546
rect 6533 250404 6549 250546
rect 6483 250388 6549 250404
rect 6903 250546 6969 250562
rect 6903 250404 6919 250546
rect 6953 250404 6969 250546
rect 6903 250388 6969 250404
rect 7323 250546 7389 250562
rect 7323 250404 7339 250546
rect 7373 250404 7389 250546
rect 7323 250388 7389 250404
rect 7743 250546 7809 250562
rect 7743 250404 7759 250546
rect 7793 250404 7809 250546
rect 7743 250388 7809 250404
rect 8163 250546 8229 250562
rect 8163 250404 8179 250546
rect 8213 250404 8229 250546
rect 8163 250388 8229 250404
rect 8583 250546 8649 250562
rect 8583 250404 8599 250546
rect 8633 250404 8649 250546
rect 8583 250388 8649 250404
rect 9003 250546 9069 250562
rect 9003 250404 9019 250546
rect 9053 250404 9069 250546
rect 9003 250388 9069 250404
rect 9423 250546 9489 250562
rect 9423 250404 9439 250546
rect 9473 250404 9489 250546
rect 9423 250388 9489 250404
rect 9843 250546 9909 250562
rect 9843 250404 9859 250546
rect 9893 250404 9909 250546
rect 9843 250388 9909 250404
rect 10263 250546 10329 250562
rect 10263 250404 10279 250546
rect 10313 250404 10329 250546
rect 10263 250388 10329 250404
rect 10683 250546 10749 250562
rect 10683 250404 10699 250546
rect 10733 250404 10749 250546
rect 10683 250388 10749 250404
rect 11103 250546 11169 250562
rect 11103 250404 11119 250546
rect 11153 250404 11169 250546
rect 11103 250388 11169 250404
rect 11523 250546 11589 250562
rect 11523 250404 11539 250546
rect 11573 250404 11589 250546
rect 11523 250388 11589 250404
rect 11943 250546 12009 250562
rect 11943 250404 11959 250546
rect 11993 250404 12009 250546
rect 11943 250388 12009 250404
rect 12363 250546 12429 250562
rect 12363 250404 12379 250546
rect 12413 250404 12429 250546
rect 12363 250388 12429 250404
rect 12783 250546 12849 250562
rect 12783 250404 12799 250546
rect 12833 250404 12849 250546
rect 12783 250388 12849 250404
rect 13203 250546 13269 250562
rect 13203 250404 13219 250546
rect 13253 250404 13269 250546
rect 13203 250388 13269 250404
rect 13623 250546 13689 250562
rect 13623 250404 13639 250546
rect 13673 250404 13689 250546
rect 13623 250388 13689 250404
rect 14043 250546 14109 250562
rect 14043 250404 14059 250546
rect 14093 250404 14109 250546
rect 14043 250388 14109 250404
rect 14463 250546 14529 250562
rect 14463 250404 14479 250546
rect 14513 250404 14529 250546
rect 14463 250388 14529 250404
rect 14883 250546 14949 250562
rect 14883 250404 14899 250546
rect 14933 250404 14949 250546
rect 14883 250388 14949 250404
rect 15303 250546 15369 250562
rect 15303 250404 15319 250546
rect 15353 250404 15369 250546
rect 15303 250388 15369 250404
rect 15723 250546 15789 250562
rect 15723 250404 15739 250546
rect 15773 250404 15789 250546
rect 15723 250388 15789 250404
rect 16143 250546 16209 250562
rect 16143 250404 16159 250546
rect 16193 250404 16209 250546
rect 16143 250388 16209 250404
rect 16563 250546 16629 250562
rect 16563 250404 16579 250546
rect 16613 250404 16629 250546
rect 16563 250388 16629 250404
rect 16983 250546 17049 250562
rect 16983 250404 16999 250546
rect 17033 250404 17049 250546
rect 16983 250388 17049 250404
rect 17403 250546 17469 250562
rect 17403 250404 17419 250546
rect 17453 250404 17469 250546
rect 17403 250388 17469 250404
rect 17823 250546 17889 250562
rect 17823 250404 17839 250546
rect 17873 250404 17889 250546
rect 17823 250388 17889 250404
rect 18243 250546 18309 250562
rect 18243 250404 18259 250546
rect 18293 250404 18309 250546
rect 18243 250388 18309 250404
rect 18663 250546 18729 250562
rect 18663 250404 18679 250546
rect 18713 250404 18729 250546
rect 18663 250388 18729 250404
rect 19083 250546 19149 250562
rect 19083 250404 19099 250546
rect 19133 250404 19149 250546
rect 19083 250388 19149 250404
rect 19503 250546 19569 250562
rect 19503 250404 19519 250546
rect 19553 250404 19569 250546
rect 19503 250388 19569 250404
rect 19923 250546 19989 250562
rect 19923 250404 19939 250546
rect 19973 250404 19989 250546
rect 19923 250388 19989 250404
rect 20343 250546 20409 250562
rect 20343 250404 20359 250546
rect 20393 250404 20409 250546
rect 20343 250388 20409 250404
rect 20763 250546 20829 250562
rect 20763 250404 20779 250546
rect 20813 250404 20829 250546
rect 20763 250388 20829 250404
rect 21183 250546 21249 250562
rect 21183 250404 21199 250546
rect 21233 250404 21249 250546
rect 21183 250388 21249 250404
rect 21603 250546 21669 250562
rect 21603 250404 21619 250546
rect 21653 250404 21669 250546
rect 21603 250388 21669 250404
rect 22023 250546 22089 250562
rect 22023 250404 22039 250546
rect 22073 250404 22089 250546
rect 22023 250388 22089 250404
rect 22443 250546 22509 250562
rect 22443 250404 22459 250546
rect 22493 250404 22509 250546
rect 22443 250388 22509 250404
rect 22863 250546 22929 250562
rect 22863 250404 22879 250546
rect 22913 250404 22929 250546
rect 22863 250388 22929 250404
rect 23283 250546 23349 250562
rect 23283 250404 23299 250546
rect 23333 250404 23349 250546
rect 23283 250388 23349 250404
rect 23703 250546 23769 250562
rect 23703 250404 23719 250546
rect 23753 250404 23769 250546
rect 23703 250388 23769 250404
rect 24123 250546 24189 250562
rect 24123 250404 24139 250546
rect 24173 250404 24189 250546
rect 24123 250388 24189 250404
rect 24543 250546 24609 250562
rect 24543 250404 24559 250546
rect 24593 250404 24609 250546
rect 24543 250388 24609 250404
rect 24963 250546 25029 250562
rect 24963 250404 24979 250546
rect 25013 250404 25029 250546
rect 24963 250388 25029 250404
rect 25383 250546 25449 250562
rect 25383 250404 25399 250546
rect 25433 250404 25449 250546
rect 25383 250388 25449 250404
rect 25803 250546 25869 250562
rect 25803 250404 25819 250546
rect 25853 250404 25869 250546
rect 25803 250388 25869 250404
rect 26223 250546 26289 250562
rect 26223 250404 26239 250546
rect 26273 250404 26289 250546
rect 26223 250388 26289 250404
rect 26643 250546 26709 250562
rect 26643 250404 26659 250546
rect 26693 250404 26709 250546
rect 26643 250388 26709 250404
rect 27063 250546 27129 250562
rect 27063 250404 27079 250546
rect 27113 250404 27129 250546
rect 27063 250388 27129 250404
rect -3999 250357 -3969 250388
rect -3789 250357 -3759 250383
rect -3579 250357 -3549 250388
rect -3369 250357 -3339 250383
rect -3159 250357 -3129 250388
rect -2949 250357 -2919 250383
rect -2739 250357 -2709 250388
rect -2529 250357 -2499 250383
rect -2319 250357 -2289 250388
rect -2109 250357 -2079 250383
rect -1899 250357 -1869 250388
rect -1689 250357 -1659 250383
rect -1479 250357 -1449 250388
rect -1269 250357 -1239 250383
rect -1059 250357 -1029 250388
rect -849 250357 -819 250383
rect -639 250357 -609 250388
rect -429 250357 -399 250383
rect -219 250357 -189 250388
rect -9 250357 21 250383
rect 201 250357 231 250388
rect 411 250357 441 250383
rect 621 250357 651 250388
rect 831 250357 861 250383
rect 1041 250357 1071 250388
rect 1251 250357 1281 250383
rect 1461 250357 1491 250388
rect 1671 250357 1701 250383
rect 1881 250357 1911 250388
rect 2091 250357 2121 250383
rect 2301 250357 2331 250388
rect 2511 250357 2541 250383
rect 2721 250357 2751 250388
rect 2931 250357 2961 250383
rect 3141 250357 3171 250388
rect 3351 250357 3381 250383
rect 3561 250357 3591 250388
rect 3771 250357 3801 250383
rect 3981 250357 4011 250388
rect 4191 250357 4221 250383
rect 4401 250357 4431 250388
rect 4611 250357 4641 250383
rect 4821 250357 4851 250388
rect 5031 250357 5061 250383
rect 5241 250357 5271 250388
rect 5451 250357 5481 250383
rect 5661 250357 5691 250388
rect 5871 250357 5901 250383
rect 6081 250357 6111 250388
rect 6291 250357 6321 250383
rect 6501 250357 6531 250388
rect 6711 250357 6741 250383
rect 6921 250357 6951 250388
rect 7131 250357 7161 250383
rect 7341 250357 7371 250388
rect 7551 250357 7581 250383
rect 7761 250357 7791 250388
rect 7971 250357 8001 250383
rect 8181 250357 8211 250388
rect 8391 250357 8421 250383
rect 8601 250357 8631 250388
rect 8811 250357 8841 250383
rect 9021 250357 9051 250388
rect 9231 250357 9261 250383
rect 9441 250357 9471 250388
rect 9651 250357 9681 250383
rect 9861 250357 9891 250388
rect 10071 250357 10101 250383
rect 10281 250357 10311 250388
rect 10491 250357 10521 250383
rect 10701 250357 10731 250388
rect 10911 250357 10941 250383
rect 11121 250357 11151 250388
rect 11331 250357 11361 250383
rect 11541 250357 11571 250388
rect 11751 250357 11781 250383
rect 11961 250357 11991 250388
rect 12171 250357 12201 250383
rect 12381 250357 12411 250388
rect 12591 250357 12621 250383
rect 12801 250357 12831 250388
rect 13011 250357 13041 250383
rect 13221 250357 13251 250388
rect 13431 250357 13461 250383
rect 13641 250357 13671 250388
rect 13851 250357 13881 250383
rect 14061 250357 14091 250388
rect 14271 250357 14301 250383
rect 14481 250357 14511 250388
rect 14691 250357 14721 250383
rect 14901 250357 14931 250388
rect 15111 250357 15141 250383
rect 15321 250357 15351 250388
rect 15531 250357 15561 250383
rect 15741 250357 15771 250388
rect 15951 250357 15981 250383
rect 16161 250357 16191 250388
rect 16371 250357 16401 250383
rect 16581 250357 16611 250388
rect 16791 250357 16821 250383
rect 17001 250357 17031 250388
rect 17211 250357 17241 250383
rect 17421 250357 17451 250388
rect 17631 250357 17661 250383
rect 17841 250357 17871 250388
rect 18051 250357 18081 250383
rect 18261 250357 18291 250388
rect 18471 250357 18501 250383
rect 18681 250357 18711 250388
rect 18891 250357 18921 250383
rect 19101 250357 19131 250388
rect 19311 250357 19341 250383
rect 19521 250357 19551 250388
rect 19731 250357 19761 250383
rect 19941 250357 19971 250388
rect 20151 250357 20181 250383
rect 20361 250357 20391 250388
rect 20571 250357 20601 250383
rect 20781 250357 20811 250388
rect 20991 250357 21021 250383
rect 21201 250357 21231 250388
rect 21411 250357 21441 250383
rect 21621 250357 21651 250388
rect 21831 250357 21861 250383
rect 22041 250357 22071 250388
rect 22251 250357 22281 250383
rect 22461 250357 22491 250388
rect 22671 250357 22701 250383
rect 22881 250357 22911 250388
rect 23091 250357 23121 250383
rect 23301 250357 23331 250388
rect 23511 250357 23541 250383
rect 23721 250357 23751 250388
rect 23931 250357 23961 250383
rect 24141 250357 24171 250388
rect 24351 250357 24381 250383
rect 24561 250357 24591 250388
rect 24771 250357 24801 250383
rect 24981 250357 25011 250388
rect 25191 250357 25221 250383
rect 25401 250357 25431 250388
rect 25611 250357 25641 250383
rect 25821 250357 25851 250388
rect 26031 250357 26061 250383
rect 26241 250357 26271 250388
rect 26451 250357 26481 250383
rect 26661 250357 26691 250388
rect 26871 250357 26901 250383
rect 27081 250357 27111 250388
rect 27291 250357 27321 250383
rect -3999 249531 -3969 249557
rect -3789 249526 -3759 249557
rect -3579 249531 -3549 249557
rect -3369 249526 -3339 249557
rect -3159 249531 -3129 249557
rect -2949 249526 -2919 249557
rect -2739 249531 -2709 249557
rect -2529 249526 -2499 249557
rect -2319 249531 -2289 249557
rect -2109 249526 -2079 249557
rect -1899 249531 -1869 249557
rect -1689 249526 -1659 249557
rect -1479 249531 -1449 249557
rect -1269 249526 -1239 249557
rect -1059 249531 -1029 249557
rect -849 249526 -819 249557
rect -639 249531 -609 249557
rect -429 249526 -399 249557
rect -219 249531 -189 249557
rect -9 249526 21 249557
rect 201 249531 231 249557
rect 411 249526 441 249557
rect 621 249531 651 249557
rect 831 249526 861 249557
rect 1041 249531 1071 249557
rect 1251 249526 1281 249557
rect 1461 249531 1491 249557
rect 1671 249526 1701 249557
rect 1881 249531 1911 249557
rect 2091 249526 2121 249557
rect 2301 249531 2331 249557
rect 2511 249526 2541 249557
rect 2721 249531 2751 249557
rect 2931 249526 2961 249557
rect 3141 249531 3171 249557
rect 3351 249526 3381 249557
rect 3561 249531 3591 249557
rect 3771 249526 3801 249557
rect 3981 249531 4011 249557
rect 4191 249526 4221 249557
rect 4401 249531 4431 249557
rect 4611 249526 4641 249557
rect 4821 249531 4851 249557
rect 5031 249526 5061 249557
rect 5241 249531 5271 249557
rect 5451 249526 5481 249557
rect 5661 249531 5691 249557
rect 5871 249526 5901 249557
rect 6081 249531 6111 249557
rect 6291 249526 6321 249557
rect 6501 249531 6531 249557
rect 6711 249526 6741 249557
rect 6921 249531 6951 249557
rect 7131 249526 7161 249557
rect 7341 249531 7371 249557
rect 7551 249526 7581 249557
rect 7761 249531 7791 249557
rect 7971 249526 8001 249557
rect 8181 249531 8211 249557
rect 8391 249526 8421 249557
rect 8601 249531 8631 249557
rect 8811 249526 8841 249557
rect 9021 249531 9051 249557
rect 9231 249526 9261 249557
rect 9441 249531 9471 249557
rect 9651 249526 9681 249557
rect 9861 249531 9891 249557
rect 10071 249526 10101 249557
rect 10281 249531 10311 249557
rect 10491 249526 10521 249557
rect 10701 249531 10731 249557
rect 10911 249526 10941 249557
rect 11121 249531 11151 249557
rect 11331 249526 11361 249557
rect 11541 249531 11571 249557
rect 11751 249526 11781 249557
rect 11961 249531 11991 249557
rect 12171 249526 12201 249557
rect 12381 249531 12411 249557
rect 12591 249526 12621 249557
rect 12801 249531 12831 249557
rect 13011 249526 13041 249557
rect 13221 249531 13251 249557
rect 13431 249526 13461 249557
rect 13641 249531 13671 249557
rect 13851 249526 13881 249557
rect 14061 249531 14091 249557
rect 14271 249526 14301 249557
rect 14481 249531 14511 249557
rect 14691 249526 14721 249557
rect 14901 249531 14931 249557
rect 15111 249526 15141 249557
rect 15321 249531 15351 249557
rect 15531 249526 15561 249557
rect 15741 249531 15771 249557
rect 15951 249526 15981 249557
rect 16161 249531 16191 249557
rect 16371 249526 16401 249557
rect 16581 249531 16611 249557
rect 16791 249526 16821 249557
rect 17001 249531 17031 249557
rect 17211 249526 17241 249557
rect 17421 249531 17451 249557
rect 17631 249526 17661 249557
rect 17841 249531 17871 249557
rect 18051 249526 18081 249557
rect 18261 249531 18291 249557
rect 18471 249526 18501 249557
rect 18681 249531 18711 249557
rect 18891 249526 18921 249557
rect 19101 249531 19131 249557
rect 19311 249526 19341 249557
rect 19521 249531 19551 249557
rect 19731 249526 19761 249557
rect 19941 249531 19971 249557
rect 20151 249526 20181 249557
rect 20361 249531 20391 249557
rect 20571 249526 20601 249557
rect 20781 249531 20811 249557
rect 20991 249526 21021 249557
rect 21201 249531 21231 249557
rect 21411 249526 21441 249557
rect 21621 249531 21651 249557
rect 21831 249526 21861 249557
rect 22041 249531 22071 249557
rect 22251 249526 22281 249557
rect 22461 249531 22491 249557
rect 22671 249526 22701 249557
rect 22881 249531 22911 249557
rect 23091 249526 23121 249557
rect 23301 249531 23331 249557
rect 23511 249526 23541 249557
rect 23721 249531 23751 249557
rect 23931 249526 23961 249557
rect 24141 249531 24171 249557
rect 24351 249526 24381 249557
rect 24561 249531 24591 249557
rect 24771 249526 24801 249557
rect 24981 249531 25011 249557
rect 25191 249526 25221 249557
rect 25401 249531 25431 249557
rect 25611 249526 25641 249557
rect 25821 249531 25851 249557
rect 26031 249526 26061 249557
rect 26241 249531 26271 249557
rect 26451 249526 26481 249557
rect 26661 249531 26691 249557
rect 26871 249526 26901 249557
rect 27081 249531 27111 249557
rect 27291 249526 27321 249557
rect -3807 249510 -3678 249526
rect -3807 249476 -3791 249510
rect -3695 249476 -3678 249510
rect -3807 249460 -3678 249476
rect -3387 249510 -3258 249526
rect -3387 249476 -3371 249510
rect -3275 249476 -3258 249510
rect -3387 249460 -3258 249476
rect -2967 249510 -2838 249526
rect -2967 249476 -2951 249510
rect -2855 249476 -2838 249510
rect -2967 249460 -2838 249476
rect -2547 249510 -2418 249526
rect -2547 249476 -2531 249510
rect -2435 249476 -2418 249510
rect -2547 249460 -2418 249476
rect -2127 249510 -1998 249526
rect -2127 249476 -2111 249510
rect -2015 249476 -1998 249510
rect -2127 249460 -1998 249476
rect -1707 249510 -1578 249526
rect -1707 249476 -1691 249510
rect -1595 249476 -1578 249510
rect -1707 249460 -1578 249476
rect -1287 249510 -1158 249526
rect -1287 249476 -1271 249510
rect -1175 249476 -1158 249510
rect -1287 249460 -1158 249476
rect -867 249510 -738 249526
rect -867 249476 -851 249510
rect -755 249476 -738 249510
rect -867 249460 -738 249476
rect -447 249510 -318 249526
rect -447 249476 -431 249510
rect -335 249476 -318 249510
rect -447 249460 -318 249476
rect -27 249510 102 249526
rect -27 249476 -11 249510
rect 85 249476 102 249510
rect -27 249460 102 249476
rect 393 249510 522 249526
rect 393 249476 409 249510
rect 505 249476 522 249510
rect 393 249460 522 249476
rect 813 249510 942 249526
rect 813 249476 829 249510
rect 925 249476 942 249510
rect 813 249460 942 249476
rect 1233 249510 1362 249526
rect 1233 249476 1249 249510
rect 1345 249476 1362 249510
rect 1233 249460 1362 249476
rect 1653 249510 1782 249526
rect 1653 249476 1669 249510
rect 1765 249476 1782 249510
rect 1653 249460 1782 249476
rect 2073 249510 2202 249526
rect 2073 249476 2089 249510
rect 2185 249476 2202 249510
rect 2073 249460 2202 249476
rect 2493 249510 2622 249526
rect 2493 249476 2509 249510
rect 2605 249476 2622 249510
rect 2493 249460 2622 249476
rect 2913 249510 3042 249526
rect 2913 249476 2929 249510
rect 3025 249476 3042 249510
rect 2913 249460 3042 249476
rect 3333 249510 3462 249526
rect 3333 249476 3349 249510
rect 3445 249476 3462 249510
rect 3333 249460 3462 249476
rect 3753 249510 3882 249526
rect 3753 249476 3769 249510
rect 3865 249476 3882 249510
rect 3753 249460 3882 249476
rect 4173 249510 4302 249526
rect 4173 249476 4189 249510
rect 4285 249476 4302 249510
rect 4173 249460 4302 249476
rect 4593 249510 4722 249526
rect 4593 249476 4609 249510
rect 4705 249476 4722 249510
rect 4593 249460 4722 249476
rect 5013 249510 5142 249526
rect 5013 249476 5029 249510
rect 5125 249476 5142 249510
rect 5013 249460 5142 249476
rect 5433 249510 5562 249526
rect 5433 249476 5449 249510
rect 5545 249476 5562 249510
rect 5433 249460 5562 249476
rect 5853 249510 5982 249526
rect 5853 249476 5869 249510
rect 5965 249476 5982 249510
rect 5853 249460 5982 249476
rect 6273 249510 6402 249526
rect 6273 249476 6289 249510
rect 6385 249476 6402 249510
rect 6273 249460 6402 249476
rect 6693 249510 6822 249526
rect 6693 249476 6709 249510
rect 6805 249476 6822 249510
rect 6693 249460 6822 249476
rect 7113 249510 7242 249526
rect 7113 249476 7129 249510
rect 7225 249476 7242 249510
rect 7113 249460 7242 249476
rect 7533 249510 7662 249526
rect 7533 249476 7549 249510
rect 7645 249476 7662 249510
rect 7533 249460 7662 249476
rect 7953 249510 8082 249526
rect 7953 249476 7969 249510
rect 8065 249476 8082 249510
rect 7953 249460 8082 249476
rect 8373 249510 8502 249526
rect 8373 249476 8389 249510
rect 8485 249476 8502 249510
rect 8373 249460 8502 249476
rect 8793 249510 8922 249526
rect 8793 249476 8809 249510
rect 8905 249476 8922 249510
rect 8793 249460 8922 249476
rect 9213 249510 9342 249526
rect 9213 249476 9229 249510
rect 9325 249476 9342 249510
rect 9213 249460 9342 249476
rect 9633 249510 9762 249526
rect 9633 249476 9649 249510
rect 9745 249476 9762 249510
rect 9633 249460 9762 249476
rect 10053 249510 10182 249526
rect 10053 249476 10069 249510
rect 10165 249476 10182 249510
rect 10053 249460 10182 249476
rect 10473 249510 10602 249526
rect 10473 249476 10489 249510
rect 10585 249476 10602 249510
rect 10473 249460 10602 249476
rect 10893 249510 11022 249526
rect 10893 249476 10909 249510
rect 11005 249476 11022 249510
rect 10893 249460 11022 249476
rect 11313 249510 11442 249526
rect 11313 249476 11329 249510
rect 11425 249476 11442 249510
rect 11313 249460 11442 249476
rect 11733 249510 11862 249526
rect 11733 249476 11749 249510
rect 11845 249476 11862 249510
rect 11733 249460 11862 249476
rect 12153 249510 12282 249526
rect 12153 249476 12169 249510
rect 12265 249476 12282 249510
rect 12153 249460 12282 249476
rect 12573 249510 12702 249526
rect 12573 249476 12589 249510
rect 12685 249476 12702 249510
rect 12573 249460 12702 249476
rect 12993 249510 13122 249526
rect 12993 249476 13009 249510
rect 13105 249476 13122 249510
rect 12993 249460 13122 249476
rect 13413 249510 13542 249526
rect 13413 249476 13429 249510
rect 13525 249476 13542 249510
rect 13413 249460 13542 249476
rect 13833 249510 13962 249526
rect 13833 249476 13849 249510
rect 13945 249476 13962 249510
rect 13833 249460 13962 249476
rect 14253 249510 14382 249526
rect 14253 249476 14269 249510
rect 14365 249476 14382 249510
rect 14253 249460 14382 249476
rect 14673 249510 14802 249526
rect 14673 249476 14689 249510
rect 14785 249476 14802 249510
rect 14673 249460 14802 249476
rect 15093 249510 15222 249526
rect 15093 249476 15109 249510
rect 15205 249476 15222 249510
rect 15093 249460 15222 249476
rect 15513 249510 15642 249526
rect 15513 249476 15529 249510
rect 15625 249476 15642 249510
rect 15513 249460 15642 249476
rect 15933 249510 16062 249526
rect 15933 249476 15949 249510
rect 16045 249476 16062 249510
rect 15933 249460 16062 249476
rect 16353 249510 16482 249526
rect 16353 249476 16369 249510
rect 16465 249476 16482 249510
rect 16353 249460 16482 249476
rect 16773 249510 16902 249526
rect 16773 249476 16789 249510
rect 16885 249476 16902 249510
rect 16773 249460 16902 249476
rect 17193 249510 17322 249526
rect 17193 249476 17209 249510
rect 17305 249476 17322 249510
rect 17193 249460 17322 249476
rect 17613 249510 17742 249526
rect 17613 249476 17629 249510
rect 17725 249476 17742 249510
rect 17613 249460 17742 249476
rect 18033 249510 18162 249526
rect 18033 249476 18049 249510
rect 18145 249476 18162 249510
rect 18033 249460 18162 249476
rect 18453 249510 18582 249526
rect 18453 249476 18469 249510
rect 18565 249476 18582 249510
rect 18453 249460 18582 249476
rect 18873 249510 19002 249526
rect 18873 249476 18889 249510
rect 18985 249476 19002 249510
rect 18873 249460 19002 249476
rect 19293 249510 19422 249526
rect 19293 249476 19309 249510
rect 19405 249476 19422 249510
rect 19293 249460 19422 249476
rect 19713 249510 19842 249526
rect 19713 249476 19729 249510
rect 19825 249476 19842 249510
rect 19713 249460 19842 249476
rect 20133 249510 20262 249526
rect 20133 249476 20149 249510
rect 20245 249476 20262 249510
rect 20133 249460 20262 249476
rect 20553 249510 20682 249526
rect 20553 249476 20569 249510
rect 20665 249476 20682 249510
rect 20553 249460 20682 249476
rect 20973 249510 21102 249526
rect 20973 249476 20989 249510
rect 21085 249476 21102 249510
rect 20973 249460 21102 249476
rect 21393 249510 21522 249526
rect 21393 249476 21409 249510
rect 21505 249476 21522 249510
rect 21393 249460 21522 249476
rect 21813 249510 21942 249526
rect 21813 249476 21829 249510
rect 21925 249476 21942 249510
rect 21813 249460 21942 249476
rect 22233 249510 22362 249526
rect 22233 249476 22249 249510
rect 22345 249476 22362 249510
rect 22233 249460 22362 249476
rect 22653 249510 22782 249526
rect 22653 249476 22669 249510
rect 22765 249476 22782 249510
rect 22653 249460 22782 249476
rect 23073 249510 23202 249526
rect 23073 249476 23089 249510
rect 23185 249476 23202 249510
rect 23073 249460 23202 249476
rect 23493 249510 23622 249526
rect 23493 249476 23509 249510
rect 23605 249476 23622 249510
rect 23493 249460 23622 249476
rect 23913 249510 24042 249526
rect 23913 249476 23929 249510
rect 24025 249476 24042 249510
rect 23913 249460 24042 249476
rect 24333 249510 24462 249526
rect 24333 249476 24349 249510
rect 24445 249476 24462 249510
rect 24333 249460 24462 249476
rect 24753 249510 24882 249526
rect 24753 249476 24769 249510
rect 24865 249476 24882 249510
rect 24753 249460 24882 249476
rect 25173 249510 25302 249526
rect 25173 249476 25189 249510
rect 25285 249476 25302 249510
rect 25173 249460 25302 249476
rect 25593 249510 25722 249526
rect 25593 249476 25609 249510
rect 25705 249476 25722 249510
rect 25593 249460 25722 249476
rect 26013 249510 26142 249526
rect 26013 249476 26029 249510
rect 26125 249476 26142 249510
rect 26013 249460 26142 249476
rect 26433 249510 26562 249526
rect 26433 249476 26449 249510
rect 26545 249476 26562 249510
rect 26433 249460 26562 249476
rect 26853 249510 26982 249526
rect 26853 249476 26869 249510
rect 26965 249476 26982 249510
rect 26853 249460 26982 249476
rect 27273 249510 27402 249526
rect 27273 249476 27289 249510
rect 27385 249476 27402 249510
rect 27273 249460 27402 249476
rect -4017 249273 -3888 249289
rect -4017 249239 -4001 249273
rect -3905 249239 -3888 249273
rect -4017 249223 -3888 249239
rect -3597 249273 -3468 249289
rect -3597 249239 -3581 249273
rect -3485 249239 -3468 249273
rect -3597 249223 -3468 249239
rect -3177 249273 -3048 249289
rect -3177 249239 -3161 249273
rect -3065 249239 -3048 249273
rect -3177 249223 -3048 249239
rect -2757 249273 -2628 249289
rect -2757 249239 -2741 249273
rect -2645 249239 -2628 249273
rect -2757 249223 -2628 249239
rect -2337 249273 -2208 249289
rect -2337 249239 -2321 249273
rect -2225 249239 -2208 249273
rect -2337 249223 -2208 249239
rect -1917 249273 -1788 249289
rect -1917 249239 -1901 249273
rect -1805 249239 -1788 249273
rect -1917 249223 -1788 249239
rect -1497 249273 -1368 249289
rect -1497 249239 -1481 249273
rect -1385 249239 -1368 249273
rect -1497 249223 -1368 249239
rect -1077 249273 -948 249289
rect -1077 249239 -1061 249273
rect -965 249239 -948 249273
rect -1077 249223 -948 249239
rect -657 249273 -528 249289
rect -657 249239 -641 249273
rect -545 249239 -528 249273
rect -657 249223 -528 249239
rect -237 249273 -108 249289
rect -237 249239 -221 249273
rect -125 249239 -108 249273
rect -237 249223 -108 249239
rect 183 249273 312 249289
rect 183 249239 199 249273
rect 295 249239 312 249273
rect 183 249223 312 249239
rect 603 249273 732 249289
rect 603 249239 619 249273
rect 715 249239 732 249273
rect 603 249223 732 249239
rect 1023 249273 1152 249289
rect 1023 249239 1039 249273
rect 1135 249239 1152 249273
rect 1023 249223 1152 249239
rect 1443 249273 1572 249289
rect 1443 249239 1459 249273
rect 1555 249239 1572 249273
rect 1443 249223 1572 249239
rect 1863 249273 1992 249289
rect 1863 249239 1879 249273
rect 1975 249239 1992 249273
rect 1863 249223 1992 249239
rect 2283 249273 2412 249289
rect 2283 249239 2299 249273
rect 2395 249239 2412 249273
rect 2283 249223 2412 249239
rect 2703 249273 2832 249289
rect 2703 249239 2719 249273
rect 2815 249239 2832 249273
rect 2703 249223 2832 249239
rect 3123 249273 3252 249289
rect 3123 249239 3139 249273
rect 3235 249239 3252 249273
rect 3123 249223 3252 249239
rect 3543 249273 3672 249289
rect 3543 249239 3559 249273
rect 3655 249239 3672 249273
rect 3543 249223 3672 249239
rect 3963 249273 4092 249289
rect 3963 249239 3979 249273
rect 4075 249239 4092 249273
rect 3963 249223 4092 249239
rect 4383 249273 4512 249289
rect 4383 249239 4399 249273
rect 4495 249239 4512 249273
rect 4383 249223 4512 249239
rect 4803 249273 4932 249289
rect 4803 249239 4819 249273
rect 4915 249239 4932 249273
rect 4803 249223 4932 249239
rect 5223 249273 5352 249289
rect 5223 249239 5239 249273
rect 5335 249239 5352 249273
rect 5223 249223 5352 249239
rect 5643 249273 5772 249289
rect 5643 249239 5659 249273
rect 5755 249239 5772 249273
rect 5643 249223 5772 249239
rect 6063 249273 6192 249289
rect 6063 249239 6079 249273
rect 6175 249239 6192 249273
rect 6063 249223 6192 249239
rect 6483 249273 6612 249289
rect 6483 249239 6499 249273
rect 6595 249239 6612 249273
rect 6483 249223 6612 249239
rect 6903 249273 7032 249289
rect 6903 249239 6919 249273
rect 7015 249239 7032 249273
rect 6903 249223 7032 249239
rect 7323 249273 7452 249289
rect 7323 249239 7339 249273
rect 7435 249239 7452 249273
rect 7323 249223 7452 249239
rect 7743 249273 7872 249289
rect 7743 249239 7759 249273
rect 7855 249239 7872 249273
rect 7743 249223 7872 249239
rect 8163 249273 8292 249289
rect 8163 249239 8179 249273
rect 8275 249239 8292 249273
rect 8163 249223 8292 249239
rect 8583 249273 8712 249289
rect 8583 249239 8599 249273
rect 8695 249239 8712 249273
rect 8583 249223 8712 249239
rect 9003 249273 9132 249289
rect 9003 249239 9019 249273
rect 9115 249239 9132 249273
rect 9003 249223 9132 249239
rect 9423 249273 9552 249289
rect 9423 249239 9439 249273
rect 9535 249239 9552 249273
rect 9423 249223 9552 249239
rect 9843 249273 9972 249289
rect 9843 249239 9859 249273
rect 9955 249239 9972 249273
rect 9843 249223 9972 249239
rect 10263 249273 10392 249289
rect 10263 249239 10279 249273
rect 10375 249239 10392 249273
rect 10263 249223 10392 249239
rect 10683 249273 10812 249289
rect 10683 249239 10699 249273
rect 10795 249239 10812 249273
rect 10683 249223 10812 249239
rect 11103 249273 11232 249289
rect 11103 249239 11119 249273
rect 11215 249239 11232 249273
rect 11103 249223 11232 249239
rect 11523 249273 11652 249289
rect 11523 249239 11539 249273
rect 11635 249239 11652 249273
rect 11523 249223 11652 249239
rect 11943 249273 12072 249289
rect 11943 249239 11959 249273
rect 12055 249239 12072 249273
rect 11943 249223 12072 249239
rect 12363 249273 12492 249289
rect 12363 249239 12379 249273
rect 12475 249239 12492 249273
rect 12363 249223 12492 249239
rect 12783 249273 12912 249289
rect 12783 249239 12799 249273
rect 12895 249239 12912 249273
rect 12783 249223 12912 249239
rect 13203 249273 13332 249289
rect 13203 249239 13219 249273
rect 13315 249239 13332 249273
rect 13203 249223 13332 249239
rect 13623 249273 13752 249289
rect 13623 249239 13639 249273
rect 13735 249239 13752 249273
rect 13623 249223 13752 249239
rect 14043 249273 14172 249289
rect 14043 249239 14059 249273
rect 14155 249239 14172 249273
rect 14043 249223 14172 249239
rect 14463 249273 14592 249289
rect 14463 249239 14479 249273
rect 14575 249239 14592 249273
rect 14463 249223 14592 249239
rect 14883 249273 15012 249289
rect 14883 249239 14899 249273
rect 14995 249239 15012 249273
rect 14883 249223 15012 249239
rect 15303 249273 15432 249289
rect 15303 249239 15319 249273
rect 15415 249239 15432 249273
rect 15303 249223 15432 249239
rect 15723 249273 15852 249289
rect 15723 249239 15739 249273
rect 15835 249239 15852 249273
rect 15723 249223 15852 249239
rect 16143 249273 16272 249289
rect 16143 249239 16159 249273
rect 16255 249239 16272 249273
rect 16143 249223 16272 249239
rect 16563 249273 16692 249289
rect 16563 249239 16579 249273
rect 16675 249239 16692 249273
rect 16563 249223 16692 249239
rect 16983 249273 17112 249289
rect 16983 249239 16999 249273
rect 17095 249239 17112 249273
rect 16983 249223 17112 249239
rect 17403 249273 17532 249289
rect 17403 249239 17419 249273
rect 17515 249239 17532 249273
rect 17403 249223 17532 249239
rect 17823 249273 17952 249289
rect 17823 249239 17839 249273
rect 17935 249239 17952 249273
rect 17823 249223 17952 249239
rect 18243 249273 18372 249289
rect 18243 249239 18259 249273
rect 18355 249239 18372 249273
rect 18243 249223 18372 249239
rect 18663 249273 18792 249289
rect 18663 249239 18679 249273
rect 18775 249239 18792 249273
rect 18663 249223 18792 249239
rect 19083 249273 19212 249289
rect 19083 249239 19099 249273
rect 19195 249239 19212 249273
rect 19083 249223 19212 249239
rect 19503 249273 19632 249289
rect 19503 249239 19519 249273
rect 19615 249239 19632 249273
rect 19503 249223 19632 249239
rect 19923 249273 20052 249289
rect 19923 249239 19939 249273
rect 20035 249239 20052 249273
rect 19923 249223 20052 249239
rect 20343 249273 20472 249289
rect 20343 249239 20359 249273
rect 20455 249239 20472 249273
rect 20343 249223 20472 249239
rect 20763 249273 20892 249289
rect 20763 249239 20779 249273
rect 20875 249239 20892 249273
rect 20763 249223 20892 249239
rect 21183 249273 21312 249289
rect 21183 249239 21199 249273
rect 21295 249239 21312 249273
rect 21183 249223 21312 249239
rect 21603 249273 21732 249289
rect 21603 249239 21619 249273
rect 21715 249239 21732 249273
rect 21603 249223 21732 249239
rect 22023 249273 22152 249289
rect 22023 249239 22039 249273
rect 22135 249239 22152 249273
rect 22023 249223 22152 249239
rect 22443 249273 22572 249289
rect 22443 249239 22459 249273
rect 22555 249239 22572 249273
rect 22443 249223 22572 249239
rect 22863 249273 22992 249289
rect 22863 249239 22879 249273
rect 22975 249239 22992 249273
rect 22863 249223 22992 249239
rect 23283 249273 23412 249289
rect 23283 249239 23299 249273
rect 23395 249239 23412 249273
rect 23283 249223 23412 249239
rect 23703 249273 23832 249289
rect 23703 249239 23719 249273
rect 23815 249239 23832 249273
rect 23703 249223 23832 249239
rect 24123 249273 24252 249289
rect 24123 249239 24139 249273
rect 24235 249239 24252 249273
rect 24123 249223 24252 249239
rect 24543 249273 24672 249289
rect 24543 249239 24559 249273
rect 24655 249239 24672 249273
rect 24543 249223 24672 249239
rect 24963 249273 25092 249289
rect 24963 249239 24979 249273
rect 25075 249239 25092 249273
rect 24963 249223 25092 249239
rect 25383 249273 25512 249289
rect 25383 249239 25399 249273
rect 25495 249239 25512 249273
rect 25383 249223 25512 249239
rect 25803 249273 25932 249289
rect 25803 249239 25819 249273
rect 25915 249239 25932 249273
rect 25803 249223 25932 249239
rect 26223 249273 26352 249289
rect 26223 249239 26239 249273
rect 26335 249239 26352 249273
rect 26223 249223 26352 249239
rect 26643 249273 26772 249289
rect 26643 249239 26659 249273
rect 26755 249239 26772 249273
rect 26643 249223 26772 249239
rect 27063 249273 27192 249289
rect 27063 249239 27079 249273
rect 27175 249239 27192 249273
rect 27063 249223 27192 249239
rect -3999 249192 -3969 249223
rect -3789 249192 -3759 249218
rect -3579 249192 -3549 249223
rect -3369 249192 -3339 249218
rect -3159 249192 -3129 249223
rect -2949 249192 -2919 249218
rect -2739 249192 -2709 249223
rect -2529 249192 -2499 249218
rect -2319 249192 -2289 249223
rect -2109 249192 -2079 249218
rect -1899 249192 -1869 249223
rect -1689 249192 -1659 249218
rect -1479 249192 -1449 249223
rect -1269 249192 -1239 249218
rect -1059 249192 -1029 249223
rect -849 249192 -819 249218
rect -639 249192 -609 249223
rect -429 249192 -399 249218
rect -219 249192 -189 249223
rect -9 249192 21 249218
rect 201 249192 231 249223
rect 411 249192 441 249218
rect 621 249192 651 249223
rect 831 249192 861 249218
rect 1041 249192 1071 249223
rect 1251 249192 1281 249218
rect 1461 249192 1491 249223
rect 1671 249192 1701 249218
rect 1881 249192 1911 249223
rect 2091 249192 2121 249218
rect 2301 249192 2331 249223
rect 2511 249192 2541 249218
rect 2721 249192 2751 249223
rect 2931 249192 2961 249218
rect 3141 249192 3171 249223
rect 3351 249192 3381 249218
rect 3561 249192 3591 249223
rect 3771 249192 3801 249218
rect 3981 249192 4011 249223
rect 4191 249192 4221 249218
rect 4401 249192 4431 249223
rect 4611 249192 4641 249218
rect 4821 249192 4851 249223
rect 5031 249192 5061 249218
rect 5241 249192 5271 249223
rect 5451 249192 5481 249218
rect 5661 249192 5691 249223
rect 5871 249192 5901 249218
rect 6081 249192 6111 249223
rect 6291 249192 6321 249218
rect 6501 249192 6531 249223
rect 6711 249192 6741 249218
rect 6921 249192 6951 249223
rect 7131 249192 7161 249218
rect 7341 249192 7371 249223
rect 7551 249192 7581 249218
rect 7761 249192 7791 249223
rect 7971 249192 8001 249218
rect 8181 249192 8211 249223
rect 8391 249192 8421 249218
rect 8601 249192 8631 249223
rect 8811 249192 8841 249218
rect 9021 249192 9051 249223
rect 9231 249192 9261 249218
rect 9441 249192 9471 249223
rect 9651 249192 9681 249218
rect 9861 249192 9891 249223
rect 10071 249192 10101 249218
rect 10281 249192 10311 249223
rect 10491 249192 10521 249218
rect 10701 249192 10731 249223
rect 10911 249192 10941 249218
rect 11121 249192 11151 249223
rect 11331 249192 11361 249218
rect 11541 249192 11571 249223
rect 11751 249192 11781 249218
rect 11961 249192 11991 249223
rect 12171 249192 12201 249218
rect 12381 249192 12411 249223
rect 12591 249192 12621 249218
rect 12801 249192 12831 249223
rect 13011 249192 13041 249218
rect 13221 249192 13251 249223
rect 13431 249192 13461 249218
rect 13641 249192 13671 249223
rect 13851 249192 13881 249218
rect 14061 249192 14091 249223
rect 14271 249192 14301 249218
rect 14481 249192 14511 249223
rect 14691 249192 14721 249218
rect 14901 249192 14931 249223
rect 15111 249192 15141 249218
rect 15321 249192 15351 249223
rect 15531 249192 15561 249218
rect 15741 249192 15771 249223
rect 15951 249192 15981 249218
rect 16161 249192 16191 249223
rect 16371 249192 16401 249218
rect 16581 249192 16611 249223
rect 16791 249192 16821 249218
rect 17001 249192 17031 249223
rect 17211 249192 17241 249218
rect 17421 249192 17451 249223
rect 17631 249192 17661 249218
rect 17841 249192 17871 249223
rect 18051 249192 18081 249218
rect 18261 249192 18291 249223
rect 18471 249192 18501 249218
rect 18681 249192 18711 249223
rect 18891 249192 18921 249218
rect 19101 249192 19131 249223
rect 19311 249192 19341 249218
rect 19521 249192 19551 249223
rect 19731 249192 19761 249218
rect 19941 249192 19971 249223
rect 20151 249192 20181 249218
rect 20361 249192 20391 249223
rect 20571 249192 20601 249218
rect 20781 249192 20811 249223
rect 20991 249192 21021 249218
rect 21201 249192 21231 249223
rect 21411 249192 21441 249218
rect 21621 249192 21651 249223
rect 21831 249192 21861 249218
rect 22041 249192 22071 249223
rect 22251 249192 22281 249218
rect 22461 249192 22491 249223
rect 22671 249192 22701 249218
rect 22881 249192 22911 249223
rect 23091 249192 23121 249218
rect 23301 249192 23331 249223
rect 23511 249192 23541 249218
rect 23721 249192 23751 249223
rect 23931 249192 23961 249218
rect 24141 249192 24171 249223
rect 24351 249192 24381 249218
rect 24561 249192 24591 249223
rect 24771 249192 24801 249218
rect 24981 249192 25011 249223
rect 25191 249192 25221 249218
rect 25401 249192 25431 249223
rect 25611 249192 25641 249218
rect 25821 249192 25851 249223
rect 26031 249192 26061 249218
rect 26241 249192 26271 249223
rect 26451 249192 26481 249218
rect 26661 249192 26691 249223
rect 26871 249192 26901 249218
rect 27081 249192 27111 249223
rect 27291 249192 27321 249218
rect -3999 248366 -3969 248392
rect -3789 248361 -3759 248392
rect -3579 248366 -3549 248392
rect -3369 248361 -3339 248392
rect -3159 248366 -3129 248392
rect -2949 248361 -2919 248392
rect -2739 248366 -2709 248392
rect -2529 248361 -2499 248392
rect -2319 248366 -2289 248392
rect -2109 248361 -2079 248392
rect -1899 248366 -1869 248392
rect -1689 248361 -1659 248392
rect -1479 248366 -1449 248392
rect -1269 248361 -1239 248392
rect -1059 248366 -1029 248392
rect -849 248361 -819 248392
rect -639 248366 -609 248392
rect -429 248361 -399 248392
rect -219 248366 -189 248392
rect -9 248361 21 248392
rect 201 248366 231 248392
rect 411 248361 441 248392
rect 621 248366 651 248392
rect 831 248361 861 248392
rect 1041 248366 1071 248392
rect 1251 248361 1281 248392
rect 1461 248366 1491 248392
rect 1671 248361 1701 248392
rect 1881 248366 1911 248392
rect 2091 248361 2121 248392
rect 2301 248366 2331 248392
rect 2511 248361 2541 248392
rect 2721 248366 2751 248392
rect 2931 248361 2961 248392
rect 3141 248366 3171 248392
rect 3351 248361 3381 248392
rect 3561 248366 3591 248392
rect 3771 248361 3801 248392
rect 3981 248366 4011 248392
rect 4191 248361 4221 248392
rect 4401 248366 4431 248392
rect 4611 248361 4641 248392
rect 4821 248366 4851 248392
rect 5031 248361 5061 248392
rect 5241 248366 5271 248392
rect 5451 248361 5481 248392
rect 5661 248366 5691 248392
rect 5871 248361 5901 248392
rect 6081 248366 6111 248392
rect 6291 248361 6321 248392
rect 6501 248366 6531 248392
rect 6711 248361 6741 248392
rect 6921 248366 6951 248392
rect 7131 248361 7161 248392
rect 7341 248366 7371 248392
rect 7551 248361 7581 248392
rect 7761 248366 7791 248392
rect 7971 248361 8001 248392
rect 8181 248366 8211 248392
rect 8391 248361 8421 248392
rect 8601 248366 8631 248392
rect 8811 248361 8841 248392
rect 9021 248366 9051 248392
rect 9231 248361 9261 248392
rect 9441 248366 9471 248392
rect 9651 248361 9681 248392
rect 9861 248366 9891 248392
rect 10071 248361 10101 248392
rect 10281 248366 10311 248392
rect 10491 248361 10521 248392
rect 10701 248366 10731 248392
rect 10911 248361 10941 248392
rect 11121 248366 11151 248392
rect 11331 248361 11361 248392
rect 11541 248366 11571 248392
rect 11751 248361 11781 248392
rect 11961 248366 11991 248392
rect 12171 248361 12201 248392
rect 12381 248366 12411 248392
rect 12591 248361 12621 248392
rect 12801 248366 12831 248392
rect 13011 248361 13041 248392
rect 13221 248366 13251 248392
rect 13431 248361 13461 248392
rect 13641 248366 13671 248392
rect 13851 248361 13881 248392
rect 14061 248366 14091 248392
rect 14271 248361 14301 248392
rect 14481 248366 14511 248392
rect 14691 248361 14721 248392
rect 14901 248366 14931 248392
rect 15111 248361 15141 248392
rect 15321 248366 15351 248392
rect 15531 248361 15561 248392
rect 15741 248366 15771 248392
rect 15951 248361 15981 248392
rect 16161 248366 16191 248392
rect 16371 248361 16401 248392
rect 16581 248366 16611 248392
rect 16791 248361 16821 248392
rect 17001 248366 17031 248392
rect 17211 248361 17241 248392
rect 17421 248366 17451 248392
rect 17631 248361 17661 248392
rect 17841 248366 17871 248392
rect 18051 248361 18081 248392
rect 18261 248366 18291 248392
rect 18471 248361 18501 248392
rect 18681 248366 18711 248392
rect 18891 248361 18921 248392
rect 19101 248366 19131 248392
rect 19311 248361 19341 248392
rect 19521 248366 19551 248392
rect 19731 248361 19761 248392
rect 19941 248366 19971 248392
rect 20151 248361 20181 248392
rect 20361 248366 20391 248392
rect 20571 248361 20601 248392
rect 20781 248366 20811 248392
rect 20991 248361 21021 248392
rect 21201 248366 21231 248392
rect 21411 248361 21441 248392
rect 21621 248366 21651 248392
rect 21831 248361 21861 248392
rect 22041 248366 22071 248392
rect 22251 248361 22281 248392
rect 22461 248366 22491 248392
rect 22671 248361 22701 248392
rect 22881 248366 22911 248392
rect 23091 248361 23121 248392
rect 23301 248366 23331 248392
rect 23511 248361 23541 248392
rect 23721 248366 23751 248392
rect 23931 248361 23961 248392
rect 24141 248366 24171 248392
rect 24351 248361 24381 248392
rect 24561 248366 24591 248392
rect 24771 248361 24801 248392
rect 24981 248366 25011 248392
rect 25191 248361 25221 248392
rect 25401 248366 25431 248392
rect 25611 248361 25641 248392
rect 25821 248366 25851 248392
rect 26031 248361 26061 248392
rect 26241 248366 26271 248392
rect 26451 248361 26481 248392
rect 26661 248366 26691 248392
rect 26871 248361 26901 248392
rect 27081 248366 27111 248392
rect 27291 248361 27321 248392
rect -3807 248345 -3741 248361
rect -3807 248203 -3791 248345
rect -3757 248203 -3741 248345
rect -3807 248187 -3741 248203
rect -3387 248345 -3321 248361
rect -3387 248203 -3371 248345
rect -3337 248203 -3321 248345
rect -3387 248187 -3321 248203
rect -2967 248345 -2901 248361
rect -2967 248203 -2951 248345
rect -2917 248203 -2901 248345
rect -2967 248187 -2901 248203
rect -2547 248345 -2481 248361
rect -2547 248203 -2531 248345
rect -2497 248203 -2481 248345
rect -2547 248187 -2481 248203
rect -2127 248345 -2061 248361
rect -2127 248203 -2111 248345
rect -2077 248203 -2061 248345
rect -2127 248187 -2061 248203
rect -1707 248345 -1641 248361
rect -1707 248203 -1691 248345
rect -1657 248203 -1641 248345
rect -1707 248187 -1641 248203
rect -1287 248345 -1221 248361
rect -1287 248203 -1271 248345
rect -1237 248203 -1221 248345
rect -1287 248187 -1221 248203
rect -867 248345 -801 248361
rect -867 248203 -851 248345
rect -817 248203 -801 248345
rect -867 248187 -801 248203
rect -447 248345 -381 248361
rect -447 248203 -431 248345
rect -397 248203 -381 248345
rect -447 248187 -381 248203
rect -27 248345 39 248361
rect -27 248203 -11 248345
rect 23 248203 39 248345
rect -27 248187 39 248203
rect 393 248345 459 248361
rect 393 248203 409 248345
rect 443 248203 459 248345
rect 393 248187 459 248203
rect 813 248345 879 248361
rect 813 248203 829 248345
rect 863 248203 879 248345
rect 813 248187 879 248203
rect 1233 248345 1299 248361
rect 1233 248203 1249 248345
rect 1283 248203 1299 248345
rect 1233 248187 1299 248203
rect 1653 248345 1719 248361
rect 1653 248203 1669 248345
rect 1703 248203 1719 248345
rect 1653 248187 1719 248203
rect 2073 248345 2139 248361
rect 2073 248203 2089 248345
rect 2123 248203 2139 248345
rect 2073 248187 2139 248203
rect 2493 248345 2559 248361
rect 2493 248203 2509 248345
rect 2543 248203 2559 248345
rect 2493 248187 2559 248203
rect 2913 248345 2979 248361
rect 2913 248203 2929 248345
rect 2963 248203 2979 248345
rect 2913 248187 2979 248203
rect 3333 248345 3399 248361
rect 3333 248203 3349 248345
rect 3383 248203 3399 248345
rect 3333 248187 3399 248203
rect 3753 248345 3819 248361
rect 3753 248203 3769 248345
rect 3803 248203 3819 248345
rect 3753 248187 3819 248203
rect 4173 248345 4239 248361
rect 4173 248203 4189 248345
rect 4223 248203 4239 248345
rect 4173 248187 4239 248203
rect 4593 248345 4659 248361
rect 4593 248203 4609 248345
rect 4643 248203 4659 248345
rect 4593 248187 4659 248203
rect 5013 248345 5079 248361
rect 5013 248203 5029 248345
rect 5063 248203 5079 248345
rect 5013 248187 5079 248203
rect 5433 248345 5499 248361
rect 5433 248203 5449 248345
rect 5483 248203 5499 248345
rect 5433 248187 5499 248203
rect 5853 248345 5919 248361
rect 5853 248203 5869 248345
rect 5903 248203 5919 248345
rect 5853 248187 5919 248203
rect 6273 248345 6339 248361
rect 6273 248203 6289 248345
rect 6323 248203 6339 248345
rect 6273 248187 6339 248203
rect 6693 248345 6759 248361
rect 6693 248203 6709 248345
rect 6743 248203 6759 248345
rect 6693 248187 6759 248203
rect 7113 248345 7179 248361
rect 7113 248203 7129 248345
rect 7163 248203 7179 248345
rect 7113 248187 7179 248203
rect 7533 248345 7599 248361
rect 7533 248203 7549 248345
rect 7583 248203 7599 248345
rect 7533 248187 7599 248203
rect 7953 248345 8019 248361
rect 7953 248203 7969 248345
rect 8003 248203 8019 248345
rect 7953 248187 8019 248203
rect 8373 248345 8439 248361
rect 8373 248203 8389 248345
rect 8423 248203 8439 248345
rect 8373 248187 8439 248203
rect 8793 248345 8859 248361
rect 8793 248203 8809 248345
rect 8843 248203 8859 248345
rect 8793 248187 8859 248203
rect 9213 248345 9279 248361
rect 9213 248203 9229 248345
rect 9263 248203 9279 248345
rect 9213 248187 9279 248203
rect 9633 248345 9699 248361
rect 9633 248203 9649 248345
rect 9683 248203 9699 248345
rect 9633 248187 9699 248203
rect 10053 248345 10119 248361
rect 10053 248203 10069 248345
rect 10103 248203 10119 248345
rect 10053 248187 10119 248203
rect 10473 248345 10539 248361
rect 10473 248203 10489 248345
rect 10523 248203 10539 248345
rect 10473 248187 10539 248203
rect 10893 248345 10959 248361
rect 10893 248203 10909 248345
rect 10943 248203 10959 248345
rect 10893 248187 10959 248203
rect 11313 248345 11379 248361
rect 11313 248203 11329 248345
rect 11363 248203 11379 248345
rect 11313 248187 11379 248203
rect 11733 248345 11799 248361
rect 11733 248203 11749 248345
rect 11783 248203 11799 248345
rect 11733 248187 11799 248203
rect 12153 248345 12219 248361
rect 12153 248203 12169 248345
rect 12203 248203 12219 248345
rect 12153 248187 12219 248203
rect 12573 248345 12639 248361
rect 12573 248203 12589 248345
rect 12623 248203 12639 248345
rect 12573 248187 12639 248203
rect 12993 248345 13059 248361
rect 12993 248203 13009 248345
rect 13043 248203 13059 248345
rect 12993 248187 13059 248203
rect 13413 248345 13479 248361
rect 13413 248203 13429 248345
rect 13463 248203 13479 248345
rect 13413 248187 13479 248203
rect 13833 248345 13899 248361
rect 13833 248203 13849 248345
rect 13883 248203 13899 248345
rect 13833 248187 13899 248203
rect 14253 248345 14319 248361
rect 14253 248203 14269 248345
rect 14303 248203 14319 248345
rect 14253 248187 14319 248203
rect 14673 248345 14739 248361
rect 14673 248203 14689 248345
rect 14723 248203 14739 248345
rect 14673 248187 14739 248203
rect 15093 248345 15159 248361
rect 15093 248203 15109 248345
rect 15143 248203 15159 248345
rect 15093 248187 15159 248203
rect 15513 248345 15579 248361
rect 15513 248203 15529 248345
rect 15563 248203 15579 248345
rect 15513 248187 15579 248203
rect 15933 248345 15999 248361
rect 15933 248203 15949 248345
rect 15983 248203 15999 248345
rect 15933 248187 15999 248203
rect 16353 248345 16419 248361
rect 16353 248203 16369 248345
rect 16403 248203 16419 248345
rect 16353 248187 16419 248203
rect 16773 248345 16839 248361
rect 16773 248203 16789 248345
rect 16823 248203 16839 248345
rect 16773 248187 16839 248203
rect 17193 248345 17259 248361
rect 17193 248203 17209 248345
rect 17243 248203 17259 248345
rect 17193 248187 17259 248203
rect 17613 248345 17679 248361
rect 17613 248203 17629 248345
rect 17663 248203 17679 248345
rect 17613 248187 17679 248203
rect 18033 248345 18099 248361
rect 18033 248203 18049 248345
rect 18083 248203 18099 248345
rect 18033 248187 18099 248203
rect 18453 248345 18519 248361
rect 18453 248203 18469 248345
rect 18503 248203 18519 248345
rect 18453 248187 18519 248203
rect 18873 248345 18939 248361
rect 18873 248203 18889 248345
rect 18923 248203 18939 248345
rect 18873 248187 18939 248203
rect 19293 248345 19359 248361
rect 19293 248203 19309 248345
rect 19343 248203 19359 248345
rect 19293 248187 19359 248203
rect 19713 248345 19779 248361
rect 19713 248203 19729 248345
rect 19763 248203 19779 248345
rect 19713 248187 19779 248203
rect 20133 248345 20199 248361
rect 20133 248203 20149 248345
rect 20183 248203 20199 248345
rect 20133 248187 20199 248203
rect 20553 248345 20619 248361
rect 20553 248203 20569 248345
rect 20603 248203 20619 248345
rect 20553 248187 20619 248203
rect 20973 248345 21039 248361
rect 20973 248203 20989 248345
rect 21023 248203 21039 248345
rect 20973 248187 21039 248203
rect 21393 248345 21459 248361
rect 21393 248203 21409 248345
rect 21443 248203 21459 248345
rect 21393 248187 21459 248203
rect 21813 248345 21879 248361
rect 21813 248203 21829 248345
rect 21863 248203 21879 248345
rect 21813 248187 21879 248203
rect 22233 248345 22299 248361
rect 22233 248203 22249 248345
rect 22283 248203 22299 248345
rect 22233 248187 22299 248203
rect 22653 248345 22719 248361
rect 22653 248203 22669 248345
rect 22703 248203 22719 248345
rect 22653 248187 22719 248203
rect 23073 248345 23139 248361
rect 23073 248203 23089 248345
rect 23123 248203 23139 248345
rect 23073 248187 23139 248203
rect 23493 248345 23559 248361
rect 23493 248203 23509 248345
rect 23543 248203 23559 248345
rect 23493 248187 23559 248203
rect 23913 248345 23979 248361
rect 23913 248203 23929 248345
rect 23963 248203 23979 248345
rect 23913 248187 23979 248203
rect 24333 248345 24399 248361
rect 24333 248203 24349 248345
rect 24383 248203 24399 248345
rect 24333 248187 24399 248203
rect 24753 248345 24819 248361
rect 24753 248203 24769 248345
rect 24803 248203 24819 248345
rect 24753 248187 24819 248203
rect 25173 248345 25239 248361
rect 25173 248203 25189 248345
rect 25223 248203 25239 248345
rect 25173 248187 25239 248203
rect 25593 248345 25659 248361
rect 25593 248203 25609 248345
rect 25643 248203 25659 248345
rect 25593 248187 25659 248203
rect 26013 248345 26079 248361
rect 26013 248203 26029 248345
rect 26063 248203 26079 248345
rect 26013 248187 26079 248203
rect 26433 248345 26499 248361
rect 26433 248203 26449 248345
rect 26483 248203 26499 248345
rect 26433 248187 26499 248203
rect 26853 248345 26919 248361
rect 26853 248203 26869 248345
rect 26903 248203 26919 248345
rect 26853 248187 26919 248203
rect 27273 248345 27339 248361
rect 27273 248203 27289 248345
rect 27323 248203 27339 248345
rect 27273 248187 27339 248203
rect -3999 248156 -3969 248182
rect -3789 248156 -3759 248187
rect -3579 248156 -3549 248182
rect -3369 248156 -3339 248187
rect -3159 248156 -3129 248182
rect -2949 248156 -2919 248187
rect -2739 248156 -2709 248182
rect -2529 248156 -2499 248187
rect -2319 248156 -2289 248182
rect -2109 248156 -2079 248187
rect -1899 248156 -1869 248182
rect -1689 248156 -1659 248187
rect -1479 248156 -1449 248182
rect -1269 248156 -1239 248187
rect -1059 248156 -1029 248182
rect -849 248156 -819 248187
rect -639 248156 -609 248182
rect -429 248156 -399 248187
rect -219 248156 -189 248182
rect -9 248156 21 248187
rect 201 248156 231 248182
rect 411 248156 441 248187
rect 621 248156 651 248182
rect 831 248156 861 248187
rect 1041 248156 1071 248182
rect 1251 248156 1281 248187
rect 1461 248156 1491 248182
rect 1671 248156 1701 248187
rect 1881 248156 1911 248182
rect 2091 248156 2121 248187
rect 2301 248156 2331 248182
rect 2511 248156 2541 248187
rect 2721 248156 2751 248182
rect 2931 248156 2961 248187
rect 3141 248156 3171 248182
rect 3351 248156 3381 248187
rect 3561 248156 3591 248182
rect 3771 248156 3801 248187
rect 3981 248156 4011 248182
rect 4191 248156 4221 248187
rect 4401 248156 4431 248182
rect 4611 248156 4641 248187
rect 4821 248156 4851 248182
rect 5031 248156 5061 248187
rect 5241 248156 5271 248182
rect 5451 248156 5481 248187
rect 5661 248156 5691 248182
rect 5871 248156 5901 248187
rect 6081 248156 6111 248182
rect 6291 248156 6321 248187
rect 6501 248156 6531 248182
rect 6711 248156 6741 248187
rect 6921 248156 6951 248182
rect 7131 248156 7161 248187
rect 7341 248156 7371 248182
rect 7551 248156 7581 248187
rect 7761 248156 7791 248182
rect 7971 248156 8001 248187
rect 8181 248156 8211 248182
rect 8391 248156 8421 248187
rect 8601 248156 8631 248182
rect 8811 248156 8841 248187
rect 9021 248156 9051 248182
rect 9231 248156 9261 248187
rect 9441 248156 9471 248182
rect 9651 248156 9681 248187
rect 9861 248156 9891 248182
rect 10071 248156 10101 248187
rect 10281 248156 10311 248182
rect 10491 248156 10521 248187
rect 10701 248156 10731 248182
rect 10911 248156 10941 248187
rect 11121 248156 11151 248182
rect 11331 248156 11361 248187
rect 11541 248156 11571 248182
rect 11751 248156 11781 248187
rect 11961 248156 11991 248182
rect 12171 248156 12201 248187
rect 12381 248156 12411 248182
rect 12591 248156 12621 248187
rect 12801 248156 12831 248182
rect 13011 248156 13041 248187
rect 13221 248156 13251 248182
rect 13431 248156 13461 248187
rect 13641 248156 13671 248182
rect 13851 248156 13881 248187
rect 14061 248156 14091 248182
rect 14271 248156 14301 248187
rect 14481 248156 14511 248182
rect 14691 248156 14721 248187
rect 14901 248156 14931 248182
rect 15111 248156 15141 248187
rect 15321 248156 15351 248182
rect 15531 248156 15561 248187
rect 15741 248156 15771 248182
rect 15951 248156 15981 248187
rect 16161 248156 16191 248182
rect 16371 248156 16401 248187
rect 16581 248156 16611 248182
rect 16791 248156 16821 248187
rect 17001 248156 17031 248182
rect 17211 248156 17241 248187
rect 17421 248156 17451 248182
rect 17631 248156 17661 248187
rect 17841 248156 17871 248182
rect 18051 248156 18081 248187
rect 18261 248156 18291 248182
rect 18471 248156 18501 248187
rect 18681 248156 18711 248182
rect 18891 248156 18921 248187
rect 19101 248156 19131 248182
rect 19311 248156 19341 248187
rect 19521 248156 19551 248182
rect 19731 248156 19761 248187
rect 19941 248156 19971 248182
rect 20151 248156 20181 248187
rect 20361 248156 20391 248182
rect 20571 248156 20601 248187
rect 20781 248156 20811 248182
rect 20991 248156 21021 248187
rect 21201 248156 21231 248182
rect 21411 248156 21441 248187
rect 21621 248156 21651 248182
rect 21831 248156 21861 248187
rect 22041 248156 22071 248182
rect 22251 248156 22281 248187
rect 22461 248156 22491 248182
rect 22671 248156 22701 248187
rect 22881 248156 22911 248182
rect 23091 248156 23121 248187
rect 23301 248156 23331 248182
rect 23511 248156 23541 248187
rect 23721 248156 23751 248182
rect 23931 248156 23961 248187
rect 24141 248156 24171 248182
rect 24351 248156 24381 248187
rect 24561 248156 24591 248182
rect 24771 248156 24801 248187
rect 24981 248156 25011 248182
rect 25191 248156 25221 248187
rect 25401 248156 25431 248182
rect 25611 248156 25641 248187
rect 25821 248156 25851 248182
rect 26031 248156 26061 248187
rect 26241 248156 26271 248182
rect 26451 248156 26481 248187
rect 26661 248156 26691 248182
rect 26871 248156 26901 248187
rect 27081 248156 27111 248182
rect 27291 248156 27321 248187
rect -3999 247325 -3969 247356
rect -3789 247330 -3759 247356
rect -3579 247325 -3549 247356
rect -3369 247330 -3339 247356
rect -3159 247325 -3129 247356
rect -2949 247330 -2919 247356
rect -2739 247325 -2709 247356
rect -2529 247330 -2499 247356
rect -2319 247325 -2289 247356
rect -2109 247330 -2079 247356
rect -1899 247325 -1869 247356
rect -1689 247330 -1659 247356
rect -1479 247325 -1449 247356
rect -1269 247330 -1239 247356
rect -1059 247325 -1029 247356
rect -849 247330 -819 247356
rect -639 247325 -609 247356
rect -429 247330 -399 247356
rect -219 247325 -189 247356
rect -9 247330 21 247356
rect 201 247325 231 247356
rect 411 247330 441 247356
rect 621 247325 651 247356
rect 831 247330 861 247356
rect 1041 247325 1071 247356
rect 1251 247330 1281 247356
rect 1461 247325 1491 247356
rect 1671 247330 1701 247356
rect 1881 247325 1911 247356
rect 2091 247330 2121 247356
rect 2301 247325 2331 247356
rect 2511 247330 2541 247356
rect 2721 247325 2751 247356
rect 2931 247330 2961 247356
rect 3141 247325 3171 247356
rect 3351 247330 3381 247356
rect 3561 247325 3591 247356
rect 3771 247330 3801 247356
rect 3981 247325 4011 247356
rect 4191 247330 4221 247356
rect 4401 247325 4431 247356
rect 4611 247330 4641 247356
rect 4821 247325 4851 247356
rect 5031 247330 5061 247356
rect 5241 247325 5271 247356
rect 5451 247330 5481 247356
rect 5661 247325 5691 247356
rect 5871 247330 5901 247356
rect 6081 247325 6111 247356
rect 6291 247330 6321 247356
rect 6501 247325 6531 247356
rect 6711 247330 6741 247356
rect 6921 247325 6951 247356
rect 7131 247330 7161 247356
rect 7341 247325 7371 247356
rect 7551 247330 7581 247356
rect 7761 247325 7791 247356
rect 7971 247330 8001 247356
rect 8181 247325 8211 247356
rect 8391 247330 8421 247356
rect 8601 247325 8631 247356
rect 8811 247330 8841 247356
rect 9021 247325 9051 247356
rect 9231 247330 9261 247356
rect 9441 247325 9471 247356
rect 9651 247330 9681 247356
rect 9861 247325 9891 247356
rect 10071 247330 10101 247356
rect 10281 247325 10311 247356
rect 10491 247330 10521 247356
rect 10701 247325 10731 247356
rect 10911 247330 10941 247356
rect 11121 247325 11151 247356
rect 11331 247330 11361 247356
rect 11541 247325 11571 247356
rect 11751 247330 11781 247356
rect 11961 247325 11991 247356
rect 12171 247330 12201 247356
rect 12381 247325 12411 247356
rect 12591 247330 12621 247356
rect 12801 247325 12831 247356
rect 13011 247330 13041 247356
rect 13221 247325 13251 247356
rect 13431 247330 13461 247356
rect 13641 247325 13671 247356
rect 13851 247330 13881 247356
rect 14061 247325 14091 247356
rect 14271 247330 14301 247356
rect 14481 247325 14511 247356
rect 14691 247330 14721 247356
rect 14901 247325 14931 247356
rect 15111 247330 15141 247356
rect 15321 247325 15351 247356
rect 15531 247330 15561 247356
rect 15741 247325 15771 247356
rect 15951 247330 15981 247356
rect 16161 247325 16191 247356
rect 16371 247330 16401 247356
rect 16581 247325 16611 247356
rect 16791 247330 16821 247356
rect 17001 247325 17031 247356
rect 17211 247330 17241 247356
rect 17421 247325 17451 247356
rect 17631 247330 17661 247356
rect 17841 247325 17871 247356
rect 18051 247330 18081 247356
rect 18261 247325 18291 247356
rect 18471 247330 18501 247356
rect 18681 247325 18711 247356
rect 18891 247330 18921 247356
rect 19101 247325 19131 247356
rect 19311 247330 19341 247356
rect 19521 247325 19551 247356
rect 19731 247330 19761 247356
rect 19941 247325 19971 247356
rect 20151 247330 20181 247356
rect 20361 247325 20391 247356
rect 20571 247330 20601 247356
rect 20781 247325 20811 247356
rect 20991 247330 21021 247356
rect 21201 247325 21231 247356
rect 21411 247330 21441 247356
rect 21621 247325 21651 247356
rect 21831 247330 21861 247356
rect 22041 247325 22071 247356
rect 22251 247330 22281 247356
rect 22461 247325 22491 247356
rect 22671 247330 22701 247356
rect 22881 247325 22911 247356
rect 23091 247330 23121 247356
rect 23301 247325 23331 247356
rect 23511 247330 23541 247356
rect 23721 247325 23751 247356
rect 23931 247330 23961 247356
rect 24141 247325 24171 247356
rect 24351 247330 24381 247356
rect 24561 247325 24591 247356
rect 24771 247330 24801 247356
rect 24981 247325 25011 247356
rect 25191 247330 25221 247356
rect 25401 247325 25431 247356
rect 25611 247330 25641 247356
rect 25821 247325 25851 247356
rect 26031 247330 26061 247356
rect 26241 247325 26271 247356
rect 26451 247330 26481 247356
rect 26661 247325 26691 247356
rect 26871 247330 26901 247356
rect 27081 247325 27111 247356
rect 27291 247330 27321 247356
rect -4017 247309 -3951 247325
rect -4017 247167 -4001 247309
rect -3967 247167 -3951 247309
rect -4017 247151 -3951 247167
rect -3597 247309 -3531 247325
rect -3597 247167 -3581 247309
rect -3547 247167 -3531 247309
rect -3597 247151 -3531 247167
rect -3177 247309 -3111 247325
rect -3177 247167 -3161 247309
rect -3127 247167 -3111 247309
rect -3177 247151 -3111 247167
rect -2757 247309 -2691 247325
rect -2757 247167 -2741 247309
rect -2707 247167 -2691 247309
rect -2757 247151 -2691 247167
rect -2337 247309 -2271 247325
rect -2337 247167 -2321 247309
rect -2287 247167 -2271 247309
rect -2337 247151 -2271 247167
rect -1917 247309 -1851 247325
rect -1917 247167 -1901 247309
rect -1867 247167 -1851 247309
rect -1917 247151 -1851 247167
rect -1497 247309 -1431 247325
rect -1497 247167 -1481 247309
rect -1447 247167 -1431 247309
rect -1497 247151 -1431 247167
rect -1077 247309 -1011 247325
rect -1077 247167 -1061 247309
rect -1027 247167 -1011 247309
rect -1077 247151 -1011 247167
rect -657 247309 -591 247325
rect -657 247167 -641 247309
rect -607 247167 -591 247309
rect -657 247151 -591 247167
rect -237 247309 -171 247325
rect -237 247167 -221 247309
rect -187 247167 -171 247309
rect -237 247151 -171 247167
rect 183 247309 249 247325
rect 183 247167 199 247309
rect 233 247167 249 247309
rect 183 247151 249 247167
rect 603 247309 669 247325
rect 603 247167 619 247309
rect 653 247167 669 247309
rect 603 247151 669 247167
rect 1023 247309 1089 247325
rect 1023 247167 1039 247309
rect 1073 247167 1089 247309
rect 1023 247151 1089 247167
rect 1443 247309 1509 247325
rect 1443 247167 1459 247309
rect 1493 247167 1509 247309
rect 1443 247151 1509 247167
rect 1863 247309 1929 247325
rect 1863 247167 1879 247309
rect 1913 247167 1929 247309
rect 1863 247151 1929 247167
rect 2283 247309 2349 247325
rect 2283 247167 2299 247309
rect 2333 247167 2349 247309
rect 2283 247151 2349 247167
rect 2703 247309 2769 247325
rect 2703 247167 2719 247309
rect 2753 247167 2769 247309
rect 2703 247151 2769 247167
rect 3123 247309 3189 247325
rect 3123 247167 3139 247309
rect 3173 247167 3189 247309
rect 3123 247151 3189 247167
rect 3543 247309 3609 247325
rect 3543 247167 3559 247309
rect 3593 247167 3609 247309
rect 3543 247151 3609 247167
rect 3963 247309 4029 247325
rect 3963 247167 3979 247309
rect 4013 247167 4029 247309
rect 3963 247151 4029 247167
rect 4383 247309 4449 247325
rect 4383 247167 4399 247309
rect 4433 247167 4449 247309
rect 4383 247151 4449 247167
rect 4803 247309 4869 247325
rect 4803 247167 4819 247309
rect 4853 247167 4869 247309
rect 4803 247151 4869 247167
rect 5223 247309 5289 247325
rect 5223 247167 5239 247309
rect 5273 247167 5289 247309
rect 5223 247151 5289 247167
rect 5643 247309 5709 247325
rect 5643 247167 5659 247309
rect 5693 247167 5709 247309
rect 5643 247151 5709 247167
rect 6063 247309 6129 247325
rect 6063 247167 6079 247309
rect 6113 247167 6129 247309
rect 6063 247151 6129 247167
rect 6483 247309 6549 247325
rect 6483 247167 6499 247309
rect 6533 247167 6549 247309
rect 6483 247151 6549 247167
rect 6903 247309 6969 247325
rect 6903 247167 6919 247309
rect 6953 247167 6969 247309
rect 6903 247151 6969 247167
rect 7323 247309 7389 247325
rect 7323 247167 7339 247309
rect 7373 247167 7389 247309
rect 7323 247151 7389 247167
rect 7743 247309 7809 247325
rect 7743 247167 7759 247309
rect 7793 247167 7809 247309
rect 7743 247151 7809 247167
rect 8163 247309 8229 247325
rect 8163 247167 8179 247309
rect 8213 247167 8229 247309
rect 8163 247151 8229 247167
rect 8583 247309 8649 247325
rect 8583 247167 8599 247309
rect 8633 247167 8649 247309
rect 8583 247151 8649 247167
rect 9003 247309 9069 247325
rect 9003 247167 9019 247309
rect 9053 247167 9069 247309
rect 9003 247151 9069 247167
rect 9423 247309 9489 247325
rect 9423 247167 9439 247309
rect 9473 247167 9489 247309
rect 9423 247151 9489 247167
rect 9843 247309 9909 247325
rect 9843 247167 9859 247309
rect 9893 247167 9909 247309
rect 9843 247151 9909 247167
rect 10263 247309 10329 247325
rect 10263 247167 10279 247309
rect 10313 247167 10329 247309
rect 10263 247151 10329 247167
rect 10683 247309 10749 247325
rect 10683 247167 10699 247309
rect 10733 247167 10749 247309
rect 10683 247151 10749 247167
rect 11103 247309 11169 247325
rect 11103 247167 11119 247309
rect 11153 247167 11169 247309
rect 11103 247151 11169 247167
rect 11523 247309 11589 247325
rect 11523 247167 11539 247309
rect 11573 247167 11589 247309
rect 11523 247151 11589 247167
rect 11943 247309 12009 247325
rect 11943 247167 11959 247309
rect 11993 247167 12009 247309
rect 11943 247151 12009 247167
rect 12363 247309 12429 247325
rect 12363 247167 12379 247309
rect 12413 247167 12429 247309
rect 12363 247151 12429 247167
rect 12783 247309 12849 247325
rect 12783 247167 12799 247309
rect 12833 247167 12849 247309
rect 12783 247151 12849 247167
rect 13203 247309 13269 247325
rect 13203 247167 13219 247309
rect 13253 247167 13269 247309
rect 13203 247151 13269 247167
rect 13623 247309 13689 247325
rect 13623 247167 13639 247309
rect 13673 247167 13689 247309
rect 13623 247151 13689 247167
rect 14043 247309 14109 247325
rect 14043 247167 14059 247309
rect 14093 247167 14109 247309
rect 14043 247151 14109 247167
rect 14463 247309 14529 247325
rect 14463 247167 14479 247309
rect 14513 247167 14529 247309
rect 14463 247151 14529 247167
rect 14883 247309 14949 247325
rect 14883 247167 14899 247309
rect 14933 247167 14949 247309
rect 14883 247151 14949 247167
rect 15303 247309 15369 247325
rect 15303 247167 15319 247309
rect 15353 247167 15369 247309
rect 15303 247151 15369 247167
rect 15723 247309 15789 247325
rect 15723 247167 15739 247309
rect 15773 247167 15789 247309
rect 15723 247151 15789 247167
rect 16143 247309 16209 247325
rect 16143 247167 16159 247309
rect 16193 247167 16209 247309
rect 16143 247151 16209 247167
rect 16563 247309 16629 247325
rect 16563 247167 16579 247309
rect 16613 247167 16629 247309
rect 16563 247151 16629 247167
rect 16983 247309 17049 247325
rect 16983 247167 16999 247309
rect 17033 247167 17049 247309
rect 16983 247151 17049 247167
rect 17403 247309 17469 247325
rect 17403 247167 17419 247309
rect 17453 247167 17469 247309
rect 17403 247151 17469 247167
rect 17823 247309 17889 247325
rect 17823 247167 17839 247309
rect 17873 247167 17889 247309
rect 17823 247151 17889 247167
rect 18243 247309 18309 247325
rect 18243 247167 18259 247309
rect 18293 247167 18309 247309
rect 18243 247151 18309 247167
rect 18663 247309 18729 247325
rect 18663 247167 18679 247309
rect 18713 247167 18729 247309
rect 18663 247151 18729 247167
rect 19083 247309 19149 247325
rect 19083 247167 19099 247309
rect 19133 247167 19149 247309
rect 19083 247151 19149 247167
rect 19503 247309 19569 247325
rect 19503 247167 19519 247309
rect 19553 247167 19569 247309
rect 19503 247151 19569 247167
rect 19923 247309 19989 247325
rect 19923 247167 19939 247309
rect 19973 247167 19989 247309
rect 19923 247151 19989 247167
rect 20343 247309 20409 247325
rect 20343 247167 20359 247309
rect 20393 247167 20409 247309
rect 20343 247151 20409 247167
rect 20763 247309 20829 247325
rect 20763 247167 20779 247309
rect 20813 247167 20829 247309
rect 20763 247151 20829 247167
rect 21183 247309 21249 247325
rect 21183 247167 21199 247309
rect 21233 247167 21249 247309
rect 21183 247151 21249 247167
rect 21603 247309 21669 247325
rect 21603 247167 21619 247309
rect 21653 247167 21669 247309
rect 21603 247151 21669 247167
rect 22023 247309 22089 247325
rect 22023 247167 22039 247309
rect 22073 247167 22089 247309
rect 22023 247151 22089 247167
rect 22443 247309 22509 247325
rect 22443 247167 22459 247309
rect 22493 247167 22509 247309
rect 22443 247151 22509 247167
rect 22863 247309 22929 247325
rect 22863 247167 22879 247309
rect 22913 247167 22929 247309
rect 22863 247151 22929 247167
rect 23283 247309 23349 247325
rect 23283 247167 23299 247309
rect 23333 247167 23349 247309
rect 23283 247151 23349 247167
rect 23703 247309 23769 247325
rect 23703 247167 23719 247309
rect 23753 247167 23769 247309
rect 23703 247151 23769 247167
rect 24123 247309 24189 247325
rect 24123 247167 24139 247309
rect 24173 247167 24189 247309
rect 24123 247151 24189 247167
rect 24543 247309 24609 247325
rect 24543 247167 24559 247309
rect 24593 247167 24609 247309
rect 24543 247151 24609 247167
rect 24963 247309 25029 247325
rect 24963 247167 24979 247309
rect 25013 247167 25029 247309
rect 24963 247151 25029 247167
rect 25383 247309 25449 247325
rect 25383 247167 25399 247309
rect 25433 247167 25449 247309
rect 25383 247151 25449 247167
rect 25803 247309 25869 247325
rect 25803 247167 25819 247309
rect 25853 247167 25869 247309
rect 25803 247151 25869 247167
rect 26223 247309 26289 247325
rect 26223 247167 26239 247309
rect 26273 247167 26289 247309
rect 26223 247151 26289 247167
rect 26643 247309 26709 247325
rect 26643 247167 26659 247309
rect 26693 247167 26709 247309
rect 26643 247151 26709 247167
rect 27063 247309 27129 247325
rect 27063 247167 27079 247309
rect 27113 247167 27129 247309
rect 27063 247151 27129 247167
rect -3999 247120 -3969 247151
rect -3789 247120 -3759 247146
rect -3579 247120 -3549 247151
rect -3369 247120 -3339 247146
rect -3159 247120 -3129 247151
rect -2949 247120 -2919 247146
rect -2739 247120 -2709 247151
rect -2529 247120 -2499 247146
rect -2319 247120 -2289 247151
rect -2109 247120 -2079 247146
rect -1899 247120 -1869 247151
rect -1689 247120 -1659 247146
rect -1479 247120 -1449 247151
rect -1269 247120 -1239 247146
rect -1059 247120 -1029 247151
rect -849 247120 -819 247146
rect -639 247120 -609 247151
rect -429 247120 -399 247146
rect -219 247120 -189 247151
rect -9 247120 21 247146
rect 201 247120 231 247151
rect 411 247120 441 247146
rect 621 247120 651 247151
rect 831 247120 861 247146
rect 1041 247120 1071 247151
rect 1251 247120 1281 247146
rect 1461 247120 1491 247151
rect 1671 247120 1701 247146
rect 1881 247120 1911 247151
rect 2091 247120 2121 247146
rect 2301 247120 2331 247151
rect 2511 247120 2541 247146
rect 2721 247120 2751 247151
rect 2931 247120 2961 247146
rect 3141 247120 3171 247151
rect 3351 247120 3381 247146
rect 3561 247120 3591 247151
rect 3771 247120 3801 247146
rect 3981 247120 4011 247151
rect 4191 247120 4221 247146
rect 4401 247120 4431 247151
rect 4611 247120 4641 247146
rect 4821 247120 4851 247151
rect 5031 247120 5061 247146
rect 5241 247120 5271 247151
rect 5451 247120 5481 247146
rect 5661 247120 5691 247151
rect 5871 247120 5901 247146
rect 6081 247120 6111 247151
rect 6291 247120 6321 247146
rect 6501 247120 6531 247151
rect 6711 247120 6741 247146
rect 6921 247120 6951 247151
rect 7131 247120 7161 247146
rect 7341 247120 7371 247151
rect 7551 247120 7581 247146
rect 7761 247120 7791 247151
rect 7971 247120 8001 247146
rect 8181 247120 8211 247151
rect 8391 247120 8421 247146
rect 8601 247120 8631 247151
rect 8811 247120 8841 247146
rect 9021 247120 9051 247151
rect 9231 247120 9261 247146
rect 9441 247120 9471 247151
rect 9651 247120 9681 247146
rect 9861 247120 9891 247151
rect 10071 247120 10101 247146
rect 10281 247120 10311 247151
rect 10491 247120 10521 247146
rect 10701 247120 10731 247151
rect 10911 247120 10941 247146
rect 11121 247120 11151 247151
rect 11331 247120 11361 247146
rect 11541 247120 11571 247151
rect 11751 247120 11781 247146
rect 11961 247120 11991 247151
rect 12171 247120 12201 247146
rect 12381 247120 12411 247151
rect 12591 247120 12621 247146
rect 12801 247120 12831 247151
rect 13011 247120 13041 247146
rect 13221 247120 13251 247151
rect 13431 247120 13461 247146
rect 13641 247120 13671 247151
rect 13851 247120 13881 247146
rect 14061 247120 14091 247151
rect 14271 247120 14301 247146
rect 14481 247120 14511 247151
rect 14691 247120 14721 247146
rect 14901 247120 14931 247151
rect 15111 247120 15141 247146
rect 15321 247120 15351 247151
rect 15531 247120 15561 247146
rect 15741 247120 15771 247151
rect 15951 247120 15981 247146
rect 16161 247120 16191 247151
rect 16371 247120 16401 247146
rect 16581 247120 16611 247151
rect 16791 247120 16821 247146
rect 17001 247120 17031 247151
rect 17211 247120 17241 247146
rect 17421 247120 17451 247151
rect 17631 247120 17661 247146
rect 17841 247120 17871 247151
rect 18051 247120 18081 247146
rect 18261 247120 18291 247151
rect 18471 247120 18501 247146
rect 18681 247120 18711 247151
rect 18891 247120 18921 247146
rect 19101 247120 19131 247151
rect 19311 247120 19341 247146
rect 19521 247120 19551 247151
rect 19731 247120 19761 247146
rect 19941 247120 19971 247151
rect 20151 247120 20181 247146
rect 20361 247120 20391 247151
rect 20571 247120 20601 247146
rect 20781 247120 20811 247151
rect 20991 247120 21021 247146
rect 21201 247120 21231 247151
rect 21411 247120 21441 247146
rect 21621 247120 21651 247151
rect 21831 247120 21861 247146
rect 22041 247120 22071 247151
rect 22251 247120 22281 247146
rect 22461 247120 22491 247151
rect 22671 247120 22701 247146
rect 22881 247120 22911 247151
rect 23091 247120 23121 247146
rect 23301 247120 23331 247151
rect 23511 247120 23541 247146
rect 23721 247120 23751 247151
rect 23931 247120 23961 247146
rect 24141 247120 24171 247151
rect 24351 247120 24381 247146
rect 24561 247120 24591 247151
rect 24771 247120 24801 247146
rect 24981 247120 25011 247151
rect 25191 247120 25221 247146
rect 25401 247120 25431 247151
rect 25611 247120 25641 247146
rect 25821 247120 25851 247151
rect 26031 247120 26061 247146
rect 26241 247120 26271 247151
rect 26451 247120 26481 247146
rect 26661 247120 26691 247151
rect 26871 247120 26901 247146
rect 27081 247120 27111 247151
rect 27291 247120 27321 247146
rect -3999 246294 -3969 246320
rect -3789 246289 -3759 246320
rect -3579 246294 -3549 246320
rect -3369 246289 -3339 246320
rect -3159 246294 -3129 246320
rect -2949 246289 -2919 246320
rect -2739 246294 -2709 246320
rect -2529 246289 -2499 246320
rect -2319 246294 -2289 246320
rect -2109 246289 -2079 246320
rect -1899 246294 -1869 246320
rect -1689 246289 -1659 246320
rect -1479 246294 -1449 246320
rect -1269 246289 -1239 246320
rect -1059 246294 -1029 246320
rect -849 246289 -819 246320
rect -639 246294 -609 246320
rect -429 246289 -399 246320
rect -219 246294 -189 246320
rect -9 246289 21 246320
rect 201 246294 231 246320
rect 411 246289 441 246320
rect 621 246294 651 246320
rect 831 246289 861 246320
rect 1041 246294 1071 246320
rect 1251 246289 1281 246320
rect 1461 246294 1491 246320
rect 1671 246289 1701 246320
rect 1881 246294 1911 246320
rect 2091 246289 2121 246320
rect 2301 246294 2331 246320
rect 2511 246289 2541 246320
rect 2721 246294 2751 246320
rect 2931 246289 2961 246320
rect 3141 246294 3171 246320
rect 3351 246289 3381 246320
rect 3561 246294 3591 246320
rect 3771 246289 3801 246320
rect 3981 246294 4011 246320
rect 4191 246289 4221 246320
rect 4401 246294 4431 246320
rect 4611 246289 4641 246320
rect 4821 246294 4851 246320
rect 5031 246289 5061 246320
rect 5241 246294 5271 246320
rect 5451 246289 5481 246320
rect 5661 246294 5691 246320
rect 5871 246289 5901 246320
rect 6081 246294 6111 246320
rect 6291 246289 6321 246320
rect 6501 246294 6531 246320
rect 6711 246289 6741 246320
rect 6921 246294 6951 246320
rect 7131 246289 7161 246320
rect 7341 246294 7371 246320
rect 7551 246289 7581 246320
rect 7761 246294 7791 246320
rect 7971 246289 8001 246320
rect 8181 246294 8211 246320
rect 8391 246289 8421 246320
rect 8601 246294 8631 246320
rect 8811 246289 8841 246320
rect 9021 246294 9051 246320
rect 9231 246289 9261 246320
rect 9441 246294 9471 246320
rect 9651 246289 9681 246320
rect 9861 246294 9891 246320
rect 10071 246289 10101 246320
rect 10281 246294 10311 246320
rect 10491 246289 10521 246320
rect 10701 246294 10731 246320
rect 10911 246289 10941 246320
rect 11121 246294 11151 246320
rect 11331 246289 11361 246320
rect 11541 246294 11571 246320
rect 11751 246289 11781 246320
rect 11961 246294 11991 246320
rect 12171 246289 12201 246320
rect 12381 246294 12411 246320
rect 12591 246289 12621 246320
rect 12801 246294 12831 246320
rect 13011 246289 13041 246320
rect 13221 246294 13251 246320
rect 13431 246289 13461 246320
rect 13641 246294 13671 246320
rect 13851 246289 13881 246320
rect 14061 246294 14091 246320
rect 14271 246289 14301 246320
rect 14481 246294 14511 246320
rect 14691 246289 14721 246320
rect 14901 246294 14931 246320
rect 15111 246289 15141 246320
rect 15321 246294 15351 246320
rect 15531 246289 15561 246320
rect 15741 246294 15771 246320
rect 15951 246289 15981 246320
rect 16161 246294 16191 246320
rect 16371 246289 16401 246320
rect 16581 246294 16611 246320
rect 16791 246289 16821 246320
rect 17001 246294 17031 246320
rect 17211 246289 17241 246320
rect 17421 246294 17451 246320
rect 17631 246289 17661 246320
rect 17841 246294 17871 246320
rect 18051 246289 18081 246320
rect 18261 246294 18291 246320
rect 18471 246289 18501 246320
rect 18681 246294 18711 246320
rect 18891 246289 18921 246320
rect 19101 246294 19131 246320
rect 19311 246289 19341 246320
rect 19521 246294 19551 246320
rect 19731 246289 19761 246320
rect 19941 246294 19971 246320
rect 20151 246289 20181 246320
rect 20361 246294 20391 246320
rect 20571 246289 20601 246320
rect 20781 246294 20811 246320
rect 20991 246289 21021 246320
rect 21201 246294 21231 246320
rect 21411 246289 21441 246320
rect 21621 246294 21651 246320
rect 21831 246289 21861 246320
rect 22041 246294 22071 246320
rect 22251 246289 22281 246320
rect 22461 246294 22491 246320
rect 22671 246289 22701 246320
rect 22881 246294 22911 246320
rect 23091 246289 23121 246320
rect 23301 246294 23331 246320
rect 23511 246289 23541 246320
rect 23721 246294 23751 246320
rect 23931 246289 23961 246320
rect 24141 246294 24171 246320
rect 24351 246289 24381 246320
rect 24561 246294 24591 246320
rect 24771 246289 24801 246320
rect 24981 246294 25011 246320
rect 25191 246289 25221 246320
rect 25401 246294 25431 246320
rect 25611 246289 25641 246320
rect 25821 246294 25851 246320
rect 26031 246289 26061 246320
rect 26241 246294 26271 246320
rect 26451 246289 26481 246320
rect 26661 246294 26691 246320
rect 26871 246289 26901 246320
rect 27081 246294 27111 246320
rect 27291 246289 27321 246320
rect -3807 246273 -3741 246289
rect -3807 246131 -3791 246273
rect -3757 246131 -3741 246273
rect -3807 246115 -3741 246131
rect -3387 246273 -3321 246289
rect -3387 246131 -3371 246273
rect -3337 246131 -3321 246273
rect -3387 246115 -3321 246131
rect -2967 246273 -2901 246289
rect -2967 246131 -2951 246273
rect -2917 246131 -2901 246273
rect -2967 246115 -2901 246131
rect -2547 246273 -2481 246289
rect -2547 246131 -2531 246273
rect -2497 246131 -2481 246273
rect -2547 246115 -2481 246131
rect -2127 246273 -2061 246289
rect -2127 246131 -2111 246273
rect -2077 246131 -2061 246273
rect -2127 246115 -2061 246131
rect -1707 246273 -1641 246289
rect -1707 246131 -1691 246273
rect -1657 246131 -1641 246273
rect -1707 246115 -1641 246131
rect -1287 246273 -1221 246289
rect -1287 246131 -1271 246273
rect -1237 246131 -1221 246273
rect -1287 246115 -1221 246131
rect -867 246273 -801 246289
rect -867 246131 -851 246273
rect -817 246131 -801 246273
rect -867 246115 -801 246131
rect -447 246273 -381 246289
rect -447 246131 -431 246273
rect -397 246131 -381 246273
rect -447 246115 -381 246131
rect -27 246273 39 246289
rect -27 246131 -11 246273
rect 23 246131 39 246273
rect -27 246115 39 246131
rect 393 246273 459 246289
rect 393 246131 409 246273
rect 443 246131 459 246273
rect 393 246115 459 246131
rect 813 246273 879 246289
rect 813 246131 829 246273
rect 863 246131 879 246273
rect 813 246115 879 246131
rect 1233 246273 1299 246289
rect 1233 246131 1249 246273
rect 1283 246131 1299 246273
rect 1233 246115 1299 246131
rect 1653 246273 1719 246289
rect 1653 246131 1669 246273
rect 1703 246131 1719 246273
rect 1653 246115 1719 246131
rect 2073 246273 2139 246289
rect 2073 246131 2089 246273
rect 2123 246131 2139 246273
rect 2073 246115 2139 246131
rect 2493 246273 2559 246289
rect 2493 246131 2509 246273
rect 2543 246131 2559 246273
rect 2493 246115 2559 246131
rect 2913 246273 2979 246289
rect 2913 246131 2929 246273
rect 2963 246131 2979 246273
rect 2913 246115 2979 246131
rect 3333 246273 3399 246289
rect 3333 246131 3349 246273
rect 3383 246131 3399 246273
rect 3333 246115 3399 246131
rect 3753 246273 3819 246289
rect 3753 246131 3769 246273
rect 3803 246131 3819 246273
rect 3753 246115 3819 246131
rect 4173 246273 4239 246289
rect 4173 246131 4189 246273
rect 4223 246131 4239 246273
rect 4173 246115 4239 246131
rect 4593 246273 4659 246289
rect 4593 246131 4609 246273
rect 4643 246131 4659 246273
rect 4593 246115 4659 246131
rect 5013 246273 5079 246289
rect 5013 246131 5029 246273
rect 5063 246131 5079 246273
rect 5013 246115 5079 246131
rect 5433 246273 5499 246289
rect 5433 246131 5449 246273
rect 5483 246131 5499 246273
rect 5433 246115 5499 246131
rect 5853 246273 5919 246289
rect 5853 246131 5869 246273
rect 5903 246131 5919 246273
rect 5853 246115 5919 246131
rect 6273 246273 6339 246289
rect 6273 246131 6289 246273
rect 6323 246131 6339 246273
rect 6273 246115 6339 246131
rect 6693 246273 6759 246289
rect 6693 246131 6709 246273
rect 6743 246131 6759 246273
rect 6693 246115 6759 246131
rect 7113 246273 7179 246289
rect 7113 246131 7129 246273
rect 7163 246131 7179 246273
rect 7113 246115 7179 246131
rect 7533 246273 7599 246289
rect 7533 246131 7549 246273
rect 7583 246131 7599 246273
rect 7533 246115 7599 246131
rect 7953 246273 8019 246289
rect 7953 246131 7969 246273
rect 8003 246131 8019 246273
rect 7953 246115 8019 246131
rect 8373 246273 8439 246289
rect 8373 246131 8389 246273
rect 8423 246131 8439 246273
rect 8373 246115 8439 246131
rect 8793 246273 8859 246289
rect 8793 246131 8809 246273
rect 8843 246131 8859 246273
rect 8793 246115 8859 246131
rect 9213 246273 9279 246289
rect 9213 246131 9229 246273
rect 9263 246131 9279 246273
rect 9213 246115 9279 246131
rect 9633 246273 9699 246289
rect 9633 246131 9649 246273
rect 9683 246131 9699 246273
rect 9633 246115 9699 246131
rect 10053 246273 10119 246289
rect 10053 246131 10069 246273
rect 10103 246131 10119 246273
rect 10053 246115 10119 246131
rect 10473 246273 10539 246289
rect 10473 246131 10489 246273
rect 10523 246131 10539 246273
rect 10473 246115 10539 246131
rect 10893 246273 10959 246289
rect 10893 246131 10909 246273
rect 10943 246131 10959 246273
rect 10893 246115 10959 246131
rect 11313 246273 11379 246289
rect 11313 246131 11329 246273
rect 11363 246131 11379 246273
rect 11313 246115 11379 246131
rect 11733 246273 11799 246289
rect 11733 246131 11749 246273
rect 11783 246131 11799 246273
rect 11733 246115 11799 246131
rect 12153 246273 12219 246289
rect 12153 246131 12169 246273
rect 12203 246131 12219 246273
rect 12153 246115 12219 246131
rect 12573 246273 12639 246289
rect 12573 246131 12589 246273
rect 12623 246131 12639 246273
rect 12573 246115 12639 246131
rect 12993 246273 13059 246289
rect 12993 246131 13009 246273
rect 13043 246131 13059 246273
rect 12993 246115 13059 246131
rect 13413 246273 13479 246289
rect 13413 246131 13429 246273
rect 13463 246131 13479 246273
rect 13413 246115 13479 246131
rect 13833 246273 13899 246289
rect 13833 246131 13849 246273
rect 13883 246131 13899 246273
rect 13833 246115 13899 246131
rect 14253 246273 14319 246289
rect 14253 246131 14269 246273
rect 14303 246131 14319 246273
rect 14253 246115 14319 246131
rect 14673 246273 14739 246289
rect 14673 246131 14689 246273
rect 14723 246131 14739 246273
rect 14673 246115 14739 246131
rect 15093 246273 15159 246289
rect 15093 246131 15109 246273
rect 15143 246131 15159 246273
rect 15093 246115 15159 246131
rect 15513 246273 15579 246289
rect 15513 246131 15529 246273
rect 15563 246131 15579 246273
rect 15513 246115 15579 246131
rect 15933 246273 15999 246289
rect 15933 246131 15949 246273
rect 15983 246131 15999 246273
rect 15933 246115 15999 246131
rect 16353 246273 16419 246289
rect 16353 246131 16369 246273
rect 16403 246131 16419 246273
rect 16353 246115 16419 246131
rect 16773 246273 16839 246289
rect 16773 246131 16789 246273
rect 16823 246131 16839 246273
rect 16773 246115 16839 246131
rect 17193 246273 17259 246289
rect 17193 246131 17209 246273
rect 17243 246131 17259 246273
rect 17193 246115 17259 246131
rect 17613 246273 17679 246289
rect 17613 246131 17629 246273
rect 17663 246131 17679 246273
rect 17613 246115 17679 246131
rect 18033 246273 18099 246289
rect 18033 246131 18049 246273
rect 18083 246131 18099 246273
rect 18033 246115 18099 246131
rect 18453 246273 18519 246289
rect 18453 246131 18469 246273
rect 18503 246131 18519 246273
rect 18453 246115 18519 246131
rect 18873 246273 18939 246289
rect 18873 246131 18889 246273
rect 18923 246131 18939 246273
rect 18873 246115 18939 246131
rect 19293 246273 19359 246289
rect 19293 246131 19309 246273
rect 19343 246131 19359 246273
rect 19293 246115 19359 246131
rect 19713 246273 19779 246289
rect 19713 246131 19729 246273
rect 19763 246131 19779 246273
rect 19713 246115 19779 246131
rect 20133 246273 20199 246289
rect 20133 246131 20149 246273
rect 20183 246131 20199 246273
rect 20133 246115 20199 246131
rect 20553 246273 20619 246289
rect 20553 246131 20569 246273
rect 20603 246131 20619 246273
rect 20553 246115 20619 246131
rect 20973 246273 21039 246289
rect 20973 246131 20989 246273
rect 21023 246131 21039 246273
rect 20973 246115 21039 246131
rect 21393 246273 21459 246289
rect 21393 246131 21409 246273
rect 21443 246131 21459 246273
rect 21393 246115 21459 246131
rect 21813 246273 21879 246289
rect 21813 246131 21829 246273
rect 21863 246131 21879 246273
rect 21813 246115 21879 246131
rect 22233 246273 22299 246289
rect 22233 246131 22249 246273
rect 22283 246131 22299 246273
rect 22233 246115 22299 246131
rect 22653 246273 22719 246289
rect 22653 246131 22669 246273
rect 22703 246131 22719 246273
rect 22653 246115 22719 246131
rect 23073 246273 23139 246289
rect 23073 246131 23089 246273
rect 23123 246131 23139 246273
rect 23073 246115 23139 246131
rect 23493 246273 23559 246289
rect 23493 246131 23509 246273
rect 23543 246131 23559 246273
rect 23493 246115 23559 246131
rect 23913 246273 23979 246289
rect 23913 246131 23929 246273
rect 23963 246131 23979 246273
rect 23913 246115 23979 246131
rect 24333 246273 24399 246289
rect 24333 246131 24349 246273
rect 24383 246131 24399 246273
rect 24333 246115 24399 246131
rect 24753 246273 24819 246289
rect 24753 246131 24769 246273
rect 24803 246131 24819 246273
rect 24753 246115 24819 246131
rect 25173 246273 25239 246289
rect 25173 246131 25189 246273
rect 25223 246131 25239 246273
rect 25173 246115 25239 246131
rect 25593 246273 25659 246289
rect 25593 246131 25609 246273
rect 25643 246131 25659 246273
rect 25593 246115 25659 246131
rect 26013 246273 26079 246289
rect 26013 246131 26029 246273
rect 26063 246131 26079 246273
rect 26013 246115 26079 246131
rect 26433 246273 26499 246289
rect 26433 246131 26449 246273
rect 26483 246131 26499 246273
rect 26433 246115 26499 246131
rect 26853 246273 26919 246289
rect 26853 246131 26869 246273
rect 26903 246131 26919 246273
rect 26853 246115 26919 246131
rect 27273 246273 27339 246289
rect 27273 246131 27289 246273
rect 27323 246131 27339 246273
rect 27273 246115 27339 246131
rect -3999 246084 -3969 246110
rect -3789 246084 -3759 246115
rect -3579 246084 -3549 246110
rect -3369 246084 -3339 246115
rect -3159 246084 -3129 246110
rect -2949 246084 -2919 246115
rect -2739 246084 -2709 246110
rect -2529 246084 -2499 246115
rect -2319 246084 -2289 246110
rect -2109 246084 -2079 246115
rect -1899 246084 -1869 246110
rect -1689 246084 -1659 246115
rect -1479 246084 -1449 246110
rect -1269 246084 -1239 246115
rect -1059 246084 -1029 246110
rect -849 246084 -819 246115
rect -639 246084 -609 246110
rect -429 246084 -399 246115
rect -219 246084 -189 246110
rect -9 246084 21 246115
rect 201 246084 231 246110
rect 411 246084 441 246115
rect 621 246084 651 246110
rect 831 246084 861 246115
rect 1041 246084 1071 246110
rect 1251 246084 1281 246115
rect 1461 246084 1491 246110
rect 1671 246084 1701 246115
rect 1881 246084 1911 246110
rect 2091 246084 2121 246115
rect 2301 246084 2331 246110
rect 2511 246084 2541 246115
rect 2721 246084 2751 246110
rect 2931 246084 2961 246115
rect 3141 246084 3171 246110
rect 3351 246084 3381 246115
rect 3561 246084 3591 246110
rect 3771 246084 3801 246115
rect 3981 246084 4011 246110
rect 4191 246084 4221 246115
rect 4401 246084 4431 246110
rect 4611 246084 4641 246115
rect 4821 246084 4851 246110
rect 5031 246084 5061 246115
rect 5241 246084 5271 246110
rect 5451 246084 5481 246115
rect 5661 246084 5691 246110
rect 5871 246084 5901 246115
rect 6081 246084 6111 246110
rect 6291 246084 6321 246115
rect 6501 246084 6531 246110
rect 6711 246084 6741 246115
rect 6921 246084 6951 246110
rect 7131 246084 7161 246115
rect 7341 246084 7371 246110
rect 7551 246084 7581 246115
rect 7761 246084 7791 246110
rect 7971 246084 8001 246115
rect 8181 246084 8211 246110
rect 8391 246084 8421 246115
rect 8601 246084 8631 246110
rect 8811 246084 8841 246115
rect 9021 246084 9051 246110
rect 9231 246084 9261 246115
rect 9441 246084 9471 246110
rect 9651 246084 9681 246115
rect 9861 246084 9891 246110
rect 10071 246084 10101 246115
rect 10281 246084 10311 246110
rect 10491 246084 10521 246115
rect 10701 246084 10731 246110
rect 10911 246084 10941 246115
rect 11121 246084 11151 246110
rect 11331 246084 11361 246115
rect 11541 246084 11571 246110
rect 11751 246084 11781 246115
rect 11961 246084 11991 246110
rect 12171 246084 12201 246115
rect 12381 246084 12411 246110
rect 12591 246084 12621 246115
rect 12801 246084 12831 246110
rect 13011 246084 13041 246115
rect 13221 246084 13251 246110
rect 13431 246084 13461 246115
rect 13641 246084 13671 246110
rect 13851 246084 13881 246115
rect 14061 246084 14091 246110
rect 14271 246084 14301 246115
rect 14481 246084 14511 246110
rect 14691 246084 14721 246115
rect 14901 246084 14931 246110
rect 15111 246084 15141 246115
rect 15321 246084 15351 246110
rect 15531 246084 15561 246115
rect 15741 246084 15771 246110
rect 15951 246084 15981 246115
rect 16161 246084 16191 246110
rect 16371 246084 16401 246115
rect 16581 246084 16611 246110
rect 16791 246084 16821 246115
rect 17001 246084 17031 246110
rect 17211 246084 17241 246115
rect 17421 246084 17451 246110
rect 17631 246084 17661 246115
rect 17841 246084 17871 246110
rect 18051 246084 18081 246115
rect 18261 246084 18291 246110
rect 18471 246084 18501 246115
rect 18681 246084 18711 246110
rect 18891 246084 18921 246115
rect 19101 246084 19131 246110
rect 19311 246084 19341 246115
rect 19521 246084 19551 246110
rect 19731 246084 19761 246115
rect 19941 246084 19971 246110
rect 20151 246084 20181 246115
rect 20361 246084 20391 246110
rect 20571 246084 20601 246115
rect 20781 246084 20811 246110
rect 20991 246084 21021 246115
rect 21201 246084 21231 246110
rect 21411 246084 21441 246115
rect 21621 246084 21651 246110
rect 21831 246084 21861 246115
rect 22041 246084 22071 246110
rect 22251 246084 22281 246115
rect 22461 246084 22491 246110
rect 22671 246084 22701 246115
rect 22881 246084 22911 246110
rect 23091 246084 23121 246115
rect 23301 246084 23331 246110
rect 23511 246084 23541 246115
rect 23721 246084 23751 246110
rect 23931 246084 23961 246115
rect 24141 246084 24171 246110
rect 24351 246084 24381 246115
rect 24561 246084 24591 246110
rect 24771 246084 24801 246115
rect 24981 246084 25011 246110
rect 25191 246084 25221 246115
rect 25401 246084 25431 246110
rect 25611 246084 25641 246115
rect 25821 246084 25851 246110
rect 26031 246084 26061 246115
rect 26241 246084 26271 246110
rect 26451 246084 26481 246115
rect 26661 246084 26691 246110
rect 26871 246084 26901 246115
rect 27081 246084 27111 246110
rect 27291 246084 27321 246115
rect -3999 245253 -3969 245284
rect -3789 245258 -3759 245284
rect -3579 245253 -3549 245284
rect -3369 245258 -3339 245284
rect -3159 245253 -3129 245284
rect -2949 245258 -2919 245284
rect -2739 245253 -2709 245284
rect -2529 245258 -2499 245284
rect -2319 245253 -2289 245284
rect -2109 245258 -2079 245284
rect -1899 245253 -1869 245284
rect -1689 245258 -1659 245284
rect -1479 245253 -1449 245284
rect -1269 245258 -1239 245284
rect -1059 245253 -1029 245284
rect -849 245258 -819 245284
rect -639 245253 -609 245284
rect -429 245258 -399 245284
rect -219 245253 -189 245284
rect -9 245258 21 245284
rect 201 245253 231 245284
rect 411 245258 441 245284
rect 621 245253 651 245284
rect 831 245258 861 245284
rect 1041 245253 1071 245284
rect 1251 245258 1281 245284
rect 1461 245253 1491 245284
rect 1671 245258 1701 245284
rect 1881 245253 1911 245284
rect 2091 245258 2121 245284
rect 2301 245253 2331 245284
rect 2511 245258 2541 245284
rect 2721 245253 2751 245284
rect 2931 245258 2961 245284
rect 3141 245253 3171 245284
rect 3351 245258 3381 245284
rect 3561 245253 3591 245284
rect 3771 245258 3801 245284
rect 3981 245253 4011 245284
rect 4191 245258 4221 245284
rect 4401 245253 4431 245284
rect 4611 245258 4641 245284
rect 4821 245253 4851 245284
rect 5031 245258 5061 245284
rect 5241 245253 5271 245284
rect 5451 245258 5481 245284
rect 5661 245253 5691 245284
rect 5871 245258 5901 245284
rect 6081 245253 6111 245284
rect 6291 245258 6321 245284
rect 6501 245253 6531 245284
rect 6711 245258 6741 245284
rect 6921 245253 6951 245284
rect 7131 245258 7161 245284
rect 7341 245253 7371 245284
rect 7551 245258 7581 245284
rect 7761 245253 7791 245284
rect 7971 245258 8001 245284
rect 8181 245253 8211 245284
rect 8391 245258 8421 245284
rect 8601 245253 8631 245284
rect 8811 245258 8841 245284
rect 9021 245253 9051 245284
rect 9231 245258 9261 245284
rect 9441 245253 9471 245284
rect 9651 245258 9681 245284
rect 9861 245253 9891 245284
rect 10071 245258 10101 245284
rect 10281 245253 10311 245284
rect 10491 245258 10521 245284
rect 10701 245253 10731 245284
rect 10911 245258 10941 245284
rect 11121 245253 11151 245284
rect 11331 245258 11361 245284
rect 11541 245253 11571 245284
rect 11751 245258 11781 245284
rect 11961 245253 11991 245284
rect 12171 245258 12201 245284
rect 12381 245253 12411 245284
rect 12591 245258 12621 245284
rect 12801 245253 12831 245284
rect 13011 245258 13041 245284
rect 13221 245253 13251 245284
rect 13431 245258 13461 245284
rect 13641 245253 13671 245284
rect 13851 245258 13881 245284
rect 14061 245253 14091 245284
rect 14271 245258 14301 245284
rect 14481 245253 14511 245284
rect 14691 245258 14721 245284
rect 14901 245253 14931 245284
rect 15111 245258 15141 245284
rect 15321 245253 15351 245284
rect 15531 245258 15561 245284
rect 15741 245253 15771 245284
rect 15951 245258 15981 245284
rect 16161 245253 16191 245284
rect 16371 245258 16401 245284
rect 16581 245253 16611 245284
rect 16791 245258 16821 245284
rect 17001 245253 17031 245284
rect 17211 245258 17241 245284
rect 17421 245253 17451 245284
rect 17631 245258 17661 245284
rect 17841 245253 17871 245284
rect 18051 245258 18081 245284
rect 18261 245253 18291 245284
rect 18471 245258 18501 245284
rect 18681 245253 18711 245284
rect 18891 245258 18921 245284
rect 19101 245253 19131 245284
rect 19311 245258 19341 245284
rect 19521 245253 19551 245284
rect 19731 245258 19761 245284
rect 19941 245253 19971 245284
rect 20151 245258 20181 245284
rect 20361 245253 20391 245284
rect 20571 245258 20601 245284
rect 20781 245253 20811 245284
rect 20991 245258 21021 245284
rect 21201 245253 21231 245284
rect 21411 245258 21441 245284
rect 21621 245253 21651 245284
rect 21831 245258 21861 245284
rect 22041 245253 22071 245284
rect 22251 245258 22281 245284
rect 22461 245253 22491 245284
rect 22671 245258 22701 245284
rect 22881 245253 22911 245284
rect 23091 245258 23121 245284
rect 23301 245253 23331 245284
rect 23511 245258 23541 245284
rect 23721 245253 23751 245284
rect 23931 245258 23961 245284
rect 24141 245253 24171 245284
rect 24351 245258 24381 245284
rect 24561 245253 24591 245284
rect 24771 245258 24801 245284
rect 24981 245253 25011 245284
rect 25191 245258 25221 245284
rect 25401 245253 25431 245284
rect 25611 245258 25641 245284
rect 25821 245253 25851 245284
rect 26031 245258 26061 245284
rect 26241 245253 26271 245284
rect 26451 245258 26481 245284
rect 26661 245253 26691 245284
rect 26871 245258 26901 245284
rect 27081 245253 27111 245284
rect 27291 245258 27321 245284
rect -4017 245237 -3951 245253
rect -4017 245095 -4001 245237
rect -3967 245095 -3951 245237
rect -4017 245079 -3951 245095
rect -3597 245237 -3531 245253
rect -3597 245095 -3581 245237
rect -3547 245095 -3531 245237
rect -3597 245079 -3531 245095
rect -3177 245237 -3111 245253
rect -3177 245095 -3161 245237
rect -3127 245095 -3111 245237
rect -3177 245079 -3111 245095
rect -2757 245237 -2691 245253
rect -2757 245095 -2741 245237
rect -2707 245095 -2691 245237
rect -2757 245079 -2691 245095
rect -2337 245237 -2271 245253
rect -2337 245095 -2321 245237
rect -2287 245095 -2271 245237
rect -2337 245079 -2271 245095
rect -1917 245237 -1851 245253
rect -1917 245095 -1901 245237
rect -1867 245095 -1851 245237
rect -1917 245079 -1851 245095
rect -1497 245237 -1431 245253
rect -1497 245095 -1481 245237
rect -1447 245095 -1431 245237
rect -1497 245079 -1431 245095
rect -1077 245237 -1011 245253
rect -1077 245095 -1061 245237
rect -1027 245095 -1011 245237
rect -1077 245079 -1011 245095
rect -657 245237 -591 245253
rect -657 245095 -641 245237
rect -607 245095 -591 245237
rect -657 245079 -591 245095
rect -237 245237 -171 245253
rect -237 245095 -221 245237
rect -187 245095 -171 245237
rect -237 245079 -171 245095
rect 183 245237 249 245253
rect 183 245095 199 245237
rect 233 245095 249 245237
rect 183 245079 249 245095
rect 603 245237 669 245253
rect 603 245095 619 245237
rect 653 245095 669 245237
rect 603 245079 669 245095
rect 1023 245237 1089 245253
rect 1023 245095 1039 245237
rect 1073 245095 1089 245237
rect 1023 245079 1089 245095
rect 1443 245237 1509 245253
rect 1443 245095 1459 245237
rect 1493 245095 1509 245237
rect 1443 245079 1509 245095
rect 1863 245237 1929 245253
rect 1863 245095 1879 245237
rect 1913 245095 1929 245237
rect 1863 245079 1929 245095
rect 2283 245237 2349 245253
rect 2283 245095 2299 245237
rect 2333 245095 2349 245237
rect 2283 245079 2349 245095
rect 2703 245237 2769 245253
rect 2703 245095 2719 245237
rect 2753 245095 2769 245237
rect 2703 245079 2769 245095
rect 3123 245237 3189 245253
rect 3123 245095 3139 245237
rect 3173 245095 3189 245237
rect 3123 245079 3189 245095
rect 3543 245237 3609 245253
rect 3543 245095 3559 245237
rect 3593 245095 3609 245237
rect 3543 245079 3609 245095
rect 3963 245237 4029 245253
rect 3963 245095 3979 245237
rect 4013 245095 4029 245237
rect 3963 245079 4029 245095
rect 4383 245237 4449 245253
rect 4383 245095 4399 245237
rect 4433 245095 4449 245237
rect 4383 245079 4449 245095
rect 4803 245237 4869 245253
rect 4803 245095 4819 245237
rect 4853 245095 4869 245237
rect 4803 245079 4869 245095
rect 5223 245237 5289 245253
rect 5223 245095 5239 245237
rect 5273 245095 5289 245237
rect 5223 245079 5289 245095
rect 5643 245237 5709 245253
rect 5643 245095 5659 245237
rect 5693 245095 5709 245237
rect 5643 245079 5709 245095
rect 6063 245237 6129 245253
rect 6063 245095 6079 245237
rect 6113 245095 6129 245237
rect 6063 245079 6129 245095
rect 6483 245237 6549 245253
rect 6483 245095 6499 245237
rect 6533 245095 6549 245237
rect 6483 245079 6549 245095
rect 6903 245237 6969 245253
rect 6903 245095 6919 245237
rect 6953 245095 6969 245237
rect 6903 245079 6969 245095
rect 7323 245237 7389 245253
rect 7323 245095 7339 245237
rect 7373 245095 7389 245237
rect 7323 245079 7389 245095
rect 7743 245237 7809 245253
rect 7743 245095 7759 245237
rect 7793 245095 7809 245237
rect 7743 245079 7809 245095
rect 8163 245237 8229 245253
rect 8163 245095 8179 245237
rect 8213 245095 8229 245237
rect 8163 245079 8229 245095
rect 8583 245237 8649 245253
rect 8583 245095 8599 245237
rect 8633 245095 8649 245237
rect 8583 245079 8649 245095
rect 9003 245237 9069 245253
rect 9003 245095 9019 245237
rect 9053 245095 9069 245237
rect 9003 245079 9069 245095
rect 9423 245237 9489 245253
rect 9423 245095 9439 245237
rect 9473 245095 9489 245237
rect 9423 245079 9489 245095
rect 9843 245237 9909 245253
rect 9843 245095 9859 245237
rect 9893 245095 9909 245237
rect 9843 245079 9909 245095
rect 10263 245237 10329 245253
rect 10263 245095 10279 245237
rect 10313 245095 10329 245237
rect 10263 245079 10329 245095
rect 10683 245237 10749 245253
rect 10683 245095 10699 245237
rect 10733 245095 10749 245237
rect 10683 245079 10749 245095
rect 11103 245237 11169 245253
rect 11103 245095 11119 245237
rect 11153 245095 11169 245237
rect 11103 245079 11169 245095
rect 11523 245237 11589 245253
rect 11523 245095 11539 245237
rect 11573 245095 11589 245237
rect 11523 245079 11589 245095
rect 11943 245237 12009 245253
rect 11943 245095 11959 245237
rect 11993 245095 12009 245237
rect 11943 245079 12009 245095
rect 12363 245237 12429 245253
rect 12363 245095 12379 245237
rect 12413 245095 12429 245237
rect 12363 245079 12429 245095
rect 12783 245237 12849 245253
rect 12783 245095 12799 245237
rect 12833 245095 12849 245237
rect 12783 245079 12849 245095
rect 13203 245237 13269 245253
rect 13203 245095 13219 245237
rect 13253 245095 13269 245237
rect 13203 245079 13269 245095
rect 13623 245237 13689 245253
rect 13623 245095 13639 245237
rect 13673 245095 13689 245237
rect 13623 245079 13689 245095
rect 14043 245237 14109 245253
rect 14043 245095 14059 245237
rect 14093 245095 14109 245237
rect 14043 245079 14109 245095
rect 14463 245237 14529 245253
rect 14463 245095 14479 245237
rect 14513 245095 14529 245237
rect 14463 245079 14529 245095
rect 14883 245237 14949 245253
rect 14883 245095 14899 245237
rect 14933 245095 14949 245237
rect 14883 245079 14949 245095
rect 15303 245237 15369 245253
rect 15303 245095 15319 245237
rect 15353 245095 15369 245237
rect 15303 245079 15369 245095
rect 15723 245237 15789 245253
rect 15723 245095 15739 245237
rect 15773 245095 15789 245237
rect 15723 245079 15789 245095
rect 16143 245237 16209 245253
rect 16143 245095 16159 245237
rect 16193 245095 16209 245237
rect 16143 245079 16209 245095
rect 16563 245237 16629 245253
rect 16563 245095 16579 245237
rect 16613 245095 16629 245237
rect 16563 245079 16629 245095
rect 16983 245237 17049 245253
rect 16983 245095 16999 245237
rect 17033 245095 17049 245237
rect 16983 245079 17049 245095
rect 17403 245237 17469 245253
rect 17403 245095 17419 245237
rect 17453 245095 17469 245237
rect 17403 245079 17469 245095
rect 17823 245237 17889 245253
rect 17823 245095 17839 245237
rect 17873 245095 17889 245237
rect 17823 245079 17889 245095
rect 18243 245237 18309 245253
rect 18243 245095 18259 245237
rect 18293 245095 18309 245237
rect 18243 245079 18309 245095
rect 18663 245237 18729 245253
rect 18663 245095 18679 245237
rect 18713 245095 18729 245237
rect 18663 245079 18729 245095
rect 19083 245237 19149 245253
rect 19083 245095 19099 245237
rect 19133 245095 19149 245237
rect 19083 245079 19149 245095
rect 19503 245237 19569 245253
rect 19503 245095 19519 245237
rect 19553 245095 19569 245237
rect 19503 245079 19569 245095
rect 19923 245237 19989 245253
rect 19923 245095 19939 245237
rect 19973 245095 19989 245237
rect 19923 245079 19989 245095
rect 20343 245237 20409 245253
rect 20343 245095 20359 245237
rect 20393 245095 20409 245237
rect 20343 245079 20409 245095
rect 20763 245237 20829 245253
rect 20763 245095 20779 245237
rect 20813 245095 20829 245237
rect 20763 245079 20829 245095
rect 21183 245237 21249 245253
rect 21183 245095 21199 245237
rect 21233 245095 21249 245237
rect 21183 245079 21249 245095
rect 21603 245237 21669 245253
rect 21603 245095 21619 245237
rect 21653 245095 21669 245237
rect 21603 245079 21669 245095
rect 22023 245237 22089 245253
rect 22023 245095 22039 245237
rect 22073 245095 22089 245237
rect 22023 245079 22089 245095
rect 22443 245237 22509 245253
rect 22443 245095 22459 245237
rect 22493 245095 22509 245237
rect 22443 245079 22509 245095
rect 22863 245237 22929 245253
rect 22863 245095 22879 245237
rect 22913 245095 22929 245237
rect 22863 245079 22929 245095
rect 23283 245237 23349 245253
rect 23283 245095 23299 245237
rect 23333 245095 23349 245237
rect 23283 245079 23349 245095
rect 23703 245237 23769 245253
rect 23703 245095 23719 245237
rect 23753 245095 23769 245237
rect 23703 245079 23769 245095
rect 24123 245237 24189 245253
rect 24123 245095 24139 245237
rect 24173 245095 24189 245237
rect 24123 245079 24189 245095
rect 24543 245237 24609 245253
rect 24543 245095 24559 245237
rect 24593 245095 24609 245237
rect 24543 245079 24609 245095
rect 24963 245237 25029 245253
rect 24963 245095 24979 245237
rect 25013 245095 25029 245237
rect 24963 245079 25029 245095
rect 25383 245237 25449 245253
rect 25383 245095 25399 245237
rect 25433 245095 25449 245237
rect 25383 245079 25449 245095
rect 25803 245237 25869 245253
rect 25803 245095 25819 245237
rect 25853 245095 25869 245237
rect 25803 245079 25869 245095
rect 26223 245237 26289 245253
rect 26223 245095 26239 245237
rect 26273 245095 26289 245237
rect 26223 245079 26289 245095
rect 26643 245237 26709 245253
rect 26643 245095 26659 245237
rect 26693 245095 26709 245237
rect 26643 245079 26709 245095
rect 27063 245237 27129 245253
rect 27063 245095 27079 245237
rect 27113 245095 27129 245237
rect 27063 245079 27129 245095
rect -3999 245048 -3969 245079
rect -3789 245048 -3759 245074
rect -3579 245048 -3549 245079
rect -3369 245048 -3339 245074
rect -3159 245048 -3129 245079
rect -2949 245048 -2919 245074
rect -2739 245048 -2709 245079
rect -2529 245048 -2499 245074
rect -2319 245048 -2289 245079
rect -2109 245048 -2079 245074
rect -1899 245048 -1869 245079
rect -1689 245048 -1659 245074
rect -1479 245048 -1449 245079
rect -1269 245048 -1239 245074
rect -1059 245048 -1029 245079
rect -849 245048 -819 245074
rect -639 245048 -609 245079
rect -429 245048 -399 245074
rect -219 245048 -189 245079
rect -9 245048 21 245074
rect 201 245048 231 245079
rect 411 245048 441 245074
rect 621 245048 651 245079
rect 831 245048 861 245074
rect 1041 245048 1071 245079
rect 1251 245048 1281 245074
rect 1461 245048 1491 245079
rect 1671 245048 1701 245074
rect 1881 245048 1911 245079
rect 2091 245048 2121 245074
rect 2301 245048 2331 245079
rect 2511 245048 2541 245074
rect 2721 245048 2751 245079
rect 2931 245048 2961 245074
rect 3141 245048 3171 245079
rect 3351 245048 3381 245074
rect 3561 245048 3591 245079
rect 3771 245048 3801 245074
rect 3981 245048 4011 245079
rect 4191 245048 4221 245074
rect 4401 245048 4431 245079
rect 4611 245048 4641 245074
rect 4821 245048 4851 245079
rect 5031 245048 5061 245074
rect 5241 245048 5271 245079
rect 5451 245048 5481 245074
rect 5661 245048 5691 245079
rect 5871 245048 5901 245074
rect 6081 245048 6111 245079
rect 6291 245048 6321 245074
rect 6501 245048 6531 245079
rect 6711 245048 6741 245074
rect 6921 245048 6951 245079
rect 7131 245048 7161 245074
rect 7341 245048 7371 245079
rect 7551 245048 7581 245074
rect 7761 245048 7791 245079
rect 7971 245048 8001 245074
rect 8181 245048 8211 245079
rect 8391 245048 8421 245074
rect 8601 245048 8631 245079
rect 8811 245048 8841 245074
rect 9021 245048 9051 245079
rect 9231 245048 9261 245074
rect 9441 245048 9471 245079
rect 9651 245048 9681 245074
rect 9861 245048 9891 245079
rect 10071 245048 10101 245074
rect 10281 245048 10311 245079
rect 10491 245048 10521 245074
rect 10701 245048 10731 245079
rect 10911 245048 10941 245074
rect 11121 245048 11151 245079
rect 11331 245048 11361 245074
rect 11541 245048 11571 245079
rect 11751 245048 11781 245074
rect 11961 245048 11991 245079
rect 12171 245048 12201 245074
rect 12381 245048 12411 245079
rect 12591 245048 12621 245074
rect 12801 245048 12831 245079
rect 13011 245048 13041 245074
rect 13221 245048 13251 245079
rect 13431 245048 13461 245074
rect 13641 245048 13671 245079
rect 13851 245048 13881 245074
rect 14061 245048 14091 245079
rect 14271 245048 14301 245074
rect 14481 245048 14511 245079
rect 14691 245048 14721 245074
rect 14901 245048 14931 245079
rect 15111 245048 15141 245074
rect 15321 245048 15351 245079
rect 15531 245048 15561 245074
rect 15741 245048 15771 245079
rect 15951 245048 15981 245074
rect 16161 245048 16191 245079
rect 16371 245048 16401 245074
rect 16581 245048 16611 245079
rect 16791 245048 16821 245074
rect 17001 245048 17031 245079
rect 17211 245048 17241 245074
rect 17421 245048 17451 245079
rect 17631 245048 17661 245074
rect 17841 245048 17871 245079
rect 18051 245048 18081 245074
rect 18261 245048 18291 245079
rect 18471 245048 18501 245074
rect 18681 245048 18711 245079
rect 18891 245048 18921 245074
rect 19101 245048 19131 245079
rect 19311 245048 19341 245074
rect 19521 245048 19551 245079
rect 19731 245048 19761 245074
rect 19941 245048 19971 245079
rect 20151 245048 20181 245074
rect 20361 245048 20391 245079
rect 20571 245048 20601 245074
rect 20781 245048 20811 245079
rect 20991 245048 21021 245074
rect 21201 245048 21231 245079
rect 21411 245048 21441 245074
rect 21621 245048 21651 245079
rect 21831 245048 21861 245074
rect 22041 245048 22071 245079
rect 22251 245048 22281 245074
rect 22461 245048 22491 245079
rect 22671 245048 22701 245074
rect 22881 245048 22911 245079
rect 23091 245048 23121 245074
rect 23301 245048 23331 245079
rect 23511 245048 23541 245074
rect 23721 245048 23751 245079
rect 23931 245048 23961 245074
rect 24141 245048 24171 245079
rect 24351 245048 24381 245074
rect 24561 245048 24591 245079
rect 24771 245048 24801 245074
rect 24981 245048 25011 245079
rect 25191 245048 25221 245074
rect 25401 245048 25431 245079
rect 25611 245048 25641 245074
rect 25821 245048 25851 245079
rect 26031 245048 26061 245074
rect 26241 245048 26271 245079
rect 26451 245048 26481 245074
rect 26661 245048 26691 245079
rect 26871 245048 26901 245074
rect 27081 245048 27111 245079
rect 27291 245048 27321 245074
rect -3999 244222 -3969 244248
rect -3789 244217 -3759 244248
rect -3579 244222 -3549 244248
rect -3369 244217 -3339 244248
rect -3159 244222 -3129 244248
rect -2949 244217 -2919 244248
rect -2739 244222 -2709 244248
rect -2529 244217 -2499 244248
rect -2319 244222 -2289 244248
rect -2109 244217 -2079 244248
rect -1899 244222 -1869 244248
rect -1689 244217 -1659 244248
rect -1479 244222 -1449 244248
rect -1269 244217 -1239 244248
rect -1059 244222 -1029 244248
rect -849 244217 -819 244248
rect -639 244222 -609 244248
rect -429 244217 -399 244248
rect -219 244222 -189 244248
rect -9 244217 21 244248
rect 201 244222 231 244248
rect 411 244217 441 244248
rect 621 244222 651 244248
rect 831 244217 861 244248
rect 1041 244222 1071 244248
rect 1251 244217 1281 244248
rect 1461 244222 1491 244248
rect 1671 244217 1701 244248
rect 1881 244222 1911 244248
rect 2091 244217 2121 244248
rect 2301 244222 2331 244248
rect 2511 244217 2541 244248
rect 2721 244222 2751 244248
rect 2931 244217 2961 244248
rect 3141 244222 3171 244248
rect 3351 244217 3381 244248
rect 3561 244222 3591 244248
rect 3771 244217 3801 244248
rect 3981 244222 4011 244248
rect 4191 244217 4221 244248
rect 4401 244222 4431 244248
rect 4611 244217 4641 244248
rect 4821 244222 4851 244248
rect 5031 244217 5061 244248
rect 5241 244222 5271 244248
rect 5451 244217 5481 244248
rect 5661 244222 5691 244248
rect 5871 244217 5901 244248
rect 6081 244222 6111 244248
rect 6291 244217 6321 244248
rect 6501 244222 6531 244248
rect 6711 244217 6741 244248
rect 6921 244222 6951 244248
rect 7131 244217 7161 244248
rect 7341 244222 7371 244248
rect 7551 244217 7581 244248
rect 7761 244222 7791 244248
rect 7971 244217 8001 244248
rect 8181 244222 8211 244248
rect 8391 244217 8421 244248
rect 8601 244222 8631 244248
rect 8811 244217 8841 244248
rect 9021 244222 9051 244248
rect 9231 244217 9261 244248
rect 9441 244222 9471 244248
rect 9651 244217 9681 244248
rect 9861 244222 9891 244248
rect 10071 244217 10101 244248
rect 10281 244222 10311 244248
rect 10491 244217 10521 244248
rect 10701 244222 10731 244248
rect 10911 244217 10941 244248
rect 11121 244222 11151 244248
rect 11331 244217 11361 244248
rect 11541 244222 11571 244248
rect 11751 244217 11781 244248
rect 11961 244222 11991 244248
rect 12171 244217 12201 244248
rect 12381 244222 12411 244248
rect 12591 244217 12621 244248
rect 12801 244222 12831 244248
rect 13011 244217 13041 244248
rect 13221 244222 13251 244248
rect 13431 244217 13461 244248
rect 13641 244222 13671 244248
rect 13851 244217 13881 244248
rect 14061 244222 14091 244248
rect 14271 244217 14301 244248
rect 14481 244222 14511 244248
rect 14691 244217 14721 244248
rect 14901 244222 14931 244248
rect 15111 244217 15141 244248
rect 15321 244222 15351 244248
rect 15531 244217 15561 244248
rect 15741 244222 15771 244248
rect 15951 244217 15981 244248
rect 16161 244222 16191 244248
rect 16371 244217 16401 244248
rect 16581 244222 16611 244248
rect 16791 244217 16821 244248
rect 17001 244222 17031 244248
rect 17211 244217 17241 244248
rect 17421 244222 17451 244248
rect 17631 244217 17661 244248
rect 17841 244222 17871 244248
rect 18051 244217 18081 244248
rect 18261 244222 18291 244248
rect 18471 244217 18501 244248
rect 18681 244222 18711 244248
rect 18891 244217 18921 244248
rect 19101 244222 19131 244248
rect 19311 244217 19341 244248
rect 19521 244222 19551 244248
rect 19731 244217 19761 244248
rect 19941 244222 19971 244248
rect 20151 244217 20181 244248
rect 20361 244222 20391 244248
rect 20571 244217 20601 244248
rect 20781 244222 20811 244248
rect 20991 244217 21021 244248
rect 21201 244222 21231 244248
rect 21411 244217 21441 244248
rect 21621 244222 21651 244248
rect 21831 244217 21861 244248
rect 22041 244222 22071 244248
rect 22251 244217 22281 244248
rect 22461 244222 22491 244248
rect 22671 244217 22701 244248
rect 22881 244222 22911 244248
rect 23091 244217 23121 244248
rect 23301 244222 23331 244248
rect 23511 244217 23541 244248
rect 23721 244222 23751 244248
rect 23931 244217 23961 244248
rect 24141 244222 24171 244248
rect 24351 244217 24381 244248
rect 24561 244222 24591 244248
rect 24771 244217 24801 244248
rect 24981 244222 25011 244248
rect 25191 244217 25221 244248
rect 25401 244222 25431 244248
rect 25611 244217 25641 244248
rect 25821 244222 25851 244248
rect 26031 244217 26061 244248
rect 26241 244222 26271 244248
rect 26451 244217 26481 244248
rect 26661 244222 26691 244248
rect 26871 244217 26901 244248
rect 27081 244222 27111 244248
rect 27291 244217 27321 244248
rect -3807 244201 -3678 244217
rect -3807 244167 -3791 244201
rect -3695 244167 -3678 244201
rect -3807 244151 -3678 244167
rect -3387 244201 -3258 244217
rect -3387 244167 -3371 244201
rect -3275 244167 -3258 244201
rect -3387 244151 -3258 244167
rect -2967 244201 -2838 244217
rect -2967 244167 -2951 244201
rect -2855 244167 -2838 244201
rect -2967 244151 -2838 244167
rect -2547 244201 -2418 244217
rect -2547 244167 -2531 244201
rect -2435 244167 -2418 244201
rect -2547 244151 -2418 244167
rect -2127 244201 -1998 244217
rect -2127 244167 -2111 244201
rect -2015 244167 -1998 244201
rect -2127 244151 -1998 244167
rect -1707 244201 -1578 244217
rect -1707 244167 -1691 244201
rect -1595 244167 -1578 244201
rect -1707 244151 -1578 244167
rect -1287 244201 -1158 244217
rect -1287 244167 -1271 244201
rect -1175 244167 -1158 244201
rect -1287 244151 -1158 244167
rect -867 244201 -738 244217
rect -867 244167 -851 244201
rect -755 244167 -738 244201
rect -867 244151 -738 244167
rect -447 244201 -318 244217
rect -447 244167 -431 244201
rect -335 244167 -318 244201
rect -447 244151 -318 244167
rect -27 244201 102 244217
rect -27 244167 -11 244201
rect 85 244167 102 244201
rect -27 244151 102 244167
rect 393 244201 522 244217
rect 393 244167 409 244201
rect 505 244167 522 244201
rect 393 244151 522 244167
rect 813 244201 942 244217
rect 813 244167 829 244201
rect 925 244167 942 244201
rect 813 244151 942 244167
rect 1233 244201 1362 244217
rect 1233 244167 1249 244201
rect 1345 244167 1362 244201
rect 1233 244151 1362 244167
rect 1653 244201 1782 244217
rect 1653 244167 1669 244201
rect 1765 244167 1782 244201
rect 1653 244151 1782 244167
rect 2073 244201 2202 244217
rect 2073 244167 2089 244201
rect 2185 244167 2202 244201
rect 2073 244151 2202 244167
rect 2493 244201 2622 244217
rect 2493 244167 2509 244201
rect 2605 244167 2622 244201
rect 2493 244151 2622 244167
rect 2913 244201 3042 244217
rect 2913 244167 2929 244201
rect 3025 244167 3042 244201
rect 2913 244151 3042 244167
rect 3333 244201 3462 244217
rect 3333 244167 3349 244201
rect 3445 244167 3462 244201
rect 3333 244151 3462 244167
rect 3753 244201 3882 244217
rect 3753 244167 3769 244201
rect 3865 244167 3882 244201
rect 3753 244151 3882 244167
rect 4173 244201 4302 244217
rect 4173 244167 4189 244201
rect 4285 244167 4302 244201
rect 4173 244151 4302 244167
rect 4593 244201 4722 244217
rect 4593 244167 4609 244201
rect 4705 244167 4722 244201
rect 4593 244151 4722 244167
rect 5013 244201 5142 244217
rect 5013 244167 5029 244201
rect 5125 244167 5142 244201
rect 5013 244151 5142 244167
rect 5433 244201 5562 244217
rect 5433 244167 5449 244201
rect 5545 244167 5562 244201
rect 5433 244151 5562 244167
rect 5853 244201 5982 244217
rect 5853 244167 5869 244201
rect 5965 244167 5982 244201
rect 5853 244151 5982 244167
rect 6273 244201 6402 244217
rect 6273 244167 6289 244201
rect 6385 244167 6402 244201
rect 6273 244151 6402 244167
rect 6693 244201 6822 244217
rect 6693 244167 6709 244201
rect 6805 244167 6822 244201
rect 6693 244151 6822 244167
rect 7113 244201 7242 244217
rect 7113 244167 7129 244201
rect 7225 244167 7242 244201
rect 7113 244151 7242 244167
rect 7533 244201 7662 244217
rect 7533 244167 7549 244201
rect 7645 244167 7662 244201
rect 7533 244151 7662 244167
rect 7953 244201 8082 244217
rect 7953 244167 7969 244201
rect 8065 244167 8082 244201
rect 7953 244151 8082 244167
rect 8373 244201 8502 244217
rect 8373 244167 8389 244201
rect 8485 244167 8502 244201
rect 8373 244151 8502 244167
rect 8793 244201 8922 244217
rect 8793 244167 8809 244201
rect 8905 244167 8922 244201
rect 8793 244151 8922 244167
rect 9213 244201 9342 244217
rect 9213 244167 9229 244201
rect 9325 244167 9342 244201
rect 9213 244151 9342 244167
rect 9633 244201 9762 244217
rect 9633 244167 9649 244201
rect 9745 244167 9762 244201
rect 9633 244151 9762 244167
rect 10053 244201 10182 244217
rect 10053 244167 10069 244201
rect 10165 244167 10182 244201
rect 10053 244151 10182 244167
rect 10473 244201 10602 244217
rect 10473 244167 10489 244201
rect 10585 244167 10602 244201
rect 10473 244151 10602 244167
rect 10893 244201 11022 244217
rect 10893 244167 10909 244201
rect 11005 244167 11022 244201
rect 10893 244151 11022 244167
rect 11313 244201 11442 244217
rect 11313 244167 11329 244201
rect 11425 244167 11442 244201
rect 11313 244151 11442 244167
rect 11733 244201 11862 244217
rect 11733 244167 11749 244201
rect 11845 244167 11862 244201
rect 11733 244151 11862 244167
rect 12153 244201 12282 244217
rect 12153 244167 12169 244201
rect 12265 244167 12282 244201
rect 12153 244151 12282 244167
rect 12573 244201 12702 244217
rect 12573 244167 12589 244201
rect 12685 244167 12702 244201
rect 12573 244151 12702 244167
rect 12993 244201 13122 244217
rect 12993 244167 13009 244201
rect 13105 244167 13122 244201
rect 12993 244151 13122 244167
rect 13413 244201 13542 244217
rect 13413 244167 13429 244201
rect 13525 244167 13542 244201
rect 13413 244151 13542 244167
rect 13833 244201 13962 244217
rect 13833 244167 13849 244201
rect 13945 244167 13962 244201
rect 13833 244151 13962 244167
rect 14253 244201 14382 244217
rect 14253 244167 14269 244201
rect 14365 244167 14382 244201
rect 14253 244151 14382 244167
rect 14673 244201 14802 244217
rect 14673 244167 14689 244201
rect 14785 244167 14802 244201
rect 14673 244151 14802 244167
rect 15093 244201 15222 244217
rect 15093 244167 15109 244201
rect 15205 244167 15222 244201
rect 15093 244151 15222 244167
rect 15513 244201 15642 244217
rect 15513 244167 15529 244201
rect 15625 244167 15642 244201
rect 15513 244151 15642 244167
rect 15933 244201 16062 244217
rect 15933 244167 15949 244201
rect 16045 244167 16062 244201
rect 15933 244151 16062 244167
rect 16353 244201 16482 244217
rect 16353 244167 16369 244201
rect 16465 244167 16482 244201
rect 16353 244151 16482 244167
rect 16773 244201 16902 244217
rect 16773 244167 16789 244201
rect 16885 244167 16902 244201
rect 16773 244151 16902 244167
rect 17193 244201 17322 244217
rect 17193 244167 17209 244201
rect 17305 244167 17322 244201
rect 17193 244151 17322 244167
rect 17613 244201 17742 244217
rect 17613 244167 17629 244201
rect 17725 244167 17742 244201
rect 17613 244151 17742 244167
rect 18033 244201 18162 244217
rect 18033 244167 18049 244201
rect 18145 244167 18162 244201
rect 18033 244151 18162 244167
rect 18453 244201 18582 244217
rect 18453 244167 18469 244201
rect 18565 244167 18582 244201
rect 18453 244151 18582 244167
rect 18873 244201 19002 244217
rect 18873 244167 18889 244201
rect 18985 244167 19002 244201
rect 18873 244151 19002 244167
rect 19293 244201 19422 244217
rect 19293 244167 19309 244201
rect 19405 244167 19422 244201
rect 19293 244151 19422 244167
rect 19713 244201 19842 244217
rect 19713 244167 19729 244201
rect 19825 244167 19842 244201
rect 19713 244151 19842 244167
rect 20133 244201 20262 244217
rect 20133 244167 20149 244201
rect 20245 244167 20262 244201
rect 20133 244151 20262 244167
rect 20553 244201 20682 244217
rect 20553 244167 20569 244201
rect 20665 244167 20682 244201
rect 20553 244151 20682 244167
rect 20973 244201 21102 244217
rect 20973 244167 20989 244201
rect 21085 244167 21102 244201
rect 20973 244151 21102 244167
rect 21393 244201 21522 244217
rect 21393 244167 21409 244201
rect 21505 244167 21522 244201
rect 21393 244151 21522 244167
rect 21813 244201 21942 244217
rect 21813 244167 21829 244201
rect 21925 244167 21942 244201
rect 21813 244151 21942 244167
rect 22233 244201 22362 244217
rect 22233 244167 22249 244201
rect 22345 244167 22362 244201
rect 22233 244151 22362 244167
rect 22653 244201 22782 244217
rect 22653 244167 22669 244201
rect 22765 244167 22782 244201
rect 22653 244151 22782 244167
rect 23073 244201 23202 244217
rect 23073 244167 23089 244201
rect 23185 244167 23202 244201
rect 23073 244151 23202 244167
rect 23493 244201 23622 244217
rect 23493 244167 23509 244201
rect 23605 244167 23622 244201
rect 23493 244151 23622 244167
rect 23913 244201 24042 244217
rect 23913 244167 23929 244201
rect 24025 244167 24042 244201
rect 23913 244151 24042 244167
rect 24333 244201 24462 244217
rect 24333 244167 24349 244201
rect 24445 244167 24462 244201
rect 24333 244151 24462 244167
rect 24753 244201 24882 244217
rect 24753 244167 24769 244201
rect 24865 244167 24882 244201
rect 24753 244151 24882 244167
rect 25173 244201 25302 244217
rect 25173 244167 25189 244201
rect 25285 244167 25302 244201
rect 25173 244151 25302 244167
rect 25593 244201 25722 244217
rect 25593 244167 25609 244201
rect 25705 244167 25722 244201
rect 25593 244151 25722 244167
rect 26013 244201 26142 244217
rect 26013 244167 26029 244201
rect 26125 244167 26142 244201
rect 26013 244151 26142 244167
rect 26433 244201 26562 244217
rect 26433 244167 26449 244201
rect 26545 244167 26562 244201
rect 26433 244151 26562 244167
rect 26853 244201 26982 244217
rect 26853 244167 26869 244201
rect 26965 244167 26982 244201
rect 26853 244151 26982 244167
rect 27273 244201 27402 244217
rect 27273 244167 27289 244201
rect 27385 244167 27402 244201
rect 27273 244151 27402 244167
<< polycont >>
rect -4001 264076 -3905 264110
rect -3581 264076 -3485 264110
rect -3161 264076 -3065 264110
rect -2741 264076 -2645 264110
rect -2321 264076 -2225 264110
rect -1901 264076 -1805 264110
rect -1481 264076 -1385 264110
rect -1061 264076 -965 264110
rect -641 264076 -545 264110
rect -221 264076 -125 264110
rect 199 264076 295 264110
rect 619 264076 715 264110
rect 1039 264076 1135 264110
rect 1459 264076 1555 264110
rect 1879 264076 1975 264110
rect 2299 264076 2395 264110
rect 2719 264076 2815 264110
rect 3139 264076 3235 264110
rect 3559 264076 3655 264110
rect 3979 264076 4075 264110
rect 4399 264076 4495 264110
rect 4819 264076 4915 264110
rect 5239 264076 5335 264110
rect 5659 264076 5755 264110
rect 6079 264076 6175 264110
rect 6499 264076 6595 264110
rect 6919 264076 7015 264110
rect 7339 264076 7435 264110
rect 7759 264076 7855 264110
rect 8179 264076 8275 264110
rect 8599 264076 8695 264110
rect 9019 264076 9115 264110
rect 9439 264076 9535 264110
rect 9859 264076 9955 264110
rect 10279 264076 10375 264110
rect 10699 264076 10795 264110
rect 11119 264076 11215 264110
rect 11539 264076 11635 264110
rect 11959 264076 12055 264110
rect 12379 264076 12475 264110
rect 12799 264076 12895 264110
rect 13219 264076 13315 264110
rect 13639 264076 13735 264110
rect 14059 264076 14155 264110
rect 14479 264076 14575 264110
rect 14899 264076 14995 264110
rect 15319 264076 15415 264110
rect 15739 264076 15835 264110
rect 16159 264076 16255 264110
rect 16579 264076 16675 264110
rect 16999 264076 17095 264110
rect 17419 264076 17515 264110
rect 17839 264076 17935 264110
rect 18259 264076 18355 264110
rect 18679 264076 18775 264110
rect 19099 264076 19195 264110
rect 19519 264076 19615 264110
rect 19939 264076 20035 264110
rect 20359 264076 20455 264110
rect 20779 264076 20875 264110
rect 21199 264076 21295 264110
rect 21619 264076 21715 264110
rect 22039 264076 22135 264110
rect 22459 264076 22555 264110
rect 22879 264076 22975 264110
rect 23299 264076 23395 264110
rect 23719 264076 23815 264110
rect 24139 264076 24235 264110
rect 24559 264076 24655 264110
rect 24979 264076 25075 264110
rect 25399 264076 25495 264110
rect 25819 264076 25915 264110
rect 26239 264076 26335 264110
rect 26659 264076 26755 264110
rect 27079 264076 27175 264110
rect -3791 263164 -3757 263198
rect -3791 263056 -3757 263090
rect -3371 263164 -3337 263198
rect -3371 263056 -3337 263090
rect -2951 263164 -2917 263198
rect -2951 263056 -2917 263090
rect -2531 263164 -2497 263198
rect -2531 263056 -2497 263090
rect -2111 263164 -2077 263198
rect -2111 263056 -2077 263090
rect -1691 263164 -1657 263198
rect -1691 263056 -1657 263090
rect -1271 263164 -1237 263198
rect -1271 263056 -1237 263090
rect -851 263164 -817 263198
rect -851 263056 -817 263090
rect -431 263164 -397 263198
rect -431 263056 -397 263090
rect -11 263164 23 263198
rect -11 263056 23 263090
rect 409 263164 443 263198
rect 409 263056 443 263090
rect 829 263164 863 263198
rect 829 263056 863 263090
rect 1249 263164 1283 263198
rect 1249 263056 1283 263090
rect 1669 263164 1703 263198
rect 1669 263056 1703 263090
rect 2089 263164 2123 263198
rect 2089 263056 2123 263090
rect 2509 263164 2543 263198
rect 2509 263056 2543 263090
rect 2929 263164 2963 263198
rect 2929 263056 2963 263090
rect 3349 263164 3383 263198
rect 3349 263056 3383 263090
rect 3769 263164 3803 263198
rect 3769 263056 3803 263090
rect 4189 263164 4223 263198
rect 4189 263056 4223 263090
rect 4609 263164 4643 263198
rect 4609 263056 4643 263090
rect 5029 263164 5063 263198
rect 5029 263056 5063 263090
rect 5449 263164 5483 263198
rect 5449 263056 5483 263090
rect 5869 263164 5903 263198
rect 5869 263056 5903 263090
rect 6289 263164 6323 263198
rect 6289 263056 6323 263090
rect 6709 263164 6743 263198
rect 6709 263056 6743 263090
rect 7129 263164 7163 263198
rect 7129 263056 7163 263090
rect 7549 263164 7583 263198
rect 7549 263056 7583 263090
rect 7969 263164 8003 263198
rect 7969 263056 8003 263090
rect 8389 263164 8423 263198
rect 8389 263056 8423 263090
rect 8809 263164 8843 263198
rect 8809 263056 8843 263090
rect 9229 263164 9263 263198
rect 9229 263056 9263 263090
rect 9649 263164 9683 263198
rect 9649 263056 9683 263090
rect 10069 263164 10103 263198
rect 10069 263056 10103 263090
rect 10489 263164 10523 263198
rect 10489 263056 10523 263090
rect 10909 263164 10943 263198
rect 10909 263056 10943 263090
rect 11329 263164 11363 263198
rect 11329 263056 11363 263090
rect 11749 263164 11783 263198
rect 11749 263056 11783 263090
rect 12169 263164 12203 263198
rect 12169 263056 12203 263090
rect 12589 263164 12623 263198
rect 12589 263056 12623 263090
rect 13009 263164 13043 263198
rect 13009 263056 13043 263090
rect 13429 263164 13463 263198
rect 13429 263056 13463 263090
rect 13849 263164 13883 263198
rect 13849 263056 13883 263090
rect 14269 263164 14303 263198
rect 14269 263056 14303 263090
rect 14689 263164 14723 263198
rect 14689 263056 14723 263090
rect 15109 263164 15143 263198
rect 15109 263056 15143 263090
rect 15529 263164 15563 263198
rect 15529 263056 15563 263090
rect 15949 263164 15983 263198
rect 15949 263056 15983 263090
rect 16369 263164 16403 263198
rect 16369 263056 16403 263090
rect 16789 263164 16823 263198
rect 16789 263056 16823 263090
rect 17209 263164 17243 263198
rect 17209 263056 17243 263090
rect 17629 263164 17663 263198
rect 17629 263056 17663 263090
rect 18049 263164 18083 263198
rect 18049 263056 18083 263090
rect 18469 263164 18503 263198
rect 18469 263056 18503 263090
rect 18889 263164 18923 263198
rect 18889 263056 18923 263090
rect 19309 263164 19343 263198
rect 19309 263056 19343 263090
rect 19729 263164 19763 263198
rect 19729 263056 19763 263090
rect 20149 263164 20183 263198
rect 20149 263056 20183 263090
rect 20569 263164 20603 263198
rect 20569 263056 20603 263090
rect 20989 263164 21023 263198
rect 20989 263056 21023 263090
rect 21409 263164 21443 263198
rect 21409 263056 21443 263090
rect 21829 263164 21863 263198
rect 21829 263056 21863 263090
rect 22249 263164 22283 263198
rect 22249 263056 22283 263090
rect 22669 263164 22703 263198
rect 22669 263056 22703 263090
rect 23089 263164 23123 263198
rect 23089 263056 23123 263090
rect 23509 263164 23543 263198
rect 23509 263056 23543 263090
rect 23929 263164 23963 263198
rect 23929 263056 23963 263090
rect 24349 263164 24383 263198
rect 24349 263056 24383 263090
rect 24769 263164 24803 263198
rect 24769 263056 24803 263090
rect 25189 263164 25223 263198
rect 25189 263056 25223 263090
rect 25609 263164 25643 263198
rect 25609 263056 25643 263090
rect 26029 263164 26063 263198
rect 26029 263056 26063 263090
rect 26449 263164 26483 263198
rect 26449 263056 26483 263090
rect 26869 263164 26903 263198
rect 26869 263056 26903 263090
rect 27289 263164 27323 263198
rect 27289 263056 27323 263090
rect -4001 262144 -3905 262178
rect -3581 262144 -3485 262178
rect -3161 262144 -3065 262178
rect -2741 262144 -2645 262178
rect -2321 262144 -2225 262178
rect -1901 262144 -1805 262178
rect -1481 262144 -1385 262178
rect -1061 262144 -965 262178
rect -641 262144 -545 262178
rect -221 262144 -125 262178
rect 199 262144 295 262178
rect 619 262144 715 262178
rect 1039 262144 1135 262178
rect 1459 262144 1555 262178
rect 1879 262144 1975 262178
rect 2299 262144 2395 262178
rect 2719 262144 2815 262178
rect 3139 262144 3235 262178
rect 3559 262144 3655 262178
rect 3979 262144 4075 262178
rect 4399 262144 4495 262178
rect 4819 262144 4915 262178
rect 5239 262144 5335 262178
rect 5659 262144 5755 262178
rect 6079 262144 6175 262178
rect 6499 262144 6595 262178
rect 6919 262144 7015 262178
rect 7339 262144 7435 262178
rect 7759 262144 7855 262178
rect 8179 262144 8275 262178
rect 8599 262144 8695 262178
rect 9019 262144 9115 262178
rect 9439 262144 9535 262178
rect 9859 262144 9955 262178
rect 10279 262144 10375 262178
rect 10699 262144 10795 262178
rect 11119 262144 11215 262178
rect 11539 262144 11635 262178
rect 11959 262144 12055 262178
rect 12379 262144 12475 262178
rect 12799 262144 12895 262178
rect 13219 262144 13315 262178
rect 13639 262144 13735 262178
rect 14059 262144 14155 262178
rect 14479 262144 14575 262178
rect 14899 262144 14995 262178
rect 15319 262144 15415 262178
rect 15739 262144 15835 262178
rect 16159 262144 16255 262178
rect 16579 262144 16675 262178
rect 16999 262144 17095 262178
rect 17419 262144 17515 262178
rect 17839 262144 17935 262178
rect 18259 262144 18355 262178
rect 18679 262144 18775 262178
rect 19099 262144 19195 262178
rect 19519 262144 19615 262178
rect 19939 262144 20035 262178
rect 20359 262144 20455 262178
rect 20779 262144 20875 262178
rect 21199 262144 21295 262178
rect 21619 262144 21715 262178
rect 22039 262144 22135 262178
rect 22459 262144 22555 262178
rect 22879 262144 22975 262178
rect 23299 262144 23395 262178
rect 23719 262144 23815 262178
rect 24139 262144 24235 262178
rect 24559 262144 24655 262178
rect 24979 262144 25075 262178
rect 25399 262144 25495 262178
rect 25819 262144 25915 262178
rect 26239 262144 26335 262178
rect 26659 262144 26755 262178
rect 27079 262144 27175 262178
rect -4001 254548 -3905 254582
rect -3581 254548 -3485 254582
rect -3161 254548 -3065 254582
rect -2741 254548 -2645 254582
rect -2321 254548 -2225 254582
rect -1901 254548 -1805 254582
rect -1481 254548 -1385 254582
rect -1061 254548 -965 254582
rect -641 254548 -545 254582
rect -221 254548 -125 254582
rect 199 254548 295 254582
rect 619 254548 715 254582
rect 1039 254548 1135 254582
rect 1459 254548 1555 254582
rect 1879 254548 1975 254582
rect 2299 254548 2395 254582
rect 2719 254548 2815 254582
rect 3139 254548 3235 254582
rect 3559 254548 3655 254582
rect 3979 254548 4075 254582
rect 4399 254548 4495 254582
rect 4819 254548 4915 254582
rect 5239 254548 5335 254582
rect 5659 254548 5755 254582
rect 6079 254548 6175 254582
rect 6499 254548 6595 254582
rect 6919 254548 7015 254582
rect 7339 254548 7435 254582
rect 7759 254548 7855 254582
rect 8179 254548 8275 254582
rect 8599 254548 8695 254582
rect 9019 254548 9115 254582
rect 9439 254548 9535 254582
rect 9859 254548 9955 254582
rect 10279 254548 10375 254582
rect 10699 254548 10795 254582
rect 11119 254548 11215 254582
rect 11539 254548 11635 254582
rect 11959 254548 12055 254582
rect 12379 254548 12475 254582
rect 12799 254548 12895 254582
rect 13219 254548 13315 254582
rect 13639 254548 13735 254582
rect 14059 254548 14155 254582
rect 14479 254548 14575 254582
rect 14899 254548 14995 254582
rect 15319 254548 15415 254582
rect 15739 254548 15835 254582
rect 16159 254548 16255 254582
rect 16579 254548 16675 254582
rect 16999 254548 17095 254582
rect 17419 254548 17515 254582
rect 17839 254548 17935 254582
rect 18259 254548 18355 254582
rect 18679 254548 18775 254582
rect 19099 254548 19195 254582
rect 19519 254548 19615 254582
rect 19939 254548 20035 254582
rect 20359 254548 20455 254582
rect 20779 254548 20875 254582
rect 21199 254548 21295 254582
rect 21619 254548 21715 254582
rect 22039 254548 22135 254582
rect 22459 254548 22555 254582
rect 22879 254548 22975 254582
rect 23299 254548 23395 254582
rect 23719 254548 23815 254582
rect 24139 254548 24235 254582
rect 24559 254548 24655 254582
rect 24979 254548 25075 254582
rect 25399 254548 25495 254582
rect 25819 254548 25915 254582
rect 26239 254548 26335 254582
rect 26659 254548 26755 254582
rect 27079 254548 27175 254582
rect -3791 253512 -3757 253654
rect -3371 253512 -3337 253654
rect -2951 253512 -2917 253654
rect -2531 253512 -2497 253654
rect -2111 253512 -2077 253654
rect -1691 253512 -1657 253654
rect -1271 253512 -1237 253654
rect -851 253512 -817 253654
rect -431 253512 -397 253654
rect -11 253512 23 253654
rect 409 253512 443 253654
rect 829 253512 863 253654
rect 1249 253512 1283 253654
rect 1669 253512 1703 253654
rect 2089 253512 2123 253654
rect 2509 253512 2543 253654
rect 2929 253512 2963 253654
rect 3349 253512 3383 253654
rect 3769 253512 3803 253654
rect 4189 253512 4223 253654
rect 4609 253512 4643 253654
rect 5029 253512 5063 253654
rect 5449 253512 5483 253654
rect 5869 253512 5903 253654
rect 6289 253512 6323 253654
rect 6709 253512 6743 253654
rect 7129 253512 7163 253654
rect 7549 253512 7583 253654
rect 7969 253512 8003 253654
rect 8389 253512 8423 253654
rect 8809 253512 8843 253654
rect 9229 253512 9263 253654
rect 9649 253512 9683 253654
rect 10069 253512 10103 253654
rect 10489 253512 10523 253654
rect 10909 253512 10943 253654
rect 11329 253512 11363 253654
rect 11749 253512 11783 253654
rect 12169 253512 12203 253654
rect 12589 253512 12623 253654
rect 13009 253512 13043 253654
rect 13429 253512 13463 253654
rect 13849 253512 13883 253654
rect 14269 253512 14303 253654
rect 14689 253512 14723 253654
rect 15109 253512 15143 253654
rect 15529 253512 15563 253654
rect 15949 253512 15983 253654
rect 16369 253512 16403 253654
rect 16789 253512 16823 253654
rect 17209 253512 17243 253654
rect 17629 253512 17663 253654
rect 18049 253512 18083 253654
rect 18469 253512 18503 253654
rect 18889 253512 18923 253654
rect 19309 253512 19343 253654
rect 19729 253512 19763 253654
rect 20149 253512 20183 253654
rect 20569 253512 20603 253654
rect 20989 253512 21023 253654
rect 21409 253512 21443 253654
rect 21829 253512 21863 253654
rect 22249 253512 22283 253654
rect 22669 253512 22703 253654
rect 23089 253512 23123 253654
rect 23509 253512 23543 253654
rect 23929 253512 23963 253654
rect 24349 253512 24383 253654
rect 24769 253512 24803 253654
rect 25189 253512 25223 253654
rect 25609 253512 25643 253654
rect 26029 253512 26063 253654
rect 26449 253512 26483 253654
rect 26869 253512 26903 253654
rect 27289 253512 27323 253654
rect -4001 252476 -3967 252618
rect -3581 252476 -3547 252618
rect -3161 252476 -3127 252618
rect -2741 252476 -2707 252618
rect -2321 252476 -2287 252618
rect -1901 252476 -1867 252618
rect -1481 252476 -1447 252618
rect -1061 252476 -1027 252618
rect -641 252476 -607 252618
rect -221 252476 -187 252618
rect 199 252476 233 252618
rect 619 252476 653 252618
rect 1039 252476 1073 252618
rect 1459 252476 1493 252618
rect 1879 252476 1913 252618
rect 2299 252476 2333 252618
rect 2719 252476 2753 252618
rect 3139 252476 3173 252618
rect 3559 252476 3593 252618
rect 3979 252476 4013 252618
rect 4399 252476 4433 252618
rect 4819 252476 4853 252618
rect 5239 252476 5273 252618
rect 5659 252476 5693 252618
rect 6079 252476 6113 252618
rect 6499 252476 6533 252618
rect 6919 252476 6953 252618
rect 7339 252476 7373 252618
rect 7759 252476 7793 252618
rect 8179 252476 8213 252618
rect 8599 252476 8633 252618
rect 9019 252476 9053 252618
rect 9439 252476 9473 252618
rect 9859 252476 9893 252618
rect 10279 252476 10313 252618
rect 10699 252476 10733 252618
rect 11119 252476 11153 252618
rect 11539 252476 11573 252618
rect 11959 252476 11993 252618
rect 12379 252476 12413 252618
rect 12799 252476 12833 252618
rect 13219 252476 13253 252618
rect 13639 252476 13673 252618
rect 14059 252476 14093 252618
rect 14479 252476 14513 252618
rect 14899 252476 14933 252618
rect 15319 252476 15353 252618
rect 15739 252476 15773 252618
rect 16159 252476 16193 252618
rect 16579 252476 16613 252618
rect 16999 252476 17033 252618
rect 17419 252476 17453 252618
rect 17839 252476 17873 252618
rect 18259 252476 18293 252618
rect 18679 252476 18713 252618
rect 19099 252476 19133 252618
rect 19519 252476 19553 252618
rect 19939 252476 19973 252618
rect 20359 252476 20393 252618
rect 20779 252476 20813 252618
rect 21199 252476 21233 252618
rect 21619 252476 21653 252618
rect 22039 252476 22073 252618
rect 22459 252476 22493 252618
rect 22879 252476 22913 252618
rect 23299 252476 23333 252618
rect 23719 252476 23753 252618
rect 24139 252476 24173 252618
rect 24559 252476 24593 252618
rect 24979 252476 25013 252618
rect 25399 252476 25433 252618
rect 25819 252476 25853 252618
rect 26239 252476 26273 252618
rect 26659 252476 26693 252618
rect 27079 252476 27113 252618
rect -3791 251440 -3757 251582
rect -3371 251440 -3337 251582
rect -2951 251440 -2917 251582
rect -2531 251440 -2497 251582
rect -2111 251440 -2077 251582
rect -1691 251440 -1657 251582
rect -1271 251440 -1237 251582
rect -851 251440 -817 251582
rect -431 251440 -397 251582
rect -11 251440 23 251582
rect 409 251440 443 251582
rect 829 251440 863 251582
rect 1249 251440 1283 251582
rect 1669 251440 1703 251582
rect 2089 251440 2123 251582
rect 2509 251440 2543 251582
rect 2929 251440 2963 251582
rect 3349 251440 3383 251582
rect 3769 251440 3803 251582
rect 4189 251440 4223 251582
rect 4609 251440 4643 251582
rect 5029 251440 5063 251582
rect 5449 251440 5483 251582
rect 5869 251440 5903 251582
rect 6289 251440 6323 251582
rect 6709 251440 6743 251582
rect 7129 251440 7163 251582
rect 7549 251440 7583 251582
rect 7969 251440 8003 251582
rect 8389 251440 8423 251582
rect 8809 251440 8843 251582
rect 9229 251440 9263 251582
rect 9649 251440 9683 251582
rect 10069 251440 10103 251582
rect 10489 251440 10523 251582
rect 10909 251440 10943 251582
rect 11329 251440 11363 251582
rect 11749 251440 11783 251582
rect 12169 251440 12203 251582
rect 12589 251440 12623 251582
rect 13009 251440 13043 251582
rect 13429 251440 13463 251582
rect 13849 251440 13883 251582
rect 14269 251440 14303 251582
rect 14689 251440 14723 251582
rect 15109 251440 15143 251582
rect 15529 251440 15563 251582
rect 15949 251440 15983 251582
rect 16369 251440 16403 251582
rect 16789 251440 16823 251582
rect 17209 251440 17243 251582
rect 17629 251440 17663 251582
rect 18049 251440 18083 251582
rect 18469 251440 18503 251582
rect 18889 251440 18923 251582
rect 19309 251440 19343 251582
rect 19729 251440 19763 251582
rect 20149 251440 20183 251582
rect 20569 251440 20603 251582
rect 20989 251440 21023 251582
rect 21409 251440 21443 251582
rect 21829 251440 21863 251582
rect 22249 251440 22283 251582
rect 22669 251440 22703 251582
rect 23089 251440 23123 251582
rect 23509 251440 23543 251582
rect 23929 251440 23963 251582
rect 24349 251440 24383 251582
rect 24769 251440 24803 251582
rect 25189 251440 25223 251582
rect 25609 251440 25643 251582
rect 26029 251440 26063 251582
rect 26449 251440 26483 251582
rect 26869 251440 26903 251582
rect 27289 251440 27323 251582
rect -4001 250404 -3967 250546
rect -3581 250404 -3547 250546
rect -3161 250404 -3127 250546
rect -2741 250404 -2707 250546
rect -2321 250404 -2287 250546
rect -1901 250404 -1867 250546
rect -1481 250404 -1447 250546
rect -1061 250404 -1027 250546
rect -641 250404 -607 250546
rect -221 250404 -187 250546
rect 199 250404 233 250546
rect 619 250404 653 250546
rect 1039 250404 1073 250546
rect 1459 250404 1493 250546
rect 1879 250404 1913 250546
rect 2299 250404 2333 250546
rect 2719 250404 2753 250546
rect 3139 250404 3173 250546
rect 3559 250404 3593 250546
rect 3979 250404 4013 250546
rect 4399 250404 4433 250546
rect 4819 250404 4853 250546
rect 5239 250404 5273 250546
rect 5659 250404 5693 250546
rect 6079 250404 6113 250546
rect 6499 250404 6533 250546
rect 6919 250404 6953 250546
rect 7339 250404 7373 250546
rect 7759 250404 7793 250546
rect 8179 250404 8213 250546
rect 8599 250404 8633 250546
rect 9019 250404 9053 250546
rect 9439 250404 9473 250546
rect 9859 250404 9893 250546
rect 10279 250404 10313 250546
rect 10699 250404 10733 250546
rect 11119 250404 11153 250546
rect 11539 250404 11573 250546
rect 11959 250404 11993 250546
rect 12379 250404 12413 250546
rect 12799 250404 12833 250546
rect 13219 250404 13253 250546
rect 13639 250404 13673 250546
rect 14059 250404 14093 250546
rect 14479 250404 14513 250546
rect 14899 250404 14933 250546
rect 15319 250404 15353 250546
rect 15739 250404 15773 250546
rect 16159 250404 16193 250546
rect 16579 250404 16613 250546
rect 16999 250404 17033 250546
rect 17419 250404 17453 250546
rect 17839 250404 17873 250546
rect 18259 250404 18293 250546
rect 18679 250404 18713 250546
rect 19099 250404 19133 250546
rect 19519 250404 19553 250546
rect 19939 250404 19973 250546
rect 20359 250404 20393 250546
rect 20779 250404 20813 250546
rect 21199 250404 21233 250546
rect 21619 250404 21653 250546
rect 22039 250404 22073 250546
rect 22459 250404 22493 250546
rect 22879 250404 22913 250546
rect 23299 250404 23333 250546
rect 23719 250404 23753 250546
rect 24139 250404 24173 250546
rect 24559 250404 24593 250546
rect 24979 250404 25013 250546
rect 25399 250404 25433 250546
rect 25819 250404 25853 250546
rect 26239 250404 26273 250546
rect 26659 250404 26693 250546
rect 27079 250404 27113 250546
rect -3791 249476 -3695 249510
rect -3371 249476 -3275 249510
rect -2951 249476 -2855 249510
rect -2531 249476 -2435 249510
rect -2111 249476 -2015 249510
rect -1691 249476 -1595 249510
rect -1271 249476 -1175 249510
rect -851 249476 -755 249510
rect -431 249476 -335 249510
rect -11 249476 85 249510
rect 409 249476 505 249510
rect 829 249476 925 249510
rect 1249 249476 1345 249510
rect 1669 249476 1765 249510
rect 2089 249476 2185 249510
rect 2509 249476 2605 249510
rect 2929 249476 3025 249510
rect 3349 249476 3445 249510
rect 3769 249476 3865 249510
rect 4189 249476 4285 249510
rect 4609 249476 4705 249510
rect 5029 249476 5125 249510
rect 5449 249476 5545 249510
rect 5869 249476 5965 249510
rect 6289 249476 6385 249510
rect 6709 249476 6805 249510
rect 7129 249476 7225 249510
rect 7549 249476 7645 249510
rect 7969 249476 8065 249510
rect 8389 249476 8485 249510
rect 8809 249476 8905 249510
rect 9229 249476 9325 249510
rect 9649 249476 9745 249510
rect 10069 249476 10165 249510
rect 10489 249476 10585 249510
rect 10909 249476 11005 249510
rect 11329 249476 11425 249510
rect 11749 249476 11845 249510
rect 12169 249476 12265 249510
rect 12589 249476 12685 249510
rect 13009 249476 13105 249510
rect 13429 249476 13525 249510
rect 13849 249476 13945 249510
rect 14269 249476 14365 249510
rect 14689 249476 14785 249510
rect 15109 249476 15205 249510
rect 15529 249476 15625 249510
rect 15949 249476 16045 249510
rect 16369 249476 16465 249510
rect 16789 249476 16885 249510
rect 17209 249476 17305 249510
rect 17629 249476 17725 249510
rect 18049 249476 18145 249510
rect 18469 249476 18565 249510
rect 18889 249476 18985 249510
rect 19309 249476 19405 249510
rect 19729 249476 19825 249510
rect 20149 249476 20245 249510
rect 20569 249476 20665 249510
rect 20989 249476 21085 249510
rect 21409 249476 21505 249510
rect 21829 249476 21925 249510
rect 22249 249476 22345 249510
rect 22669 249476 22765 249510
rect 23089 249476 23185 249510
rect 23509 249476 23605 249510
rect 23929 249476 24025 249510
rect 24349 249476 24445 249510
rect 24769 249476 24865 249510
rect 25189 249476 25285 249510
rect 25609 249476 25705 249510
rect 26029 249476 26125 249510
rect 26449 249476 26545 249510
rect 26869 249476 26965 249510
rect 27289 249476 27385 249510
rect -4001 249239 -3905 249273
rect -3581 249239 -3485 249273
rect -3161 249239 -3065 249273
rect -2741 249239 -2645 249273
rect -2321 249239 -2225 249273
rect -1901 249239 -1805 249273
rect -1481 249239 -1385 249273
rect -1061 249239 -965 249273
rect -641 249239 -545 249273
rect -221 249239 -125 249273
rect 199 249239 295 249273
rect 619 249239 715 249273
rect 1039 249239 1135 249273
rect 1459 249239 1555 249273
rect 1879 249239 1975 249273
rect 2299 249239 2395 249273
rect 2719 249239 2815 249273
rect 3139 249239 3235 249273
rect 3559 249239 3655 249273
rect 3979 249239 4075 249273
rect 4399 249239 4495 249273
rect 4819 249239 4915 249273
rect 5239 249239 5335 249273
rect 5659 249239 5755 249273
rect 6079 249239 6175 249273
rect 6499 249239 6595 249273
rect 6919 249239 7015 249273
rect 7339 249239 7435 249273
rect 7759 249239 7855 249273
rect 8179 249239 8275 249273
rect 8599 249239 8695 249273
rect 9019 249239 9115 249273
rect 9439 249239 9535 249273
rect 9859 249239 9955 249273
rect 10279 249239 10375 249273
rect 10699 249239 10795 249273
rect 11119 249239 11215 249273
rect 11539 249239 11635 249273
rect 11959 249239 12055 249273
rect 12379 249239 12475 249273
rect 12799 249239 12895 249273
rect 13219 249239 13315 249273
rect 13639 249239 13735 249273
rect 14059 249239 14155 249273
rect 14479 249239 14575 249273
rect 14899 249239 14995 249273
rect 15319 249239 15415 249273
rect 15739 249239 15835 249273
rect 16159 249239 16255 249273
rect 16579 249239 16675 249273
rect 16999 249239 17095 249273
rect 17419 249239 17515 249273
rect 17839 249239 17935 249273
rect 18259 249239 18355 249273
rect 18679 249239 18775 249273
rect 19099 249239 19195 249273
rect 19519 249239 19615 249273
rect 19939 249239 20035 249273
rect 20359 249239 20455 249273
rect 20779 249239 20875 249273
rect 21199 249239 21295 249273
rect 21619 249239 21715 249273
rect 22039 249239 22135 249273
rect 22459 249239 22555 249273
rect 22879 249239 22975 249273
rect 23299 249239 23395 249273
rect 23719 249239 23815 249273
rect 24139 249239 24235 249273
rect 24559 249239 24655 249273
rect 24979 249239 25075 249273
rect 25399 249239 25495 249273
rect 25819 249239 25915 249273
rect 26239 249239 26335 249273
rect 26659 249239 26755 249273
rect 27079 249239 27175 249273
rect -3791 248203 -3757 248345
rect -3371 248203 -3337 248345
rect -2951 248203 -2917 248345
rect -2531 248203 -2497 248345
rect -2111 248203 -2077 248345
rect -1691 248203 -1657 248345
rect -1271 248203 -1237 248345
rect -851 248203 -817 248345
rect -431 248203 -397 248345
rect -11 248203 23 248345
rect 409 248203 443 248345
rect 829 248203 863 248345
rect 1249 248203 1283 248345
rect 1669 248203 1703 248345
rect 2089 248203 2123 248345
rect 2509 248203 2543 248345
rect 2929 248203 2963 248345
rect 3349 248203 3383 248345
rect 3769 248203 3803 248345
rect 4189 248203 4223 248345
rect 4609 248203 4643 248345
rect 5029 248203 5063 248345
rect 5449 248203 5483 248345
rect 5869 248203 5903 248345
rect 6289 248203 6323 248345
rect 6709 248203 6743 248345
rect 7129 248203 7163 248345
rect 7549 248203 7583 248345
rect 7969 248203 8003 248345
rect 8389 248203 8423 248345
rect 8809 248203 8843 248345
rect 9229 248203 9263 248345
rect 9649 248203 9683 248345
rect 10069 248203 10103 248345
rect 10489 248203 10523 248345
rect 10909 248203 10943 248345
rect 11329 248203 11363 248345
rect 11749 248203 11783 248345
rect 12169 248203 12203 248345
rect 12589 248203 12623 248345
rect 13009 248203 13043 248345
rect 13429 248203 13463 248345
rect 13849 248203 13883 248345
rect 14269 248203 14303 248345
rect 14689 248203 14723 248345
rect 15109 248203 15143 248345
rect 15529 248203 15563 248345
rect 15949 248203 15983 248345
rect 16369 248203 16403 248345
rect 16789 248203 16823 248345
rect 17209 248203 17243 248345
rect 17629 248203 17663 248345
rect 18049 248203 18083 248345
rect 18469 248203 18503 248345
rect 18889 248203 18923 248345
rect 19309 248203 19343 248345
rect 19729 248203 19763 248345
rect 20149 248203 20183 248345
rect 20569 248203 20603 248345
rect 20989 248203 21023 248345
rect 21409 248203 21443 248345
rect 21829 248203 21863 248345
rect 22249 248203 22283 248345
rect 22669 248203 22703 248345
rect 23089 248203 23123 248345
rect 23509 248203 23543 248345
rect 23929 248203 23963 248345
rect 24349 248203 24383 248345
rect 24769 248203 24803 248345
rect 25189 248203 25223 248345
rect 25609 248203 25643 248345
rect 26029 248203 26063 248345
rect 26449 248203 26483 248345
rect 26869 248203 26903 248345
rect 27289 248203 27323 248345
rect -4001 247167 -3967 247309
rect -3581 247167 -3547 247309
rect -3161 247167 -3127 247309
rect -2741 247167 -2707 247309
rect -2321 247167 -2287 247309
rect -1901 247167 -1867 247309
rect -1481 247167 -1447 247309
rect -1061 247167 -1027 247309
rect -641 247167 -607 247309
rect -221 247167 -187 247309
rect 199 247167 233 247309
rect 619 247167 653 247309
rect 1039 247167 1073 247309
rect 1459 247167 1493 247309
rect 1879 247167 1913 247309
rect 2299 247167 2333 247309
rect 2719 247167 2753 247309
rect 3139 247167 3173 247309
rect 3559 247167 3593 247309
rect 3979 247167 4013 247309
rect 4399 247167 4433 247309
rect 4819 247167 4853 247309
rect 5239 247167 5273 247309
rect 5659 247167 5693 247309
rect 6079 247167 6113 247309
rect 6499 247167 6533 247309
rect 6919 247167 6953 247309
rect 7339 247167 7373 247309
rect 7759 247167 7793 247309
rect 8179 247167 8213 247309
rect 8599 247167 8633 247309
rect 9019 247167 9053 247309
rect 9439 247167 9473 247309
rect 9859 247167 9893 247309
rect 10279 247167 10313 247309
rect 10699 247167 10733 247309
rect 11119 247167 11153 247309
rect 11539 247167 11573 247309
rect 11959 247167 11993 247309
rect 12379 247167 12413 247309
rect 12799 247167 12833 247309
rect 13219 247167 13253 247309
rect 13639 247167 13673 247309
rect 14059 247167 14093 247309
rect 14479 247167 14513 247309
rect 14899 247167 14933 247309
rect 15319 247167 15353 247309
rect 15739 247167 15773 247309
rect 16159 247167 16193 247309
rect 16579 247167 16613 247309
rect 16999 247167 17033 247309
rect 17419 247167 17453 247309
rect 17839 247167 17873 247309
rect 18259 247167 18293 247309
rect 18679 247167 18713 247309
rect 19099 247167 19133 247309
rect 19519 247167 19553 247309
rect 19939 247167 19973 247309
rect 20359 247167 20393 247309
rect 20779 247167 20813 247309
rect 21199 247167 21233 247309
rect 21619 247167 21653 247309
rect 22039 247167 22073 247309
rect 22459 247167 22493 247309
rect 22879 247167 22913 247309
rect 23299 247167 23333 247309
rect 23719 247167 23753 247309
rect 24139 247167 24173 247309
rect 24559 247167 24593 247309
rect 24979 247167 25013 247309
rect 25399 247167 25433 247309
rect 25819 247167 25853 247309
rect 26239 247167 26273 247309
rect 26659 247167 26693 247309
rect 27079 247167 27113 247309
rect -3791 246131 -3757 246273
rect -3371 246131 -3337 246273
rect -2951 246131 -2917 246273
rect -2531 246131 -2497 246273
rect -2111 246131 -2077 246273
rect -1691 246131 -1657 246273
rect -1271 246131 -1237 246273
rect -851 246131 -817 246273
rect -431 246131 -397 246273
rect -11 246131 23 246273
rect 409 246131 443 246273
rect 829 246131 863 246273
rect 1249 246131 1283 246273
rect 1669 246131 1703 246273
rect 2089 246131 2123 246273
rect 2509 246131 2543 246273
rect 2929 246131 2963 246273
rect 3349 246131 3383 246273
rect 3769 246131 3803 246273
rect 4189 246131 4223 246273
rect 4609 246131 4643 246273
rect 5029 246131 5063 246273
rect 5449 246131 5483 246273
rect 5869 246131 5903 246273
rect 6289 246131 6323 246273
rect 6709 246131 6743 246273
rect 7129 246131 7163 246273
rect 7549 246131 7583 246273
rect 7969 246131 8003 246273
rect 8389 246131 8423 246273
rect 8809 246131 8843 246273
rect 9229 246131 9263 246273
rect 9649 246131 9683 246273
rect 10069 246131 10103 246273
rect 10489 246131 10523 246273
rect 10909 246131 10943 246273
rect 11329 246131 11363 246273
rect 11749 246131 11783 246273
rect 12169 246131 12203 246273
rect 12589 246131 12623 246273
rect 13009 246131 13043 246273
rect 13429 246131 13463 246273
rect 13849 246131 13883 246273
rect 14269 246131 14303 246273
rect 14689 246131 14723 246273
rect 15109 246131 15143 246273
rect 15529 246131 15563 246273
rect 15949 246131 15983 246273
rect 16369 246131 16403 246273
rect 16789 246131 16823 246273
rect 17209 246131 17243 246273
rect 17629 246131 17663 246273
rect 18049 246131 18083 246273
rect 18469 246131 18503 246273
rect 18889 246131 18923 246273
rect 19309 246131 19343 246273
rect 19729 246131 19763 246273
rect 20149 246131 20183 246273
rect 20569 246131 20603 246273
rect 20989 246131 21023 246273
rect 21409 246131 21443 246273
rect 21829 246131 21863 246273
rect 22249 246131 22283 246273
rect 22669 246131 22703 246273
rect 23089 246131 23123 246273
rect 23509 246131 23543 246273
rect 23929 246131 23963 246273
rect 24349 246131 24383 246273
rect 24769 246131 24803 246273
rect 25189 246131 25223 246273
rect 25609 246131 25643 246273
rect 26029 246131 26063 246273
rect 26449 246131 26483 246273
rect 26869 246131 26903 246273
rect 27289 246131 27323 246273
rect -4001 245095 -3967 245237
rect -3581 245095 -3547 245237
rect -3161 245095 -3127 245237
rect -2741 245095 -2707 245237
rect -2321 245095 -2287 245237
rect -1901 245095 -1867 245237
rect -1481 245095 -1447 245237
rect -1061 245095 -1027 245237
rect -641 245095 -607 245237
rect -221 245095 -187 245237
rect 199 245095 233 245237
rect 619 245095 653 245237
rect 1039 245095 1073 245237
rect 1459 245095 1493 245237
rect 1879 245095 1913 245237
rect 2299 245095 2333 245237
rect 2719 245095 2753 245237
rect 3139 245095 3173 245237
rect 3559 245095 3593 245237
rect 3979 245095 4013 245237
rect 4399 245095 4433 245237
rect 4819 245095 4853 245237
rect 5239 245095 5273 245237
rect 5659 245095 5693 245237
rect 6079 245095 6113 245237
rect 6499 245095 6533 245237
rect 6919 245095 6953 245237
rect 7339 245095 7373 245237
rect 7759 245095 7793 245237
rect 8179 245095 8213 245237
rect 8599 245095 8633 245237
rect 9019 245095 9053 245237
rect 9439 245095 9473 245237
rect 9859 245095 9893 245237
rect 10279 245095 10313 245237
rect 10699 245095 10733 245237
rect 11119 245095 11153 245237
rect 11539 245095 11573 245237
rect 11959 245095 11993 245237
rect 12379 245095 12413 245237
rect 12799 245095 12833 245237
rect 13219 245095 13253 245237
rect 13639 245095 13673 245237
rect 14059 245095 14093 245237
rect 14479 245095 14513 245237
rect 14899 245095 14933 245237
rect 15319 245095 15353 245237
rect 15739 245095 15773 245237
rect 16159 245095 16193 245237
rect 16579 245095 16613 245237
rect 16999 245095 17033 245237
rect 17419 245095 17453 245237
rect 17839 245095 17873 245237
rect 18259 245095 18293 245237
rect 18679 245095 18713 245237
rect 19099 245095 19133 245237
rect 19519 245095 19553 245237
rect 19939 245095 19973 245237
rect 20359 245095 20393 245237
rect 20779 245095 20813 245237
rect 21199 245095 21233 245237
rect 21619 245095 21653 245237
rect 22039 245095 22073 245237
rect 22459 245095 22493 245237
rect 22879 245095 22913 245237
rect 23299 245095 23333 245237
rect 23719 245095 23753 245237
rect 24139 245095 24173 245237
rect 24559 245095 24593 245237
rect 24979 245095 25013 245237
rect 25399 245095 25433 245237
rect 25819 245095 25853 245237
rect 26239 245095 26273 245237
rect 26659 245095 26693 245237
rect 27079 245095 27113 245237
rect -3791 244167 -3695 244201
rect -3371 244167 -3275 244201
rect -2951 244167 -2855 244201
rect -2531 244167 -2435 244201
rect -2111 244167 -2015 244201
rect -1691 244167 -1595 244201
rect -1271 244167 -1175 244201
rect -851 244167 -755 244201
rect -431 244167 -335 244201
rect -11 244167 85 244201
rect 409 244167 505 244201
rect 829 244167 925 244201
rect 1249 244167 1345 244201
rect 1669 244167 1765 244201
rect 2089 244167 2185 244201
rect 2509 244167 2605 244201
rect 2929 244167 3025 244201
rect 3349 244167 3445 244201
rect 3769 244167 3865 244201
rect 4189 244167 4285 244201
rect 4609 244167 4705 244201
rect 5029 244167 5125 244201
rect 5449 244167 5545 244201
rect 5869 244167 5965 244201
rect 6289 244167 6385 244201
rect 6709 244167 6805 244201
rect 7129 244167 7225 244201
rect 7549 244167 7645 244201
rect 7969 244167 8065 244201
rect 8389 244167 8485 244201
rect 8809 244167 8905 244201
rect 9229 244167 9325 244201
rect 9649 244167 9745 244201
rect 10069 244167 10165 244201
rect 10489 244167 10585 244201
rect 10909 244167 11005 244201
rect 11329 244167 11425 244201
rect 11749 244167 11845 244201
rect 12169 244167 12265 244201
rect 12589 244167 12685 244201
rect 13009 244167 13105 244201
rect 13429 244167 13525 244201
rect 13849 244167 13945 244201
rect 14269 244167 14365 244201
rect 14689 244167 14785 244201
rect 15109 244167 15205 244201
rect 15529 244167 15625 244201
rect 15949 244167 16045 244201
rect 16369 244167 16465 244201
rect 16789 244167 16885 244201
rect 17209 244167 17305 244201
rect 17629 244167 17725 244201
rect 18049 244167 18145 244201
rect 18469 244167 18565 244201
rect 18889 244167 18985 244201
rect 19309 244167 19405 244201
rect 19729 244167 19825 244201
rect 20149 244167 20245 244201
rect 20569 244167 20665 244201
rect 20989 244167 21085 244201
rect 21409 244167 21505 244201
rect 21829 244167 21925 244201
rect 22249 244167 22345 244201
rect 22669 244167 22765 244201
rect 23089 244167 23185 244201
rect 23509 244167 23605 244201
rect 23929 244167 24025 244201
rect 24349 244167 24445 244201
rect 24769 244167 24865 244201
rect 25189 244167 25285 244201
rect 25609 244167 25705 244201
rect 26029 244167 26125 244201
rect 26449 244167 26545 244201
rect 26869 244167 26965 244201
rect 27289 244167 27385 244201
<< locali >>
rect -4163 264178 -4067 264212
rect 27389 264178 27485 264212
rect -4163 264116 -4129 264178
rect 27451 264116 27485 264178
rect -4017 264076 -4001 264110
rect -3905 264076 -3889 264110
rect -3597 264076 -3581 264110
rect -3485 264076 -3469 264110
rect -3177 264076 -3161 264110
rect -3065 264076 -3049 264110
rect -2757 264076 -2741 264110
rect -2645 264076 -2629 264110
rect -2337 264076 -2321 264110
rect -2225 264076 -2209 264110
rect -1917 264076 -1901 264110
rect -1805 264076 -1789 264110
rect -1497 264076 -1481 264110
rect -1385 264076 -1369 264110
rect -1077 264076 -1061 264110
rect -965 264076 -949 264110
rect -657 264076 -641 264110
rect -545 264076 -529 264110
rect -237 264076 -221 264110
rect -125 264076 -109 264110
rect 183 264076 199 264110
rect 295 264076 311 264110
rect 603 264076 619 264110
rect 715 264076 731 264110
rect 1023 264076 1039 264110
rect 1135 264076 1151 264110
rect 1443 264076 1459 264110
rect 1555 264076 1571 264110
rect 1863 264076 1879 264110
rect 1975 264076 1991 264110
rect 2283 264076 2299 264110
rect 2395 264076 2411 264110
rect 2703 264076 2719 264110
rect 2815 264076 2831 264110
rect 3123 264076 3139 264110
rect 3235 264076 3251 264110
rect 3543 264076 3559 264110
rect 3655 264076 3671 264110
rect 3963 264076 3979 264110
rect 4075 264076 4091 264110
rect 4383 264076 4399 264110
rect 4495 264076 4511 264110
rect 4803 264076 4819 264110
rect 4915 264076 4931 264110
rect 5223 264076 5239 264110
rect 5335 264076 5351 264110
rect 5643 264076 5659 264110
rect 5755 264076 5771 264110
rect 6063 264076 6079 264110
rect 6175 264076 6191 264110
rect 6483 264076 6499 264110
rect 6595 264076 6611 264110
rect 6903 264076 6919 264110
rect 7015 264076 7031 264110
rect 7323 264076 7339 264110
rect 7435 264076 7451 264110
rect 7743 264076 7759 264110
rect 7855 264076 7871 264110
rect 8163 264076 8179 264110
rect 8275 264076 8291 264110
rect 8583 264076 8599 264110
rect 8695 264076 8711 264110
rect 9003 264076 9019 264110
rect 9115 264076 9131 264110
rect 9423 264076 9439 264110
rect 9535 264076 9551 264110
rect 9843 264076 9859 264110
rect 9955 264076 9971 264110
rect 10263 264076 10279 264110
rect 10375 264076 10391 264110
rect 10683 264076 10699 264110
rect 10795 264076 10811 264110
rect 11103 264076 11119 264110
rect 11215 264076 11231 264110
rect 11523 264076 11539 264110
rect 11635 264076 11651 264110
rect 11943 264076 11959 264110
rect 12055 264076 12071 264110
rect 12363 264076 12379 264110
rect 12475 264076 12491 264110
rect 12783 264076 12799 264110
rect 12895 264076 12911 264110
rect 13203 264076 13219 264110
rect 13315 264076 13331 264110
rect 13623 264076 13639 264110
rect 13735 264076 13751 264110
rect 14043 264076 14059 264110
rect 14155 264076 14171 264110
rect 14463 264076 14479 264110
rect 14575 264076 14591 264110
rect 14883 264076 14899 264110
rect 14995 264076 15011 264110
rect 15303 264076 15319 264110
rect 15415 264076 15431 264110
rect 15723 264076 15739 264110
rect 15835 264076 15851 264110
rect 16143 264076 16159 264110
rect 16255 264076 16271 264110
rect 16563 264076 16579 264110
rect 16675 264076 16691 264110
rect 16983 264076 16999 264110
rect 17095 264076 17111 264110
rect 17403 264076 17419 264110
rect 17515 264076 17531 264110
rect 17823 264076 17839 264110
rect 17935 264076 17951 264110
rect 18243 264076 18259 264110
rect 18355 264076 18371 264110
rect 18663 264076 18679 264110
rect 18775 264076 18791 264110
rect 19083 264076 19099 264110
rect 19195 264076 19211 264110
rect 19503 264076 19519 264110
rect 19615 264076 19631 264110
rect 19923 264076 19939 264110
rect 20035 264076 20051 264110
rect 20343 264076 20359 264110
rect 20455 264076 20471 264110
rect 20763 264076 20779 264110
rect 20875 264076 20891 264110
rect 21183 264076 21199 264110
rect 21295 264076 21311 264110
rect 21603 264076 21619 264110
rect 21715 264076 21731 264110
rect 22023 264076 22039 264110
rect 22135 264076 22151 264110
rect 22443 264076 22459 264110
rect 22555 264076 22571 264110
rect 22863 264076 22879 264110
rect 22975 264076 22991 264110
rect 23283 264076 23299 264110
rect 23395 264076 23411 264110
rect 23703 264076 23719 264110
rect 23815 264076 23831 264110
rect 24123 264076 24139 264110
rect 24235 264076 24251 264110
rect 24543 264076 24559 264110
rect 24655 264076 24671 264110
rect 24963 264076 24979 264110
rect 25075 264076 25091 264110
rect 25383 264076 25399 264110
rect 25495 264076 25511 264110
rect 25803 264076 25819 264110
rect 25915 264076 25931 264110
rect 26223 264076 26239 264110
rect 26335 264076 26351 264110
rect 26643 264076 26659 264110
rect 26755 264076 26771 264110
rect 27063 264076 27079 264110
rect 27175 264076 27191 264110
rect -4049 264026 -4015 264042
rect -4049 263234 -4015 263250
rect -3953 264026 -3919 264042
rect -3953 263234 -3919 263250
rect -3839 264026 -3805 264042
rect -3839 263234 -3805 263250
rect -3743 264026 -3709 264042
rect -3743 263234 -3709 263250
rect -3629 264026 -3595 264042
rect -3629 263234 -3595 263250
rect -3533 264026 -3499 264042
rect -3533 263234 -3499 263250
rect -3419 264026 -3385 264042
rect -3419 263234 -3385 263250
rect -3323 264026 -3289 264042
rect -3323 263234 -3289 263250
rect -3209 264026 -3175 264042
rect -3209 263234 -3175 263250
rect -3113 264026 -3079 264042
rect -3113 263234 -3079 263250
rect -2999 264026 -2965 264042
rect -2999 263234 -2965 263250
rect -2903 264026 -2869 264042
rect -2903 263234 -2869 263250
rect -2789 264026 -2755 264042
rect -2789 263234 -2755 263250
rect -2693 264026 -2659 264042
rect -2693 263234 -2659 263250
rect -2579 264026 -2545 264042
rect -2579 263234 -2545 263250
rect -2483 264026 -2449 264042
rect -2483 263234 -2449 263250
rect -2369 264026 -2335 264042
rect -2369 263234 -2335 263250
rect -2273 264026 -2239 264042
rect -2273 263234 -2239 263250
rect -2159 264026 -2125 264042
rect -2159 263234 -2125 263250
rect -2063 264026 -2029 264042
rect -2063 263234 -2029 263250
rect -1949 264026 -1915 264042
rect -1949 263234 -1915 263250
rect -1853 264026 -1819 264042
rect -1853 263234 -1819 263250
rect -1739 264026 -1705 264042
rect -1739 263234 -1705 263250
rect -1643 264026 -1609 264042
rect -1643 263234 -1609 263250
rect -1529 264026 -1495 264042
rect -1529 263234 -1495 263250
rect -1433 264026 -1399 264042
rect -1433 263234 -1399 263250
rect -1319 264026 -1285 264042
rect -1319 263234 -1285 263250
rect -1223 264026 -1189 264042
rect -1223 263234 -1189 263250
rect -1109 264026 -1075 264042
rect -1109 263234 -1075 263250
rect -1013 264026 -979 264042
rect -1013 263234 -979 263250
rect -899 264026 -865 264042
rect -899 263234 -865 263250
rect -803 264026 -769 264042
rect -803 263234 -769 263250
rect -689 264026 -655 264042
rect -689 263234 -655 263250
rect -593 264026 -559 264042
rect -593 263234 -559 263250
rect -479 264026 -445 264042
rect -479 263234 -445 263250
rect -383 264026 -349 264042
rect -383 263234 -349 263250
rect -269 264026 -235 264042
rect -269 263234 -235 263250
rect -173 264026 -139 264042
rect -173 263234 -139 263250
rect -59 264026 -25 264042
rect -59 263234 -25 263250
rect 37 264026 71 264042
rect 37 263234 71 263250
rect 151 264026 185 264042
rect 151 263234 185 263250
rect 247 264026 281 264042
rect 247 263234 281 263250
rect 361 264026 395 264042
rect 361 263234 395 263250
rect 457 264026 491 264042
rect 457 263234 491 263250
rect 571 264026 605 264042
rect 571 263234 605 263250
rect 667 264026 701 264042
rect 667 263234 701 263250
rect 781 264026 815 264042
rect 781 263234 815 263250
rect 877 264026 911 264042
rect 877 263234 911 263250
rect 991 264026 1025 264042
rect 991 263234 1025 263250
rect 1087 264026 1121 264042
rect 1087 263234 1121 263250
rect 1201 264026 1235 264042
rect 1201 263234 1235 263250
rect 1297 264026 1331 264042
rect 1297 263234 1331 263250
rect 1411 264026 1445 264042
rect 1411 263234 1445 263250
rect 1507 264026 1541 264042
rect 1507 263234 1541 263250
rect 1621 264026 1655 264042
rect 1621 263234 1655 263250
rect 1717 264026 1751 264042
rect 1717 263234 1751 263250
rect 1831 264026 1865 264042
rect 1831 263234 1865 263250
rect 1927 264026 1961 264042
rect 1927 263234 1961 263250
rect 2041 264026 2075 264042
rect 2041 263234 2075 263250
rect 2137 264026 2171 264042
rect 2137 263234 2171 263250
rect 2251 264026 2285 264042
rect 2251 263234 2285 263250
rect 2347 264026 2381 264042
rect 2347 263234 2381 263250
rect 2461 264026 2495 264042
rect 2461 263234 2495 263250
rect 2557 264026 2591 264042
rect 2557 263234 2591 263250
rect 2671 264026 2705 264042
rect 2671 263234 2705 263250
rect 2767 264026 2801 264042
rect 2767 263234 2801 263250
rect 2881 264026 2915 264042
rect 2881 263234 2915 263250
rect 2977 264026 3011 264042
rect 2977 263234 3011 263250
rect 3091 264026 3125 264042
rect 3091 263234 3125 263250
rect 3187 264026 3221 264042
rect 3187 263234 3221 263250
rect 3301 264026 3335 264042
rect 3301 263234 3335 263250
rect 3397 264026 3431 264042
rect 3397 263234 3431 263250
rect 3511 264026 3545 264042
rect 3511 263234 3545 263250
rect 3607 264026 3641 264042
rect 3607 263234 3641 263250
rect 3721 264026 3755 264042
rect 3721 263234 3755 263250
rect 3817 264026 3851 264042
rect 3817 263234 3851 263250
rect 3931 264026 3965 264042
rect 3931 263234 3965 263250
rect 4027 264026 4061 264042
rect 4027 263234 4061 263250
rect 4141 264026 4175 264042
rect 4141 263234 4175 263250
rect 4237 264026 4271 264042
rect 4237 263234 4271 263250
rect 4351 264026 4385 264042
rect 4351 263234 4385 263250
rect 4447 264026 4481 264042
rect 4447 263234 4481 263250
rect 4561 264026 4595 264042
rect 4561 263234 4595 263250
rect 4657 264026 4691 264042
rect 4657 263234 4691 263250
rect 4771 264026 4805 264042
rect 4771 263234 4805 263250
rect 4867 264026 4901 264042
rect 4867 263234 4901 263250
rect 4981 264026 5015 264042
rect 4981 263234 5015 263250
rect 5077 264026 5111 264042
rect 5077 263234 5111 263250
rect 5191 264026 5225 264042
rect 5191 263234 5225 263250
rect 5287 264026 5321 264042
rect 5287 263234 5321 263250
rect 5401 264026 5435 264042
rect 5401 263234 5435 263250
rect 5497 264026 5531 264042
rect 5497 263234 5531 263250
rect 5611 264026 5645 264042
rect 5611 263234 5645 263250
rect 5707 264026 5741 264042
rect 5707 263234 5741 263250
rect 5821 264026 5855 264042
rect 5821 263234 5855 263250
rect 5917 264026 5951 264042
rect 5917 263234 5951 263250
rect 6031 264026 6065 264042
rect 6031 263234 6065 263250
rect 6127 264026 6161 264042
rect 6127 263234 6161 263250
rect 6241 264026 6275 264042
rect 6241 263234 6275 263250
rect 6337 264026 6371 264042
rect 6337 263234 6371 263250
rect 6451 264026 6485 264042
rect 6451 263234 6485 263250
rect 6547 264026 6581 264042
rect 6547 263234 6581 263250
rect 6661 264026 6695 264042
rect 6661 263234 6695 263250
rect 6757 264026 6791 264042
rect 6757 263234 6791 263250
rect 6871 264026 6905 264042
rect 6871 263234 6905 263250
rect 6967 264026 7001 264042
rect 6967 263234 7001 263250
rect 7081 264026 7115 264042
rect 7081 263234 7115 263250
rect 7177 264026 7211 264042
rect 7177 263234 7211 263250
rect 7291 264026 7325 264042
rect 7291 263234 7325 263250
rect 7387 264026 7421 264042
rect 7387 263234 7421 263250
rect 7501 264026 7535 264042
rect 7501 263234 7535 263250
rect 7597 264026 7631 264042
rect 7597 263234 7631 263250
rect 7711 264026 7745 264042
rect 7711 263234 7745 263250
rect 7807 264026 7841 264042
rect 7807 263234 7841 263250
rect 7921 264026 7955 264042
rect 7921 263234 7955 263250
rect 8017 264026 8051 264042
rect 8017 263234 8051 263250
rect 8131 264026 8165 264042
rect 8131 263234 8165 263250
rect 8227 264026 8261 264042
rect 8227 263234 8261 263250
rect 8341 264026 8375 264042
rect 8341 263234 8375 263250
rect 8437 264026 8471 264042
rect 8437 263234 8471 263250
rect 8551 264026 8585 264042
rect 8551 263234 8585 263250
rect 8647 264026 8681 264042
rect 8647 263234 8681 263250
rect 8761 264026 8795 264042
rect 8761 263234 8795 263250
rect 8857 264026 8891 264042
rect 8857 263234 8891 263250
rect 8971 264026 9005 264042
rect 8971 263234 9005 263250
rect 9067 264026 9101 264042
rect 9067 263234 9101 263250
rect 9181 264026 9215 264042
rect 9181 263234 9215 263250
rect 9277 264026 9311 264042
rect 9277 263234 9311 263250
rect 9391 264026 9425 264042
rect 9391 263234 9425 263250
rect 9487 264026 9521 264042
rect 9487 263234 9521 263250
rect 9601 264026 9635 264042
rect 9601 263234 9635 263250
rect 9697 264026 9731 264042
rect 9697 263234 9731 263250
rect 9811 264026 9845 264042
rect 9811 263234 9845 263250
rect 9907 264026 9941 264042
rect 9907 263234 9941 263250
rect 10021 264026 10055 264042
rect 10021 263234 10055 263250
rect 10117 264026 10151 264042
rect 10117 263234 10151 263250
rect 10231 264026 10265 264042
rect 10231 263234 10265 263250
rect 10327 264026 10361 264042
rect 10327 263234 10361 263250
rect 10441 264026 10475 264042
rect 10441 263234 10475 263250
rect 10537 264026 10571 264042
rect 10537 263234 10571 263250
rect 10651 264026 10685 264042
rect 10651 263234 10685 263250
rect 10747 264026 10781 264042
rect 10747 263234 10781 263250
rect 10861 264026 10895 264042
rect 10861 263234 10895 263250
rect 10957 264026 10991 264042
rect 10957 263234 10991 263250
rect 11071 264026 11105 264042
rect 11071 263234 11105 263250
rect 11167 264026 11201 264042
rect 11167 263234 11201 263250
rect 11281 264026 11315 264042
rect 11281 263234 11315 263250
rect 11377 264026 11411 264042
rect 11377 263234 11411 263250
rect 11491 264026 11525 264042
rect 11491 263234 11525 263250
rect 11587 264026 11621 264042
rect 11587 263234 11621 263250
rect 11701 264026 11735 264042
rect 11701 263234 11735 263250
rect 11797 264026 11831 264042
rect 11797 263234 11831 263250
rect 11911 264026 11945 264042
rect 11911 263234 11945 263250
rect 12007 264026 12041 264042
rect 12007 263234 12041 263250
rect 12121 264026 12155 264042
rect 12121 263234 12155 263250
rect 12217 264026 12251 264042
rect 12217 263234 12251 263250
rect 12331 264026 12365 264042
rect 12331 263234 12365 263250
rect 12427 264026 12461 264042
rect 12427 263234 12461 263250
rect 12541 264026 12575 264042
rect 12541 263234 12575 263250
rect 12637 264026 12671 264042
rect 12637 263234 12671 263250
rect 12751 264026 12785 264042
rect 12751 263234 12785 263250
rect 12847 264026 12881 264042
rect 12847 263234 12881 263250
rect 12961 264026 12995 264042
rect 12961 263234 12995 263250
rect 13057 264026 13091 264042
rect 13057 263234 13091 263250
rect 13171 264026 13205 264042
rect 13171 263234 13205 263250
rect 13267 264026 13301 264042
rect 13267 263234 13301 263250
rect 13381 264026 13415 264042
rect 13381 263234 13415 263250
rect 13477 264026 13511 264042
rect 13477 263234 13511 263250
rect 13591 264026 13625 264042
rect 13591 263234 13625 263250
rect 13687 264026 13721 264042
rect 13687 263234 13721 263250
rect 13801 264026 13835 264042
rect 13801 263234 13835 263250
rect 13897 264026 13931 264042
rect 13897 263234 13931 263250
rect 14011 264026 14045 264042
rect 14011 263234 14045 263250
rect 14107 264026 14141 264042
rect 14107 263234 14141 263250
rect 14221 264026 14255 264042
rect 14221 263234 14255 263250
rect 14317 264026 14351 264042
rect 14317 263234 14351 263250
rect 14431 264026 14465 264042
rect 14431 263234 14465 263250
rect 14527 264026 14561 264042
rect 14527 263234 14561 263250
rect 14641 264026 14675 264042
rect 14641 263234 14675 263250
rect 14737 264026 14771 264042
rect 14737 263234 14771 263250
rect 14851 264026 14885 264042
rect 14851 263234 14885 263250
rect 14947 264026 14981 264042
rect 14947 263234 14981 263250
rect 15061 264026 15095 264042
rect 15061 263234 15095 263250
rect 15157 264026 15191 264042
rect 15157 263234 15191 263250
rect 15271 264026 15305 264042
rect 15271 263234 15305 263250
rect 15367 264026 15401 264042
rect 15367 263234 15401 263250
rect 15481 264026 15515 264042
rect 15481 263234 15515 263250
rect 15577 264026 15611 264042
rect 15577 263234 15611 263250
rect 15691 264026 15725 264042
rect 15691 263234 15725 263250
rect 15787 264026 15821 264042
rect 15787 263234 15821 263250
rect 15901 264026 15935 264042
rect 15901 263234 15935 263250
rect 15997 264026 16031 264042
rect 15997 263234 16031 263250
rect 16111 264026 16145 264042
rect 16111 263234 16145 263250
rect 16207 264026 16241 264042
rect 16207 263234 16241 263250
rect 16321 264026 16355 264042
rect 16321 263234 16355 263250
rect 16417 264026 16451 264042
rect 16417 263234 16451 263250
rect 16531 264026 16565 264042
rect 16531 263234 16565 263250
rect 16627 264026 16661 264042
rect 16627 263234 16661 263250
rect 16741 264026 16775 264042
rect 16741 263234 16775 263250
rect 16837 264026 16871 264042
rect 16837 263234 16871 263250
rect 16951 264026 16985 264042
rect 16951 263234 16985 263250
rect 17047 264026 17081 264042
rect 17047 263234 17081 263250
rect 17161 264026 17195 264042
rect 17161 263234 17195 263250
rect 17257 264026 17291 264042
rect 17257 263234 17291 263250
rect 17371 264026 17405 264042
rect 17371 263234 17405 263250
rect 17467 264026 17501 264042
rect 17467 263234 17501 263250
rect 17581 264026 17615 264042
rect 17581 263234 17615 263250
rect 17677 264026 17711 264042
rect 17677 263234 17711 263250
rect 17791 264026 17825 264042
rect 17791 263234 17825 263250
rect 17887 264026 17921 264042
rect 17887 263234 17921 263250
rect 18001 264026 18035 264042
rect 18001 263234 18035 263250
rect 18097 264026 18131 264042
rect 18097 263234 18131 263250
rect 18211 264026 18245 264042
rect 18211 263234 18245 263250
rect 18307 264026 18341 264042
rect 18307 263234 18341 263250
rect 18421 264026 18455 264042
rect 18421 263234 18455 263250
rect 18517 264026 18551 264042
rect 18517 263234 18551 263250
rect 18631 264026 18665 264042
rect 18631 263234 18665 263250
rect 18727 264026 18761 264042
rect 18727 263234 18761 263250
rect 18841 264026 18875 264042
rect 18841 263234 18875 263250
rect 18937 264026 18971 264042
rect 18937 263234 18971 263250
rect 19051 264026 19085 264042
rect 19051 263234 19085 263250
rect 19147 264026 19181 264042
rect 19147 263234 19181 263250
rect 19261 264026 19295 264042
rect 19261 263234 19295 263250
rect 19357 264026 19391 264042
rect 19357 263234 19391 263250
rect 19471 264026 19505 264042
rect 19471 263234 19505 263250
rect 19567 264026 19601 264042
rect 19567 263234 19601 263250
rect 19681 264026 19715 264042
rect 19681 263234 19715 263250
rect 19777 264026 19811 264042
rect 19777 263234 19811 263250
rect 19891 264026 19925 264042
rect 19891 263234 19925 263250
rect 19987 264026 20021 264042
rect 19987 263234 20021 263250
rect 20101 264026 20135 264042
rect 20101 263234 20135 263250
rect 20197 264026 20231 264042
rect 20197 263234 20231 263250
rect 20311 264026 20345 264042
rect 20311 263234 20345 263250
rect 20407 264026 20441 264042
rect 20407 263234 20441 263250
rect 20521 264026 20555 264042
rect 20521 263234 20555 263250
rect 20617 264026 20651 264042
rect 20617 263234 20651 263250
rect 20731 264026 20765 264042
rect 20731 263234 20765 263250
rect 20827 264026 20861 264042
rect 20827 263234 20861 263250
rect 20941 264026 20975 264042
rect 20941 263234 20975 263250
rect 21037 264026 21071 264042
rect 21037 263234 21071 263250
rect 21151 264026 21185 264042
rect 21151 263234 21185 263250
rect 21247 264026 21281 264042
rect 21247 263234 21281 263250
rect 21361 264026 21395 264042
rect 21361 263234 21395 263250
rect 21457 264026 21491 264042
rect 21457 263234 21491 263250
rect 21571 264026 21605 264042
rect 21571 263234 21605 263250
rect 21667 264026 21701 264042
rect 21667 263234 21701 263250
rect 21781 264026 21815 264042
rect 21781 263234 21815 263250
rect 21877 264026 21911 264042
rect 21877 263234 21911 263250
rect 21991 264026 22025 264042
rect 21991 263234 22025 263250
rect 22087 264026 22121 264042
rect 22087 263234 22121 263250
rect 22201 264026 22235 264042
rect 22201 263234 22235 263250
rect 22297 264026 22331 264042
rect 22297 263234 22331 263250
rect 22411 264026 22445 264042
rect 22411 263234 22445 263250
rect 22507 264026 22541 264042
rect 22507 263234 22541 263250
rect 22621 264026 22655 264042
rect 22621 263234 22655 263250
rect 22717 264026 22751 264042
rect 22717 263234 22751 263250
rect 22831 264026 22865 264042
rect 22831 263234 22865 263250
rect 22927 264026 22961 264042
rect 22927 263234 22961 263250
rect 23041 264026 23075 264042
rect 23041 263234 23075 263250
rect 23137 264026 23171 264042
rect 23137 263234 23171 263250
rect 23251 264026 23285 264042
rect 23251 263234 23285 263250
rect 23347 264026 23381 264042
rect 23347 263234 23381 263250
rect 23461 264026 23495 264042
rect 23461 263234 23495 263250
rect 23557 264026 23591 264042
rect 23557 263234 23591 263250
rect 23671 264026 23705 264042
rect 23671 263234 23705 263250
rect 23767 264026 23801 264042
rect 23767 263234 23801 263250
rect 23881 264026 23915 264042
rect 23881 263234 23915 263250
rect 23977 264026 24011 264042
rect 23977 263234 24011 263250
rect 24091 264026 24125 264042
rect 24091 263234 24125 263250
rect 24187 264026 24221 264042
rect 24187 263234 24221 263250
rect 24301 264026 24335 264042
rect 24301 263234 24335 263250
rect 24397 264026 24431 264042
rect 24397 263234 24431 263250
rect 24511 264026 24545 264042
rect 24511 263234 24545 263250
rect 24607 264026 24641 264042
rect 24607 263234 24641 263250
rect 24721 264026 24755 264042
rect 24721 263234 24755 263250
rect 24817 264026 24851 264042
rect 24817 263234 24851 263250
rect 24931 264026 24965 264042
rect 24931 263234 24965 263250
rect 25027 264026 25061 264042
rect 25027 263234 25061 263250
rect 25141 264026 25175 264042
rect 25141 263234 25175 263250
rect 25237 264026 25271 264042
rect 25237 263234 25271 263250
rect 25351 264026 25385 264042
rect 25351 263234 25385 263250
rect 25447 264026 25481 264042
rect 25447 263234 25481 263250
rect 25561 264026 25595 264042
rect 25561 263234 25595 263250
rect 25657 264026 25691 264042
rect 25657 263234 25691 263250
rect 25771 264026 25805 264042
rect 25771 263234 25805 263250
rect 25867 264026 25901 264042
rect 25867 263234 25901 263250
rect 25981 264026 26015 264042
rect 25981 263234 26015 263250
rect 26077 264026 26111 264042
rect 26077 263234 26111 263250
rect 26191 264026 26225 264042
rect 26191 263234 26225 263250
rect 26287 264026 26321 264042
rect 26287 263234 26321 263250
rect 26401 264026 26435 264042
rect 26401 263234 26435 263250
rect 26497 264026 26531 264042
rect 26497 263234 26531 263250
rect 26611 264026 26645 264042
rect 26611 263234 26645 263250
rect 26707 264026 26741 264042
rect 26707 263234 26741 263250
rect 26821 264026 26855 264042
rect 26821 263234 26855 263250
rect 26917 264026 26951 264042
rect 26917 263234 26951 263250
rect 27031 264026 27065 264042
rect 27031 263234 27065 263250
rect 27127 264026 27161 264042
rect 27127 263234 27161 263250
rect 27241 264026 27275 264042
rect 27241 263234 27275 263250
rect 27337 264026 27371 264042
rect 27337 263234 27371 263250
rect -3807 263164 -3791 263198
rect -3757 263164 -3741 263198
rect -3387 263164 -3371 263198
rect -3337 263164 -3321 263198
rect -2967 263164 -2951 263198
rect -2917 263164 -2901 263198
rect -2547 263164 -2531 263198
rect -2497 263164 -2481 263198
rect -2127 263164 -2111 263198
rect -2077 263164 -2061 263198
rect -1707 263164 -1691 263198
rect -1657 263164 -1641 263198
rect -1287 263164 -1271 263198
rect -1237 263164 -1221 263198
rect -867 263164 -851 263198
rect -817 263164 -801 263198
rect -447 263164 -431 263198
rect -397 263164 -381 263198
rect -27 263164 -11 263198
rect 23 263164 39 263198
rect 393 263164 409 263198
rect 443 263164 459 263198
rect 813 263164 829 263198
rect 863 263164 879 263198
rect 1233 263164 1249 263198
rect 1283 263164 1299 263198
rect 1653 263164 1669 263198
rect 1703 263164 1719 263198
rect 2073 263164 2089 263198
rect 2123 263164 2139 263198
rect 2493 263164 2509 263198
rect 2543 263164 2559 263198
rect 2913 263164 2929 263198
rect 2963 263164 2979 263198
rect 3333 263164 3349 263198
rect 3383 263164 3399 263198
rect 3753 263164 3769 263198
rect 3803 263164 3819 263198
rect 4173 263164 4189 263198
rect 4223 263164 4239 263198
rect 4593 263164 4609 263198
rect 4643 263164 4659 263198
rect 5013 263164 5029 263198
rect 5063 263164 5079 263198
rect 5433 263164 5449 263198
rect 5483 263164 5499 263198
rect 5853 263164 5869 263198
rect 5903 263164 5919 263198
rect 6273 263164 6289 263198
rect 6323 263164 6339 263198
rect 6693 263164 6709 263198
rect 6743 263164 6759 263198
rect 7113 263164 7129 263198
rect 7163 263164 7179 263198
rect 7533 263164 7549 263198
rect 7583 263164 7599 263198
rect 7953 263164 7969 263198
rect 8003 263164 8019 263198
rect 8373 263164 8389 263198
rect 8423 263164 8439 263198
rect 8793 263164 8809 263198
rect 8843 263164 8859 263198
rect 9213 263164 9229 263198
rect 9263 263164 9279 263198
rect 9633 263164 9649 263198
rect 9683 263164 9699 263198
rect 10053 263164 10069 263198
rect 10103 263164 10119 263198
rect 10473 263164 10489 263198
rect 10523 263164 10539 263198
rect 10893 263164 10909 263198
rect 10943 263164 10959 263198
rect 11313 263164 11329 263198
rect 11363 263164 11379 263198
rect 11733 263164 11749 263198
rect 11783 263164 11799 263198
rect 12153 263164 12169 263198
rect 12203 263164 12219 263198
rect 12573 263164 12589 263198
rect 12623 263164 12639 263198
rect 12993 263164 13009 263198
rect 13043 263164 13059 263198
rect 13413 263164 13429 263198
rect 13463 263164 13479 263198
rect 13833 263164 13849 263198
rect 13883 263164 13899 263198
rect 14253 263164 14269 263198
rect 14303 263164 14319 263198
rect 14673 263164 14689 263198
rect 14723 263164 14739 263198
rect 15093 263164 15109 263198
rect 15143 263164 15159 263198
rect 15513 263164 15529 263198
rect 15563 263164 15579 263198
rect 15933 263164 15949 263198
rect 15983 263164 15999 263198
rect 16353 263164 16369 263198
rect 16403 263164 16419 263198
rect 16773 263164 16789 263198
rect 16823 263164 16839 263198
rect 17193 263164 17209 263198
rect 17243 263164 17259 263198
rect 17613 263164 17629 263198
rect 17663 263164 17679 263198
rect 18033 263164 18049 263198
rect 18083 263164 18099 263198
rect 18453 263164 18469 263198
rect 18503 263164 18519 263198
rect 18873 263164 18889 263198
rect 18923 263164 18939 263198
rect 19293 263164 19309 263198
rect 19343 263164 19359 263198
rect 19713 263164 19729 263198
rect 19763 263164 19779 263198
rect 20133 263164 20149 263198
rect 20183 263164 20199 263198
rect 20553 263164 20569 263198
rect 20603 263164 20619 263198
rect 20973 263164 20989 263198
rect 21023 263164 21039 263198
rect 21393 263164 21409 263198
rect 21443 263164 21459 263198
rect 21813 263164 21829 263198
rect 21863 263164 21879 263198
rect 22233 263164 22249 263198
rect 22283 263164 22299 263198
rect 22653 263164 22669 263198
rect 22703 263164 22719 263198
rect 23073 263164 23089 263198
rect 23123 263164 23139 263198
rect 23493 263164 23509 263198
rect 23543 263164 23559 263198
rect 23913 263164 23929 263198
rect 23963 263164 23979 263198
rect 24333 263164 24349 263198
rect 24383 263164 24399 263198
rect 24753 263164 24769 263198
rect 24803 263164 24819 263198
rect 25173 263164 25189 263198
rect 25223 263164 25239 263198
rect 25593 263164 25609 263198
rect 25643 263164 25659 263198
rect 26013 263164 26029 263198
rect 26063 263164 26079 263198
rect 26433 263164 26449 263198
rect 26483 263164 26499 263198
rect 26853 263164 26869 263198
rect 26903 263164 26919 263198
rect 27273 263164 27289 263198
rect 27323 263164 27339 263198
rect -3807 263056 -3791 263090
rect -3757 263056 -3741 263090
rect -3387 263056 -3371 263090
rect -3337 263056 -3321 263090
rect -2967 263056 -2951 263090
rect -2917 263056 -2901 263090
rect -2547 263056 -2531 263090
rect -2497 263056 -2481 263090
rect -2127 263056 -2111 263090
rect -2077 263056 -2061 263090
rect -1707 263056 -1691 263090
rect -1657 263056 -1641 263090
rect -1287 263056 -1271 263090
rect -1237 263056 -1221 263090
rect -867 263056 -851 263090
rect -817 263056 -801 263090
rect -447 263056 -431 263090
rect -397 263056 -381 263090
rect -27 263056 -11 263090
rect 23 263056 39 263090
rect 393 263056 409 263090
rect 443 263056 459 263090
rect 813 263056 829 263090
rect 863 263056 879 263090
rect 1233 263056 1249 263090
rect 1283 263056 1299 263090
rect 1653 263056 1669 263090
rect 1703 263056 1719 263090
rect 2073 263056 2089 263090
rect 2123 263056 2139 263090
rect 2493 263056 2509 263090
rect 2543 263056 2559 263090
rect 2913 263056 2929 263090
rect 2963 263056 2979 263090
rect 3333 263056 3349 263090
rect 3383 263056 3399 263090
rect 3753 263056 3769 263090
rect 3803 263056 3819 263090
rect 4173 263056 4189 263090
rect 4223 263056 4239 263090
rect 4593 263056 4609 263090
rect 4643 263056 4659 263090
rect 5013 263056 5029 263090
rect 5063 263056 5079 263090
rect 5433 263056 5449 263090
rect 5483 263056 5499 263090
rect 5853 263056 5869 263090
rect 5903 263056 5919 263090
rect 6273 263056 6289 263090
rect 6323 263056 6339 263090
rect 6693 263056 6709 263090
rect 6743 263056 6759 263090
rect 7113 263056 7129 263090
rect 7163 263056 7179 263090
rect 7533 263056 7549 263090
rect 7583 263056 7599 263090
rect 7953 263056 7969 263090
rect 8003 263056 8019 263090
rect 8373 263056 8389 263090
rect 8423 263056 8439 263090
rect 8793 263056 8809 263090
rect 8843 263056 8859 263090
rect 9213 263056 9229 263090
rect 9263 263056 9279 263090
rect 9633 263056 9649 263090
rect 9683 263056 9699 263090
rect 10053 263056 10069 263090
rect 10103 263056 10119 263090
rect 10473 263056 10489 263090
rect 10523 263056 10539 263090
rect 10893 263056 10909 263090
rect 10943 263056 10959 263090
rect 11313 263056 11329 263090
rect 11363 263056 11379 263090
rect 11733 263056 11749 263090
rect 11783 263056 11799 263090
rect 12153 263056 12169 263090
rect 12203 263056 12219 263090
rect 12573 263056 12589 263090
rect 12623 263056 12639 263090
rect 12993 263056 13009 263090
rect 13043 263056 13059 263090
rect 13413 263056 13429 263090
rect 13463 263056 13479 263090
rect 13833 263056 13849 263090
rect 13883 263056 13899 263090
rect 14253 263056 14269 263090
rect 14303 263056 14319 263090
rect 14673 263056 14689 263090
rect 14723 263056 14739 263090
rect 15093 263056 15109 263090
rect 15143 263056 15159 263090
rect 15513 263056 15529 263090
rect 15563 263056 15579 263090
rect 15933 263056 15949 263090
rect 15983 263056 15999 263090
rect 16353 263056 16369 263090
rect 16403 263056 16419 263090
rect 16773 263056 16789 263090
rect 16823 263056 16839 263090
rect 17193 263056 17209 263090
rect 17243 263056 17259 263090
rect 17613 263056 17629 263090
rect 17663 263056 17679 263090
rect 18033 263056 18049 263090
rect 18083 263056 18099 263090
rect 18453 263056 18469 263090
rect 18503 263056 18519 263090
rect 18873 263056 18889 263090
rect 18923 263056 18939 263090
rect 19293 263056 19309 263090
rect 19343 263056 19359 263090
rect 19713 263056 19729 263090
rect 19763 263056 19779 263090
rect 20133 263056 20149 263090
rect 20183 263056 20199 263090
rect 20553 263056 20569 263090
rect 20603 263056 20619 263090
rect 20973 263056 20989 263090
rect 21023 263056 21039 263090
rect 21393 263056 21409 263090
rect 21443 263056 21459 263090
rect 21813 263056 21829 263090
rect 21863 263056 21879 263090
rect 22233 263056 22249 263090
rect 22283 263056 22299 263090
rect 22653 263056 22669 263090
rect 22703 263056 22719 263090
rect 23073 263056 23089 263090
rect 23123 263056 23139 263090
rect 23493 263056 23509 263090
rect 23543 263056 23559 263090
rect 23913 263056 23929 263090
rect 23963 263056 23979 263090
rect 24333 263056 24349 263090
rect 24383 263056 24399 263090
rect 24753 263056 24769 263090
rect 24803 263056 24819 263090
rect 25173 263056 25189 263090
rect 25223 263056 25239 263090
rect 25593 263056 25609 263090
rect 25643 263056 25659 263090
rect 26013 263056 26029 263090
rect 26063 263056 26079 263090
rect 26433 263056 26449 263090
rect 26483 263056 26499 263090
rect 26853 263056 26869 263090
rect 26903 263056 26919 263090
rect 27273 263056 27289 263090
rect 27323 263056 27339 263090
rect -4049 263004 -4015 263020
rect -4049 262212 -4015 262228
rect -3953 263004 -3919 263020
rect -3953 262212 -3919 262228
rect -3839 263004 -3805 263020
rect -3839 262212 -3805 262228
rect -3743 263004 -3709 263020
rect -3743 262212 -3709 262228
rect -3629 263004 -3595 263020
rect -3629 262212 -3595 262228
rect -3533 263004 -3499 263020
rect -3533 262212 -3499 262228
rect -3419 263004 -3385 263020
rect -3419 262212 -3385 262228
rect -3323 263004 -3289 263020
rect -3323 262212 -3289 262228
rect -3209 263004 -3175 263020
rect -3209 262212 -3175 262228
rect -3113 263004 -3079 263020
rect -3113 262212 -3079 262228
rect -2999 263004 -2965 263020
rect -2999 262212 -2965 262228
rect -2903 263004 -2869 263020
rect -2903 262212 -2869 262228
rect -2789 263004 -2755 263020
rect -2789 262212 -2755 262228
rect -2693 263004 -2659 263020
rect -2693 262212 -2659 262228
rect -2579 263004 -2545 263020
rect -2579 262212 -2545 262228
rect -2483 263004 -2449 263020
rect -2483 262212 -2449 262228
rect -2369 263004 -2335 263020
rect -2369 262212 -2335 262228
rect -2273 263004 -2239 263020
rect -2273 262212 -2239 262228
rect -2159 263004 -2125 263020
rect -2159 262212 -2125 262228
rect -2063 263004 -2029 263020
rect -2063 262212 -2029 262228
rect -1949 263004 -1915 263020
rect -1949 262212 -1915 262228
rect -1853 263004 -1819 263020
rect -1853 262212 -1819 262228
rect -1739 263004 -1705 263020
rect -1739 262212 -1705 262228
rect -1643 263004 -1609 263020
rect -1643 262212 -1609 262228
rect -1529 263004 -1495 263020
rect -1529 262212 -1495 262228
rect -1433 263004 -1399 263020
rect -1433 262212 -1399 262228
rect -1319 263004 -1285 263020
rect -1319 262212 -1285 262228
rect -1223 263004 -1189 263020
rect -1223 262212 -1189 262228
rect -1109 263004 -1075 263020
rect -1109 262212 -1075 262228
rect -1013 263004 -979 263020
rect -1013 262212 -979 262228
rect -899 263004 -865 263020
rect -899 262212 -865 262228
rect -803 263004 -769 263020
rect -803 262212 -769 262228
rect -689 263004 -655 263020
rect -689 262212 -655 262228
rect -593 263004 -559 263020
rect -593 262212 -559 262228
rect -479 263004 -445 263020
rect -479 262212 -445 262228
rect -383 263004 -349 263020
rect -383 262212 -349 262228
rect -269 263004 -235 263020
rect -269 262212 -235 262228
rect -173 263004 -139 263020
rect -173 262212 -139 262228
rect -59 263004 -25 263020
rect -59 262212 -25 262228
rect 37 263004 71 263020
rect 37 262212 71 262228
rect 151 263004 185 263020
rect 151 262212 185 262228
rect 247 263004 281 263020
rect 247 262212 281 262228
rect 361 263004 395 263020
rect 361 262212 395 262228
rect 457 263004 491 263020
rect 457 262212 491 262228
rect 571 263004 605 263020
rect 571 262212 605 262228
rect 667 263004 701 263020
rect 667 262212 701 262228
rect 781 263004 815 263020
rect 781 262212 815 262228
rect 877 263004 911 263020
rect 877 262212 911 262228
rect 991 263004 1025 263020
rect 991 262212 1025 262228
rect 1087 263004 1121 263020
rect 1087 262212 1121 262228
rect 1201 263004 1235 263020
rect 1201 262212 1235 262228
rect 1297 263004 1331 263020
rect 1297 262212 1331 262228
rect 1411 263004 1445 263020
rect 1411 262212 1445 262228
rect 1507 263004 1541 263020
rect 1507 262212 1541 262228
rect 1621 263004 1655 263020
rect 1621 262212 1655 262228
rect 1717 263004 1751 263020
rect 1717 262212 1751 262228
rect 1831 263004 1865 263020
rect 1831 262212 1865 262228
rect 1927 263004 1961 263020
rect 1927 262212 1961 262228
rect 2041 263004 2075 263020
rect 2041 262212 2075 262228
rect 2137 263004 2171 263020
rect 2137 262212 2171 262228
rect 2251 263004 2285 263020
rect 2251 262212 2285 262228
rect 2347 263004 2381 263020
rect 2347 262212 2381 262228
rect 2461 263004 2495 263020
rect 2461 262212 2495 262228
rect 2557 263004 2591 263020
rect 2557 262212 2591 262228
rect 2671 263004 2705 263020
rect 2671 262212 2705 262228
rect 2767 263004 2801 263020
rect 2767 262212 2801 262228
rect 2881 263004 2915 263020
rect 2881 262212 2915 262228
rect 2977 263004 3011 263020
rect 2977 262212 3011 262228
rect 3091 263004 3125 263020
rect 3091 262212 3125 262228
rect 3187 263004 3221 263020
rect 3187 262212 3221 262228
rect 3301 263004 3335 263020
rect 3301 262212 3335 262228
rect 3397 263004 3431 263020
rect 3397 262212 3431 262228
rect 3511 263004 3545 263020
rect 3511 262212 3545 262228
rect 3607 263004 3641 263020
rect 3607 262212 3641 262228
rect 3721 263004 3755 263020
rect 3721 262212 3755 262228
rect 3817 263004 3851 263020
rect 3817 262212 3851 262228
rect 3931 263004 3965 263020
rect 3931 262212 3965 262228
rect 4027 263004 4061 263020
rect 4027 262212 4061 262228
rect 4141 263004 4175 263020
rect 4141 262212 4175 262228
rect 4237 263004 4271 263020
rect 4237 262212 4271 262228
rect 4351 263004 4385 263020
rect 4351 262212 4385 262228
rect 4447 263004 4481 263020
rect 4447 262212 4481 262228
rect 4561 263004 4595 263020
rect 4561 262212 4595 262228
rect 4657 263004 4691 263020
rect 4657 262212 4691 262228
rect 4771 263004 4805 263020
rect 4771 262212 4805 262228
rect 4867 263004 4901 263020
rect 4867 262212 4901 262228
rect 4981 263004 5015 263020
rect 4981 262212 5015 262228
rect 5077 263004 5111 263020
rect 5077 262212 5111 262228
rect 5191 263004 5225 263020
rect 5191 262212 5225 262228
rect 5287 263004 5321 263020
rect 5287 262212 5321 262228
rect 5401 263004 5435 263020
rect 5401 262212 5435 262228
rect 5497 263004 5531 263020
rect 5497 262212 5531 262228
rect 5611 263004 5645 263020
rect 5611 262212 5645 262228
rect 5707 263004 5741 263020
rect 5707 262212 5741 262228
rect 5821 263004 5855 263020
rect 5821 262212 5855 262228
rect 5917 263004 5951 263020
rect 5917 262212 5951 262228
rect 6031 263004 6065 263020
rect 6031 262212 6065 262228
rect 6127 263004 6161 263020
rect 6127 262212 6161 262228
rect 6241 263004 6275 263020
rect 6241 262212 6275 262228
rect 6337 263004 6371 263020
rect 6337 262212 6371 262228
rect 6451 263004 6485 263020
rect 6451 262212 6485 262228
rect 6547 263004 6581 263020
rect 6547 262212 6581 262228
rect 6661 263004 6695 263020
rect 6661 262212 6695 262228
rect 6757 263004 6791 263020
rect 6757 262212 6791 262228
rect 6871 263004 6905 263020
rect 6871 262212 6905 262228
rect 6967 263004 7001 263020
rect 6967 262212 7001 262228
rect 7081 263004 7115 263020
rect 7081 262212 7115 262228
rect 7177 263004 7211 263020
rect 7177 262212 7211 262228
rect 7291 263004 7325 263020
rect 7291 262212 7325 262228
rect 7387 263004 7421 263020
rect 7387 262212 7421 262228
rect 7501 263004 7535 263020
rect 7501 262212 7535 262228
rect 7597 263004 7631 263020
rect 7597 262212 7631 262228
rect 7711 263004 7745 263020
rect 7711 262212 7745 262228
rect 7807 263004 7841 263020
rect 7807 262212 7841 262228
rect 7921 263004 7955 263020
rect 7921 262212 7955 262228
rect 8017 263004 8051 263020
rect 8017 262212 8051 262228
rect 8131 263004 8165 263020
rect 8131 262212 8165 262228
rect 8227 263004 8261 263020
rect 8227 262212 8261 262228
rect 8341 263004 8375 263020
rect 8341 262212 8375 262228
rect 8437 263004 8471 263020
rect 8437 262212 8471 262228
rect 8551 263004 8585 263020
rect 8551 262212 8585 262228
rect 8647 263004 8681 263020
rect 8647 262212 8681 262228
rect 8761 263004 8795 263020
rect 8761 262212 8795 262228
rect 8857 263004 8891 263020
rect 8857 262212 8891 262228
rect 8971 263004 9005 263020
rect 8971 262212 9005 262228
rect 9067 263004 9101 263020
rect 9067 262212 9101 262228
rect 9181 263004 9215 263020
rect 9181 262212 9215 262228
rect 9277 263004 9311 263020
rect 9277 262212 9311 262228
rect 9391 263004 9425 263020
rect 9391 262212 9425 262228
rect 9487 263004 9521 263020
rect 9487 262212 9521 262228
rect 9601 263004 9635 263020
rect 9601 262212 9635 262228
rect 9697 263004 9731 263020
rect 9697 262212 9731 262228
rect 9811 263004 9845 263020
rect 9811 262212 9845 262228
rect 9907 263004 9941 263020
rect 9907 262212 9941 262228
rect 10021 263004 10055 263020
rect 10021 262212 10055 262228
rect 10117 263004 10151 263020
rect 10117 262212 10151 262228
rect 10231 263004 10265 263020
rect 10231 262212 10265 262228
rect 10327 263004 10361 263020
rect 10327 262212 10361 262228
rect 10441 263004 10475 263020
rect 10441 262212 10475 262228
rect 10537 263004 10571 263020
rect 10537 262212 10571 262228
rect 10651 263004 10685 263020
rect 10651 262212 10685 262228
rect 10747 263004 10781 263020
rect 10747 262212 10781 262228
rect 10861 263004 10895 263020
rect 10861 262212 10895 262228
rect 10957 263004 10991 263020
rect 10957 262212 10991 262228
rect 11071 263004 11105 263020
rect 11071 262212 11105 262228
rect 11167 263004 11201 263020
rect 11167 262212 11201 262228
rect 11281 263004 11315 263020
rect 11281 262212 11315 262228
rect 11377 263004 11411 263020
rect 11377 262212 11411 262228
rect 11491 263004 11525 263020
rect 11491 262212 11525 262228
rect 11587 263004 11621 263020
rect 11587 262212 11621 262228
rect 11701 263004 11735 263020
rect 11701 262212 11735 262228
rect 11797 263004 11831 263020
rect 11797 262212 11831 262228
rect 11911 263004 11945 263020
rect 11911 262212 11945 262228
rect 12007 263004 12041 263020
rect 12007 262212 12041 262228
rect 12121 263004 12155 263020
rect 12121 262212 12155 262228
rect 12217 263004 12251 263020
rect 12217 262212 12251 262228
rect 12331 263004 12365 263020
rect 12331 262212 12365 262228
rect 12427 263004 12461 263020
rect 12427 262212 12461 262228
rect 12541 263004 12575 263020
rect 12541 262212 12575 262228
rect 12637 263004 12671 263020
rect 12637 262212 12671 262228
rect 12751 263004 12785 263020
rect 12751 262212 12785 262228
rect 12847 263004 12881 263020
rect 12847 262212 12881 262228
rect 12961 263004 12995 263020
rect 12961 262212 12995 262228
rect 13057 263004 13091 263020
rect 13057 262212 13091 262228
rect 13171 263004 13205 263020
rect 13171 262212 13205 262228
rect 13267 263004 13301 263020
rect 13267 262212 13301 262228
rect 13381 263004 13415 263020
rect 13381 262212 13415 262228
rect 13477 263004 13511 263020
rect 13477 262212 13511 262228
rect 13591 263004 13625 263020
rect 13591 262212 13625 262228
rect 13687 263004 13721 263020
rect 13687 262212 13721 262228
rect 13801 263004 13835 263020
rect 13801 262212 13835 262228
rect 13897 263004 13931 263020
rect 13897 262212 13931 262228
rect 14011 263004 14045 263020
rect 14011 262212 14045 262228
rect 14107 263004 14141 263020
rect 14107 262212 14141 262228
rect 14221 263004 14255 263020
rect 14221 262212 14255 262228
rect 14317 263004 14351 263020
rect 14317 262212 14351 262228
rect 14431 263004 14465 263020
rect 14431 262212 14465 262228
rect 14527 263004 14561 263020
rect 14527 262212 14561 262228
rect 14641 263004 14675 263020
rect 14641 262212 14675 262228
rect 14737 263004 14771 263020
rect 14737 262212 14771 262228
rect 14851 263004 14885 263020
rect 14851 262212 14885 262228
rect 14947 263004 14981 263020
rect 14947 262212 14981 262228
rect 15061 263004 15095 263020
rect 15061 262212 15095 262228
rect 15157 263004 15191 263020
rect 15157 262212 15191 262228
rect 15271 263004 15305 263020
rect 15271 262212 15305 262228
rect 15367 263004 15401 263020
rect 15367 262212 15401 262228
rect 15481 263004 15515 263020
rect 15481 262212 15515 262228
rect 15577 263004 15611 263020
rect 15577 262212 15611 262228
rect 15691 263004 15725 263020
rect 15691 262212 15725 262228
rect 15787 263004 15821 263020
rect 15787 262212 15821 262228
rect 15901 263004 15935 263020
rect 15901 262212 15935 262228
rect 15997 263004 16031 263020
rect 15997 262212 16031 262228
rect 16111 263004 16145 263020
rect 16111 262212 16145 262228
rect 16207 263004 16241 263020
rect 16207 262212 16241 262228
rect 16321 263004 16355 263020
rect 16321 262212 16355 262228
rect 16417 263004 16451 263020
rect 16417 262212 16451 262228
rect 16531 263004 16565 263020
rect 16531 262212 16565 262228
rect 16627 263004 16661 263020
rect 16627 262212 16661 262228
rect 16741 263004 16775 263020
rect 16741 262212 16775 262228
rect 16837 263004 16871 263020
rect 16837 262212 16871 262228
rect 16951 263004 16985 263020
rect 16951 262212 16985 262228
rect 17047 263004 17081 263020
rect 17047 262212 17081 262228
rect 17161 263004 17195 263020
rect 17161 262212 17195 262228
rect 17257 263004 17291 263020
rect 17257 262212 17291 262228
rect 17371 263004 17405 263020
rect 17371 262212 17405 262228
rect 17467 263004 17501 263020
rect 17467 262212 17501 262228
rect 17581 263004 17615 263020
rect 17581 262212 17615 262228
rect 17677 263004 17711 263020
rect 17677 262212 17711 262228
rect 17791 263004 17825 263020
rect 17791 262212 17825 262228
rect 17887 263004 17921 263020
rect 17887 262212 17921 262228
rect 18001 263004 18035 263020
rect 18001 262212 18035 262228
rect 18097 263004 18131 263020
rect 18097 262212 18131 262228
rect 18211 263004 18245 263020
rect 18211 262212 18245 262228
rect 18307 263004 18341 263020
rect 18307 262212 18341 262228
rect 18421 263004 18455 263020
rect 18421 262212 18455 262228
rect 18517 263004 18551 263020
rect 18517 262212 18551 262228
rect 18631 263004 18665 263020
rect 18631 262212 18665 262228
rect 18727 263004 18761 263020
rect 18727 262212 18761 262228
rect 18841 263004 18875 263020
rect 18841 262212 18875 262228
rect 18937 263004 18971 263020
rect 18937 262212 18971 262228
rect 19051 263004 19085 263020
rect 19051 262212 19085 262228
rect 19147 263004 19181 263020
rect 19147 262212 19181 262228
rect 19261 263004 19295 263020
rect 19261 262212 19295 262228
rect 19357 263004 19391 263020
rect 19357 262212 19391 262228
rect 19471 263004 19505 263020
rect 19471 262212 19505 262228
rect 19567 263004 19601 263020
rect 19567 262212 19601 262228
rect 19681 263004 19715 263020
rect 19681 262212 19715 262228
rect 19777 263004 19811 263020
rect 19777 262212 19811 262228
rect 19891 263004 19925 263020
rect 19891 262212 19925 262228
rect 19987 263004 20021 263020
rect 19987 262212 20021 262228
rect 20101 263004 20135 263020
rect 20101 262212 20135 262228
rect 20197 263004 20231 263020
rect 20197 262212 20231 262228
rect 20311 263004 20345 263020
rect 20311 262212 20345 262228
rect 20407 263004 20441 263020
rect 20407 262212 20441 262228
rect 20521 263004 20555 263020
rect 20521 262212 20555 262228
rect 20617 263004 20651 263020
rect 20617 262212 20651 262228
rect 20731 263004 20765 263020
rect 20731 262212 20765 262228
rect 20827 263004 20861 263020
rect 20827 262212 20861 262228
rect 20941 263004 20975 263020
rect 20941 262212 20975 262228
rect 21037 263004 21071 263020
rect 21037 262212 21071 262228
rect 21151 263004 21185 263020
rect 21151 262212 21185 262228
rect 21247 263004 21281 263020
rect 21247 262212 21281 262228
rect 21361 263004 21395 263020
rect 21361 262212 21395 262228
rect 21457 263004 21491 263020
rect 21457 262212 21491 262228
rect 21571 263004 21605 263020
rect 21571 262212 21605 262228
rect 21667 263004 21701 263020
rect 21667 262212 21701 262228
rect 21781 263004 21815 263020
rect 21781 262212 21815 262228
rect 21877 263004 21911 263020
rect 21877 262212 21911 262228
rect 21991 263004 22025 263020
rect 21991 262212 22025 262228
rect 22087 263004 22121 263020
rect 22087 262212 22121 262228
rect 22201 263004 22235 263020
rect 22201 262212 22235 262228
rect 22297 263004 22331 263020
rect 22297 262212 22331 262228
rect 22411 263004 22445 263020
rect 22411 262212 22445 262228
rect 22507 263004 22541 263020
rect 22507 262212 22541 262228
rect 22621 263004 22655 263020
rect 22621 262212 22655 262228
rect 22717 263004 22751 263020
rect 22717 262212 22751 262228
rect 22831 263004 22865 263020
rect 22831 262212 22865 262228
rect 22927 263004 22961 263020
rect 22927 262212 22961 262228
rect 23041 263004 23075 263020
rect 23041 262212 23075 262228
rect 23137 263004 23171 263020
rect 23137 262212 23171 262228
rect 23251 263004 23285 263020
rect 23251 262212 23285 262228
rect 23347 263004 23381 263020
rect 23347 262212 23381 262228
rect 23461 263004 23495 263020
rect 23461 262212 23495 262228
rect 23557 263004 23591 263020
rect 23557 262212 23591 262228
rect 23671 263004 23705 263020
rect 23671 262212 23705 262228
rect 23767 263004 23801 263020
rect 23767 262212 23801 262228
rect 23881 263004 23915 263020
rect 23881 262212 23915 262228
rect 23977 263004 24011 263020
rect 23977 262212 24011 262228
rect 24091 263004 24125 263020
rect 24091 262212 24125 262228
rect 24187 263004 24221 263020
rect 24187 262212 24221 262228
rect 24301 263004 24335 263020
rect 24301 262212 24335 262228
rect 24397 263004 24431 263020
rect 24397 262212 24431 262228
rect 24511 263004 24545 263020
rect 24511 262212 24545 262228
rect 24607 263004 24641 263020
rect 24607 262212 24641 262228
rect 24721 263004 24755 263020
rect 24721 262212 24755 262228
rect 24817 263004 24851 263020
rect 24817 262212 24851 262228
rect 24931 263004 24965 263020
rect 24931 262212 24965 262228
rect 25027 263004 25061 263020
rect 25027 262212 25061 262228
rect 25141 263004 25175 263020
rect 25141 262212 25175 262228
rect 25237 263004 25271 263020
rect 25237 262212 25271 262228
rect 25351 263004 25385 263020
rect 25351 262212 25385 262228
rect 25447 263004 25481 263020
rect 25447 262212 25481 262228
rect 25561 263004 25595 263020
rect 25561 262212 25595 262228
rect 25657 263004 25691 263020
rect 25657 262212 25691 262228
rect 25771 263004 25805 263020
rect 25771 262212 25805 262228
rect 25867 263004 25901 263020
rect 25867 262212 25901 262228
rect 25981 263004 26015 263020
rect 25981 262212 26015 262228
rect 26077 263004 26111 263020
rect 26077 262212 26111 262228
rect 26191 263004 26225 263020
rect 26191 262212 26225 262228
rect 26287 263004 26321 263020
rect 26287 262212 26321 262228
rect 26401 263004 26435 263020
rect 26401 262212 26435 262228
rect 26497 263004 26531 263020
rect 26497 262212 26531 262228
rect 26611 263004 26645 263020
rect 26611 262212 26645 262228
rect 26707 263004 26741 263020
rect 26707 262212 26741 262228
rect 26821 263004 26855 263020
rect 26821 262212 26855 262228
rect 26917 263004 26951 263020
rect 26917 262212 26951 262228
rect 27031 263004 27065 263020
rect 27031 262212 27065 262228
rect 27127 263004 27161 263020
rect 27127 262212 27161 262228
rect 27241 263004 27275 263020
rect 27241 262212 27275 262228
rect 27337 263004 27371 263020
rect 27337 262212 27371 262228
rect -4017 262144 -4001 262178
rect -3905 262144 -3889 262178
rect -3597 262144 -3581 262178
rect -3485 262144 -3469 262178
rect -3177 262144 -3161 262178
rect -3065 262144 -3049 262178
rect -2757 262144 -2741 262178
rect -2645 262144 -2629 262178
rect -2337 262144 -2321 262178
rect -2225 262144 -2209 262178
rect -1917 262144 -1901 262178
rect -1805 262144 -1789 262178
rect -1497 262144 -1481 262178
rect -1385 262144 -1369 262178
rect -1077 262144 -1061 262178
rect -965 262144 -949 262178
rect -657 262144 -641 262178
rect -545 262144 -529 262178
rect -237 262144 -221 262178
rect -125 262144 -109 262178
rect 183 262144 199 262178
rect 295 262144 311 262178
rect 603 262144 619 262178
rect 715 262144 731 262178
rect 1023 262144 1039 262178
rect 1135 262144 1151 262178
rect 1443 262144 1459 262178
rect 1555 262144 1571 262178
rect 1863 262144 1879 262178
rect 1975 262144 1991 262178
rect 2283 262144 2299 262178
rect 2395 262144 2411 262178
rect 2703 262144 2719 262178
rect 2815 262144 2831 262178
rect 3123 262144 3139 262178
rect 3235 262144 3251 262178
rect 3543 262144 3559 262178
rect 3655 262144 3671 262178
rect 3963 262144 3979 262178
rect 4075 262144 4091 262178
rect 4383 262144 4399 262178
rect 4495 262144 4511 262178
rect 4803 262144 4819 262178
rect 4915 262144 4931 262178
rect 5223 262144 5239 262178
rect 5335 262144 5351 262178
rect 5643 262144 5659 262178
rect 5755 262144 5771 262178
rect 6063 262144 6079 262178
rect 6175 262144 6191 262178
rect 6483 262144 6499 262178
rect 6595 262144 6611 262178
rect 6903 262144 6919 262178
rect 7015 262144 7031 262178
rect 7323 262144 7339 262178
rect 7435 262144 7451 262178
rect 7743 262144 7759 262178
rect 7855 262144 7871 262178
rect 8163 262144 8179 262178
rect 8275 262144 8291 262178
rect 8583 262144 8599 262178
rect 8695 262144 8711 262178
rect 9003 262144 9019 262178
rect 9115 262144 9131 262178
rect 9423 262144 9439 262178
rect 9535 262144 9551 262178
rect 9843 262144 9859 262178
rect 9955 262144 9971 262178
rect 10263 262144 10279 262178
rect 10375 262144 10391 262178
rect 10683 262144 10699 262178
rect 10795 262144 10811 262178
rect 11103 262144 11119 262178
rect 11215 262144 11231 262178
rect 11523 262144 11539 262178
rect 11635 262144 11651 262178
rect 11943 262144 11959 262178
rect 12055 262144 12071 262178
rect 12363 262144 12379 262178
rect 12475 262144 12491 262178
rect 12783 262144 12799 262178
rect 12895 262144 12911 262178
rect 13203 262144 13219 262178
rect 13315 262144 13331 262178
rect 13623 262144 13639 262178
rect 13735 262144 13751 262178
rect 14043 262144 14059 262178
rect 14155 262144 14171 262178
rect 14463 262144 14479 262178
rect 14575 262144 14591 262178
rect 14883 262144 14899 262178
rect 14995 262144 15011 262178
rect 15303 262144 15319 262178
rect 15415 262144 15431 262178
rect 15723 262144 15739 262178
rect 15835 262144 15851 262178
rect 16143 262144 16159 262178
rect 16255 262144 16271 262178
rect 16563 262144 16579 262178
rect 16675 262144 16691 262178
rect 16983 262144 16999 262178
rect 17095 262144 17111 262178
rect 17403 262144 17419 262178
rect 17515 262144 17531 262178
rect 17823 262144 17839 262178
rect 17935 262144 17951 262178
rect 18243 262144 18259 262178
rect 18355 262144 18371 262178
rect 18663 262144 18679 262178
rect 18775 262144 18791 262178
rect 19083 262144 19099 262178
rect 19195 262144 19211 262178
rect 19503 262144 19519 262178
rect 19615 262144 19631 262178
rect 19923 262144 19939 262178
rect 20035 262144 20051 262178
rect 20343 262144 20359 262178
rect 20455 262144 20471 262178
rect 20763 262144 20779 262178
rect 20875 262144 20891 262178
rect 21183 262144 21199 262178
rect 21295 262144 21311 262178
rect 21603 262144 21619 262178
rect 21715 262144 21731 262178
rect 22023 262144 22039 262178
rect 22135 262144 22151 262178
rect 22443 262144 22459 262178
rect 22555 262144 22571 262178
rect 22863 262144 22879 262178
rect 22975 262144 22991 262178
rect 23283 262144 23299 262178
rect 23395 262144 23411 262178
rect 23703 262144 23719 262178
rect 23815 262144 23831 262178
rect 24123 262144 24139 262178
rect 24235 262144 24251 262178
rect 24543 262144 24559 262178
rect 24655 262144 24671 262178
rect 24963 262144 24979 262178
rect 25075 262144 25091 262178
rect 25383 262144 25399 262178
rect 25495 262144 25511 262178
rect 25803 262144 25819 262178
rect 25915 262144 25931 262178
rect 26223 262144 26239 262178
rect 26335 262144 26351 262178
rect 26643 262144 26659 262178
rect 26755 262144 26771 262178
rect 27063 262144 27079 262178
rect 27175 262144 27191 262178
rect -4163 262076 -4129 262138
rect 27451 262076 27485 262138
rect -4163 262042 -4067 262076
rect 27389 262042 27485 262076
rect -4163 254650 -4067 254684
rect 27389 254650 27485 254684
rect -4163 254588 -4129 254650
rect 27451 254588 27485 254650
rect -4017 254548 -4001 254582
rect -3905 254548 -3889 254582
rect -3597 254548 -3581 254582
rect -3485 254548 -3469 254582
rect -3177 254548 -3161 254582
rect -3065 254548 -3049 254582
rect -2757 254548 -2741 254582
rect -2645 254548 -2629 254582
rect -2337 254548 -2321 254582
rect -2225 254548 -2209 254582
rect -1917 254548 -1901 254582
rect -1805 254548 -1789 254582
rect -1497 254548 -1481 254582
rect -1385 254548 -1369 254582
rect -1077 254548 -1061 254582
rect -965 254548 -949 254582
rect -657 254548 -641 254582
rect -545 254548 -529 254582
rect -237 254548 -221 254582
rect -125 254548 -109 254582
rect 183 254548 199 254582
rect 295 254548 311 254582
rect 603 254548 619 254582
rect 715 254548 731 254582
rect 1023 254548 1039 254582
rect 1135 254548 1151 254582
rect 1443 254548 1459 254582
rect 1555 254548 1571 254582
rect 1863 254548 1879 254582
rect 1975 254548 1991 254582
rect 2283 254548 2299 254582
rect 2395 254548 2411 254582
rect 2703 254548 2719 254582
rect 2815 254548 2831 254582
rect 3123 254548 3139 254582
rect 3235 254548 3251 254582
rect 3543 254548 3559 254582
rect 3655 254548 3671 254582
rect 3963 254548 3979 254582
rect 4075 254548 4091 254582
rect 4383 254548 4399 254582
rect 4495 254548 4511 254582
rect 4803 254548 4819 254582
rect 4915 254548 4931 254582
rect 5223 254548 5239 254582
rect 5335 254548 5351 254582
rect 5643 254548 5659 254582
rect 5755 254548 5771 254582
rect 6063 254548 6079 254582
rect 6175 254548 6191 254582
rect 6483 254548 6499 254582
rect 6595 254548 6611 254582
rect 6903 254548 6919 254582
rect 7015 254548 7031 254582
rect 7323 254548 7339 254582
rect 7435 254548 7451 254582
rect 7743 254548 7759 254582
rect 7855 254548 7871 254582
rect 8163 254548 8179 254582
rect 8275 254548 8291 254582
rect 8583 254548 8599 254582
rect 8695 254548 8711 254582
rect 9003 254548 9019 254582
rect 9115 254548 9131 254582
rect 9423 254548 9439 254582
rect 9535 254548 9551 254582
rect 9843 254548 9859 254582
rect 9955 254548 9971 254582
rect 10263 254548 10279 254582
rect 10375 254548 10391 254582
rect 10683 254548 10699 254582
rect 10795 254548 10811 254582
rect 11103 254548 11119 254582
rect 11215 254548 11231 254582
rect 11523 254548 11539 254582
rect 11635 254548 11651 254582
rect 11943 254548 11959 254582
rect 12055 254548 12071 254582
rect 12363 254548 12379 254582
rect 12475 254548 12491 254582
rect 12783 254548 12799 254582
rect 12895 254548 12911 254582
rect 13203 254548 13219 254582
rect 13315 254548 13331 254582
rect 13623 254548 13639 254582
rect 13735 254548 13751 254582
rect 14043 254548 14059 254582
rect 14155 254548 14171 254582
rect 14463 254548 14479 254582
rect 14575 254548 14591 254582
rect 14883 254548 14899 254582
rect 14995 254548 15011 254582
rect 15303 254548 15319 254582
rect 15415 254548 15431 254582
rect 15723 254548 15739 254582
rect 15835 254548 15851 254582
rect 16143 254548 16159 254582
rect 16255 254548 16271 254582
rect 16563 254548 16579 254582
rect 16675 254548 16691 254582
rect 16983 254548 16999 254582
rect 17095 254548 17111 254582
rect 17403 254548 17419 254582
rect 17515 254548 17531 254582
rect 17823 254548 17839 254582
rect 17935 254548 17951 254582
rect 18243 254548 18259 254582
rect 18355 254548 18371 254582
rect 18663 254548 18679 254582
rect 18775 254548 18791 254582
rect 19083 254548 19099 254582
rect 19195 254548 19211 254582
rect 19503 254548 19519 254582
rect 19615 254548 19631 254582
rect 19923 254548 19939 254582
rect 20035 254548 20051 254582
rect 20343 254548 20359 254582
rect 20455 254548 20471 254582
rect 20763 254548 20779 254582
rect 20875 254548 20891 254582
rect 21183 254548 21199 254582
rect 21295 254548 21311 254582
rect 21603 254548 21619 254582
rect 21715 254548 21731 254582
rect 22023 254548 22039 254582
rect 22135 254548 22151 254582
rect 22443 254548 22459 254582
rect 22555 254548 22571 254582
rect 22863 254548 22879 254582
rect 22975 254548 22991 254582
rect 23283 254548 23299 254582
rect 23395 254548 23411 254582
rect 23703 254548 23719 254582
rect 23815 254548 23831 254582
rect 24123 254548 24139 254582
rect 24235 254548 24251 254582
rect 24543 254548 24559 254582
rect 24655 254548 24671 254582
rect 24963 254548 24979 254582
rect 25075 254548 25091 254582
rect 25383 254548 25399 254582
rect 25495 254548 25511 254582
rect 25803 254548 25819 254582
rect 25915 254548 25931 254582
rect 26223 254548 26239 254582
rect 26335 254548 26351 254582
rect 26643 254548 26659 254582
rect 26755 254548 26771 254582
rect 27063 254548 27079 254582
rect 27175 254548 27191 254582
rect -4049 254489 -4015 254505
rect -4049 253697 -4015 253713
rect -3953 254489 -3919 254505
rect -3953 253697 -3919 253713
rect -3839 254489 -3805 254505
rect -3839 253697 -3805 253713
rect -3743 254489 -3709 254505
rect -3743 253697 -3709 253713
rect -3629 254489 -3595 254505
rect -3629 253697 -3595 253713
rect -3533 254489 -3499 254505
rect -3533 253697 -3499 253713
rect -3419 254489 -3385 254505
rect -3419 253697 -3385 253713
rect -3323 254489 -3289 254505
rect -3323 253697 -3289 253713
rect -3209 254489 -3175 254505
rect -3209 253697 -3175 253713
rect -3113 254489 -3079 254505
rect -3113 253697 -3079 253713
rect -2999 254489 -2965 254505
rect -2999 253697 -2965 253713
rect -2903 254489 -2869 254505
rect -2903 253697 -2869 253713
rect -2789 254489 -2755 254505
rect -2789 253697 -2755 253713
rect -2693 254489 -2659 254505
rect -2693 253697 -2659 253713
rect -2579 254489 -2545 254505
rect -2579 253697 -2545 253713
rect -2483 254489 -2449 254505
rect -2483 253697 -2449 253713
rect -2369 254489 -2335 254505
rect -2369 253697 -2335 253713
rect -2273 254489 -2239 254505
rect -2273 253697 -2239 253713
rect -2159 254489 -2125 254505
rect -2159 253697 -2125 253713
rect -2063 254489 -2029 254505
rect -2063 253697 -2029 253713
rect -1949 254489 -1915 254505
rect -1949 253697 -1915 253713
rect -1853 254489 -1819 254505
rect -1853 253697 -1819 253713
rect -1739 254489 -1705 254505
rect -1739 253697 -1705 253713
rect -1643 254489 -1609 254505
rect -1643 253697 -1609 253713
rect -1529 254489 -1495 254505
rect -1529 253697 -1495 253713
rect -1433 254489 -1399 254505
rect -1433 253697 -1399 253713
rect -1319 254489 -1285 254505
rect -1319 253697 -1285 253713
rect -1223 254489 -1189 254505
rect -1223 253697 -1189 253713
rect -1109 254489 -1075 254505
rect -1109 253697 -1075 253713
rect -1013 254489 -979 254505
rect -1013 253697 -979 253713
rect -899 254489 -865 254505
rect -899 253697 -865 253713
rect -803 254489 -769 254505
rect -803 253697 -769 253713
rect -689 254489 -655 254505
rect -689 253697 -655 253713
rect -593 254489 -559 254505
rect -593 253697 -559 253713
rect -479 254489 -445 254505
rect -479 253697 -445 253713
rect -383 254489 -349 254505
rect -383 253697 -349 253713
rect -269 254489 -235 254505
rect -269 253697 -235 253713
rect -173 254489 -139 254505
rect -173 253697 -139 253713
rect -59 254489 -25 254505
rect -59 253697 -25 253713
rect 37 254489 71 254505
rect 37 253697 71 253713
rect 151 254489 185 254505
rect 151 253697 185 253713
rect 247 254489 281 254505
rect 247 253697 281 253713
rect 361 254489 395 254505
rect 361 253697 395 253713
rect 457 254489 491 254505
rect 457 253697 491 253713
rect 571 254489 605 254505
rect 571 253697 605 253713
rect 667 254489 701 254505
rect 667 253697 701 253713
rect 781 254489 815 254505
rect 781 253697 815 253713
rect 877 254489 911 254505
rect 877 253697 911 253713
rect 991 254489 1025 254505
rect 991 253697 1025 253713
rect 1087 254489 1121 254505
rect 1087 253697 1121 253713
rect 1201 254489 1235 254505
rect 1201 253697 1235 253713
rect 1297 254489 1331 254505
rect 1297 253697 1331 253713
rect 1411 254489 1445 254505
rect 1411 253697 1445 253713
rect 1507 254489 1541 254505
rect 1507 253697 1541 253713
rect 1621 254489 1655 254505
rect 1621 253697 1655 253713
rect 1717 254489 1751 254505
rect 1717 253697 1751 253713
rect 1831 254489 1865 254505
rect 1831 253697 1865 253713
rect 1927 254489 1961 254505
rect 1927 253697 1961 253713
rect 2041 254489 2075 254505
rect 2041 253697 2075 253713
rect 2137 254489 2171 254505
rect 2137 253697 2171 253713
rect 2251 254489 2285 254505
rect 2251 253697 2285 253713
rect 2347 254489 2381 254505
rect 2347 253697 2381 253713
rect 2461 254489 2495 254505
rect 2461 253697 2495 253713
rect 2557 254489 2591 254505
rect 2557 253697 2591 253713
rect 2671 254489 2705 254505
rect 2671 253697 2705 253713
rect 2767 254489 2801 254505
rect 2767 253697 2801 253713
rect 2881 254489 2915 254505
rect 2881 253697 2915 253713
rect 2977 254489 3011 254505
rect 2977 253697 3011 253713
rect 3091 254489 3125 254505
rect 3091 253697 3125 253713
rect 3187 254489 3221 254505
rect 3187 253697 3221 253713
rect 3301 254489 3335 254505
rect 3301 253697 3335 253713
rect 3397 254489 3431 254505
rect 3397 253697 3431 253713
rect 3511 254489 3545 254505
rect 3511 253697 3545 253713
rect 3607 254489 3641 254505
rect 3607 253697 3641 253713
rect 3721 254489 3755 254505
rect 3721 253697 3755 253713
rect 3817 254489 3851 254505
rect 3817 253697 3851 253713
rect 3931 254489 3965 254505
rect 3931 253697 3965 253713
rect 4027 254489 4061 254505
rect 4027 253697 4061 253713
rect 4141 254489 4175 254505
rect 4141 253697 4175 253713
rect 4237 254489 4271 254505
rect 4237 253697 4271 253713
rect 4351 254489 4385 254505
rect 4351 253697 4385 253713
rect 4447 254489 4481 254505
rect 4447 253697 4481 253713
rect 4561 254489 4595 254505
rect 4561 253697 4595 253713
rect 4657 254489 4691 254505
rect 4657 253697 4691 253713
rect 4771 254489 4805 254505
rect 4771 253697 4805 253713
rect 4867 254489 4901 254505
rect 4867 253697 4901 253713
rect 4981 254489 5015 254505
rect 4981 253697 5015 253713
rect 5077 254489 5111 254505
rect 5077 253697 5111 253713
rect 5191 254489 5225 254505
rect 5191 253697 5225 253713
rect 5287 254489 5321 254505
rect 5287 253697 5321 253713
rect 5401 254489 5435 254505
rect 5401 253697 5435 253713
rect 5497 254489 5531 254505
rect 5497 253697 5531 253713
rect 5611 254489 5645 254505
rect 5611 253697 5645 253713
rect 5707 254489 5741 254505
rect 5707 253697 5741 253713
rect 5821 254489 5855 254505
rect 5821 253697 5855 253713
rect 5917 254489 5951 254505
rect 5917 253697 5951 253713
rect 6031 254489 6065 254505
rect 6031 253697 6065 253713
rect 6127 254489 6161 254505
rect 6127 253697 6161 253713
rect 6241 254489 6275 254505
rect 6241 253697 6275 253713
rect 6337 254489 6371 254505
rect 6337 253697 6371 253713
rect 6451 254489 6485 254505
rect 6451 253697 6485 253713
rect 6547 254489 6581 254505
rect 6547 253697 6581 253713
rect 6661 254489 6695 254505
rect 6661 253697 6695 253713
rect 6757 254489 6791 254505
rect 6757 253697 6791 253713
rect 6871 254489 6905 254505
rect 6871 253697 6905 253713
rect 6967 254489 7001 254505
rect 6967 253697 7001 253713
rect 7081 254489 7115 254505
rect 7081 253697 7115 253713
rect 7177 254489 7211 254505
rect 7177 253697 7211 253713
rect 7291 254489 7325 254505
rect 7291 253697 7325 253713
rect 7387 254489 7421 254505
rect 7387 253697 7421 253713
rect 7501 254489 7535 254505
rect 7501 253697 7535 253713
rect 7597 254489 7631 254505
rect 7597 253697 7631 253713
rect 7711 254489 7745 254505
rect 7711 253697 7745 253713
rect 7807 254489 7841 254505
rect 7807 253697 7841 253713
rect 7921 254489 7955 254505
rect 7921 253697 7955 253713
rect 8017 254489 8051 254505
rect 8017 253697 8051 253713
rect 8131 254489 8165 254505
rect 8131 253697 8165 253713
rect 8227 254489 8261 254505
rect 8227 253697 8261 253713
rect 8341 254489 8375 254505
rect 8341 253697 8375 253713
rect 8437 254489 8471 254505
rect 8437 253697 8471 253713
rect 8551 254489 8585 254505
rect 8551 253697 8585 253713
rect 8647 254489 8681 254505
rect 8647 253697 8681 253713
rect 8761 254489 8795 254505
rect 8761 253697 8795 253713
rect 8857 254489 8891 254505
rect 8857 253697 8891 253713
rect 8971 254489 9005 254505
rect 8971 253697 9005 253713
rect 9067 254489 9101 254505
rect 9067 253697 9101 253713
rect 9181 254489 9215 254505
rect 9181 253697 9215 253713
rect 9277 254489 9311 254505
rect 9277 253697 9311 253713
rect 9391 254489 9425 254505
rect 9391 253697 9425 253713
rect 9487 254489 9521 254505
rect 9487 253697 9521 253713
rect 9601 254489 9635 254505
rect 9601 253697 9635 253713
rect 9697 254489 9731 254505
rect 9697 253697 9731 253713
rect 9811 254489 9845 254505
rect 9811 253697 9845 253713
rect 9907 254489 9941 254505
rect 9907 253697 9941 253713
rect 10021 254489 10055 254505
rect 10021 253697 10055 253713
rect 10117 254489 10151 254505
rect 10117 253697 10151 253713
rect 10231 254489 10265 254505
rect 10231 253697 10265 253713
rect 10327 254489 10361 254505
rect 10327 253697 10361 253713
rect 10441 254489 10475 254505
rect 10441 253697 10475 253713
rect 10537 254489 10571 254505
rect 10537 253697 10571 253713
rect 10651 254489 10685 254505
rect 10651 253697 10685 253713
rect 10747 254489 10781 254505
rect 10747 253697 10781 253713
rect 10861 254489 10895 254505
rect 10861 253697 10895 253713
rect 10957 254489 10991 254505
rect 10957 253697 10991 253713
rect 11071 254489 11105 254505
rect 11071 253697 11105 253713
rect 11167 254489 11201 254505
rect 11167 253697 11201 253713
rect 11281 254489 11315 254505
rect 11281 253697 11315 253713
rect 11377 254489 11411 254505
rect 11377 253697 11411 253713
rect 11491 254489 11525 254505
rect 11491 253697 11525 253713
rect 11587 254489 11621 254505
rect 11587 253697 11621 253713
rect 11701 254489 11735 254505
rect 11701 253697 11735 253713
rect 11797 254489 11831 254505
rect 11797 253697 11831 253713
rect 11911 254489 11945 254505
rect 11911 253697 11945 253713
rect 12007 254489 12041 254505
rect 12007 253697 12041 253713
rect 12121 254489 12155 254505
rect 12121 253697 12155 253713
rect 12217 254489 12251 254505
rect 12217 253697 12251 253713
rect 12331 254489 12365 254505
rect 12331 253697 12365 253713
rect 12427 254489 12461 254505
rect 12427 253697 12461 253713
rect 12541 254489 12575 254505
rect 12541 253697 12575 253713
rect 12637 254489 12671 254505
rect 12637 253697 12671 253713
rect 12751 254489 12785 254505
rect 12751 253697 12785 253713
rect 12847 254489 12881 254505
rect 12847 253697 12881 253713
rect 12961 254489 12995 254505
rect 12961 253697 12995 253713
rect 13057 254489 13091 254505
rect 13057 253697 13091 253713
rect 13171 254489 13205 254505
rect 13171 253697 13205 253713
rect 13267 254489 13301 254505
rect 13267 253697 13301 253713
rect 13381 254489 13415 254505
rect 13381 253697 13415 253713
rect 13477 254489 13511 254505
rect 13477 253697 13511 253713
rect 13591 254489 13625 254505
rect 13591 253697 13625 253713
rect 13687 254489 13721 254505
rect 13687 253697 13721 253713
rect 13801 254489 13835 254505
rect 13801 253697 13835 253713
rect 13897 254489 13931 254505
rect 13897 253697 13931 253713
rect 14011 254489 14045 254505
rect 14011 253697 14045 253713
rect 14107 254489 14141 254505
rect 14107 253697 14141 253713
rect 14221 254489 14255 254505
rect 14221 253697 14255 253713
rect 14317 254489 14351 254505
rect 14317 253697 14351 253713
rect 14431 254489 14465 254505
rect 14431 253697 14465 253713
rect 14527 254489 14561 254505
rect 14527 253697 14561 253713
rect 14641 254489 14675 254505
rect 14641 253697 14675 253713
rect 14737 254489 14771 254505
rect 14737 253697 14771 253713
rect 14851 254489 14885 254505
rect 14851 253697 14885 253713
rect 14947 254489 14981 254505
rect 14947 253697 14981 253713
rect 15061 254489 15095 254505
rect 15061 253697 15095 253713
rect 15157 254489 15191 254505
rect 15157 253697 15191 253713
rect 15271 254489 15305 254505
rect 15271 253697 15305 253713
rect 15367 254489 15401 254505
rect 15367 253697 15401 253713
rect 15481 254489 15515 254505
rect 15481 253697 15515 253713
rect 15577 254489 15611 254505
rect 15577 253697 15611 253713
rect 15691 254489 15725 254505
rect 15691 253697 15725 253713
rect 15787 254489 15821 254505
rect 15787 253697 15821 253713
rect 15901 254489 15935 254505
rect 15901 253697 15935 253713
rect 15997 254489 16031 254505
rect 15997 253697 16031 253713
rect 16111 254489 16145 254505
rect 16111 253697 16145 253713
rect 16207 254489 16241 254505
rect 16207 253697 16241 253713
rect 16321 254489 16355 254505
rect 16321 253697 16355 253713
rect 16417 254489 16451 254505
rect 16417 253697 16451 253713
rect 16531 254489 16565 254505
rect 16531 253697 16565 253713
rect 16627 254489 16661 254505
rect 16627 253697 16661 253713
rect 16741 254489 16775 254505
rect 16741 253697 16775 253713
rect 16837 254489 16871 254505
rect 16837 253697 16871 253713
rect 16951 254489 16985 254505
rect 16951 253697 16985 253713
rect 17047 254489 17081 254505
rect 17047 253697 17081 253713
rect 17161 254489 17195 254505
rect 17161 253697 17195 253713
rect 17257 254489 17291 254505
rect 17257 253697 17291 253713
rect 17371 254489 17405 254505
rect 17371 253697 17405 253713
rect 17467 254489 17501 254505
rect 17467 253697 17501 253713
rect 17581 254489 17615 254505
rect 17581 253697 17615 253713
rect 17677 254489 17711 254505
rect 17677 253697 17711 253713
rect 17791 254489 17825 254505
rect 17791 253697 17825 253713
rect 17887 254489 17921 254505
rect 17887 253697 17921 253713
rect 18001 254489 18035 254505
rect 18001 253697 18035 253713
rect 18097 254489 18131 254505
rect 18097 253697 18131 253713
rect 18211 254489 18245 254505
rect 18211 253697 18245 253713
rect 18307 254489 18341 254505
rect 18307 253697 18341 253713
rect 18421 254489 18455 254505
rect 18421 253697 18455 253713
rect 18517 254489 18551 254505
rect 18517 253697 18551 253713
rect 18631 254489 18665 254505
rect 18631 253697 18665 253713
rect 18727 254489 18761 254505
rect 18727 253697 18761 253713
rect 18841 254489 18875 254505
rect 18841 253697 18875 253713
rect 18937 254489 18971 254505
rect 18937 253697 18971 253713
rect 19051 254489 19085 254505
rect 19051 253697 19085 253713
rect 19147 254489 19181 254505
rect 19147 253697 19181 253713
rect 19261 254489 19295 254505
rect 19261 253697 19295 253713
rect 19357 254489 19391 254505
rect 19357 253697 19391 253713
rect 19471 254489 19505 254505
rect 19471 253697 19505 253713
rect 19567 254489 19601 254505
rect 19567 253697 19601 253713
rect 19681 254489 19715 254505
rect 19681 253697 19715 253713
rect 19777 254489 19811 254505
rect 19777 253697 19811 253713
rect 19891 254489 19925 254505
rect 19891 253697 19925 253713
rect 19987 254489 20021 254505
rect 19987 253697 20021 253713
rect 20101 254489 20135 254505
rect 20101 253697 20135 253713
rect 20197 254489 20231 254505
rect 20197 253697 20231 253713
rect 20311 254489 20345 254505
rect 20311 253697 20345 253713
rect 20407 254489 20441 254505
rect 20407 253697 20441 253713
rect 20521 254489 20555 254505
rect 20521 253697 20555 253713
rect 20617 254489 20651 254505
rect 20617 253697 20651 253713
rect 20731 254489 20765 254505
rect 20731 253697 20765 253713
rect 20827 254489 20861 254505
rect 20827 253697 20861 253713
rect 20941 254489 20975 254505
rect 20941 253697 20975 253713
rect 21037 254489 21071 254505
rect 21037 253697 21071 253713
rect 21151 254489 21185 254505
rect 21151 253697 21185 253713
rect 21247 254489 21281 254505
rect 21247 253697 21281 253713
rect 21361 254489 21395 254505
rect 21361 253697 21395 253713
rect 21457 254489 21491 254505
rect 21457 253697 21491 253713
rect 21571 254489 21605 254505
rect 21571 253697 21605 253713
rect 21667 254489 21701 254505
rect 21667 253697 21701 253713
rect 21781 254489 21815 254505
rect 21781 253697 21815 253713
rect 21877 254489 21911 254505
rect 21877 253697 21911 253713
rect 21991 254489 22025 254505
rect 21991 253697 22025 253713
rect 22087 254489 22121 254505
rect 22087 253697 22121 253713
rect 22201 254489 22235 254505
rect 22201 253697 22235 253713
rect 22297 254489 22331 254505
rect 22297 253697 22331 253713
rect 22411 254489 22445 254505
rect 22411 253697 22445 253713
rect 22507 254489 22541 254505
rect 22507 253697 22541 253713
rect 22621 254489 22655 254505
rect 22621 253697 22655 253713
rect 22717 254489 22751 254505
rect 22717 253697 22751 253713
rect 22831 254489 22865 254505
rect 22831 253697 22865 253713
rect 22927 254489 22961 254505
rect 22927 253697 22961 253713
rect 23041 254489 23075 254505
rect 23041 253697 23075 253713
rect 23137 254489 23171 254505
rect 23137 253697 23171 253713
rect 23251 254489 23285 254505
rect 23251 253697 23285 253713
rect 23347 254489 23381 254505
rect 23347 253697 23381 253713
rect 23461 254489 23495 254505
rect 23461 253697 23495 253713
rect 23557 254489 23591 254505
rect 23557 253697 23591 253713
rect 23671 254489 23705 254505
rect 23671 253697 23705 253713
rect 23767 254489 23801 254505
rect 23767 253697 23801 253713
rect 23881 254489 23915 254505
rect 23881 253697 23915 253713
rect 23977 254489 24011 254505
rect 23977 253697 24011 253713
rect 24091 254489 24125 254505
rect 24091 253697 24125 253713
rect 24187 254489 24221 254505
rect 24187 253697 24221 253713
rect 24301 254489 24335 254505
rect 24301 253697 24335 253713
rect 24397 254489 24431 254505
rect 24397 253697 24431 253713
rect 24511 254489 24545 254505
rect 24511 253697 24545 253713
rect 24607 254489 24641 254505
rect 24607 253697 24641 253713
rect 24721 254489 24755 254505
rect 24721 253697 24755 253713
rect 24817 254489 24851 254505
rect 24817 253697 24851 253713
rect 24931 254489 24965 254505
rect 24931 253697 24965 253713
rect 25027 254489 25061 254505
rect 25027 253697 25061 253713
rect 25141 254489 25175 254505
rect 25141 253697 25175 253713
rect 25237 254489 25271 254505
rect 25237 253697 25271 253713
rect 25351 254489 25385 254505
rect 25351 253697 25385 253713
rect 25447 254489 25481 254505
rect 25447 253697 25481 253713
rect 25561 254489 25595 254505
rect 25561 253697 25595 253713
rect 25657 254489 25691 254505
rect 25657 253697 25691 253713
rect 25771 254489 25805 254505
rect 25771 253697 25805 253713
rect 25867 254489 25901 254505
rect 25867 253697 25901 253713
rect 25981 254489 26015 254505
rect 25981 253697 26015 253713
rect 26077 254489 26111 254505
rect 26077 253697 26111 253713
rect 26191 254489 26225 254505
rect 26191 253697 26225 253713
rect 26287 254489 26321 254505
rect 26287 253697 26321 253713
rect 26401 254489 26435 254505
rect 26401 253697 26435 253713
rect 26497 254489 26531 254505
rect 26497 253697 26531 253713
rect 26611 254489 26645 254505
rect 26611 253697 26645 253713
rect 26707 254489 26741 254505
rect 26707 253697 26741 253713
rect 26821 254489 26855 254505
rect 26821 253697 26855 253713
rect 26917 254489 26951 254505
rect 26917 253697 26951 253713
rect 27031 254489 27065 254505
rect 27031 253697 27065 253713
rect 27127 254489 27161 254505
rect 27127 253697 27161 253713
rect 27241 254489 27275 254505
rect 27241 253697 27275 253713
rect 27337 254489 27371 254505
rect 27337 253697 27371 253713
rect -3807 253620 -3791 253654
rect -3807 253512 -3791 253546
rect -3757 253620 -3741 253654
rect -3387 253620 -3371 253654
rect -3757 253512 -3741 253546
rect -3387 253512 -3371 253546
rect -3337 253620 -3321 253654
rect -2967 253620 -2951 253654
rect -3337 253512 -3321 253546
rect -2967 253512 -2951 253546
rect -2917 253620 -2901 253654
rect -2547 253620 -2531 253654
rect -2917 253512 -2901 253546
rect -2547 253512 -2531 253546
rect -2497 253620 -2481 253654
rect -2127 253620 -2111 253654
rect -2497 253512 -2481 253546
rect -2127 253512 -2111 253546
rect -2077 253620 -2061 253654
rect -1707 253620 -1691 253654
rect -2077 253512 -2061 253546
rect -1707 253512 -1691 253546
rect -1657 253620 -1641 253654
rect -1287 253620 -1271 253654
rect -1657 253512 -1641 253546
rect -1287 253512 -1271 253546
rect -1237 253620 -1221 253654
rect -867 253620 -851 253654
rect -1237 253512 -1221 253546
rect -867 253512 -851 253546
rect -817 253620 -801 253654
rect -447 253620 -431 253654
rect -817 253512 -801 253546
rect -447 253512 -431 253546
rect -397 253620 -381 253654
rect -27 253620 -11 253654
rect -397 253512 -381 253546
rect -27 253512 -11 253546
rect 23 253620 39 253654
rect 393 253620 409 253654
rect 23 253512 39 253546
rect 393 253512 409 253546
rect 443 253620 459 253654
rect 813 253620 829 253654
rect 443 253512 459 253546
rect 813 253512 829 253546
rect 863 253620 879 253654
rect 1233 253620 1249 253654
rect 863 253512 879 253546
rect 1233 253512 1249 253546
rect 1283 253620 1299 253654
rect 1653 253620 1669 253654
rect 1283 253512 1299 253546
rect 1653 253512 1669 253546
rect 1703 253620 1719 253654
rect 2073 253620 2089 253654
rect 1703 253512 1719 253546
rect 2073 253512 2089 253546
rect 2123 253620 2139 253654
rect 2493 253620 2509 253654
rect 2123 253512 2139 253546
rect 2493 253512 2509 253546
rect 2543 253620 2559 253654
rect 2913 253620 2929 253654
rect 2543 253512 2559 253546
rect 2913 253512 2929 253546
rect 2963 253620 2979 253654
rect 3333 253620 3349 253654
rect 2963 253512 2979 253546
rect 3333 253512 3349 253546
rect 3383 253620 3399 253654
rect 3753 253620 3769 253654
rect 3383 253512 3399 253546
rect 3753 253512 3769 253546
rect 3803 253620 3819 253654
rect 4173 253620 4189 253654
rect 3803 253512 3819 253546
rect 4173 253512 4189 253546
rect 4223 253620 4239 253654
rect 4593 253620 4609 253654
rect 4223 253512 4239 253546
rect 4593 253512 4609 253546
rect 4643 253620 4659 253654
rect 5013 253620 5029 253654
rect 4643 253512 4659 253546
rect 5013 253512 5029 253546
rect 5063 253620 5079 253654
rect 5433 253620 5449 253654
rect 5063 253512 5079 253546
rect 5433 253512 5449 253546
rect 5483 253620 5499 253654
rect 5853 253620 5869 253654
rect 5483 253512 5499 253546
rect 5853 253512 5869 253546
rect 5903 253620 5919 253654
rect 6273 253620 6289 253654
rect 5903 253512 5919 253546
rect 6273 253512 6289 253546
rect 6323 253620 6339 253654
rect 6693 253620 6709 253654
rect 6323 253512 6339 253546
rect 6693 253512 6709 253546
rect 6743 253620 6759 253654
rect 7113 253620 7129 253654
rect 6743 253512 6759 253546
rect 7113 253512 7129 253546
rect 7163 253620 7179 253654
rect 7533 253620 7549 253654
rect 7163 253512 7179 253546
rect 7533 253512 7549 253546
rect 7583 253620 7599 253654
rect 7953 253620 7969 253654
rect 7583 253512 7599 253546
rect 7953 253512 7969 253546
rect 8003 253620 8019 253654
rect 8373 253620 8389 253654
rect 8003 253512 8019 253546
rect 8373 253512 8389 253546
rect 8423 253620 8439 253654
rect 8793 253620 8809 253654
rect 8423 253512 8439 253546
rect 8793 253512 8809 253546
rect 8843 253620 8859 253654
rect 9213 253620 9229 253654
rect 8843 253512 8859 253546
rect 9213 253512 9229 253546
rect 9263 253620 9279 253654
rect 9633 253620 9649 253654
rect 9263 253512 9279 253546
rect 9633 253512 9649 253546
rect 9683 253620 9699 253654
rect 10053 253620 10069 253654
rect 9683 253512 9699 253546
rect 10053 253512 10069 253546
rect 10103 253620 10119 253654
rect 10473 253620 10489 253654
rect 10103 253512 10119 253546
rect 10473 253512 10489 253546
rect 10523 253620 10539 253654
rect 10893 253620 10909 253654
rect 10523 253512 10539 253546
rect 10893 253512 10909 253546
rect 10943 253620 10959 253654
rect 11313 253620 11329 253654
rect 10943 253512 10959 253546
rect 11313 253512 11329 253546
rect 11363 253620 11379 253654
rect 11733 253620 11749 253654
rect 11363 253512 11379 253546
rect 11733 253512 11749 253546
rect 11783 253620 11799 253654
rect 12153 253620 12169 253654
rect 11783 253512 11799 253546
rect 12153 253512 12169 253546
rect 12203 253620 12219 253654
rect 12573 253620 12589 253654
rect 12203 253512 12219 253546
rect 12573 253512 12589 253546
rect 12623 253620 12639 253654
rect 12993 253620 13009 253654
rect 12623 253512 12639 253546
rect 12993 253512 13009 253546
rect 13043 253620 13059 253654
rect 13413 253620 13429 253654
rect 13043 253512 13059 253546
rect 13413 253512 13429 253546
rect 13463 253620 13479 253654
rect 13833 253620 13849 253654
rect 13463 253512 13479 253546
rect 13833 253512 13849 253546
rect 13883 253620 13899 253654
rect 14253 253620 14269 253654
rect 13883 253512 13899 253546
rect 14253 253512 14269 253546
rect 14303 253620 14319 253654
rect 14673 253620 14689 253654
rect 14303 253512 14319 253546
rect 14673 253512 14689 253546
rect 14723 253620 14739 253654
rect 15093 253620 15109 253654
rect 14723 253512 14739 253546
rect 15093 253512 15109 253546
rect 15143 253620 15159 253654
rect 15513 253620 15529 253654
rect 15143 253512 15159 253546
rect 15513 253512 15529 253546
rect 15563 253620 15579 253654
rect 15933 253620 15949 253654
rect 15563 253512 15579 253546
rect 15933 253512 15949 253546
rect 15983 253620 15999 253654
rect 16353 253620 16369 253654
rect 15983 253512 15999 253546
rect 16353 253512 16369 253546
rect 16403 253620 16419 253654
rect 16773 253620 16789 253654
rect 16403 253512 16419 253546
rect 16773 253512 16789 253546
rect 16823 253620 16839 253654
rect 17193 253620 17209 253654
rect 16823 253512 16839 253546
rect 17193 253512 17209 253546
rect 17243 253620 17259 253654
rect 17613 253620 17629 253654
rect 17243 253512 17259 253546
rect 17613 253512 17629 253546
rect 17663 253620 17679 253654
rect 18033 253620 18049 253654
rect 17663 253512 17679 253546
rect 18033 253512 18049 253546
rect 18083 253620 18099 253654
rect 18453 253620 18469 253654
rect 18083 253512 18099 253546
rect 18453 253512 18469 253546
rect 18503 253620 18519 253654
rect 18873 253620 18889 253654
rect 18503 253512 18519 253546
rect 18873 253512 18889 253546
rect 18923 253620 18939 253654
rect 19293 253620 19309 253654
rect 18923 253512 18939 253546
rect 19293 253512 19309 253546
rect 19343 253620 19359 253654
rect 19713 253620 19729 253654
rect 19343 253512 19359 253546
rect 19713 253512 19729 253546
rect 19763 253620 19779 253654
rect 20133 253620 20149 253654
rect 19763 253512 19779 253546
rect 20133 253512 20149 253546
rect 20183 253620 20199 253654
rect 20553 253620 20569 253654
rect 20183 253512 20199 253546
rect 20553 253512 20569 253546
rect 20603 253620 20619 253654
rect 20973 253620 20989 253654
rect 20603 253512 20619 253546
rect 20973 253512 20989 253546
rect 21023 253620 21039 253654
rect 21393 253620 21409 253654
rect 21023 253512 21039 253546
rect 21393 253512 21409 253546
rect 21443 253620 21459 253654
rect 21813 253620 21829 253654
rect 21443 253512 21459 253546
rect 21813 253512 21829 253546
rect 21863 253620 21879 253654
rect 22233 253620 22249 253654
rect 21863 253512 21879 253546
rect 22233 253512 22249 253546
rect 22283 253620 22299 253654
rect 22653 253620 22669 253654
rect 22283 253512 22299 253546
rect 22653 253512 22669 253546
rect 22703 253620 22719 253654
rect 23073 253620 23089 253654
rect 22703 253512 22719 253546
rect 23073 253512 23089 253546
rect 23123 253620 23139 253654
rect 23493 253620 23509 253654
rect 23123 253512 23139 253546
rect 23493 253512 23509 253546
rect 23543 253620 23559 253654
rect 23913 253620 23929 253654
rect 23543 253512 23559 253546
rect 23913 253512 23929 253546
rect 23963 253620 23979 253654
rect 24333 253620 24349 253654
rect 23963 253512 23979 253546
rect 24333 253512 24349 253546
rect 24383 253620 24399 253654
rect 24753 253620 24769 253654
rect 24383 253512 24399 253546
rect 24753 253512 24769 253546
rect 24803 253620 24819 253654
rect 25173 253620 25189 253654
rect 24803 253512 24819 253546
rect 25173 253512 25189 253546
rect 25223 253620 25239 253654
rect 25593 253620 25609 253654
rect 25223 253512 25239 253546
rect 25593 253512 25609 253546
rect 25643 253620 25659 253654
rect 26013 253620 26029 253654
rect 25643 253512 25659 253546
rect 26013 253512 26029 253546
rect 26063 253620 26079 253654
rect 26433 253620 26449 253654
rect 26063 253512 26079 253546
rect 26433 253512 26449 253546
rect 26483 253620 26499 253654
rect 26853 253620 26869 253654
rect 26483 253512 26499 253546
rect 26853 253512 26869 253546
rect 26903 253620 26919 253654
rect 27273 253620 27289 253654
rect 26903 253512 26919 253546
rect 27273 253512 27289 253546
rect 27323 253620 27339 253654
rect 27323 253512 27339 253546
rect -4049 253453 -4015 253469
rect -4049 252661 -4015 252677
rect -3953 253453 -3919 253469
rect -3953 252661 -3919 252677
rect -3839 253453 -3805 253469
rect -3839 252661 -3805 252677
rect -3743 253453 -3709 253469
rect -3743 252661 -3709 252677
rect -3629 253453 -3595 253469
rect -3629 252661 -3595 252677
rect -3533 253453 -3499 253469
rect -3533 252661 -3499 252677
rect -3419 253453 -3385 253469
rect -3419 252661 -3385 252677
rect -3323 253453 -3289 253469
rect -3323 252661 -3289 252677
rect -3209 253453 -3175 253469
rect -3209 252661 -3175 252677
rect -3113 253453 -3079 253469
rect -3113 252661 -3079 252677
rect -2999 253453 -2965 253469
rect -2999 252661 -2965 252677
rect -2903 253453 -2869 253469
rect -2903 252661 -2869 252677
rect -2789 253453 -2755 253469
rect -2789 252661 -2755 252677
rect -2693 253453 -2659 253469
rect -2693 252661 -2659 252677
rect -2579 253453 -2545 253469
rect -2579 252661 -2545 252677
rect -2483 253453 -2449 253469
rect -2483 252661 -2449 252677
rect -2369 253453 -2335 253469
rect -2369 252661 -2335 252677
rect -2273 253453 -2239 253469
rect -2273 252661 -2239 252677
rect -2159 253453 -2125 253469
rect -2159 252661 -2125 252677
rect -2063 253453 -2029 253469
rect -2063 252661 -2029 252677
rect -1949 253453 -1915 253469
rect -1949 252661 -1915 252677
rect -1853 253453 -1819 253469
rect -1853 252661 -1819 252677
rect -1739 253453 -1705 253469
rect -1739 252661 -1705 252677
rect -1643 253453 -1609 253469
rect -1643 252661 -1609 252677
rect -1529 253453 -1495 253469
rect -1529 252661 -1495 252677
rect -1433 253453 -1399 253469
rect -1433 252661 -1399 252677
rect -1319 253453 -1285 253469
rect -1319 252661 -1285 252677
rect -1223 253453 -1189 253469
rect -1223 252661 -1189 252677
rect -1109 253453 -1075 253469
rect -1109 252661 -1075 252677
rect -1013 253453 -979 253469
rect -1013 252661 -979 252677
rect -899 253453 -865 253469
rect -899 252661 -865 252677
rect -803 253453 -769 253469
rect -803 252661 -769 252677
rect -689 253453 -655 253469
rect -689 252661 -655 252677
rect -593 253453 -559 253469
rect -593 252661 -559 252677
rect -479 253453 -445 253469
rect -479 252661 -445 252677
rect -383 253453 -349 253469
rect -383 252661 -349 252677
rect -269 253453 -235 253469
rect -269 252661 -235 252677
rect -173 253453 -139 253469
rect -173 252661 -139 252677
rect -59 253453 -25 253469
rect -59 252661 -25 252677
rect 37 253453 71 253469
rect 37 252661 71 252677
rect 151 253453 185 253469
rect 151 252661 185 252677
rect 247 253453 281 253469
rect 247 252661 281 252677
rect 361 253453 395 253469
rect 361 252661 395 252677
rect 457 253453 491 253469
rect 457 252661 491 252677
rect 571 253453 605 253469
rect 571 252661 605 252677
rect 667 253453 701 253469
rect 667 252661 701 252677
rect 781 253453 815 253469
rect 781 252661 815 252677
rect 877 253453 911 253469
rect 877 252661 911 252677
rect 991 253453 1025 253469
rect 991 252661 1025 252677
rect 1087 253453 1121 253469
rect 1087 252661 1121 252677
rect 1201 253453 1235 253469
rect 1201 252661 1235 252677
rect 1297 253453 1331 253469
rect 1297 252661 1331 252677
rect 1411 253453 1445 253469
rect 1411 252661 1445 252677
rect 1507 253453 1541 253469
rect 1507 252661 1541 252677
rect 1621 253453 1655 253469
rect 1621 252661 1655 252677
rect 1717 253453 1751 253469
rect 1717 252661 1751 252677
rect 1831 253453 1865 253469
rect 1831 252661 1865 252677
rect 1927 253453 1961 253469
rect 1927 252661 1961 252677
rect 2041 253453 2075 253469
rect 2041 252661 2075 252677
rect 2137 253453 2171 253469
rect 2137 252661 2171 252677
rect 2251 253453 2285 253469
rect 2251 252661 2285 252677
rect 2347 253453 2381 253469
rect 2347 252661 2381 252677
rect 2461 253453 2495 253469
rect 2461 252661 2495 252677
rect 2557 253453 2591 253469
rect 2557 252661 2591 252677
rect 2671 253453 2705 253469
rect 2671 252661 2705 252677
rect 2767 253453 2801 253469
rect 2767 252661 2801 252677
rect 2881 253453 2915 253469
rect 2881 252661 2915 252677
rect 2977 253453 3011 253469
rect 2977 252661 3011 252677
rect 3091 253453 3125 253469
rect 3091 252661 3125 252677
rect 3187 253453 3221 253469
rect 3187 252661 3221 252677
rect 3301 253453 3335 253469
rect 3301 252661 3335 252677
rect 3397 253453 3431 253469
rect 3397 252661 3431 252677
rect 3511 253453 3545 253469
rect 3511 252661 3545 252677
rect 3607 253453 3641 253469
rect 3607 252661 3641 252677
rect 3721 253453 3755 253469
rect 3721 252661 3755 252677
rect 3817 253453 3851 253469
rect 3817 252661 3851 252677
rect 3931 253453 3965 253469
rect 3931 252661 3965 252677
rect 4027 253453 4061 253469
rect 4027 252661 4061 252677
rect 4141 253453 4175 253469
rect 4141 252661 4175 252677
rect 4237 253453 4271 253469
rect 4237 252661 4271 252677
rect 4351 253453 4385 253469
rect 4351 252661 4385 252677
rect 4447 253453 4481 253469
rect 4447 252661 4481 252677
rect 4561 253453 4595 253469
rect 4561 252661 4595 252677
rect 4657 253453 4691 253469
rect 4657 252661 4691 252677
rect 4771 253453 4805 253469
rect 4771 252661 4805 252677
rect 4867 253453 4901 253469
rect 4867 252661 4901 252677
rect 4981 253453 5015 253469
rect 4981 252661 5015 252677
rect 5077 253453 5111 253469
rect 5077 252661 5111 252677
rect 5191 253453 5225 253469
rect 5191 252661 5225 252677
rect 5287 253453 5321 253469
rect 5287 252661 5321 252677
rect 5401 253453 5435 253469
rect 5401 252661 5435 252677
rect 5497 253453 5531 253469
rect 5497 252661 5531 252677
rect 5611 253453 5645 253469
rect 5611 252661 5645 252677
rect 5707 253453 5741 253469
rect 5707 252661 5741 252677
rect 5821 253453 5855 253469
rect 5821 252661 5855 252677
rect 5917 253453 5951 253469
rect 5917 252661 5951 252677
rect 6031 253453 6065 253469
rect 6031 252661 6065 252677
rect 6127 253453 6161 253469
rect 6127 252661 6161 252677
rect 6241 253453 6275 253469
rect 6241 252661 6275 252677
rect 6337 253453 6371 253469
rect 6337 252661 6371 252677
rect 6451 253453 6485 253469
rect 6451 252661 6485 252677
rect 6547 253453 6581 253469
rect 6547 252661 6581 252677
rect 6661 253453 6695 253469
rect 6661 252661 6695 252677
rect 6757 253453 6791 253469
rect 6757 252661 6791 252677
rect 6871 253453 6905 253469
rect 6871 252661 6905 252677
rect 6967 253453 7001 253469
rect 6967 252661 7001 252677
rect 7081 253453 7115 253469
rect 7081 252661 7115 252677
rect 7177 253453 7211 253469
rect 7177 252661 7211 252677
rect 7291 253453 7325 253469
rect 7291 252661 7325 252677
rect 7387 253453 7421 253469
rect 7387 252661 7421 252677
rect 7501 253453 7535 253469
rect 7501 252661 7535 252677
rect 7597 253453 7631 253469
rect 7597 252661 7631 252677
rect 7711 253453 7745 253469
rect 7711 252661 7745 252677
rect 7807 253453 7841 253469
rect 7807 252661 7841 252677
rect 7921 253453 7955 253469
rect 7921 252661 7955 252677
rect 8017 253453 8051 253469
rect 8017 252661 8051 252677
rect 8131 253453 8165 253469
rect 8131 252661 8165 252677
rect 8227 253453 8261 253469
rect 8227 252661 8261 252677
rect 8341 253453 8375 253469
rect 8341 252661 8375 252677
rect 8437 253453 8471 253469
rect 8437 252661 8471 252677
rect 8551 253453 8585 253469
rect 8551 252661 8585 252677
rect 8647 253453 8681 253469
rect 8647 252661 8681 252677
rect 8761 253453 8795 253469
rect 8761 252661 8795 252677
rect 8857 253453 8891 253469
rect 8857 252661 8891 252677
rect 8971 253453 9005 253469
rect 8971 252661 9005 252677
rect 9067 253453 9101 253469
rect 9067 252661 9101 252677
rect 9181 253453 9215 253469
rect 9181 252661 9215 252677
rect 9277 253453 9311 253469
rect 9277 252661 9311 252677
rect 9391 253453 9425 253469
rect 9391 252661 9425 252677
rect 9487 253453 9521 253469
rect 9487 252661 9521 252677
rect 9601 253453 9635 253469
rect 9601 252661 9635 252677
rect 9697 253453 9731 253469
rect 9697 252661 9731 252677
rect 9811 253453 9845 253469
rect 9811 252661 9845 252677
rect 9907 253453 9941 253469
rect 9907 252661 9941 252677
rect 10021 253453 10055 253469
rect 10021 252661 10055 252677
rect 10117 253453 10151 253469
rect 10117 252661 10151 252677
rect 10231 253453 10265 253469
rect 10231 252661 10265 252677
rect 10327 253453 10361 253469
rect 10327 252661 10361 252677
rect 10441 253453 10475 253469
rect 10441 252661 10475 252677
rect 10537 253453 10571 253469
rect 10537 252661 10571 252677
rect 10651 253453 10685 253469
rect 10651 252661 10685 252677
rect 10747 253453 10781 253469
rect 10747 252661 10781 252677
rect 10861 253453 10895 253469
rect 10861 252661 10895 252677
rect 10957 253453 10991 253469
rect 10957 252661 10991 252677
rect 11071 253453 11105 253469
rect 11071 252661 11105 252677
rect 11167 253453 11201 253469
rect 11167 252661 11201 252677
rect 11281 253453 11315 253469
rect 11281 252661 11315 252677
rect 11377 253453 11411 253469
rect 11377 252661 11411 252677
rect 11491 253453 11525 253469
rect 11491 252661 11525 252677
rect 11587 253453 11621 253469
rect 11587 252661 11621 252677
rect 11701 253453 11735 253469
rect 11701 252661 11735 252677
rect 11797 253453 11831 253469
rect 11797 252661 11831 252677
rect 11911 253453 11945 253469
rect 11911 252661 11945 252677
rect 12007 253453 12041 253469
rect 12007 252661 12041 252677
rect 12121 253453 12155 253469
rect 12121 252661 12155 252677
rect 12217 253453 12251 253469
rect 12217 252661 12251 252677
rect 12331 253453 12365 253469
rect 12331 252661 12365 252677
rect 12427 253453 12461 253469
rect 12427 252661 12461 252677
rect 12541 253453 12575 253469
rect 12541 252661 12575 252677
rect 12637 253453 12671 253469
rect 12637 252661 12671 252677
rect 12751 253453 12785 253469
rect 12751 252661 12785 252677
rect 12847 253453 12881 253469
rect 12847 252661 12881 252677
rect 12961 253453 12995 253469
rect 12961 252661 12995 252677
rect 13057 253453 13091 253469
rect 13057 252661 13091 252677
rect 13171 253453 13205 253469
rect 13171 252661 13205 252677
rect 13267 253453 13301 253469
rect 13267 252661 13301 252677
rect 13381 253453 13415 253469
rect 13381 252661 13415 252677
rect 13477 253453 13511 253469
rect 13477 252661 13511 252677
rect 13591 253453 13625 253469
rect 13591 252661 13625 252677
rect 13687 253453 13721 253469
rect 13687 252661 13721 252677
rect 13801 253453 13835 253469
rect 13801 252661 13835 252677
rect 13897 253453 13931 253469
rect 13897 252661 13931 252677
rect 14011 253453 14045 253469
rect 14011 252661 14045 252677
rect 14107 253453 14141 253469
rect 14107 252661 14141 252677
rect 14221 253453 14255 253469
rect 14221 252661 14255 252677
rect 14317 253453 14351 253469
rect 14317 252661 14351 252677
rect 14431 253453 14465 253469
rect 14431 252661 14465 252677
rect 14527 253453 14561 253469
rect 14527 252661 14561 252677
rect 14641 253453 14675 253469
rect 14641 252661 14675 252677
rect 14737 253453 14771 253469
rect 14737 252661 14771 252677
rect 14851 253453 14885 253469
rect 14851 252661 14885 252677
rect 14947 253453 14981 253469
rect 14947 252661 14981 252677
rect 15061 253453 15095 253469
rect 15061 252661 15095 252677
rect 15157 253453 15191 253469
rect 15157 252661 15191 252677
rect 15271 253453 15305 253469
rect 15271 252661 15305 252677
rect 15367 253453 15401 253469
rect 15367 252661 15401 252677
rect 15481 253453 15515 253469
rect 15481 252661 15515 252677
rect 15577 253453 15611 253469
rect 15577 252661 15611 252677
rect 15691 253453 15725 253469
rect 15691 252661 15725 252677
rect 15787 253453 15821 253469
rect 15787 252661 15821 252677
rect 15901 253453 15935 253469
rect 15901 252661 15935 252677
rect 15997 253453 16031 253469
rect 15997 252661 16031 252677
rect 16111 253453 16145 253469
rect 16111 252661 16145 252677
rect 16207 253453 16241 253469
rect 16207 252661 16241 252677
rect 16321 253453 16355 253469
rect 16321 252661 16355 252677
rect 16417 253453 16451 253469
rect 16417 252661 16451 252677
rect 16531 253453 16565 253469
rect 16531 252661 16565 252677
rect 16627 253453 16661 253469
rect 16627 252661 16661 252677
rect 16741 253453 16775 253469
rect 16741 252661 16775 252677
rect 16837 253453 16871 253469
rect 16837 252661 16871 252677
rect 16951 253453 16985 253469
rect 16951 252661 16985 252677
rect 17047 253453 17081 253469
rect 17047 252661 17081 252677
rect 17161 253453 17195 253469
rect 17161 252661 17195 252677
rect 17257 253453 17291 253469
rect 17257 252661 17291 252677
rect 17371 253453 17405 253469
rect 17371 252661 17405 252677
rect 17467 253453 17501 253469
rect 17467 252661 17501 252677
rect 17581 253453 17615 253469
rect 17581 252661 17615 252677
rect 17677 253453 17711 253469
rect 17677 252661 17711 252677
rect 17791 253453 17825 253469
rect 17791 252661 17825 252677
rect 17887 253453 17921 253469
rect 17887 252661 17921 252677
rect 18001 253453 18035 253469
rect 18001 252661 18035 252677
rect 18097 253453 18131 253469
rect 18097 252661 18131 252677
rect 18211 253453 18245 253469
rect 18211 252661 18245 252677
rect 18307 253453 18341 253469
rect 18307 252661 18341 252677
rect 18421 253453 18455 253469
rect 18421 252661 18455 252677
rect 18517 253453 18551 253469
rect 18517 252661 18551 252677
rect 18631 253453 18665 253469
rect 18631 252661 18665 252677
rect 18727 253453 18761 253469
rect 18727 252661 18761 252677
rect 18841 253453 18875 253469
rect 18841 252661 18875 252677
rect 18937 253453 18971 253469
rect 18937 252661 18971 252677
rect 19051 253453 19085 253469
rect 19051 252661 19085 252677
rect 19147 253453 19181 253469
rect 19147 252661 19181 252677
rect 19261 253453 19295 253469
rect 19261 252661 19295 252677
rect 19357 253453 19391 253469
rect 19357 252661 19391 252677
rect 19471 253453 19505 253469
rect 19471 252661 19505 252677
rect 19567 253453 19601 253469
rect 19567 252661 19601 252677
rect 19681 253453 19715 253469
rect 19681 252661 19715 252677
rect 19777 253453 19811 253469
rect 19777 252661 19811 252677
rect 19891 253453 19925 253469
rect 19891 252661 19925 252677
rect 19987 253453 20021 253469
rect 19987 252661 20021 252677
rect 20101 253453 20135 253469
rect 20101 252661 20135 252677
rect 20197 253453 20231 253469
rect 20197 252661 20231 252677
rect 20311 253453 20345 253469
rect 20311 252661 20345 252677
rect 20407 253453 20441 253469
rect 20407 252661 20441 252677
rect 20521 253453 20555 253469
rect 20521 252661 20555 252677
rect 20617 253453 20651 253469
rect 20617 252661 20651 252677
rect 20731 253453 20765 253469
rect 20731 252661 20765 252677
rect 20827 253453 20861 253469
rect 20827 252661 20861 252677
rect 20941 253453 20975 253469
rect 20941 252661 20975 252677
rect 21037 253453 21071 253469
rect 21037 252661 21071 252677
rect 21151 253453 21185 253469
rect 21151 252661 21185 252677
rect 21247 253453 21281 253469
rect 21247 252661 21281 252677
rect 21361 253453 21395 253469
rect 21361 252661 21395 252677
rect 21457 253453 21491 253469
rect 21457 252661 21491 252677
rect 21571 253453 21605 253469
rect 21571 252661 21605 252677
rect 21667 253453 21701 253469
rect 21667 252661 21701 252677
rect 21781 253453 21815 253469
rect 21781 252661 21815 252677
rect 21877 253453 21911 253469
rect 21877 252661 21911 252677
rect 21991 253453 22025 253469
rect 21991 252661 22025 252677
rect 22087 253453 22121 253469
rect 22087 252661 22121 252677
rect 22201 253453 22235 253469
rect 22201 252661 22235 252677
rect 22297 253453 22331 253469
rect 22297 252661 22331 252677
rect 22411 253453 22445 253469
rect 22411 252661 22445 252677
rect 22507 253453 22541 253469
rect 22507 252661 22541 252677
rect 22621 253453 22655 253469
rect 22621 252661 22655 252677
rect 22717 253453 22751 253469
rect 22717 252661 22751 252677
rect 22831 253453 22865 253469
rect 22831 252661 22865 252677
rect 22927 253453 22961 253469
rect 22927 252661 22961 252677
rect 23041 253453 23075 253469
rect 23041 252661 23075 252677
rect 23137 253453 23171 253469
rect 23137 252661 23171 252677
rect 23251 253453 23285 253469
rect 23251 252661 23285 252677
rect 23347 253453 23381 253469
rect 23347 252661 23381 252677
rect 23461 253453 23495 253469
rect 23461 252661 23495 252677
rect 23557 253453 23591 253469
rect 23557 252661 23591 252677
rect 23671 253453 23705 253469
rect 23671 252661 23705 252677
rect 23767 253453 23801 253469
rect 23767 252661 23801 252677
rect 23881 253453 23915 253469
rect 23881 252661 23915 252677
rect 23977 253453 24011 253469
rect 23977 252661 24011 252677
rect 24091 253453 24125 253469
rect 24091 252661 24125 252677
rect 24187 253453 24221 253469
rect 24187 252661 24221 252677
rect 24301 253453 24335 253469
rect 24301 252661 24335 252677
rect 24397 253453 24431 253469
rect 24397 252661 24431 252677
rect 24511 253453 24545 253469
rect 24511 252661 24545 252677
rect 24607 253453 24641 253469
rect 24607 252661 24641 252677
rect 24721 253453 24755 253469
rect 24721 252661 24755 252677
rect 24817 253453 24851 253469
rect 24817 252661 24851 252677
rect 24931 253453 24965 253469
rect 24931 252661 24965 252677
rect 25027 253453 25061 253469
rect 25027 252661 25061 252677
rect 25141 253453 25175 253469
rect 25141 252661 25175 252677
rect 25237 253453 25271 253469
rect 25237 252661 25271 252677
rect 25351 253453 25385 253469
rect 25351 252661 25385 252677
rect 25447 253453 25481 253469
rect 25447 252661 25481 252677
rect 25561 253453 25595 253469
rect 25561 252661 25595 252677
rect 25657 253453 25691 253469
rect 25657 252661 25691 252677
rect 25771 253453 25805 253469
rect 25771 252661 25805 252677
rect 25867 253453 25901 253469
rect 25867 252661 25901 252677
rect 25981 253453 26015 253469
rect 25981 252661 26015 252677
rect 26077 253453 26111 253469
rect 26077 252661 26111 252677
rect 26191 253453 26225 253469
rect 26191 252661 26225 252677
rect 26287 253453 26321 253469
rect 26287 252661 26321 252677
rect 26401 253453 26435 253469
rect 26401 252661 26435 252677
rect 26497 253453 26531 253469
rect 26497 252661 26531 252677
rect 26611 253453 26645 253469
rect 26611 252661 26645 252677
rect 26707 253453 26741 253469
rect 26707 252661 26741 252677
rect 26821 253453 26855 253469
rect 26821 252661 26855 252677
rect 26917 253453 26951 253469
rect 26917 252661 26951 252677
rect 27031 253453 27065 253469
rect 27031 252661 27065 252677
rect 27127 253453 27161 253469
rect 27127 252661 27161 252677
rect 27241 253453 27275 253469
rect 27241 252661 27275 252677
rect 27337 253453 27371 253469
rect 27337 252661 27371 252677
rect -4017 252584 -4001 252618
rect -4017 252476 -4001 252510
rect -3967 252584 -3951 252618
rect -3597 252584 -3581 252618
rect -3967 252476 -3951 252510
rect -3597 252476 -3581 252510
rect -3547 252584 -3531 252618
rect -3177 252584 -3161 252618
rect -3547 252476 -3531 252510
rect -3177 252476 -3161 252510
rect -3127 252584 -3111 252618
rect -2757 252584 -2741 252618
rect -3127 252476 -3111 252510
rect -2757 252476 -2741 252510
rect -2707 252584 -2691 252618
rect -2337 252584 -2321 252618
rect -2707 252476 -2691 252510
rect -2337 252476 -2321 252510
rect -2287 252584 -2271 252618
rect -1917 252584 -1901 252618
rect -2287 252476 -2271 252510
rect -1917 252476 -1901 252510
rect -1867 252584 -1851 252618
rect -1497 252584 -1481 252618
rect -1867 252476 -1851 252510
rect -1497 252476 -1481 252510
rect -1447 252584 -1431 252618
rect -1077 252584 -1061 252618
rect -1447 252476 -1431 252510
rect -1077 252476 -1061 252510
rect -1027 252584 -1011 252618
rect -657 252584 -641 252618
rect -1027 252476 -1011 252510
rect -657 252476 -641 252510
rect -607 252584 -591 252618
rect -237 252584 -221 252618
rect -607 252476 -591 252510
rect -237 252476 -221 252510
rect -187 252584 -171 252618
rect 183 252584 199 252618
rect -187 252476 -171 252510
rect 183 252476 199 252510
rect 233 252584 249 252618
rect 603 252584 619 252618
rect 233 252476 249 252510
rect 603 252476 619 252510
rect 653 252584 669 252618
rect 1023 252584 1039 252618
rect 653 252476 669 252510
rect 1023 252476 1039 252510
rect 1073 252584 1089 252618
rect 1443 252584 1459 252618
rect 1073 252476 1089 252510
rect 1443 252476 1459 252510
rect 1493 252584 1509 252618
rect 1863 252584 1879 252618
rect 1493 252476 1509 252510
rect 1863 252476 1879 252510
rect 1913 252584 1929 252618
rect 2283 252584 2299 252618
rect 1913 252476 1929 252510
rect 2283 252476 2299 252510
rect 2333 252584 2349 252618
rect 2703 252584 2719 252618
rect 2333 252476 2349 252510
rect 2703 252476 2719 252510
rect 2753 252584 2769 252618
rect 3123 252584 3139 252618
rect 2753 252476 2769 252510
rect 3123 252476 3139 252510
rect 3173 252584 3189 252618
rect 3543 252584 3559 252618
rect 3173 252476 3189 252510
rect 3543 252476 3559 252510
rect 3593 252584 3609 252618
rect 3963 252584 3979 252618
rect 3593 252476 3609 252510
rect 3963 252476 3979 252510
rect 4013 252584 4029 252618
rect 4383 252584 4399 252618
rect 4013 252476 4029 252510
rect 4383 252476 4399 252510
rect 4433 252584 4449 252618
rect 4803 252584 4819 252618
rect 4433 252476 4449 252510
rect 4803 252476 4819 252510
rect 4853 252584 4869 252618
rect 5223 252584 5239 252618
rect 4853 252476 4869 252510
rect 5223 252476 5239 252510
rect 5273 252584 5289 252618
rect 5643 252584 5659 252618
rect 5273 252476 5289 252510
rect 5643 252476 5659 252510
rect 5693 252584 5709 252618
rect 6063 252584 6079 252618
rect 5693 252476 5709 252510
rect 6063 252476 6079 252510
rect 6113 252584 6129 252618
rect 6483 252584 6499 252618
rect 6113 252476 6129 252510
rect 6483 252476 6499 252510
rect 6533 252584 6549 252618
rect 6903 252584 6919 252618
rect 6533 252476 6549 252510
rect 6903 252476 6919 252510
rect 6953 252584 6969 252618
rect 7323 252584 7339 252618
rect 6953 252476 6969 252510
rect 7323 252476 7339 252510
rect 7373 252584 7389 252618
rect 7743 252584 7759 252618
rect 7373 252476 7389 252510
rect 7743 252476 7759 252510
rect 7793 252584 7809 252618
rect 8163 252584 8179 252618
rect 7793 252476 7809 252510
rect 8163 252476 8179 252510
rect 8213 252584 8229 252618
rect 8583 252584 8599 252618
rect 8213 252476 8229 252510
rect 8583 252476 8599 252510
rect 8633 252584 8649 252618
rect 9003 252584 9019 252618
rect 8633 252476 8649 252510
rect 9003 252476 9019 252510
rect 9053 252584 9069 252618
rect 9423 252584 9439 252618
rect 9053 252476 9069 252510
rect 9423 252476 9439 252510
rect 9473 252584 9489 252618
rect 9843 252584 9859 252618
rect 9473 252476 9489 252510
rect 9843 252476 9859 252510
rect 9893 252584 9909 252618
rect 10263 252584 10279 252618
rect 9893 252476 9909 252510
rect 10263 252476 10279 252510
rect 10313 252584 10329 252618
rect 10683 252584 10699 252618
rect 10313 252476 10329 252510
rect 10683 252476 10699 252510
rect 10733 252584 10749 252618
rect 11103 252584 11119 252618
rect 10733 252476 10749 252510
rect 11103 252476 11119 252510
rect 11153 252584 11169 252618
rect 11523 252584 11539 252618
rect 11153 252476 11169 252510
rect 11523 252476 11539 252510
rect 11573 252584 11589 252618
rect 11943 252584 11959 252618
rect 11573 252476 11589 252510
rect 11943 252476 11959 252510
rect 11993 252584 12009 252618
rect 12363 252584 12379 252618
rect 11993 252476 12009 252510
rect 12363 252476 12379 252510
rect 12413 252584 12429 252618
rect 12783 252584 12799 252618
rect 12413 252476 12429 252510
rect 12783 252476 12799 252510
rect 12833 252584 12849 252618
rect 13203 252584 13219 252618
rect 12833 252476 12849 252510
rect 13203 252476 13219 252510
rect 13253 252584 13269 252618
rect 13623 252584 13639 252618
rect 13253 252476 13269 252510
rect 13623 252476 13639 252510
rect 13673 252584 13689 252618
rect 14043 252584 14059 252618
rect 13673 252476 13689 252510
rect 14043 252476 14059 252510
rect 14093 252584 14109 252618
rect 14463 252584 14479 252618
rect 14093 252476 14109 252510
rect 14463 252476 14479 252510
rect 14513 252584 14529 252618
rect 14883 252584 14899 252618
rect 14513 252476 14529 252510
rect 14883 252476 14899 252510
rect 14933 252584 14949 252618
rect 15303 252584 15319 252618
rect 14933 252476 14949 252510
rect 15303 252476 15319 252510
rect 15353 252584 15369 252618
rect 15723 252584 15739 252618
rect 15353 252476 15369 252510
rect 15723 252476 15739 252510
rect 15773 252584 15789 252618
rect 16143 252584 16159 252618
rect 15773 252476 15789 252510
rect 16143 252476 16159 252510
rect 16193 252584 16209 252618
rect 16563 252584 16579 252618
rect 16193 252476 16209 252510
rect 16563 252476 16579 252510
rect 16613 252584 16629 252618
rect 16983 252584 16999 252618
rect 16613 252476 16629 252510
rect 16983 252476 16999 252510
rect 17033 252584 17049 252618
rect 17403 252584 17419 252618
rect 17033 252476 17049 252510
rect 17403 252476 17419 252510
rect 17453 252584 17469 252618
rect 17823 252584 17839 252618
rect 17453 252476 17469 252510
rect 17823 252476 17839 252510
rect 17873 252584 17889 252618
rect 18243 252584 18259 252618
rect 17873 252476 17889 252510
rect 18243 252476 18259 252510
rect 18293 252584 18309 252618
rect 18663 252584 18679 252618
rect 18293 252476 18309 252510
rect 18663 252476 18679 252510
rect 18713 252584 18729 252618
rect 19083 252584 19099 252618
rect 18713 252476 18729 252510
rect 19083 252476 19099 252510
rect 19133 252584 19149 252618
rect 19503 252584 19519 252618
rect 19133 252476 19149 252510
rect 19503 252476 19519 252510
rect 19553 252584 19569 252618
rect 19923 252584 19939 252618
rect 19553 252476 19569 252510
rect 19923 252476 19939 252510
rect 19973 252584 19989 252618
rect 20343 252584 20359 252618
rect 19973 252476 19989 252510
rect 20343 252476 20359 252510
rect 20393 252584 20409 252618
rect 20763 252584 20779 252618
rect 20393 252476 20409 252510
rect 20763 252476 20779 252510
rect 20813 252584 20829 252618
rect 21183 252584 21199 252618
rect 20813 252476 20829 252510
rect 21183 252476 21199 252510
rect 21233 252584 21249 252618
rect 21603 252584 21619 252618
rect 21233 252476 21249 252510
rect 21603 252476 21619 252510
rect 21653 252584 21669 252618
rect 22023 252584 22039 252618
rect 21653 252476 21669 252510
rect 22023 252476 22039 252510
rect 22073 252584 22089 252618
rect 22443 252584 22459 252618
rect 22073 252476 22089 252510
rect 22443 252476 22459 252510
rect 22493 252584 22509 252618
rect 22863 252584 22879 252618
rect 22493 252476 22509 252510
rect 22863 252476 22879 252510
rect 22913 252584 22929 252618
rect 23283 252584 23299 252618
rect 22913 252476 22929 252510
rect 23283 252476 23299 252510
rect 23333 252584 23349 252618
rect 23703 252584 23719 252618
rect 23333 252476 23349 252510
rect 23703 252476 23719 252510
rect 23753 252584 23769 252618
rect 24123 252584 24139 252618
rect 23753 252476 23769 252510
rect 24123 252476 24139 252510
rect 24173 252584 24189 252618
rect 24543 252584 24559 252618
rect 24173 252476 24189 252510
rect 24543 252476 24559 252510
rect 24593 252584 24609 252618
rect 24963 252584 24979 252618
rect 24593 252476 24609 252510
rect 24963 252476 24979 252510
rect 25013 252584 25029 252618
rect 25383 252584 25399 252618
rect 25013 252476 25029 252510
rect 25383 252476 25399 252510
rect 25433 252584 25449 252618
rect 25803 252584 25819 252618
rect 25433 252476 25449 252510
rect 25803 252476 25819 252510
rect 25853 252584 25869 252618
rect 26223 252584 26239 252618
rect 25853 252476 25869 252510
rect 26223 252476 26239 252510
rect 26273 252584 26289 252618
rect 26643 252584 26659 252618
rect 26273 252476 26289 252510
rect 26643 252476 26659 252510
rect 26693 252584 26709 252618
rect 27063 252584 27079 252618
rect 26693 252476 26709 252510
rect 27063 252476 27079 252510
rect 27113 252584 27129 252618
rect 27113 252476 27129 252510
rect -4049 252417 -4015 252433
rect -4049 251625 -4015 251641
rect -3953 252417 -3919 252433
rect -3953 251625 -3919 251641
rect -3839 252417 -3805 252433
rect -3839 251625 -3805 251641
rect -3743 252417 -3709 252433
rect -3743 251625 -3709 251641
rect -3629 252417 -3595 252433
rect -3629 251625 -3595 251641
rect -3533 252417 -3499 252433
rect -3533 251625 -3499 251641
rect -3419 252417 -3385 252433
rect -3419 251625 -3385 251641
rect -3323 252417 -3289 252433
rect -3323 251625 -3289 251641
rect -3209 252417 -3175 252433
rect -3209 251625 -3175 251641
rect -3113 252417 -3079 252433
rect -3113 251625 -3079 251641
rect -2999 252417 -2965 252433
rect -2999 251625 -2965 251641
rect -2903 252417 -2869 252433
rect -2903 251625 -2869 251641
rect -2789 252417 -2755 252433
rect -2789 251625 -2755 251641
rect -2693 252417 -2659 252433
rect -2693 251625 -2659 251641
rect -2579 252417 -2545 252433
rect -2579 251625 -2545 251641
rect -2483 252417 -2449 252433
rect -2483 251625 -2449 251641
rect -2369 252417 -2335 252433
rect -2369 251625 -2335 251641
rect -2273 252417 -2239 252433
rect -2273 251625 -2239 251641
rect -2159 252417 -2125 252433
rect -2159 251625 -2125 251641
rect -2063 252417 -2029 252433
rect -2063 251625 -2029 251641
rect -1949 252417 -1915 252433
rect -1949 251625 -1915 251641
rect -1853 252417 -1819 252433
rect -1853 251625 -1819 251641
rect -1739 252417 -1705 252433
rect -1739 251625 -1705 251641
rect -1643 252417 -1609 252433
rect -1643 251625 -1609 251641
rect -1529 252417 -1495 252433
rect -1529 251625 -1495 251641
rect -1433 252417 -1399 252433
rect -1433 251625 -1399 251641
rect -1319 252417 -1285 252433
rect -1319 251625 -1285 251641
rect -1223 252417 -1189 252433
rect -1223 251625 -1189 251641
rect -1109 252417 -1075 252433
rect -1109 251625 -1075 251641
rect -1013 252417 -979 252433
rect -1013 251625 -979 251641
rect -899 252417 -865 252433
rect -899 251625 -865 251641
rect -803 252417 -769 252433
rect -803 251625 -769 251641
rect -689 252417 -655 252433
rect -689 251625 -655 251641
rect -593 252417 -559 252433
rect -593 251625 -559 251641
rect -479 252417 -445 252433
rect -479 251625 -445 251641
rect -383 252417 -349 252433
rect -383 251625 -349 251641
rect -269 252417 -235 252433
rect -269 251625 -235 251641
rect -173 252417 -139 252433
rect -173 251625 -139 251641
rect -59 252417 -25 252433
rect -59 251625 -25 251641
rect 37 252417 71 252433
rect 37 251625 71 251641
rect 151 252417 185 252433
rect 151 251625 185 251641
rect 247 252417 281 252433
rect 247 251625 281 251641
rect 361 252417 395 252433
rect 361 251625 395 251641
rect 457 252417 491 252433
rect 457 251625 491 251641
rect 571 252417 605 252433
rect 571 251625 605 251641
rect 667 252417 701 252433
rect 667 251625 701 251641
rect 781 252417 815 252433
rect 781 251625 815 251641
rect 877 252417 911 252433
rect 877 251625 911 251641
rect 991 252417 1025 252433
rect 991 251625 1025 251641
rect 1087 252417 1121 252433
rect 1087 251625 1121 251641
rect 1201 252417 1235 252433
rect 1201 251625 1235 251641
rect 1297 252417 1331 252433
rect 1297 251625 1331 251641
rect 1411 252417 1445 252433
rect 1411 251625 1445 251641
rect 1507 252417 1541 252433
rect 1507 251625 1541 251641
rect 1621 252417 1655 252433
rect 1621 251625 1655 251641
rect 1717 252417 1751 252433
rect 1717 251625 1751 251641
rect 1831 252417 1865 252433
rect 1831 251625 1865 251641
rect 1927 252417 1961 252433
rect 1927 251625 1961 251641
rect 2041 252417 2075 252433
rect 2041 251625 2075 251641
rect 2137 252417 2171 252433
rect 2137 251625 2171 251641
rect 2251 252417 2285 252433
rect 2251 251625 2285 251641
rect 2347 252417 2381 252433
rect 2347 251625 2381 251641
rect 2461 252417 2495 252433
rect 2461 251625 2495 251641
rect 2557 252417 2591 252433
rect 2557 251625 2591 251641
rect 2671 252417 2705 252433
rect 2671 251625 2705 251641
rect 2767 252417 2801 252433
rect 2767 251625 2801 251641
rect 2881 252417 2915 252433
rect 2881 251625 2915 251641
rect 2977 252417 3011 252433
rect 2977 251625 3011 251641
rect 3091 252417 3125 252433
rect 3091 251625 3125 251641
rect 3187 252417 3221 252433
rect 3187 251625 3221 251641
rect 3301 252417 3335 252433
rect 3301 251625 3335 251641
rect 3397 252417 3431 252433
rect 3397 251625 3431 251641
rect 3511 252417 3545 252433
rect 3511 251625 3545 251641
rect 3607 252417 3641 252433
rect 3607 251625 3641 251641
rect 3721 252417 3755 252433
rect 3721 251625 3755 251641
rect 3817 252417 3851 252433
rect 3817 251625 3851 251641
rect 3931 252417 3965 252433
rect 3931 251625 3965 251641
rect 4027 252417 4061 252433
rect 4027 251625 4061 251641
rect 4141 252417 4175 252433
rect 4141 251625 4175 251641
rect 4237 252417 4271 252433
rect 4237 251625 4271 251641
rect 4351 252417 4385 252433
rect 4351 251625 4385 251641
rect 4447 252417 4481 252433
rect 4447 251625 4481 251641
rect 4561 252417 4595 252433
rect 4561 251625 4595 251641
rect 4657 252417 4691 252433
rect 4657 251625 4691 251641
rect 4771 252417 4805 252433
rect 4771 251625 4805 251641
rect 4867 252417 4901 252433
rect 4867 251625 4901 251641
rect 4981 252417 5015 252433
rect 4981 251625 5015 251641
rect 5077 252417 5111 252433
rect 5077 251625 5111 251641
rect 5191 252417 5225 252433
rect 5191 251625 5225 251641
rect 5287 252417 5321 252433
rect 5287 251625 5321 251641
rect 5401 252417 5435 252433
rect 5401 251625 5435 251641
rect 5497 252417 5531 252433
rect 5497 251625 5531 251641
rect 5611 252417 5645 252433
rect 5611 251625 5645 251641
rect 5707 252417 5741 252433
rect 5707 251625 5741 251641
rect 5821 252417 5855 252433
rect 5821 251625 5855 251641
rect 5917 252417 5951 252433
rect 5917 251625 5951 251641
rect 6031 252417 6065 252433
rect 6031 251625 6065 251641
rect 6127 252417 6161 252433
rect 6127 251625 6161 251641
rect 6241 252417 6275 252433
rect 6241 251625 6275 251641
rect 6337 252417 6371 252433
rect 6337 251625 6371 251641
rect 6451 252417 6485 252433
rect 6451 251625 6485 251641
rect 6547 252417 6581 252433
rect 6547 251625 6581 251641
rect 6661 252417 6695 252433
rect 6661 251625 6695 251641
rect 6757 252417 6791 252433
rect 6757 251625 6791 251641
rect 6871 252417 6905 252433
rect 6871 251625 6905 251641
rect 6967 252417 7001 252433
rect 6967 251625 7001 251641
rect 7081 252417 7115 252433
rect 7081 251625 7115 251641
rect 7177 252417 7211 252433
rect 7177 251625 7211 251641
rect 7291 252417 7325 252433
rect 7291 251625 7325 251641
rect 7387 252417 7421 252433
rect 7387 251625 7421 251641
rect 7501 252417 7535 252433
rect 7501 251625 7535 251641
rect 7597 252417 7631 252433
rect 7597 251625 7631 251641
rect 7711 252417 7745 252433
rect 7711 251625 7745 251641
rect 7807 252417 7841 252433
rect 7807 251625 7841 251641
rect 7921 252417 7955 252433
rect 7921 251625 7955 251641
rect 8017 252417 8051 252433
rect 8017 251625 8051 251641
rect 8131 252417 8165 252433
rect 8131 251625 8165 251641
rect 8227 252417 8261 252433
rect 8227 251625 8261 251641
rect 8341 252417 8375 252433
rect 8341 251625 8375 251641
rect 8437 252417 8471 252433
rect 8437 251625 8471 251641
rect 8551 252417 8585 252433
rect 8551 251625 8585 251641
rect 8647 252417 8681 252433
rect 8647 251625 8681 251641
rect 8761 252417 8795 252433
rect 8761 251625 8795 251641
rect 8857 252417 8891 252433
rect 8857 251625 8891 251641
rect 8971 252417 9005 252433
rect 8971 251625 9005 251641
rect 9067 252417 9101 252433
rect 9067 251625 9101 251641
rect 9181 252417 9215 252433
rect 9181 251625 9215 251641
rect 9277 252417 9311 252433
rect 9277 251625 9311 251641
rect 9391 252417 9425 252433
rect 9391 251625 9425 251641
rect 9487 252417 9521 252433
rect 9487 251625 9521 251641
rect 9601 252417 9635 252433
rect 9601 251625 9635 251641
rect 9697 252417 9731 252433
rect 9697 251625 9731 251641
rect 9811 252417 9845 252433
rect 9811 251625 9845 251641
rect 9907 252417 9941 252433
rect 9907 251625 9941 251641
rect 10021 252417 10055 252433
rect 10021 251625 10055 251641
rect 10117 252417 10151 252433
rect 10117 251625 10151 251641
rect 10231 252417 10265 252433
rect 10231 251625 10265 251641
rect 10327 252417 10361 252433
rect 10327 251625 10361 251641
rect 10441 252417 10475 252433
rect 10441 251625 10475 251641
rect 10537 252417 10571 252433
rect 10537 251625 10571 251641
rect 10651 252417 10685 252433
rect 10651 251625 10685 251641
rect 10747 252417 10781 252433
rect 10747 251625 10781 251641
rect 10861 252417 10895 252433
rect 10861 251625 10895 251641
rect 10957 252417 10991 252433
rect 10957 251625 10991 251641
rect 11071 252417 11105 252433
rect 11071 251625 11105 251641
rect 11167 252417 11201 252433
rect 11167 251625 11201 251641
rect 11281 252417 11315 252433
rect 11281 251625 11315 251641
rect 11377 252417 11411 252433
rect 11377 251625 11411 251641
rect 11491 252417 11525 252433
rect 11491 251625 11525 251641
rect 11587 252417 11621 252433
rect 11587 251625 11621 251641
rect 11701 252417 11735 252433
rect 11701 251625 11735 251641
rect 11797 252417 11831 252433
rect 11797 251625 11831 251641
rect 11911 252417 11945 252433
rect 11911 251625 11945 251641
rect 12007 252417 12041 252433
rect 12007 251625 12041 251641
rect 12121 252417 12155 252433
rect 12121 251625 12155 251641
rect 12217 252417 12251 252433
rect 12217 251625 12251 251641
rect 12331 252417 12365 252433
rect 12331 251625 12365 251641
rect 12427 252417 12461 252433
rect 12427 251625 12461 251641
rect 12541 252417 12575 252433
rect 12541 251625 12575 251641
rect 12637 252417 12671 252433
rect 12637 251625 12671 251641
rect 12751 252417 12785 252433
rect 12751 251625 12785 251641
rect 12847 252417 12881 252433
rect 12847 251625 12881 251641
rect 12961 252417 12995 252433
rect 12961 251625 12995 251641
rect 13057 252417 13091 252433
rect 13057 251625 13091 251641
rect 13171 252417 13205 252433
rect 13171 251625 13205 251641
rect 13267 252417 13301 252433
rect 13267 251625 13301 251641
rect 13381 252417 13415 252433
rect 13381 251625 13415 251641
rect 13477 252417 13511 252433
rect 13477 251625 13511 251641
rect 13591 252417 13625 252433
rect 13591 251625 13625 251641
rect 13687 252417 13721 252433
rect 13687 251625 13721 251641
rect 13801 252417 13835 252433
rect 13801 251625 13835 251641
rect 13897 252417 13931 252433
rect 13897 251625 13931 251641
rect 14011 252417 14045 252433
rect 14011 251625 14045 251641
rect 14107 252417 14141 252433
rect 14107 251625 14141 251641
rect 14221 252417 14255 252433
rect 14221 251625 14255 251641
rect 14317 252417 14351 252433
rect 14317 251625 14351 251641
rect 14431 252417 14465 252433
rect 14431 251625 14465 251641
rect 14527 252417 14561 252433
rect 14527 251625 14561 251641
rect 14641 252417 14675 252433
rect 14641 251625 14675 251641
rect 14737 252417 14771 252433
rect 14737 251625 14771 251641
rect 14851 252417 14885 252433
rect 14851 251625 14885 251641
rect 14947 252417 14981 252433
rect 14947 251625 14981 251641
rect 15061 252417 15095 252433
rect 15061 251625 15095 251641
rect 15157 252417 15191 252433
rect 15157 251625 15191 251641
rect 15271 252417 15305 252433
rect 15271 251625 15305 251641
rect 15367 252417 15401 252433
rect 15367 251625 15401 251641
rect 15481 252417 15515 252433
rect 15481 251625 15515 251641
rect 15577 252417 15611 252433
rect 15577 251625 15611 251641
rect 15691 252417 15725 252433
rect 15691 251625 15725 251641
rect 15787 252417 15821 252433
rect 15787 251625 15821 251641
rect 15901 252417 15935 252433
rect 15901 251625 15935 251641
rect 15997 252417 16031 252433
rect 15997 251625 16031 251641
rect 16111 252417 16145 252433
rect 16111 251625 16145 251641
rect 16207 252417 16241 252433
rect 16207 251625 16241 251641
rect 16321 252417 16355 252433
rect 16321 251625 16355 251641
rect 16417 252417 16451 252433
rect 16417 251625 16451 251641
rect 16531 252417 16565 252433
rect 16531 251625 16565 251641
rect 16627 252417 16661 252433
rect 16627 251625 16661 251641
rect 16741 252417 16775 252433
rect 16741 251625 16775 251641
rect 16837 252417 16871 252433
rect 16837 251625 16871 251641
rect 16951 252417 16985 252433
rect 16951 251625 16985 251641
rect 17047 252417 17081 252433
rect 17047 251625 17081 251641
rect 17161 252417 17195 252433
rect 17161 251625 17195 251641
rect 17257 252417 17291 252433
rect 17257 251625 17291 251641
rect 17371 252417 17405 252433
rect 17371 251625 17405 251641
rect 17467 252417 17501 252433
rect 17467 251625 17501 251641
rect 17581 252417 17615 252433
rect 17581 251625 17615 251641
rect 17677 252417 17711 252433
rect 17677 251625 17711 251641
rect 17791 252417 17825 252433
rect 17791 251625 17825 251641
rect 17887 252417 17921 252433
rect 17887 251625 17921 251641
rect 18001 252417 18035 252433
rect 18001 251625 18035 251641
rect 18097 252417 18131 252433
rect 18097 251625 18131 251641
rect 18211 252417 18245 252433
rect 18211 251625 18245 251641
rect 18307 252417 18341 252433
rect 18307 251625 18341 251641
rect 18421 252417 18455 252433
rect 18421 251625 18455 251641
rect 18517 252417 18551 252433
rect 18517 251625 18551 251641
rect 18631 252417 18665 252433
rect 18631 251625 18665 251641
rect 18727 252417 18761 252433
rect 18727 251625 18761 251641
rect 18841 252417 18875 252433
rect 18841 251625 18875 251641
rect 18937 252417 18971 252433
rect 18937 251625 18971 251641
rect 19051 252417 19085 252433
rect 19051 251625 19085 251641
rect 19147 252417 19181 252433
rect 19147 251625 19181 251641
rect 19261 252417 19295 252433
rect 19261 251625 19295 251641
rect 19357 252417 19391 252433
rect 19357 251625 19391 251641
rect 19471 252417 19505 252433
rect 19471 251625 19505 251641
rect 19567 252417 19601 252433
rect 19567 251625 19601 251641
rect 19681 252417 19715 252433
rect 19681 251625 19715 251641
rect 19777 252417 19811 252433
rect 19777 251625 19811 251641
rect 19891 252417 19925 252433
rect 19891 251625 19925 251641
rect 19987 252417 20021 252433
rect 19987 251625 20021 251641
rect 20101 252417 20135 252433
rect 20101 251625 20135 251641
rect 20197 252417 20231 252433
rect 20197 251625 20231 251641
rect 20311 252417 20345 252433
rect 20311 251625 20345 251641
rect 20407 252417 20441 252433
rect 20407 251625 20441 251641
rect 20521 252417 20555 252433
rect 20521 251625 20555 251641
rect 20617 252417 20651 252433
rect 20617 251625 20651 251641
rect 20731 252417 20765 252433
rect 20731 251625 20765 251641
rect 20827 252417 20861 252433
rect 20827 251625 20861 251641
rect 20941 252417 20975 252433
rect 20941 251625 20975 251641
rect 21037 252417 21071 252433
rect 21037 251625 21071 251641
rect 21151 252417 21185 252433
rect 21151 251625 21185 251641
rect 21247 252417 21281 252433
rect 21247 251625 21281 251641
rect 21361 252417 21395 252433
rect 21361 251625 21395 251641
rect 21457 252417 21491 252433
rect 21457 251625 21491 251641
rect 21571 252417 21605 252433
rect 21571 251625 21605 251641
rect 21667 252417 21701 252433
rect 21667 251625 21701 251641
rect 21781 252417 21815 252433
rect 21781 251625 21815 251641
rect 21877 252417 21911 252433
rect 21877 251625 21911 251641
rect 21991 252417 22025 252433
rect 21991 251625 22025 251641
rect 22087 252417 22121 252433
rect 22087 251625 22121 251641
rect 22201 252417 22235 252433
rect 22201 251625 22235 251641
rect 22297 252417 22331 252433
rect 22297 251625 22331 251641
rect 22411 252417 22445 252433
rect 22411 251625 22445 251641
rect 22507 252417 22541 252433
rect 22507 251625 22541 251641
rect 22621 252417 22655 252433
rect 22621 251625 22655 251641
rect 22717 252417 22751 252433
rect 22717 251625 22751 251641
rect 22831 252417 22865 252433
rect 22831 251625 22865 251641
rect 22927 252417 22961 252433
rect 22927 251625 22961 251641
rect 23041 252417 23075 252433
rect 23041 251625 23075 251641
rect 23137 252417 23171 252433
rect 23137 251625 23171 251641
rect 23251 252417 23285 252433
rect 23251 251625 23285 251641
rect 23347 252417 23381 252433
rect 23347 251625 23381 251641
rect 23461 252417 23495 252433
rect 23461 251625 23495 251641
rect 23557 252417 23591 252433
rect 23557 251625 23591 251641
rect 23671 252417 23705 252433
rect 23671 251625 23705 251641
rect 23767 252417 23801 252433
rect 23767 251625 23801 251641
rect 23881 252417 23915 252433
rect 23881 251625 23915 251641
rect 23977 252417 24011 252433
rect 23977 251625 24011 251641
rect 24091 252417 24125 252433
rect 24091 251625 24125 251641
rect 24187 252417 24221 252433
rect 24187 251625 24221 251641
rect 24301 252417 24335 252433
rect 24301 251625 24335 251641
rect 24397 252417 24431 252433
rect 24397 251625 24431 251641
rect 24511 252417 24545 252433
rect 24511 251625 24545 251641
rect 24607 252417 24641 252433
rect 24607 251625 24641 251641
rect 24721 252417 24755 252433
rect 24721 251625 24755 251641
rect 24817 252417 24851 252433
rect 24817 251625 24851 251641
rect 24931 252417 24965 252433
rect 24931 251625 24965 251641
rect 25027 252417 25061 252433
rect 25027 251625 25061 251641
rect 25141 252417 25175 252433
rect 25141 251625 25175 251641
rect 25237 252417 25271 252433
rect 25237 251625 25271 251641
rect 25351 252417 25385 252433
rect 25351 251625 25385 251641
rect 25447 252417 25481 252433
rect 25447 251625 25481 251641
rect 25561 252417 25595 252433
rect 25561 251625 25595 251641
rect 25657 252417 25691 252433
rect 25657 251625 25691 251641
rect 25771 252417 25805 252433
rect 25771 251625 25805 251641
rect 25867 252417 25901 252433
rect 25867 251625 25901 251641
rect 25981 252417 26015 252433
rect 25981 251625 26015 251641
rect 26077 252417 26111 252433
rect 26077 251625 26111 251641
rect 26191 252417 26225 252433
rect 26191 251625 26225 251641
rect 26287 252417 26321 252433
rect 26287 251625 26321 251641
rect 26401 252417 26435 252433
rect 26401 251625 26435 251641
rect 26497 252417 26531 252433
rect 26497 251625 26531 251641
rect 26611 252417 26645 252433
rect 26611 251625 26645 251641
rect 26707 252417 26741 252433
rect 26707 251625 26741 251641
rect 26821 252417 26855 252433
rect 26821 251625 26855 251641
rect 26917 252417 26951 252433
rect 26917 251625 26951 251641
rect 27031 252417 27065 252433
rect 27031 251625 27065 251641
rect 27127 252417 27161 252433
rect 27127 251625 27161 251641
rect 27241 252417 27275 252433
rect 27241 251625 27275 251641
rect 27337 252417 27371 252433
rect 27337 251625 27371 251641
rect -3807 251548 -3791 251582
rect -3807 251440 -3791 251474
rect -3757 251548 -3741 251582
rect -3387 251548 -3371 251582
rect -3757 251440 -3741 251474
rect -3387 251440 -3371 251474
rect -3337 251548 -3321 251582
rect -2967 251548 -2951 251582
rect -3337 251440 -3321 251474
rect -2967 251440 -2951 251474
rect -2917 251548 -2901 251582
rect -2547 251548 -2531 251582
rect -2917 251440 -2901 251474
rect -2547 251440 -2531 251474
rect -2497 251548 -2481 251582
rect -2127 251548 -2111 251582
rect -2497 251440 -2481 251474
rect -2127 251440 -2111 251474
rect -2077 251548 -2061 251582
rect -1707 251548 -1691 251582
rect -2077 251440 -2061 251474
rect -1707 251440 -1691 251474
rect -1657 251548 -1641 251582
rect -1287 251548 -1271 251582
rect -1657 251440 -1641 251474
rect -1287 251440 -1271 251474
rect -1237 251548 -1221 251582
rect -867 251548 -851 251582
rect -1237 251440 -1221 251474
rect -867 251440 -851 251474
rect -817 251548 -801 251582
rect -447 251548 -431 251582
rect -817 251440 -801 251474
rect -447 251440 -431 251474
rect -397 251548 -381 251582
rect -27 251548 -11 251582
rect -397 251440 -381 251474
rect -27 251440 -11 251474
rect 23 251548 39 251582
rect 393 251548 409 251582
rect 23 251440 39 251474
rect 393 251440 409 251474
rect 443 251548 459 251582
rect 813 251548 829 251582
rect 443 251440 459 251474
rect 813 251440 829 251474
rect 863 251548 879 251582
rect 1233 251548 1249 251582
rect 863 251440 879 251474
rect 1233 251440 1249 251474
rect 1283 251548 1299 251582
rect 1653 251548 1669 251582
rect 1283 251440 1299 251474
rect 1653 251440 1669 251474
rect 1703 251548 1719 251582
rect 2073 251548 2089 251582
rect 1703 251440 1719 251474
rect 2073 251440 2089 251474
rect 2123 251548 2139 251582
rect 2493 251548 2509 251582
rect 2123 251440 2139 251474
rect 2493 251440 2509 251474
rect 2543 251548 2559 251582
rect 2913 251548 2929 251582
rect 2543 251440 2559 251474
rect 2913 251440 2929 251474
rect 2963 251548 2979 251582
rect 3333 251548 3349 251582
rect 2963 251440 2979 251474
rect 3333 251440 3349 251474
rect 3383 251548 3399 251582
rect 3753 251548 3769 251582
rect 3383 251440 3399 251474
rect 3753 251440 3769 251474
rect 3803 251548 3819 251582
rect 4173 251548 4189 251582
rect 3803 251440 3819 251474
rect 4173 251440 4189 251474
rect 4223 251548 4239 251582
rect 4593 251548 4609 251582
rect 4223 251440 4239 251474
rect 4593 251440 4609 251474
rect 4643 251548 4659 251582
rect 5013 251548 5029 251582
rect 4643 251440 4659 251474
rect 5013 251440 5029 251474
rect 5063 251548 5079 251582
rect 5433 251548 5449 251582
rect 5063 251440 5079 251474
rect 5433 251440 5449 251474
rect 5483 251548 5499 251582
rect 5853 251548 5869 251582
rect 5483 251440 5499 251474
rect 5853 251440 5869 251474
rect 5903 251548 5919 251582
rect 6273 251548 6289 251582
rect 5903 251440 5919 251474
rect 6273 251440 6289 251474
rect 6323 251548 6339 251582
rect 6693 251548 6709 251582
rect 6323 251440 6339 251474
rect 6693 251440 6709 251474
rect 6743 251548 6759 251582
rect 7113 251548 7129 251582
rect 6743 251440 6759 251474
rect 7113 251440 7129 251474
rect 7163 251548 7179 251582
rect 7533 251548 7549 251582
rect 7163 251440 7179 251474
rect 7533 251440 7549 251474
rect 7583 251548 7599 251582
rect 7953 251548 7969 251582
rect 7583 251440 7599 251474
rect 7953 251440 7969 251474
rect 8003 251548 8019 251582
rect 8373 251548 8389 251582
rect 8003 251440 8019 251474
rect 8373 251440 8389 251474
rect 8423 251548 8439 251582
rect 8793 251548 8809 251582
rect 8423 251440 8439 251474
rect 8793 251440 8809 251474
rect 8843 251548 8859 251582
rect 9213 251548 9229 251582
rect 8843 251440 8859 251474
rect 9213 251440 9229 251474
rect 9263 251548 9279 251582
rect 9633 251548 9649 251582
rect 9263 251440 9279 251474
rect 9633 251440 9649 251474
rect 9683 251548 9699 251582
rect 10053 251548 10069 251582
rect 9683 251440 9699 251474
rect 10053 251440 10069 251474
rect 10103 251548 10119 251582
rect 10473 251548 10489 251582
rect 10103 251440 10119 251474
rect 10473 251440 10489 251474
rect 10523 251548 10539 251582
rect 10893 251548 10909 251582
rect 10523 251440 10539 251474
rect 10893 251440 10909 251474
rect 10943 251548 10959 251582
rect 11313 251548 11329 251582
rect 10943 251440 10959 251474
rect 11313 251440 11329 251474
rect 11363 251548 11379 251582
rect 11733 251548 11749 251582
rect 11363 251440 11379 251474
rect 11733 251440 11749 251474
rect 11783 251548 11799 251582
rect 12153 251548 12169 251582
rect 11783 251440 11799 251474
rect 12153 251440 12169 251474
rect 12203 251548 12219 251582
rect 12573 251548 12589 251582
rect 12203 251440 12219 251474
rect 12573 251440 12589 251474
rect 12623 251548 12639 251582
rect 12993 251548 13009 251582
rect 12623 251440 12639 251474
rect 12993 251440 13009 251474
rect 13043 251548 13059 251582
rect 13413 251548 13429 251582
rect 13043 251440 13059 251474
rect 13413 251440 13429 251474
rect 13463 251548 13479 251582
rect 13833 251548 13849 251582
rect 13463 251440 13479 251474
rect 13833 251440 13849 251474
rect 13883 251548 13899 251582
rect 14253 251548 14269 251582
rect 13883 251440 13899 251474
rect 14253 251440 14269 251474
rect 14303 251548 14319 251582
rect 14673 251548 14689 251582
rect 14303 251440 14319 251474
rect 14673 251440 14689 251474
rect 14723 251548 14739 251582
rect 15093 251548 15109 251582
rect 14723 251440 14739 251474
rect 15093 251440 15109 251474
rect 15143 251548 15159 251582
rect 15513 251548 15529 251582
rect 15143 251440 15159 251474
rect 15513 251440 15529 251474
rect 15563 251548 15579 251582
rect 15933 251548 15949 251582
rect 15563 251440 15579 251474
rect 15933 251440 15949 251474
rect 15983 251548 15999 251582
rect 16353 251548 16369 251582
rect 15983 251440 15999 251474
rect 16353 251440 16369 251474
rect 16403 251548 16419 251582
rect 16773 251548 16789 251582
rect 16403 251440 16419 251474
rect 16773 251440 16789 251474
rect 16823 251548 16839 251582
rect 17193 251548 17209 251582
rect 16823 251440 16839 251474
rect 17193 251440 17209 251474
rect 17243 251548 17259 251582
rect 17613 251548 17629 251582
rect 17243 251440 17259 251474
rect 17613 251440 17629 251474
rect 17663 251548 17679 251582
rect 18033 251548 18049 251582
rect 17663 251440 17679 251474
rect 18033 251440 18049 251474
rect 18083 251548 18099 251582
rect 18453 251548 18469 251582
rect 18083 251440 18099 251474
rect 18453 251440 18469 251474
rect 18503 251548 18519 251582
rect 18873 251548 18889 251582
rect 18503 251440 18519 251474
rect 18873 251440 18889 251474
rect 18923 251548 18939 251582
rect 19293 251548 19309 251582
rect 18923 251440 18939 251474
rect 19293 251440 19309 251474
rect 19343 251548 19359 251582
rect 19713 251548 19729 251582
rect 19343 251440 19359 251474
rect 19713 251440 19729 251474
rect 19763 251548 19779 251582
rect 20133 251548 20149 251582
rect 19763 251440 19779 251474
rect 20133 251440 20149 251474
rect 20183 251548 20199 251582
rect 20553 251548 20569 251582
rect 20183 251440 20199 251474
rect 20553 251440 20569 251474
rect 20603 251548 20619 251582
rect 20973 251548 20989 251582
rect 20603 251440 20619 251474
rect 20973 251440 20989 251474
rect 21023 251548 21039 251582
rect 21393 251548 21409 251582
rect 21023 251440 21039 251474
rect 21393 251440 21409 251474
rect 21443 251548 21459 251582
rect 21813 251548 21829 251582
rect 21443 251440 21459 251474
rect 21813 251440 21829 251474
rect 21863 251548 21879 251582
rect 22233 251548 22249 251582
rect 21863 251440 21879 251474
rect 22233 251440 22249 251474
rect 22283 251548 22299 251582
rect 22653 251548 22669 251582
rect 22283 251440 22299 251474
rect 22653 251440 22669 251474
rect 22703 251548 22719 251582
rect 23073 251548 23089 251582
rect 22703 251440 22719 251474
rect 23073 251440 23089 251474
rect 23123 251548 23139 251582
rect 23493 251548 23509 251582
rect 23123 251440 23139 251474
rect 23493 251440 23509 251474
rect 23543 251548 23559 251582
rect 23913 251548 23929 251582
rect 23543 251440 23559 251474
rect 23913 251440 23929 251474
rect 23963 251548 23979 251582
rect 24333 251548 24349 251582
rect 23963 251440 23979 251474
rect 24333 251440 24349 251474
rect 24383 251548 24399 251582
rect 24753 251548 24769 251582
rect 24383 251440 24399 251474
rect 24753 251440 24769 251474
rect 24803 251548 24819 251582
rect 25173 251548 25189 251582
rect 24803 251440 24819 251474
rect 25173 251440 25189 251474
rect 25223 251548 25239 251582
rect 25593 251548 25609 251582
rect 25223 251440 25239 251474
rect 25593 251440 25609 251474
rect 25643 251548 25659 251582
rect 26013 251548 26029 251582
rect 25643 251440 25659 251474
rect 26013 251440 26029 251474
rect 26063 251548 26079 251582
rect 26433 251548 26449 251582
rect 26063 251440 26079 251474
rect 26433 251440 26449 251474
rect 26483 251548 26499 251582
rect 26853 251548 26869 251582
rect 26483 251440 26499 251474
rect 26853 251440 26869 251474
rect 26903 251548 26919 251582
rect 27273 251548 27289 251582
rect 26903 251440 26919 251474
rect 27273 251440 27289 251474
rect 27323 251548 27339 251582
rect 27323 251440 27339 251474
rect -4049 251381 -4015 251397
rect -4049 250589 -4015 250605
rect -3953 251381 -3919 251397
rect -3953 250589 -3919 250605
rect -3839 251381 -3805 251397
rect -3839 250589 -3805 250605
rect -3743 251381 -3709 251397
rect -3743 250589 -3709 250605
rect -3629 251381 -3595 251397
rect -3629 250589 -3595 250605
rect -3533 251381 -3499 251397
rect -3533 250589 -3499 250605
rect -3419 251381 -3385 251397
rect -3419 250589 -3385 250605
rect -3323 251381 -3289 251397
rect -3323 250589 -3289 250605
rect -3209 251381 -3175 251397
rect -3209 250589 -3175 250605
rect -3113 251381 -3079 251397
rect -3113 250589 -3079 250605
rect -2999 251381 -2965 251397
rect -2999 250589 -2965 250605
rect -2903 251381 -2869 251397
rect -2903 250589 -2869 250605
rect -2789 251381 -2755 251397
rect -2789 250589 -2755 250605
rect -2693 251381 -2659 251397
rect -2693 250589 -2659 250605
rect -2579 251381 -2545 251397
rect -2579 250589 -2545 250605
rect -2483 251381 -2449 251397
rect -2483 250589 -2449 250605
rect -2369 251381 -2335 251397
rect -2369 250589 -2335 250605
rect -2273 251381 -2239 251397
rect -2273 250589 -2239 250605
rect -2159 251381 -2125 251397
rect -2159 250589 -2125 250605
rect -2063 251381 -2029 251397
rect -2063 250589 -2029 250605
rect -1949 251381 -1915 251397
rect -1949 250589 -1915 250605
rect -1853 251381 -1819 251397
rect -1853 250589 -1819 250605
rect -1739 251381 -1705 251397
rect -1739 250589 -1705 250605
rect -1643 251381 -1609 251397
rect -1643 250589 -1609 250605
rect -1529 251381 -1495 251397
rect -1529 250589 -1495 250605
rect -1433 251381 -1399 251397
rect -1433 250589 -1399 250605
rect -1319 251381 -1285 251397
rect -1319 250589 -1285 250605
rect -1223 251381 -1189 251397
rect -1223 250589 -1189 250605
rect -1109 251381 -1075 251397
rect -1109 250589 -1075 250605
rect -1013 251381 -979 251397
rect -1013 250589 -979 250605
rect -899 251381 -865 251397
rect -899 250589 -865 250605
rect -803 251381 -769 251397
rect -803 250589 -769 250605
rect -689 251381 -655 251397
rect -689 250589 -655 250605
rect -593 251381 -559 251397
rect -593 250589 -559 250605
rect -479 251381 -445 251397
rect -479 250589 -445 250605
rect -383 251381 -349 251397
rect -383 250589 -349 250605
rect -269 251381 -235 251397
rect -269 250589 -235 250605
rect -173 251381 -139 251397
rect -173 250589 -139 250605
rect -59 251381 -25 251397
rect -59 250589 -25 250605
rect 37 251381 71 251397
rect 37 250589 71 250605
rect 151 251381 185 251397
rect 151 250589 185 250605
rect 247 251381 281 251397
rect 247 250589 281 250605
rect 361 251381 395 251397
rect 361 250589 395 250605
rect 457 251381 491 251397
rect 457 250589 491 250605
rect 571 251381 605 251397
rect 571 250589 605 250605
rect 667 251381 701 251397
rect 667 250589 701 250605
rect 781 251381 815 251397
rect 781 250589 815 250605
rect 877 251381 911 251397
rect 877 250589 911 250605
rect 991 251381 1025 251397
rect 991 250589 1025 250605
rect 1087 251381 1121 251397
rect 1087 250589 1121 250605
rect 1201 251381 1235 251397
rect 1201 250589 1235 250605
rect 1297 251381 1331 251397
rect 1297 250589 1331 250605
rect 1411 251381 1445 251397
rect 1411 250589 1445 250605
rect 1507 251381 1541 251397
rect 1507 250589 1541 250605
rect 1621 251381 1655 251397
rect 1621 250589 1655 250605
rect 1717 251381 1751 251397
rect 1717 250589 1751 250605
rect 1831 251381 1865 251397
rect 1831 250589 1865 250605
rect 1927 251381 1961 251397
rect 1927 250589 1961 250605
rect 2041 251381 2075 251397
rect 2041 250589 2075 250605
rect 2137 251381 2171 251397
rect 2137 250589 2171 250605
rect 2251 251381 2285 251397
rect 2251 250589 2285 250605
rect 2347 251381 2381 251397
rect 2347 250589 2381 250605
rect 2461 251381 2495 251397
rect 2461 250589 2495 250605
rect 2557 251381 2591 251397
rect 2557 250589 2591 250605
rect 2671 251381 2705 251397
rect 2671 250589 2705 250605
rect 2767 251381 2801 251397
rect 2767 250589 2801 250605
rect 2881 251381 2915 251397
rect 2881 250589 2915 250605
rect 2977 251381 3011 251397
rect 2977 250589 3011 250605
rect 3091 251381 3125 251397
rect 3091 250589 3125 250605
rect 3187 251381 3221 251397
rect 3187 250589 3221 250605
rect 3301 251381 3335 251397
rect 3301 250589 3335 250605
rect 3397 251381 3431 251397
rect 3397 250589 3431 250605
rect 3511 251381 3545 251397
rect 3511 250589 3545 250605
rect 3607 251381 3641 251397
rect 3607 250589 3641 250605
rect 3721 251381 3755 251397
rect 3721 250589 3755 250605
rect 3817 251381 3851 251397
rect 3817 250589 3851 250605
rect 3931 251381 3965 251397
rect 3931 250589 3965 250605
rect 4027 251381 4061 251397
rect 4027 250589 4061 250605
rect 4141 251381 4175 251397
rect 4141 250589 4175 250605
rect 4237 251381 4271 251397
rect 4237 250589 4271 250605
rect 4351 251381 4385 251397
rect 4351 250589 4385 250605
rect 4447 251381 4481 251397
rect 4447 250589 4481 250605
rect 4561 251381 4595 251397
rect 4561 250589 4595 250605
rect 4657 251381 4691 251397
rect 4657 250589 4691 250605
rect 4771 251381 4805 251397
rect 4771 250589 4805 250605
rect 4867 251381 4901 251397
rect 4867 250589 4901 250605
rect 4981 251381 5015 251397
rect 4981 250589 5015 250605
rect 5077 251381 5111 251397
rect 5077 250589 5111 250605
rect 5191 251381 5225 251397
rect 5191 250589 5225 250605
rect 5287 251381 5321 251397
rect 5287 250589 5321 250605
rect 5401 251381 5435 251397
rect 5401 250589 5435 250605
rect 5497 251381 5531 251397
rect 5497 250589 5531 250605
rect 5611 251381 5645 251397
rect 5611 250589 5645 250605
rect 5707 251381 5741 251397
rect 5707 250589 5741 250605
rect 5821 251381 5855 251397
rect 5821 250589 5855 250605
rect 5917 251381 5951 251397
rect 5917 250589 5951 250605
rect 6031 251381 6065 251397
rect 6031 250589 6065 250605
rect 6127 251381 6161 251397
rect 6127 250589 6161 250605
rect 6241 251381 6275 251397
rect 6241 250589 6275 250605
rect 6337 251381 6371 251397
rect 6337 250589 6371 250605
rect 6451 251381 6485 251397
rect 6451 250589 6485 250605
rect 6547 251381 6581 251397
rect 6547 250589 6581 250605
rect 6661 251381 6695 251397
rect 6661 250589 6695 250605
rect 6757 251381 6791 251397
rect 6757 250589 6791 250605
rect 6871 251381 6905 251397
rect 6871 250589 6905 250605
rect 6967 251381 7001 251397
rect 6967 250589 7001 250605
rect 7081 251381 7115 251397
rect 7081 250589 7115 250605
rect 7177 251381 7211 251397
rect 7177 250589 7211 250605
rect 7291 251381 7325 251397
rect 7291 250589 7325 250605
rect 7387 251381 7421 251397
rect 7387 250589 7421 250605
rect 7501 251381 7535 251397
rect 7501 250589 7535 250605
rect 7597 251381 7631 251397
rect 7597 250589 7631 250605
rect 7711 251381 7745 251397
rect 7711 250589 7745 250605
rect 7807 251381 7841 251397
rect 7807 250589 7841 250605
rect 7921 251381 7955 251397
rect 7921 250589 7955 250605
rect 8017 251381 8051 251397
rect 8017 250589 8051 250605
rect 8131 251381 8165 251397
rect 8131 250589 8165 250605
rect 8227 251381 8261 251397
rect 8227 250589 8261 250605
rect 8341 251381 8375 251397
rect 8341 250589 8375 250605
rect 8437 251381 8471 251397
rect 8437 250589 8471 250605
rect 8551 251381 8585 251397
rect 8551 250589 8585 250605
rect 8647 251381 8681 251397
rect 8647 250589 8681 250605
rect 8761 251381 8795 251397
rect 8761 250589 8795 250605
rect 8857 251381 8891 251397
rect 8857 250589 8891 250605
rect 8971 251381 9005 251397
rect 8971 250589 9005 250605
rect 9067 251381 9101 251397
rect 9067 250589 9101 250605
rect 9181 251381 9215 251397
rect 9181 250589 9215 250605
rect 9277 251381 9311 251397
rect 9277 250589 9311 250605
rect 9391 251381 9425 251397
rect 9391 250589 9425 250605
rect 9487 251381 9521 251397
rect 9487 250589 9521 250605
rect 9601 251381 9635 251397
rect 9601 250589 9635 250605
rect 9697 251381 9731 251397
rect 9697 250589 9731 250605
rect 9811 251381 9845 251397
rect 9811 250589 9845 250605
rect 9907 251381 9941 251397
rect 9907 250589 9941 250605
rect 10021 251381 10055 251397
rect 10021 250589 10055 250605
rect 10117 251381 10151 251397
rect 10117 250589 10151 250605
rect 10231 251381 10265 251397
rect 10231 250589 10265 250605
rect 10327 251381 10361 251397
rect 10327 250589 10361 250605
rect 10441 251381 10475 251397
rect 10441 250589 10475 250605
rect 10537 251381 10571 251397
rect 10537 250589 10571 250605
rect 10651 251381 10685 251397
rect 10651 250589 10685 250605
rect 10747 251381 10781 251397
rect 10747 250589 10781 250605
rect 10861 251381 10895 251397
rect 10861 250589 10895 250605
rect 10957 251381 10991 251397
rect 10957 250589 10991 250605
rect 11071 251381 11105 251397
rect 11071 250589 11105 250605
rect 11167 251381 11201 251397
rect 11167 250589 11201 250605
rect 11281 251381 11315 251397
rect 11281 250589 11315 250605
rect 11377 251381 11411 251397
rect 11377 250589 11411 250605
rect 11491 251381 11525 251397
rect 11491 250589 11525 250605
rect 11587 251381 11621 251397
rect 11587 250589 11621 250605
rect 11701 251381 11735 251397
rect 11701 250589 11735 250605
rect 11797 251381 11831 251397
rect 11797 250589 11831 250605
rect 11911 251381 11945 251397
rect 11911 250589 11945 250605
rect 12007 251381 12041 251397
rect 12007 250589 12041 250605
rect 12121 251381 12155 251397
rect 12121 250589 12155 250605
rect 12217 251381 12251 251397
rect 12217 250589 12251 250605
rect 12331 251381 12365 251397
rect 12331 250589 12365 250605
rect 12427 251381 12461 251397
rect 12427 250589 12461 250605
rect 12541 251381 12575 251397
rect 12541 250589 12575 250605
rect 12637 251381 12671 251397
rect 12637 250589 12671 250605
rect 12751 251381 12785 251397
rect 12751 250589 12785 250605
rect 12847 251381 12881 251397
rect 12847 250589 12881 250605
rect 12961 251381 12995 251397
rect 12961 250589 12995 250605
rect 13057 251381 13091 251397
rect 13057 250589 13091 250605
rect 13171 251381 13205 251397
rect 13171 250589 13205 250605
rect 13267 251381 13301 251397
rect 13267 250589 13301 250605
rect 13381 251381 13415 251397
rect 13381 250589 13415 250605
rect 13477 251381 13511 251397
rect 13477 250589 13511 250605
rect 13591 251381 13625 251397
rect 13591 250589 13625 250605
rect 13687 251381 13721 251397
rect 13687 250589 13721 250605
rect 13801 251381 13835 251397
rect 13801 250589 13835 250605
rect 13897 251381 13931 251397
rect 13897 250589 13931 250605
rect 14011 251381 14045 251397
rect 14011 250589 14045 250605
rect 14107 251381 14141 251397
rect 14107 250589 14141 250605
rect 14221 251381 14255 251397
rect 14221 250589 14255 250605
rect 14317 251381 14351 251397
rect 14317 250589 14351 250605
rect 14431 251381 14465 251397
rect 14431 250589 14465 250605
rect 14527 251381 14561 251397
rect 14527 250589 14561 250605
rect 14641 251381 14675 251397
rect 14641 250589 14675 250605
rect 14737 251381 14771 251397
rect 14737 250589 14771 250605
rect 14851 251381 14885 251397
rect 14851 250589 14885 250605
rect 14947 251381 14981 251397
rect 14947 250589 14981 250605
rect 15061 251381 15095 251397
rect 15061 250589 15095 250605
rect 15157 251381 15191 251397
rect 15157 250589 15191 250605
rect 15271 251381 15305 251397
rect 15271 250589 15305 250605
rect 15367 251381 15401 251397
rect 15367 250589 15401 250605
rect 15481 251381 15515 251397
rect 15481 250589 15515 250605
rect 15577 251381 15611 251397
rect 15577 250589 15611 250605
rect 15691 251381 15725 251397
rect 15691 250589 15725 250605
rect 15787 251381 15821 251397
rect 15787 250589 15821 250605
rect 15901 251381 15935 251397
rect 15901 250589 15935 250605
rect 15997 251381 16031 251397
rect 15997 250589 16031 250605
rect 16111 251381 16145 251397
rect 16111 250589 16145 250605
rect 16207 251381 16241 251397
rect 16207 250589 16241 250605
rect 16321 251381 16355 251397
rect 16321 250589 16355 250605
rect 16417 251381 16451 251397
rect 16417 250589 16451 250605
rect 16531 251381 16565 251397
rect 16531 250589 16565 250605
rect 16627 251381 16661 251397
rect 16627 250589 16661 250605
rect 16741 251381 16775 251397
rect 16741 250589 16775 250605
rect 16837 251381 16871 251397
rect 16837 250589 16871 250605
rect 16951 251381 16985 251397
rect 16951 250589 16985 250605
rect 17047 251381 17081 251397
rect 17047 250589 17081 250605
rect 17161 251381 17195 251397
rect 17161 250589 17195 250605
rect 17257 251381 17291 251397
rect 17257 250589 17291 250605
rect 17371 251381 17405 251397
rect 17371 250589 17405 250605
rect 17467 251381 17501 251397
rect 17467 250589 17501 250605
rect 17581 251381 17615 251397
rect 17581 250589 17615 250605
rect 17677 251381 17711 251397
rect 17677 250589 17711 250605
rect 17791 251381 17825 251397
rect 17791 250589 17825 250605
rect 17887 251381 17921 251397
rect 17887 250589 17921 250605
rect 18001 251381 18035 251397
rect 18001 250589 18035 250605
rect 18097 251381 18131 251397
rect 18097 250589 18131 250605
rect 18211 251381 18245 251397
rect 18211 250589 18245 250605
rect 18307 251381 18341 251397
rect 18307 250589 18341 250605
rect 18421 251381 18455 251397
rect 18421 250589 18455 250605
rect 18517 251381 18551 251397
rect 18517 250589 18551 250605
rect 18631 251381 18665 251397
rect 18631 250589 18665 250605
rect 18727 251381 18761 251397
rect 18727 250589 18761 250605
rect 18841 251381 18875 251397
rect 18841 250589 18875 250605
rect 18937 251381 18971 251397
rect 18937 250589 18971 250605
rect 19051 251381 19085 251397
rect 19051 250589 19085 250605
rect 19147 251381 19181 251397
rect 19147 250589 19181 250605
rect 19261 251381 19295 251397
rect 19261 250589 19295 250605
rect 19357 251381 19391 251397
rect 19357 250589 19391 250605
rect 19471 251381 19505 251397
rect 19471 250589 19505 250605
rect 19567 251381 19601 251397
rect 19567 250589 19601 250605
rect 19681 251381 19715 251397
rect 19681 250589 19715 250605
rect 19777 251381 19811 251397
rect 19777 250589 19811 250605
rect 19891 251381 19925 251397
rect 19891 250589 19925 250605
rect 19987 251381 20021 251397
rect 19987 250589 20021 250605
rect 20101 251381 20135 251397
rect 20101 250589 20135 250605
rect 20197 251381 20231 251397
rect 20197 250589 20231 250605
rect 20311 251381 20345 251397
rect 20311 250589 20345 250605
rect 20407 251381 20441 251397
rect 20407 250589 20441 250605
rect 20521 251381 20555 251397
rect 20521 250589 20555 250605
rect 20617 251381 20651 251397
rect 20617 250589 20651 250605
rect 20731 251381 20765 251397
rect 20731 250589 20765 250605
rect 20827 251381 20861 251397
rect 20827 250589 20861 250605
rect 20941 251381 20975 251397
rect 20941 250589 20975 250605
rect 21037 251381 21071 251397
rect 21037 250589 21071 250605
rect 21151 251381 21185 251397
rect 21151 250589 21185 250605
rect 21247 251381 21281 251397
rect 21247 250589 21281 250605
rect 21361 251381 21395 251397
rect 21361 250589 21395 250605
rect 21457 251381 21491 251397
rect 21457 250589 21491 250605
rect 21571 251381 21605 251397
rect 21571 250589 21605 250605
rect 21667 251381 21701 251397
rect 21667 250589 21701 250605
rect 21781 251381 21815 251397
rect 21781 250589 21815 250605
rect 21877 251381 21911 251397
rect 21877 250589 21911 250605
rect 21991 251381 22025 251397
rect 21991 250589 22025 250605
rect 22087 251381 22121 251397
rect 22087 250589 22121 250605
rect 22201 251381 22235 251397
rect 22201 250589 22235 250605
rect 22297 251381 22331 251397
rect 22297 250589 22331 250605
rect 22411 251381 22445 251397
rect 22411 250589 22445 250605
rect 22507 251381 22541 251397
rect 22507 250589 22541 250605
rect 22621 251381 22655 251397
rect 22621 250589 22655 250605
rect 22717 251381 22751 251397
rect 22717 250589 22751 250605
rect 22831 251381 22865 251397
rect 22831 250589 22865 250605
rect 22927 251381 22961 251397
rect 22927 250589 22961 250605
rect 23041 251381 23075 251397
rect 23041 250589 23075 250605
rect 23137 251381 23171 251397
rect 23137 250589 23171 250605
rect 23251 251381 23285 251397
rect 23251 250589 23285 250605
rect 23347 251381 23381 251397
rect 23347 250589 23381 250605
rect 23461 251381 23495 251397
rect 23461 250589 23495 250605
rect 23557 251381 23591 251397
rect 23557 250589 23591 250605
rect 23671 251381 23705 251397
rect 23671 250589 23705 250605
rect 23767 251381 23801 251397
rect 23767 250589 23801 250605
rect 23881 251381 23915 251397
rect 23881 250589 23915 250605
rect 23977 251381 24011 251397
rect 23977 250589 24011 250605
rect 24091 251381 24125 251397
rect 24091 250589 24125 250605
rect 24187 251381 24221 251397
rect 24187 250589 24221 250605
rect 24301 251381 24335 251397
rect 24301 250589 24335 250605
rect 24397 251381 24431 251397
rect 24397 250589 24431 250605
rect 24511 251381 24545 251397
rect 24511 250589 24545 250605
rect 24607 251381 24641 251397
rect 24607 250589 24641 250605
rect 24721 251381 24755 251397
rect 24721 250589 24755 250605
rect 24817 251381 24851 251397
rect 24817 250589 24851 250605
rect 24931 251381 24965 251397
rect 24931 250589 24965 250605
rect 25027 251381 25061 251397
rect 25027 250589 25061 250605
rect 25141 251381 25175 251397
rect 25141 250589 25175 250605
rect 25237 251381 25271 251397
rect 25237 250589 25271 250605
rect 25351 251381 25385 251397
rect 25351 250589 25385 250605
rect 25447 251381 25481 251397
rect 25447 250589 25481 250605
rect 25561 251381 25595 251397
rect 25561 250589 25595 250605
rect 25657 251381 25691 251397
rect 25657 250589 25691 250605
rect 25771 251381 25805 251397
rect 25771 250589 25805 250605
rect 25867 251381 25901 251397
rect 25867 250589 25901 250605
rect 25981 251381 26015 251397
rect 25981 250589 26015 250605
rect 26077 251381 26111 251397
rect 26077 250589 26111 250605
rect 26191 251381 26225 251397
rect 26191 250589 26225 250605
rect 26287 251381 26321 251397
rect 26287 250589 26321 250605
rect 26401 251381 26435 251397
rect 26401 250589 26435 250605
rect 26497 251381 26531 251397
rect 26497 250589 26531 250605
rect 26611 251381 26645 251397
rect 26611 250589 26645 250605
rect 26707 251381 26741 251397
rect 26707 250589 26741 250605
rect 26821 251381 26855 251397
rect 26821 250589 26855 250605
rect 26917 251381 26951 251397
rect 26917 250589 26951 250605
rect 27031 251381 27065 251397
rect 27031 250589 27065 250605
rect 27127 251381 27161 251397
rect 27127 250589 27161 250605
rect 27241 251381 27275 251397
rect 27241 250589 27275 250605
rect 27337 251381 27371 251397
rect 27337 250589 27371 250605
rect -4017 250512 -4001 250546
rect -4017 250404 -4001 250438
rect -3967 250512 -3951 250546
rect -3597 250512 -3581 250546
rect -3967 250404 -3951 250438
rect -3597 250404 -3581 250438
rect -3547 250512 -3531 250546
rect -3177 250512 -3161 250546
rect -3547 250404 -3531 250438
rect -3177 250404 -3161 250438
rect -3127 250512 -3111 250546
rect -2757 250512 -2741 250546
rect -3127 250404 -3111 250438
rect -2757 250404 -2741 250438
rect -2707 250512 -2691 250546
rect -2337 250512 -2321 250546
rect -2707 250404 -2691 250438
rect -2337 250404 -2321 250438
rect -2287 250512 -2271 250546
rect -1917 250512 -1901 250546
rect -2287 250404 -2271 250438
rect -1917 250404 -1901 250438
rect -1867 250512 -1851 250546
rect -1497 250512 -1481 250546
rect -1867 250404 -1851 250438
rect -1497 250404 -1481 250438
rect -1447 250512 -1431 250546
rect -1077 250512 -1061 250546
rect -1447 250404 -1431 250438
rect -1077 250404 -1061 250438
rect -1027 250512 -1011 250546
rect -657 250512 -641 250546
rect -1027 250404 -1011 250438
rect -657 250404 -641 250438
rect -607 250512 -591 250546
rect -237 250512 -221 250546
rect -607 250404 -591 250438
rect -237 250404 -221 250438
rect -187 250512 -171 250546
rect 183 250512 199 250546
rect -187 250404 -171 250438
rect 183 250404 199 250438
rect 233 250512 249 250546
rect 603 250512 619 250546
rect 233 250404 249 250438
rect 603 250404 619 250438
rect 653 250512 669 250546
rect 1023 250512 1039 250546
rect 653 250404 669 250438
rect 1023 250404 1039 250438
rect 1073 250512 1089 250546
rect 1443 250512 1459 250546
rect 1073 250404 1089 250438
rect 1443 250404 1459 250438
rect 1493 250512 1509 250546
rect 1863 250512 1879 250546
rect 1493 250404 1509 250438
rect 1863 250404 1879 250438
rect 1913 250512 1929 250546
rect 2283 250512 2299 250546
rect 1913 250404 1929 250438
rect 2283 250404 2299 250438
rect 2333 250512 2349 250546
rect 2703 250512 2719 250546
rect 2333 250404 2349 250438
rect 2703 250404 2719 250438
rect 2753 250512 2769 250546
rect 3123 250512 3139 250546
rect 2753 250404 2769 250438
rect 3123 250404 3139 250438
rect 3173 250512 3189 250546
rect 3543 250512 3559 250546
rect 3173 250404 3189 250438
rect 3543 250404 3559 250438
rect 3593 250512 3609 250546
rect 3963 250512 3979 250546
rect 3593 250404 3609 250438
rect 3963 250404 3979 250438
rect 4013 250512 4029 250546
rect 4383 250512 4399 250546
rect 4013 250404 4029 250438
rect 4383 250404 4399 250438
rect 4433 250512 4449 250546
rect 4803 250512 4819 250546
rect 4433 250404 4449 250438
rect 4803 250404 4819 250438
rect 4853 250512 4869 250546
rect 5223 250512 5239 250546
rect 4853 250404 4869 250438
rect 5223 250404 5239 250438
rect 5273 250512 5289 250546
rect 5643 250512 5659 250546
rect 5273 250404 5289 250438
rect 5643 250404 5659 250438
rect 5693 250512 5709 250546
rect 6063 250512 6079 250546
rect 5693 250404 5709 250438
rect 6063 250404 6079 250438
rect 6113 250512 6129 250546
rect 6483 250512 6499 250546
rect 6113 250404 6129 250438
rect 6483 250404 6499 250438
rect 6533 250512 6549 250546
rect 6903 250512 6919 250546
rect 6533 250404 6549 250438
rect 6903 250404 6919 250438
rect 6953 250512 6969 250546
rect 7323 250512 7339 250546
rect 6953 250404 6969 250438
rect 7323 250404 7339 250438
rect 7373 250512 7389 250546
rect 7743 250512 7759 250546
rect 7373 250404 7389 250438
rect 7743 250404 7759 250438
rect 7793 250512 7809 250546
rect 8163 250512 8179 250546
rect 7793 250404 7809 250438
rect 8163 250404 8179 250438
rect 8213 250512 8229 250546
rect 8583 250512 8599 250546
rect 8213 250404 8229 250438
rect 8583 250404 8599 250438
rect 8633 250512 8649 250546
rect 9003 250512 9019 250546
rect 8633 250404 8649 250438
rect 9003 250404 9019 250438
rect 9053 250512 9069 250546
rect 9423 250512 9439 250546
rect 9053 250404 9069 250438
rect 9423 250404 9439 250438
rect 9473 250512 9489 250546
rect 9843 250512 9859 250546
rect 9473 250404 9489 250438
rect 9843 250404 9859 250438
rect 9893 250512 9909 250546
rect 10263 250512 10279 250546
rect 9893 250404 9909 250438
rect 10263 250404 10279 250438
rect 10313 250512 10329 250546
rect 10683 250512 10699 250546
rect 10313 250404 10329 250438
rect 10683 250404 10699 250438
rect 10733 250512 10749 250546
rect 11103 250512 11119 250546
rect 10733 250404 10749 250438
rect 11103 250404 11119 250438
rect 11153 250512 11169 250546
rect 11523 250512 11539 250546
rect 11153 250404 11169 250438
rect 11523 250404 11539 250438
rect 11573 250512 11589 250546
rect 11943 250512 11959 250546
rect 11573 250404 11589 250438
rect 11943 250404 11959 250438
rect 11993 250512 12009 250546
rect 12363 250512 12379 250546
rect 11993 250404 12009 250438
rect 12363 250404 12379 250438
rect 12413 250512 12429 250546
rect 12783 250512 12799 250546
rect 12413 250404 12429 250438
rect 12783 250404 12799 250438
rect 12833 250512 12849 250546
rect 13203 250512 13219 250546
rect 12833 250404 12849 250438
rect 13203 250404 13219 250438
rect 13253 250512 13269 250546
rect 13623 250512 13639 250546
rect 13253 250404 13269 250438
rect 13623 250404 13639 250438
rect 13673 250512 13689 250546
rect 14043 250512 14059 250546
rect 13673 250404 13689 250438
rect 14043 250404 14059 250438
rect 14093 250512 14109 250546
rect 14463 250512 14479 250546
rect 14093 250404 14109 250438
rect 14463 250404 14479 250438
rect 14513 250512 14529 250546
rect 14883 250512 14899 250546
rect 14513 250404 14529 250438
rect 14883 250404 14899 250438
rect 14933 250512 14949 250546
rect 15303 250512 15319 250546
rect 14933 250404 14949 250438
rect 15303 250404 15319 250438
rect 15353 250512 15369 250546
rect 15723 250512 15739 250546
rect 15353 250404 15369 250438
rect 15723 250404 15739 250438
rect 15773 250512 15789 250546
rect 16143 250512 16159 250546
rect 15773 250404 15789 250438
rect 16143 250404 16159 250438
rect 16193 250512 16209 250546
rect 16563 250512 16579 250546
rect 16193 250404 16209 250438
rect 16563 250404 16579 250438
rect 16613 250512 16629 250546
rect 16983 250512 16999 250546
rect 16613 250404 16629 250438
rect 16983 250404 16999 250438
rect 17033 250512 17049 250546
rect 17403 250512 17419 250546
rect 17033 250404 17049 250438
rect 17403 250404 17419 250438
rect 17453 250512 17469 250546
rect 17823 250512 17839 250546
rect 17453 250404 17469 250438
rect 17823 250404 17839 250438
rect 17873 250512 17889 250546
rect 18243 250512 18259 250546
rect 17873 250404 17889 250438
rect 18243 250404 18259 250438
rect 18293 250512 18309 250546
rect 18663 250512 18679 250546
rect 18293 250404 18309 250438
rect 18663 250404 18679 250438
rect 18713 250512 18729 250546
rect 19083 250512 19099 250546
rect 18713 250404 18729 250438
rect 19083 250404 19099 250438
rect 19133 250512 19149 250546
rect 19503 250512 19519 250546
rect 19133 250404 19149 250438
rect 19503 250404 19519 250438
rect 19553 250512 19569 250546
rect 19923 250512 19939 250546
rect 19553 250404 19569 250438
rect 19923 250404 19939 250438
rect 19973 250512 19989 250546
rect 20343 250512 20359 250546
rect 19973 250404 19989 250438
rect 20343 250404 20359 250438
rect 20393 250512 20409 250546
rect 20763 250512 20779 250546
rect 20393 250404 20409 250438
rect 20763 250404 20779 250438
rect 20813 250512 20829 250546
rect 21183 250512 21199 250546
rect 20813 250404 20829 250438
rect 21183 250404 21199 250438
rect 21233 250512 21249 250546
rect 21603 250512 21619 250546
rect 21233 250404 21249 250438
rect 21603 250404 21619 250438
rect 21653 250512 21669 250546
rect 22023 250512 22039 250546
rect 21653 250404 21669 250438
rect 22023 250404 22039 250438
rect 22073 250512 22089 250546
rect 22443 250512 22459 250546
rect 22073 250404 22089 250438
rect 22443 250404 22459 250438
rect 22493 250512 22509 250546
rect 22863 250512 22879 250546
rect 22493 250404 22509 250438
rect 22863 250404 22879 250438
rect 22913 250512 22929 250546
rect 23283 250512 23299 250546
rect 22913 250404 22929 250438
rect 23283 250404 23299 250438
rect 23333 250512 23349 250546
rect 23703 250512 23719 250546
rect 23333 250404 23349 250438
rect 23703 250404 23719 250438
rect 23753 250512 23769 250546
rect 24123 250512 24139 250546
rect 23753 250404 23769 250438
rect 24123 250404 24139 250438
rect 24173 250512 24189 250546
rect 24543 250512 24559 250546
rect 24173 250404 24189 250438
rect 24543 250404 24559 250438
rect 24593 250512 24609 250546
rect 24963 250512 24979 250546
rect 24593 250404 24609 250438
rect 24963 250404 24979 250438
rect 25013 250512 25029 250546
rect 25383 250512 25399 250546
rect 25013 250404 25029 250438
rect 25383 250404 25399 250438
rect 25433 250512 25449 250546
rect 25803 250512 25819 250546
rect 25433 250404 25449 250438
rect 25803 250404 25819 250438
rect 25853 250512 25869 250546
rect 26223 250512 26239 250546
rect 25853 250404 25869 250438
rect 26223 250404 26239 250438
rect 26273 250512 26289 250546
rect 26643 250512 26659 250546
rect 26273 250404 26289 250438
rect 26643 250404 26659 250438
rect 26693 250512 26709 250546
rect 27063 250512 27079 250546
rect 26693 250404 26709 250438
rect 27063 250404 27079 250438
rect 27113 250512 27129 250546
rect 27113 250404 27129 250438
rect -4049 250345 -4015 250361
rect -4049 249553 -4015 249569
rect -3953 250345 -3919 250361
rect -3953 249553 -3919 249569
rect -3839 250345 -3805 250361
rect -3839 249553 -3805 249569
rect -3743 250345 -3709 250361
rect -3743 249553 -3709 249569
rect -3629 250345 -3595 250361
rect -3629 249553 -3595 249569
rect -3533 250345 -3499 250361
rect -3533 249553 -3499 249569
rect -3419 250345 -3385 250361
rect -3419 249553 -3385 249569
rect -3323 250345 -3289 250361
rect -3323 249553 -3289 249569
rect -3209 250345 -3175 250361
rect -3209 249553 -3175 249569
rect -3113 250345 -3079 250361
rect -3113 249553 -3079 249569
rect -2999 250345 -2965 250361
rect -2999 249553 -2965 249569
rect -2903 250345 -2869 250361
rect -2903 249553 -2869 249569
rect -2789 250345 -2755 250361
rect -2789 249553 -2755 249569
rect -2693 250345 -2659 250361
rect -2693 249553 -2659 249569
rect -2579 250345 -2545 250361
rect -2579 249553 -2545 249569
rect -2483 250345 -2449 250361
rect -2483 249553 -2449 249569
rect -2369 250345 -2335 250361
rect -2369 249553 -2335 249569
rect -2273 250345 -2239 250361
rect -2273 249553 -2239 249569
rect -2159 250345 -2125 250361
rect -2159 249553 -2125 249569
rect -2063 250345 -2029 250361
rect -2063 249553 -2029 249569
rect -1949 250345 -1915 250361
rect -1949 249553 -1915 249569
rect -1853 250345 -1819 250361
rect -1853 249553 -1819 249569
rect -1739 250345 -1705 250361
rect -1739 249553 -1705 249569
rect -1643 250345 -1609 250361
rect -1643 249553 -1609 249569
rect -1529 250345 -1495 250361
rect -1529 249553 -1495 249569
rect -1433 250345 -1399 250361
rect -1433 249553 -1399 249569
rect -1319 250345 -1285 250361
rect -1319 249553 -1285 249569
rect -1223 250345 -1189 250361
rect -1223 249553 -1189 249569
rect -1109 250345 -1075 250361
rect -1109 249553 -1075 249569
rect -1013 250345 -979 250361
rect -1013 249553 -979 249569
rect -899 250345 -865 250361
rect -899 249553 -865 249569
rect -803 250345 -769 250361
rect -803 249553 -769 249569
rect -689 250345 -655 250361
rect -689 249553 -655 249569
rect -593 250345 -559 250361
rect -593 249553 -559 249569
rect -479 250345 -445 250361
rect -479 249553 -445 249569
rect -383 250345 -349 250361
rect -383 249553 -349 249569
rect -269 250345 -235 250361
rect -269 249553 -235 249569
rect -173 250345 -139 250361
rect -173 249553 -139 249569
rect -59 250345 -25 250361
rect -59 249553 -25 249569
rect 37 250345 71 250361
rect 37 249553 71 249569
rect 151 250345 185 250361
rect 151 249553 185 249569
rect 247 250345 281 250361
rect 247 249553 281 249569
rect 361 250345 395 250361
rect 361 249553 395 249569
rect 457 250345 491 250361
rect 457 249553 491 249569
rect 571 250345 605 250361
rect 571 249553 605 249569
rect 667 250345 701 250361
rect 667 249553 701 249569
rect 781 250345 815 250361
rect 781 249553 815 249569
rect 877 250345 911 250361
rect 877 249553 911 249569
rect 991 250345 1025 250361
rect 991 249553 1025 249569
rect 1087 250345 1121 250361
rect 1087 249553 1121 249569
rect 1201 250345 1235 250361
rect 1201 249553 1235 249569
rect 1297 250345 1331 250361
rect 1297 249553 1331 249569
rect 1411 250345 1445 250361
rect 1411 249553 1445 249569
rect 1507 250345 1541 250361
rect 1507 249553 1541 249569
rect 1621 250345 1655 250361
rect 1621 249553 1655 249569
rect 1717 250345 1751 250361
rect 1717 249553 1751 249569
rect 1831 250345 1865 250361
rect 1831 249553 1865 249569
rect 1927 250345 1961 250361
rect 1927 249553 1961 249569
rect 2041 250345 2075 250361
rect 2041 249553 2075 249569
rect 2137 250345 2171 250361
rect 2137 249553 2171 249569
rect 2251 250345 2285 250361
rect 2251 249553 2285 249569
rect 2347 250345 2381 250361
rect 2347 249553 2381 249569
rect 2461 250345 2495 250361
rect 2461 249553 2495 249569
rect 2557 250345 2591 250361
rect 2557 249553 2591 249569
rect 2671 250345 2705 250361
rect 2671 249553 2705 249569
rect 2767 250345 2801 250361
rect 2767 249553 2801 249569
rect 2881 250345 2915 250361
rect 2881 249553 2915 249569
rect 2977 250345 3011 250361
rect 2977 249553 3011 249569
rect 3091 250345 3125 250361
rect 3091 249553 3125 249569
rect 3187 250345 3221 250361
rect 3187 249553 3221 249569
rect 3301 250345 3335 250361
rect 3301 249553 3335 249569
rect 3397 250345 3431 250361
rect 3397 249553 3431 249569
rect 3511 250345 3545 250361
rect 3511 249553 3545 249569
rect 3607 250345 3641 250361
rect 3607 249553 3641 249569
rect 3721 250345 3755 250361
rect 3721 249553 3755 249569
rect 3817 250345 3851 250361
rect 3817 249553 3851 249569
rect 3931 250345 3965 250361
rect 3931 249553 3965 249569
rect 4027 250345 4061 250361
rect 4027 249553 4061 249569
rect 4141 250345 4175 250361
rect 4141 249553 4175 249569
rect 4237 250345 4271 250361
rect 4237 249553 4271 249569
rect 4351 250345 4385 250361
rect 4351 249553 4385 249569
rect 4447 250345 4481 250361
rect 4447 249553 4481 249569
rect 4561 250345 4595 250361
rect 4561 249553 4595 249569
rect 4657 250345 4691 250361
rect 4657 249553 4691 249569
rect 4771 250345 4805 250361
rect 4771 249553 4805 249569
rect 4867 250345 4901 250361
rect 4867 249553 4901 249569
rect 4981 250345 5015 250361
rect 4981 249553 5015 249569
rect 5077 250345 5111 250361
rect 5077 249553 5111 249569
rect 5191 250345 5225 250361
rect 5191 249553 5225 249569
rect 5287 250345 5321 250361
rect 5287 249553 5321 249569
rect 5401 250345 5435 250361
rect 5401 249553 5435 249569
rect 5497 250345 5531 250361
rect 5497 249553 5531 249569
rect 5611 250345 5645 250361
rect 5611 249553 5645 249569
rect 5707 250345 5741 250361
rect 5707 249553 5741 249569
rect 5821 250345 5855 250361
rect 5821 249553 5855 249569
rect 5917 250345 5951 250361
rect 5917 249553 5951 249569
rect 6031 250345 6065 250361
rect 6031 249553 6065 249569
rect 6127 250345 6161 250361
rect 6127 249553 6161 249569
rect 6241 250345 6275 250361
rect 6241 249553 6275 249569
rect 6337 250345 6371 250361
rect 6337 249553 6371 249569
rect 6451 250345 6485 250361
rect 6451 249553 6485 249569
rect 6547 250345 6581 250361
rect 6547 249553 6581 249569
rect 6661 250345 6695 250361
rect 6661 249553 6695 249569
rect 6757 250345 6791 250361
rect 6757 249553 6791 249569
rect 6871 250345 6905 250361
rect 6871 249553 6905 249569
rect 6967 250345 7001 250361
rect 6967 249553 7001 249569
rect 7081 250345 7115 250361
rect 7081 249553 7115 249569
rect 7177 250345 7211 250361
rect 7177 249553 7211 249569
rect 7291 250345 7325 250361
rect 7291 249553 7325 249569
rect 7387 250345 7421 250361
rect 7387 249553 7421 249569
rect 7501 250345 7535 250361
rect 7501 249553 7535 249569
rect 7597 250345 7631 250361
rect 7597 249553 7631 249569
rect 7711 250345 7745 250361
rect 7711 249553 7745 249569
rect 7807 250345 7841 250361
rect 7807 249553 7841 249569
rect 7921 250345 7955 250361
rect 7921 249553 7955 249569
rect 8017 250345 8051 250361
rect 8017 249553 8051 249569
rect 8131 250345 8165 250361
rect 8131 249553 8165 249569
rect 8227 250345 8261 250361
rect 8227 249553 8261 249569
rect 8341 250345 8375 250361
rect 8341 249553 8375 249569
rect 8437 250345 8471 250361
rect 8437 249553 8471 249569
rect 8551 250345 8585 250361
rect 8551 249553 8585 249569
rect 8647 250345 8681 250361
rect 8647 249553 8681 249569
rect 8761 250345 8795 250361
rect 8761 249553 8795 249569
rect 8857 250345 8891 250361
rect 8857 249553 8891 249569
rect 8971 250345 9005 250361
rect 8971 249553 9005 249569
rect 9067 250345 9101 250361
rect 9067 249553 9101 249569
rect 9181 250345 9215 250361
rect 9181 249553 9215 249569
rect 9277 250345 9311 250361
rect 9277 249553 9311 249569
rect 9391 250345 9425 250361
rect 9391 249553 9425 249569
rect 9487 250345 9521 250361
rect 9487 249553 9521 249569
rect 9601 250345 9635 250361
rect 9601 249553 9635 249569
rect 9697 250345 9731 250361
rect 9697 249553 9731 249569
rect 9811 250345 9845 250361
rect 9811 249553 9845 249569
rect 9907 250345 9941 250361
rect 9907 249553 9941 249569
rect 10021 250345 10055 250361
rect 10021 249553 10055 249569
rect 10117 250345 10151 250361
rect 10117 249553 10151 249569
rect 10231 250345 10265 250361
rect 10231 249553 10265 249569
rect 10327 250345 10361 250361
rect 10327 249553 10361 249569
rect 10441 250345 10475 250361
rect 10441 249553 10475 249569
rect 10537 250345 10571 250361
rect 10537 249553 10571 249569
rect 10651 250345 10685 250361
rect 10651 249553 10685 249569
rect 10747 250345 10781 250361
rect 10747 249553 10781 249569
rect 10861 250345 10895 250361
rect 10861 249553 10895 249569
rect 10957 250345 10991 250361
rect 10957 249553 10991 249569
rect 11071 250345 11105 250361
rect 11071 249553 11105 249569
rect 11167 250345 11201 250361
rect 11167 249553 11201 249569
rect 11281 250345 11315 250361
rect 11281 249553 11315 249569
rect 11377 250345 11411 250361
rect 11377 249553 11411 249569
rect 11491 250345 11525 250361
rect 11491 249553 11525 249569
rect 11587 250345 11621 250361
rect 11587 249553 11621 249569
rect 11701 250345 11735 250361
rect 11701 249553 11735 249569
rect 11797 250345 11831 250361
rect 11797 249553 11831 249569
rect 11911 250345 11945 250361
rect 11911 249553 11945 249569
rect 12007 250345 12041 250361
rect 12007 249553 12041 249569
rect 12121 250345 12155 250361
rect 12121 249553 12155 249569
rect 12217 250345 12251 250361
rect 12217 249553 12251 249569
rect 12331 250345 12365 250361
rect 12331 249553 12365 249569
rect 12427 250345 12461 250361
rect 12427 249553 12461 249569
rect 12541 250345 12575 250361
rect 12541 249553 12575 249569
rect 12637 250345 12671 250361
rect 12637 249553 12671 249569
rect 12751 250345 12785 250361
rect 12751 249553 12785 249569
rect 12847 250345 12881 250361
rect 12847 249553 12881 249569
rect 12961 250345 12995 250361
rect 12961 249553 12995 249569
rect 13057 250345 13091 250361
rect 13057 249553 13091 249569
rect 13171 250345 13205 250361
rect 13171 249553 13205 249569
rect 13267 250345 13301 250361
rect 13267 249553 13301 249569
rect 13381 250345 13415 250361
rect 13381 249553 13415 249569
rect 13477 250345 13511 250361
rect 13477 249553 13511 249569
rect 13591 250345 13625 250361
rect 13591 249553 13625 249569
rect 13687 250345 13721 250361
rect 13687 249553 13721 249569
rect 13801 250345 13835 250361
rect 13801 249553 13835 249569
rect 13897 250345 13931 250361
rect 13897 249553 13931 249569
rect 14011 250345 14045 250361
rect 14011 249553 14045 249569
rect 14107 250345 14141 250361
rect 14107 249553 14141 249569
rect 14221 250345 14255 250361
rect 14221 249553 14255 249569
rect 14317 250345 14351 250361
rect 14317 249553 14351 249569
rect 14431 250345 14465 250361
rect 14431 249553 14465 249569
rect 14527 250345 14561 250361
rect 14527 249553 14561 249569
rect 14641 250345 14675 250361
rect 14641 249553 14675 249569
rect 14737 250345 14771 250361
rect 14737 249553 14771 249569
rect 14851 250345 14885 250361
rect 14851 249553 14885 249569
rect 14947 250345 14981 250361
rect 14947 249553 14981 249569
rect 15061 250345 15095 250361
rect 15061 249553 15095 249569
rect 15157 250345 15191 250361
rect 15157 249553 15191 249569
rect 15271 250345 15305 250361
rect 15271 249553 15305 249569
rect 15367 250345 15401 250361
rect 15367 249553 15401 249569
rect 15481 250345 15515 250361
rect 15481 249553 15515 249569
rect 15577 250345 15611 250361
rect 15577 249553 15611 249569
rect 15691 250345 15725 250361
rect 15691 249553 15725 249569
rect 15787 250345 15821 250361
rect 15787 249553 15821 249569
rect 15901 250345 15935 250361
rect 15901 249553 15935 249569
rect 15997 250345 16031 250361
rect 15997 249553 16031 249569
rect 16111 250345 16145 250361
rect 16111 249553 16145 249569
rect 16207 250345 16241 250361
rect 16207 249553 16241 249569
rect 16321 250345 16355 250361
rect 16321 249553 16355 249569
rect 16417 250345 16451 250361
rect 16417 249553 16451 249569
rect 16531 250345 16565 250361
rect 16531 249553 16565 249569
rect 16627 250345 16661 250361
rect 16627 249553 16661 249569
rect 16741 250345 16775 250361
rect 16741 249553 16775 249569
rect 16837 250345 16871 250361
rect 16837 249553 16871 249569
rect 16951 250345 16985 250361
rect 16951 249553 16985 249569
rect 17047 250345 17081 250361
rect 17047 249553 17081 249569
rect 17161 250345 17195 250361
rect 17161 249553 17195 249569
rect 17257 250345 17291 250361
rect 17257 249553 17291 249569
rect 17371 250345 17405 250361
rect 17371 249553 17405 249569
rect 17467 250345 17501 250361
rect 17467 249553 17501 249569
rect 17581 250345 17615 250361
rect 17581 249553 17615 249569
rect 17677 250345 17711 250361
rect 17677 249553 17711 249569
rect 17791 250345 17825 250361
rect 17791 249553 17825 249569
rect 17887 250345 17921 250361
rect 17887 249553 17921 249569
rect 18001 250345 18035 250361
rect 18001 249553 18035 249569
rect 18097 250345 18131 250361
rect 18097 249553 18131 249569
rect 18211 250345 18245 250361
rect 18211 249553 18245 249569
rect 18307 250345 18341 250361
rect 18307 249553 18341 249569
rect 18421 250345 18455 250361
rect 18421 249553 18455 249569
rect 18517 250345 18551 250361
rect 18517 249553 18551 249569
rect 18631 250345 18665 250361
rect 18631 249553 18665 249569
rect 18727 250345 18761 250361
rect 18727 249553 18761 249569
rect 18841 250345 18875 250361
rect 18841 249553 18875 249569
rect 18937 250345 18971 250361
rect 18937 249553 18971 249569
rect 19051 250345 19085 250361
rect 19051 249553 19085 249569
rect 19147 250345 19181 250361
rect 19147 249553 19181 249569
rect 19261 250345 19295 250361
rect 19261 249553 19295 249569
rect 19357 250345 19391 250361
rect 19357 249553 19391 249569
rect 19471 250345 19505 250361
rect 19471 249553 19505 249569
rect 19567 250345 19601 250361
rect 19567 249553 19601 249569
rect 19681 250345 19715 250361
rect 19681 249553 19715 249569
rect 19777 250345 19811 250361
rect 19777 249553 19811 249569
rect 19891 250345 19925 250361
rect 19891 249553 19925 249569
rect 19987 250345 20021 250361
rect 19987 249553 20021 249569
rect 20101 250345 20135 250361
rect 20101 249553 20135 249569
rect 20197 250345 20231 250361
rect 20197 249553 20231 249569
rect 20311 250345 20345 250361
rect 20311 249553 20345 249569
rect 20407 250345 20441 250361
rect 20407 249553 20441 249569
rect 20521 250345 20555 250361
rect 20521 249553 20555 249569
rect 20617 250345 20651 250361
rect 20617 249553 20651 249569
rect 20731 250345 20765 250361
rect 20731 249553 20765 249569
rect 20827 250345 20861 250361
rect 20827 249553 20861 249569
rect 20941 250345 20975 250361
rect 20941 249553 20975 249569
rect 21037 250345 21071 250361
rect 21037 249553 21071 249569
rect 21151 250345 21185 250361
rect 21151 249553 21185 249569
rect 21247 250345 21281 250361
rect 21247 249553 21281 249569
rect 21361 250345 21395 250361
rect 21361 249553 21395 249569
rect 21457 250345 21491 250361
rect 21457 249553 21491 249569
rect 21571 250345 21605 250361
rect 21571 249553 21605 249569
rect 21667 250345 21701 250361
rect 21667 249553 21701 249569
rect 21781 250345 21815 250361
rect 21781 249553 21815 249569
rect 21877 250345 21911 250361
rect 21877 249553 21911 249569
rect 21991 250345 22025 250361
rect 21991 249553 22025 249569
rect 22087 250345 22121 250361
rect 22087 249553 22121 249569
rect 22201 250345 22235 250361
rect 22201 249553 22235 249569
rect 22297 250345 22331 250361
rect 22297 249553 22331 249569
rect 22411 250345 22445 250361
rect 22411 249553 22445 249569
rect 22507 250345 22541 250361
rect 22507 249553 22541 249569
rect 22621 250345 22655 250361
rect 22621 249553 22655 249569
rect 22717 250345 22751 250361
rect 22717 249553 22751 249569
rect 22831 250345 22865 250361
rect 22831 249553 22865 249569
rect 22927 250345 22961 250361
rect 22927 249553 22961 249569
rect 23041 250345 23075 250361
rect 23041 249553 23075 249569
rect 23137 250345 23171 250361
rect 23137 249553 23171 249569
rect 23251 250345 23285 250361
rect 23251 249553 23285 249569
rect 23347 250345 23381 250361
rect 23347 249553 23381 249569
rect 23461 250345 23495 250361
rect 23461 249553 23495 249569
rect 23557 250345 23591 250361
rect 23557 249553 23591 249569
rect 23671 250345 23705 250361
rect 23671 249553 23705 249569
rect 23767 250345 23801 250361
rect 23767 249553 23801 249569
rect 23881 250345 23915 250361
rect 23881 249553 23915 249569
rect 23977 250345 24011 250361
rect 23977 249553 24011 249569
rect 24091 250345 24125 250361
rect 24091 249553 24125 249569
rect 24187 250345 24221 250361
rect 24187 249553 24221 249569
rect 24301 250345 24335 250361
rect 24301 249553 24335 249569
rect 24397 250345 24431 250361
rect 24397 249553 24431 249569
rect 24511 250345 24545 250361
rect 24511 249553 24545 249569
rect 24607 250345 24641 250361
rect 24607 249553 24641 249569
rect 24721 250345 24755 250361
rect 24721 249553 24755 249569
rect 24817 250345 24851 250361
rect 24817 249553 24851 249569
rect 24931 250345 24965 250361
rect 24931 249553 24965 249569
rect 25027 250345 25061 250361
rect 25027 249553 25061 249569
rect 25141 250345 25175 250361
rect 25141 249553 25175 249569
rect 25237 250345 25271 250361
rect 25237 249553 25271 249569
rect 25351 250345 25385 250361
rect 25351 249553 25385 249569
rect 25447 250345 25481 250361
rect 25447 249553 25481 249569
rect 25561 250345 25595 250361
rect 25561 249553 25595 249569
rect 25657 250345 25691 250361
rect 25657 249553 25691 249569
rect 25771 250345 25805 250361
rect 25771 249553 25805 249569
rect 25867 250345 25901 250361
rect 25867 249553 25901 249569
rect 25981 250345 26015 250361
rect 25981 249553 26015 249569
rect 26077 250345 26111 250361
rect 26077 249553 26111 249569
rect 26191 250345 26225 250361
rect 26191 249553 26225 249569
rect 26287 250345 26321 250361
rect 26287 249553 26321 249569
rect 26401 250345 26435 250361
rect 26401 249553 26435 249569
rect 26497 250345 26531 250361
rect 26497 249553 26531 249569
rect 26611 250345 26645 250361
rect 26611 249553 26645 249569
rect 26707 250345 26741 250361
rect 26707 249553 26741 249569
rect 26821 250345 26855 250361
rect 26821 249553 26855 249569
rect 26917 250345 26951 250361
rect 26917 249553 26951 249569
rect 27031 250345 27065 250361
rect 27031 249553 27065 249569
rect 27127 250345 27161 250361
rect 27127 249553 27161 249569
rect 27241 250345 27275 250361
rect 27241 249553 27275 249569
rect 27337 250345 27371 250361
rect 27337 249553 27371 249569
rect -3807 249476 -3791 249510
rect -3695 249476 -3679 249510
rect -3387 249476 -3371 249510
rect -3275 249476 -3259 249510
rect -2967 249476 -2951 249510
rect -2855 249476 -2839 249510
rect -2547 249476 -2531 249510
rect -2435 249476 -2419 249510
rect -2127 249476 -2111 249510
rect -2015 249476 -1999 249510
rect -1707 249476 -1691 249510
rect -1595 249476 -1579 249510
rect -1287 249476 -1271 249510
rect -1175 249476 -1159 249510
rect -867 249476 -851 249510
rect -755 249476 -739 249510
rect -447 249476 -431 249510
rect -335 249476 -319 249510
rect -27 249476 -11 249510
rect 85 249476 101 249510
rect 393 249476 409 249510
rect 505 249476 521 249510
rect 813 249476 829 249510
rect 925 249476 941 249510
rect 1233 249476 1249 249510
rect 1345 249476 1361 249510
rect 1653 249476 1669 249510
rect 1765 249476 1781 249510
rect 2073 249476 2089 249510
rect 2185 249476 2201 249510
rect 2493 249476 2509 249510
rect 2605 249476 2621 249510
rect 2913 249476 2929 249510
rect 3025 249476 3041 249510
rect 3333 249476 3349 249510
rect 3445 249476 3461 249510
rect 3753 249476 3769 249510
rect 3865 249476 3881 249510
rect 4173 249476 4189 249510
rect 4285 249476 4301 249510
rect 4593 249476 4609 249510
rect 4705 249476 4721 249510
rect 5013 249476 5029 249510
rect 5125 249476 5141 249510
rect 5433 249476 5449 249510
rect 5545 249476 5561 249510
rect 5853 249476 5869 249510
rect 5965 249476 5981 249510
rect 6273 249476 6289 249510
rect 6385 249476 6401 249510
rect 6693 249476 6709 249510
rect 6805 249476 6821 249510
rect 7113 249476 7129 249510
rect 7225 249476 7241 249510
rect 7533 249476 7549 249510
rect 7645 249476 7661 249510
rect 7953 249476 7969 249510
rect 8065 249476 8081 249510
rect 8373 249476 8389 249510
rect 8485 249476 8501 249510
rect 8793 249476 8809 249510
rect 8905 249476 8921 249510
rect 9213 249476 9229 249510
rect 9325 249476 9341 249510
rect 9633 249476 9649 249510
rect 9745 249476 9761 249510
rect 10053 249476 10069 249510
rect 10165 249476 10181 249510
rect 10473 249476 10489 249510
rect 10585 249476 10601 249510
rect 10893 249476 10909 249510
rect 11005 249476 11021 249510
rect 11313 249476 11329 249510
rect 11425 249476 11441 249510
rect 11733 249476 11749 249510
rect 11845 249476 11861 249510
rect 12153 249476 12169 249510
rect 12265 249476 12281 249510
rect 12573 249476 12589 249510
rect 12685 249476 12701 249510
rect 12993 249476 13009 249510
rect 13105 249476 13121 249510
rect 13413 249476 13429 249510
rect 13525 249476 13541 249510
rect 13833 249476 13849 249510
rect 13945 249476 13961 249510
rect 14253 249476 14269 249510
rect 14365 249476 14381 249510
rect 14673 249476 14689 249510
rect 14785 249476 14801 249510
rect 15093 249476 15109 249510
rect 15205 249476 15221 249510
rect 15513 249476 15529 249510
rect 15625 249476 15641 249510
rect 15933 249476 15949 249510
rect 16045 249476 16061 249510
rect 16353 249476 16369 249510
rect 16465 249476 16481 249510
rect 16773 249476 16789 249510
rect 16885 249476 16901 249510
rect 17193 249476 17209 249510
rect 17305 249476 17321 249510
rect 17613 249476 17629 249510
rect 17725 249476 17741 249510
rect 18033 249476 18049 249510
rect 18145 249476 18161 249510
rect 18453 249476 18469 249510
rect 18565 249476 18581 249510
rect 18873 249476 18889 249510
rect 18985 249476 19001 249510
rect 19293 249476 19309 249510
rect 19405 249476 19421 249510
rect 19713 249476 19729 249510
rect 19825 249476 19841 249510
rect 20133 249476 20149 249510
rect 20245 249476 20261 249510
rect 20553 249476 20569 249510
rect 20665 249476 20681 249510
rect 20973 249476 20989 249510
rect 21085 249476 21101 249510
rect 21393 249476 21409 249510
rect 21505 249476 21521 249510
rect 21813 249476 21829 249510
rect 21925 249476 21941 249510
rect 22233 249476 22249 249510
rect 22345 249476 22361 249510
rect 22653 249476 22669 249510
rect 22765 249476 22781 249510
rect 23073 249476 23089 249510
rect 23185 249476 23201 249510
rect 23493 249476 23509 249510
rect 23605 249476 23621 249510
rect 23913 249476 23929 249510
rect 24025 249476 24041 249510
rect 24333 249476 24349 249510
rect 24445 249476 24461 249510
rect 24753 249476 24769 249510
rect 24865 249476 24881 249510
rect 25173 249476 25189 249510
rect 25285 249476 25301 249510
rect 25593 249476 25609 249510
rect 25705 249476 25721 249510
rect 26013 249476 26029 249510
rect 26125 249476 26141 249510
rect 26433 249476 26449 249510
rect 26545 249476 26561 249510
rect 26853 249476 26869 249510
rect 26965 249476 26981 249510
rect 27273 249476 27289 249510
rect 27385 249476 27401 249510
rect -4163 249408 -4129 249470
rect 27451 249408 27485 249470
rect -4163 249341 -4067 249408
rect 27389 249375 27485 249408
rect 27389 249341 27485 249374
rect -4163 249279 -4129 249341
rect 27451 249279 27485 249341
rect -4017 249239 -4001 249273
rect -3905 249239 -3889 249273
rect -3597 249239 -3581 249273
rect -3485 249239 -3469 249273
rect -3177 249239 -3161 249273
rect -3065 249239 -3049 249273
rect -2757 249239 -2741 249273
rect -2645 249239 -2629 249273
rect -2337 249239 -2321 249273
rect -2225 249239 -2209 249273
rect -1917 249239 -1901 249273
rect -1805 249239 -1789 249273
rect -1497 249239 -1481 249273
rect -1385 249239 -1369 249273
rect -1077 249239 -1061 249273
rect -965 249239 -949 249273
rect -657 249239 -641 249273
rect -545 249239 -529 249273
rect -237 249239 -221 249273
rect -125 249239 -109 249273
rect 183 249239 199 249273
rect 295 249239 311 249273
rect 603 249239 619 249273
rect 715 249239 731 249273
rect 1023 249239 1039 249273
rect 1135 249239 1151 249273
rect 1443 249239 1459 249273
rect 1555 249239 1571 249273
rect 1863 249239 1879 249273
rect 1975 249239 1991 249273
rect 2283 249239 2299 249273
rect 2395 249239 2411 249273
rect 2703 249239 2719 249273
rect 2815 249239 2831 249273
rect 3123 249239 3139 249273
rect 3235 249239 3251 249273
rect 3543 249239 3559 249273
rect 3655 249239 3671 249273
rect 3963 249239 3979 249273
rect 4075 249239 4091 249273
rect 4383 249239 4399 249273
rect 4495 249239 4511 249273
rect 4803 249239 4819 249273
rect 4915 249239 4931 249273
rect 5223 249239 5239 249273
rect 5335 249239 5351 249273
rect 5643 249239 5659 249273
rect 5755 249239 5771 249273
rect 6063 249239 6079 249273
rect 6175 249239 6191 249273
rect 6483 249239 6499 249273
rect 6595 249239 6611 249273
rect 6903 249239 6919 249273
rect 7015 249239 7031 249273
rect 7323 249239 7339 249273
rect 7435 249239 7451 249273
rect 7743 249239 7759 249273
rect 7855 249239 7871 249273
rect 8163 249239 8179 249273
rect 8275 249239 8291 249273
rect 8583 249239 8599 249273
rect 8695 249239 8711 249273
rect 9003 249239 9019 249273
rect 9115 249239 9131 249273
rect 9423 249239 9439 249273
rect 9535 249239 9551 249273
rect 9843 249239 9859 249273
rect 9955 249239 9971 249273
rect 10263 249239 10279 249273
rect 10375 249239 10391 249273
rect 10683 249239 10699 249273
rect 10795 249239 10811 249273
rect 11103 249239 11119 249273
rect 11215 249239 11231 249273
rect 11523 249239 11539 249273
rect 11635 249239 11651 249273
rect 11943 249239 11959 249273
rect 12055 249239 12071 249273
rect 12363 249239 12379 249273
rect 12475 249239 12491 249273
rect 12783 249239 12799 249273
rect 12895 249239 12911 249273
rect 13203 249239 13219 249273
rect 13315 249239 13331 249273
rect 13623 249239 13639 249273
rect 13735 249239 13751 249273
rect 14043 249239 14059 249273
rect 14155 249239 14171 249273
rect 14463 249239 14479 249273
rect 14575 249239 14591 249273
rect 14883 249239 14899 249273
rect 14995 249239 15011 249273
rect 15303 249239 15319 249273
rect 15415 249239 15431 249273
rect 15723 249239 15739 249273
rect 15835 249239 15851 249273
rect 16143 249239 16159 249273
rect 16255 249239 16271 249273
rect 16563 249239 16579 249273
rect 16675 249239 16691 249273
rect 16983 249239 16999 249273
rect 17095 249239 17111 249273
rect 17403 249239 17419 249273
rect 17515 249239 17531 249273
rect 17823 249239 17839 249273
rect 17935 249239 17951 249273
rect 18243 249239 18259 249273
rect 18355 249239 18371 249273
rect 18663 249239 18679 249273
rect 18775 249239 18791 249273
rect 19083 249239 19099 249273
rect 19195 249239 19211 249273
rect 19503 249239 19519 249273
rect 19615 249239 19631 249273
rect 19923 249239 19939 249273
rect 20035 249239 20051 249273
rect 20343 249239 20359 249273
rect 20455 249239 20471 249273
rect 20763 249239 20779 249273
rect 20875 249239 20891 249273
rect 21183 249239 21199 249273
rect 21295 249239 21311 249273
rect 21603 249239 21619 249273
rect 21715 249239 21731 249273
rect 22023 249239 22039 249273
rect 22135 249239 22151 249273
rect 22443 249239 22459 249273
rect 22555 249239 22571 249273
rect 22863 249239 22879 249273
rect 22975 249239 22991 249273
rect 23283 249239 23299 249273
rect 23395 249239 23411 249273
rect 23703 249239 23719 249273
rect 23815 249239 23831 249273
rect 24123 249239 24139 249273
rect 24235 249239 24251 249273
rect 24543 249239 24559 249273
rect 24655 249239 24671 249273
rect 24963 249239 24979 249273
rect 25075 249239 25091 249273
rect 25383 249239 25399 249273
rect 25495 249239 25511 249273
rect 25803 249239 25819 249273
rect 25915 249239 25931 249273
rect 26223 249239 26239 249273
rect 26335 249239 26351 249273
rect 26643 249239 26659 249273
rect 26755 249239 26771 249273
rect 27063 249239 27079 249273
rect 27175 249239 27191 249273
rect -4049 249180 -4015 249196
rect -4049 248388 -4015 248404
rect -3953 249180 -3919 249196
rect -3953 248388 -3919 248404
rect -3839 249180 -3805 249196
rect -3839 248388 -3805 248404
rect -3743 249180 -3709 249196
rect -3743 248388 -3709 248404
rect -3629 249180 -3595 249196
rect -3629 248388 -3595 248404
rect -3533 249180 -3499 249196
rect -3533 248388 -3499 248404
rect -3419 249180 -3385 249196
rect -3419 248388 -3385 248404
rect -3323 249180 -3289 249196
rect -3323 248388 -3289 248404
rect -3209 249180 -3175 249196
rect -3209 248388 -3175 248404
rect -3113 249180 -3079 249196
rect -3113 248388 -3079 248404
rect -2999 249180 -2965 249196
rect -2999 248388 -2965 248404
rect -2903 249180 -2869 249196
rect -2903 248388 -2869 248404
rect -2789 249180 -2755 249196
rect -2789 248388 -2755 248404
rect -2693 249180 -2659 249196
rect -2693 248388 -2659 248404
rect -2579 249180 -2545 249196
rect -2579 248388 -2545 248404
rect -2483 249180 -2449 249196
rect -2483 248388 -2449 248404
rect -2369 249180 -2335 249196
rect -2369 248388 -2335 248404
rect -2273 249180 -2239 249196
rect -2273 248388 -2239 248404
rect -2159 249180 -2125 249196
rect -2159 248388 -2125 248404
rect -2063 249180 -2029 249196
rect -2063 248388 -2029 248404
rect -1949 249180 -1915 249196
rect -1949 248388 -1915 248404
rect -1853 249180 -1819 249196
rect -1853 248388 -1819 248404
rect -1739 249180 -1705 249196
rect -1739 248388 -1705 248404
rect -1643 249180 -1609 249196
rect -1643 248388 -1609 248404
rect -1529 249180 -1495 249196
rect -1529 248388 -1495 248404
rect -1433 249180 -1399 249196
rect -1433 248388 -1399 248404
rect -1319 249180 -1285 249196
rect -1319 248388 -1285 248404
rect -1223 249180 -1189 249196
rect -1223 248388 -1189 248404
rect -1109 249180 -1075 249196
rect -1109 248388 -1075 248404
rect -1013 249180 -979 249196
rect -1013 248388 -979 248404
rect -899 249180 -865 249196
rect -899 248388 -865 248404
rect -803 249180 -769 249196
rect -803 248388 -769 248404
rect -689 249180 -655 249196
rect -689 248388 -655 248404
rect -593 249180 -559 249196
rect -593 248388 -559 248404
rect -479 249180 -445 249196
rect -479 248388 -445 248404
rect -383 249180 -349 249196
rect -383 248388 -349 248404
rect -269 249180 -235 249196
rect -269 248388 -235 248404
rect -173 249180 -139 249196
rect -173 248388 -139 248404
rect -59 249180 -25 249196
rect -59 248388 -25 248404
rect 37 249180 71 249196
rect 37 248388 71 248404
rect 151 249180 185 249196
rect 151 248388 185 248404
rect 247 249180 281 249196
rect 247 248388 281 248404
rect 361 249180 395 249196
rect 361 248388 395 248404
rect 457 249180 491 249196
rect 457 248388 491 248404
rect 571 249180 605 249196
rect 571 248388 605 248404
rect 667 249180 701 249196
rect 667 248388 701 248404
rect 781 249180 815 249196
rect 781 248388 815 248404
rect 877 249180 911 249196
rect 877 248388 911 248404
rect 991 249180 1025 249196
rect 991 248388 1025 248404
rect 1087 249180 1121 249196
rect 1087 248388 1121 248404
rect 1201 249180 1235 249196
rect 1201 248388 1235 248404
rect 1297 249180 1331 249196
rect 1297 248388 1331 248404
rect 1411 249180 1445 249196
rect 1411 248388 1445 248404
rect 1507 249180 1541 249196
rect 1507 248388 1541 248404
rect 1621 249180 1655 249196
rect 1621 248388 1655 248404
rect 1717 249180 1751 249196
rect 1717 248388 1751 248404
rect 1831 249180 1865 249196
rect 1831 248388 1865 248404
rect 1927 249180 1961 249196
rect 1927 248388 1961 248404
rect 2041 249180 2075 249196
rect 2041 248388 2075 248404
rect 2137 249180 2171 249196
rect 2137 248388 2171 248404
rect 2251 249180 2285 249196
rect 2251 248388 2285 248404
rect 2347 249180 2381 249196
rect 2347 248388 2381 248404
rect 2461 249180 2495 249196
rect 2461 248388 2495 248404
rect 2557 249180 2591 249196
rect 2557 248388 2591 248404
rect 2671 249180 2705 249196
rect 2671 248388 2705 248404
rect 2767 249180 2801 249196
rect 2767 248388 2801 248404
rect 2881 249180 2915 249196
rect 2881 248388 2915 248404
rect 2977 249180 3011 249196
rect 2977 248388 3011 248404
rect 3091 249180 3125 249196
rect 3091 248388 3125 248404
rect 3187 249180 3221 249196
rect 3187 248388 3221 248404
rect 3301 249180 3335 249196
rect 3301 248388 3335 248404
rect 3397 249180 3431 249196
rect 3397 248388 3431 248404
rect 3511 249180 3545 249196
rect 3511 248388 3545 248404
rect 3607 249180 3641 249196
rect 3607 248388 3641 248404
rect 3721 249180 3755 249196
rect 3721 248388 3755 248404
rect 3817 249180 3851 249196
rect 3817 248388 3851 248404
rect 3931 249180 3965 249196
rect 3931 248388 3965 248404
rect 4027 249180 4061 249196
rect 4027 248388 4061 248404
rect 4141 249180 4175 249196
rect 4141 248388 4175 248404
rect 4237 249180 4271 249196
rect 4237 248388 4271 248404
rect 4351 249180 4385 249196
rect 4351 248388 4385 248404
rect 4447 249180 4481 249196
rect 4447 248388 4481 248404
rect 4561 249180 4595 249196
rect 4561 248388 4595 248404
rect 4657 249180 4691 249196
rect 4657 248388 4691 248404
rect 4771 249180 4805 249196
rect 4771 248388 4805 248404
rect 4867 249180 4901 249196
rect 4867 248388 4901 248404
rect 4981 249180 5015 249196
rect 4981 248388 5015 248404
rect 5077 249180 5111 249196
rect 5077 248388 5111 248404
rect 5191 249180 5225 249196
rect 5191 248388 5225 248404
rect 5287 249180 5321 249196
rect 5287 248388 5321 248404
rect 5401 249180 5435 249196
rect 5401 248388 5435 248404
rect 5497 249180 5531 249196
rect 5497 248388 5531 248404
rect 5611 249180 5645 249196
rect 5611 248388 5645 248404
rect 5707 249180 5741 249196
rect 5707 248388 5741 248404
rect 5821 249180 5855 249196
rect 5821 248388 5855 248404
rect 5917 249180 5951 249196
rect 5917 248388 5951 248404
rect 6031 249180 6065 249196
rect 6031 248388 6065 248404
rect 6127 249180 6161 249196
rect 6127 248388 6161 248404
rect 6241 249180 6275 249196
rect 6241 248388 6275 248404
rect 6337 249180 6371 249196
rect 6337 248388 6371 248404
rect 6451 249180 6485 249196
rect 6451 248388 6485 248404
rect 6547 249180 6581 249196
rect 6547 248388 6581 248404
rect 6661 249180 6695 249196
rect 6661 248388 6695 248404
rect 6757 249180 6791 249196
rect 6757 248388 6791 248404
rect 6871 249180 6905 249196
rect 6871 248388 6905 248404
rect 6967 249180 7001 249196
rect 6967 248388 7001 248404
rect 7081 249180 7115 249196
rect 7081 248388 7115 248404
rect 7177 249180 7211 249196
rect 7177 248388 7211 248404
rect 7291 249180 7325 249196
rect 7291 248388 7325 248404
rect 7387 249180 7421 249196
rect 7387 248388 7421 248404
rect 7501 249180 7535 249196
rect 7501 248388 7535 248404
rect 7597 249180 7631 249196
rect 7597 248388 7631 248404
rect 7711 249180 7745 249196
rect 7711 248388 7745 248404
rect 7807 249180 7841 249196
rect 7807 248388 7841 248404
rect 7921 249180 7955 249196
rect 7921 248388 7955 248404
rect 8017 249180 8051 249196
rect 8017 248388 8051 248404
rect 8131 249180 8165 249196
rect 8131 248388 8165 248404
rect 8227 249180 8261 249196
rect 8227 248388 8261 248404
rect 8341 249180 8375 249196
rect 8341 248388 8375 248404
rect 8437 249180 8471 249196
rect 8437 248388 8471 248404
rect 8551 249180 8585 249196
rect 8551 248388 8585 248404
rect 8647 249180 8681 249196
rect 8647 248388 8681 248404
rect 8761 249180 8795 249196
rect 8761 248388 8795 248404
rect 8857 249180 8891 249196
rect 8857 248388 8891 248404
rect 8971 249180 9005 249196
rect 8971 248388 9005 248404
rect 9067 249180 9101 249196
rect 9067 248388 9101 248404
rect 9181 249180 9215 249196
rect 9181 248388 9215 248404
rect 9277 249180 9311 249196
rect 9277 248388 9311 248404
rect 9391 249180 9425 249196
rect 9391 248388 9425 248404
rect 9487 249180 9521 249196
rect 9487 248388 9521 248404
rect 9601 249180 9635 249196
rect 9601 248388 9635 248404
rect 9697 249180 9731 249196
rect 9697 248388 9731 248404
rect 9811 249180 9845 249196
rect 9811 248388 9845 248404
rect 9907 249180 9941 249196
rect 9907 248388 9941 248404
rect 10021 249180 10055 249196
rect 10021 248388 10055 248404
rect 10117 249180 10151 249196
rect 10117 248388 10151 248404
rect 10231 249180 10265 249196
rect 10231 248388 10265 248404
rect 10327 249180 10361 249196
rect 10327 248388 10361 248404
rect 10441 249180 10475 249196
rect 10441 248388 10475 248404
rect 10537 249180 10571 249196
rect 10537 248388 10571 248404
rect 10651 249180 10685 249196
rect 10651 248388 10685 248404
rect 10747 249180 10781 249196
rect 10747 248388 10781 248404
rect 10861 249180 10895 249196
rect 10861 248388 10895 248404
rect 10957 249180 10991 249196
rect 10957 248388 10991 248404
rect 11071 249180 11105 249196
rect 11071 248388 11105 248404
rect 11167 249180 11201 249196
rect 11167 248388 11201 248404
rect 11281 249180 11315 249196
rect 11281 248388 11315 248404
rect 11377 249180 11411 249196
rect 11377 248388 11411 248404
rect 11491 249180 11525 249196
rect 11491 248388 11525 248404
rect 11587 249180 11621 249196
rect 11587 248388 11621 248404
rect 11701 249180 11735 249196
rect 11701 248388 11735 248404
rect 11797 249180 11831 249196
rect 11797 248388 11831 248404
rect 11911 249180 11945 249196
rect 11911 248388 11945 248404
rect 12007 249180 12041 249196
rect 12007 248388 12041 248404
rect 12121 249180 12155 249196
rect 12121 248388 12155 248404
rect 12217 249180 12251 249196
rect 12217 248388 12251 248404
rect 12331 249180 12365 249196
rect 12331 248388 12365 248404
rect 12427 249180 12461 249196
rect 12427 248388 12461 248404
rect 12541 249180 12575 249196
rect 12541 248388 12575 248404
rect 12637 249180 12671 249196
rect 12637 248388 12671 248404
rect 12751 249180 12785 249196
rect 12751 248388 12785 248404
rect 12847 249180 12881 249196
rect 12847 248388 12881 248404
rect 12961 249180 12995 249196
rect 12961 248388 12995 248404
rect 13057 249180 13091 249196
rect 13057 248388 13091 248404
rect 13171 249180 13205 249196
rect 13171 248388 13205 248404
rect 13267 249180 13301 249196
rect 13267 248388 13301 248404
rect 13381 249180 13415 249196
rect 13381 248388 13415 248404
rect 13477 249180 13511 249196
rect 13477 248388 13511 248404
rect 13591 249180 13625 249196
rect 13591 248388 13625 248404
rect 13687 249180 13721 249196
rect 13687 248388 13721 248404
rect 13801 249180 13835 249196
rect 13801 248388 13835 248404
rect 13897 249180 13931 249196
rect 13897 248388 13931 248404
rect 14011 249180 14045 249196
rect 14011 248388 14045 248404
rect 14107 249180 14141 249196
rect 14107 248388 14141 248404
rect 14221 249180 14255 249196
rect 14221 248388 14255 248404
rect 14317 249180 14351 249196
rect 14317 248388 14351 248404
rect 14431 249180 14465 249196
rect 14431 248388 14465 248404
rect 14527 249180 14561 249196
rect 14527 248388 14561 248404
rect 14641 249180 14675 249196
rect 14641 248388 14675 248404
rect 14737 249180 14771 249196
rect 14737 248388 14771 248404
rect 14851 249180 14885 249196
rect 14851 248388 14885 248404
rect 14947 249180 14981 249196
rect 14947 248388 14981 248404
rect 15061 249180 15095 249196
rect 15061 248388 15095 248404
rect 15157 249180 15191 249196
rect 15157 248388 15191 248404
rect 15271 249180 15305 249196
rect 15271 248388 15305 248404
rect 15367 249180 15401 249196
rect 15367 248388 15401 248404
rect 15481 249180 15515 249196
rect 15481 248388 15515 248404
rect 15577 249180 15611 249196
rect 15577 248388 15611 248404
rect 15691 249180 15725 249196
rect 15691 248388 15725 248404
rect 15787 249180 15821 249196
rect 15787 248388 15821 248404
rect 15901 249180 15935 249196
rect 15901 248388 15935 248404
rect 15997 249180 16031 249196
rect 15997 248388 16031 248404
rect 16111 249180 16145 249196
rect 16111 248388 16145 248404
rect 16207 249180 16241 249196
rect 16207 248388 16241 248404
rect 16321 249180 16355 249196
rect 16321 248388 16355 248404
rect 16417 249180 16451 249196
rect 16417 248388 16451 248404
rect 16531 249180 16565 249196
rect 16531 248388 16565 248404
rect 16627 249180 16661 249196
rect 16627 248388 16661 248404
rect 16741 249180 16775 249196
rect 16741 248388 16775 248404
rect 16837 249180 16871 249196
rect 16837 248388 16871 248404
rect 16951 249180 16985 249196
rect 16951 248388 16985 248404
rect 17047 249180 17081 249196
rect 17047 248388 17081 248404
rect 17161 249180 17195 249196
rect 17161 248388 17195 248404
rect 17257 249180 17291 249196
rect 17257 248388 17291 248404
rect 17371 249180 17405 249196
rect 17371 248388 17405 248404
rect 17467 249180 17501 249196
rect 17467 248388 17501 248404
rect 17581 249180 17615 249196
rect 17581 248388 17615 248404
rect 17677 249180 17711 249196
rect 17677 248388 17711 248404
rect 17791 249180 17825 249196
rect 17791 248388 17825 248404
rect 17887 249180 17921 249196
rect 17887 248388 17921 248404
rect 18001 249180 18035 249196
rect 18001 248388 18035 248404
rect 18097 249180 18131 249196
rect 18097 248388 18131 248404
rect 18211 249180 18245 249196
rect 18211 248388 18245 248404
rect 18307 249180 18341 249196
rect 18307 248388 18341 248404
rect 18421 249180 18455 249196
rect 18421 248388 18455 248404
rect 18517 249180 18551 249196
rect 18517 248388 18551 248404
rect 18631 249180 18665 249196
rect 18631 248388 18665 248404
rect 18727 249180 18761 249196
rect 18727 248388 18761 248404
rect 18841 249180 18875 249196
rect 18841 248388 18875 248404
rect 18937 249180 18971 249196
rect 18937 248388 18971 248404
rect 19051 249180 19085 249196
rect 19051 248388 19085 248404
rect 19147 249180 19181 249196
rect 19147 248388 19181 248404
rect 19261 249180 19295 249196
rect 19261 248388 19295 248404
rect 19357 249180 19391 249196
rect 19357 248388 19391 248404
rect 19471 249180 19505 249196
rect 19471 248388 19505 248404
rect 19567 249180 19601 249196
rect 19567 248388 19601 248404
rect 19681 249180 19715 249196
rect 19681 248388 19715 248404
rect 19777 249180 19811 249196
rect 19777 248388 19811 248404
rect 19891 249180 19925 249196
rect 19891 248388 19925 248404
rect 19987 249180 20021 249196
rect 19987 248388 20021 248404
rect 20101 249180 20135 249196
rect 20101 248388 20135 248404
rect 20197 249180 20231 249196
rect 20197 248388 20231 248404
rect 20311 249180 20345 249196
rect 20311 248388 20345 248404
rect 20407 249180 20441 249196
rect 20407 248388 20441 248404
rect 20521 249180 20555 249196
rect 20521 248388 20555 248404
rect 20617 249180 20651 249196
rect 20617 248388 20651 248404
rect 20731 249180 20765 249196
rect 20731 248388 20765 248404
rect 20827 249180 20861 249196
rect 20827 248388 20861 248404
rect 20941 249180 20975 249196
rect 20941 248388 20975 248404
rect 21037 249180 21071 249196
rect 21037 248388 21071 248404
rect 21151 249180 21185 249196
rect 21151 248388 21185 248404
rect 21247 249180 21281 249196
rect 21247 248388 21281 248404
rect 21361 249180 21395 249196
rect 21361 248388 21395 248404
rect 21457 249180 21491 249196
rect 21457 248388 21491 248404
rect 21571 249180 21605 249196
rect 21571 248388 21605 248404
rect 21667 249180 21701 249196
rect 21667 248388 21701 248404
rect 21781 249180 21815 249196
rect 21781 248388 21815 248404
rect 21877 249180 21911 249196
rect 21877 248388 21911 248404
rect 21991 249180 22025 249196
rect 21991 248388 22025 248404
rect 22087 249180 22121 249196
rect 22087 248388 22121 248404
rect 22201 249180 22235 249196
rect 22201 248388 22235 248404
rect 22297 249180 22331 249196
rect 22297 248388 22331 248404
rect 22411 249180 22445 249196
rect 22411 248388 22445 248404
rect 22507 249180 22541 249196
rect 22507 248388 22541 248404
rect 22621 249180 22655 249196
rect 22621 248388 22655 248404
rect 22717 249180 22751 249196
rect 22717 248388 22751 248404
rect 22831 249180 22865 249196
rect 22831 248388 22865 248404
rect 22927 249180 22961 249196
rect 22927 248388 22961 248404
rect 23041 249180 23075 249196
rect 23041 248388 23075 248404
rect 23137 249180 23171 249196
rect 23137 248388 23171 248404
rect 23251 249180 23285 249196
rect 23251 248388 23285 248404
rect 23347 249180 23381 249196
rect 23347 248388 23381 248404
rect 23461 249180 23495 249196
rect 23461 248388 23495 248404
rect 23557 249180 23591 249196
rect 23557 248388 23591 248404
rect 23671 249180 23705 249196
rect 23671 248388 23705 248404
rect 23767 249180 23801 249196
rect 23767 248388 23801 248404
rect 23881 249180 23915 249196
rect 23881 248388 23915 248404
rect 23977 249180 24011 249196
rect 23977 248388 24011 248404
rect 24091 249180 24125 249196
rect 24091 248388 24125 248404
rect 24187 249180 24221 249196
rect 24187 248388 24221 248404
rect 24301 249180 24335 249196
rect 24301 248388 24335 248404
rect 24397 249180 24431 249196
rect 24397 248388 24431 248404
rect 24511 249180 24545 249196
rect 24511 248388 24545 248404
rect 24607 249180 24641 249196
rect 24607 248388 24641 248404
rect 24721 249180 24755 249196
rect 24721 248388 24755 248404
rect 24817 249180 24851 249196
rect 24817 248388 24851 248404
rect 24931 249180 24965 249196
rect 24931 248388 24965 248404
rect 25027 249180 25061 249196
rect 25027 248388 25061 248404
rect 25141 249180 25175 249196
rect 25141 248388 25175 248404
rect 25237 249180 25271 249196
rect 25237 248388 25271 248404
rect 25351 249180 25385 249196
rect 25351 248388 25385 248404
rect 25447 249180 25481 249196
rect 25447 248388 25481 248404
rect 25561 249180 25595 249196
rect 25561 248388 25595 248404
rect 25657 249180 25691 249196
rect 25657 248388 25691 248404
rect 25771 249180 25805 249196
rect 25771 248388 25805 248404
rect 25867 249180 25901 249196
rect 25867 248388 25901 248404
rect 25981 249180 26015 249196
rect 25981 248388 26015 248404
rect 26077 249180 26111 249196
rect 26077 248388 26111 248404
rect 26191 249180 26225 249196
rect 26191 248388 26225 248404
rect 26287 249180 26321 249196
rect 26287 248388 26321 248404
rect 26401 249180 26435 249196
rect 26401 248388 26435 248404
rect 26497 249180 26531 249196
rect 26497 248388 26531 248404
rect 26611 249180 26645 249196
rect 26611 248388 26645 248404
rect 26707 249180 26741 249196
rect 26707 248388 26741 248404
rect 26821 249180 26855 249196
rect 26821 248388 26855 248404
rect 26917 249180 26951 249196
rect 26917 248388 26951 248404
rect 27031 249180 27065 249196
rect 27031 248388 27065 248404
rect 27127 249180 27161 249196
rect 27127 248388 27161 248404
rect 27241 249180 27275 249196
rect 27241 248388 27275 248404
rect 27337 249180 27371 249196
rect 27337 248388 27371 248404
rect -3807 248311 -3791 248345
rect -3807 248203 -3791 248237
rect -3757 248311 -3741 248345
rect -3387 248311 -3371 248345
rect -3757 248203 -3741 248237
rect -3387 248203 -3371 248237
rect -3337 248311 -3321 248345
rect -2967 248311 -2951 248345
rect -3337 248203 -3321 248237
rect -2967 248203 -2951 248237
rect -2917 248311 -2901 248345
rect -2547 248311 -2531 248345
rect -2917 248203 -2901 248237
rect -2547 248203 -2531 248237
rect -2497 248311 -2481 248345
rect -2127 248311 -2111 248345
rect -2497 248203 -2481 248237
rect -2127 248203 -2111 248237
rect -2077 248311 -2061 248345
rect -1707 248311 -1691 248345
rect -2077 248203 -2061 248237
rect -1707 248203 -1691 248237
rect -1657 248311 -1641 248345
rect -1287 248311 -1271 248345
rect -1657 248203 -1641 248237
rect -1287 248203 -1271 248237
rect -1237 248311 -1221 248345
rect -867 248311 -851 248345
rect -1237 248203 -1221 248237
rect -867 248203 -851 248237
rect -817 248311 -801 248345
rect -447 248311 -431 248345
rect -817 248203 -801 248237
rect -447 248203 -431 248237
rect -397 248311 -381 248345
rect -27 248311 -11 248345
rect -397 248203 -381 248237
rect -27 248203 -11 248237
rect 23 248311 39 248345
rect 393 248311 409 248345
rect 23 248203 39 248237
rect 393 248203 409 248237
rect 443 248311 459 248345
rect 813 248311 829 248345
rect 443 248203 459 248237
rect 813 248203 829 248237
rect 863 248311 879 248345
rect 1233 248311 1249 248345
rect 863 248203 879 248237
rect 1233 248203 1249 248237
rect 1283 248311 1299 248345
rect 1653 248311 1669 248345
rect 1283 248203 1299 248237
rect 1653 248203 1669 248237
rect 1703 248311 1719 248345
rect 2073 248311 2089 248345
rect 1703 248203 1719 248237
rect 2073 248203 2089 248237
rect 2123 248311 2139 248345
rect 2493 248311 2509 248345
rect 2123 248203 2139 248237
rect 2493 248203 2509 248237
rect 2543 248311 2559 248345
rect 2913 248311 2929 248345
rect 2543 248203 2559 248237
rect 2913 248203 2929 248237
rect 2963 248311 2979 248345
rect 3333 248311 3349 248345
rect 2963 248203 2979 248237
rect 3333 248203 3349 248237
rect 3383 248311 3399 248345
rect 3753 248311 3769 248345
rect 3383 248203 3399 248237
rect 3753 248203 3769 248237
rect 3803 248311 3819 248345
rect 4173 248311 4189 248345
rect 3803 248203 3819 248237
rect 4173 248203 4189 248237
rect 4223 248311 4239 248345
rect 4593 248311 4609 248345
rect 4223 248203 4239 248237
rect 4593 248203 4609 248237
rect 4643 248311 4659 248345
rect 5013 248311 5029 248345
rect 4643 248203 4659 248237
rect 5013 248203 5029 248237
rect 5063 248311 5079 248345
rect 5433 248311 5449 248345
rect 5063 248203 5079 248237
rect 5433 248203 5449 248237
rect 5483 248311 5499 248345
rect 5853 248311 5869 248345
rect 5483 248203 5499 248237
rect 5853 248203 5869 248237
rect 5903 248311 5919 248345
rect 6273 248311 6289 248345
rect 5903 248203 5919 248237
rect 6273 248203 6289 248237
rect 6323 248311 6339 248345
rect 6693 248311 6709 248345
rect 6323 248203 6339 248237
rect 6693 248203 6709 248237
rect 6743 248311 6759 248345
rect 7113 248311 7129 248345
rect 6743 248203 6759 248237
rect 7113 248203 7129 248237
rect 7163 248311 7179 248345
rect 7533 248311 7549 248345
rect 7163 248203 7179 248237
rect 7533 248203 7549 248237
rect 7583 248311 7599 248345
rect 7953 248311 7969 248345
rect 7583 248203 7599 248237
rect 7953 248203 7969 248237
rect 8003 248311 8019 248345
rect 8373 248311 8389 248345
rect 8003 248203 8019 248237
rect 8373 248203 8389 248237
rect 8423 248311 8439 248345
rect 8793 248311 8809 248345
rect 8423 248203 8439 248237
rect 8793 248203 8809 248237
rect 8843 248311 8859 248345
rect 9213 248311 9229 248345
rect 8843 248203 8859 248237
rect 9213 248203 9229 248237
rect 9263 248311 9279 248345
rect 9633 248311 9649 248345
rect 9263 248203 9279 248237
rect 9633 248203 9649 248237
rect 9683 248311 9699 248345
rect 10053 248311 10069 248345
rect 9683 248203 9699 248237
rect 10053 248203 10069 248237
rect 10103 248311 10119 248345
rect 10473 248311 10489 248345
rect 10103 248203 10119 248237
rect 10473 248203 10489 248237
rect 10523 248311 10539 248345
rect 10893 248311 10909 248345
rect 10523 248203 10539 248237
rect 10893 248203 10909 248237
rect 10943 248311 10959 248345
rect 11313 248311 11329 248345
rect 10943 248203 10959 248237
rect 11313 248203 11329 248237
rect 11363 248311 11379 248345
rect 11733 248311 11749 248345
rect 11363 248203 11379 248237
rect 11733 248203 11749 248237
rect 11783 248311 11799 248345
rect 12153 248311 12169 248345
rect 11783 248203 11799 248237
rect 12153 248203 12169 248237
rect 12203 248311 12219 248345
rect 12573 248311 12589 248345
rect 12203 248203 12219 248237
rect 12573 248203 12589 248237
rect 12623 248311 12639 248345
rect 12993 248311 13009 248345
rect 12623 248203 12639 248237
rect 12993 248203 13009 248237
rect 13043 248311 13059 248345
rect 13413 248311 13429 248345
rect 13043 248203 13059 248237
rect 13413 248203 13429 248237
rect 13463 248311 13479 248345
rect 13833 248311 13849 248345
rect 13463 248203 13479 248237
rect 13833 248203 13849 248237
rect 13883 248311 13899 248345
rect 14253 248311 14269 248345
rect 13883 248203 13899 248237
rect 14253 248203 14269 248237
rect 14303 248311 14319 248345
rect 14673 248311 14689 248345
rect 14303 248203 14319 248237
rect 14673 248203 14689 248237
rect 14723 248311 14739 248345
rect 15093 248311 15109 248345
rect 14723 248203 14739 248237
rect 15093 248203 15109 248237
rect 15143 248311 15159 248345
rect 15513 248311 15529 248345
rect 15143 248203 15159 248237
rect 15513 248203 15529 248237
rect 15563 248311 15579 248345
rect 15933 248311 15949 248345
rect 15563 248203 15579 248237
rect 15933 248203 15949 248237
rect 15983 248311 15999 248345
rect 16353 248311 16369 248345
rect 15983 248203 15999 248237
rect 16353 248203 16369 248237
rect 16403 248311 16419 248345
rect 16773 248311 16789 248345
rect 16403 248203 16419 248237
rect 16773 248203 16789 248237
rect 16823 248311 16839 248345
rect 17193 248311 17209 248345
rect 16823 248203 16839 248237
rect 17193 248203 17209 248237
rect 17243 248311 17259 248345
rect 17613 248311 17629 248345
rect 17243 248203 17259 248237
rect 17613 248203 17629 248237
rect 17663 248311 17679 248345
rect 18033 248311 18049 248345
rect 17663 248203 17679 248237
rect 18033 248203 18049 248237
rect 18083 248311 18099 248345
rect 18453 248311 18469 248345
rect 18083 248203 18099 248237
rect 18453 248203 18469 248237
rect 18503 248311 18519 248345
rect 18873 248311 18889 248345
rect 18503 248203 18519 248237
rect 18873 248203 18889 248237
rect 18923 248311 18939 248345
rect 19293 248311 19309 248345
rect 18923 248203 18939 248237
rect 19293 248203 19309 248237
rect 19343 248311 19359 248345
rect 19713 248311 19729 248345
rect 19343 248203 19359 248237
rect 19713 248203 19729 248237
rect 19763 248311 19779 248345
rect 20133 248311 20149 248345
rect 19763 248203 19779 248237
rect 20133 248203 20149 248237
rect 20183 248311 20199 248345
rect 20553 248311 20569 248345
rect 20183 248203 20199 248237
rect 20553 248203 20569 248237
rect 20603 248311 20619 248345
rect 20973 248311 20989 248345
rect 20603 248203 20619 248237
rect 20973 248203 20989 248237
rect 21023 248311 21039 248345
rect 21393 248311 21409 248345
rect 21023 248203 21039 248237
rect 21393 248203 21409 248237
rect 21443 248311 21459 248345
rect 21813 248311 21829 248345
rect 21443 248203 21459 248237
rect 21813 248203 21829 248237
rect 21863 248311 21879 248345
rect 22233 248311 22249 248345
rect 21863 248203 21879 248237
rect 22233 248203 22249 248237
rect 22283 248311 22299 248345
rect 22653 248311 22669 248345
rect 22283 248203 22299 248237
rect 22653 248203 22669 248237
rect 22703 248311 22719 248345
rect 23073 248311 23089 248345
rect 22703 248203 22719 248237
rect 23073 248203 23089 248237
rect 23123 248311 23139 248345
rect 23493 248311 23509 248345
rect 23123 248203 23139 248237
rect 23493 248203 23509 248237
rect 23543 248311 23559 248345
rect 23913 248311 23929 248345
rect 23543 248203 23559 248237
rect 23913 248203 23929 248237
rect 23963 248311 23979 248345
rect 24333 248311 24349 248345
rect 23963 248203 23979 248237
rect 24333 248203 24349 248237
rect 24383 248311 24399 248345
rect 24753 248311 24769 248345
rect 24383 248203 24399 248237
rect 24753 248203 24769 248237
rect 24803 248311 24819 248345
rect 25173 248311 25189 248345
rect 24803 248203 24819 248237
rect 25173 248203 25189 248237
rect 25223 248311 25239 248345
rect 25593 248311 25609 248345
rect 25223 248203 25239 248237
rect 25593 248203 25609 248237
rect 25643 248311 25659 248345
rect 26013 248311 26029 248345
rect 25643 248203 25659 248237
rect 26013 248203 26029 248237
rect 26063 248311 26079 248345
rect 26433 248311 26449 248345
rect 26063 248203 26079 248237
rect 26433 248203 26449 248237
rect 26483 248311 26499 248345
rect 26853 248311 26869 248345
rect 26483 248203 26499 248237
rect 26853 248203 26869 248237
rect 26903 248311 26919 248345
rect 27273 248311 27289 248345
rect 26903 248203 26919 248237
rect 27273 248203 27289 248237
rect 27323 248311 27339 248345
rect 27323 248203 27339 248237
rect -4049 248144 -4015 248160
rect -4049 247352 -4015 247368
rect -3953 248144 -3919 248160
rect -3953 247352 -3919 247368
rect -3839 248144 -3805 248160
rect -3839 247352 -3805 247368
rect -3743 248144 -3709 248160
rect -3743 247352 -3709 247368
rect -3629 248144 -3595 248160
rect -3629 247352 -3595 247368
rect -3533 248144 -3499 248160
rect -3533 247352 -3499 247368
rect -3419 248144 -3385 248160
rect -3419 247352 -3385 247368
rect -3323 248144 -3289 248160
rect -3323 247352 -3289 247368
rect -3209 248144 -3175 248160
rect -3209 247352 -3175 247368
rect -3113 248144 -3079 248160
rect -3113 247352 -3079 247368
rect -2999 248144 -2965 248160
rect -2999 247352 -2965 247368
rect -2903 248144 -2869 248160
rect -2903 247352 -2869 247368
rect -2789 248144 -2755 248160
rect -2789 247352 -2755 247368
rect -2693 248144 -2659 248160
rect -2693 247352 -2659 247368
rect -2579 248144 -2545 248160
rect -2579 247352 -2545 247368
rect -2483 248144 -2449 248160
rect -2483 247352 -2449 247368
rect -2369 248144 -2335 248160
rect -2369 247352 -2335 247368
rect -2273 248144 -2239 248160
rect -2273 247352 -2239 247368
rect -2159 248144 -2125 248160
rect -2159 247352 -2125 247368
rect -2063 248144 -2029 248160
rect -2063 247352 -2029 247368
rect -1949 248144 -1915 248160
rect -1949 247352 -1915 247368
rect -1853 248144 -1819 248160
rect -1853 247352 -1819 247368
rect -1739 248144 -1705 248160
rect -1739 247352 -1705 247368
rect -1643 248144 -1609 248160
rect -1643 247352 -1609 247368
rect -1529 248144 -1495 248160
rect -1529 247352 -1495 247368
rect -1433 248144 -1399 248160
rect -1433 247352 -1399 247368
rect -1319 248144 -1285 248160
rect -1319 247352 -1285 247368
rect -1223 248144 -1189 248160
rect -1223 247352 -1189 247368
rect -1109 248144 -1075 248160
rect -1109 247352 -1075 247368
rect -1013 248144 -979 248160
rect -1013 247352 -979 247368
rect -899 248144 -865 248160
rect -899 247352 -865 247368
rect -803 248144 -769 248160
rect -803 247352 -769 247368
rect -689 248144 -655 248160
rect -689 247352 -655 247368
rect -593 248144 -559 248160
rect -593 247352 -559 247368
rect -479 248144 -445 248160
rect -479 247352 -445 247368
rect -383 248144 -349 248160
rect -383 247352 -349 247368
rect -269 248144 -235 248160
rect -269 247352 -235 247368
rect -173 248144 -139 248160
rect -173 247352 -139 247368
rect -59 248144 -25 248160
rect -59 247352 -25 247368
rect 37 248144 71 248160
rect 37 247352 71 247368
rect 151 248144 185 248160
rect 151 247352 185 247368
rect 247 248144 281 248160
rect 247 247352 281 247368
rect 361 248144 395 248160
rect 361 247352 395 247368
rect 457 248144 491 248160
rect 457 247352 491 247368
rect 571 248144 605 248160
rect 571 247352 605 247368
rect 667 248144 701 248160
rect 667 247352 701 247368
rect 781 248144 815 248160
rect 781 247352 815 247368
rect 877 248144 911 248160
rect 877 247352 911 247368
rect 991 248144 1025 248160
rect 991 247352 1025 247368
rect 1087 248144 1121 248160
rect 1087 247352 1121 247368
rect 1201 248144 1235 248160
rect 1201 247352 1235 247368
rect 1297 248144 1331 248160
rect 1297 247352 1331 247368
rect 1411 248144 1445 248160
rect 1411 247352 1445 247368
rect 1507 248144 1541 248160
rect 1507 247352 1541 247368
rect 1621 248144 1655 248160
rect 1621 247352 1655 247368
rect 1717 248144 1751 248160
rect 1717 247352 1751 247368
rect 1831 248144 1865 248160
rect 1831 247352 1865 247368
rect 1927 248144 1961 248160
rect 1927 247352 1961 247368
rect 2041 248144 2075 248160
rect 2041 247352 2075 247368
rect 2137 248144 2171 248160
rect 2137 247352 2171 247368
rect 2251 248144 2285 248160
rect 2251 247352 2285 247368
rect 2347 248144 2381 248160
rect 2347 247352 2381 247368
rect 2461 248144 2495 248160
rect 2461 247352 2495 247368
rect 2557 248144 2591 248160
rect 2557 247352 2591 247368
rect 2671 248144 2705 248160
rect 2671 247352 2705 247368
rect 2767 248144 2801 248160
rect 2767 247352 2801 247368
rect 2881 248144 2915 248160
rect 2881 247352 2915 247368
rect 2977 248144 3011 248160
rect 2977 247352 3011 247368
rect 3091 248144 3125 248160
rect 3091 247352 3125 247368
rect 3187 248144 3221 248160
rect 3187 247352 3221 247368
rect 3301 248144 3335 248160
rect 3301 247352 3335 247368
rect 3397 248144 3431 248160
rect 3397 247352 3431 247368
rect 3511 248144 3545 248160
rect 3511 247352 3545 247368
rect 3607 248144 3641 248160
rect 3607 247352 3641 247368
rect 3721 248144 3755 248160
rect 3721 247352 3755 247368
rect 3817 248144 3851 248160
rect 3817 247352 3851 247368
rect 3931 248144 3965 248160
rect 3931 247352 3965 247368
rect 4027 248144 4061 248160
rect 4027 247352 4061 247368
rect 4141 248144 4175 248160
rect 4141 247352 4175 247368
rect 4237 248144 4271 248160
rect 4237 247352 4271 247368
rect 4351 248144 4385 248160
rect 4351 247352 4385 247368
rect 4447 248144 4481 248160
rect 4447 247352 4481 247368
rect 4561 248144 4595 248160
rect 4561 247352 4595 247368
rect 4657 248144 4691 248160
rect 4657 247352 4691 247368
rect 4771 248144 4805 248160
rect 4771 247352 4805 247368
rect 4867 248144 4901 248160
rect 4867 247352 4901 247368
rect 4981 248144 5015 248160
rect 4981 247352 5015 247368
rect 5077 248144 5111 248160
rect 5077 247352 5111 247368
rect 5191 248144 5225 248160
rect 5191 247352 5225 247368
rect 5287 248144 5321 248160
rect 5287 247352 5321 247368
rect 5401 248144 5435 248160
rect 5401 247352 5435 247368
rect 5497 248144 5531 248160
rect 5497 247352 5531 247368
rect 5611 248144 5645 248160
rect 5611 247352 5645 247368
rect 5707 248144 5741 248160
rect 5707 247352 5741 247368
rect 5821 248144 5855 248160
rect 5821 247352 5855 247368
rect 5917 248144 5951 248160
rect 5917 247352 5951 247368
rect 6031 248144 6065 248160
rect 6031 247352 6065 247368
rect 6127 248144 6161 248160
rect 6127 247352 6161 247368
rect 6241 248144 6275 248160
rect 6241 247352 6275 247368
rect 6337 248144 6371 248160
rect 6337 247352 6371 247368
rect 6451 248144 6485 248160
rect 6451 247352 6485 247368
rect 6547 248144 6581 248160
rect 6547 247352 6581 247368
rect 6661 248144 6695 248160
rect 6661 247352 6695 247368
rect 6757 248144 6791 248160
rect 6757 247352 6791 247368
rect 6871 248144 6905 248160
rect 6871 247352 6905 247368
rect 6967 248144 7001 248160
rect 6967 247352 7001 247368
rect 7081 248144 7115 248160
rect 7081 247352 7115 247368
rect 7177 248144 7211 248160
rect 7177 247352 7211 247368
rect 7291 248144 7325 248160
rect 7291 247352 7325 247368
rect 7387 248144 7421 248160
rect 7387 247352 7421 247368
rect 7501 248144 7535 248160
rect 7501 247352 7535 247368
rect 7597 248144 7631 248160
rect 7597 247352 7631 247368
rect 7711 248144 7745 248160
rect 7711 247352 7745 247368
rect 7807 248144 7841 248160
rect 7807 247352 7841 247368
rect 7921 248144 7955 248160
rect 7921 247352 7955 247368
rect 8017 248144 8051 248160
rect 8017 247352 8051 247368
rect 8131 248144 8165 248160
rect 8131 247352 8165 247368
rect 8227 248144 8261 248160
rect 8227 247352 8261 247368
rect 8341 248144 8375 248160
rect 8341 247352 8375 247368
rect 8437 248144 8471 248160
rect 8437 247352 8471 247368
rect 8551 248144 8585 248160
rect 8551 247352 8585 247368
rect 8647 248144 8681 248160
rect 8647 247352 8681 247368
rect 8761 248144 8795 248160
rect 8761 247352 8795 247368
rect 8857 248144 8891 248160
rect 8857 247352 8891 247368
rect 8971 248144 9005 248160
rect 8971 247352 9005 247368
rect 9067 248144 9101 248160
rect 9067 247352 9101 247368
rect 9181 248144 9215 248160
rect 9181 247352 9215 247368
rect 9277 248144 9311 248160
rect 9277 247352 9311 247368
rect 9391 248144 9425 248160
rect 9391 247352 9425 247368
rect 9487 248144 9521 248160
rect 9487 247352 9521 247368
rect 9601 248144 9635 248160
rect 9601 247352 9635 247368
rect 9697 248144 9731 248160
rect 9697 247352 9731 247368
rect 9811 248144 9845 248160
rect 9811 247352 9845 247368
rect 9907 248144 9941 248160
rect 9907 247352 9941 247368
rect 10021 248144 10055 248160
rect 10021 247352 10055 247368
rect 10117 248144 10151 248160
rect 10117 247352 10151 247368
rect 10231 248144 10265 248160
rect 10231 247352 10265 247368
rect 10327 248144 10361 248160
rect 10327 247352 10361 247368
rect 10441 248144 10475 248160
rect 10441 247352 10475 247368
rect 10537 248144 10571 248160
rect 10537 247352 10571 247368
rect 10651 248144 10685 248160
rect 10651 247352 10685 247368
rect 10747 248144 10781 248160
rect 10747 247352 10781 247368
rect 10861 248144 10895 248160
rect 10861 247352 10895 247368
rect 10957 248144 10991 248160
rect 10957 247352 10991 247368
rect 11071 248144 11105 248160
rect 11071 247352 11105 247368
rect 11167 248144 11201 248160
rect 11167 247352 11201 247368
rect 11281 248144 11315 248160
rect 11281 247352 11315 247368
rect 11377 248144 11411 248160
rect 11377 247352 11411 247368
rect 11491 248144 11525 248160
rect 11491 247352 11525 247368
rect 11587 248144 11621 248160
rect 11587 247352 11621 247368
rect 11701 248144 11735 248160
rect 11701 247352 11735 247368
rect 11797 248144 11831 248160
rect 11797 247352 11831 247368
rect 11911 248144 11945 248160
rect 11911 247352 11945 247368
rect 12007 248144 12041 248160
rect 12007 247352 12041 247368
rect 12121 248144 12155 248160
rect 12121 247352 12155 247368
rect 12217 248144 12251 248160
rect 12217 247352 12251 247368
rect 12331 248144 12365 248160
rect 12331 247352 12365 247368
rect 12427 248144 12461 248160
rect 12427 247352 12461 247368
rect 12541 248144 12575 248160
rect 12541 247352 12575 247368
rect 12637 248144 12671 248160
rect 12637 247352 12671 247368
rect 12751 248144 12785 248160
rect 12751 247352 12785 247368
rect 12847 248144 12881 248160
rect 12847 247352 12881 247368
rect 12961 248144 12995 248160
rect 12961 247352 12995 247368
rect 13057 248144 13091 248160
rect 13057 247352 13091 247368
rect 13171 248144 13205 248160
rect 13171 247352 13205 247368
rect 13267 248144 13301 248160
rect 13267 247352 13301 247368
rect 13381 248144 13415 248160
rect 13381 247352 13415 247368
rect 13477 248144 13511 248160
rect 13477 247352 13511 247368
rect 13591 248144 13625 248160
rect 13591 247352 13625 247368
rect 13687 248144 13721 248160
rect 13687 247352 13721 247368
rect 13801 248144 13835 248160
rect 13801 247352 13835 247368
rect 13897 248144 13931 248160
rect 13897 247352 13931 247368
rect 14011 248144 14045 248160
rect 14011 247352 14045 247368
rect 14107 248144 14141 248160
rect 14107 247352 14141 247368
rect 14221 248144 14255 248160
rect 14221 247352 14255 247368
rect 14317 248144 14351 248160
rect 14317 247352 14351 247368
rect 14431 248144 14465 248160
rect 14431 247352 14465 247368
rect 14527 248144 14561 248160
rect 14527 247352 14561 247368
rect 14641 248144 14675 248160
rect 14641 247352 14675 247368
rect 14737 248144 14771 248160
rect 14737 247352 14771 247368
rect 14851 248144 14885 248160
rect 14851 247352 14885 247368
rect 14947 248144 14981 248160
rect 14947 247352 14981 247368
rect 15061 248144 15095 248160
rect 15061 247352 15095 247368
rect 15157 248144 15191 248160
rect 15157 247352 15191 247368
rect 15271 248144 15305 248160
rect 15271 247352 15305 247368
rect 15367 248144 15401 248160
rect 15367 247352 15401 247368
rect 15481 248144 15515 248160
rect 15481 247352 15515 247368
rect 15577 248144 15611 248160
rect 15577 247352 15611 247368
rect 15691 248144 15725 248160
rect 15691 247352 15725 247368
rect 15787 248144 15821 248160
rect 15787 247352 15821 247368
rect 15901 248144 15935 248160
rect 15901 247352 15935 247368
rect 15997 248144 16031 248160
rect 15997 247352 16031 247368
rect 16111 248144 16145 248160
rect 16111 247352 16145 247368
rect 16207 248144 16241 248160
rect 16207 247352 16241 247368
rect 16321 248144 16355 248160
rect 16321 247352 16355 247368
rect 16417 248144 16451 248160
rect 16417 247352 16451 247368
rect 16531 248144 16565 248160
rect 16531 247352 16565 247368
rect 16627 248144 16661 248160
rect 16627 247352 16661 247368
rect 16741 248144 16775 248160
rect 16741 247352 16775 247368
rect 16837 248144 16871 248160
rect 16837 247352 16871 247368
rect 16951 248144 16985 248160
rect 16951 247352 16985 247368
rect 17047 248144 17081 248160
rect 17047 247352 17081 247368
rect 17161 248144 17195 248160
rect 17161 247352 17195 247368
rect 17257 248144 17291 248160
rect 17257 247352 17291 247368
rect 17371 248144 17405 248160
rect 17371 247352 17405 247368
rect 17467 248144 17501 248160
rect 17467 247352 17501 247368
rect 17581 248144 17615 248160
rect 17581 247352 17615 247368
rect 17677 248144 17711 248160
rect 17677 247352 17711 247368
rect 17791 248144 17825 248160
rect 17791 247352 17825 247368
rect 17887 248144 17921 248160
rect 17887 247352 17921 247368
rect 18001 248144 18035 248160
rect 18001 247352 18035 247368
rect 18097 248144 18131 248160
rect 18097 247352 18131 247368
rect 18211 248144 18245 248160
rect 18211 247352 18245 247368
rect 18307 248144 18341 248160
rect 18307 247352 18341 247368
rect 18421 248144 18455 248160
rect 18421 247352 18455 247368
rect 18517 248144 18551 248160
rect 18517 247352 18551 247368
rect 18631 248144 18665 248160
rect 18631 247352 18665 247368
rect 18727 248144 18761 248160
rect 18727 247352 18761 247368
rect 18841 248144 18875 248160
rect 18841 247352 18875 247368
rect 18937 248144 18971 248160
rect 18937 247352 18971 247368
rect 19051 248144 19085 248160
rect 19051 247352 19085 247368
rect 19147 248144 19181 248160
rect 19147 247352 19181 247368
rect 19261 248144 19295 248160
rect 19261 247352 19295 247368
rect 19357 248144 19391 248160
rect 19357 247352 19391 247368
rect 19471 248144 19505 248160
rect 19471 247352 19505 247368
rect 19567 248144 19601 248160
rect 19567 247352 19601 247368
rect 19681 248144 19715 248160
rect 19681 247352 19715 247368
rect 19777 248144 19811 248160
rect 19777 247352 19811 247368
rect 19891 248144 19925 248160
rect 19891 247352 19925 247368
rect 19987 248144 20021 248160
rect 19987 247352 20021 247368
rect 20101 248144 20135 248160
rect 20101 247352 20135 247368
rect 20197 248144 20231 248160
rect 20197 247352 20231 247368
rect 20311 248144 20345 248160
rect 20311 247352 20345 247368
rect 20407 248144 20441 248160
rect 20407 247352 20441 247368
rect 20521 248144 20555 248160
rect 20521 247352 20555 247368
rect 20617 248144 20651 248160
rect 20617 247352 20651 247368
rect 20731 248144 20765 248160
rect 20731 247352 20765 247368
rect 20827 248144 20861 248160
rect 20827 247352 20861 247368
rect 20941 248144 20975 248160
rect 20941 247352 20975 247368
rect 21037 248144 21071 248160
rect 21037 247352 21071 247368
rect 21151 248144 21185 248160
rect 21151 247352 21185 247368
rect 21247 248144 21281 248160
rect 21247 247352 21281 247368
rect 21361 248144 21395 248160
rect 21361 247352 21395 247368
rect 21457 248144 21491 248160
rect 21457 247352 21491 247368
rect 21571 248144 21605 248160
rect 21571 247352 21605 247368
rect 21667 248144 21701 248160
rect 21667 247352 21701 247368
rect 21781 248144 21815 248160
rect 21781 247352 21815 247368
rect 21877 248144 21911 248160
rect 21877 247352 21911 247368
rect 21991 248144 22025 248160
rect 21991 247352 22025 247368
rect 22087 248144 22121 248160
rect 22087 247352 22121 247368
rect 22201 248144 22235 248160
rect 22201 247352 22235 247368
rect 22297 248144 22331 248160
rect 22297 247352 22331 247368
rect 22411 248144 22445 248160
rect 22411 247352 22445 247368
rect 22507 248144 22541 248160
rect 22507 247352 22541 247368
rect 22621 248144 22655 248160
rect 22621 247352 22655 247368
rect 22717 248144 22751 248160
rect 22717 247352 22751 247368
rect 22831 248144 22865 248160
rect 22831 247352 22865 247368
rect 22927 248144 22961 248160
rect 22927 247352 22961 247368
rect 23041 248144 23075 248160
rect 23041 247352 23075 247368
rect 23137 248144 23171 248160
rect 23137 247352 23171 247368
rect 23251 248144 23285 248160
rect 23251 247352 23285 247368
rect 23347 248144 23381 248160
rect 23347 247352 23381 247368
rect 23461 248144 23495 248160
rect 23461 247352 23495 247368
rect 23557 248144 23591 248160
rect 23557 247352 23591 247368
rect 23671 248144 23705 248160
rect 23671 247352 23705 247368
rect 23767 248144 23801 248160
rect 23767 247352 23801 247368
rect 23881 248144 23915 248160
rect 23881 247352 23915 247368
rect 23977 248144 24011 248160
rect 23977 247352 24011 247368
rect 24091 248144 24125 248160
rect 24091 247352 24125 247368
rect 24187 248144 24221 248160
rect 24187 247352 24221 247368
rect 24301 248144 24335 248160
rect 24301 247352 24335 247368
rect 24397 248144 24431 248160
rect 24397 247352 24431 247368
rect 24511 248144 24545 248160
rect 24511 247352 24545 247368
rect 24607 248144 24641 248160
rect 24607 247352 24641 247368
rect 24721 248144 24755 248160
rect 24721 247352 24755 247368
rect 24817 248144 24851 248160
rect 24817 247352 24851 247368
rect 24931 248144 24965 248160
rect 24931 247352 24965 247368
rect 25027 248144 25061 248160
rect 25027 247352 25061 247368
rect 25141 248144 25175 248160
rect 25141 247352 25175 247368
rect 25237 248144 25271 248160
rect 25237 247352 25271 247368
rect 25351 248144 25385 248160
rect 25351 247352 25385 247368
rect 25447 248144 25481 248160
rect 25447 247352 25481 247368
rect 25561 248144 25595 248160
rect 25561 247352 25595 247368
rect 25657 248144 25691 248160
rect 25657 247352 25691 247368
rect 25771 248144 25805 248160
rect 25771 247352 25805 247368
rect 25867 248144 25901 248160
rect 25867 247352 25901 247368
rect 25981 248144 26015 248160
rect 25981 247352 26015 247368
rect 26077 248144 26111 248160
rect 26077 247352 26111 247368
rect 26191 248144 26225 248160
rect 26191 247352 26225 247368
rect 26287 248144 26321 248160
rect 26287 247352 26321 247368
rect 26401 248144 26435 248160
rect 26401 247352 26435 247368
rect 26497 248144 26531 248160
rect 26497 247352 26531 247368
rect 26611 248144 26645 248160
rect 26611 247352 26645 247368
rect 26707 248144 26741 248160
rect 26707 247352 26741 247368
rect 26821 248144 26855 248160
rect 26821 247352 26855 247368
rect 26917 248144 26951 248160
rect 26917 247352 26951 247368
rect 27031 248144 27065 248160
rect 27031 247352 27065 247368
rect 27127 248144 27161 248160
rect 27127 247352 27161 247368
rect 27241 248144 27275 248160
rect 27241 247352 27275 247368
rect 27337 248144 27371 248160
rect 27337 247352 27371 247368
rect -4017 247275 -4001 247309
rect -4017 247167 -4001 247201
rect -3967 247275 -3951 247309
rect -3597 247275 -3581 247309
rect -3967 247167 -3951 247201
rect -3597 247167 -3581 247201
rect -3547 247275 -3531 247309
rect -3177 247275 -3161 247309
rect -3547 247167 -3531 247201
rect -3177 247167 -3161 247201
rect -3127 247275 -3111 247309
rect -2757 247275 -2741 247309
rect -3127 247167 -3111 247201
rect -2757 247167 -2741 247201
rect -2707 247275 -2691 247309
rect -2337 247275 -2321 247309
rect -2707 247167 -2691 247201
rect -2337 247167 -2321 247201
rect -2287 247275 -2271 247309
rect -1917 247275 -1901 247309
rect -2287 247167 -2271 247201
rect -1917 247167 -1901 247201
rect -1867 247275 -1851 247309
rect -1497 247275 -1481 247309
rect -1867 247167 -1851 247201
rect -1497 247167 -1481 247201
rect -1447 247275 -1431 247309
rect -1077 247275 -1061 247309
rect -1447 247167 -1431 247201
rect -1077 247167 -1061 247201
rect -1027 247275 -1011 247309
rect -657 247275 -641 247309
rect -1027 247167 -1011 247201
rect -657 247167 -641 247201
rect -607 247275 -591 247309
rect -237 247275 -221 247309
rect -607 247167 -591 247201
rect -237 247167 -221 247201
rect -187 247275 -171 247309
rect 183 247275 199 247309
rect -187 247167 -171 247201
rect 183 247167 199 247201
rect 233 247275 249 247309
rect 603 247275 619 247309
rect 233 247167 249 247201
rect 603 247167 619 247201
rect 653 247275 669 247309
rect 1023 247275 1039 247309
rect 653 247167 669 247201
rect 1023 247167 1039 247201
rect 1073 247275 1089 247309
rect 1443 247275 1459 247309
rect 1073 247167 1089 247201
rect 1443 247167 1459 247201
rect 1493 247275 1509 247309
rect 1863 247275 1879 247309
rect 1493 247167 1509 247201
rect 1863 247167 1879 247201
rect 1913 247275 1929 247309
rect 2283 247275 2299 247309
rect 1913 247167 1929 247201
rect 2283 247167 2299 247201
rect 2333 247275 2349 247309
rect 2703 247275 2719 247309
rect 2333 247167 2349 247201
rect 2703 247167 2719 247201
rect 2753 247275 2769 247309
rect 3123 247275 3139 247309
rect 2753 247167 2769 247201
rect 3123 247167 3139 247201
rect 3173 247275 3189 247309
rect 3543 247275 3559 247309
rect 3173 247167 3189 247201
rect 3543 247167 3559 247201
rect 3593 247275 3609 247309
rect 3963 247275 3979 247309
rect 3593 247167 3609 247201
rect 3963 247167 3979 247201
rect 4013 247275 4029 247309
rect 4383 247275 4399 247309
rect 4013 247167 4029 247201
rect 4383 247167 4399 247201
rect 4433 247275 4449 247309
rect 4803 247275 4819 247309
rect 4433 247167 4449 247201
rect 4803 247167 4819 247201
rect 4853 247275 4869 247309
rect 5223 247275 5239 247309
rect 4853 247167 4869 247201
rect 5223 247167 5239 247201
rect 5273 247275 5289 247309
rect 5643 247275 5659 247309
rect 5273 247167 5289 247201
rect 5643 247167 5659 247201
rect 5693 247275 5709 247309
rect 6063 247275 6079 247309
rect 5693 247167 5709 247201
rect 6063 247167 6079 247201
rect 6113 247275 6129 247309
rect 6483 247275 6499 247309
rect 6113 247167 6129 247201
rect 6483 247167 6499 247201
rect 6533 247275 6549 247309
rect 6903 247275 6919 247309
rect 6533 247167 6549 247201
rect 6903 247167 6919 247201
rect 6953 247275 6969 247309
rect 7323 247275 7339 247309
rect 6953 247167 6969 247201
rect 7323 247167 7339 247201
rect 7373 247275 7389 247309
rect 7743 247275 7759 247309
rect 7373 247167 7389 247201
rect 7743 247167 7759 247201
rect 7793 247275 7809 247309
rect 8163 247275 8179 247309
rect 7793 247167 7809 247201
rect 8163 247167 8179 247201
rect 8213 247275 8229 247309
rect 8583 247275 8599 247309
rect 8213 247167 8229 247201
rect 8583 247167 8599 247201
rect 8633 247275 8649 247309
rect 9003 247275 9019 247309
rect 8633 247167 8649 247201
rect 9003 247167 9019 247201
rect 9053 247275 9069 247309
rect 9423 247275 9439 247309
rect 9053 247167 9069 247201
rect 9423 247167 9439 247201
rect 9473 247275 9489 247309
rect 9843 247275 9859 247309
rect 9473 247167 9489 247201
rect 9843 247167 9859 247201
rect 9893 247275 9909 247309
rect 10263 247275 10279 247309
rect 9893 247167 9909 247201
rect 10263 247167 10279 247201
rect 10313 247275 10329 247309
rect 10683 247275 10699 247309
rect 10313 247167 10329 247201
rect 10683 247167 10699 247201
rect 10733 247275 10749 247309
rect 11103 247275 11119 247309
rect 10733 247167 10749 247201
rect 11103 247167 11119 247201
rect 11153 247275 11169 247309
rect 11523 247275 11539 247309
rect 11153 247167 11169 247201
rect 11523 247167 11539 247201
rect 11573 247275 11589 247309
rect 11943 247275 11959 247309
rect 11573 247167 11589 247201
rect 11943 247167 11959 247201
rect 11993 247275 12009 247309
rect 12363 247275 12379 247309
rect 11993 247167 12009 247201
rect 12363 247167 12379 247201
rect 12413 247275 12429 247309
rect 12783 247275 12799 247309
rect 12413 247167 12429 247201
rect 12783 247167 12799 247201
rect 12833 247275 12849 247309
rect 13203 247275 13219 247309
rect 12833 247167 12849 247201
rect 13203 247167 13219 247201
rect 13253 247275 13269 247309
rect 13623 247275 13639 247309
rect 13253 247167 13269 247201
rect 13623 247167 13639 247201
rect 13673 247275 13689 247309
rect 14043 247275 14059 247309
rect 13673 247167 13689 247201
rect 14043 247167 14059 247201
rect 14093 247275 14109 247309
rect 14463 247275 14479 247309
rect 14093 247167 14109 247201
rect 14463 247167 14479 247201
rect 14513 247275 14529 247309
rect 14883 247275 14899 247309
rect 14513 247167 14529 247201
rect 14883 247167 14899 247201
rect 14933 247275 14949 247309
rect 15303 247275 15319 247309
rect 14933 247167 14949 247201
rect 15303 247167 15319 247201
rect 15353 247275 15369 247309
rect 15723 247275 15739 247309
rect 15353 247167 15369 247201
rect 15723 247167 15739 247201
rect 15773 247275 15789 247309
rect 16143 247275 16159 247309
rect 15773 247167 15789 247201
rect 16143 247167 16159 247201
rect 16193 247275 16209 247309
rect 16563 247275 16579 247309
rect 16193 247167 16209 247201
rect 16563 247167 16579 247201
rect 16613 247275 16629 247309
rect 16983 247275 16999 247309
rect 16613 247167 16629 247201
rect 16983 247167 16999 247201
rect 17033 247275 17049 247309
rect 17403 247275 17419 247309
rect 17033 247167 17049 247201
rect 17403 247167 17419 247201
rect 17453 247275 17469 247309
rect 17823 247275 17839 247309
rect 17453 247167 17469 247201
rect 17823 247167 17839 247201
rect 17873 247275 17889 247309
rect 18243 247275 18259 247309
rect 17873 247167 17889 247201
rect 18243 247167 18259 247201
rect 18293 247275 18309 247309
rect 18663 247275 18679 247309
rect 18293 247167 18309 247201
rect 18663 247167 18679 247201
rect 18713 247275 18729 247309
rect 19083 247275 19099 247309
rect 18713 247167 18729 247201
rect 19083 247167 19099 247201
rect 19133 247275 19149 247309
rect 19503 247275 19519 247309
rect 19133 247167 19149 247201
rect 19503 247167 19519 247201
rect 19553 247275 19569 247309
rect 19923 247275 19939 247309
rect 19553 247167 19569 247201
rect 19923 247167 19939 247201
rect 19973 247275 19989 247309
rect 20343 247275 20359 247309
rect 19973 247167 19989 247201
rect 20343 247167 20359 247201
rect 20393 247275 20409 247309
rect 20763 247275 20779 247309
rect 20393 247167 20409 247201
rect 20763 247167 20779 247201
rect 20813 247275 20829 247309
rect 21183 247275 21199 247309
rect 20813 247167 20829 247201
rect 21183 247167 21199 247201
rect 21233 247275 21249 247309
rect 21603 247275 21619 247309
rect 21233 247167 21249 247201
rect 21603 247167 21619 247201
rect 21653 247275 21669 247309
rect 22023 247275 22039 247309
rect 21653 247167 21669 247201
rect 22023 247167 22039 247201
rect 22073 247275 22089 247309
rect 22443 247275 22459 247309
rect 22073 247167 22089 247201
rect 22443 247167 22459 247201
rect 22493 247275 22509 247309
rect 22863 247275 22879 247309
rect 22493 247167 22509 247201
rect 22863 247167 22879 247201
rect 22913 247275 22929 247309
rect 23283 247275 23299 247309
rect 22913 247167 22929 247201
rect 23283 247167 23299 247201
rect 23333 247275 23349 247309
rect 23703 247275 23719 247309
rect 23333 247167 23349 247201
rect 23703 247167 23719 247201
rect 23753 247275 23769 247309
rect 24123 247275 24139 247309
rect 23753 247167 23769 247201
rect 24123 247167 24139 247201
rect 24173 247275 24189 247309
rect 24543 247275 24559 247309
rect 24173 247167 24189 247201
rect 24543 247167 24559 247201
rect 24593 247275 24609 247309
rect 24963 247275 24979 247309
rect 24593 247167 24609 247201
rect 24963 247167 24979 247201
rect 25013 247275 25029 247309
rect 25383 247275 25399 247309
rect 25013 247167 25029 247201
rect 25383 247167 25399 247201
rect 25433 247275 25449 247309
rect 25803 247275 25819 247309
rect 25433 247167 25449 247201
rect 25803 247167 25819 247201
rect 25853 247275 25869 247309
rect 26223 247275 26239 247309
rect 25853 247167 25869 247201
rect 26223 247167 26239 247201
rect 26273 247275 26289 247309
rect 26643 247275 26659 247309
rect 26273 247167 26289 247201
rect 26643 247167 26659 247201
rect 26693 247275 26709 247309
rect 27063 247275 27079 247309
rect 26693 247167 26709 247201
rect 27063 247167 27079 247201
rect 27113 247275 27129 247309
rect 27113 247167 27129 247201
rect -4049 247108 -4015 247124
rect -4049 246316 -4015 246332
rect -3953 247108 -3919 247124
rect -3953 246316 -3919 246332
rect -3839 247108 -3805 247124
rect -3839 246316 -3805 246332
rect -3743 247108 -3709 247124
rect -3743 246316 -3709 246332
rect -3629 247108 -3595 247124
rect -3629 246316 -3595 246332
rect -3533 247108 -3499 247124
rect -3533 246316 -3499 246332
rect -3419 247108 -3385 247124
rect -3419 246316 -3385 246332
rect -3323 247108 -3289 247124
rect -3323 246316 -3289 246332
rect -3209 247108 -3175 247124
rect -3209 246316 -3175 246332
rect -3113 247108 -3079 247124
rect -3113 246316 -3079 246332
rect -2999 247108 -2965 247124
rect -2999 246316 -2965 246332
rect -2903 247108 -2869 247124
rect -2903 246316 -2869 246332
rect -2789 247108 -2755 247124
rect -2789 246316 -2755 246332
rect -2693 247108 -2659 247124
rect -2693 246316 -2659 246332
rect -2579 247108 -2545 247124
rect -2579 246316 -2545 246332
rect -2483 247108 -2449 247124
rect -2483 246316 -2449 246332
rect -2369 247108 -2335 247124
rect -2369 246316 -2335 246332
rect -2273 247108 -2239 247124
rect -2273 246316 -2239 246332
rect -2159 247108 -2125 247124
rect -2159 246316 -2125 246332
rect -2063 247108 -2029 247124
rect -2063 246316 -2029 246332
rect -1949 247108 -1915 247124
rect -1949 246316 -1915 246332
rect -1853 247108 -1819 247124
rect -1853 246316 -1819 246332
rect -1739 247108 -1705 247124
rect -1739 246316 -1705 246332
rect -1643 247108 -1609 247124
rect -1643 246316 -1609 246332
rect -1529 247108 -1495 247124
rect -1529 246316 -1495 246332
rect -1433 247108 -1399 247124
rect -1433 246316 -1399 246332
rect -1319 247108 -1285 247124
rect -1319 246316 -1285 246332
rect -1223 247108 -1189 247124
rect -1223 246316 -1189 246332
rect -1109 247108 -1075 247124
rect -1109 246316 -1075 246332
rect -1013 247108 -979 247124
rect -1013 246316 -979 246332
rect -899 247108 -865 247124
rect -899 246316 -865 246332
rect -803 247108 -769 247124
rect -803 246316 -769 246332
rect -689 247108 -655 247124
rect -689 246316 -655 246332
rect -593 247108 -559 247124
rect -593 246316 -559 246332
rect -479 247108 -445 247124
rect -479 246316 -445 246332
rect -383 247108 -349 247124
rect -383 246316 -349 246332
rect -269 247108 -235 247124
rect -269 246316 -235 246332
rect -173 247108 -139 247124
rect -173 246316 -139 246332
rect -59 247108 -25 247124
rect -59 246316 -25 246332
rect 37 247108 71 247124
rect 37 246316 71 246332
rect 151 247108 185 247124
rect 151 246316 185 246332
rect 247 247108 281 247124
rect 247 246316 281 246332
rect 361 247108 395 247124
rect 361 246316 395 246332
rect 457 247108 491 247124
rect 457 246316 491 246332
rect 571 247108 605 247124
rect 571 246316 605 246332
rect 667 247108 701 247124
rect 667 246316 701 246332
rect 781 247108 815 247124
rect 781 246316 815 246332
rect 877 247108 911 247124
rect 877 246316 911 246332
rect 991 247108 1025 247124
rect 991 246316 1025 246332
rect 1087 247108 1121 247124
rect 1087 246316 1121 246332
rect 1201 247108 1235 247124
rect 1201 246316 1235 246332
rect 1297 247108 1331 247124
rect 1297 246316 1331 246332
rect 1411 247108 1445 247124
rect 1411 246316 1445 246332
rect 1507 247108 1541 247124
rect 1507 246316 1541 246332
rect 1621 247108 1655 247124
rect 1621 246316 1655 246332
rect 1717 247108 1751 247124
rect 1717 246316 1751 246332
rect 1831 247108 1865 247124
rect 1831 246316 1865 246332
rect 1927 247108 1961 247124
rect 1927 246316 1961 246332
rect 2041 247108 2075 247124
rect 2041 246316 2075 246332
rect 2137 247108 2171 247124
rect 2137 246316 2171 246332
rect 2251 247108 2285 247124
rect 2251 246316 2285 246332
rect 2347 247108 2381 247124
rect 2347 246316 2381 246332
rect 2461 247108 2495 247124
rect 2461 246316 2495 246332
rect 2557 247108 2591 247124
rect 2557 246316 2591 246332
rect 2671 247108 2705 247124
rect 2671 246316 2705 246332
rect 2767 247108 2801 247124
rect 2767 246316 2801 246332
rect 2881 247108 2915 247124
rect 2881 246316 2915 246332
rect 2977 247108 3011 247124
rect 2977 246316 3011 246332
rect 3091 247108 3125 247124
rect 3091 246316 3125 246332
rect 3187 247108 3221 247124
rect 3187 246316 3221 246332
rect 3301 247108 3335 247124
rect 3301 246316 3335 246332
rect 3397 247108 3431 247124
rect 3397 246316 3431 246332
rect 3511 247108 3545 247124
rect 3511 246316 3545 246332
rect 3607 247108 3641 247124
rect 3607 246316 3641 246332
rect 3721 247108 3755 247124
rect 3721 246316 3755 246332
rect 3817 247108 3851 247124
rect 3817 246316 3851 246332
rect 3931 247108 3965 247124
rect 3931 246316 3965 246332
rect 4027 247108 4061 247124
rect 4027 246316 4061 246332
rect 4141 247108 4175 247124
rect 4141 246316 4175 246332
rect 4237 247108 4271 247124
rect 4237 246316 4271 246332
rect 4351 247108 4385 247124
rect 4351 246316 4385 246332
rect 4447 247108 4481 247124
rect 4447 246316 4481 246332
rect 4561 247108 4595 247124
rect 4561 246316 4595 246332
rect 4657 247108 4691 247124
rect 4657 246316 4691 246332
rect 4771 247108 4805 247124
rect 4771 246316 4805 246332
rect 4867 247108 4901 247124
rect 4867 246316 4901 246332
rect 4981 247108 5015 247124
rect 4981 246316 5015 246332
rect 5077 247108 5111 247124
rect 5077 246316 5111 246332
rect 5191 247108 5225 247124
rect 5191 246316 5225 246332
rect 5287 247108 5321 247124
rect 5287 246316 5321 246332
rect 5401 247108 5435 247124
rect 5401 246316 5435 246332
rect 5497 247108 5531 247124
rect 5497 246316 5531 246332
rect 5611 247108 5645 247124
rect 5611 246316 5645 246332
rect 5707 247108 5741 247124
rect 5707 246316 5741 246332
rect 5821 247108 5855 247124
rect 5821 246316 5855 246332
rect 5917 247108 5951 247124
rect 5917 246316 5951 246332
rect 6031 247108 6065 247124
rect 6031 246316 6065 246332
rect 6127 247108 6161 247124
rect 6127 246316 6161 246332
rect 6241 247108 6275 247124
rect 6241 246316 6275 246332
rect 6337 247108 6371 247124
rect 6337 246316 6371 246332
rect 6451 247108 6485 247124
rect 6451 246316 6485 246332
rect 6547 247108 6581 247124
rect 6547 246316 6581 246332
rect 6661 247108 6695 247124
rect 6661 246316 6695 246332
rect 6757 247108 6791 247124
rect 6757 246316 6791 246332
rect 6871 247108 6905 247124
rect 6871 246316 6905 246332
rect 6967 247108 7001 247124
rect 6967 246316 7001 246332
rect 7081 247108 7115 247124
rect 7081 246316 7115 246332
rect 7177 247108 7211 247124
rect 7177 246316 7211 246332
rect 7291 247108 7325 247124
rect 7291 246316 7325 246332
rect 7387 247108 7421 247124
rect 7387 246316 7421 246332
rect 7501 247108 7535 247124
rect 7501 246316 7535 246332
rect 7597 247108 7631 247124
rect 7597 246316 7631 246332
rect 7711 247108 7745 247124
rect 7711 246316 7745 246332
rect 7807 247108 7841 247124
rect 7807 246316 7841 246332
rect 7921 247108 7955 247124
rect 7921 246316 7955 246332
rect 8017 247108 8051 247124
rect 8017 246316 8051 246332
rect 8131 247108 8165 247124
rect 8131 246316 8165 246332
rect 8227 247108 8261 247124
rect 8227 246316 8261 246332
rect 8341 247108 8375 247124
rect 8341 246316 8375 246332
rect 8437 247108 8471 247124
rect 8437 246316 8471 246332
rect 8551 247108 8585 247124
rect 8551 246316 8585 246332
rect 8647 247108 8681 247124
rect 8647 246316 8681 246332
rect 8761 247108 8795 247124
rect 8761 246316 8795 246332
rect 8857 247108 8891 247124
rect 8857 246316 8891 246332
rect 8971 247108 9005 247124
rect 8971 246316 9005 246332
rect 9067 247108 9101 247124
rect 9067 246316 9101 246332
rect 9181 247108 9215 247124
rect 9181 246316 9215 246332
rect 9277 247108 9311 247124
rect 9277 246316 9311 246332
rect 9391 247108 9425 247124
rect 9391 246316 9425 246332
rect 9487 247108 9521 247124
rect 9487 246316 9521 246332
rect 9601 247108 9635 247124
rect 9601 246316 9635 246332
rect 9697 247108 9731 247124
rect 9697 246316 9731 246332
rect 9811 247108 9845 247124
rect 9811 246316 9845 246332
rect 9907 247108 9941 247124
rect 9907 246316 9941 246332
rect 10021 247108 10055 247124
rect 10021 246316 10055 246332
rect 10117 247108 10151 247124
rect 10117 246316 10151 246332
rect 10231 247108 10265 247124
rect 10231 246316 10265 246332
rect 10327 247108 10361 247124
rect 10327 246316 10361 246332
rect 10441 247108 10475 247124
rect 10441 246316 10475 246332
rect 10537 247108 10571 247124
rect 10537 246316 10571 246332
rect 10651 247108 10685 247124
rect 10651 246316 10685 246332
rect 10747 247108 10781 247124
rect 10747 246316 10781 246332
rect 10861 247108 10895 247124
rect 10861 246316 10895 246332
rect 10957 247108 10991 247124
rect 10957 246316 10991 246332
rect 11071 247108 11105 247124
rect 11071 246316 11105 246332
rect 11167 247108 11201 247124
rect 11167 246316 11201 246332
rect 11281 247108 11315 247124
rect 11281 246316 11315 246332
rect 11377 247108 11411 247124
rect 11377 246316 11411 246332
rect 11491 247108 11525 247124
rect 11491 246316 11525 246332
rect 11587 247108 11621 247124
rect 11587 246316 11621 246332
rect 11701 247108 11735 247124
rect 11701 246316 11735 246332
rect 11797 247108 11831 247124
rect 11797 246316 11831 246332
rect 11911 247108 11945 247124
rect 11911 246316 11945 246332
rect 12007 247108 12041 247124
rect 12007 246316 12041 246332
rect 12121 247108 12155 247124
rect 12121 246316 12155 246332
rect 12217 247108 12251 247124
rect 12217 246316 12251 246332
rect 12331 247108 12365 247124
rect 12331 246316 12365 246332
rect 12427 247108 12461 247124
rect 12427 246316 12461 246332
rect 12541 247108 12575 247124
rect 12541 246316 12575 246332
rect 12637 247108 12671 247124
rect 12637 246316 12671 246332
rect 12751 247108 12785 247124
rect 12751 246316 12785 246332
rect 12847 247108 12881 247124
rect 12847 246316 12881 246332
rect 12961 247108 12995 247124
rect 12961 246316 12995 246332
rect 13057 247108 13091 247124
rect 13057 246316 13091 246332
rect 13171 247108 13205 247124
rect 13171 246316 13205 246332
rect 13267 247108 13301 247124
rect 13267 246316 13301 246332
rect 13381 247108 13415 247124
rect 13381 246316 13415 246332
rect 13477 247108 13511 247124
rect 13477 246316 13511 246332
rect 13591 247108 13625 247124
rect 13591 246316 13625 246332
rect 13687 247108 13721 247124
rect 13687 246316 13721 246332
rect 13801 247108 13835 247124
rect 13801 246316 13835 246332
rect 13897 247108 13931 247124
rect 13897 246316 13931 246332
rect 14011 247108 14045 247124
rect 14011 246316 14045 246332
rect 14107 247108 14141 247124
rect 14107 246316 14141 246332
rect 14221 247108 14255 247124
rect 14221 246316 14255 246332
rect 14317 247108 14351 247124
rect 14317 246316 14351 246332
rect 14431 247108 14465 247124
rect 14431 246316 14465 246332
rect 14527 247108 14561 247124
rect 14527 246316 14561 246332
rect 14641 247108 14675 247124
rect 14641 246316 14675 246332
rect 14737 247108 14771 247124
rect 14737 246316 14771 246332
rect 14851 247108 14885 247124
rect 14851 246316 14885 246332
rect 14947 247108 14981 247124
rect 14947 246316 14981 246332
rect 15061 247108 15095 247124
rect 15061 246316 15095 246332
rect 15157 247108 15191 247124
rect 15157 246316 15191 246332
rect 15271 247108 15305 247124
rect 15271 246316 15305 246332
rect 15367 247108 15401 247124
rect 15367 246316 15401 246332
rect 15481 247108 15515 247124
rect 15481 246316 15515 246332
rect 15577 247108 15611 247124
rect 15577 246316 15611 246332
rect 15691 247108 15725 247124
rect 15691 246316 15725 246332
rect 15787 247108 15821 247124
rect 15787 246316 15821 246332
rect 15901 247108 15935 247124
rect 15901 246316 15935 246332
rect 15997 247108 16031 247124
rect 15997 246316 16031 246332
rect 16111 247108 16145 247124
rect 16111 246316 16145 246332
rect 16207 247108 16241 247124
rect 16207 246316 16241 246332
rect 16321 247108 16355 247124
rect 16321 246316 16355 246332
rect 16417 247108 16451 247124
rect 16417 246316 16451 246332
rect 16531 247108 16565 247124
rect 16531 246316 16565 246332
rect 16627 247108 16661 247124
rect 16627 246316 16661 246332
rect 16741 247108 16775 247124
rect 16741 246316 16775 246332
rect 16837 247108 16871 247124
rect 16837 246316 16871 246332
rect 16951 247108 16985 247124
rect 16951 246316 16985 246332
rect 17047 247108 17081 247124
rect 17047 246316 17081 246332
rect 17161 247108 17195 247124
rect 17161 246316 17195 246332
rect 17257 247108 17291 247124
rect 17257 246316 17291 246332
rect 17371 247108 17405 247124
rect 17371 246316 17405 246332
rect 17467 247108 17501 247124
rect 17467 246316 17501 246332
rect 17581 247108 17615 247124
rect 17581 246316 17615 246332
rect 17677 247108 17711 247124
rect 17677 246316 17711 246332
rect 17791 247108 17825 247124
rect 17791 246316 17825 246332
rect 17887 247108 17921 247124
rect 17887 246316 17921 246332
rect 18001 247108 18035 247124
rect 18001 246316 18035 246332
rect 18097 247108 18131 247124
rect 18097 246316 18131 246332
rect 18211 247108 18245 247124
rect 18211 246316 18245 246332
rect 18307 247108 18341 247124
rect 18307 246316 18341 246332
rect 18421 247108 18455 247124
rect 18421 246316 18455 246332
rect 18517 247108 18551 247124
rect 18517 246316 18551 246332
rect 18631 247108 18665 247124
rect 18631 246316 18665 246332
rect 18727 247108 18761 247124
rect 18727 246316 18761 246332
rect 18841 247108 18875 247124
rect 18841 246316 18875 246332
rect 18937 247108 18971 247124
rect 18937 246316 18971 246332
rect 19051 247108 19085 247124
rect 19051 246316 19085 246332
rect 19147 247108 19181 247124
rect 19147 246316 19181 246332
rect 19261 247108 19295 247124
rect 19261 246316 19295 246332
rect 19357 247108 19391 247124
rect 19357 246316 19391 246332
rect 19471 247108 19505 247124
rect 19471 246316 19505 246332
rect 19567 247108 19601 247124
rect 19567 246316 19601 246332
rect 19681 247108 19715 247124
rect 19681 246316 19715 246332
rect 19777 247108 19811 247124
rect 19777 246316 19811 246332
rect 19891 247108 19925 247124
rect 19891 246316 19925 246332
rect 19987 247108 20021 247124
rect 19987 246316 20021 246332
rect 20101 247108 20135 247124
rect 20101 246316 20135 246332
rect 20197 247108 20231 247124
rect 20197 246316 20231 246332
rect 20311 247108 20345 247124
rect 20311 246316 20345 246332
rect 20407 247108 20441 247124
rect 20407 246316 20441 246332
rect 20521 247108 20555 247124
rect 20521 246316 20555 246332
rect 20617 247108 20651 247124
rect 20617 246316 20651 246332
rect 20731 247108 20765 247124
rect 20731 246316 20765 246332
rect 20827 247108 20861 247124
rect 20827 246316 20861 246332
rect 20941 247108 20975 247124
rect 20941 246316 20975 246332
rect 21037 247108 21071 247124
rect 21037 246316 21071 246332
rect 21151 247108 21185 247124
rect 21151 246316 21185 246332
rect 21247 247108 21281 247124
rect 21247 246316 21281 246332
rect 21361 247108 21395 247124
rect 21361 246316 21395 246332
rect 21457 247108 21491 247124
rect 21457 246316 21491 246332
rect 21571 247108 21605 247124
rect 21571 246316 21605 246332
rect 21667 247108 21701 247124
rect 21667 246316 21701 246332
rect 21781 247108 21815 247124
rect 21781 246316 21815 246332
rect 21877 247108 21911 247124
rect 21877 246316 21911 246332
rect 21991 247108 22025 247124
rect 21991 246316 22025 246332
rect 22087 247108 22121 247124
rect 22087 246316 22121 246332
rect 22201 247108 22235 247124
rect 22201 246316 22235 246332
rect 22297 247108 22331 247124
rect 22297 246316 22331 246332
rect 22411 247108 22445 247124
rect 22411 246316 22445 246332
rect 22507 247108 22541 247124
rect 22507 246316 22541 246332
rect 22621 247108 22655 247124
rect 22621 246316 22655 246332
rect 22717 247108 22751 247124
rect 22717 246316 22751 246332
rect 22831 247108 22865 247124
rect 22831 246316 22865 246332
rect 22927 247108 22961 247124
rect 22927 246316 22961 246332
rect 23041 247108 23075 247124
rect 23041 246316 23075 246332
rect 23137 247108 23171 247124
rect 23137 246316 23171 246332
rect 23251 247108 23285 247124
rect 23251 246316 23285 246332
rect 23347 247108 23381 247124
rect 23347 246316 23381 246332
rect 23461 247108 23495 247124
rect 23461 246316 23495 246332
rect 23557 247108 23591 247124
rect 23557 246316 23591 246332
rect 23671 247108 23705 247124
rect 23671 246316 23705 246332
rect 23767 247108 23801 247124
rect 23767 246316 23801 246332
rect 23881 247108 23915 247124
rect 23881 246316 23915 246332
rect 23977 247108 24011 247124
rect 23977 246316 24011 246332
rect 24091 247108 24125 247124
rect 24091 246316 24125 246332
rect 24187 247108 24221 247124
rect 24187 246316 24221 246332
rect 24301 247108 24335 247124
rect 24301 246316 24335 246332
rect 24397 247108 24431 247124
rect 24397 246316 24431 246332
rect 24511 247108 24545 247124
rect 24511 246316 24545 246332
rect 24607 247108 24641 247124
rect 24607 246316 24641 246332
rect 24721 247108 24755 247124
rect 24721 246316 24755 246332
rect 24817 247108 24851 247124
rect 24817 246316 24851 246332
rect 24931 247108 24965 247124
rect 24931 246316 24965 246332
rect 25027 247108 25061 247124
rect 25027 246316 25061 246332
rect 25141 247108 25175 247124
rect 25141 246316 25175 246332
rect 25237 247108 25271 247124
rect 25237 246316 25271 246332
rect 25351 247108 25385 247124
rect 25351 246316 25385 246332
rect 25447 247108 25481 247124
rect 25447 246316 25481 246332
rect 25561 247108 25595 247124
rect 25561 246316 25595 246332
rect 25657 247108 25691 247124
rect 25657 246316 25691 246332
rect 25771 247108 25805 247124
rect 25771 246316 25805 246332
rect 25867 247108 25901 247124
rect 25867 246316 25901 246332
rect 25981 247108 26015 247124
rect 25981 246316 26015 246332
rect 26077 247108 26111 247124
rect 26077 246316 26111 246332
rect 26191 247108 26225 247124
rect 26191 246316 26225 246332
rect 26287 247108 26321 247124
rect 26287 246316 26321 246332
rect 26401 247108 26435 247124
rect 26401 246316 26435 246332
rect 26497 247108 26531 247124
rect 26497 246316 26531 246332
rect 26611 247108 26645 247124
rect 26611 246316 26645 246332
rect 26707 247108 26741 247124
rect 26707 246316 26741 246332
rect 26821 247108 26855 247124
rect 26821 246316 26855 246332
rect 26917 247108 26951 247124
rect 26917 246316 26951 246332
rect 27031 247108 27065 247124
rect 27031 246316 27065 246332
rect 27127 247108 27161 247124
rect 27127 246316 27161 246332
rect 27241 247108 27275 247124
rect 27241 246316 27275 246332
rect 27337 247108 27371 247124
rect 27337 246316 27371 246332
rect -3807 246239 -3791 246273
rect -3807 246131 -3791 246165
rect -3757 246239 -3741 246273
rect -3387 246239 -3371 246273
rect -3757 246131 -3741 246165
rect -3387 246131 -3371 246165
rect -3337 246239 -3321 246273
rect -2967 246239 -2951 246273
rect -3337 246131 -3321 246165
rect -2967 246131 -2951 246165
rect -2917 246239 -2901 246273
rect -2547 246239 -2531 246273
rect -2917 246131 -2901 246165
rect -2547 246131 -2531 246165
rect -2497 246239 -2481 246273
rect -2127 246239 -2111 246273
rect -2497 246131 -2481 246165
rect -2127 246131 -2111 246165
rect -2077 246239 -2061 246273
rect -1707 246239 -1691 246273
rect -2077 246131 -2061 246165
rect -1707 246131 -1691 246165
rect -1657 246239 -1641 246273
rect -1287 246239 -1271 246273
rect -1657 246131 -1641 246165
rect -1287 246131 -1271 246165
rect -1237 246239 -1221 246273
rect -867 246239 -851 246273
rect -1237 246131 -1221 246165
rect -867 246131 -851 246165
rect -817 246239 -801 246273
rect -447 246239 -431 246273
rect -817 246131 -801 246165
rect -447 246131 -431 246165
rect -397 246239 -381 246273
rect -27 246239 -11 246273
rect -397 246131 -381 246165
rect -27 246131 -11 246165
rect 23 246239 39 246273
rect 393 246239 409 246273
rect 23 246131 39 246165
rect 393 246131 409 246165
rect 443 246239 459 246273
rect 813 246239 829 246273
rect 443 246131 459 246165
rect 813 246131 829 246165
rect 863 246239 879 246273
rect 1233 246239 1249 246273
rect 863 246131 879 246165
rect 1233 246131 1249 246165
rect 1283 246239 1299 246273
rect 1653 246239 1669 246273
rect 1283 246131 1299 246165
rect 1653 246131 1669 246165
rect 1703 246239 1719 246273
rect 2073 246239 2089 246273
rect 1703 246131 1719 246165
rect 2073 246131 2089 246165
rect 2123 246239 2139 246273
rect 2493 246239 2509 246273
rect 2123 246131 2139 246165
rect 2493 246131 2509 246165
rect 2543 246239 2559 246273
rect 2913 246239 2929 246273
rect 2543 246131 2559 246165
rect 2913 246131 2929 246165
rect 2963 246239 2979 246273
rect 3333 246239 3349 246273
rect 2963 246131 2979 246165
rect 3333 246131 3349 246165
rect 3383 246239 3399 246273
rect 3753 246239 3769 246273
rect 3383 246131 3399 246165
rect 3753 246131 3769 246165
rect 3803 246239 3819 246273
rect 4173 246239 4189 246273
rect 3803 246131 3819 246165
rect 4173 246131 4189 246165
rect 4223 246239 4239 246273
rect 4593 246239 4609 246273
rect 4223 246131 4239 246165
rect 4593 246131 4609 246165
rect 4643 246239 4659 246273
rect 5013 246239 5029 246273
rect 4643 246131 4659 246165
rect 5013 246131 5029 246165
rect 5063 246239 5079 246273
rect 5433 246239 5449 246273
rect 5063 246131 5079 246165
rect 5433 246131 5449 246165
rect 5483 246239 5499 246273
rect 5853 246239 5869 246273
rect 5483 246131 5499 246165
rect 5853 246131 5869 246165
rect 5903 246239 5919 246273
rect 6273 246239 6289 246273
rect 5903 246131 5919 246165
rect 6273 246131 6289 246165
rect 6323 246239 6339 246273
rect 6693 246239 6709 246273
rect 6323 246131 6339 246165
rect 6693 246131 6709 246165
rect 6743 246239 6759 246273
rect 7113 246239 7129 246273
rect 6743 246131 6759 246165
rect 7113 246131 7129 246165
rect 7163 246239 7179 246273
rect 7533 246239 7549 246273
rect 7163 246131 7179 246165
rect 7533 246131 7549 246165
rect 7583 246239 7599 246273
rect 7953 246239 7969 246273
rect 7583 246131 7599 246165
rect 7953 246131 7969 246165
rect 8003 246239 8019 246273
rect 8373 246239 8389 246273
rect 8003 246131 8019 246165
rect 8373 246131 8389 246165
rect 8423 246239 8439 246273
rect 8793 246239 8809 246273
rect 8423 246131 8439 246165
rect 8793 246131 8809 246165
rect 8843 246239 8859 246273
rect 9213 246239 9229 246273
rect 8843 246131 8859 246165
rect 9213 246131 9229 246165
rect 9263 246239 9279 246273
rect 9633 246239 9649 246273
rect 9263 246131 9279 246165
rect 9633 246131 9649 246165
rect 9683 246239 9699 246273
rect 10053 246239 10069 246273
rect 9683 246131 9699 246165
rect 10053 246131 10069 246165
rect 10103 246239 10119 246273
rect 10473 246239 10489 246273
rect 10103 246131 10119 246165
rect 10473 246131 10489 246165
rect 10523 246239 10539 246273
rect 10893 246239 10909 246273
rect 10523 246131 10539 246165
rect 10893 246131 10909 246165
rect 10943 246239 10959 246273
rect 11313 246239 11329 246273
rect 10943 246131 10959 246165
rect 11313 246131 11329 246165
rect 11363 246239 11379 246273
rect 11733 246239 11749 246273
rect 11363 246131 11379 246165
rect 11733 246131 11749 246165
rect 11783 246239 11799 246273
rect 12153 246239 12169 246273
rect 11783 246131 11799 246165
rect 12153 246131 12169 246165
rect 12203 246239 12219 246273
rect 12573 246239 12589 246273
rect 12203 246131 12219 246165
rect 12573 246131 12589 246165
rect 12623 246239 12639 246273
rect 12993 246239 13009 246273
rect 12623 246131 12639 246165
rect 12993 246131 13009 246165
rect 13043 246239 13059 246273
rect 13413 246239 13429 246273
rect 13043 246131 13059 246165
rect 13413 246131 13429 246165
rect 13463 246239 13479 246273
rect 13833 246239 13849 246273
rect 13463 246131 13479 246165
rect 13833 246131 13849 246165
rect 13883 246239 13899 246273
rect 14253 246239 14269 246273
rect 13883 246131 13899 246165
rect 14253 246131 14269 246165
rect 14303 246239 14319 246273
rect 14673 246239 14689 246273
rect 14303 246131 14319 246165
rect 14673 246131 14689 246165
rect 14723 246239 14739 246273
rect 15093 246239 15109 246273
rect 14723 246131 14739 246165
rect 15093 246131 15109 246165
rect 15143 246239 15159 246273
rect 15513 246239 15529 246273
rect 15143 246131 15159 246165
rect 15513 246131 15529 246165
rect 15563 246239 15579 246273
rect 15933 246239 15949 246273
rect 15563 246131 15579 246165
rect 15933 246131 15949 246165
rect 15983 246239 15999 246273
rect 16353 246239 16369 246273
rect 15983 246131 15999 246165
rect 16353 246131 16369 246165
rect 16403 246239 16419 246273
rect 16773 246239 16789 246273
rect 16403 246131 16419 246165
rect 16773 246131 16789 246165
rect 16823 246239 16839 246273
rect 17193 246239 17209 246273
rect 16823 246131 16839 246165
rect 17193 246131 17209 246165
rect 17243 246239 17259 246273
rect 17613 246239 17629 246273
rect 17243 246131 17259 246165
rect 17613 246131 17629 246165
rect 17663 246239 17679 246273
rect 18033 246239 18049 246273
rect 17663 246131 17679 246165
rect 18033 246131 18049 246165
rect 18083 246239 18099 246273
rect 18453 246239 18469 246273
rect 18083 246131 18099 246165
rect 18453 246131 18469 246165
rect 18503 246239 18519 246273
rect 18873 246239 18889 246273
rect 18503 246131 18519 246165
rect 18873 246131 18889 246165
rect 18923 246239 18939 246273
rect 19293 246239 19309 246273
rect 18923 246131 18939 246165
rect 19293 246131 19309 246165
rect 19343 246239 19359 246273
rect 19713 246239 19729 246273
rect 19343 246131 19359 246165
rect 19713 246131 19729 246165
rect 19763 246239 19779 246273
rect 20133 246239 20149 246273
rect 19763 246131 19779 246165
rect 20133 246131 20149 246165
rect 20183 246239 20199 246273
rect 20553 246239 20569 246273
rect 20183 246131 20199 246165
rect 20553 246131 20569 246165
rect 20603 246239 20619 246273
rect 20973 246239 20989 246273
rect 20603 246131 20619 246165
rect 20973 246131 20989 246165
rect 21023 246239 21039 246273
rect 21393 246239 21409 246273
rect 21023 246131 21039 246165
rect 21393 246131 21409 246165
rect 21443 246239 21459 246273
rect 21813 246239 21829 246273
rect 21443 246131 21459 246165
rect 21813 246131 21829 246165
rect 21863 246239 21879 246273
rect 22233 246239 22249 246273
rect 21863 246131 21879 246165
rect 22233 246131 22249 246165
rect 22283 246239 22299 246273
rect 22653 246239 22669 246273
rect 22283 246131 22299 246165
rect 22653 246131 22669 246165
rect 22703 246239 22719 246273
rect 23073 246239 23089 246273
rect 22703 246131 22719 246165
rect 23073 246131 23089 246165
rect 23123 246239 23139 246273
rect 23493 246239 23509 246273
rect 23123 246131 23139 246165
rect 23493 246131 23509 246165
rect 23543 246239 23559 246273
rect 23913 246239 23929 246273
rect 23543 246131 23559 246165
rect 23913 246131 23929 246165
rect 23963 246239 23979 246273
rect 24333 246239 24349 246273
rect 23963 246131 23979 246165
rect 24333 246131 24349 246165
rect 24383 246239 24399 246273
rect 24753 246239 24769 246273
rect 24383 246131 24399 246165
rect 24753 246131 24769 246165
rect 24803 246239 24819 246273
rect 25173 246239 25189 246273
rect 24803 246131 24819 246165
rect 25173 246131 25189 246165
rect 25223 246239 25239 246273
rect 25593 246239 25609 246273
rect 25223 246131 25239 246165
rect 25593 246131 25609 246165
rect 25643 246239 25659 246273
rect 26013 246239 26029 246273
rect 25643 246131 25659 246165
rect 26013 246131 26029 246165
rect 26063 246239 26079 246273
rect 26433 246239 26449 246273
rect 26063 246131 26079 246165
rect 26433 246131 26449 246165
rect 26483 246239 26499 246273
rect 26853 246239 26869 246273
rect 26483 246131 26499 246165
rect 26853 246131 26869 246165
rect 26903 246239 26919 246273
rect 27273 246239 27289 246273
rect 26903 246131 26919 246165
rect 27273 246131 27289 246165
rect 27323 246239 27339 246273
rect 27323 246131 27339 246165
rect -4049 246072 -4015 246088
rect -4049 245280 -4015 245296
rect -3953 246072 -3919 246088
rect -3953 245280 -3919 245296
rect -3839 246072 -3805 246088
rect -3839 245280 -3805 245296
rect -3743 246072 -3709 246088
rect -3743 245280 -3709 245296
rect -3629 246072 -3595 246088
rect -3629 245280 -3595 245296
rect -3533 246072 -3499 246088
rect -3533 245280 -3499 245296
rect -3419 246072 -3385 246088
rect -3419 245280 -3385 245296
rect -3323 246072 -3289 246088
rect -3323 245280 -3289 245296
rect -3209 246072 -3175 246088
rect -3209 245280 -3175 245296
rect -3113 246072 -3079 246088
rect -3113 245280 -3079 245296
rect -2999 246072 -2965 246088
rect -2999 245280 -2965 245296
rect -2903 246072 -2869 246088
rect -2903 245280 -2869 245296
rect -2789 246072 -2755 246088
rect -2789 245280 -2755 245296
rect -2693 246072 -2659 246088
rect -2693 245280 -2659 245296
rect -2579 246072 -2545 246088
rect -2579 245280 -2545 245296
rect -2483 246072 -2449 246088
rect -2483 245280 -2449 245296
rect -2369 246072 -2335 246088
rect -2369 245280 -2335 245296
rect -2273 246072 -2239 246088
rect -2273 245280 -2239 245296
rect -2159 246072 -2125 246088
rect -2159 245280 -2125 245296
rect -2063 246072 -2029 246088
rect -2063 245280 -2029 245296
rect -1949 246072 -1915 246088
rect -1949 245280 -1915 245296
rect -1853 246072 -1819 246088
rect -1853 245280 -1819 245296
rect -1739 246072 -1705 246088
rect -1739 245280 -1705 245296
rect -1643 246072 -1609 246088
rect -1643 245280 -1609 245296
rect -1529 246072 -1495 246088
rect -1529 245280 -1495 245296
rect -1433 246072 -1399 246088
rect -1433 245280 -1399 245296
rect -1319 246072 -1285 246088
rect -1319 245280 -1285 245296
rect -1223 246072 -1189 246088
rect -1223 245280 -1189 245296
rect -1109 246072 -1075 246088
rect -1109 245280 -1075 245296
rect -1013 246072 -979 246088
rect -1013 245280 -979 245296
rect -899 246072 -865 246088
rect -899 245280 -865 245296
rect -803 246072 -769 246088
rect -803 245280 -769 245296
rect -689 246072 -655 246088
rect -689 245280 -655 245296
rect -593 246072 -559 246088
rect -593 245280 -559 245296
rect -479 246072 -445 246088
rect -479 245280 -445 245296
rect -383 246072 -349 246088
rect -383 245280 -349 245296
rect -269 246072 -235 246088
rect -269 245280 -235 245296
rect -173 246072 -139 246088
rect -173 245280 -139 245296
rect -59 246072 -25 246088
rect -59 245280 -25 245296
rect 37 246072 71 246088
rect 37 245280 71 245296
rect 151 246072 185 246088
rect 151 245280 185 245296
rect 247 246072 281 246088
rect 247 245280 281 245296
rect 361 246072 395 246088
rect 361 245280 395 245296
rect 457 246072 491 246088
rect 457 245280 491 245296
rect 571 246072 605 246088
rect 571 245280 605 245296
rect 667 246072 701 246088
rect 667 245280 701 245296
rect 781 246072 815 246088
rect 781 245280 815 245296
rect 877 246072 911 246088
rect 877 245280 911 245296
rect 991 246072 1025 246088
rect 991 245280 1025 245296
rect 1087 246072 1121 246088
rect 1087 245280 1121 245296
rect 1201 246072 1235 246088
rect 1201 245280 1235 245296
rect 1297 246072 1331 246088
rect 1297 245280 1331 245296
rect 1411 246072 1445 246088
rect 1411 245280 1445 245296
rect 1507 246072 1541 246088
rect 1507 245280 1541 245296
rect 1621 246072 1655 246088
rect 1621 245280 1655 245296
rect 1717 246072 1751 246088
rect 1717 245280 1751 245296
rect 1831 246072 1865 246088
rect 1831 245280 1865 245296
rect 1927 246072 1961 246088
rect 1927 245280 1961 245296
rect 2041 246072 2075 246088
rect 2041 245280 2075 245296
rect 2137 246072 2171 246088
rect 2137 245280 2171 245296
rect 2251 246072 2285 246088
rect 2251 245280 2285 245296
rect 2347 246072 2381 246088
rect 2347 245280 2381 245296
rect 2461 246072 2495 246088
rect 2461 245280 2495 245296
rect 2557 246072 2591 246088
rect 2557 245280 2591 245296
rect 2671 246072 2705 246088
rect 2671 245280 2705 245296
rect 2767 246072 2801 246088
rect 2767 245280 2801 245296
rect 2881 246072 2915 246088
rect 2881 245280 2915 245296
rect 2977 246072 3011 246088
rect 2977 245280 3011 245296
rect 3091 246072 3125 246088
rect 3091 245280 3125 245296
rect 3187 246072 3221 246088
rect 3187 245280 3221 245296
rect 3301 246072 3335 246088
rect 3301 245280 3335 245296
rect 3397 246072 3431 246088
rect 3397 245280 3431 245296
rect 3511 246072 3545 246088
rect 3511 245280 3545 245296
rect 3607 246072 3641 246088
rect 3607 245280 3641 245296
rect 3721 246072 3755 246088
rect 3721 245280 3755 245296
rect 3817 246072 3851 246088
rect 3817 245280 3851 245296
rect 3931 246072 3965 246088
rect 3931 245280 3965 245296
rect 4027 246072 4061 246088
rect 4027 245280 4061 245296
rect 4141 246072 4175 246088
rect 4141 245280 4175 245296
rect 4237 246072 4271 246088
rect 4237 245280 4271 245296
rect 4351 246072 4385 246088
rect 4351 245280 4385 245296
rect 4447 246072 4481 246088
rect 4447 245280 4481 245296
rect 4561 246072 4595 246088
rect 4561 245280 4595 245296
rect 4657 246072 4691 246088
rect 4657 245280 4691 245296
rect 4771 246072 4805 246088
rect 4771 245280 4805 245296
rect 4867 246072 4901 246088
rect 4867 245280 4901 245296
rect 4981 246072 5015 246088
rect 4981 245280 5015 245296
rect 5077 246072 5111 246088
rect 5077 245280 5111 245296
rect 5191 246072 5225 246088
rect 5191 245280 5225 245296
rect 5287 246072 5321 246088
rect 5287 245280 5321 245296
rect 5401 246072 5435 246088
rect 5401 245280 5435 245296
rect 5497 246072 5531 246088
rect 5497 245280 5531 245296
rect 5611 246072 5645 246088
rect 5611 245280 5645 245296
rect 5707 246072 5741 246088
rect 5707 245280 5741 245296
rect 5821 246072 5855 246088
rect 5821 245280 5855 245296
rect 5917 246072 5951 246088
rect 5917 245280 5951 245296
rect 6031 246072 6065 246088
rect 6031 245280 6065 245296
rect 6127 246072 6161 246088
rect 6127 245280 6161 245296
rect 6241 246072 6275 246088
rect 6241 245280 6275 245296
rect 6337 246072 6371 246088
rect 6337 245280 6371 245296
rect 6451 246072 6485 246088
rect 6451 245280 6485 245296
rect 6547 246072 6581 246088
rect 6547 245280 6581 245296
rect 6661 246072 6695 246088
rect 6661 245280 6695 245296
rect 6757 246072 6791 246088
rect 6757 245280 6791 245296
rect 6871 246072 6905 246088
rect 6871 245280 6905 245296
rect 6967 246072 7001 246088
rect 6967 245280 7001 245296
rect 7081 246072 7115 246088
rect 7081 245280 7115 245296
rect 7177 246072 7211 246088
rect 7177 245280 7211 245296
rect 7291 246072 7325 246088
rect 7291 245280 7325 245296
rect 7387 246072 7421 246088
rect 7387 245280 7421 245296
rect 7501 246072 7535 246088
rect 7501 245280 7535 245296
rect 7597 246072 7631 246088
rect 7597 245280 7631 245296
rect 7711 246072 7745 246088
rect 7711 245280 7745 245296
rect 7807 246072 7841 246088
rect 7807 245280 7841 245296
rect 7921 246072 7955 246088
rect 7921 245280 7955 245296
rect 8017 246072 8051 246088
rect 8017 245280 8051 245296
rect 8131 246072 8165 246088
rect 8131 245280 8165 245296
rect 8227 246072 8261 246088
rect 8227 245280 8261 245296
rect 8341 246072 8375 246088
rect 8341 245280 8375 245296
rect 8437 246072 8471 246088
rect 8437 245280 8471 245296
rect 8551 246072 8585 246088
rect 8551 245280 8585 245296
rect 8647 246072 8681 246088
rect 8647 245280 8681 245296
rect 8761 246072 8795 246088
rect 8761 245280 8795 245296
rect 8857 246072 8891 246088
rect 8857 245280 8891 245296
rect 8971 246072 9005 246088
rect 8971 245280 9005 245296
rect 9067 246072 9101 246088
rect 9067 245280 9101 245296
rect 9181 246072 9215 246088
rect 9181 245280 9215 245296
rect 9277 246072 9311 246088
rect 9277 245280 9311 245296
rect 9391 246072 9425 246088
rect 9391 245280 9425 245296
rect 9487 246072 9521 246088
rect 9487 245280 9521 245296
rect 9601 246072 9635 246088
rect 9601 245280 9635 245296
rect 9697 246072 9731 246088
rect 9697 245280 9731 245296
rect 9811 246072 9845 246088
rect 9811 245280 9845 245296
rect 9907 246072 9941 246088
rect 9907 245280 9941 245296
rect 10021 246072 10055 246088
rect 10021 245280 10055 245296
rect 10117 246072 10151 246088
rect 10117 245280 10151 245296
rect 10231 246072 10265 246088
rect 10231 245280 10265 245296
rect 10327 246072 10361 246088
rect 10327 245280 10361 245296
rect 10441 246072 10475 246088
rect 10441 245280 10475 245296
rect 10537 246072 10571 246088
rect 10537 245280 10571 245296
rect 10651 246072 10685 246088
rect 10651 245280 10685 245296
rect 10747 246072 10781 246088
rect 10747 245280 10781 245296
rect 10861 246072 10895 246088
rect 10861 245280 10895 245296
rect 10957 246072 10991 246088
rect 10957 245280 10991 245296
rect 11071 246072 11105 246088
rect 11071 245280 11105 245296
rect 11167 246072 11201 246088
rect 11167 245280 11201 245296
rect 11281 246072 11315 246088
rect 11281 245280 11315 245296
rect 11377 246072 11411 246088
rect 11377 245280 11411 245296
rect 11491 246072 11525 246088
rect 11491 245280 11525 245296
rect 11587 246072 11621 246088
rect 11587 245280 11621 245296
rect 11701 246072 11735 246088
rect 11701 245280 11735 245296
rect 11797 246072 11831 246088
rect 11797 245280 11831 245296
rect 11911 246072 11945 246088
rect 11911 245280 11945 245296
rect 12007 246072 12041 246088
rect 12007 245280 12041 245296
rect 12121 246072 12155 246088
rect 12121 245280 12155 245296
rect 12217 246072 12251 246088
rect 12217 245280 12251 245296
rect 12331 246072 12365 246088
rect 12331 245280 12365 245296
rect 12427 246072 12461 246088
rect 12427 245280 12461 245296
rect 12541 246072 12575 246088
rect 12541 245280 12575 245296
rect 12637 246072 12671 246088
rect 12637 245280 12671 245296
rect 12751 246072 12785 246088
rect 12751 245280 12785 245296
rect 12847 246072 12881 246088
rect 12847 245280 12881 245296
rect 12961 246072 12995 246088
rect 12961 245280 12995 245296
rect 13057 246072 13091 246088
rect 13057 245280 13091 245296
rect 13171 246072 13205 246088
rect 13171 245280 13205 245296
rect 13267 246072 13301 246088
rect 13267 245280 13301 245296
rect 13381 246072 13415 246088
rect 13381 245280 13415 245296
rect 13477 246072 13511 246088
rect 13477 245280 13511 245296
rect 13591 246072 13625 246088
rect 13591 245280 13625 245296
rect 13687 246072 13721 246088
rect 13687 245280 13721 245296
rect 13801 246072 13835 246088
rect 13801 245280 13835 245296
rect 13897 246072 13931 246088
rect 13897 245280 13931 245296
rect 14011 246072 14045 246088
rect 14011 245280 14045 245296
rect 14107 246072 14141 246088
rect 14107 245280 14141 245296
rect 14221 246072 14255 246088
rect 14221 245280 14255 245296
rect 14317 246072 14351 246088
rect 14317 245280 14351 245296
rect 14431 246072 14465 246088
rect 14431 245280 14465 245296
rect 14527 246072 14561 246088
rect 14527 245280 14561 245296
rect 14641 246072 14675 246088
rect 14641 245280 14675 245296
rect 14737 246072 14771 246088
rect 14737 245280 14771 245296
rect 14851 246072 14885 246088
rect 14851 245280 14885 245296
rect 14947 246072 14981 246088
rect 14947 245280 14981 245296
rect 15061 246072 15095 246088
rect 15061 245280 15095 245296
rect 15157 246072 15191 246088
rect 15157 245280 15191 245296
rect 15271 246072 15305 246088
rect 15271 245280 15305 245296
rect 15367 246072 15401 246088
rect 15367 245280 15401 245296
rect 15481 246072 15515 246088
rect 15481 245280 15515 245296
rect 15577 246072 15611 246088
rect 15577 245280 15611 245296
rect 15691 246072 15725 246088
rect 15691 245280 15725 245296
rect 15787 246072 15821 246088
rect 15787 245280 15821 245296
rect 15901 246072 15935 246088
rect 15901 245280 15935 245296
rect 15997 246072 16031 246088
rect 15997 245280 16031 245296
rect 16111 246072 16145 246088
rect 16111 245280 16145 245296
rect 16207 246072 16241 246088
rect 16207 245280 16241 245296
rect 16321 246072 16355 246088
rect 16321 245280 16355 245296
rect 16417 246072 16451 246088
rect 16417 245280 16451 245296
rect 16531 246072 16565 246088
rect 16531 245280 16565 245296
rect 16627 246072 16661 246088
rect 16627 245280 16661 245296
rect 16741 246072 16775 246088
rect 16741 245280 16775 245296
rect 16837 246072 16871 246088
rect 16837 245280 16871 245296
rect 16951 246072 16985 246088
rect 16951 245280 16985 245296
rect 17047 246072 17081 246088
rect 17047 245280 17081 245296
rect 17161 246072 17195 246088
rect 17161 245280 17195 245296
rect 17257 246072 17291 246088
rect 17257 245280 17291 245296
rect 17371 246072 17405 246088
rect 17371 245280 17405 245296
rect 17467 246072 17501 246088
rect 17467 245280 17501 245296
rect 17581 246072 17615 246088
rect 17581 245280 17615 245296
rect 17677 246072 17711 246088
rect 17677 245280 17711 245296
rect 17791 246072 17825 246088
rect 17791 245280 17825 245296
rect 17887 246072 17921 246088
rect 17887 245280 17921 245296
rect 18001 246072 18035 246088
rect 18001 245280 18035 245296
rect 18097 246072 18131 246088
rect 18097 245280 18131 245296
rect 18211 246072 18245 246088
rect 18211 245280 18245 245296
rect 18307 246072 18341 246088
rect 18307 245280 18341 245296
rect 18421 246072 18455 246088
rect 18421 245280 18455 245296
rect 18517 246072 18551 246088
rect 18517 245280 18551 245296
rect 18631 246072 18665 246088
rect 18631 245280 18665 245296
rect 18727 246072 18761 246088
rect 18727 245280 18761 245296
rect 18841 246072 18875 246088
rect 18841 245280 18875 245296
rect 18937 246072 18971 246088
rect 18937 245280 18971 245296
rect 19051 246072 19085 246088
rect 19051 245280 19085 245296
rect 19147 246072 19181 246088
rect 19147 245280 19181 245296
rect 19261 246072 19295 246088
rect 19261 245280 19295 245296
rect 19357 246072 19391 246088
rect 19357 245280 19391 245296
rect 19471 246072 19505 246088
rect 19471 245280 19505 245296
rect 19567 246072 19601 246088
rect 19567 245280 19601 245296
rect 19681 246072 19715 246088
rect 19681 245280 19715 245296
rect 19777 246072 19811 246088
rect 19777 245280 19811 245296
rect 19891 246072 19925 246088
rect 19891 245280 19925 245296
rect 19987 246072 20021 246088
rect 19987 245280 20021 245296
rect 20101 246072 20135 246088
rect 20101 245280 20135 245296
rect 20197 246072 20231 246088
rect 20197 245280 20231 245296
rect 20311 246072 20345 246088
rect 20311 245280 20345 245296
rect 20407 246072 20441 246088
rect 20407 245280 20441 245296
rect 20521 246072 20555 246088
rect 20521 245280 20555 245296
rect 20617 246072 20651 246088
rect 20617 245280 20651 245296
rect 20731 246072 20765 246088
rect 20731 245280 20765 245296
rect 20827 246072 20861 246088
rect 20827 245280 20861 245296
rect 20941 246072 20975 246088
rect 20941 245280 20975 245296
rect 21037 246072 21071 246088
rect 21037 245280 21071 245296
rect 21151 246072 21185 246088
rect 21151 245280 21185 245296
rect 21247 246072 21281 246088
rect 21247 245280 21281 245296
rect 21361 246072 21395 246088
rect 21361 245280 21395 245296
rect 21457 246072 21491 246088
rect 21457 245280 21491 245296
rect 21571 246072 21605 246088
rect 21571 245280 21605 245296
rect 21667 246072 21701 246088
rect 21667 245280 21701 245296
rect 21781 246072 21815 246088
rect 21781 245280 21815 245296
rect 21877 246072 21911 246088
rect 21877 245280 21911 245296
rect 21991 246072 22025 246088
rect 21991 245280 22025 245296
rect 22087 246072 22121 246088
rect 22087 245280 22121 245296
rect 22201 246072 22235 246088
rect 22201 245280 22235 245296
rect 22297 246072 22331 246088
rect 22297 245280 22331 245296
rect 22411 246072 22445 246088
rect 22411 245280 22445 245296
rect 22507 246072 22541 246088
rect 22507 245280 22541 245296
rect 22621 246072 22655 246088
rect 22621 245280 22655 245296
rect 22717 246072 22751 246088
rect 22717 245280 22751 245296
rect 22831 246072 22865 246088
rect 22831 245280 22865 245296
rect 22927 246072 22961 246088
rect 22927 245280 22961 245296
rect 23041 246072 23075 246088
rect 23041 245280 23075 245296
rect 23137 246072 23171 246088
rect 23137 245280 23171 245296
rect 23251 246072 23285 246088
rect 23251 245280 23285 245296
rect 23347 246072 23381 246088
rect 23347 245280 23381 245296
rect 23461 246072 23495 246088
rect 23461 245280 23495 245296
rect 23557 246072 23591 246088
rect 23557 245280 23591 245296
rect 23671 246072 23705 246088
rect 23671 245280 23705 245296
rect 23767 246072 23801 246088
rect 23767 245280 23801 245296
rect 23881 246072 23915 246088
rect 23881 245280 23915 245296
rect 23977 246072 24011 246088
rect 23977 245280 24011 245296
rect 24091 246072 24125 246088
rect 24091 245280 24125 245296
rect 24187 246072 24221 246088
rect 24187 245280 24221 245296
rect 24301 246072 24335 246088
rect 24301 245280 24335 245296
rect 24397 246072 24431 246088
rect 24397 245280 24431 245296
rect 24511 246072 24545 246088
rect 24511 245280 24545 245296
rect 24607 246072 24641 246088
rect 24607 245280 24641 245296
rect 24721 246072 24755 246088
rect 24721 245280 24755 245296
rect 24817 246072 24851 246088
rect 24817 245280 24851 245296
rect 24931 246072 24965 246088
rect 24931 245280 24965 245296
rect 25027 246072 25061 246088
rect 25027 245280 25061 245296
rect 25141 246072 25175 246088
rect 25141 245280 25175 245296
rect 25237 246072 25271 246088
rect 25237 245280 25271 245296
rect 25351 246072 25385 246088
rect 25351 245280 25385 245296
rect 25447 246072 25481 246088
rect 25447 245280 25481 245296
rect 25561 246072 25595 246088
rect 25561 245280 25595 245296
rect 25657 246072 25691 246088
rect 25657 245280 25691 245296
rect 25771 246072 25805 246088
rect 25771 245280 25805 245296
rect 25867 246072 25901 246088
rect 25867 245280 25901 245296
rect 25981 246072 26015 246088
rect 25981 245280 26015 245296
rect 26077 246072 26111 246088
rect 26077 245280 26111 245296
rect 26191 246072 26225 246088
rect 26191 245280 26225 245296
rect 26287 246072 26321 246088
rect 26287 245280 26321 245296
rect 26401 246072 26435 246088
rect 26401 245280 26435 245296
rect 26497 246072 26531 246088
rect 26497 245280 26531 245296
rect 26611 246072 26645 246088
rect 26611 245280 26645 245296
rect 26707 246072 26741 246088
rect 26707 245280 26741 245296
rect 26821 246072 26855 246088
rect 26821 245280 26855 245296
rect 26917 246072 26951 246088
rect 26917 245280 26951 245296
rect 27031 246072 27065 246088
rect 27031 245280 27065 245296
rect 27127 246072 27161 246088
rect 27127 245280 27161 245296
rect 27241 246072 27275 246088
rect 27241 245280 27275 245296
rect 27337 246072 27371 246088
rect 27337 245280 27371 245296
rect -4017 245203 -4001 245237
rect -4017 245095 -4001 245129
rect -3967 245203 -3951 245237
rect -3597 245203 -3581 245237
rect -3967 245095 -3951 245129
rect -3597 245095 -3581 245129
rect -3547 245203 -3531 245237
rect -3177 245203 -3161 245237
rect -3547 245095 -3531 245129
rect -3177 245095 -3161 245129
rect -3127 245203 -3111 245237
rect -2757 245203 -2741 245237
rect -3127 245095 -3111 245129
rect -2757 245095 -2741 245129
rect -2707 245203 -2691 245237
rect -2337 245203 -2321 245237
rect -2707 245095 -2691 245129
rect -2337 245095 -2321 245129
rect -2287 245203 -2271 245237
rect -1917 245203 -1901 245237
rect -2287 245095 -2271 245129
rect -1917 245095 -1901 245129
rect -1867 245203 -1851 245237
rect -1497 245203 -1481 245237
rect -1867 245095 -1851 245129
rect -1497 245095 -1481 245129
rect -1447 245203 -1431 245237
rect -1077 245203 -1061 245237
rect -1447 245095 -1431 245129
rect -1077 245095 -1061 245129
rect -1027 245203 -1011 245237
rect -657 245203 -641 245237
rect -1027 245095 -1011 245129
rect -657 245095 -641 245129
rect -607 245203 -591 245237
rect -237 245203 -221 245237
rect -607 245095 -591 245129
rect -237 245095 -221 245129
rect -187 245203 -171 245237
rect 183 245203 199 245237
rect -187 245095 -171 245129
rect 183 245095 199 245129
rect 233 245203 249 245237
rect 603 245203 619 245237
rect 233 245095 249 245129
rect 603 245095 619 245129
rect 653 245203 669 245237
rect 1023 245203 1039 245237
rect 653 245095 669 245129
rect 1023 245095 1039 245129
rect 1073 245203 1089 245237
rect 1443 245203 1459 245237
rect 1073 245095 1089 245129
rect 1443 245095 1459 245129
rect 1493 245203 1509 245237
rect 1863 245203 1879 245237
rect 1493 245095 1509 245129
rect 1863 245095 1879 245129
rect 1913 245203 1929 245237
rect 2283 245203 2299 245237
rect 1913 245095 1929 245129
rect 2283 245095 2299 245129
rect 2333 245203 2349 245237
rect 2703 245203 2719 245237
rect 2333 245095 2349 245129
rect 2703 245095 2719 245129
rect 2753 245203 2769 245237
rect 3123 245203 3139 245237
rect 2753 245095 2769 245129
rect 3123 245095 3139 245129
rect 3173 245203 3189 245237
rect 3543 245203 3559 245237
rect 3173 245095 3189 245129
rect 3543 245095 3559 245129
rect 3593 245203 3609 245237
rect 3963 245203 3979 245237
rect 3593 245095 3609 245129
rect 3963 245095 3979 245129
rect 4013 245203 4029 245237
rect 4383 245203 4399 245237
rect 4013 245095 4029 245129
rect 4383 245095 4399 245129
rect 4433 245203 4449 245237
rect 4803 245203 4819 245237
rect 4433 245095 4449 245129
rect 4803 245095 4819 245129
rect 4853 245203 4869 245237
rect 5223 245203 5239 245237
rect 4853 245095 4869 245129
rect 5223 245095 5239 245129
rect 5273 245203 5289 245237
rect 5643 245203 5659 245237
rect 5273 245095 5289 245129
rect 5643 245095 5659 245129
rect 5693 245203 5709 245237
rect 6063 245203 6079 245237
rect 5693 245095 5709 245129
rect 6063 245095 6079 245129
rect 6113 245203 6129 245237
rect 6483 245203 6499 245237
rect 6113 245095 6129 245129
rect 6483 245095 6499 245129
rect 6533 245203 6549 245237
rect 6903 245203 6919 245237
rect 6533 245095 6549 245129
rect 6903 245095 6919 245129
rect 6953 245203 6969 245237
rect 7323 245203 7339 245237
rect 6953 245095 6969 245129
rect 7323 245095 7339 245129
rect 7373 245203 7389 245237
rect 7743 245203 7759 245237
rect 7373 245095 7389 245129
rect 7743 245095 7759 245129
rect 7793 245203 7809 245237
rect 8163 245203 8179 245237
rect 7793 245095 7809 245129
rect 8163 245095 8179 245129
rect 8213 245203 8229 245237
rect 8583 245203 8599 245237
rect 8213 245095 8229 245129
rect 8583 245095 8599 245129
rect 8633 245203 8649 245237
rect 9003 245203 9019 245237
rect 8633 245095 8649 245129
rect 9003 245095 9019 245129
rect 9053 245203 9069 245237
rect 9423 245203 9439 245237
rect 9053 245095 9069 245129
rect 9423 245095 9439 245129
rect 9473 245203 9489 245237
rect 9843 245203 9859 245237
rect 9473 245095 9489 245129
rect 9843 245095 9859 245129
rect 9893 245203 9909 245237
rect 10263 245203 10279 245237
rect 9893 245095 9909 245129
rect 10263 245095 10279 245129
rect 10313 245203 10329 245237
rect 10683 245203 10699 245237
rect 10313 245095 10329 245129
rect 10683 245095 10699 245129
rect 10733 245203 10749 245237
rect 11103 245203 11119 245237
rect 10733 245095 10749 245129
rect 11103 245095 11119 245129
rect 11153 245203 11169 245237
rect 11523 245203 11539 245237
rect 11153 245095 11169 245129
rect 11523 245095 11539 245129
rect 11573 245203 11589 245237
rect 11943 245203 11959 245237
rect 11573 245095 11589 245129
rect 11943 245095 11959 245129
rect 11993 245203 12009 245237
rect 12363 245203 12379 245237
rect 11993 245095 12009 245129
rect 12363 245095 12379 245129
rect 12413 245203 12429 245237
rect 12783 245203 12799 245237
rect 12413 245095 12429 245129
rect 12783 245095 12799 245129
rect 12833 245203 12849 245237
rect 13203 245203 13219 245237
rect 12833 245095 12849 245129
rect 13203 245095 13219 245129
rect 13253 245203 13269 245237
rect 13623 245203 13639 245237
rect 13253 245095 13269 245129
rect 13623 245095 13639 245129
rect 13673 245203 13689 245237
rect 14043 245203 14059 245237
rect 13673 245095 13689 245129
rect 14043 245095 14059 245129
rect 14093 245203 14109 245237
rect 14463 245203 14479 245237
rect 14093 245095 14109 245129
rect 14463 245095 14479 245129
rect 14513 245203 14529 245237
rect 14883 245203 14899 245237
rect 14513 245095 14529 245129
rect 14883 245095 14899 245129
rect 14933 245203 14949 245237
rect 15303 245203 15319 245237
rect 14933 245095 14949 245129
rect 15303 245095 15319 245129
rect 15353 245203 15369 245237
rect 15723 245203 15739 245237
rect 15353 245095 15369 245129
rect 15723 245095 15739 245129
rect 15773 245203 15789 245237
rect 16143 245203 16159 245237
rect 15773 245095 15789 245129
rect 16143 245095 16159 245129
rect 16193 245203 16209 245237
rect 16563 245203 16579 245237
rect 16193 245095 16209 245129
rect 16563 245095 16579 245129
rect 16613 245203 16629 245237
rect 16983 245203 16999 245237
rect 16613 245095 16629 245129
rect 16983 245095 16999 245129
rect 17033 245203 17049 245237
rect 17403 245203 17419 245237
rect 17033 245095 17049 245129
rect 17403 245095 17419 245129
rect 17453 245203 17469 245237
rect 17823 245203 17839 245237
rect 17453 245095 17469 245129
rect 17823 245095 17839 245129
rect 17873 245203 17889 245237
rect 18243 245203 18259 245237
rect 17873 245095 17889 245129
rect 18243 245095 18259 245129
rect 18293 245203 18309 245237
rect 18663 245203 18679 245237
rect 18293 245095 18309 245129
rect 18663 245095 18679 245129
rect 18713 245203 18729 245237
rect 19083 245203 19099 245237
rect 18713 245095 18729 245129
rect 19083 245095 19099 245129
rect 19133 245203 19149 245237
rect 19503 245203 19519 245237
rect 19133 245095 19149 245129
rect 19503 245095 19519 245129
rect 19553 245203 19569 245237
rect 19923 245203 19939 245237
rect 19553 245095 19569 245129
rect 19923 245095 19939 245129
rect 19973 245203 19989 245237
rect 20343 245203 20359 245237
rect 19973 245095 19989 245129
rect 20343 245095 20359 245129
rect 20393 245203 20409 245237
rect 20763 245203 20779 245237
rect 20393 245095 20409 245129
rect 20763 245095 20779 245129
rect 20813 245203 20829 245237
rect 21183 245203 21199 245237
rect 20813 245095 20829 245129
rect 21183 245095 21199 245129
rect 21233 245203 21249 245237
rect 21603 245203 21619 245237
rect 21233 245095 21249 245129
rect 21603 245095 21619 245129
rect 21653 245203 21669 245237
rect 22023 245203 22039 245237
rect 21653 245095 21669 245129
rect 22023 245095 22039 245129
rect 22073 245203 22089 245237
rect 22443 245203 22459 245237
rect 22073 245095 22089 245129
rect 22443 245095 22459 245129
rect 22493 245203 22509 245237
rect 22863 245203 22879 245237
rect 22493 245095 22509 245129
rect 22863 245095 22879 245129
rect 22913 245203 22929 245237
rect 23283 245203 23299 245237
rect 22913 245095 22929 245129
rect 23283 245095 23299 245129
rect 23333 245203 23349 245237
rect 23703 245203 23719 245237
rect 23333 245095 23349 245129
rect 23703 245095 23719 245129
rect 23753 245203 23769 245237
rect 24123 245203 24139 245237
rect 23753 245095 23769 245129
rect 24123 245095 24139 245129
rect 24173 245203 24189 245237
rect 24543 245203 24559 245237
rect 24173 245095 24189 245129
rect 24543 245095 24559 245129
rect 24593 245203 24609 245237
rect 24963 245203 24979 245237
rect 24593 245095 24609 245129
rect 24963 245095 24979 245129
rect 25013 245203 25029 245237
rect 25383 245203 25399 245237
rect 25013 245095 25029 245129
rect 25383 245095 25399 245129
rect 25433 245203 25449 245237
rect 25803 245203 25819 245237
rect 25433 245095 25449 245129
rect 25803 245095 25819 245129
rect 25853 245203 25869 245237
rect 26223 245203 26239 245237
rect 25853 245095 25869 245129
rect 26223 245095 26239 245129
rect 26273 245203 26289 245237
rect 26643 245203 26659 245237
rect 26273 245095 26289 245129
rect 26643 245095 26659 245129
rect 26693 245203 26709 245237
rect 27063 245203 27079 245237
rect 26693 245095 26709 245129
rect 27063 245095 27079 245129
rect 27113 245203 27129 245237
rect 27113 245095 27129 245129
rect -4049 245036 -4015 245052
rect -4049 244244 -4015 244260
rect -3953 245036 -3919 245052
rect -3953 244244 -3919 244260
rect -3839 245036 -3805 245052
rect -3839 244244 -3805 244260
rect -3743 245036 -3709 245052
rect -3743 244244 -3709 244260
rect -3629 245036 -3595 245052
rect -3629 244244 -3595 244260
rect -3533 245036 -3499 245052
rect -3533 244244 -3499 244260
rect -3419 245036 -3385 245052
rect -3419 244244 -3385 244260
rect -3323 245036 -3289 245052
rect -3323 244244 -3289 244260
rect -3209 245036 -3175 245052
rect -3209 244244 -3175 244260
rect -3113 245036 -3079 245052
rect -3113 244244 -3079 244260
rect -2999 245036 -2965 245052
rect -2999 244244 -2965 244260
rect -2903 245036 -2869 245052
rect -2903 244244 -2869 244260
rect -2789 245036 -2755 245052
rect -2789 244244 -2755 244260
rect -2693 245036 -2659 245052
rect -2693 244244 -2659 244260
rect -2579 245036 -2545 245052
rect -2579 244244 -2545 244260
rect -2483 245036 -2449 245052
rect -2483 244244 -2449 244260
rect -2369 245036 -2335 245052
rect -2369 244244 -2335 244260
rect -2273 245036 -2239 245052
rect -2273 244244 -2239 244260
rect -2159 245036 -2125 245052
rect -2159 244244 -2125 244260
rect -2063 245036 -2029 245052
rect -2063 244244 -2029 244260
rect -1949 245036 -1915 245052
rect -1949 244244 -1915 244260
rect -1853 245036 -1819 245052
rect -1853 244244 -1819 244260
rect -1739 245036 -1705 245052
rect -1739 244244 -1705 244260
rect -1643 245036 -1609 245052
rect -1643 244244 -1609 244260
rect -1529 245036 -1495 245052
rect -1529 244244 -1495 244260
rect -1433 245036 -1399 245052
rect -1433 244244 -1399 244260
rect -1319 245036 -1285 245052
rect -1319 244244 -1285 244260
rect -1223 245036 -1189 245052
rect -1223 244244 -1189 244260
rect -1109 245036 -1075 245052
rect -1109 244244 -1075 244260
rect -1013 245036 -979 245052
rect -1013 244244 -979 244260
rect -899 245036 -865 245052
rect -899 244244 -865 244260
rect -803 245036 -769 245052
rect -803 244244 -769 244260
rect -689 245036 -655 245052
rect -689 244244 -655 244260
rect -593 245036 -559 245052
rect -593 244244 -559 244260
rect -479 245036 -445 245052
rect -479 244244 -445 244260
rect -383 245036 -349 245052
rect -383 244244 -349 244260
rect -269 245036 -235 245052
rect -269 244244 -235 244260
rect -173 245036 -139 245052
rect -173 244244 -139 244260
rect -59 245036 -25 245052
rect -59 244244 -25 244260
rect 37 245036 71 245052
rect 37 244244 71 244260
rect 151 245036 185 245052
rect 151 244244 185 244260
rect 247 245036 281 245052
rect 247 244244 281 244260
rect 361 245036 395 245052
rect 361 244244 395 244260
rect 457 245036 491 245052
rect 457 244244 491 244260
rect 571 245036 605 245052
rect 571 244244 605 244260
rect 667 245036 701 245052
rect 667 244244 701 244260
rect 781 245036 815 245052
rect 781 244244 815 244260
rect 877 245036 911 245052
rect 877 244244 911 244260
rect 991 245036 1025 245052
rect 991 244244 1025 244260
rect 1087 245036 1121 245052
rect 1087 244244 1121 244260
rect 1201 245036 1235 245052
rect 1201 244244 1235 244260
rect 1297 245036 1331 245052
rect 1297 244244 1331 244260
rect 1411 245036 1445 245052
rect 1411 244244 1445 244260
rect 1507 245036 1541 245052
rect 1507 244244 1541 244260
rect 1621 245036 1655 245052
rect 1621 244244 1655 244260
rect 1717 245036 1751 245052
rect 1717 244244 1751 244260
rect 1831 245036 1865 245052
rect 1831 244244 1865 244260
rect 1927 245036 1961 245052
rect 1927 244244 1961 244260
rect 2041 245036 2075 245052
rect 2041 244244 2075 244260
rect 2137 245036 2171 245052
rect 2137 244244 2171 244260
rect 2251 245036 2285 245052
rect 2251 244244 2285 244260
rect 2347 245036 2381 245052
rect 2347 244244 2381 244260
rect 2461 245036 2495 245052
rect 2461 244244 2495 244260
rect 2557 245036 2591 245052
rect 2557 244244 2591 244260
rect 2671 245036 2705 245052
rect 2671 244244 2705 244260
rect 2767 245036 2801 245052
rect 2767 244244 2801 244260
rect 2881 245036 2915 245052
rect 2881 244244 2915 244260
rect 2977 245036 3011 245052
rect 2977 244244 3011 244260
rect 3091 245036 3125 245052
rect 3091 244244 3125 244260
rect 3187 245036 3221 245052
rect 3187 244244 3221 244260
rect 3301 245036 3335 245052
rect 3301 244244 3335 244260
rect 3397 245036 3431 245052
rect 3397 244244 3431 244260
rect 3511 245036 3545 245052
rect 3511 244244 3545 244260
rect 3607 245036 3641 245052
rect 3607 244244 3641 244260
rect 3721 245036 3755 245052
rect 3721 244244 3755 244260
rect 3817 245036 3851 245052
rect 3817 244244 3851 244260
rect 3931 245036 3965 245052
rect 3931 244244 3965 244260
rect 4027 245036 4061 245052
rect 4027 244244 4061 244260
rect 4141 245036 4175 245052
rect 4141 244244 4175 244260
rect 4237 245036 4271 245052
rect 4237 244244 4271 244260
rect 4351 245036 4385 245052
rect 4351 244244 4385 244260
rect 4447 245036 4481 245052
rect 4447 244244 4481 244260
rect 4561 245036 4595 245052
rect 4561 244244 4595 244260
rect 4657 245036 4691 245052
rect 4657 244244 4691 244260
rect 4771 245036 4805 245052
rect 4771 244244 4805 244260
rect 4867 245036 4901 245052
rect 4867 244244 4901 244260
rect 4981 245036 5015 245052
rect 4981 244244 5015 244260
rect 5077 245036 5111 245052
rect 5077 244244 5111 244260
rect 5191 245036 5225 245052
rect 5191 244244 5225 244260
rect 5287 245036 5321 245052
rect 5287 244244 5321 244260
rect 5401 245036 5435 245052
rect 5401 244244 5435 244260
rect 5497 245036 5531 245052
rect 5497 244244 5531 244260
rect 5611 245036 5645 245052
rect 5611 244244 5645 244260
rect 5707 245036 5741 245052
rect 5707 244244 5741 244260
rect 5821 245036 5855 245052
rect 5821 244244 5855 244260
rect 5917 245036 5951 245052
rect 5917 244244 5951 244260
rect 6031 245036 6065 245052
rect 6031 244244 6065 244260
rect 6127 245036 6161 245052
rect 6127 244244 6161 244260
rect 6241 245036 6275 245052
rect 6241 244244 6275 244260
rect 6337 245036 6371 245052
rect 6337 244244 6371 244260
rect 6451 245036 6485 245052
rect 6451 244244 6485 244260
rect 6547 245036 6581 245052
rect 6547 244244 6581 244260
rect 6661 245036 6695 245052
rect 6661 244244 6695 244260
rect 6757 245036 6791 245052
rect 6757 244244 6791 244260
rect 6871 245036 6905 245052
rect 6871 244244 6905 244260
rect 6967 245036 7001 245052
rect 6967 244244 7001 244260
rect 7081 245036 7115 245052
rect 7081 244244 7115 244260
rect 7177 245036 7211 245052
rect 7177 244244 7211 244260
rect 7291 245036 7325 245052
rect 7291 244244 7325 244260
rect 7387 245036 7421 245052
rect 7387 244244 7421 244260
rect 7501 245036 7535 245052
rect 7501 244244 7535 244260
rect 7597 245036 7631 245052
rect 7597 244244 7631 244260
rect 7711 245036 7745 245052
rect 7711 244244 7745 244260
rect 7807 245036 7841 245052
rect 7807 244244 7841 244260
rect 7921 245036 7955 245052
rect 7921 244244 7955 244260
rect 8017 245036 8051 245052
rect 8017 244244 8051 244260
rect 8131 245036 8165 245052
rect 8131 244244 8165 244260
rect 8227 245036 8261 245052
rect 8227 244244 8261 244260
rect 8341 245036 8375 245052
rect 8341 244244 8375 244260
rect 8437 245036 8471 245052
rect 8437 244244 8471 244260
rect 8551 245036 8585 245052
rect 8551 244244 8585 244260
rect 8647 245036 8681 245052
rect 8647 244244 8681 244260
rect 8761 245036 8795 245052
rect 8761 244244 8795 244260
rect 8857 245036 8891 245052
rect 8857 244244 8891 244260
rect 8971 245036 9005 245052
rect 8971 244244 9005 244260
rect 9067 245036 9101 245052
rect 9067 244244 9101 244260
rect 9181 245036 9215 245052
rect 9181 244244 9215 244260
rect 9277 245036 9311 245052
rect 9277 244244 9311 244260
rect 9391 245036 9425 245052
rect 9391 244244 9425 244260
rect 9487 245036 9521 245052
rect 9487 244244 9521 244260
rect 9601 245036 9635 245052
rect 9601 244244 9635 244260
rect 9697 245036 9731 245052
rect 9697 244244 9731 244260
rect 9811 245036 9845 245052
rect 9811 244244 9845 244260
rect 9907 245036 9941 245052
rect 9907 244244 9941 244260
rect 10021 245036 10055 245052
rect 10021 244244 10055 244260
rect 10117 245036 10151 245052
rect 10117 244244 10151 244260
rect 10231 245036 10265 245052
rect 10231 244244 10265 244260
rect 10327 245036 10361 245052
rect 10327 244244 10361 244260
rect 10441 245036 10475 245052
rect 10441 244244 10475 244260
rect 10537 245036 10571 245052
rect 10537 244244 10571 244260
rect 10651 245036 10685 245052
rect 10651 244244 10685 244260
rect 10747 245036 10781 245052
rect 10747 244244 10781 244260
rect 10861 245036 10895 245052
rect 10861 244244 10895 244260
rect 10957 245036 10991 245052
rect 10957 244244 10991 244260
rect 11071 245036 11105 245052
rect 11071 244244 11105 244260
rect 11167 245036 11201 245052
rect 11167 244244 11201 244260
rect 11281 245036 11315 245052
rect 11281 244244 11315 244260
rect 11377 245036 11411 245052
rect 11377 244244 11411 244260
rect 11491 245036 11525 245052
rect 11491 244244 11525 244260
rect 11587 245036 11621 245052
rect 11587 244244 11621 244260
rect 11701 245036 11735 245052
rect 11701 244244 11735 244260
rect 11797 245036 11831 245052
rect 11797 244244 11831 244260
rect 11911 245036 11945 245052
rect 11911 244244 11945 244260
rect 12007 245036 12041 245052
rect 12007 244244 12041 244260
rect 12121 245036 12155 245052
rect 12121 244244 12155 244260
rect 12217 245036 12251 245052
rect 12217 244244 12251 244260
rect 12331 245036 12365 245052
rect 12331 244244 12365 244260
rect 12427 245036 12461 245052
rect 12427 244244 12461 244260
rect 12541 245036 12575 245052
rect 12541 244244 12575 244260
rect 12637 245036 12671 245052
rect 12637 244244 12671 244260
rect 12751 245036 12785 245052
rect 12751 244244 12785 244260
rect 12847 245036 12881 245052
rect 12847 244244 12881 244260
rect 12961 245036 12995 245052
rect 12961 244244 12995 244260
rect 13057 245036 13091 245052
rect 13057 244244 13091 244260
rect 13171 245036 13205 245052
rect 13171 244244 13205 244260
rect 13267 245036 13301 245052
rect 13267 244244 13301 244260
rect 13381 245036 13415 245052
rect 13381 244244 13415 244260
rect 13477 245036 13511 245052
rect 13477 244244 13511 244260
rect 13591 245036 13625 245052
rect 13591 244244 13625 244260
rect 13687 245036 13721 245052
rect 13687 244244 13721 244260
rect 13801 245036 13835 245052
rect 13801 244244 13835 244260
rect 13897 245036 13931 245052
rect 13897 244244 13931 244260
rect 14011 245036 14045 245052
rect 14011 244244 14045 244260
rect 14107 245036 14141 245052
rect 14107 244244 14141 244260
rect 14221 245036 14255 245052
rect 14221 244244 14255 244260
rect 14317 245036 14351 245052
rect 14317 244244 14351 244260
rect 14431 245036 14465 245052
rect 14431 244244 14465 244260
rect 14527 245036 14561 245052
rect 14527 244244 14561 244260
rect 14641 245036 14675 245052
rect 14641 244244 14675 244260
rect 14737 245036 14771 245052
rect 14737 244244 14771 244260
rect 14851 245036 14885 245052
rect 14851 244244 14885 244260
rect 14947 245036 14981 245052
rect 14947 244244 14981 244260
rect 15061 245036 15095 245052
rect 15061 244244 15095 244260
rect 15157 245036 15191 245052
rect 15157 244244 15191 244260
rect 15271 245036 15305 245052
rect 15271 244244 15305 244260
rect 15367 245036 15401 245052
rect 15367 244244 15401 244260
rect 15481 245036 15515 245052
rect 15481 244244 15515 244260
rect 15577 245036 15611 245052
rect 15577 244244 15611 244260
rect 15691 245036 15725 245052
rect 15691 244244 15725 244260
rect 15787 245036 15821 245052
rect 15787 244244 15821 244260
rect 15901 245036 15935 245052
rect 15901 244244 15935 244260
rect 15997 245036 16031 245052
rect 15997 244244 16031 244260
rect 16111 245036 16145 245052
rect 16111 244244 16145 244260
rect 16207 245036 16241 245052
rect 16207 244244 16241 244260
rect 16321 245036 16355 245052
rect 16321 244244 16355 244260
rect 16417 245036 16451 245052
rect 16417 244244 16451 244260
rect 16531 245036 16565 245052
rect 16531 244244 16565 244260
rect 16627 245036 16661 245052
rect 16627 244244 16661 244260
rect 16741 245036 16775 245052
rect 16741 244244 16775 244260
rect 16837 245036 16871 245052
rect 16837 244244 16871 244260
rect 16951 245036 16985 245052
rect 16951 244244 16985 244260
rect 17047 245036 17081 245052
rect 17047 244244 17081 244260
rect 17161 245036 17195 245052
rect 17161 244244 17195 244260
rect 17257 245036 17291 245052
rect 17257 244244 17291 244260
rect 17371 245036 17405 245052
rect 17371 244244 17405 244260
rect 17467 245036 17501 245052
rect 17467 244244 17501 244260
rect 17581 245036 17615 245052
rect 17581 244244 17615 244260
rect 17677 245036 17711 245052
rect 17677 244244 17711 244260
rect 17791 245036 17825 245052
rect 17791 244244 17825 244260
rect 17887 245036 17921 245052
rect 17887 244244 17921 244260
rect 18001 245036 18035 245052
rect 18001 244244 18035 244260
rect 18097 245036 18131 245052
rect 18097 244244 18131 244260
rect 18211 245036 18245 245052
rect 18211 244244 18245 244260
rect 18307 245036 18341 245052
rect 18307 244244 18341 244260
rect 18421 245036 18455 245052
rect 18421 244244 18455 244260
rect 18517 245036 18551 245052
rect 18517 244244 18551 244260
rect 18631 245036 18665 245052
rect 18631 244244 18665 244260
rect 18727 245036 18761 245052
rect 18727 244244 18761 244260
rect 18841 245036 18875 245052
rect 18841 244244 18875 244260
rect 18937 245036 18971 245052
rect 18937 244244 18971 244260
rect 19051 245036 19085 245052
rect 19051 244244 19085 244260
rect 19147 245036 19181 245052
rect 19147 244244 19181 244260
rect 19261 245036 19295 245052
rect 19261 244244 19295 244260
rect 19357 245036 19391 245052
rect 19357 244244 19391 244260
rect 19471 245036 19505 245052
rect 19471 244244 19505 244260
rect 19567 245036 19601 245052
rect 19567 244244 19601 244260
rect 19681 245036 19715 245052
rect 19681 244244 19715 244260
rect 19777 245036 19811 245052
rect 19777 244244 19811 244260
rect 19891 245036 19925 245052
rect 19891 244244 19925 244260
rect 19987 245036 20021 245052
rect 19987 244244 20021 244260
rect 20101 245036 20135 245052
rect 20101 244244 20135 244260
rect 20197 245036 20231 245052
rect 20197 244244 20231 244260
rect 20311 245036 20345 245052
rect 20311 244244 20345 244260
rect 20407 245036 20441 245052
rect 20407 244244 20441 244260
rect 20521 245036 20555 245052
rect 20521 244244 20555 244260
rect 20617 245036 20651 245052
rect 20617 244244 20651 244260
rect 20731 245036 20765 245052
rect 20731 244244 20765 244260
rect 20827 245036 20861 245052
rect 20827 244244 20861 244260
rect 20941 245036 20975 245052
rect 20941 244244 20975 244260
rect 21037 245036 21071 245052
rect 21037 244244 21071 244260
rect 21151 245036 21185 245052
rect 21151 244244 21185 244260
rect 21247 245036 21281 245052
rect 21247 244244 21281 244260
rect 21361 245036 21395 245052
rect 21361 244244 21395 244260
rect 21457 245036 21491 245052
rect 21457 244244 21491 244260
rect 21571 245036 21605 245052
rect 21571 244244 21605 244260
rect 21667 245036 21701 245052
rect 21667 244244 21701 244260
rect 21781 245036 21815 245052
rect 21781 244244 21815 244260
rect 21877 245036 21911 245052
rect 21877 244244 21911 244260
rect 21991 245036 22025 245052
rect 21991 244244 22025 244260
rect 22087 245036 22121 245052
rect 22087 244244 22121 244260
rect 22201 245036 22235 245052
rect 22201 244244 22235 244260
rect 22297 245036 22331 245052
rect 22297 244244 22331 244260
rect 22411 245036 22445 245052
rect 22411 244244 22445 244260
rect 22507 245036 22541 245052
rect 22507 244244 22541 244260
rect 22621 245036 22655 245052
rect 22621 244244 22655 244260
rect 22717 245036 22751 245052
rect 22717 244244 22751 244260
rect 22831 245036 22865 245052
rect 22831 244244 22865 244260
rect 22927 245036 22961 245052
rect 22927 244244 22961 244260
rect 23041 245036 23075 245052
rect 23041 244244 23075 244260
rect 23137 245036 23171 245052
rect 23137 244244 23171 244260
rect 23251 245036 23285 245052
rect 23251 244244 23285 244260
rect 23347 245036 23381 245052
rect 23347 244244 23381 244260
rect 23461 245036 23495 245052
rect 23461 244244 23495 244260
rect 23557 245036 23591 245052
rect 23557 244244 23591 244260
rect 23671 245036 23705 245052
rect 23671 244244 23705 244260
rect 23767 245036 23801 245052
rect 23767 244244 23801 244260
rect 23881 245036 23915 245052
rect 23881 244244 23915 244260
rect 23977 245036 24011 245052
rect 23977 244244 24011 244260
rect 24091 245036 24125 245052
rect 24091 244244 24125 244260
rect 24187 245036 24221 245052
rect 24187 244244 24221 244260
rect 24301 245036 24335 245052
rect 24301 244244 24335 244260
rect 24397 245036 24431 245052
rect 24397 244244 24431 244260
rect 24511 245036 24545 245052
rect 24511 244244 24545 244260
rect 24607 245036 24641 245052
rect 24607 244244 24641 244260
rect 24721 245036 24755 245052
rect 24721 244244 24755 244260
rect 24817 245036 24851 245052
rect 24817 244244 24851 244260
rect 24931 245036 24965 245052
rect 24931 244244 24965 244260
rect 25027 245036 25061 245052
rect 25027 244244 25061 244260
rect 25141 245036 25175 245052
rect 25141 244244 25175 244260
rect 25237 245036 25271 245052
rect 25237 244244 25271 244260
rect 25351 245036 25385 245052
rect 25351 244244 25385 244260
rect 25447 245036 25481 245052
rect 25447 244244 25481 244260
rect 25561 245036 25595 245052
rect 25561 244244 25595 244260
rect 25657 245036 25691 245052
rect 25657 244244 25691 244260
rect 25771 245036 25805 245052
rect 25771 244244 25805 244260
rect 25867 245036 25901 245052
rect 25867 244244 25901 244260
rect 25981 245036 26015 245052
rect 25981 244244 26015 244260
rect 26077 245036 26111 245052
rect 26077 244244 26111 244260
rect 26191 245036 26225 245052
rect 26191 244244 26225 244260
rect 26287 245036 26321 245052
rect 26287 244244 26321 244260
rect 26401 245036 26435 245052
rect 26401 244244 26435 244260
rect 26497 245036 26531 245052
rect 26497 244244 26531 244260
rect 26611 245036 26645 245052
rect 26611 244244 26645 244260
rect 26707 245036 26741 245052
rect 26707 244244 26741 244260
rect 26821 245036 26855 245052
rect 26821 244244 26855 244260
rect 26917 245036 26951 245052
rect 26917 244244 26951 244260
rect 27031 245036 27065 245052
rect 27031 244244 27065 244260
rect 27127 245036 27161 245052
rect 27127 244244 27161 244260
rect 27241 245036 27275 245052
rect 27241 244244 27275 244260
rect 27337 245036 27371 245052
rect 27337 244244 27371 244260
rect -3807 244167 -3791 244201
rect -3695 244167 -3679 244201
rect -3387 244167 -3371 244201
rect -3275 244167 -3259 244201
rect -2967 244167 -2951 244201
rect -2855 244167 -2839 244201
rect -2547 244167 -2531 244201
rect -2435 244167 -2419 244201
rect -2127 244167 -2111 244201
rect -2015 244167 -1999 244201
rect -1707 244167 -1691 244201
rect -1595 244167 -1579 244201
rect -1287 244167 -1271 244201
rect -1175 244167 -1159 244201
rect -867 244167 -851 244201
rect -755 244167 -739 244201
rect -447 244167 -431 244201
rect -335 244167 -319 244201
rect -27 244167 -11 244201
rect 85 244167 101 244201
rect 393 244167 409 244201
rect 505 244167 521 244201
rect 813 244167 829 244201
rect 925 244167 941 244201
rect 1233 244167 1249 244201
rect 1345 244167 1361 244201
rect 1653 244167 1669 244201
rect 1765 244167 1781 244201
rect 2073 244167 2089 244201
rect 2185 244167 2201 244201
rect 2493 244167 2509 244201
rect 2605 244167 2621 244201
rect 2913 244167 2929 244201
rect 3025 244167 3041 244201
rect 3333 244167 3349 244201
rect 3445 244167 3461 244201
rect 3753 244167 3769 244201
rect 3865 244167 3881 244201
rect 4173 244167 4189 244201
rect 4285 244167 4301 244201
rect 4593 244167 4609 244201
rect 4705 244167 4721 244201
rect 5013 244167 5029 244201
rect 5125 244167 5141 244201
rect 5433 244167 5449 244201
rect 5545 244167 5561 244201
rect 5853 244167 5869 244201
rect 5965 244167 5981 244201
rect 6273 244167 6289 244201
rect 6385 244167 6401 244201
rect 6693 244167 6709 244201
rect 6805 244167 6821 244201
rect 7113 244167 7129 244201
rect 7225 244167 7241 244201
rect 7533 244167 7549 244201
rect 7645 244167 7661 244201
rect 7953 244167 7969 244201
rect 8065 244167 8081 244201
rect 8373 244167 8389 244201
rect 8485 244167 8501 244201
rect 8793 244167 8809 244201
rect 8905 244167 8921 244201
rect 9213 244167 9229 244201
rect 9325 244167 9341 244201
rect 9633 244167 9649 244201
rect 9745 244167 9761 244201
rect 10053 244167 10069 244201
rect 10165 244167 10181 244201
rect 10473 244167 10489 244201
rect 10585 244167 10601 244201
rect 10893 244167 10909 244201
rect 11005 244167 11021 244201
rect 11313 244167 11329 244201
rect 11425 244167 11441 244201
rect 11733 244167 11749 244201
rect 11845 244167 11861 244201
rect 12153 244167 12169 244201
rect 12265 244167 12281 244201
rect 12573 244167 12589 244201
rect 12685 244167 12701 244201
rect 12993 244167 13009 244201
rect 13105 244167 13121 244201
rect 13413 244167 13429 244201
rect 13525 244167 13541 244201
rect 13833 244167 13849 244201
rect 13945 244167 13961 244201
rect 14253 244167 14269 244201
rect 14365 244167 14381 244201
rect 14673 244167 14689 244201
rect 14785 244167 14801 244201
rect 15093 244167 15109 244201
rect 15205 244167 15221 244201
rect 15513 244167 15529 244201
rect 15625 244167 15641 244201
rect 15933 244167 15949 244201
rect 16045 244167 16061 244201
rect 16353 244167 16369 244201
rect 16465 244167 16481 244201
rect 16773 244167 16789 244201
rect 16885 244167 16901 244201
rect 17193 244167 17209 244201
rect 17305 244167 17321 244201
rect 17613 244167 17629 244201
rect 17725 244167 17741 244201
rect 18033 244167 18049 244201
rect 18145 244167 18161 244201
rect 18453 244167 18469 244201
rect 18565 244167 18581 244201
rect 18873 244167 18889 244201
rect 18985 244167 19001 244201
rect 19293 244167 19309 244201
rect 19405 244167 19421 244201
rect 19713 244167 19729 244201
rect 19825 244167 19841 244201
rect 20133 244167 20149 244201
rect 20245 244167 20261 244201
rect 20553 244167 20569 244201
rect 20665 244167 20681 244201
rect 20973 244167 20989 244201
rect 21085 244167 21101 244201
rect 21393 244167 21409 244201
rect 21505 244167 21521 244201
rect 21813 244167 21829 244201
rect 21925 244167 21941 244201
rect 22233 244167 22249 244201
rect 22345 244167 22361 244201
rect 22653 244167 22669 244201
rect 22765 244167 22781 244201
rect 23073 244167 23089 244201
rect 23185 244167 23201 244201
rect 23493 244167 23509 244201
rect 23605 244167 23621 244201
rect 23913 244167 23929 244201
rect 24025 244167 24041 244201
rect 24333 244167 24349 244201
rect 24445 244167 24461 244201
rect 24753 244167 24769 244201
rect 24865 244167 24881 244201
rect 25173 244167 25189 244201
rect 25285 244167 25301 244201
rect 25593 244167 25609 244201
rect 25705 244167 25721 244201
rect 26013 244167 26029 244201
rect 26125 244167 26141 244201
rect 26433 244167 26449 244201
rect 26545 244167 26561 244201
rect 26853 244167 26869 244201
rect 26965 244167 26981 244201
rect 27273 244167 27289 244201
rect 27385 244167 27401 244201
rect -4163 244099 -4129 244161
rect 27451 244099 27485 244161
rect -4163 244065 -4067 244099
rect 27389 244065 27485 244099
<< viali >>
rect -4163 264212 27486 264317
rect -4001 264076 -3905 264110
rect -3581 264076 -3485 264110
rect -3161 264076 -3065 264110
rect -2741 264076 -2645 264110
rect -2321 264076 -2225 264110
rect -1901 264076 -1805 264110
rect -1481 264076 -1385 264110
rect -1061 264076 -965 264110
rect -641 264076 -545 264110
rect -221 264076 -125 264110
rect 199 264076 295 264110
rect 619 264076 715 264110
rect 1039 264076 1135 264110
rect 1459 264076 1555 264110
rect 1879 264076 1975 264110
rect 2299 264076 2395 264110
rect 2719 264076 2815 264110
rect 3139 264076 3235 264110
rect 3559 264076 3655 264110
rect 3979 264076 4075 264110
rect 4399 264076 4495 264110
rect 4819 264076 4915 264110
rect 5239 264076 5335 264110
rect 5659 264076 5755 264110
rect 6079 264076 6175 264110
rect 6499 264076 6595 264110
rect 6919 264076 7015 264110
rect 7339 264076 7435 264110
rect 7759 264076 7855 264110
rect 8179 264076 8275 264110
rect 8599 264076 8695 264110
rect 9019 264076 9115 264110
rect 9439 264076 9535 264110
rect 9859 264076 9955 264110
rect 10279 264076 10375 264110
rect 10699 264076 10795 264110
rect 11119 264076 11215 264110
rect 11539 264076 11635 264110
rect 11959 264076 12055 264110
rect 12379 264076 12475 264110
rect 12799 264076 12895 264110
rect 13219 264076 13315 264110
rect 13639 264076 13735 264110
rect 14059 264076 14155 264110
rect 14479 264076 14575 264110
rect 14899 264076 14995 264110
rect 15319 264076 15415 264110
rect 15739 264076 15835 264110
rect 16159 264076 16255 264110
rect 16579 264076 16675 264110
rect 16999 264076 17095 264110
rect 17419 264076 17515 264110
rect 17839 264076 17935 264110
rect 18259 264076 18355 264110
rect 18679 264076 18775 264110
rect 19099 264076 19195 264110
rect 19519 264076 19615 264110
rect 19939 264076 20035 264110
rect 20359 264076 20455 264110
rect 20779 264076 20875 264110
rect 21199 264076 21295 264110
rect 21619 264076 21715 264110
rect 22039 264076 22135 264110
rect 22459 264076 22555 264110
rect 22879 264076 22975 264110
rect 23299 264076 23395 264110
rect 23719 264076 23815 264110
rect 24139 264076 24235 264110
rect 24559 264076 24655 264110
rect 24979 264076 25075 264110
rect 25399 264076 25495 264110
rect 25819 264076 25915 264110
rect 26239 264076 26335 264110
rect 26659 264076 26755 264110
rect 27079 264076 27175 264110
rect -4049 263250 -4015 264026
rect -3953 263250 -3919 264026
rect -3839 263250 -3805 264026
rect -3743 263250 -3709 264026
rect -3629 263250 -3595 264026
rect -3533 263250 -3499 264026
rect -3419 263250 -3385 264026
rect -3323 263250 -3289 264026
rect -3209 263250 -3175 264026
rect -3113 263250 -3079 264026
rect -2999 263250 -2965 264026
rect -2903 263250 -2869 264026
rect -2789 263250 -2755 264026
rect -2693 263250 -2659 264026
rect -2579 263250 -2545 264026
rect -2483 263250 -2449 264026
rect -2369 263250 -2335 264026
rect -2273 263250 -2239 264026
rect -2159 263250 -2125 264026
rect -2063 263250 -2029 264026
rect -1949 263250 -1915 264026
rect -1853 263250 -1819 264026
rect -1739 263250 -1705 264026
rect -1643 263250 -1609 264026
rect -1529 263250 -1495 264026
rect -1433 263250 -1399 264026
rect -1319 263250 -1285 264026
rect -1223 263250 -1189 264026
rect -1109 263250 -1075 264026
rect -1013 263250 -979 264026
rect -899 263250 -865 264026
rect -803 263250 -769 264026
rect -689 263250 -655 264026
rect -593 263250 -559 264026
rect -479 263250 -445 264026
rect -383 263250 -349 264026
rect -269 263250 -235 264026
rect -173 263250 -139 264026
rect -59 263250 -25 264026
rect 37 263250 71 264026
rect 151 263250 185 264026
rect 247 263250 281 264026
rect 361 263250 395 264026
rect 457 263250 491 264026
rect 571 263250 605 264026
rect 667 263250 701 264026
rect 781 263250 815 264026
rect 877 263250 911 264026
rect 991 263250 1025 264026
rect 1087 263250 1121 264026
rect 1201 263250 1235 264026
rect 1297 263250 1331 264026
rect 1411 263250 1445 264026
rect 1507 263250 1541 264026
rect 1621 263250 1655 264026
rect 1717 263250 1751 264026
rect 1831 263250 1865 264026
rect 1927 263250 1961 264026
rect 2041 263250 2075 264026
rect 2137 263250 2171 264026
rect 2251 263250 2285 264026
rect 2347 263250 2381 264026
rect 2461 263250 2495 264026
rect 2557 263250 2591 264026
rect 2671 263250 2705 264026
rect 2767 263250 2801 264026
rect 2881 263250 2915 264026
rect 2977 263250 3011 264026
rect 3091 263250 3125 264026
rect 3187 263250 3221 264026
rect 3301 263250 3335 264026
rect 3397 263250 3431 264026
rect 3511 263250 3545 264026
rect 3607 263250 3641 264026
rect 3721 263250 3755 264026
rect 3817 263250 3851 264026
rect 3931 263250 3965 264026
rect 4027 263250 4061 264026
rect 4141 263250 4175 264026
rect 4237 263250 4271 264026
rect 4351 263250 4385 264026
rect 4447 263250 4481 264026
rect 4561 263250 4595 264026
rect 4657 263250 4691 264026
rect 4771 263250 4805 264026
rect 4867 263250 4901 264026
rect 4981 263250 5015 264026
rect 5077 263250 5111 264026
rect 5191 263250 5225 264026
rect 5287 263250 5321 264026
rect 5401 263250 5435 264026
rect 5497 263250 5531 264026
rect 5611 263250 5645 264026
rect 5707 263250 5741 264026
rect 5821 263250 5855 264026
rect 5917 263250 5951 264026
rect 6031 263250 6065 264026
rect 6127 263250 6161 264026
rect 6241 263250 6275 264026
rect 6337 263250 6371 264026
rect 6451 263250 6485 264026
rect 6547 263250 6581 264026
rect 6661 263250 6695 264026
rect 6757 263250 6791 264026
rect 6871 263250 6905 264026
rect 6967 263250 7001 264026
rect 7081 263250 7115 264026
rect 7177 263250 7211 264026
rect 7291 263250 7325 264026
rect 7387 263250 7421 264026
rect 7501 263250 7535 264026
rect 7597 263250 7631 264026
rect 7711 263250 7745 264026
rect 7807 263250 7841 264026
rect 7921 263250 7955 264026
rect 8017 263250 8051 264026
rect 8131 263250 8165 264026
rect 8227 263250 8261 264026
rect 8341 263250 8375 264026
rect 8437 263250 8471 264026
rect 8551 263250 8585 264026
rect 8647 263250 8681 264026
rect 8761 263250 8795 264026
rect 8857 263250 8891 264026
rect 8971 263250 9005 264026
rect 9067 263250 9101 264026
rect 9181 263250 9215 264026
rect 9277 263250 9311 264026
rect 9391 263250 9425 264026
rect 9487 263250 9521 264026
rect 9601 263250 9635 264026
rect 9697 263250 9731 264026
rect 9811 263250 9845 264026
rect 9907 263250 9941 264026
rect 10021 263250 10055 264026
rect 10117 263250 10151 264026
rect 10231 263250 10265 264026
rect 10327 263250 10361 264026
rect 10441 263250 10475 264026
rect 10537 263250 10571 264026
rect 10651 263250 10685 264026
rect 10747 263250 10781 264026
rect 10861 263250 10895 264026
rect 10957 263250 10991 264026
rect 11071 263250 11105 264026
rect 11167 263250 11201 264026
rect 11281 263250 11315 264026
rect 11377 263250 11411 264026
rect 11491 263250 11525 264026
rect 11587 263250 11621 264026
rect 11701 263250 11735 264026
rect 11797 263250 11831 264026
rect 11911 263250 11945 264026
rect 12007 263250 12041 264026
rect 12121 263250 12155 264026
rect 12217 263250 12251 264026
rect 12331 263250 12365 264026
rect 12427 263250 12461 264026
rect 12541 263250 12575 264026
rect 12637 263250 12671 264026
rect 12751 263250 12785 264026
rect 12847 263250 12881 264026
rect 12961 263250 12995 264026
rect 13057 263250 13091 264026
rect 13171 263250 13205 264026
rect 13267 263250 13301 264026
rect 13381 263250 13415 264026
rect 13477 263250 13511 264026
rect 13591 263250 13625 264026
rect 13687 263250 13721 264026
rect 13801 263250 13835 264026
rect 13897 263250 13931 264026
rect 14011 263250 14045 264026
rect 14107 263250 14141 264026
rect 14221 263250 14255 264026
rect 14317 263250 14351 264026
rect 14431 263250 14465 264026
rect 14527 263250 14561 264026
rect 14641 263250 14675 264026
rect 14737 263250 14771 264026
rect 14851 263250 14885 264026
rect 14947 263250 14981 264026
rect 15061 263250 15095 264026
rect 15157 263250 15191 264026
rect 15271 263250 15305 264026
rect 15367 263250 15401 264026
rect 15481 263250 15515 264026
rect 15577 263250 15611 264026
rect 15691 263250 15725 264026
rect 15787 263250 15821 264026
rect 15901 263250 15935 264026
rect 15997 263250 16031 264026
rect 16111 263250 16145 264026
rect 16207 263250 16241 264026
rect 16321 263250 16355 264026
rect 16417 263250 16451 264026
rect 16531 263250 16565 264026
rect 16627 263250 16661 264026
rect 16741 263250 16775 264026
rect 16837 263250 16871 264026
rect 16951 263250 16985 264026
rect 17047 263250 17081 264026
rect 17161 263250 17195 264026
rect 17257 263250 17291 264026
rect 17371 263250 17405 264026
rect 17467 263250 17501 264026
rect 17581 263250 17615 264026
rect 17677 263250 17711 264026
rect 17791 263250 17825 264026
rect 17887 263250 17921 264026
rect 18001 263250 18035 264026
rect 18097 263250 18131 264026
rect 18211 263250 18245 264026
rect 18307 263250 18341 264026
rect 18421 263250 18455 264026
rect 18517 263250 18551 264026
rect 18631 263250 18665 264026
rect 18727 263250 18761 264026
rect 18841 263250 18875 264026
rect 18937 263250 18971 264026
rect 19051 263250 19085 264026
rect 19147 263250 19181 264026
rect 19261 263250 19295 264026
rect 19357 263250 19391 264026
rect 19471 263250 19505 264026
rect 19567 263250 19601 264026
rect 19681 263250 19715 264026
rect 19777 263250 19811 264026
rect 19891 263250 19925 264026
rect 19987 263250 20021 264026
rect 20101 263250 20135 264026
rect 20197 263250 20231 264026
rect 20311 263250 20345 264026
rect 20407 263250 20441 264026
rect 20521 263250 20555 264026
rect 20617 263250 20651 264026
rect 20731 263250 20765 264026
rect 20827 263250 20861 264026
rect 20941 263250 20975 264026
rect 21037 263250 21071 264026
rect 21151 263250 21185 264026
rect 21247 263250 21281 264026
rect 21361 263250 21395 264026
rect 21457 263250 21491 264026
rect 21571 263250 21605 264026
rect 21667 263250 21701 264026
rect 21781 263250 21815 264026
rect 21877 263250 21911 264026
rect 21991 263250 22025 264026
rect 22087 263250 22121 264026
rect 22201 263250 22235 264026
rect 22297 263250 22331 264026
rect 22411 263250 22445 264026
rect 22507 263250 22541 264026
rect 22621 263250 22655 264026
rect 22717 263250 22751 264026
rect 22831 263250 22865 264026
rect 22927 263250 22961 264026
rect 23041 263250 23075 264026
rect 23137 263250 23171 264026
rect 23251 263250 23285 264026
rect 23347 263250 23381 264026
rect 23461 263250 23495 264026
rect 23557 263250 23591 264026
rect 23671 263250 23705 264026
rect 23767 263250 23801 264026
rect 23881 263250 23915 264026
rect 23977 263250 24011 264026
rect 24091 263250 24125 264026
rect 24187 263250 24221 264026
rect 24301 263250 24335 264026
rect 24397 263250 24431 264026
rect 24511 263250 24545 264026
rect 24607 263250 24641 264026
rect 24721 263250 24755 264026
rect 24817 263250 24851 264026
rect 24931 263250 24965 264026
rect 25027 263250 25061 264026
rect 25141 263250 25175 264026
rect 25237 263250 25271 264026
rect 25351 263250 25385 264026
rect 25447 263250 25481 264026
rect 25561 263250 25595 264026
rect 25657 263250 25691 264026
rect 25771 263250 25805 264026
rect 25867 263250 25901 264026
rect 25981 263250 26015 264026
rect 26077 263250 26111 264026
rect 26191 263250 26225 264026
rect 26287 263250 26321 264026
rect 26401 263250 26435 264026
rect 26497 263250 26531 264026
rect 26611 263250 26645 264026
rect 26707 263250 26741 264026
rect 26821 263250 26855 264026
rect 26917 263250 26951 264026
rect 27031 263250 27065 264026
rect 27127 263250 27161 264026
rect 27241 263250 27275 264026
rect 27337 263250 27371 264026
rect -3791 263164 -3757 263198
rect -3371 263164 -3337 263198
rect -2951 263164 -2917 263198
rect -2531 263164 -2497 263198
rect -2111 263164 -2077 263198
rect -1691 263164 -1657 263198
rect -1271 263164 -1237 263198
rect -851 263164 -817 263198
rect -431 263164 -397 263198
rect -11 263164 23 263198
rect 409 263164 443 263198
rect 829 263164 863 263198
rect 1249 263164 1283 263198
rect 1669 263164 1703 263198
rect 2089 263164 2123 263198
rect 2509 263164 2543 263198
rect 2929 263164 2963 263198
rect 3349 263164 3383 263198
rect 3769 263164 3803 263198
rect 4189 263164 4223 263198
rect 4609 263164 4643 263198
rect 5029 263164 5063 263198
rect 5449 263164 5483 263198
rect 5869 263164 5903 263198
rect 6289 263164 6323 263198
rect 6709 263164 6743 263198
rect 7129 263164 7163 263198
rect 7549 263164 7583 263198
rect 7969 263164 8003 263198
rect 8389 263164 8423 263198
rect 8809 263164 8843 263198
rect 9229 263164 9263 263198
rect 9649 263164 9683 263198
rect 10069 263164 10103 263198
rect 10489 263164 10523 263198
rect 10909 263164 10943 263198
rect 11329 263164 11363 263198
rect 11749 263164 11783 263198
rect 12169 263164 12203 263198
rect 12589 263164 12623 263198
rect 13009 263164 13043 263198
rect 13429 263164 13463 263198
rect 13849 263164 13883 263198
rect 14269 263164 14303 263198
rect 14689 263164 14723 263198
rect 15109 263164 15143 263198
rect 15529 263164 15563 263198
rect 15949 263164 15983 263198
rect 16369 263164 16403 263198
rect 16789 263164 16823 263198
rect 17209 263164 17243 263198
rect 17629 263164 17663 263198
rect 18049 263164 18083 263198
rect 18469 263164 18503 263198
rect 18889 263164 18923 263198
rect 19309 263164 19343 263198
rect 19729 263164 19763 263198
rect 20149 263164 20183 263198
rect 20569 263164 20603 263198
rect 20989 263164 21023 263198
rect 21409 263164 21443 263198
rect 21829 263164 21863 263198
rect 22249 263164 22283 263198
rect 22669 263164 22703 263198
rect 23089 263164 23123 263198
rect 23509 263164 23543 263198
rect 23929 263164 23963 263198
rect 24349 263164 24383 263198
rect 24769 263164 24803 263198
rect 25189 263164 25223 263198
rect 25609 263164 25643 263198
rect 26029 263164 26063 263198
rect 26449 263164 26483 263198
rect 26869 263164 26903 263198
rect 27289 263164 27323 263198
rect -3791 263090 -3757 263164
rect -3371 263090 -3337 263164
rect -2951 263090 -2917 263164
rect -2531 263090 -2497 263164
rect -2111 263090 -2077 263164
rect -1691 263090 -1657 263164
rect -1271 263090 -1237 263164
rect -851 263090 -817 263164
rect -431 263090 -397 263164
rect -11 263090 23 263164
rect 409 263090 443 263164
rect 829 263090 863 263164
rect 1249 263090 1283 263164
rect 1669 263090 1703 263164
rect 2089 263090 2123 263164
rect 2509 263090 2543 263164
rect 2929 263090 2963 263164
rect 3349 263090 3383 263164
rect 3769 263090 3803 263164
rect 4189 263090 4223 263164
rect 4609 263090 4643 263164
rect 5029 263090 5063 263164
rect 5449 263090 5483 263164
rect 5869 263090 5903 263164
rect 6289 263090 6323 263164
rect 6709 263090 6743 263164
rect 7129 263090 7163 263164
rect 7549 263090 7583 263164
rect 7969 263090 8003 263164
rect 8389 263090 8423 263164
rect 8809 263090 8843 263164
rect 9229 263090 9263 263164
rect 9649 263090 9683 263164
rect 10069 263090 10103 263164
rect 10489 263090 10523 263164
rect 10909 263090 10943 263164
rect 11329 263090 11363 263164
rect 11749 263090 11783 263164
rect 12169 263090 12203 263164
rect 12589 263090 12623 263164
rect 13009 263090 13043 263164
rect 13429 263090 13463 263164
rect 13849 263090 13883 263164
rect 14269 263090 14303 263164
rect 14689 263090 14723 263164
rect 15109 263090 15143 263164
rect 15529 263090 15563 263164
rect 15949 263090 15983 263164
rect 16369 263090 16403 263164
rect 16789 263090 16823 263164
rect 17209 263090 17243 263164
rect 17629 263090 17663 263164
rect 18049 263090 18083 263164
rect 18469 263090 18503 263164
rect 18889 263090 18923 263164
rect 19309 263090 19343 263164
rect 19729 263090 19763 263164
rect 20149 263090 20183 263164
rect 20569 263090 20603 263164
rect 20989 263090 21023 263164
rect 21409 263090 21443 263164
rect 21829 263090 21863 263164
rect 22249 263090 22283 263164
rect 22669 263090 22703 263164
rect 23089 263090 23123 263164
rect 23509 263090 23543 263164
rect 23929 263090 23963 263164
rect 24349 263090 24383 263164
rect 24769 263090 24803 263164
rect 25189 263090 25223 263164
rect 25609 263090 25643 263164
rect 26029 263090 26063 263164
rect 26449 263090 26483 263164
rect 26869 263090 26903 263164
rect 27289 263090 27323 263164
rect -3791 263056 -3757 263090
rect -3371 263056 -3337 263090
rect -2951 263056 -2917 263090
rect -2531 263056 -2497 263090
rect -2111 263056 -2077 263090
rect -1691 263056 -1657 263090
rect -1271 263056 -1237 263090
rect -851 263056 -817 263090
rect -431 263056 -397 263090
rect -11 263056 23 263090
rect 409 263056 443 263090
rect 829 263056 863 263090
rect 1249 263056 1283 263090
rect 1669 263056 1703 263090
rect 2089 263056 2123 263090
rect 2509 263056 2543 263090
rect 2929 263056 2963 263090
rect 3349 263056 3383 263090
rect 3769 263056 3803 263090
rect 4189 263056 4223 263090
rect 4609 263056 4643 263090
rect 5029 263056 5063 263090
rect 5449 263056 5483 263090
rect 5869 263056 5903 263090
rect 6289 263056 6323 263090
rect 6709 263056 6743 263090
rect 7129 263056 7163 263090
rect 7549 263056 7583 263090
rect 7969 263056 8003 263090
rect 8389 263056 8423 263090
rect 8809 263056 8843 263090
rect 9229 263056 9263 263090
rect 9649 263056 9683 263090
rect 10069 263056 10103 263090
rect 10489 263056 10523 263090
rect 10909 263056 10943 263090
rect 11329 263056 11363 263090
rect 11749 263056 11783 263090
rect 12169 263056 12203 263090
rect 12589 263056 12623 263090
rect 13009 263056 13043 263090
rect 13429 263056 13463 263090
rect 13849 263056 13883 263090
rect 14269 263056 14303 263090
rect 14689 263056 14723 263090
rect 15109 263056 15143 263090
rect 15529 263056 15563 263090
rect 15949 263056 15983 263090
rect 16369 263056 16403 263090
rect 16789 263056 16823 263090
rect 17209 263056 17243 263090
rect 17629 263056 17663 263090
rect 18049 263056 18083 263090
rect 18469 263056 18503 263090
rect 18889 263056 18923 263090
rect 19309 263056 19343 263090
rect 19729 263056 19763 263090
rect 20149 263056 20183 263090
rect 20569 263056 20603 263090
rect 20989 263056 21023 263090
rect 21409 263056 21443 263090
rect 21829 263056 21863 263090
rect 22249 263056 22283 263090
rect 22669 263056 22703 263090
rect 23089 263056 23123 263090
rect 23509 263056 23543 263090
rect 23929 263056 23963 263090
rect 24349 263056 24383 263090
rect 24769 263056 24803 263090
rect 25189 263056 25223 263090
rect 25609 263056 25643 263090
rect 26029 263056 26063 263090
rect 26449 263056 26483 263090
rect 26869 263056 26903 263090
rect 27289 263056 27323 263090
rect -4049 262228 -4015 263004
rect -3953 262228 -3919 263004
rect -3839 262228 -3805 263004
rect -3743 262228 -3709 263004
rect -3629 262228 -3595 263004
rect -3533 262228 -3499 263004
rect -3419 262228 -3385 263004
rect -3323 262228 -3289 263004
rect -3209 262228 -3175 263004
rect -3113 262228 -3079 263004
rect -2999 262228 -2965 263004
rect -2903 262228 -2869 263004
rect -2789 262228 -2755 263004
rect -2693 262228 -2659 263004
rect -2579 262228 -2545 263004
rect -2483 262228 -2449 263004
rect -2369 262228 -2335 263004
rect -2273 262228 -2239 263004
rect -2159 262228 -2125 263004
rect -2063 262228 -2029 263004
rect -1949 262228 -1915 263004
rect -1853 262228 -1819 263004
rect -1739 262228 -1705 263004
rect -1643 262228 -1609 263004
rect -1529 262228 -1495 263004
rect -1433 262228 -1399 263004
rect -1319 262228 -1285 263004
rect -1223 262228 -1189 263004
rect -1109 262228 -1075 263004
rect -1013 262228 -979 263004
rect -899 262228 -865 263004
rect -803 262228 -769 263004
rect -689 262228 -655 263004
rect -593 262228 -559 263004
rect -479 262228 -445 263004
rect -383 262228 -349 263004
rect -269 262228 -235 263004
rect -173 262228 -139 263004
rect -59 262228 -25 263004
rect 37 262228 71 263004
rect 151 262228 185 263004
rect 247 262228 281 263004
rect 361 262228 395 263004
rect 457 262228 491 263004
rect 571 262228 605 263004
rect 667 262228 701 263004
rect 781 262228 815 263004
rect 877 262228 911 263004
rect 991 262228 1025 263004
rect 1087 262228 1121 263004
rect 1201 262228 1235 263004
rect 1297 262228 1331 263004
rect 1411 262228 1445 263004
rect 1507 262228 1541 263004
rect 1621 262228 1655 263004
rect 1717 262228 1751 263004
rect 1831 262228 1865 263004
rect 1927 262228 1961 263004
rect 2041 262228 2075 263004
rect 2137 262228 2171 263004
rect 2251 262228 2285 263004
rect 2347 262228 2381 263004
rect 2461 262228 2495 263004
rect 2557 262228 2591 263004
rect 2671 262228 2705 263004
rect 2767 262228 2801 263004
rect 2881 262228 2915 263004
rect 2977 262228 3011 263004
rect 3091 262228 3125 263004
rect 3187 262228 3221 263004
rect 3301 262228 3335 263004
rect 3397 262228 3431 263004
rect 3511 262228 3545 263004
rect 3607 262228 3641 263004
rect 3721 262228 3755 263004
rect 3817 262228 3851 263004
rect 3931 262228 3965 263004
rect 4027 262228 4061 263004
rect 4141 262228 4175 263004
rect 4237 262228 4271 263004
rect 4351 262228 4385 263004
rect 4447 262228 4481 263004
rect 4561 262228 4595 263004
rect 4657 262228 4691 263004
rect 4771 262228 4805 263004
rect 4867 262228 4901 263004
rect 4981 262228 5015 263004
rect 5077 262228 5111 263004
rect 5191 262228 5225 263004
rect 5287 262228 5321 263004
rect 5401 262228 5435 263004
rect 5497 262228 5531 263004
rect 5611 262228 5645 263004
rect 5707 262228 5741 263004
rect 5821 262228 5855 263004
rect 5917 262228 5951 263004
rect 6031 262228 6065 263004
rect 6127 262228 6161 263004
rect 6241 262228 6275 263004
rect 6337 262228 6371 263004
rect 6451 262228 6485 263004
rect 6547 262228 6581 263004
rect 6661 262228 6695 263004
rect 6757 262228 6791 263004
rect 6871 262228 6905 263004
rect 6967 262228 7001 263004
rect 7081 262228 7115 263004
rect 7177 262228 7211 263004
rect 7291 262228 7325 263004
rect 7387 262228 7421 263004
rect 7501 262228 7535 263004
rect 7597 262228 7631 263004
rect 7711 262228 7745 263004
rect 7807 262228 7841 263004
rect 7921 262228 7955 263004
rect 8017 262228 8051 263004
rect 8131 262228 8165 263004
rect 8227 262228 8261 263004
rect 8341 262228 8375 263004
rect 8437 262228 8471 263004
rect 8551 262228 8585 263004
rect 8647 262228 8681 263004
rect 8761 262228 8795 263004
rect 8857 262228 8891 263004
rect 8971 262228 9005 263004
rect 9067 262228 9101 263004
rect 9181 262228 9215 263004
rect 9277 262228 9311 263004
rect 9391 262228 9425 263004
rect 9487 262228 9521 263004
rect 9601 262228 9635 263004
rect 9697 262228 9731 263004
rect 9811 262228 9845 263004
rect 9907 262228 9941 263004
rect 10021 262228 10055 263004
rect 10117 262228 10151 263004
rect 10231 262228 10265 263004
rect 10327 262228 10361 263004
rect 10441 262228 10475 263004
rect 10537 262228 10571 263004
rect 10651 262228 10685 263004
rect 10747 262228 10781 263004
rect 10861 262228 10895 263004
rect 10957 262228 10991 263004
rect 11071 262228 11105 263004
rect 11167 262228 11201 263004
rect 11281 262228 11315 263004
rect 11377 262228 11411 263004
rect 11491 262228 11525 263004
rect 11587 262228 11621 263004
rect 11701 262228 11735 263004
rect 11797 262228 11831 263004
rect 11911 262228 11945 263004
rect 12007 262228 12041 263004
rect 12121 262228 12155 263004
rect 12217 262228 12251 263004
rect 12331 262228 12365 263004
rect 12427 262228 12461 263004
rect 12541 262228 12575 263004
rect 12637 262228 12671 263004
rect 12751 262228 12785 263004
rect 12847 262228 12881 263004
rect 12961 262228 12995 263004
rect 13057 262228 13091 263004
rect 13171 262228 13205 263004
rect 13267 262228 13301 263004
rect 13381 262228 13415 263004
rect 13477 262228 13511 263004
rect 13591 262228 13625 263004
rect 13687 262228 13721 263004
rect 13801 262228 13835 263004
rect 13897 262228 13931 263004
rect 14011 262228 14045 263004
rect 14107 262228 14141 263004
rect 14221 262228 14255 263004
rect 14317 262228 14351 263004
rect 14431 262228 14465 263004
rect 14527 262228 14561 263004
rect 14641 262228 14675 263004
rect 14737 262228 14771 263004
rect 14851 262228 14885 263004
rect 14947 262228 14981 263004
rect 15061 262228 15095 263004
rect 15157 262228 15191 263004
rect 15271 262228 15305 263004
rect 15367 262228 15401 263004
rect 15481 262228 15515 263004
rect 15577 262228 15611 263004
rect 15691 262228 15725 263004
rect 15787 262228 15821 263004
rect 15901 262228 15935 263004
rect 15997 262228 16031 263004
rect 16111 262228 16145 263004
rect 16207 262228 16241 263004
rect 16321 262228 16355 263004
rect 16417 262228 16451 263004
rect 16531 262228 16565 263004
rect 16627 262228 16661 263004
rect 16741 262228 16775 263004
rect 16837 262228 16871 263004
rect 16951 262228 16985 263004
rect 17047 262228 17081 263004
rect 17161 262228 17195 263004
rect 17257 262228 17291 263004
rect 17371 262228 17405 263004
rect 17467 262228 17501 263004
rect 17581 262228 17615 263004
rect 17677 262228 17711 263004
rect 17791 262228 17825 263004
rect 17887 262228 17921 263004
rect 18001 262228 18035 263004
rect 18097 262228 18131 263004
rect 18211 262228 18245 263004
rect 18307 262228 18341 263004
rect 18421 262228 18455 263004
rect 18517 262228 18551 263004
rect 18631 262228 18665 263004
rect 18727 262228 18761 263004
rect 18841 262228 18875 263004
rect 18937 262228 18971 263004
rect 19051 262228 19085 263004
rect 19147 262228 19181 263004
rect 19261 262228 19295 263004
rect 19357 262228 19391 263004
rect 19471 262228 19505 263004
rect 19567 262228 19601 263004
rect 19681 262228 19715 263004
rect 19777 262228 19811 263004
rect 19891 262228 19925 263004
rect 19987 262228 20021 263004
rect 20101 262228 20135 263004
rect 20197 262228 20231 263004
rect 20311 262228 20345 263004
rect 20407 262228 20441 263004
rect 20521 262228 20555 263004
rect 20617 262228 20651 263004
rect 20731 262228 20765 263004
rect 20827 262228 20861 263004
rect 20941 262228 20975 263004
rect 21037 262228 21071 263004
rect 21151 262228 21185 263004
rect 21247 262228 21281 263004
rect 21361 262228 21395 263004
rect 21457 262228 21491 263004
rect 21571 262228 21605 263004
rect 21667 262228 21701 263004
rect 21781 262228 21815 263004
rect 21877 262228 21911 263004
rect 21991 262228 22025 263004
rect 22087 262228 22121 263004
rect 22201 262228 22235 263004
rect 22297 262228 22331 263004
rect 22411 262228 22445 263004
rect 22507 262228 22541 263004
rect 22621 262228 22655 263004
rect 22717 262228 22751 263004
rect 22831 262228 22865 263004
rect 22927 262228 22961 263004
rect 23041 262228 23075 263004
rect 23137 262228 23171 263004
rect 23251 262228 23285 263004
rect 23347 262228 23381 263004
rect 23461 262228 23495 263004
rect 23557 262228 23591 263004
rect 23671 262228 23705 263004
rect 23767 262228 23801 263004
rect 23881 262228 23915 263004
rect 23977 262228 24011 263004
rect 24091 262228 24125 263004
rect 24187 262228 24221 263004
rect 24301 262228 24335 263004
rect 24397 262228 24431 263004
rect 24511 262228 24545 263004
rect 24607 262228 24641 263004
rect 24721 262228 24755 263004
rect 24817 262228 24851 263004
rect 24931 262228 24965 263004
rect 25027 262228 25061 263004
rect 25141 262228 25175 263004
rect 25237 262228 25271 263004
rect 25351 262228 25385 263004
rect 25447 262228 25481 263004
rect 25561 262228 25595 263004
rect 25657 262228 25691 263004
rect 25771 262228 25805 263004
rect 25867 262228 25901 263004
rect 25981 262228 26015 263004
rect 26077 262228 26111 263004
rect 26191 262228 26225 263004
rect 26287 262228 26321 263004
rect 26401 262228 26435 263004
rect 26497 262228 26531 263004
rect 26611 262228 26645 263004
rect 26707 262228 26741 263004
rect 26821 262228 26855 263004
rect 26917 262228 26951 263004
rect 27031 262228 27065 263004
rect 27127 262228 27161 263004
rect 27241 262228 27275 263004
rect 27337 262228 27371 263004
rect -4001 262144 -3905 262178
rect -3581 262144 -3485 262178
rect -3161 262144 -3065 262178
rect -2741 262144 -2645 262178
rect -2321 262144 -2225 262178
rect -1901 262144 -1805 262178
rect -1481 262144 -1385 262178
rect -1061 262144 -965 262178
rect -641 262144 -545 262178
rect -221 262144 -125 262178
rect 199 262144 295 262178
rect 619 262144 715 262178
rect 1039 262144 1135 262178
rect 1459 262144 1555 262178
rect 1879 262144 1975 262178
rect 2299 262144 2395 262178
rect 2719 262144 2815 262178
rect 3139 262144 3235 262178
rect 3559 262144 3655 262178
rect 3979 262144 4075 262178
rect 4399 262144 4495 262178
rect 4819 262144 4915 262178
rect 5239 262144 5335 262178
rect 5659 262144 5755 262178
rect 6079 262144 6175 262178
rect 6499 262144 6595 262178
rect 6919 262144 7015 262178
rect 7339 262144 7435 262178
rect 7759 262144 7855 262178
rect 8179 262144 8275 262178
rect 8599 262144 8695 262178
rect 9019 262144 9115 262178
rect 9439 262144 9535 262178
rect 9859 262144 9955 262178
rect 10279 262144 10375 262178
rect 10699 262144 10795 262178
rect 11119 262144 11215 262178
rect 11539 262144 11635 262178
rect 11959 262144 12055 262178
rect 12379 262144 12475 262178
rect 12799 262144 12895 262178
rect 13219 262144 13315 262178
rect 13639 262144 13735 262178
rect 14059 262144 14155 262178
rect 14479 262144 14575 262178
rect 14899 262144 14995 262178
rect 15319 262144 15415 262178
rect 15739 262144 15835 262178
rect 16159 262144 16255 262178
rect 16579 262144 16675 262178
rect 16999 262144 17095 262178
rect 17419 262144 17515 262178
rect 17839 262144 17935 262178
rect 18259 262144 18355 262178
rect 18679 262144 18775 262178
rect 19099 262144 19195 262178
rect 19519 262144 19615 262178
rect 19939 262144 20035 262178
rect 20359 262144 20455 262178
rect 20779 262144 20875 262178
rect 21199 262144 21295 262178
rect 21619 262144 21715 262178
rect 22039 262144 22135 262178
rect 22459 262144 22555 262178
rect 22879 262144 22975 262178
rect 23299 262144 23395 262178
rect 23719 262144 23815 262178
rect 24139 262144 24235 262178
rect 24559 262144 24655 262178
rect 24979 262144 25075 262178
rect 25399 262144 25495 262178
rect 25819 262144 25915 262178
rect 26239 262144 26335 262178
rect 26659 262144 26755 262178
rect 27079 262144 27175 262178
rect -4001 254548 -3905 254582
rect -3581 254548 -3485 254582
rect -3161 254548 -3065 254582
rect -2741 254548 -2645 254582
rect -2321 254548 -2225 254582
rect -1901 254548 -1805 254582
rect -1481 254548 -1385 254582
rect -1061 254548 -965 254582
rect -641 254548 -545 254582
rect -221 254548 -125 254582
rect 199 254548 295 254582
rect 619 254548 715 254582
rect 1039 254548 1135 254582
rect 1459 254548 1555 254582
rect 1879 254548 1975 254582
rect 2299 254548 2395 254582
rect 2719 254548 2815 254582
rect 3139 254548 3235 254582
rect 3559 254548 3655 254582
rect 3979 254548 4075 254582
rect 4399 254548 4495 254582
rect 4819 254548 4915 254582
rect 5239 254548 5335 254582
rect 5659 254548 5755 254582
rect 6079 254548 6175 254582
rect 6499 254548 6595 254582
rect 6919 254548 7015 254582
rect 7339 254548 7435 254582
rect 7759 254548 7855 254582
rect 8179 254548 8275 254582
rect 8599 254548 8695 254582
rect 9019 254548 9115 254582
rect 9439 254548 9535 254582
rect 9859 254548 9955 254582
rect 10279 254548 10375 254582
rect 10699 254548 10795 254582
rect 11119 254548 11215 254582
rect 11539 254548 11635 254582
rect 11959 254548 12055 254582
rect 12379 254548 12475 254582
rect 12799 254548 12895 254582
rect 13219 254548 13315 254582
rect 13639 254548 13735 254582
rect 14059 254548 14155 254582
rect 14479 254548 14575 254582
rect 14899 254548 14995 254582
rect 15319 254548 15415 254582
rect 15739 254548 15835 254582
rect 16159 254548 16255 254582
rect 16579 254548 16675 254582
rect 16999 254548 17095 254582
rect 17419 254548 17515 254582
rect 17839 254548 17935 254582
rect 18259 254548 18355 254582
rect 18679 254548 18775 254582
rect 19099 254548 19195 254582
rect 19519 254548 19615 254582
rect 19939 254548 20035 254582
rect 20359 254548 20455 254582
rect 20779 254548 20875 254582
rect 21199 254548 21295 254582
rect 21619 254548 21715 254582
rect 22039 254548 22135 254582
rect 22459 254548 22555 254582
rect 22879 254548 22975 254582
rect 23299 254548 23395 254582
rect 23719 254548 23815 254582
rect 24139 254548 24235 254582
rect 24559 254548 24655 254582
rect 24979 254548 25075 254582
rect 25399 254548 25495 254582
rect 25819 254548 25915 254582
rect 26239 254548 26335 254582
rect 26659 254548 26755 254582
rect 27079 254548 27175 254582
rect -4049 253713 -4015 254489
rect -3953 253713 -3919 254489
rect -3839 253713 -3805 254489
rect -3743 253713 -3709 254489
rect -3629 253713 -3595 254489
rect -3533 253713 -3499 254489
rect -3419 253713 -3385 254489
rect -3323 253713 -3289 254489
rect -3209 253713 -3175 254489
rect -3113 253713 -3079 254489
rect -2999 253713 -2965 254489
rect -2903 253713 -2869 254489
rect -2789 253713 -2755 254489
rect -2693 253713 -2659 254489
rect -2579 253713 -2545 254489
rect -2483 253713 -2449 254489
rect -2369 253713 -2335 254489
rect -2273 253713 -2239 254489
rect -2159 253713 -2125 254489
rect -2063 253713 -2029 254489
rect -1949 253713 -1915 254489
rect -1853 253713 -1819 254489
rect -1739 253713 -1705 254489
rect -1643 253713 -1609 254489
rect -1529 253713 -1495 254489
rect -1433 253713 -1399 254489
rect -1319 253713 -1285 254489
rect -1223 253713 -1189 254489
rect -1109 253713 -1075 254489
rect -1013 253713 -979 254489
rect -899 253713 -865 254489
rect -803 253713 -769 254489
rect -689 253713 -655 254489
rect -593 253713 -559 254489
rect -479 253713 -445 254489
rect -383 253713 -349 254489
rect -269 253713 -235 254489
rect -173 253713 -139 254489
rect -59 253713 -25 254489
rect 37 253713 71 254489
rect 151 253713 185 254489
rect 247 253713 281 254489
rect 361 253713 395 254489
rect 457 253713 491 254489
rect 571 253713 605 254489
rect 667 253713 701 254489
rect 781 253713 815 254489
rect 877 253713 911 254489
rect 991 253713 1025 254489
rect 1087 253713 1121 254489
rect 1201 253713 1235 254489
rect 1297 253713 1331 254489
rect 1411 253713 1445 254489
rect 1507 253713 1541 254489
rect 1621 253713 1655 254489
rect 1717 253713 1751 254489
rect 1831 253713 1865 254489
rect 1927 253713 1961 254489
rect 2041 253713 2075 254489
rect 2137 253713 2171 254489
rect 2251 253713 2285 254489
rect 2347 253713 2381 254489
rect 2461 253713 2495 254489
rect 2557 253713 2591 254489
rect 2671 253713 2705 254489
rect 2767 253713 2801 254489
rect 2881 253713 2915 254489
rect 2977 253713 3011 254489
rect 3091 253713 3125 254489
rect 3187 253713 3221 254489
rect 3301 253713 3335 254489
rect 3397 253713 3431 254489
rect 3511 253713 3545 254489
rect 3607 253713 3641 254489
rect 3721 253713 3755 254489
rect 3817 253713 3851 254489
rect 3931 253713 3965 254489
rect 4027 253713 4061 254489
rect 4141 253713 4175 254489
rect 4237 253713 4271 254489
rect 4351 253713 4385 254489
rect 4447 253713 4481 254489
rect 4561 253713 4595 254489
rect 4657 253713 4691 254489
rect 4771 253713 4805 254489
rect 4867 253713 4901 254489
rect 4981 253713 5015 254489
rect 5077 253713 5111 254489
rect 5191 253713 5225 254489
rect 5287 253713 5321 254489
rect 5401 253713 5435 254489
rect 5497 253713 5531 254489
rect 5611 253713 5645 254489
rect 5707 253713 5741 254489
rect 5821 253713 5855 254489
rect 5917 253713 5951 254489
rect 6031 253713 6065 254489
rect 6127 253713 6161 254489
rect 6241 253713 6275 254489
rect 6337 253713 6371 254489
rect 6451 253713 6485 254489
rect 6547 253713 6581 254489
rect 6661 253713 6695 254489
rect 6757 253713 6791 254489
rect 6871 253713 6905 254489
rect 6967 253713 7001 254489
rect 7081 253713 7115 254489
rect 7177 253713 7211 254489
rect 7291 253713 7325 254489
rect 7387 253713 7421 254489
rect 7501 253713 7535 254489
rect 7597 253713 7631 254489
rect 7711 253713 7745 254489
rect 7807 253713 7841 254489
rect 7921 253713 7955 254489
rect 8017 253713 8051 254489
rect 8131 253713 8165 254489
rect 8227 253713 8261 254489
rect 8341 253713 8375 254489
rect 8437 253713 8471 254489
rect 8551 253713 8585 254489
rect 8647 253713 8681 254489
rect 8761 253713 8795 254489
rect 8857 253713 8891 254489
rect 8971 253713 9005 254489
rect 9067 253713 9101 254489
rect 9181 253713 9215 254489
rect 9277 253713 9311 254489
rect 9391 253713 9425 254489
rect 9487 253713 9521 254489
rect 9601 253713 9635 254489
rect 9697 253713 9731 254489
rect 9811 253713 9845 254489
rect 9907 253713 9941 254489
rect 10021 253713 10055 254489
rect 10117 253713 10151 254489
rect 10231 253713 10265 254489
rect 10327 253713 10361 254489
rect 10441 253713 10475 254489
rect 10537 253713 10571 254489
rect 10651 253713 10685 254489
rect 10747 253713 10781 254489
rect 10861 253713 10895 254489
rect 10957 253713 10991 254489
rect 11071 253713 11105 254489
rect 11167 253713 11201 254489
rect 11281 253713 11315 254489
rect 11377 253713 11411 254489
rect 11491 253713 11525 254489
rect 11587 253713 11621 254489
rect 11701 253713 11735 254489
rect 11797 253713 11831 254489
rect 11911 253713 11945 254489
rect 12007 253713 12041 254489
rect 12121 253713 12155 254489
rect 12217 253713 12251 254489
rect 12331 253713 12365 254489
rect 12427 253713 12461 254489
rect 12541 253713 12575 254489
rect 12637 253713 12671 254489
rect 12751 253713 12785 254489
rect 12847 253713 12881 254489
rect 12961 253713 12995 254489
rect 13057 253713 13091 254489
rect 13171 253713 13205 254489
rect 13267 253713 13301 254489
rect 13381 253713 13415 254489
rect 13477 253713 13511 254489
rect 13591 253713 13625 254489
rect 13687 253713 13721 254489
rect 13801 253713 13835 254489
rect 13897 253713 13931 254489
rect 14011 253713 14045 254489
rect 14107 253713 14141 254489
rect 14221 253713 14255 254489
rect 14317 253713 14351 254489
rect 14431 253713 14465 254489
rect 14527 253713 14561 254489
rect 14641 253713 14675 254489
rect 14737 253713 14771 254489
rect 14851 253713 14885 254489
rect 14947 253713 14981 254489
rect 15061 253713 15095 254489
rect 15157 253713 15191 254489
rect 15271 253713 15305 254489
rect 15367 253713 15401 254489
rect 15481 253713 15515 254489
rect 15577 253713 15611 254489
rect 15691 253713 15725 254489
rect 15787 253713 15821 254489
rect 15901 253713 15935 254489
rect 15997 253713 16031 254489
rect 16111 253713 16145 254489
rect 16207 253713 16241 254489
rect 16321 253713 16355 254489
rect 16417 253713 16451 254489
rect 16531 253713 16565 254489
rect 16627 253713 16661 254489
rect 16741 253713 16775 254489
rect 16837 253713 16871 254489
rect 16951 253713 16985 254489
rect 17047 253713 17081 254489
rect 17161 253713 17195 254489
rect 17257 253713 17291 254489
rect 17371 253713 17405 254489
rect 17467 253713 17501 254489
rect 17581 253713 17615 254489
rect 17677 253713 17711 254489
rect 17791 253713 17825 254489
rect 17887 253713 17921 254489
rect 18001 253713 18035 254489
rect 18097 253713 18131 254489
rect 18211 253713 18245 254489
rect 18307 253713 18341 254489
rect 18421 253713 18455 254489
rect 18517 253713 18551 254489
rect 18631 253713 18665 254489
rect 18727 253713 18761 254489
rect 18841 253713 18875 254489
rect 18937 253713 18971 254489
rect 19051 253713 19085 254489
rect 19147 253713 19181 254489
rect 19261 253713 19295 254489
rect 19357 253713 19391 254489
rect 19471 253713 19505 254489
rect 19567 253713 19601 254489
rect 19681 253713 19715 254489
rect 19777 253713 19811 254489
rect 19891 253713 19925 254489
rect 19987 253713 20021 254489
rect 20101 253713 20135 254489
rect 20197 253713 20231 254489
rect 20311 253713 20345 254489
rect 20407 253713 20441 254489
rect 20521 253713 20555 254489
rect 20617 253713 20651 254489
rect 20731 253713 20765 254489
rect 20827 253713 20861 254489
rect 20941 253713 20975 254489
rect 21037 253713 21071 254489
rect 21151 253713 21185 254489
rect 21247 253713 21281 254489
rect 21361 253713 21395 254489
rect 21457 253713 21491 254489
rect 21571 253713 21605 254489
rect 21667 253713 21701 254489
rect 21781 253713 21815 254489
rect 21877 253713 21911 254489
rect 21991 253713 22025 254489
rect 22087 253713 22121 254489
rect 22201 253713 22235 254489
rect 22297 253713 22331 254489
rect 22411 253713 22445 254489
rect 22507 253713 22541 254489
rect 22621 253713 22655 254489
rect 22717 253713 22751 254489
rect 22831 253713 22865 254489
rect 22927 253713 22961 254489
rect 23041 253713 23075 254489
rect 23137 253713 23171 254489
rect 23251 253713 23285 254489
rect 23347 253713 23381 254489
rect 23461 253713 23495 254489
rect 23557 253713 23591 254489
rect 23671 253713 23705 254489
rect 23767 253713 23801 254489
rect 23881 253713 23915 254489
rect 23977 253713 24011 254489
rect 24091 253713 24125 254489
rect 24187 253713 24221 254489
rect 24301 253713 24335 254489
rect 24397 253713 24431 254489
rect 24511 253713 24545 254489
rect 24607 253713 24641 254489
rect 24721 253713 24755 254489
rect 24817 253713 24851 254489
rect 24931 253713 24965 254489
rect 25027 253713 25061 254489
rect 25141 253713 25175 254489
rect 25237 253713 25271 254489
rect 25351 253713 25385 254489
rect 25447 253713 25481 254489
rect 25561 253713 25595 254489
rect 25657 253713 25691 254489
rect 25771 253713 25805 254489
rect 25867 253713 25901 254489
rect 25981 253713 26015 254489
rect 26077 253713 26111 254489
rect 26191 253713 26225 254489
rect 26287 253713 26321 254489
rect 26401 253713 26435 254489
rect 26497 253713 26531 254489
rect 26611 253713 26645 254489
rect 26707 253713 26741 254489
rect 26821 253713 26855 254489
rect 26917 253713 26951 254489
rect 27031 253713 27065 254489
rect 27127 253713 27161 254489
rect 27241 253713 27275 254489
rect 27337 253713 27371 254489
rect -3791 253512 -3757 253654
rect -3371 253512 -3337 253654
rect -2951 253512 -2917 253654
rect -2531 253512 -2497 253654
rect -2111 253512 -2077 253654
rect -1691 253512 -1657 253654
rect -1271 253512 -1237 253654
rect -851 253512 -817 253654
rect -431 253512 -397 253654
rect -11 253512 23 253654
rect 409 253512 443 253654
rect 829 253512 863 253654
rect 1249 253512 1283 253654
rect 1669 253512 1703 253654
rect 2089 253512 2123 253654
rect 2509 253512 2543 253654
rect 2929 253512 2963 253654
rect 3349 253512 3383 253654
rect 3769 253512 3803 253654
rect 4189 253512 4223 253654
rect 4609 253512 4643 253654
rect 5029 253512 5063 253654
rect 5449 253512 5483 253654
rect 5869 253512 5903 253654
rect 6289 253512 6323 253654
rect 6709 253512 6743 253654
rect 7129 253512 7163 253654
rect 7549 253512 7583 253654
rect 7969 253512 8003 253654
rect 8389 253512 8423 253654
rect 8809 253512 8843 253654
rect 9229 253512 9263 253654
rect 9649 253512 9683 253654
rect 10069 253512 10103 253654
rect 10489 253512 10523 253654
rect 10909 253512 10943 253654
rect 11329 253512 11363 253654
rect 11749 253512 11783 253654
rect 12169 253512 12203 253654
rect 12589 253512 12623 253654
rect 13009 253512 13043 253654
rect 13429 253512 13463 253654
rect 13849 253512 13883 253654
rect 14269 253512 14303 253654
rect 14689 253512 14723 253654
rect 15109 253512 15143 253654
rect 15529 253512 15563 253654
rect 15949 253512 15983 253654
rect 16369 253512 16403 253654
rect 16789 253512 16823 253654
rect 17209 253512 17243 253654
rect 17629 253512 17663 253654
rect 18049 253512 18083 253654
rect 18469 253512 18503 253654
rect 18889 253512 18923 253654
rect 19309 253512 19343 253654
rect 19729 253512 19763 253654
rect 20149 253512 20183 253654
rect 20569 253512 20603 253654
rect 20989 253512 21023 253654
rect 21409 253512 21443 253654
rect 21829 253512 21863 253654
rect 22249 253512 22283 253654
rect 22669 253512 22703 253654
rect 23089 253512 23123 253654
rect 23509 253512 23543 253654
rect 23929 253512 23963 253654
rect 24349 253512 24383 253654
rect 24769 253512 24803 253654
rect 25189 253512 25223 253654
rect 25609 253512 25643 253654
rect 26029 253512 26063 253654
rect 26449 253512 26483 253654
rect 26869 253512 26903 253654
rect 27289 253512 27323 253654
rect -4049 252677 -4015 253453
rect -3953 252677 -3919 253453
rect -3839 252677 -3805 253453
rect -3743 252677 -3709 253453
rect -3629 252677 -3595 253453
rect -3533 252677 -3499 253453
rect -3419 252677 -3385 253453
rect -3323 252677 -3289 253453
rect -3209 252677 -3175 253453
rect -3113 252677 -3079 253453
rect -2999 252677 -2965 253453
rect -2903 252677 -2869 253453
rect -2789 252677 -2755 253453
rect -2693 252677 -2659 253453
rect -2579 252677 -2545 253453
rect -2483 252677 -2449 253453
rect -2369 252677 -2335 253453
rect -2273 252677 -2239 253453
rect -2159 252677 -2125 253453
rect -2063 252677 -2029 253453
rect -1949 252677 -1915 253453
rect -1853 252677 -1819 253453
rect -1739 252677 -1705 253453
rect -1643 252677 -1609 253453
rect -1529 252677 -1495 253453
rect -1433 252677 -1399 253453
rect -1319 252677 -1285 253453
rect -1223 252677 -1189 253453
rect -1109 252677 -1075 253453
rect -1013 252677 -979 253453
rect -899 252677 -865 253453
rect -803 252677 -769 253453
rect -689 252677 -655 253453
rect -593 252677 -559 253453
rect -479 252677 -445 253453
rect -383 252677 -349 253453
rect -269 252677 -235 253453
rect -173 252677 -139 253453
rect -59 252677 -25 253453
rect 37 252677 71 253453
rect 151 252677 185 253453
rect 247 252677 281 253453
rect 361 252677 395 253453
rect 457 252677 491 253453
rect 571 252677 605 253453
rect 667 252677 701 253453
rect 781 252677 815 253453
rect 877 252677 911 253453
rect 991 252677 1025 253453
rect 1087 252677 1121 253453
rect 1201 252677 1235 253453
rect 1297 252677 1331 253453
rect 1411 252677 1445 253453
rect 1507 252677 1541 253453
rect 1621 252677 1655 253453
rect 1717 252677 1751 253453
rect 1831 252677 1865 253453
rect 1927 252677 1961 253453
rect 2041 252677 2075 253453
rect 2137 252677 2171 253453
rect 2251 252677 2285 253453
rect 2347 252677 2381 253453
rect 2461 252677 2495 253453
rect 2557 252677 2591 253453
rect 2671 252677 2705 253453
rect 2767 252677 2801 253453
rect 2881 252677 2915 253453
rect 2977 252677 3011 253453
rect 3091 252677 3125 253453
rect 3187 252677 3221 253453
rect 3301 252677 3335 253453
rect 3397 252677 3431 253453
rect 3511 252677 3545 253453
rect 3607 252677 3641 253453
rect 3721 252677 3755 253453
rect 3817 252677 3851 253453
rect 3931 252677 3965 253453
rect 4027 252677 4061 253453
rect 4141 252677 4175 253453
rect 4237 252677 4271 253453
rect 4351 252677 4385 253453
rect 4447 252677 4481 253453
rect 4561 252677 4595 253453
rect 4657 252677 4691 253453
rect 4771 252677 4805 253453
rect 4867 252677 4901 253453
rect 4981 252677 5015 253453
rect 5077 252677 5111 253453
rect 5191 252677 5225 253453
rect 5287 252677 5321 253453
rect 5401 252677 5435 253453
rect 5497 252677 5531 253453
rect 5611 252677 5645 253453
rect 5707 252677 5741 253453
rect 5821 252677 5855 253453
rect 5917 252677 5951 253453
rect 6031 252677 6065 253453
rect 6127 252677 6161 253453
rect 6241 252677 6275 253453
rect 6337 252677 6371 253453
rect 6451 252677 6485 253453
rect 6547 252677 6581 253453
rect 6661 252677 6695 253453
rect 6757 252677 6791 253453
rect 6871 252677 6905 253453
rect 6967 252677 7001 253453
rect 7081 252677 7115 253453
rect 7177 252677 7211 253453
rect 7291 252677 7325 253453
rect 7387 252677 7421 253453
rect 7501 252677 7535 253453
rect 7597 252677 7631 253453
rect 7711 252677 7745 253453
rect 7807 252677 7841 253453
rect 7921 252677 7955 253453
rect 8017 252677 8051 253453
rect 8131 252677 8165 253453
rect 8227 252677 8261 253453
rect 8341 252677 8375 253453
rect 8437 252677 8471 253453
rect 8551 252677 8585 253453
rect 8647 252677 8681 253453
rect 8761 252677 8795 253453
rect 8857 252677 8891 253453
rect 8971 252677 9005 253453
rect 9067 252677 9101 253453
rect 9181 252677 9215 253453
rect 9277 252677 9311 253453
rect 9391 252677 9425 253453
rect 9487 252677 9521 253453
rect 9601 252677 9635 253453
rect 9697 252677 9731 253453
rect 9811 252677 9845 253453
rect 9907 252677 9941 253453
rect 10021 252677 10055 253453
rect 10117 252677 10151 253453
rect 10231 252677 10265 253453
rect 10327 252677 10361 253453
rect 10441 252677 10475 253453
rect 10537 252677 10571 253453
rect 10651 252677 10685 253453
rect 10747 252677 10781 253453
rect 10861 252677 10895 253453
rect 10957 252677 10991 253453
rect 11071 252677 11105 253453
rect 11167 252677 11201 253453
rect 11281 252677 11315 253453
rect 11377 252677 11411 253453
rect 11491 252677 11525 253453
rect 11587 252677 11621 253453
rect 11701 252677 11735 253453
rect 11797 252677 11831 253453
rect 11911 252677 11945 253453
rect 12007 252677 12041 253453
rect 12121 252677 12155 253453
rect 12217 252677 12251 253453
rect 12331 252677 12365 253453
rect 12427 252677 12461 253453
rect 12541 252677 12575 253453
rect 12637 252677 12671 253453
rect 12751 252677 12785 253453
rect 12847 252677 12881 253453
rect 12961 252677 12995 253453
rect 13057 252677 13091 253453
rect 13171 252677 13205 253453
rect 13267 252677 13301 253453
rect 13381 252677 13415 253453
rect 13477 252677 13511 253453
rect 13591 252677 13625 253453
rect 13687 252677 13721 253453
rect 13801 252677 13835 253453
rect 13897 252677 13931 253453
rect 14011 252677 14045 253453
rect 14107 252677 14141 253453
rect 14221 252677 14255 253453
rect 14317 252677 14351 253453
rect 14431 252677 14465 253453
rect 14527 252677 14561 253453
rect 14641 252677 14675 253453
rect 14737 252677 14771 253453
rect 14851 252677 14885 253453
rect 14947 252677 14981 253453
rect 15061 252677 15095 253453
rect 15157 252677 15191 253453
rect 15271 252677 15305 253453
rect 15367 252677 15401 253453
rect 15481 252677 15515 253453
rect 15577 252677 15611 253453
rect 15691 252677 15725 253453
rect 15787 252677 15821 253453
rect 15901 252677 15935 253453
rect 15997 252677 16031 253453
rect 16111 252677 16145 253453
rect 16207 252677 16241 253453
rect 16321 252677 16355 253453
rect 16417 252677 16451 253453
rect 16531 252677 16565 253453
rect 16627 252677 16661 253453
rect 16741 252677 16775 253453
rect 16837 252677 16871 253453
rect 16951 252677 16985 253453
rect 17047 252677 17081 253453
rect 17161 252677 17195 253453
rect 17257 252677 17291 253453
rect 17371 252677 17405 253453
rect 17467 252677 17501 253453
rect 17581 252677 17615 253453
rect 17677 252677 17711 253453
rect 17791 252677 17825 253453
rect 17887 252677 17921 253453
rect 18001 252677 18035 253453
rect 18097 252677 18131 253453
rect 18211 252677 18245 253453
rect 18307 252677 18341 253453
rect 18421 252677 18455 253453
rect 18517 252677 18551 253453
rect 18631 252677 18665 253453
rect 18727 252677 18761 253453
rect 18841 252677 18875 253453
rect 18937 252677 18971 253453
rect 19051 252677 19085 253453
rect 19147 252677 19181 253453
rect 19261 252677 19295 253453
rect 19357 252677 19391 253453
rect 19471 252677 19505 253453
rect 19567 252677 19601 253453
rect 19681 252677 19715 253453
rect 19777 252677 19811 253453
rect 19891 252677 19925 253453
rect 19987 252677 20021 253453
rect 20101 252677 20135 253453
rect 20197 252677 20231 253453
rect 20311 252677 20345 253453
rect 20407 252677 20441 253453
rect 20521 252677 20555 253453
rect 20617 252677 20651 253453
rect 20731 252677 20765 253453
rect 20827 252677 20861 253453
rect 20941 252677 20975 253453
rect 21037 252677 21071 253453
rect 21151 252677 21185 253453
rect 21247 252677 21281 253453
rect 21361 252677 21395 253453
rect 21457 252677 21491 253453
rect 21571 252677 21605 253453
rect 21667 252677 21701 253453
rect 21781 252677 21815 253453
rect 21877 252677 21911 253453
rect 21991 252677 22025 253453
rect 22087 252677 22121 253453
rect 22201 252677 22235 253453
rect 22297 252677 22331 253453
rect 22411 252677 22445 253453
rect 22507 252677 22541 253453
rect 22621 252677 22655 253453
rect 22717 252677 22751 253453
rect 22831 252677 22865 253453
rect 22927 252677 22961 253453
rect 23041 252677 23075 253453
rect 23137 252677 23171 253453
rect 23251 252677 23285 253453
rect 23347 252677 23381 253453
rect 23461 252677 23495 253453
rect 23557 252677 23591 253453
rect 23671 252677 23705 253453
rect 23767 252677 23801 253453
rect 23881 252677 23915 253453
rect 23977 252677 24011 253453
rect 24091 252677 24125 253453
rect 24187 252677 24221 253453
rect 24301 252677 24335 253453
rect 24397 252677 24431 253453
rect 24511 252677 24545 253453
rect 24607 252677 24641 253453
rect 24721 252677 24755 253453
rect 24817 252677 24851 253453
rect 24931 252677 24965 253453
rect 25027 252677 25061 253453
rect 25141 252677 25175 253453
rect 25237 252677 25271 253453
rect 25351 252677 25385 253453
rect 25447 252677 25481 253453
rect 25561 252677 25595 253453
rect 25657 252677 25691 253453
rect 25771 252677 25805 253453
rect 25867 252677 25901 253453
rect 25981 252677 26015 253453
rect 26077 252677 26111 253453
rect 26191 252677 26225 253453
rect 26287 252677 26321 253453
rect 26401 252677 26435 253453
rect 26497 252677 26531 253453
rect 26611 252677 26645 253453
rect 26707 252677 26741 253453
rect 26821 252677 26855 253453
rect 26917 252677 26951 253453
rect 27031 252677 27065 253453
rect 27127 252677 27161 253453
rect 27241 252677 27275 253453
rect 27337 252677 27371 253453
rect -4001 252476 -3967 252618
rect -3581 252476 -3547 252618
rect -3161 252476 -3127 252618
rect -2741 252476 -2707 252618
rect -2321 252476 -2287 252618
rect -1901 252476 -1867 252618
rect -1481 252476 -1447 252618
rect -1061 252476 -1027 252618
rect -641 252476 -607 252618
rect -221 252476 -187 252618
rect 199 252476 233 252618
rect 619 252476 653 252618
rect 1039 252476 1073 252618
rect 1459 252476 1493 252618
rect 1879 252476 1913 252618
rect 2299 252476 2333 252618
rect 2719 252476 2753 252618
rect 3139 252476 3173 252618
rect 3559 252476 3593 252618
rect 3979 252476 4013 252618
rect 4399 252476 4433 252618
rect 4819 252476 4853 252618
rect 5239 252476 5273 252618
rect 5659 252476 5693 252618
rect 6079 252476 6113 252618
rect 6499 252476 6533 252618
rect 6919 252476 6953 252618
rect 7339 252476 7373 252618
rect 7759 252476 7793 252618
rect 8179 252476 8213 252618
rect 8599 252476 8633 252618
rect 9019 252476 9053 252618
rect 9439 252476 9473 252618
rect 9859 252476 9893 252618
rect 10279 252476 10313 252618
rect 10699 252476 10733 252618
rect 11119 252476 11153 252618
rect 11539 252476 11573 252618
rect 11959 252476 11993 252618
rect 12379 252476 12413 252618
rect 12799 252476 12833 252618
rect 13219 252476 13253 252618
rect 13639 252476 13673 252618
rect 14059 252476 14093 252618
rect 14479 252476 14513 252618
rect 14899 252476 14933 252618
rect 15319 252476 15353 252618
rect 15739 252476 15773 252618
rect 16159 252476 16193 252618
rect 16579 252476 16613 252618
rect 16999 252476 17033 252618
rect 17419 252476 17453 252618
rect 17839 252476 17873 252618
rect 18259 252476 18293 252618
rect 18679 252476 18713 252618
rect 19099 252476 19133 252618
rect 19519 252476 19553 252618
rect 19939 252476 19973 252618
rect 20359 252476 20393 252618
rect 20779 252476 20813 252618
rect 21199 252476 21233 252618
rect 21619 252476 21653 252618
rect 22039 252476 22073 252618
rect 22459 252476 22493 252618
rect 22879 252476 22913 252618
rect 23299 252476 23333 252618
rect 23719 252476 23753 252618
rect 24139 252476 24173 252618
rect 24559 252476 24593 252618
rect 24979 252476 25013 252618
rect 25399 252476 25433 252618
rect 25819 252476 25853 252618
rect 26239 252476 26273 252618
rect 26659 252476 26693 252618
rect 27079 252476 27113 252618
rect -4049 251641 -4015 252417
rect -3953 251641 -3919 252417
rect -3839 251641 -3805 252417
rect -3743 251641 -3709 252417
rect -3629 251641 -3595 252417
rect -3533 251641 -3499 252417
rect -3419 251641 -3385 252417
rect -3323 251641 -3289 252417
rect -3209 251641 -3175 252417
rect -3113 251641 -3079 252417
rect -2999 251641 -2965 252417
rect -2903 251641 -2869 252417
rect -2789 251641 -2755 252417
rect -2693 251641 -2659 252417
rect -2579 251641 -2545 252417
rect -2483 251641 -2449 252417
rect -2369 251641 -2335 252417
rect -2273 251641 -2239 252417
rect -2159 251641 -2125 252417
rect -2063 251641 -2029 252417
rect -1949 251641 -1915 252417
rect -1853 251641 -1819 252417
rect -1739 251641 -1705 252417
rect -1643 251641 -1609 252417
rect -1529 251641 -1495 252417
rect -1433 251641 -1399 252417
rect -1319 251641 -1285 252417
rect -1223 251641 -1189 252417
rect -1109 251641 -1075 252417
rect -1013 251641 -979 252417
rect -899 251641 -865 252417
rect -803 251641 -769 252417
rect -689 251641 -655 252417
rect -593 251641 -559 252417
rect -479 251641 -445 252417
rect -383 251641 -349 252417
rect -269 251641 -235 252417
rect -173 251641 -139 252417
rect -59 251641 -25 252417
rect 37 251641 71 252417
rect 151 251641 185 252417
rect 247 251641 281 252417
rect 361 251641 395 252417
rect 457 251641 491 252417
rect 571 251641 605 252417
rect 667 251641 701 252417
rect 781 251641 815 252417
rect 877 251641 911 252417
rect 991 251641 1025 252417
rect 1087 251641 1121 252417
rect 1201 251641 1235 252417
rect 1297 251641 1331 252417
rect 1411 251641 1445 252417
rect 1507 251641 1541 252417
rect 1621 251641 1655 252417
rect 1717 251641 1751 252417
rect 1831 251641 1865 252417
rect 1927 251641 1961 252417
rect 2041 251641 2075 252417
rect 2137 251641 2171 252417
rect 2251 251641 2285 252417
rect 2347 251641 2381 252417
rect 2461 251641 2495 252417
rect 2557 251641 2591 252417
rect 2671 251641 2705 252417
rect 2767 251641 2801 252417
rect 2881 251641 2915 252417
rect 2977 251641 3011 252417
rect 3091 251641 3125 252417
rect 3187 251641 3221 252417
rect 3301 251641 3335 252417
rect 3397 251641 3431 252417
rect 3511 251641 3545 252417
rect 3607 251641 3641 252417
rect 3721 251641 3755 252417
rect 3817 251641 3851 252417
rect 3931 251641 3965 252417
rect 4027 251641 4061 252417
rect 4141 251641 4175 252417
rect 4237 251641 4271 252417
rect 4351 251641 4385 252417
rect 4447 251641 4481 252417
rect 4561 251641 4595 252417
rect 4657 251641 4691 252417
rect 4771 251641 4805 252417
rect 4867 251641 4901 252417
rect 4981 251641 5015 252417
rect 5077 251641 5111 252417
rect 5191 251641 5225 252417
rect 5287 251641 5321 252417
rect 5401 251641 5435 252417
rect 5497 251641 5531 252417
rect 5611 251641 5645 252417
rect 5707 251641 5741 252417
rect 5821 251641 5855 252417
rect 5917 251641 5951 252417
rect 6031 251641 6065 252417
rect 6127 251641 6161 252417
rect 6241 251641 6275 252417
rect 6337 251641 6371 252417
rect 6451 251641 6485 252417
rect 6547 251641 6581 252417
rect 6661 251641 6695 252417
rect 6757 251641 6791 252417
rect 6871 251641 6905 252417
rect 6967 251641 7001 252417
rect 7081 251641 7115 252417
rect 7177 251641 7211 252417
rect 7291 251641 7325 252417
rect 7387 251641 7421 252417
rect 7501 251641 7535 252417
rect 7597 251641 7631 252417
rect 7711 251641 7745 252417
rect 7807 251641 7841 252417
rect 7921 251641 7955 252417
rect 8017 251641 8051 252417
rect 8131 251641 8165 252417
rect 8227 251641 8261 252417
rect 8341 251641 8375 252417
rect 8437 251641 8471 252417
rect 8551 251641 8585 252417
rect 8647 251641 8681 252417
rect 8761 251641 8795 252417
rect 8857 251641 8891 252417
rect 8971 251641 9005 252417
rect 9067 251641 9101 252417
rect 9181 251641 9215 252417
rect 9277 251641 9311 252417
rect 9391 251641 9425 252417
rect 9487 251641 9521 252417
rect 9601 251641 9635 252417
rect 9697 251641 9731 252417
rect 9811 251641 9845 252417
rect 9907 251641 9941 252417
rect 10021 251641 10055 252417
rect 10117 251641 10151 252417
rect 10231 251641 10265 252417
rect 10327 251641 10361 252417
rect 10441 251641 10475 252417
rect 10537 251641 10571 252417
rect 10651 251641 10685 252417
rect 10747 251641 10781 252417
rect 10861 251641 10895 252417
rect 10957 251641 10991 252417
rect 11071 251641 11105 252417
rect 11167 251641 11201 252417
rect 11281 251641 11315 252417
rect 11377 251641 11411 252417
rect 11491 251641 11525 252417
rect 11587 251641 11621 252417
rect 11701 251641 11735 252417
rect 11797 251641 11831 252417
rect 11911 251641 11945 252417
rect 12007 251641 12041 252417
rect 12121 251641 12155 252417
rect 12217 251641 12251 252417
rect 12331 251641 12365 252417
rect 12427 251641 12461 252417
rect 12541 251641 12575 252417
rect 12637 251641 12671 252417
rect 12751 251641 12785 252417
rect 12847 251641 12881 252417
rect 12961 251641 12995 252417
rect 13057 251641 13091 252417
rect 13171 251641 13205 252417
rect 13267 251641 13301 252417
rect 13381 251641 13415 252417
rect 13477 251641 13511 252417
rect 13591 251641 13625 252417
rect 13687 251641 13721 252417
rect 13801 251641 13835 252417
rect 13897 251641 13931 252417
rect 14011 251641 14045 252417
rect 14107 251641 14141 252417
rect 14221 251641 14255 252417
rect 14317 251641 14351 252417
rect 14431 251641 14465 252417
rect 14527 251641 14561 252417
rect 14641 251641 14675 252417
rect 14737 251641 14771 252417
rect 14851 251641 14885 252417
rect 14947 251641 14981 252417
rect 15061 251641 15095 252417
rect 15157 251641 15191 252417
rect 15271 251641 15305 252417
rect 15367 251641 15401 252417
rect 15481 251641 15515 252417
rect 15577 251641 15611 252417
rect 15691 251641 15725 252417
rect 15787 251641 15821 252417
rect 15901 251641 15935 252417
rect 15997 251641 16031 252417
rect 16111 251641 16145 252417
rect 16207 251641 16241 252417
rect 16321 251641 16355 252417
rect 16417 251641 16451 252417
rect 16531 251641 16565 252417
rect 16627 251641 16661 252417
rect 16741 251641 16775 252417
rect 16837 251641 16871 252417
rect 16951 251641 16985 252417
rect 17047 251641 17081 252417
rect 17161 251641 17195 252417
rect 17257 251641 17291 252417
rect 17371 251641 17405 252417
rect 17467 251641 17501 252417
rect 17581 251641 17615 252417
rect 17677 251641 17711 252417
rect 17791 251641 17825 252417
rect 17887 251641 17921 252417
rect 18001 251641 18035 252417
rect 18097 251641 18131 252417
rect 18211 251641 18245 252417
rect 18307 251641 18341 252417
rect 18421 251641 18455 252417
rect 18517 251641 18551 252417
rect 18631 251641 18665 252417
rect 18727 251641 18761 252417
rect 18841 251641 18875 252417
rect 18937 251641 18971 252417
rect 19051 251641 19085 252417
rect 19147 251641 19181 252417
rect 19261 251641 19295 252417
rect 19357 251641 19391 252417
rect 19471 251641 19505 252417
rect 19567 251641 19601 252417
rect 19681 251641 19715 252417
rect 19777 251641 19811 252417
rect 19891 251641 19925 252417
rect 19987 251641 20021 252417
rect 20101 251641 20135 252417
rect 20197 251641 20231 252417
rect 20311 251641 20345 252417
rect 20407 251641 20441 252417
rect 20521 251641 20555 252417
rect 20617 251641 20651 252417
rect 20731 251641 20765 252417
rect 20827 251641 20861 252417
rect 20941 251641 20975 252417
rect 21037 251641 21071 252417
rect 21151 251641 21185 252417
rect 21247 251641 21281 252417
rect 21361 251641 21395 252417
rect 21457 251641 21491 252417
rect 21571 251641 21605 252417
rect 21667 251641 21701 252417
rect 21781 251641 21815 252417
rect 21877 251641 21911 252417
rect 21991 251641 22025 252417
rect 22087 251641 22121 252417
rect 22201 251641 22235 252417
rect 22297 251641 22331 252417
rect 22411 251641 22445 252417
rect 22507 251641 22541 252417
rect 22621 251641 22655 252417
rect 22717 251641 22751 252417
rect 22831 251641 22865 252417
rect 22927 251641 22961 252417
rect 23041 251641 23075 252417
rect 23137 251641 23171 252417
rect 23251 251641 23285 252417
rect 23347 251641 23381 252417
rect 23461 251641 23495 252417
rect 23557 251641 23591 252417
rect 23671 251641 23705 252417
rect 23767 251641 23801 252417
rect 23881 251641 23915 252417
rect 23977 251641 24011 252417
rect 24091 251641 24125 252417
rect 24187 251641 24221 252417
rect 24301 251641 24335 252417
rect 24397 251641 24431 252417
rect 24511 251641 24545 252417
rect 24607 251641 24641 252417
rect 24721 251641 24755 252417
rect 24817 251641 24851 252417
rect 24931 251641 24965 252417
rect 25027 251641 25061 252417
rect 25141 251641 25175 252417
rect 25237 251641 25271 252417
rect 25351 251641 25385 252417
rect 25447 251641 25481 252417
rect 25561 251641 25595 252417
rect 25657 251641 25691 252417
rect 25771 251641 25805 252417
rect 25867 251641 25901 252417
rect 25981 251641 26015 252417
rect 26077 251641 26111 252417
rect 26191 251641 26225 252417
rect 26287 251641 26321 252417
rect 26401 251641 26435 252417
rect 26497 251641 26531 252417
rect 26611 251641 26645 252417
rect 26707 251641 26741 252417
rect 26821 251641 26855 252417
rect 26917 251641 26951 252417
rect 27031 251641 27065 252417
rect 27127 251641 27161 252417
rect 27241 251641 27275 252417
rect 27337 251641 27371 252417
rect -3791 251440 -3757 251582
rect -3371 251440 -3337 251582
rect -2951 251440 -2917 251582
rect -2531 251440 -2497 251582
rect -2111 251440 -2077 251582
rect -1691 251440 -1657 251582
rect -1271 251440 -1237 251582
rect -851 251440 -817 251582
rect -431 251440 -397 251582
rect -11 251440 23 251582
rect 409 251440 443 251582
rect 829 251440 863 251582
rect 1249 251440 1283 251582
rect 1669 251440 1703 251582
rect 2089 251440 2123 251582
rect 2509 251440 2543 251582
rect 2929 251440 2963 251582
rect 3349 251440 3383 251582
rect 3769 251440 3803 251582
rect 4189 251440 4223 251582
rect 4609 251440 4643 251582
rect 5029 251440 5063 251582
rect 5449 251440 5483 251582
rect 5869 251440 5903 251582
rect 6289 251440 6323 251582
rect 6709 251440 6743 251582
rect 7129 251440 7163 251582
rect 7549 251440 7583 251582
rect 7969 251440 8003 251582
rect 8389 251440 8423 251582
rect 8809 251440 8843 251582
rect 9229 251440 9263 251582
rect 9649 251440 9683 251582
rect 10069 251440 10103 251582
rect 10489 251440 10523 251582
rect 10909 251440 10943 251582
rect 11329 251440 11363 251582
rect 11749 251440 11783 251582
rect 12169 251440 12203 251582
rect 12589 251440 12623 251582
rect 13009 251440 13043 251582
rect 13429 251440 13463 251582
rect 13849 251440 13883 251582
rect 14269 251440 14303 251582
rect 14689 251440 14723 251582
rect 15109 251440 15143 251582
rect 15529 251440 15563 251582
rect 15949 251440 15983 251582
rect 16369 251440 16403 251582
rect 16789 251440 16823 251582
rect 17209 251440 17243 251582
rect 17629 251440 17663 251582
rect 18049 251440 18083 251582
rect 18469 251440 18503 251582
rect 18889 251440 18923 251582
rect 19309 251440 19343 251582
rect 19729 251440 19763 251582
rect 20149 251440 20183 251582
rect 20569 251440 20603 251582
rect 20989 251440 21023 251582
rect 21409 251440 21443 251582
rect 21829 251440 21863 251582
rect 22249 251440 22283 251582
rect 22669 251440 22703 251582
rect 23089 251440 23123 251582
rect 23509 251440 23543 251582
rect 23929 251440 23963 251582
rect 24349 251440 24383 251582
rect 24769 251440 24803 251582
rect 25189 251440 25223 251582
rect 25609 251440 25643 251582
rect 26029 251440 26063 251582
rect 26449 251440 26483 251582
rect 26869 251440 26903 251582
rect 27289 251440 27323 251582
rect -4049 250605 -4015 251381
rect -3953 250605 -3919 251381
rect -3839 250605 -3805 251381
rect -3743 250605 -3709 251381
rect -3629 250605 -3595 251381
rect -3533 250605 -3499 251381
rect -3419 250605 -3385 251381
rect -3323 250605 -3289 251381
rect -3209 250605 -3175 251381
rect -3113 250605 -3079 251381
rect -2999 250605 -2965 251381
rect -2903 250605 -2869 251381
rect -2789 250605 -2755 251381
rect -2693 250605 -2659 251381
rect -2579 250605 -2545 251381
rect -2483 250605 -2449 251381
rect -2369 250605 -2335 251381
rect -2273 250605 -2239 251381
rect -2159 250605 -2125 251381
rect -2063 250605 -2029 251381
rect -1949 250605 -1915 251381
rect -1853 250605 -1819 251381
rect -1739 250605 -1705 251381
rect -1643 250605 -1609 251381
rect -1529 250605 -1495 251381
rect -1433 250605 -1399 251381
rect -1319 250605 -1285 251381
rect -1223 250605 -1189 251381
rect -1109 250605 -1075 251381
rect -1013 250605 -979 251381
rect -899 250605 -865 251381
rect -803 250605 -769 251381
rect -689 250605 -655 251381
rect -593 250605 -559 251381
rect -479 250605 -445 251381
rect -383 250605 -349 251381
rect -269 250605 -235 251381
rect -173 250605 -139 251381
rect -59 250605 -25 251381
rect 37 250605 71 251381
rect 151 250605 185 251381
rect 247 250605 281 251381
rect 361 250605 395 251381
rect 457 250605 491 251381
rect 571 250605 605 251381
rect 667 250605 701 251381
rect 781 250605 815 251381
rect 877 250605 911 251381
rect 991 250605 1025 251381
rect 1087 250605 1121 251381
rect 1201 250605 1235 251381
rect 1297 250605 1331 251381
rect 1411 250605 1445 251381
rect 1507 250605 1541 251381
rect 1621 250605 1655 251381
rect 1717 250605 1751 251381
rect 1831 250605 1865 251381
rect 1927 250605 1961 251381
rect 2041 250605 2075 251381
rect 2137 250605 2171 251381
rect 2251 250605 2285 251381
rect 2347 250605 2381 251381
rect 2461 250605 2495 251381
rect 2557 250605 2591 251381
rect 2671 250605 2705 251381
rect 2767 250605 2801 251381
rect 2881 250605 2915 251381
rect 2977 250605 3011 251381
rect 3091 250605 3125 251381
rect 3187 250605 3221 251381
rect 3301 250605 3335 251381
rect 3397 250605 3431 251381
rect 3511 250605 3545 251381
rect 3607 250605 3641 251381
rect 3721 250605 3755 251381
rect 3817 250605 3851 251381
rect 3931 250605 3965 251381
rect 4027 250605 4061 251381
rect 4141 250605 4175 251381
rect 4237 250605 4271 251381
rect 4351 250605 4385 251381
rect 4447 250605 4481 251381
rect 4561 250605 4595 251381
rect 4657 250605 4691 251381
rect 4771 250605 4805 251381
rect 4867 250605 4901 251381
rect 4981 250605 5015 251381
rect 5077 250605 5111 251381
rect 5191 250605 5225 251381
rect 5287 250605 5321 251381
rect 5401 250605 5435 251381
rect 5497 250605 5531 251381
rect 5611 250605 5645 251381
rect 5707 250605 5741 251381
rect 5821 250605 5855 251381
rect 5917 250605 5951 251381
rect 6031 250605 6065 251381
rect 6127 250605 6161 251381
rect 6241 250605 6275 251381
rect 6337 250605 6371 251381
rect 6451 250605 6485 251381
rect 6547 250605 6581 251381
rect 6661 250605 6695 251381
rect 6757 250605 6791 251381
rect 6871 250605 6905 251381
rect 6967 250605 7001 251381
rect 7081 250605 7115 251381
rect 7177 250605 7211 251381
rect 7291 250605 7325 251381
rect 7387 250605 7421 251381
rect 7501 250605 7535 251381
rect 7597 250605 7631 251381
rect 7711 250605 7745 251381
rect 7807 250605 7841 251381
rect 7921 250605 7955 251381
rect 8017 250605 8051 251381
rect 8131 250605 8165 251381
rect 8227 250605 8261 251381
rect 8341 250605 8375 251381
rect 8437 250605 8471 251381
rect 8551 250605 8585 251381
rect 8647 250605 8681 251381
rect 8761 250605 8795 251381
rect 8857 250605 8891 251381
rect 8971 250605 9005 251381
rect 9067 250605 9101 251381
rect 9181 250605 9215 251381
rect 9277 250605 9311 251381
rect 9391 250605 9425 251381
rect 9487 250605 9521 251381
rect 9601 250605 9635 251381
rect 9697 250605 9731 251381
rect 9811 250605 9845 251381
rect 9907 250605 9941 251381
rect 10021 250605 10055 251381
rect 10117 250605 10151 251381
rect 10231 250605 10265 251381
rect 10327 250605 10361 251381
rect 10441 250605 10475 251381
rect 10537 250605 10571 251381
rect 10651 250605 10685 251381
rect 10747 250605 10781 251381
rect 10861 250605 10895 251381
rect 10957 250605 10991 251381
rect 11071 250605 11105 251381
rect 11167 250605 11201 251381
rect 11281 250605 11315 251381
rect 11377 250605 11411 251381
rect 11491 250605 11525 251381
rect 11587 250605 11621 251381
rect 11701 250605 11735 251381
rect 11797 250605 11831 251381
rect 11911 250605 11945 251381
rect 12007 250605 12041 251381
rect 12121 250605 12155 251381
rect 12217 250605 12251 251381
rect 12331 250605 12365 251381
rect 12427 250605 12461 251381
rect 12541 250605 12575 251381
rect 12637 250605 12671 251381
rect 12751 250605 12785 251381
rect 12847 250605 12881 251381
rect 12961 250605 12995 251381
rect 13057 250605 13091 251381
rect 13171 250605 13205 251381
rect 13267 250605 13301 251381
rect 13381 250605 13415 251381
rect 13477 250605 13511 251381
rect 13591 250605 13625 251381
rect 13687 250605 13721 251381
rect 13801 250605 13835 251381
rect 13897 250605 13931 251381
rect 14011 250605 14045 251381
rect 14107 250605 14141 251381
rect 14221 250605 14255 251381
rect 14317 250605 14351 251381
rect 14431 250605 14465 251381
rect 14527 250605 14561 251381
rect 14641 250605 14675 251381
rect 14737 250605 14771 251381
rect 14851 250605 14885 251381
rect 14947 250605 14981 251381
rect 15061 250605 15095 251381
rect 15157 250605 15191 251381
rect 15271 250605 15305 251381
rect 15367 250605 15401 251381
rect 15481 250605 15515 251381
rect 15577 250605 15611 251381
rect 15691 250605 15725 251381
rect 15787 250605 15821 251381
rect 15901 250605 15935 251381
rect 15997 250605 16031 251381
rect 16111 250605 16145 251381
rect 16207 250605 16241 251381
rect 16321 250605 16355 251381
rect 16417 250605 16451 251381
rect 16531 250605 16565 251381
rect 16627 250605 16661 251381
rect 16741 250605 16775 251381
rect 16837 250605 16871 251381
rect 16951 250605 16985 251381
rect 17047 250605 17081 251381
rect 17161 250605 17195 251381
rect 17257 250605 17291 251381
rect 17371 250605 17405 251381
rect 17467 250605 17501 251381
rect 17581 250605 17615 251381
rect 17677 250605 17711 251381
rect 17791 250605 17825 251381
rect 17887 250605 17921 251381
rect 18001 250605 18035 251381
rect 18097 250605 18131 251381
rect 18211 250605 18245 251381
rect 18307 250605 18341 251381
rect 18421 250605 18455 251381
rect 18517 250605 18551 251381
rect 18631 250605 18665 251381
rect 18727 250605 18761 251381
rect 18841 250605 18875 251381
rect 18937 250605 18971 251381
rect 19051 250605 19085 251381
rect 19147 250605 19181 251381
rect 19261 250605 19295 251381
rect 19357 250605 19391 251381
rect 19471 250605 19505 251381
rect 19567 250605 19601 251381
rect 19681 250605 19715 251381
rect 19777 250605 19811 251381
rect 19891 250605 19925 251381
rect 19987 250605 20021 251381
rect 20101 250605 20135 251381
rect 20197 250605 20231 251381
rect 20311 250605 20345 251381
rect 20407 250605 20441 251381
rect 20521 250605 20555 251381
rect 20617 250605 20651 251381
rect 20731 250605 20765 251381
rect 20827 250605 20861 251381
rect 20941 250605 20975 251381
rect 21037 250605 21071 251381
rect 21151 250605 21185 251381
rect 21247 250605 21281 251381
rect 21361 250605 21395 251381
rect 21457 250605 21491 251381
rect 21571 250605 21605 251381
rect 21667 250605 21701 251381
rect 21781 250605 21815 251381
rect 21877 250605 21911 251381
rect 21991 250605 22025 251381
rect 22087 250605 22121 251381
rect 22201 250605 22235 251381
rect 22297 250605 22331 251381
rect 22411 250605 22445 251381
rect 22507 250605 22541 251381
rect 22621 250605 22655 251381
rect 22717 250605 22751 251381
rect 22831 250605 22865 251381
rect 22927 250605 22961 251381
rect 23041 250605 23075 251381
rect 23137 250605 23171 251381
rect 23251 250605 23285 251381
rect 23347 250605 23381 251381
rect 23461 250605 23495 251381
rect 23557 250605 23591 251381
rect 23671 250605 23705 251381
rect 23767 250605 23801 251381
rect 23881 250605 23915 251381
rect 23977 250605 24011 251381
rect 24091 250605 24125 251381
rect 24187 250605 24221 251381
rect 24301 250605 24335 251381
rect 24397 250605 24431 251381
rect 24511 250605 24545 251381
rect 24607 250605 24641 251381
rect 24721 250605 24755 251381
rect 24817 250605 24851 251381
rect 24931 250605 24965 251381
rect 25027 250605 25061 251381
rect 25141 250605 25175 251381
rect 25237 250605 25271 251381
rect 25351 250605 25385 251381
rect 25447 250605 25481 251381
rect 25561 250605 25595 251381
rect 25657 250605 25691 251381
rect 25771 250605 25805 251381
rect 25867 250605 25901 251381
rect 25981 250605 26015 251381
rect 26077 250605 26111 251381
rect 26191 250605 26225 251381
rect 26287 250605 26321 251381
rect 26401 250605 26435 251381
rect 26497 250605 26531 251381
rect 26611 250605 26645 251381
rect 26707 250605 26741 251381
rect 26821 250605 26855 251381
rect 26917 250605 26951 251381
rect 27031 250605 27065 251381
rect 27127 250605 27161 251381
rect 27241 250605 27275 251381
rect 27337 250605 27371 251381
rect -4001 250404 -3967 250546
rect -3581 250404 -3547 250546
rect -3161 250404 -3127 250546
rect -2741 250404 -2707 250546
rect -2321 250404 -2287 250546
rect -1901 250404 -1867 250546
rect -1481 250404 -1447 250546
rect -1061 250404 -1027 250546
rect -641 250404 -607 250546
rect -221 250404 -187 250546
rect 199 250404 233 250546
rect 619 250404 653 250546
rect 1039 250404 1073 250546
rect 1459 250404 1493 250546
rect 1879 250404 1913 250546
rect 2299 250404 2333 250546
rect 2719 250404 2753 250546
rect 3139 250404 3173 250546
rect 3559 250404 3593 250546
rect 3979 250404 4013 250546
rect 4399 250404 4433 250546
rect 4819 250404 4853 250546
rect 5239 250404 5273 250546
rect 5659 250404 5693 250546
rect 6079 250404 6113 250546
rect 6499 250404 6533 250546
rect 6919 250404 6953 250546
rect 7339 250404 7373 250546
rect 7759 250404 7793 250546
rect 8179 250404 8213 250546
rect 8599 250404 8633 250546
rect 9019 250404 9053 250546
rect 9439 250404 9473 250546
rect 9859 250404 9893 250546
rect 10279 250404 10313 250546
rect 10699 250404 10733 250546
rect 11119 250404 11153 250546
rect 11539 250404 11573 250546
rect 11959 250404 11993 250546
rect 12379 250404 12413 250546
rect 12799 250404 12833 250546
rect 13219 250404 13253 250546
rect 13639 250404 13673 250546
rect 14059 250404 14093 250546
rect 14479 250404 14513 250546
rect 14899 250404 14933 250546
rect 15319 250404 15353 250546
rect 15739 250404 15773 250546
rect 16159 250404 16193 250546
rect 16579 250404 16613 250546
rect 16999 250404 17033 250546
rect 17419 250404 17453 250546
rect 17839 250404 17873 250546
rect 18259 250404 18293 250546
rect 18679 250404 18713 250546
rect 19099 250404 19133 250546
rect 19519 250404 19553 250546
rect 19939 250404 19973 250546
rect 20359 250404 20393 250546
rect 20779 250404 20813 250546
rect 21199 250404 21233 250546
rect 21619 250404 21653 250546
rect 22039 250404 22073 250546
rect 22459 250404 22493 250546
rect 22879 250404 22913 250546
rect 23299 250404 23333 250546
rect 23719 250404 23753 250546
rect 24139 250404 24173 250546
rect 24559 250404 24593 250546
rect 24979 250404 25013 250546
rect 25399 250404 25433 250546
rect 25819 250404 25853 250546
rect 26239 250404 26273 250546
rect 26659 250404 26693 250546
rect 27079 250404 27113 250546
rect -4049 249569 -4015 250345
rect -3953 249569 -3919 250345
rect -3839 249569 -3805 250345
rect -3743 249569 -3709 250345
rect -3629 249569 -3595 250345
rect -3533 249569 -3499 250345
rect -3419 249569 -3385 250345
rect -3323 249569 -3289 250345
rect -3209 249569 -3175 250345
rect -3113 249569 -3079 250345
rect -2999 249569 -2965 250345
rect -2903 249569 -2869 250345
rect -2789 249569 -2755 250345
rect -2693 249569 -2659 250345
rect -2579 249569 -2545 250345
rect -2483 249569 -2449 250345
rect -2369 249569 -2335 250345
rect -2273 249569 -2239 250345
rect -2159 249569 -2125 250345
rect -2063 249569 -2029 250345
rect -1949 249569 -1915 250345
rect -1853 249569 -1819 250345
rect -1739 249569 -1705 250345
rect -1643 249569 -1609 250345
rect -1529 249569 -1495 250345
rect -1433 249569 -1399 250345
rect -1319 249569 -1285 250345
rect -1223 249569 -1189 250345
rect -1109 249569 -1075 250345
rect -1013 249569 -979 250345
rect -899 249569 -865 250345
rect -803 249569 -769 250345
rect -689 249569 -655 250345
rect -593 249569 -559 250345
rect -479 249569 -445 250345
rect -383 249569 -349 250345
rect -269 249569 -235 250345
rect -173 249569 -139 250345
rect -59 249569 -25 250345
rect 37 249569 71 250345
rect 151 249569 185 250345
rect 247 249569 281 250345
rect 361 249569 395 250345
rect 457 249569 491 250345
rect 571 249569 605 250345
rect 667 249569 701 250345
rect 781 249569 815 250345
rect 877 249569 911 250345
rect 991 249569 1025 250345
rect 1087 249569 1121 250345
rect 1201 249569 1235 250345
rect 1297 249569 1331 250345
rect 1411 249569 1445 250345
rect 1507 249569 1541 250345
rect 1621 249569 1655 250345
rect 1717 249569 1751 250345
rect 1831 249569 1865 250345
rect 1927 249569 1961 250345
rect 2041 249569 2075 250345
rect 2137 249569 2171 250345
rect 2251 249569 2285 250345
rect 2347 249569 2381 250345
rect 2461 249569 2495 250345
rect 2557 249569 2591 250345
rect 2671 249569 2705 250345
rect 2767 249569 2801 250345
rect 2881 249569 2915 250345
rect 2977 249569 3011 250345
rect 3091 249569 3125 250345
rect 3187 249569 3221 250345
rect 3301 249569 3335 250345
rect 3397 249569 3431 250345
rect 3511 249569 3545 250345
rect 3607 249569 3641 250345
rect 3721 249569 3755 250345
rect 3817 249569 3851 250345
rect 3931 249569 3965 250345
rect 4027 249569 4061 250345
rect 4141 249569 4175 250345
rect 4237 249569 4271 250345
rect 4351 249569 4385 250345
rect 4447 249569 4481 250345
rect 4561 249569 4595 250345
rect 4657 249569 4691 250345
rect 4771 249569 4805 250345
rect 4867 249569 4901 250345
rect 4981 249569 5015 250345
rect 5077 249569 5111 250345
rect 5191 249569 5225 250345
rect 5287 249569 5321 250345
rect 5401 249569 5435 250345
rect 5497 249569 5531 250345
rect 5611 249569 5645 250345
rect 5707 249569 5741 250345
rect 5821 249569 5855 250345
rect 5917 249569 5951 250345
rect 6031 249569 6065 250345
rect 6127 249569 6161 250345
rect 6241 249569 6275 250345
rect 6337 249569 6371 250345
rect 6451 249569 6485 250345
rect 6547 249569 6581 250345
rect 6661 249569 6695 250345
rect 6757 249569 6791 250345
rect 6871 249569 6905 250345
rect 6967 249569 7001 250345
rect 7081 249569 7115 250345
rect 7177 249569 7211 250345
rect 7291 249569 7325 250345
rect 7387 249569 7421 250345
rect 7501 249569 7535 250345
rect 7597 249569 7631 250345
rect 7711 249569 7745 250345
rect 7807 249569 7841 250345
rect 7921 249569 7955 250345
rect 8017 249569 8051 250345
rect 8131 249569 8165 250345
rect 8227 249569 8261 250345
rect 8341 249569 8375 250345
rect 8437 249569 8471 250345
rect 8551 249569 8585 250345
rect 8647 249569 8681 250345
rect 8761 249569 8795 250345
rect 8857 249569 8891 250345
rect 8971 249569 9005 250345
rect 9067 249569 9101 250345
rect 9181 249569 9215 250345
rect 9277 249569 9311 250345
rect 9391 249569 9425 250345
rect 9487 249569 9521 250345
rect 9601 249569 9635 250345
rect 9697 249569 9731 250345
rect 9811 249569 9845 250345
rect 9907 249569 9941 250345
rect 10021 249569 10055 250345
rect 10117 249569 10151 250345
rect 10231 249569 10265 250345
rect 10327 249569 10361 250345
rect 10441 249569 10475 250345
rect 10537 249569 10571 250345
rect 10651 249569 10685 250345
rect 10747 249569 10781 250345
rect 10861 249569 10895 250345
rect 10957 249569 10991 250345
rect 11071 249569 11105 250345
rect 11167 249569 11201 250345
rect 11281 249569 11315 250345
rect 11377 249569 11411 250345
rect 11491 249569 11525 250345
rect 11587 249569 11621 250345
rect 11701 249569 11735 250345
rect 11797 249569 11831 250345
rect 11911 249569 11945 250345
rect 12007 249569 12041 250345
rect 12121 249569 12155 250345
rect 12217 249569 12251 250345
rect 12331 249569 12365 250345
rect 12427 249569 12461 250345
rect 12541 249569 12575 250345
rect 12637 249569 12671 250345
rect 12751 249569 12785 250345
rect 12847 249569 12881 250345
rect 12961 249569 12995 250345
rect 13057 249569 13091 250345
rect 13171 249569 13205 250345
rect 13267 249569 13301 250345
rect 13381 249569 13415 250345
rect 13477 249569 13511 250345
rect 13591 249569 13625 250345
rect 13687 249569 13721 250345
rect 13801 249569 13835 250345
rect 13897 249569 13931 250345
rect 14011 249569 14045 250345
rect 14107 249569 14141 250345
rect 14221 249569 14255 250345
rect 14317 249569 14351 250345
rect 14431 249569 14465 250345
rect 14527 249569 14561 250345
rect 14641 249569 14675 250345
rect 14737 249569 14771 250345
rect 14851 249569 14885 250345
rect 14947 249569 14981 250345
rect 15061 249569 15095 250345
rect 15157 249569 15191 250345
rect 15271 249569 15305 250345
rect 15367 249569 15401 250345
rect 15481 249569 15515 250345
rect 15577 249569 15611 250345
rect 15691 249569 15725 250345
rect 15787 249569 15821 250345
rect 15901 249569 15935 250345
rect 15997 249569 16031 250345
rect 16111 249569 16145 250345
rect 16207 249569 16241 250345
rect 16321 249569 16355 250345
rect 16417 249569 16451 250345
rect 16531 249569 16565 250345
rect 16627 249569 16661 250345
rect 16741 249569 16775 250345
rect 16837 249569 16871 250345
rect 16951 249569 16985 250345
rect 17047 249569 17081 250345
rect 17161 249569 17195 250345
rect 17257 249569 17291 250345
rect 17371 249569 17405 250345
rect 17467 249569 17501 250345
rect 17581 249569 17615 250345
rect 17677 249569 17711 250345
rect 17791 249569 17825 250345
rect 17887 249569 17921 250345
rect 18001 249569 18035 250345
rect 18097 249569 18131 250345
rect 18211 249569 18245 250345
rect 18307 249569 18341 250345
rect 18421 249569 18455 250345
rect 18517 249569 18551 250345
rect 18631 249569 18665 250345
rect 18727 249569 18761 250345
rect 18841 249569 18875 250345
rect 18937 249569 18971 250345
rect 19051 249569 19085 250345
rect 19147 249569 19181 250345
rect 19261 249569 19295 250345
rect 19357 249569 19391 250345
rect 19471 249569 19505 250345
rect 19567 249569 19601 250345
rect 19681 249569 19715 250345
rect 19777 249569 19811 250345
rect 19891 249569 19925 250345
rect 19987 249569 20021 250345
rect 20101 249569 20135 250345
rect 20197 249569 20231 250345
rect 20311 249569 20345 250345
rect 20407 249569 20441 250345
rect 20521 249569 20555 250345
rect 20617 249569 20651 250345
rect 20731 249569 20765 250345
rect 20827 249569 20861 250345
rect 20941 249569 20975 250345
rect 21037 249569 21071 250345
rect 21151 249569 21185 250345
rect 21247 249569 21281 250345
rect 21361 249569 21395 250345
rect 21457 249569 21491 250345
rect 21571 249569 21605 250345
rect 21667 249569 21701 250345
rect 21781 249569 21815 250345
rect 21877 249569 21911 250345
rect 21991 249569 22025 250345
rect 22087 249569 22121 250345
rect 22201 249569 22235 250345
rect 22297 249569 22331 250345
rect 22411 249569 22445 250345
rect 22507 249569 22541 250345
rect 22621 249569 22655 250345
rect 22717 249569 22751 250345
rect 22831 249569 22865 250345
rect 22927 249569 22961 250345
rect 23041 249569 23075 250345
rect 23137 249569 23171 250345
rect 23251 249569 23285 250345
rect 23347 249569 23381 250345
rect 23461 249569 23495 250345
rect 23557 249569 23591 250345
rect 23671 249569 23705 250345
rect 23767 249569 23801 250345
rect 23881 249569 23915 250345
rect 23977 249569 24011 250345
rect 24091 249569 24125 250345
rect 24187 249569 24221 250345
rect 24301 249569 24335 250345
rect 24397 249569 24431 250345
rect 24511 249569 24545 250345
rect 24607 249569 24641 250345
rect 24721 249569 24755 250345
rect 24817 249569 24851 250345
rect 24931 249569 24965 250345
rect 25027 249569 25061 250345
rect 25141 249569 25175 250345
rect 25237 249569 25271 250345
rect 25351 249569 25385 250345
rect 25447 249569 25481 250345
rect 25561 249569 25595 250345
rect 25657 249569 25691 250345
rect 25771 249569 25805 250345
rect 25867 249569 25901 250345
rect 25981 249569 26015 250345
rect 26077 249569 26111 250345
rect 26191 249569 26225 250345
rect 26287 249569 26321 250345
rect 26401 249569 26435 250345
rect 26497 249569 26531 250345
rect 26611 249569 26645 250345
rect 26707 249569 26741 250345
rect 26821 249569 26855 250345
rect 26917 249569 26951 250345
rect 27031 249569 27065 250345
rect 27127 249569 27161 250345
rect 27241 249569 27275 250345
rect 27337 249569 27371 250345
rect -3791 249476 -3695 249510
rect -3371 249476 -3275 249510
rect -2951 249476 -2855 249510
rect -2531 249476 -2435 249510
rect -2111 249476 -2015 249510
rect -1691 249476 -1595 249510
rect -1271 249476 -1175 249510
rect -851 249476 -755 249510
rect -431 249476 -335 249510
rect -11 249476 85 249510
rect 409 249476 505 249510
rect 829 249476 925 249510
rect 1249 249476 1345 249510
rect 1669 249476 1765 249510
rect 2089 249476 2185 249510
rect 2509 249476 2605 249510
rect 2929 249476 3025 249510
rect 3349 249476 3445 249510
rect 3769 249476 3865 249510
rect 4189 249476 4285 249510
rect 4609 249476 4705 249510
rect 5029 249476 5125 249510
rect 5449 249476 5545 249510
rect 5869 249476 5965 249510
rect 6289 249476 6385 249510
rect 6709 249476 6805 249510
rect 7129 249476 7225 249510
rect 7549 249476 7645 249510
rect 7969 249476 8065 249510
rect 8389 249476 8485 249510
rect 8809 249476 8905 249510
rect 9229 249476 9325 249510
rect 9649 249476 9745 249510
rect 10069 249476 10165 249510
rect 10489 249476 10585 249510
rect 10909 249476 11005 249510
rect 11329 249476 11425 249510
rect 11749 249476 11845 249510
rect 12169 249476 12265 249510
rect 12589 249476 12685 249510
rect 13009 249476 13105 249510
rect 13429 249476 13525 249510
rect 13849 249476 13945 249510
rect 14269 249476 14365 249510
rect 14689 249476 14785 249510
rect 15109 249476 15205 249510
rect 15529 249476 15625 249510
rect 15949 249476 16045 249510
rect 16369 249476 16465 249510
rect 16789 249476 16885 249510
rect 17209 249476 17305 249510
rect 17629 249476 17725 249510
rect 18049 249476 18145 249510
rect 18469 249476 18565 249510
rect 18889 249476 18985 249510
rect 19309 249476 19405 249510
rect 19729 249476 19825 249510
rect 20149 249476 20245 249510
rect 20569 249476 20665 249510
rect 20989 249476 21085 249510
rect 21409 249476 21505 249510
rect 21829 249476 21925 249510
rect 22249 249476 22345 249510
rect 22669 249476 22765 249510
rect 23089 249476 23185 249510
rect 23509 249476 23605 249510
rect 23929 249476 24025 249510
rect 24349 249476 24445 249510
rect 24769 249476 24865 249510
rect 25189 249476 25285 249510
rect 25609 249476 25705 249510
rect 26029 249476 26125 249510
rect 26449 249476 26545 249510
rect 26869 249476 26965 249510
rect 27289 249476 27385 249510
rect -4001 249239 -3905 249273
rect -3581 249239 -3485 249273
rect -3161 249239 -3065 249273
rect -2741 249239 -2645 249273
rect -2321 249239 -2225 249273
rect -1901 249239 -1805 249273
rect -1481 249239 -1385 249273
rect -1061 249239 -965 249273
rect -641 249239 -545 249273
rect -221 249239 -125 249273
rect 199 249239 295 249273
rect 619 249239 715 249273
rect 1039 249239 1135 249273
rect 1459 249239 1555 249273
rect 1879 249239 1975 249273
rect 2299 249239 2395 249273
rect 2719 249239 2815 249273
rect 3139 249239 3235 249273
rect 3559 249239 3655 249273
rect 3979 249239 4075 249273
rect 4399 249239 4495 249273
rect 4819 249239 4915 249273
rect 5239 249239 5335 249273
rect 5659 249239 5755 249273
rect 6079 249239 6175 249273
rect 6499 249239 6595 249273
rect 6919 249239 7015 249273
rect 7339 249239 7435 249273
rect 7759 249239 7855 249273
rect 8179 249239 8275 249273
rect 8599 249239 8695 249273
rect 9019 249239 9115 249273
rect 9439 249239 9535 249273
rect 9859 249239 9955 249273
rect 10279 249239 10375 249273
rect 10699 249239 10795 249273
rect 11119 249239 11215 249273
rect 11539 249239 11635 249273
rect 11959 249239 12055 249273
rect 12379 249239 12475 249273
rect 12799 249239 12895 249273
rect 13219 249239 13315 249273
rect 13639 249239 13735 249273
rect 14059 249239 14155 249273
rect 14479 249239 14575 249273
rect 14899 249239 14995 249273
rect 15319 249239 15415 249273
rect 15739 249239 15835 249273
rect 16159 249239 16255 249273
rect 16579 249239 16675 249273
rect 16999 249239 17095 249273
rect 17419 249239 17515 249273
rect 17839 249239 17935 249273
rect 18259 249239 18355 249273
rect 18679 249239 18775 249273
rect 19099 249239 19195 249273
rect 19519 249239 19615 249273
rect 19939 249239 20035 249273
rect 20359 249239 20455 249273
rect 20779 249239 20875 249273
rect 21199 249239 21295 249273
rect 21619 249239 21715 249273
rect 22039 249239 22135 249273
rect 22459 249239 22555 249273
rect 22879 249239 22975 249273
rect 23299 249239 23395 249273
rect 23719 249239 23815 249273
rect 24139 249239 24235 249273
rect 24559 249239 24655 249273
rect 24979 249239 25075 249273
rect 25399 249239 25495 249273
rect 25819 249239 25915 249273
rect 26239 249239 26335 249273
rect 26659 249239 26755 249273
rect 27079 249239 27175 249273
rect -4049 248404 -4015 249180
rect -3953 248404 -3919 249180
rect -3839 248404 -3805 249180
rect -3743 248404 -3709 249180
rect -3629 248404 -3595 249180
rect -3533 248404 -3499 249180
rect -3419 248404 -3385 249180
rect -3323 248404 -3289 249180
rect -3209 248404 -3175 249180
rect -3113 248404 -3079 249180
rect -2999 248404 -2965 249180
rect -2903 248404 -2869 249180
rect -2789 248404 -2755 249180
rect -2693 248404 -2659 249180
rect -2579 248404 -2545 249180
rect -2483 248404 -2449 249180
rect -2369 248404 -2335 249180
rect -2273 248404 -2239 249180
rect -2159 248404 -2125 249180
rect -2063 248404 -2029 249180
rect -1949 248404 -1915 249180
rect -1853 248404 -1819 249180
rect -1739 248404 -1705 249180
rect -1643 248404 -1609 249180
rect -1529 248404 -1495 249180
rect -1433 248404 -1399 249180
rect -1319 248404 -1285 249180
rect -1223 248404 -1189 249180
rect -1109 248404 -1075 249180
rect -1013 248404 -979 249180
rect -899 248404 -865 249180
rect -803 248404 -769 249180
rect -689 248404 -655 249180
rect -593 248404 -559 249180
rect -479 248404 -445 249180
rect -383 248404 -349 249180
rect -269 248404 -235 249180
rect -173 248404 -139 249180
rect -59 248404 -25 249180
rect 37 248404 71 249180
rect 151 248404 185 249180
rect 247 248404 281 249180
rect 361 248404 395 249180
rect 457 248404 491 249180
rect 571 248404 605 249180
rect 667 248404 701 249180
rect 781 248404 815 249180
rect 877 248404 911 249180
rect 991 248404 1025 249180
rect 1087 248404 1121 249180
rect 1201 248404 1235 249180
rect 1297 248404 1331 249180
rect 1411 248404 1445 249180
rect 1507 248404 1541 249180
rect 1621 248404 1655 249180
rect 1717 248404 1751 249180
rect 1831 248404 1865 249180
rect 1927 248404 1961 249180
rect 2041 248404 2075 249180
rect 2137 248404 2171 249180
rect 2251 248404 2285 249180
rect 2347 248404 2381 249180
rect 2461 248404 2495 249180
rect 2557 248404 2591 249180
rect 2671 248404 2705 249180
rect 2767 248404 2801 249180
rect 2881 248404 2915 249180
rect 2977 248404 3011 249180
rect 3091 248404 3125 249180
rect 3187 248404 3221 249180
rect 3301 248404 3335 249180
rect 3397 248404 3431 249180
rect 3511 248404 3545 249180
rect 3607 248404 3641 249180
rect 3721 248404 3755 249180
rect 3817 248404 3851 249180
rect 3931 248404 3965 249180
rect 4027 248404 4061 249180
rect 4141 248404 4175 249180
rect 4237 248404 4271 249180
rect 4351 248404 4385 249180
rect 4447 248404 4481 249180
rect 4561 248404 4595 249180
rect 4657 248404 4691 249180
rect 4771 248404 4805 249180
rect 4867 248404 4901 249180
rect 4981 248404 5015 249180
rect 5077 248404 5111 249180
rect 5191 248404 5225 249180
rect 5287 248404 5321 249180
rect 5401 248404 5435 249180
rect 5497 248404 5531 249180
rect 5611 248404 5645 249180
rect 5707 248404 5741 249180
rect 5821 248404 5855 249180
rect 5917 248404 5951 249180
rect 6031 248404 6065 249180
rect 6127 248404 6161 249180
rect 6241 248404 6275 249180
rect 6337 248404 6371 249180
rect 6451 248404 6485 249180
rect 6547 248404 6581 249180
rect 6661 248404 6695 249180
rect 6757 248404 6791 249180
rect 6871 248404 6905 249180
rect 6967 248404 7001 249180
rect 7081 248404 7115 249180
rect 7177 248404 7211 249180
rect 7291 248404 7325 249180
rect 7387 248404 7421 249180
rect 7501 248404 7535 249180
rect 7597 248404 7631 249180
rect 7711 248404 7745 249180
rect 7807 248404 7841 249180
rect 7921 248404 7955 249180
rect 8017 248404 8051 249180
rect 8131 248404 8165 249180
rect 8227 248404 8261 249180
rect 8341 248404 8375 249180
rect 8437 248404 8471 249180
rect 8551 248404 8585 249180
rect 8647 248404 8681 249180
rect 8761 248404 8795 249180
rect 8857 248404 8891 249180
rect 8971 248404 9005 249180
rect 9067 248404 9101 249180
rect 9181 248404 9215 249180
rect 9277 248404 9311 249180
rect 9391 248404 9425 249180
rect 9487 248404 9521 249180
rect 9601 248404 9635 249180
rect 9697 248404 9731 249180
rect 9811 248404 9845 249180
rect 9907 248404 9941 249180
rect 10021 248404 10055 249180
rect 10117 248404 10151 249180
rect 10231 248404 10265 249180
rect 10327 248404 10361 249180
rect 10441 248404 10475 249180
rect 10537 248404 10571 249180
rect 10651 248404 10685 249180
rect 10747 248404 10781 249180
rect 10861 248404 10895 249180
rect 10957 248404 10991 249180
rect 11071 248404 11105 249180
rect 11167 248404 11201 249180
rect 11281 248404 11315 249180
rect 11377 248404 11411 249180
rect 11491 248404 11525 249180
rect 11587 248404 11621 249180
rect 11701 248404 11735 249180
rect 11797 248404 11831 249180
rect 11911 248404 11945 249180
rect 12007 248404 12041 249180
rect 12121 248404 12155 249180
rect 12217 248404 12251 249180
rect 12331 248404 12365 249180
rect 12427 248404 12461 249180
rect 12541 248404 12575 249180
rect 12637 248404 12671 249180
rect 12751 248404 12785 249180
rect 12847 248404 12881 249180
rect 12961 248404 12995 249180
rect 13057 248404 13091 249180
rect 13171 248404 13205 249180
rect 13267 248404 13301 249180
rect 13381 248404 13415 249180
rect 13477 248404 13511 249180
rect 13591 248404 13625 249180
rect 13687 248404 13721 249180
rect 13801 248404 13835 249180
rect 13897 248404 13931 249180
rect 14011 248404 14045 249180
rect 14107 248404 14141 249180
rect 14221 248404 14255 249180
rect 14317 248404 14351 249180
rect 14431 248404 14465 249180
rect 14527 248404 14561 249180
rect 14641 248404 14675 249180
rect 14737 248404 14771 249180
rect 14851 248404 14885 249180
rect 14947 248404 14981 249180
rect 15061 248404 15095 249180
rect 15157 248404 15191 249180
rect 15271 248404 15305 249180
rect 15367 248404 15401 249180
rect 15481 248404 15515 249180
rect 15577 248404 15611 249180
rect 15691 248404 15725 249180
rect 15787 248404 15821 249180
rect 15901 248404 15935 249180
rect 15997 248404 16031 249180
rect 16111 248404 16145 249180
rect 16207 248404 16241 249180
rect 16321 248404 16355 249180
rect 16417 248404 16451 249180
rect 16531 248404 16565 249180
rect 16627 248404 16661 249180
rect 16741 248404 16775 249180
rect 16837 248404 16871 249180
rect 16951 248404 16985 249180
rect 17047 248404 17081 249180
rect 17161 248404 17195 249180
rect 17257 248404 17291 249180
rect 17371 248404 17405 249180
rect 17467 248404 17501 249180
rect 17581 248404 17615 249180
rect 17677 248404 17711 249180
rect 17791 248404 17825 249180
rect 17887 248404 17921 249180
rect 18001 248404 18035 249180
rect 18097 248404 18131 249180
rect 18211 248404 18245 249180
rect 18307 248404 18341 249180
rect 18421 248404 18455 249180
rect 18517 248404 18551 249180
rect 18631 248404 18665 249180
rect 18727 248404 18761 249180
rect 18841 248404 18875 249180
rect 18937 248404 18971 249180
rect 19051 248404 19085 249180
rect 19147 248404 19181 249180
rect 19261 248404 19295 249180
rect 19357 248404 19391 249180
rect 19471 248404 19505 249180
rect 19567 248404 19601 249180
rect 19681 248404 19715 249180
rect 19777 248404 19811 249180
rect 19891 248404 19925 249180
rect 19987 248404 20021 249180
rect 20101 248404 20135 249180
rect 20197 248404 20231 249180
rect 20311 248404 20345 249180
rect 20407 248404 20441 249180
rect 20521 248404 20555 249180
rect 20617 248404 20651 249180
rect 20731 248404 20765 249180
rect 20827 248404 20861 249180
rect 20941 248404 20975 249180
rect 21037 248404 21071 249180
rect 21151 248404 21185 249180
rect 21247 248404 21281 249180
rect 21361 248404 21395 249180
rect 21457 248404 21491 249180
rect 21571 248404 21605 249180
rect 21667 248404 21701 249180
rect 21781 248404 21815 249180
rect 21877 248404 21911 249180
rect 21991 248404 22025 249180
rect 22087 248404 22121 249180
rect 22201 248404 22235 249180
rect 22297 248404 22331 249180
rect 22411 248404 22445 249180
rect 22507 248404 22541 249180
rect 22621 248404 22655 249180
rect 22717 248404 22751 249180
rect 22831 248404 22865 249180
rect 22927 248404 22961 249180
rect 23041 248404 23075 249180
rect 23137 248404 23171 249180
rect 23251 248404 23285 249180
rect 23347 248404 23381 249180
rect 23461 248404 23495 249180
rect 23557 248404 23591 249180
rect 23671 248404 23705 249180
rect 23767 248404 23801 249180
rect 23881 248404 23915 249180
rect 23977 248404 24011 249180
rect 24091 248404 24125 249180
rect 24187 248404 24221 249180
rect 24301 248404 24335 249180
rect 24397 248404 24431 249180
rect 24511 248404 24545 249180
rect 24607 248404 24641 249180
rect 24721 248404 24755 249180
rect 24817 248404 24851 249180
rect 24931 248404 24965 249180
rect 25027 248404 25061 249180
rect 25141 248404 25175 249180
rect 25237 248404 25271 249180
rect 25351 248404 25385 249180
rect 25447 248404 25481 249180
rect 25561 248404 25595 249180
rect 25657 248404 25691 249180
rect 25771 248404 25805 249180
rect 25867 248404 25901 249180
rect 25981 248404 26015 249180
rect 26077 248404 26111 249180
rect 26191 248404 26225 249180
rect 26287 248404 26321 249180
rect 26401 248404 26435 249180
rect 26497 248404 26531 249180
rect 26611 248404 26645 249180
rect 26707 248404 26741 249180
rect 26821 248404 26855 249180
rect 26917 248404 26951 249180
rect 27031 248404 27065 249180
rect 27127 248404 27161 249180
rect 27241 248404 27275 249180
rect 27337 248404 27371 249180
rect -3791 248203 -3757 248345
rect -3371 248203 -3337 248345
rect -2951 248203 -2917 248345
rect -2531 248203 -2497 248345
rect -2111 248203 -2077 248345
rect -1691 248203 -1657 248345
rect -1271 248203 -1237 248345
rect -851 248203 -817 248345
rect -431 248203 -397 248345
rect -11 248203 23 248345
rect 409 248203 443 248345
rect 829 248203 863 248345
rect 1249 248203 1283 248345
rect 1669 248203 1703 248345
rect 2089 248203 2123 248345
rect 2509 248203 2543 248345
rect 2929 248203 2963 248345
rect 3349 248203 3383 248345
rect 3769 248203 3803 248345
rect 4189 248203 4223 248345
rect 4609 248203 4643 248345
rect 5029 248203 5063 248345
rect 5449 248203 5483 248345
rect 5869 248203 5903 248345
rect 6289 248203 6323 248345
rect 6709 248203 6743 248345
rect 7129 248203 7163 248345
rect 7549 248203 7583 248345
rect 7969 248203 8003 248345
rect 8389 248203 8423 248345
rect 8809 248203 8843 248345
rect 9229 248203 9263 248345
rect 9649 248203 9683 248345
rect 10069 248203 10103 248345
rect 10489 248203 10523 248345
rect 10909 248203 10943 248345
rect 11329 248203 11363 248345
rect 11749 248203 11783 248345
rect 12169 248203 12203 248345
rect 12589 248203 12623 248345
rect 13009 248203 13043 248345
rect 13429 248203 13463 248345
rect 13849 248203 13883 248345
rect 14269 248203 14303 248345
rect 14689 248203 14723 248345
rect 15109 248203 15143 248345
rect 15529 248203 15563 248345
rect 15949 248203 15983 248345
rect 16369 248203 16403 248345
rect 16789 248203 16823 248345
rect 17209 248203 17243 248345
rect 17629 248203 17663 248345
rect 18049 248203 18083 248345
rect 18469 248203 18503 248345
rect 18889 248203 18923 248345
rect 19309 248203 19343 248345
rect 19729 248203 19763 248345
rect 20149 248203 20183 248345
rect 20569 248203 20603 248345
rect 20989 248203 21023 248345
rect 21409 248203 21443 248345
rect 21829 248203 21863 248345
rect 22249 248203 22283 248345
rect 22669 248203 22703 248345
rect 23089 248203 23123 248345
rect 23509 248203 23543 248345
rect 23929 248203 23963 248345
rect 24349 248203 24383 248345
rect 24769 248203 24803 248345
rect 25189 248203 25223 248345
rect 25609 248203 25643 248345
rect 26029 248203 26063 248345
rect 26449 248203 26483 248345
rect 26869 248203 26903 248345
rect 27289 248203 27323 248345
rect -4049 247368 -4015 248144
rect -3953 247368 -3919 248144
rect -3839 247368 -3805 248144
rect -3743 247368 -3709 248144
rect -3629 247368 -3595 248144
rect -3533 247368 -3499 248144
rect -3419 247368 -3385 248144
rect -3323 247368 -3289 248144
rect -3209 247368 -3175 248144
rect -3113 247368 -3079 248144
rect -2999 247368 -2965 248144
rect -2903 247368 -2869 248144
rect -2789 247368 -2755 248144
rect -2693 247368 -2659 248144
rect -2579 247368 -2545 248144
rect -2483 247368 -2449 248144
rect -2369 247368 -2335 248144
rect -2273 247368 -2239 248144
rect -2159 247368 -2125 248144
rect -2063 247368 -2029 248144
rect -1949 247368 -1915 248144
rect -1853 247368 -1819 248144
rect -1739 247368 -1705 248144
rect -1643 247368 -1609 248144
rect -1529 247368 -1495 248144
rect -1433 247368 -1399 248144
rect -1319 247368 -1285 248144
rect -1223 247368 -1189 248144
rect -1109 247368 -1075 248144
rect -1013 247368 -979 248144
rect -899 247368 -865 248144
rect -803 247368 -769 248144
rect -689 247368 -655 248144
rect -593 247368 -559 248144
rect -479 247368 -445 248144
rect -383 247368 -349 248144
rect -269 247368 -235 248144
rect -173 247368 -139 248144
rect -59 247368 -25 248144
rect 37 247368 71 248144
rect 151 247368 185 248144
rect 247 247368 281 248144
rect 361 247368 395 248144
rect 457 247368 491 248144
rect 571 247368 605 248144
rect 667 247368 701 248144
rect 781 247368 815 248144
rect 877 247368 911 248144
rect 991 247368 1025 248144
rect 1087 247368 1121 248144
rect 1201 247368 1235 248144
rect 1297 247368 1331 248144
rect 1411 247368 1445 248144
rect 1507 247368 1541 248144
rect 1621 247368 1655 248144
rect 1717 247368 1751 248144
rect 1831 247368 1865 248144
rect 1927 247368 1961 248144
rect 2041 247368 2075 248144
rect 2137 247368 2171 248144
rect 2251 247368 2285 248144
rect 2347 247368 2381 248144
rect 2461 247368 2495 248144
rect 2557 247368 2591 248144
rect 2671 247368 2705 248144
rect 2767 247368 2801 248144
rect 2881 247368 2915 248144
rect 2977 247368 3011 248144
rect 3091 247368 3125 248144
rect 3187 247368 3221 248144
rect 3301 247368 3335 248144
rect 3397 247368 3431 248144
rect 3511 247368 3545 248144
rect 3607 247368 3641 248144
rect 3721 247368 3755 248144
rect 3817 247368 3851 248144
rect 3931 247368 3965 248144
rect 4027 247368 4061 248144
rect 4141 247368 4175 248144
rect 4237 247368 4271 248144
rect 4351 247368 4385 248144
rect 4447 247368 4481 248144
rect 4561 247368 4595 248144
rect 4657 247368 4691 248144
rect 4771 247368 4805 248144
rect 4867 247368 4901 248144
rect 4981 247368 5015 248144
rect 5077 247368 5111 248144
rect 5191 247368 5225 248144
rect 5287 247368 5321 248144
rect 5401 247368 5435 248144
rect 5497 247368 5531 248144
rect 5611 247368 5645 248144
rect 5707 247368 5741 248144
rect 5821 247368 5855 248144
rect 5917 247368 5951 248144
rect 6031 247368 6065 248144
rect 6127 247368 6161 248144
rect 6241 247368 6275 248144
rect 6337 247368 6371 248144
rect 6451 247368 6485 248144
rect 6547 247368 6581 248144
rect 6661 247368 6695 248144
rect 6757 247368 6791 248144
rect 6871 247368 6905 248144
rect 6967 247368 7001 248144
rect 7081 247368 7115 248144
rect 7177 247368 7211 248144
rect 7291 247368 7325 248144
rect 7387 247368 7421 248144
rect 7501 247368 7535 248144
rect 7597 247368 7631 248144
rect 7711 247368 7745 248144
rect 7807 247368 7841 248144
rect 7921 247368 7955 248144
rect 8017 247368 8051 248144
rect 8131 247368 8165 248144
rect 8227 247368 8261 248144
rect 8341 247368 8375 248144
rect 8437 247368 8471 248144
rect 8551 247368 8585 248144
rect 8647 247368 8681 248144
rect 8761 247368 8795 248144
rect 8857 247368 8891 248144
rect 8971 247368 9005 248144
rect 9067 247368 9101 248144
rect 9181 247368 9215 248144
rect 9277 247368 9311 248144
rect 9391 247368 9425 248144
rect 9487 247368 9521 248144
rect 9601 247368 9635 248144
rect 9697 247368 9731 248144
rect 9811 247368 9845 248144
rect 9907 247368 9941 248144
rect 10021 247368 10055 248144
rect 10117 247368 10151 248144
rect 10231 247368 10265 248144
rect 10327 247368 10361 248144
rect 10441 247368 10475 248144
rect 10537 247368 10571 248144
rect 10651 247368 10685 248144
rect 10747 247368 10781 248144
rect 10861 247368 10895 248144
rect 10957 247368 10991 248144
rect 11071 247368 11105 248144
rect 11167 247368 11201 248144
rect 11281 247368 11315 248144
rect 11377 247368 11411 248144
rect 11491 247368 11525 248144
rect 11587 247368 11621 248144
rect 11701 247368 11735 248144
rect 11797 247368 11831 248144
rect 11911 247368 11945 248144
rect 12007 247368 12041 248144
rect 12121 247368 12155 248144
rect 12217 247368 12251 248144
rect 12331 247368 12365 248144
rect 12427 247368 12461 248144
rect 12541 247368 12575 248144
rect 12637 247368 12671 248144
rect 12751 247368 12785 248144
rect 12847 247368 12881 248144
rect 12961 247368 12995 248144
rect 13057 247368 13091 248144
rect 13171 247368 13205 248144
rect 13267 247368 13301 248144
rect 13381 247368 13415 248144
rect 13477 247368 13511 248144
rect 13591 247368 13625 248144
rect 13687 247368 13721 248144
rect 13801 247368 13835 248144
rect 13897 247368 13931 248144
rect 14011 247368 14045 248144
rect 14107 247368 14141 248144
rect 14221 247368 14255 248144
rect 14317 247368 14351 248144
rect 14431 247368 14465 248144
rect 14527 247368 14561 248144
rect 14641 247368 14675 248144
rect 14737 247368 14771 248144
rect 14851 247368 14885 248144
rect 14947 247368 14981 248144
rect 15061 247368 15095 248144
rect 15157 247368 15191 248144
rect 15271 247368 15305 248144
rect 15367 247368 15401 248144
rect 15481 247368 15515 248144
rect 15577 247368 15611 248144
rect 15691 247368 15725 248144
rect 15787 247368 15821 248144
rect 15901 247368 15935 248144
rect 15997 247368 16031 248144
rect 16111 247368 16145 248144
rect 16207 247368 16241 248144
rect 16321 247368 16355 248144
rect 16417 247368 16451 248144
rect 16531 247368 16565 248144
rect 16627 247368 16661 248144
rect 16741 247368 16775 248144
rect 16837 247368 16871 248144
rect 16951 247368 16985 248144
rect 17047 247368 17081 248144
rect 17161 247368 17195 248144
rect 17257 247368 17291 248144
rect 17371 247368 17405 248144
rect 17467 247368 17501 248144
rect 17581 247368 17615 248144
rect 17677 247368 17711 248144
rect 17791 247368 17825 248144
rect 17887 247368 17921 248144
rect 18001 247368 18035 248144
rect 18097 247368 18131 248144
rect 18211 247368 18245 248144
rect 18307 247368 18341 248144
rect 18421 247368 18455 248144
rect 18517 247368 18551 248144
rect 18631 247368 18665 248144
rect 18727 247368 18761 248144
rect 18841 247368 18875 248144
rect 18937 247368 18971 248144
rect 19051 247368 19085 248144
rect 19147 247368 19181 248144
rect 19261 247368 19295 248144
rect 19357 247368 19391 248144
rect 19471 247368 19505 248144
rect 19567 247368 19601 248144
rect 19681 247368 19715 248144
rect 19777 247368 19811 248144
rect 19891 247368 19925 248144
rect 19987 247368 20021 248144
rect 20101 247368 20135 248144
rect 20197 247368 20231 248144
rect 20311 247368 20345 248144
rect 20407 247368 20441 248144
rect 20521 247368 20555 248144
rect 20617 247368 20651 248144
rect 20731 247368 20765 248144
rect 20827 247368 20861 248144
rect 20941 247368 20975 248144
rect 21037 247368 21071 248144
rect 21151 247368 21185 248144
rect 21247 247368 21281 248144
rect 21361 247368 21395 248144
rect 21457 247368 21491 248144
rect 21571 247368 21605 248144
rect 21667 247368 21701 248144
rect 21781 247368 21815 248144
rect 21877 247368 21911 248144
rect 21991 247368 22025 248144
rect 22087 247368 22121 248144
rect 22201 247368 22235 248144
rect 22297 247368 22331 248144
rect 22411 247368 22445 248144
rect 22507 247368 22541 248144
rect 22621 247368 22655 248144
rect 22717 247368 22751 248144
rect 22831 247368 22865 248144
rect 22927 247368 22961 248144
rect 23041 247368 23075 248144
rect 23137 247368 23171 248144
rect 23251 247368 23285 248144
rect 23347 247368 23381 248144
rect 23461 247368 23495 248144
rect 23557 247368 23591 248144
rect 23671 247368 23705 248144
rect 23767 247368 23801 248144
rect 23881 247368 23915 248144
rect 23977 247368 24011 248144
rect 24091 247368 24125 248144
rect 24187 247368 24221 248144
rect 24301 247368 24335 248144
rect 24397 247368 24431 248144
rect 24511 247368 24545 248144
rect 24607 247368 24641 248144
rect 24721 247368 24755 248144
rect 24817 247368 24851 248144
rect 24931 247368 24965 248144
rect 25027 247368 25061 248144
rect 25141 247368 25175 248144
rect 25237 247368 25271 248144
rect 25351 247368 25385 248144
rect 25447 247368 25481 248144
rect 25561 247368 25595 248144
rect 25657 247368 25691 248144
rect 25771 247368 25805 248144
rect 25867 247368 25901 248144
rect 25981 247368 26015 248144
rect 26077 247368 26111 248144
rect 26191 247368 26225 248144
rect 26287 247368 26321 248144
rect 26401 247368 26435 248144
rect 26497 247368 26531 248144
rect 26611 247368 26645 248144
rect 26707 247368 26741 248144
rect 26821 247368 26855 248144
rect 26917 247368 26951 248144
rect 27031 247368 27065 248144
rect 27127 247368 27161 248144
rect 27241 247368 27275 248144
rect 27337 247368 27371 248144
rect -4001 247167 -3967 247309
rect -3581 247167 -3547 247309
rect -3161 247167 -3127 247309
rect -2741 247167 -2707 247309
rect -2321 247167 -2287 247309
rect -1901 247167 -1867 247309
rect -1481 247167 -1447 247309
rect -1061 247167 -1027 247309
rect -641 247167 -607 247309
rect -221 247167 -187 247309
rect 199 247167 233 247309
rect 619 247167 653 247309
rect 1039 247167 1073 247309
rect 1459 247167 1493 247309
rect 1879 247167 1913 247309
rect 2299 247167 2333 247309
rect 2719 247167 2753 247309
rect 3139 247167 3173 247309
rect 3559 247167 3593 247309
rect 3979 247167 4013 247309
rect 4399 247167 4433 247309
rect 4819 247167 4853 247309
rect 5239 247167 5273 247309
rect 5659 247167 5693 247309
rect 6079 247167 6113 247309
rect 6499 247167 6533 247309
rect 6919 247167 6953 247309
rect 7339 247167 7373 247309
rect 7759 247167 7793 247309
rect 8179 247167 8213 247309
rect 8599 247167 8633 247309
rect 9019 247167 9053 247309
rect 9439 247167 9473 247309
rect 9859 247167 9893 247309
rect 10279 247167 10313 247309
rect 10699 247167 10733 247309
rect 11119 247167 11153 247309
rect 11539 247167 11573 247309
rect 11959 247167 11993 247309
rect 12379 247167 12413 247309
rect 12799 247167 12833 247309
rect 13219 247167 13253 247309
rect 13639 247167 13673 247309
rect 14059 247167 14093 247309
rect 14479 247167 14513 247309
rect 14899 247167 14933 247309
rect 15319 247167 15353 247309
rect 15739 247167 15773 247309
rect 16159 247167 16193 247309
rect 16579 247167 16613 247309
rect 16999 247167 17033 247309
rect 17419 247167 17453 247309
rect 17839 247167 17873 247309
rect 18259 247167 18293 247309
rect 18679 247167 18713 247309
rect 19099 247167 19133 247309
rect 19519 247167 19553 247309
rect 19939 247167 19973 247309
rect 20359 247167 20393 247309
rect 20779 247167 20813 247309
rect 21199 247167 21233 247309
rect 21619 247167 21653 247309
rect 22039 247167 22073 247309
rect 22459 247167 22493 247309
rect 22879 247167 22913 247309
rect 23299 247167 23333 247309
rect 23719 247167 23753 247309
rect 24139 247167 24173 247309
rect 24559 247167 24593 247309
rect 24979 247167 25013 247309
rect 25399 247167 25433 247309
rect 25819 247167 25853 247309
rect 26239 247167 26273 247309
rect 26659 247167 26693 247309
rect 27079 247167 27113 247309
rect -4049 246332 -4015 247108
rect -3953 246332 -3919 247108
rect -3839 246332 -3805 247108
rect -3743 246332 -3709 247108
rect -3629 246332 -3595 247108
rect -3533 246332 -3499 247108
rect -3419 246332 -3385 247108
rect -3323 246332 -3289 247108
rect -3209 246332 -3175 247108
rect -3113 246332 -3079 247108
rect -2999 246332 -2965 247108
rect -2903 246332 -2869 247108
rect -2789 246332 -2755 247108
rect -2693 246332 -2659 247108
rect -2579 246332 -2545 247108
rect -2483 246332 -2449 247108
rect -2369 246332 -2335 247108
rect -2273 246332 -2239 247108
rect -2159 246332 -2125 247108
rect -2063 246332 -2029 247108
rect -1949 246332 -1915 247108
rect -1853 246332 -1819 247108
rect -1739 246332 -1705 247108
rect -1643 246332 -1609 247108
rect -1529 246332 -1495 247108
rect -1433 246332 -1399 247108
rect -1319 246332 -1285 247108
rect -1223 246332 -1189 247108
rect -1109 246332 -1075 247108
rect -1013 246332 -979 247108
rect -899 246332 -865 247108
rect -803 246332 -769 247108
rect -689 246332 -655 247108
rect -593 246332 -559 247108
rect -479 246332 -445 247108
rect -383 246332 -349 247108
rect -269 246332 -235 247108
rect -173 246332 -139 247108
rect -59 246332 -25 247108
rect 37 246332 71 247108
rect 151 246332 185 247108
rect 247 246332 281 247108
rect 361 246332 395 247108
rect 457 246332 491 247108
rect 571 246332 605 247108
rect 667 246332 701 247108
rect 781 246332 815 247108
rect 877 246332 911 247108
rect 991 246332 1025 247108
rect 1087 246332 1121 247108
rect 1201 246332 1235 247108
rect 1297 246332 1331 247108
rect 1411 246332 1445 247108
rect 1507 246332 1541 247108
rect 1621 246332 1655 247108
rect 1717 246332 1751 247108
rect 1831 246332 1865 247108
rect 1927 246332 1961 247108
rect 2041 246332 2075 247108
rect 2137 246332 2171 247108
rect 2251 246332 2285 247108
rect 2347 246332 2381 247108
rect 2461 246332 2495 247108
rect 2557 246332 2591 247108
rect 2671 246332 2705 247108
rect 2767 246332 2801 247108
rect 2881 246332 2915 247108
rect 2977 246332 3011 247108
rect 3091 246332 3125 247108
rect 3187 246332 3221 247108
rect 3301 246332 3335 247108
rect 3397 246332 3431 247108
rect 3511 246332 3545 247108
rect 3607 246332 3641 247108
rect 3721 246332 3755 247108
rect 3817 246332 3851 247108
rect 3931 246332 3965 247108
rect 4027 246332 4061 247108
rect 4141 246332 4175 247108
rect 4237 246332 4271 247108
rect 4351 246332 4385 247108
rect 4447 246332 4481 247108
rect 4561 246332 4595 247108
rect 4657 246332 4691 247108
rect 4771 246332 4805 247108
rect 4867 246332 4901 247108
rect 4981 246332 5015 247108
rect 5077 246332 5111 247108
rect 5191 246332 5225 247108
rect 5287 246332 5321 247108
rect 5401 246332 5435 247108
rect 5497 246332 5531 247108
rect 5611 246332 5645 247108
rect 5707 246332 5741 247108
rect 5821 246332 5855 247108
rect 5917 246332 5951 247108
rect 6031 246332 6065 247108
rect 6127 246332 6161 247108
rect 6241 246332 6275 247108
rect 6337 246332 6371 247108
rect 6451 246332 6485 247108
rect 6547 246332 6581 247108
rect 6661 246332 6695 247108
rect 6757 246332 6791 247108
rect 6871 246332 6905 247108
rect 6967 246332 7001 247108
rect 7081 246332 7115 247108
rect 7177 246332 7211 247108
rect 7291 246332 7325 247108
rect 7387 246332 7421 247108
rect 7501 246332 7535 247108
rect 7597 246332 7631 247108
rect 7711 246332 7745 247108
rect 7807 246332 7841 247108
rect 7921 246332 7955 247108
rect 8017 246332 8051 247108
rect 8131 246332 8165 247108
rect 8227 246332 8261 247108
rect 8341 246332 8375 247108
rect 8437 246332 8471 247108
rect 8551 246332 8585 247108
rect 8647 246332 8681 247108
rect 8761 246332 8795 247108
rect 8857 246332 8891 247108
rect 8971 246332 9005 247108
rect 9067 246332 9101 247108
rect 9181 246332 9215 247108
rect 9277 246332 9311 247108
rect 9391 246332 9425 247108
rect 9487 246332 9521 247108
rect 9601 246332 9635 247108
rect 9697 246332 9731 247108
rect 9811 246332 9845 247108
rect 9907 246332 9941 247108
rect 10021 246332 10055 247108
rect 10117 246332 10151 247108
rect 10231 246332 10265 247108
rect 10327 246332 10361 247108
rect 10441 246332 10475 247108
rect 10537 246332 10571 247108
rect 10651 246332 10685 247108
rect 10747 246332 10781 247108
rect 10861 246332 10895 247108
rect 10957 246332 10991 247108
rect 11071 246332 11105 247108
rect 11167 246332 11201 247108
rect 11281 246332 11315 247108
rect 11377 246332 11411 247108
rect 11491 246332 11525 247108
rect 11587 246332 11621 247108
rect 11701 246332 11735 247108
rect 11797 246332 11831 247108
rect 11911 246332 11945 247108
rect 12007 246332 12041 247108
rect 12121 246332 12155 247108
rect 12217 246332 12251 247108
rect 12331 246332 12365 247108
rect 12427 246332 12461 247108
rect 12541 246332 12575 247108
rect 12637 246332 12671 247108
rect 12751 246332 12785 247108
rect 12847 246332 12881 247108
rect 12961 246332 12995 247108
rect 13057 246332 13091 247108
rect 13171 246332 13205 247108
rect 13267 246332 13301 247108
rect 13381 246332 13415 247108
rect 13477 246332 13511 247108
rect 13591 246332 13625 247108
rect 13687 246332 13721 247108
rect 13801 246332 13835 247108
rect 13897 246332 13931 247108
rect 14011 246332 14045 247108
rect 14107 246332 14141 247108
rect 14221 246332 14255 247108
rect 14317 246332 14351 247108
rect 14431 246332 14465 247108
rect 14527 246332 14561 247108
rect 14641 246332 14675 247108
rect 14737 246332 14771 247108
rect 14851 246332 14885 247108
rect 14947 246332 14981 247108
rect 15061 246332 15095 247108
rect 15157 246332 15191 247108
rect 15271 246332 15305 247108
rect 15367 246332 15401 247108
rect 15481 246332 15515 247108
rect 15577 246332 15611 247108
rect 15691 246332 15725 247108
rect 15787 246332 15821 247108
rect 15901 246332 15935 247108
rect 15997 246332 16031 247108
rect 16111 246332 16145 247108
rect 16207 246332 16241 247108
rect 16321 246332 16355 247108
rect 16417 246332 16451 247108
rect 16531 246332 16565 247108
rect 16627 246332 16661 247108
rect 16741 246332 16775 247108
rect 16837 246332 16871 247108
rect 16951 246332 16985 247108
rect 17047 246332 17081 247108
rect 17161 246332 17195 247108
rect 17257 246332 17291 247108
rect 17371 246332 17405 247108
rect 17467 246332 17501 247108
rect 17581 246332 17615 247108
rect 17677 246332 17711 247108
rect 17791 246332 17825 247108
rect 17887 246332 17921 247108
rect 18001 246332 18035 247108
rect 18097 246332 18131 247108
rect 18211 246332 18245 247108
rect 18307 246332 18341 247108
rect 18421 246332 18455 247108
rect 18517 246332 18551 247108
rect 18631 246332 18665 247108
rect 18727 246332 18761 247108
rect 18841 246332 18875 247108
rect 18937 246332 18971 247108
rect 19051 246332 19085 247108
rect 19147 246332 19181 247108
rect 19261 246332 19295 247108
rect 19357 246332 19391 247108
rect 19471 246332 19505 247108
rect 19567 246332 19601 247108
rect 19681 246332 19715 247108
rect 19777 246332 19811 247108
rect 19891 246332 19925 247108
rect 19987 246332 20021 247108
rect 20101 246332 20135 247108
rect 20197 246332 20231 247108
rect 20311 246332 20345 247108
rect 20407 246332 20441 247108
rect 20521 246332 20555 247108
rect 20617 246332 20651 247108
rect 20731 246332 20765 247108
rect 20827 246332 20861 247108
rect 20941 246332 20975 247108
rect 21037 246332 21071 247108
rect 21151 246332 21185 247108
rect 21247 246332 21281 247108
rect 21361 246332 21395 247108
rect 21457 246332 21491 247108
rect 21571 246332 21605 247108
rect 21667 246332 21701 247108
rect 21781 246332 21815 247108
rect 21877 246332 21911 247108
rect 21991 246332 22025 247108
rect 22087 246332 22121 247108
rect 22201 246332 22235 247108
rect 22297 246332 22331 247108
rect 22411 246332 22445 247108
rect 22507 246332 22541 247108
rect 22621 246332 22655 247108
rect 22717 246332 22751 247108
rect 22831 246332 22865 247108
rect 22927 246332 22961 247108
rect 23041 246332 23075 247108
rect 23137 246332 23171 247108
rect 23251 246332 23285 247108
rect 23347 246332 23381 247108
rect 23461 246332 23495 247108
rect 23557 246332 23591 247108
rect 23671 246332 23705 247108
rect 23767 246332 23801 247108
rect 23881 246332 23915 247108
rect 23977 246332 24011 247108
rect 24091 246332 24125 247108
rect 24187 246332 24221 247108
rect 24301 246332 24335 247108
rect 24397 246332 24431 247108
rect 24511 246332 24545 247108
rect 24607 246332 24641 247108
rect 24721 246332 24755 247108
rect 24817 246332 24851 247108
rect 24931 246332 24965 247108
rect 25027 246332 25061 247108
rect 25141 246332 25175 247108
rect 25237 246332 25271 247108
rect 25351 246332 25385 247108
rect 25447 246332 25481 247108
rect 25561 246332 25595 247108
rect 25657 246332 25691 247108
rect 25771 246332 25805 247108
rect 25867 246332 25901 247108
rect 25981 246332 26015 247108
rect 26077 246332 26111 247108
rect 26191 246332 26225 247108
rect 26287 246332 26321 247108
rect 26401 246332 26435 247108
rect 26497 246332 26531 247108
rect 26611 246332 26645 247108
rect 26707 246332 26741 247108
rect 26821 246332 26855 247108
rect 26917 246332 26951 247108
rect 27031 246332 27065 247108
rect 27127 246332 27161 247108
rect 27241 246332 27275 247108
rect 27337 246332 27371 247108
rect -3791 246131 -3757 246273
rect -3371 246131 -3337 246273
rect -2951 246131 -2917 246273
rect -2531 246131 -2497 246273
rect -2111 246131 -2077 246273
rect -1691 246131 -1657 246273
rect -1271 246131 -1237 246273
rect -851 246131 -817 246273
rect -431 246131 -397 246273
rect -11 246131 23 246273
rect 409 246131 443 246273
rect 829 246131 863 246273
rect 1249 246131 1283 246273
rect 1669 246131 1703 246273
rect 2089 246131 2123 246273
rect 2509 246131 2543 246273
rect 2929 246131 2963 246273
rect 3349 246131 3383 246273
rect 3769 246131 3803 246273
rect 4189 246131 4223 246273
rect 4609 246131 4643 246273
rect 5029 246131 5063 246273
rect 5449 246131 5483 246273
rect 5869 246131 5903 246273
rect 6289 246131 6323 246273
rect 6709 246131 6743 246273
rect 7129 246131 7163 246273
rect 7549 246131 7583 246273
rect 7969 246131 8003 246273
rect 8389 246131 8423 246273
rect 8809 246131 8843 246273
rect 9229 246131 9263 246273
rect 9649 246131 9683 246273
rect 10069 246131 10103 246273
rect 10489 246131 10523 246273
rect 10909 246131 10943 246273
rect 11329 246131 11363 246273
rect 11749 246131 11783 246273
rect 12169 246131 12203 246273
rect 12589 246131 12623 246273
rect 13009 246131 13043 246273
rect 13429 246131 13463 246273
rect 13849 246131 13883 246273
rect 14269 246131 14303 246273
rect 14689 246131 14723 246273
rect 15109 246131 15143 246273
rect 15529 246131 15563 246273
rect 15949 246131 15983 246273
rect 16369 246131 16403 246273
rect 16789 246131 16823 246273
rect 17209 246131 17243 246273
rect 17629 246131 17663 246273
rect 18049 246131 18083 246273
rect 18469 246131 18503 246273
rect 18889 246131 18923 246273
rect 19309 246131 19343 246273
rect 19729 246131 19763 246273
rect 20149 246131 20183 246273
rect 20569 246131 20603 246273
rect 20989 246131 21023 246273
rect 21409 246131 21443 246273
rect 21829 246131 21863 246273
rect 22249 246131 22283 246273
rect 22669 246131 22703 246273
rect 23089 246131 23123 246273
rect 23509 246131 23543 246273
rect 23929 246131 23963 246273
rect 24349 246131 24383 246273
rect 24769 246131 24803 246273
rect 25189 246131 25223 246273
rect 25609 246131 25643 246273
rect 26029 246131 26063 246273
rect 26449 246131 26483 246273
rect 26869 246131 26903 246273
rect 27289 246131 27323 246273
rect -4049 245296 -4015 246072
rect -3953 245296 -3919 246072
rect -3839 245296 -3805 246072
rect -3743 245296 -3709 246072
rect -3629 245296 -3595 246072
rect -3533 245296 -3499 246072
rect -3419 245296 -3385 246072
rect -3323 245296 -3289 246072
rect -3209 245296 -3175 246072
rect -3113 245296 -3079 246072
rect -2999 245296 -2965 246072
rect -2903 245296 -2869 246072
rect -2789 245296 -2755 246072
rect -2693 245296 -2659 246072
rect -2579 245296 -2545 246072
rect -2483 245296 -2449 246072
rect -2369 245296 -2335 246072
rect -2273 245296 -2239 246072
rect -2159 245296 -2125 246072
rect -2063 245296 -2029 246072
rect -1949 245296 -1915 246072
rect -1853 245296 -1819 246072
rect -1739 245296 -1705 246072
rect -1643 245296 -1609 246072
rect -1529 245296 -1495 246072
rect -1433 245296 -1399 246072
rect -1319 245296 -1285 246072
rect -1223 245296 -1189 246072
rect -1109 245296 -1075 246072
rect -1013 245296 -979 246072
rect -899 245296 -865 246072
rect -803 245296 -769 246072
rect -689 245296 -655 246072
rect -593 245296 -559 246072
rect -479 245296 -445 246072
rect -383 245296 -349 246072
rect -269 245296 -235 246072
rect -173 245296 -139 246072
rect -59 245296 -25 246072
rect 37 245296 71 246072
rect 151 245296 185 246072
rect 247 245296 281 246072
rect 361 245296 395 246072
rect 457 245296 491 246072
rect 571 245296 605 246072
rect 667 245296 701 246072
rect 781 245296 815 246072
rect 877 245296 911 246072
rect 991 245296 1025 246072
rect 1087 245296 1121 246072
rect 1201 245296 1235 246072
rect 1297 245296 1331 246072
rect 1411 245296 1445 246072
rect 1507 245296 1541 246072
rect 1621 245296 1655 246072
rect 1717 245296 1751 246072
rect 1831 245296 1865 246072
rect 1927 245296 1961 246072
rect 2041 245296 2075 246072
rect 2137 245296 2171 246072
rect 2251 245296 2285 246072
rect 2347 245296 2381 246072
rect 2461 245296 2495 246072
rect 2557 245296 2591 246072
rect 2671 245296 2705 246072
rect 2767 245296 2801 246072
rect 2881 245296 2915 246072
rect 2977 245296 3011 246072
rect 3091 245296 3125 246072
rect 3187 245296 3221 246072
rect 3301 245296 3335 246072
rect 3397 245296 3431 246072
rect 3511 245296 3545 246072
rect 3607 245296 3641 246072
rect 3721 245296 3755 246072
rect 3817 245296 3851 246072
rect 3931 245296 3965 246072
rect 4027 245296 4061 246072
rect 4141 245296 4175 246072
rect 4237 245296 4271 246072
rect 4351 245296 4385 246072
rect 4447 245296 4481 246072
rect 4561 245296 4595 246072
rect 4657 245296 4691 246072
rect 4771 245296 4805 246072
rect 4867 245296 4901 246072
rect 4981 245296 5015 246072
rect 5077 245296 5111 246072
rect 5191 245296 5225 246072
rect 5287 245296 5321 246072
rect 5401 245296 5435 246072
rect 5497 245296 5531 246072
rect 5611 245296 5645 246072
rect 5707 245296 5741 246072
rect 5821 245296 5855 246072
rect 5917 245296 5951 246072
rect 6031 245296 6065 246072
rect 6127 245296 6161 246072
rect 6241 245296 6275 246072
rect 6337 245296 6371 246072
rect 6451 245296 6485 246072
rect 6547 245296 6581 246072
rect 6661 245296 6695 246072
rect 6757 245296 6791 246072
rect 6871 245296 6905 246072
rect 6967 245296 7001 246072
rect 7081 245296 7115 246072
rect 7177 245296 7211 246072
rect 7291 245296 7325 246072
rect 7387 245296 7421 246072
rect 7501 245296 7535 246072
rect 7597 245296 7631 246072
rect 7711 245296 7745 246072
rect 7807 245296 7841 246072
rect 7921 245296 7955 246072
rect 8017 245296 8051 246072
rect 8131 245296 8165 246072
rect 8227 245296 8261 246072
rect 8341 245296 8375 246072
rect 8437 245296 8471 246072
rect 8551 245296 8585 246072
rect 8647 245296 8681 246072
rect 8761 245296 8795 246072
rect 8857 245296 8891 246072
rect 8971 245296 9005 246072
rect 9067 245296 9101 246072
rect 9181 245296 9215 246072
rect 9277 245296 9311 246072
rect 9391 245296 9425 246072
rect 9487 245296 9521 246072
rect 9601 245296 9635 246072
rect 9697 245296 9731 246072
rect 9811 245296 9845 246072
rect 9907 245296 9941 246072
rect 10021 245296 10055 246072
rect 10117 245296 10151 246072
rect 10231 245296 10265 246072
rect 10327 245296 10361 246072
rect 10441 245296 10475 246072
rect 10537 245296 10571 246072
rect 10651 245296 10685 246072
rect 10747 245296 10781 246072
rect 10861 245296 10895 246072
rect 10957 245296 10991 246072
rect 11071 245296 11105 246072
rect 11167 245296 11201 246072
rect 11281 245296 11315 246072
rect 11377 245296 11411 246072
rect 11491 245296 11525 246072
rect 11587 245296 11621 246072
rect 11701 245296 11735 246072
rect 11797 245296 11831 246072
rect 11911 245296 11945 246072
rect 12007 245296 12041 246072
rect 12121 245296 12155 246072
rect 12217 245296 12251 246072
rect 12331 245296 12365 246072
rect 12427 245296 12461 246072
rect 12541 245296 12575 246072
rect 12637 245296 12671 246072
rect 12751 245296 12785 246072
rect 12847 245296 12881 246072
rect 12961 245296 12995 246072
rect 13057 245296 13091 246072
rect 13171 245296 13205 246072
rect 13267 245296 13301 246072
rect 13381 245296 13415 246072
rect 13477 245296 13511 246072
rect 13591 245296 13625 246072
rect 13687 245296 13721 246072
rect 13801 245296 13835 246072
rect 13897 245296 13931 246072
rect 14011 245296 14045 246072
rect 14107 245296 14141 246072
rect 14221 245296 14255 246072
rect 14317 245296 14351 246072
rect 14431 245296 14465 246072
rect 14527 245296 14561 246072
rect 14641 245296 14675 246072
rect 14737 245296 14771 246072
rect 14851 245296 14885 246072
rect 14947 245296 14981 246072
rect 15061 245296 15095 246072
rect 15157 245296 15191 246072
rect 15271 245296 15305 246072
rect 15367 245296 15401 246072
rect 15481 245296 15515 246072
rect 15577 245296 15611 246072
rect 15691 245296 15725 246072
rect 15787 245296 15821 246072
rect 15901 245296 15935 246072
rect 15997 245296 16031 246072
rect 16111 245296 16145 246072
rect 16207 245296 16241 246072
rect 16321 245296 16355 246072
rect 16417 245296 16451 246072
rect 16531 245296 16565 246072
rect 16627 245296 16661 246072
rect 16741 245296 16775 246072
rect 16837 245296 16871 246072
rect 16951 245296 16985 246072
rect 17047 245296 17081 246072
rect 17161 245296 17195 246072
rect 17257 245296 17291 246072
rect 17371 245296 17405 246072
rect 17467 245296 17501 246072
rect 17581 245296 17615 246072
rect 17677 245296 17711 246072
rect 17791 245296 17825 246072
rect 17887 245296 17921 246072
rect 18001 245296 18035 246072
rect 18097 245296 18131 246072
rect 18211 245296 18245 246072
rect 18307 245296 18341 246072
rect 18421 245296 18455 246072
rect 18517 245296 18551 246072
rect 18631 245296 18665 246072
rect 18727 245296 18761 246072
rect 18841 245296 18875 246072
rect 18937 245296 18971 246072
rect 19051 245296 19085 246072
rect 19147 245296 19181 246072
rect 19261 245296 19295 246072
rect 19357 245296 19391 246072
rect 19471 245296 19505 246072
rect 19567 245296 19601 246072
rect 19681 245296 19715 246072
rect 19777 245296 19811 246072
rect 19891 245296 19925 246072
rect 19987 245296 20021 246072
rect 20101 245296 20135 246072
rect 20197 245296 20231 246072
rect 20311 245296 20345 246072
rect 20407 245296 20441 246072
rect 20521 245296 20555 246072
rect 20617 245296 20651 246072
rect 20731 245296 20765 246072
rect 20827 245296 20861 246072
rect 20941 245296 20975 246072
rect 21037 245296 21071 246072
rect 21151 245296 21185 246072
rect 21247 245296 21281 246072
rect 21361 245296 21395 246072
rect 21457 245296 21491 246072
rect 21571 245296 21605 246072
rect 21667 245296 21701 246072
rect 21781 245296 21815 246072
rect 21877 245296 21911 246072
rect 21991 245296 22025 246072
rect 22087 245296 22121 246072
rect 22201 245296 22235 246072
rect 22297 245296 22331 246072
rect 22411 245296 22445 246072
rect 22507 245296 22541 246072
rect 22621 245296 22655 246072
rect 22717 245296 22751 246072
rect 22831 245296 22865 246072
rect 22927 245296 22961 246072
rect 23041 245296 23075 246072
rect 23137 245296 23171 246072
rect 23251 245296 23285 246072
rect 23347 245296 23381 246072
rect 23461 245296 23495 246072
rect 23557 245296 23591 246072
rect 23671 245296 23705 246072
rect 23767 245296 23801 246072
rect 23881 245296 23915 246072
rect 23977 245296 24011 246072
rect 24091 245296 24125 246072
rect 24187 245296 24221 246072
rect 24301 245296 24335 246072
rect 24397 245296 24431 246072
rect 24511 245296 24545 246072
rect 24607 245296 24641 246072
rect 24721 245296 24755 246072
rect 24817 245296 24851 246072
rect 24931 245296 24965 246072
rect 25027 245296 25061 246072
rect 25141 245296 25175 246072
rect 25237 245296 25271 246072
rect 25351 245296 25385 246072
rect 25447 245296 25481 246072
rect 25561 245296 25595 246072
rect 25657 245296 25691 246072
rect 25771 245296 25805 246072
rect 25867 245296 25901 246072
rect 25981 245296 26015 246072
rect 26077 245296 26111 246072
rect 26191 245296 26225 246072
rect 26287 245296 26321 246072
rect 26401 245296 26435 246072
rect 26497 245296 26531 246072
rect 26611 245296 26645 246072
rect 26707 245296 26741 246072
rect 26821 245296 26855 246072
rect 26917 245296 26951 246072
rect 27031 245296 27065 246072
rect 27127 245296 27161 246072
rect 27241 245296 27275 246072
rect 27337 245296 27371 246072
rect -4001 245095 -3967 245237
rect -3581 245095 -3547 245237
rect -3161 245095 -3127 245237
rect -2741 245095 -2707 245237
rect -2321 245095 -2287 245237
rect -1901 245095 -1867 245237
rect -1481 245095 -1447 245237
rect -1061 245095 -1027 245237
rect -641 245095 -607 245237
rect -221 245095 -187 245237
rect 199 245095 233 245237
rect 619 245095 653 245237
rect 1039 245095 1073 245237
rect 1459 245095 1493 245237
rect 1879 245095 1913 245237
rect 2299 245095 2333 245237
rect 2719 245095 2753 245237
rect 3139 245095 3173 245237
rect 3559 245095 3593 245237
rect 3979 245095 4013 245237
rect 4399 245095 4433 245237
rect 4819 245095 4853 245237
rect 5239 245095 5273 245237
rect 5659 245095 5693 245237
rect 6079 245095 6113 245237
rect 6499 245095 6533 245237
rect 6919 245095 6953 245237
rect 7339 245095 7373 245237
rect 7759 245095 7793 245237
rect 8179 245095 8213 245237
rect 8599 245095 8633 245237
rect 9019 245095 9053 245237
rect 9439 245095 9473 245237
rect 9859 245095 9893 245237
rect 10279 245095 10313 245237
rect 10699 245095 10733 245237
rect 11119 245095 11153 245237
rect 11539 245095 11573 245237
rect 11959 245095 11993 245237
rect 12379 245095 12413 245237
rect 12799 245095 12833 245237
rect 13219 245095 13253 245237
rect 13639 245095 13673 245237
rect 14059 245095 14093 245237
rect 14479 245095 14513 245237
rect 14899 245095 14933 245237
rect 15319 245095 15353 245237
rect 15739 245095 15773 245237
rect 16159 245095 16193 245237
rect 16579 245095 16613 245237
rect 16999 245095 17033 245237
rect 17419 245095 17453 245237
rect 17839 245095 17873 245237
rect 18259 245095 18293 245237
rect 18679 245095 18713 245237
rect 19099 245095 19133 245237
rect 19519 245095 19553 245237
rect 19939 245095 19973 245237
rect 20359 245095 20393 245237
rect 20779 245095 20813 245237
rect 21199 245095 21233 245237
rect 21619 245095 21653 245237
rect 22039 245095 22073 245237
rect 22459 245095 22493 245237
rect 22879 245095 22913 245237
rect 23299 245095 23333 245237
rect 23719 245095 23753 245237
rect 24139 245095 24173 245237
rect 24559 245095 24593 245237
rect 24979 245095 25013 245237
rect 25399 245095 25433 245237
rect 25819 245095 25853 245237
rect 26239 245095 26273 245237
rect 26659 245095 26693 245237
rect 27079 245095 27113 245237
rect -4049 244260 -4015 245036
rect -3953 244260 -3919 245036
rect -3839 244260 -3805 245036
rect -3743 244260 -3709 245036
rect -3629 244260 -3595 245036
rect -3533 244260 -3499 245036
rect -3419 244260 -3385 245036
rect -3323 244260 -3289 245036
rect -3209 244260 -3175 245036
rect -3113 244260 -3079 245036
rect -2999 244260 -2965 245036
rect -2903 244260 -2869 245036
rect -2789 244260 -2755 245036
rect -2693 244260 -2659 245036
rect -2579 244260 -2545 245036
rect -2483 244260 -2449 245036
rect -2369 244260 -2335 245036
rect -2273 244260 -2239 245036
rect -2159 244260 -2125 245036
rect -2063 244260 -2029 245036
rect -1949 244260 -1915 245036
rect -1853 244260 -1819 245036
rect -1739 244260 -1705 245036
rect -1643 244260 -1609 245036
rect -1529 244260 -1495 245036
rect -1433 244260 -1399 245036
rect -1319 244260 -1285 245036
rect -1223 244260 -1189 245036
rect -1109 244260 -1075 245036
rect -1013 244260 -979 245036
rect -899 244260 -865 245036
rect -803 244260 -769 245036
rect -689 244260 -655 245036
rect -593 244260 -559 245036
rect -479 244260 -445 245036
rect -383 244260 -349 245036
rect -269 244260 -235 245036
rect -173 244260 -139 245036
rect -59 244260 -25 245036
rect 37 244260 71 245036
rect 151 244260 185 245036
rect 247 244260 281 245036
rect 361 244260 395 245036
rect 457 244260 491 245036
rect 571 244260 605 245036
rect 667 244260 701 245036
rect 781 244260 815 245036
rect 877 244260 911 245036
rect 991 244260 1025 245036
rect 1087 244260 1121 245036
rect 1201 244260 1235 245036
rect 1297 244260 1331 245036
rect 1411 244260 1445 245036
rect 1507 244260 1541 245036
rect 1621 244260 1655 245036
rect 1717 244260 1751 245036
rect 1831 244260 1865 245036
rect 1927 244260 1961 245036
rect 2041 244260 2075 245036
rect 2137 244260 2171 245036
rect 2251 244260 2285 245036
rect 2347 244260 2381 245036
rect 2461 244260 2495 245036
rect 2557 244260 2591 245036
rect 2671 244260 2705 245036
rect 2767 244260 2801 245036
rect 2881 244260 2915 245036
rect 2977 244260 3011 245036
rect 3091 244260 3125 245036
rect 3187 244260 3221 245036
rect 3301 244260 3335 245036
rect 3397 244260 3431 245036
rect 3511 244260 3545 245036
rect 3607 244260 3641 245036
rect 3721 244260 3755 245036
rect 3817 244260 3851 245036
rect 3931 244260 3965 245036
rect 4027 244260 4061 245036
rect 4141 244260 4175 245036
rect 4237 244260 4271 245036
rect 4351 244260 4385 245036
rect 4447 244260 4481 245036
rect 4561 244260 4595 245036
rect 4657 244260 4691 245036
rect 4771 244260 4805 245036
rect 4867 244260 4901 245036
rect 4981 244260 5015 245036
rect 5077 244260 5111 245036
rect 5191 244260 5225 245036
rect 5287 244260 5321 245036
rect 5401 244260 5435 245036
rect 5497 244260 5531 245036
rect 5611 244260 5645 245036
rect 5707 244260 5741 245036
rect 5821 244260 5855 245036
rect 5917 244260 5951 245036
rect 6031 244260 6065 245036
rect 6127 244260 6161 245036
rect 6241 244260 6275 245036
rect 6337 244260 6371 245036
rect 6451 244260 6485 245036
rect 6547 244260 6581 245036
rect 6661 244260 6695 245036
rect 6757 244260 6791 245036
rect 6871 244260 6905 245036
rect 6967 244260 7001 245036
rect 7081 244260 7115 245036
rect 7177 244260 7211 245036
rect 7291 244260 7325 245036
rect 7387 244260 7421 245036
rect 7501 244260 7535 245036
rect 7597 244260 7631 245036
rect 7711 244260 7745 245036
rect 7807 244260 7841 245036
rect 7921 244260 7955 245036
rect 8017 244260 8051 245036
rect 8131 244260 8165 245036
rect 8227 244260 8261 245036
rect 8341 244260 8375 245036
rect 8437 244260 8471 245036
rect 8551 244260 8585 245036
rect 8647 244260 8681 245036
rect 8761 244260 8795 245036
rect 8857 244260 8891 245036
rect 8971 244260 9005 245036
rect 9067 244260 9101 245036
rect 9181 244260 9215 245036
rect 9277 244260 9311 245036
rect 9391 244260 9425 245036
rect 9487 244260 9521 245036
rect 9601 244260 9635 245036
rect 9697 244260 9731 245036
rect 9811 244260 9845 245036
rect 9907 244260 9941 245036
rect 10021 244260 10055 245036
rect 10117 244260 10151 245036
rect 10231 244260 10265 245036
rect 10327 244260 10361 245036
rect 10441 244260 10475 245036
rect 10537 244260 10571 245036
rect 10651 244260 10685 245036
rect 10747 244260 10781 245036
rect 10861 244260 10895 245036
rect 10957 244260 10991 245036
rect 11071 244260 11105 245036
rect 11167 244260 11201 245036
rect 11281 244260 11315 245036
rect 11377 244260 11411 245036
rect 11491 244260 11525 245036
rect 11587 244260 11621 245036
rect 11701 244260 11735 245036
rect 11797 244260 11831 245036
rect 11911 244260 11945 245036
rect 12007 244260 12041 245036
rect 12121 244260 12155 245036
rect 12217 244260 12251 245036
rect 12331 244260 12365 245036
rect 12427 244260 12461 245036
rect 12541 244260 12575 245036
rect 12637 244260 12671 245036
rect 12751 244260 12785 245036
rect 12847 244260 12881 245036
rect 12961 244260 12995 245036
rect 13057 244260 13091 245036
rect 13171 244260 13205 245036
rect 13267 244260 13301 245036
rect 13381 244260 13415 245036
rect 13477 244260 13511 245036
rect 13591 244260 13625 245036
rect 13687 244260 13721 245036
rect 13801 244260 13835 245036
rect 13897 244260 13931 245036
rect 14011 244260 14045 245036
rect 14107 244260 14141 245036
rect 14221 244260 14255 245036
rect 14317 244260 14351 245036
rect 14431 244260 14465 245036
rect 14527 244260 14561 245036
rect 14641 244260 14675 245036
rect 14737 244260 14771 245036
rect 14851 244260 14885 245036
rect 14947 244260 14981 245036
rect 15061 244260 15095 245036
rect 15157 244260 15191 245036
rect 15271 244260 15305 245036
rect 15367 244260 15401 245036
rect 15481 244260 15515 245036
rect 15577 244260 15611 245036
rect 15691 244260 15725 245036
rect 15787 244260 15821 245036
rect 15901 244260 15935 245036
rect 15997 244260 16031 245036
rect 16111 244260 16145 245036
rect 16207 244260 16241 245036
rect 16321 244260 16355 245036
rect 16417 244260 16451 245036
rect 16531 244260 16565 245036
rect 16627 244260 16661 245036
rect 16741 244260 16775 245036
rect 16837 244260 16871 245036
rect 16951 244260 16985 245036
rect 17047 244260 17081 245036
rect 17161 244260 17195 245036
rect 17257 244260 17291 245036
rect 17371 244260 17405 245036
rect 17467 244260 17501 245036
rect 17581 244260 17615 245036
rect 17677 244260 17711 245036
rect 17791 244260 17825 245036
rect 17887 244260 17921 245036
rect 18001 244260 18035 245036
rect 18097 244260 18131 245036
rect 18211 244260 18245 245036
rect 18307 244260 18341 245036
rect 18421 244260 18455 245036
rect 18517 244260 18551 245036
rect 18631 244260 18665 245036
rect 18727 244260 18761 245036
rect 18841 244260 18875 245036
rect 18937 244260 18971 245036
rect 19051 244260 19085 245036
rect 19147 244260 19181 245036
rect 19261 244260 19295 245036
rect 19357 244260 19391 245036
rect 19471 244260 19505 245036
rect 19567 244260 19601 245036
rect 19681 244260 19715 245036
rect 19777 244260 19811 245036
rect 19891 244260 19925 245036
rect 19987 244260 20021 245036
rect 20101 244260 20135 245036
rect 20197 244260 20231 245036
rect 20311 244260 20345 245036
rect 20407 244260 20441 245036
rect 20521 244260 20555 245036
rect 20617 244260 20651 245036
rect 20731 244260 20765 245036
rect 20827 244260 20861 245036
rect 20941 244260 20975 245036
rect 21037 244260 21071 245036
rect 21151 244260 21185 245036
rect 21247 244260 21281 245036
rect 21361 244260 21395 245036
rect 21457 244260 21491 245036
rect 21571 244260 21605 245036
rect 21667 244260 21701 245036
rect 21781 244260 21815 245036
rect 21877 244260 21911 245036
rect 21991 244260 22025 245036
rect 22087 244260 22121 245036
rect 22201 244260 22235 245036
rect 22297 244260 22331 245036
rect 22411 244260 22445 245036
rect 22507 244260 22541 245036
rect 22621 244260 22655 245036
rect 22717 244260 22751 245036
rect 22831 244260 22865 245036
rect 22927 244260 22961 245036
rect 23041 244260 23075 245036
rect 23137 244260 23171 245036
rect 23251 244260 23285 245036
rect 23347 244260 23381 245036
rect 23461 244260 23495 245036
rect 23557 244260 23591 245036
rect 23671 244260 23705 245036
rect 23767 244260 23801 245036
rect 23881 244260 23915 245036
rect 23977 244260 24011 245036
rect 24091 244260 24125 245036
rect 24187 244260 24221 245036
rect 24301 244260 24335 245036
rect 24397 244260 24431 245036
rect 24511 244260 24545 245036
rect 24607 244260 24641 245036
rect 24721 244260 24755 245036
rect 24817 244260 24851 245036
rect 24931 244260 24965 245036
rect 25027 244260 25061 245036
rect 25141 244260 25175 245036
rect 25237 244260 25271 245036
rect 25351 244260 25385 245036
rect 25447 244260 25481 245036
rect 25561 244260 25595 245036
rect 25657 244260 25691 245036
rect 25771 244260 25805 245036
rect 25867 244260 25901 245036
rect 25981 244260 26015 245036
rect 26077 244260 26111 245036
rect 26191 244260 26225 245036
rect 26287 244260 26321 245036
rect 26401 244260 26435 245036
rect 26497 244260 26531 245036
rect 26611 244260 26645 245036
rect 26707 244260 26741 245036
rect 26821 244260 26855 245036
rect 26917 244260 26951 245036
rect 27031 244260 27065 245036
rect 27127 244260 27161 245036
rect 27241 244260 27275 245036
rect 27337 244260 27371 245036
rect -3791 244167 -3695 244201
rect -3371 244167 -3275 244201
rect -2951 244167 -2855 244201
rect -2531 244167 -2435 244201
rect -2111 244167 -2015 244201
rect -1691 244167 -1595 244201
rect -1271 244167 -1175 244201
rect -851 244167 -755 244201
rect -431 244167 -335 244201
rect -11 244167 85 244201
rect 409 244167 505 244201
rect 829 244167 925 244201
rect 1249 244167 1345 244201
rect 1669 244167 1765 244201
rect 2089 244167 2185 244201
rect 2509 244167 2605 244201
rect 2929 244167 3025 244201
rect 3349 244167 3445 244201
rect 3769 244167 3865 244201
rect 4189 244167 4285 244201
rect 4609 244167 4705 244201
rect 5029 244167 5125 244201
rect 5449 244167 5545 244201
rect 5869 244167 5965 244201
rect 6289 244167 6385 244201
rect 6709 244167 6805 244201
rect 7129 244167 7225 244201
rect 7549 244167 7645 244201
rect 7969 244167 8065 244201
rect 8389 244167 8485 244201
rect 8809 244167 8905 244201
rect 9229 244167 9325 244201
rect 9649 244167 9745 244201
rect 10069 244167 10165 244201
rect 10489 244167 10585 244201
rect 10909 244167 11005 244201
rect 11329 244167 11425 244201
rect 11749 244167 11845 244201
rect 12169 244167 12265 244201
rect 12589 244167 12685 244201
rect 13009 244167 13105 244201
rect 13429 244167 13525 244201
rect 13849 244167 13945 244201
rect 14269 244167 14365 244201
rect 14689 244167 14785 244201
rect 15109 244167 15205 244201
rect 15529 244167 15625 244201
rect 15949 244167 16045 244201
rect 16369 244167 16465 244201
rect 16789 244167 16885 244201
rect 17209 244167 17305 244201
rect 17629 244167 17725 244201
rect 18049 244167 18145 244201
rect 18469 244167 18565 244201
rect 18889 244167 18985 244201
rect 19309 244167 19405 244201
rect 19729 244167 19825 244201
rect 20149 244167 20245 244201
rect 20569 244167 20665 244201
rect 20989 244167 21085 244201
rect 21409 244167 21505 244201
rect 21829 244167 21925 244201
rect 22249 244167 22345 244201
rect 22669 244167 22765 244201
rect 23089 244167 23185 244201
rect 23509 244167 23605 244201
rect 23929 244167 24025 244201
rect 24349 244167 24445 244201
rect 24769 244167 24865 244201
rect 25189 244167 25285 244201
rect 25609 244167 25705 244201
rect 26029 244167 26125 244201
rect 26449 244167 26545 244201
rect 26869 244167 26965 244201
rect 27289 244167 27385 244201
rect -4163 243960 27485 244065
<< metal1 >>
rect 27300 264323 27310 264430
rect -4175 264317 27310 264323
rect -4175 264212 -4163 264317
rect 27510 264230 27520 264430
rect 27486 264212 27498 264230
rect -4175 264206 27498 264212
rect -5008 264110 27192 264116
rect -5008 264076 -4001 264110
rect -3905 264076 -3581 264110
rect -3485 264076 -3161 264110
rect -3065 264076 -2741 264110
rect -2645 264076 -2321 264110
rect -2225 264076 -1901 264110
rect -1805 264076 -1481 264110
rect -1385 264076 -1061 264110
rect -965 264076 -641 264110
rect -545 264076 -221 264110
rect -125 264076 199 264110
rect 295 264076 619 264110
rect 715 264076 1039 264110
rect 1135 264076 1459 264110
rect 1555 264076 1879 264110
rect 1975 264076 2299 264110
rect 2395 264076 2719 264110
rect 2815 264076 3139 264110
rect 3235 264076 3559 264110
rect 3655 264076 3979 264110
rect 4075 264076 4399 264110
rect 4495 264076 4819 264110
rect 4915 264076 5239 264110
rect 5335 264076 5659 264110
rect 5755 264076 6079 264110
rect 6175 264076 6499 264110
rect 6595 264076 6919 264110
rect 7015 264076 7339 264110
rect 7435 264076 7759 264110
rect 7855 264076 8179 264110
rect 8275 264076 8599 264110
rect 8695 264076 9019 264110
rect 9115 264076 9439 264110
rect 9535 264076 9859 264110
rect 9955 264076 10279 264110
rect 10375 264076 10699 264110
rect 10795 264076 11119 264110
rect 11215 264076 11539 264110
rect 11635 264076 11959 264110
rect 12055 264076 12379 264110
rect 12475 264076 12799 264110
rect 12895 264076 13219 264110
rect 13315 264076 13639 264110
rect 13735 264076 14059 264110
rect 14155 264076 14479 264110
rect 14575 264076 14899 264110
rect 14995 264076 15319 264110
rect 15415 264076 15739 264110
rect 15835 264076 16159 264110
rect 16255 264076 16579 264110
rect 16675 264076 16999 264110
rect 17095 264076 17419 264110
rect 17515 264076 17839 264110
rect 17935 264076 18259 264110
rect 18355 264076 18679 264110
rect 18775 264076 19099 264110
rect 19195 264076 19519 264110
rect 19615 264076 19939 264110
rect 20035 264076 20359 264110
rect 20455 264076 20779 264110
rect 20875 264076 21199 264110
rect 21295 264076 21619 264110
rect 21715 264076 22039 264110
rect 22135 264076 22459 264110
rect 22555 264076 22879 264110
rect 22975 264076 23299 264110
rect 23395 264076 23719 264110
rect 23815 264076 24139 264110
rect 24235 264076 24559 264110
rect 24655 264076 24979 264110
rect 25075 264076 25399 264110
rect 25495 264076 25819 264110
rect 25915 264076 26239 264110
rect 26335 264076 26659 264110
rect 26755 264076 27079 264110
rect 27175 264076 27192 264110
rect -5008 264070 27192 264076
rect -5008 263198 -4244 264070
rect 27375 264038 27423 264206
rect -4040 264036 -4009 264038
rect -4070 264026 -4009 264036
rect -3959 264026 -3913 264038
rect -3845 264026 -3799 264038
rect -3749 264026 -3703 264038
rect -3635 264026 -3589 264038
rect -3539 264026 -3493 264038
rect -3425 264026 -3379 264038
rect -3329 264026 -3283 264038
rect -3215 264026 -3169 264038
rect -3119 264026 -3073 264038
rect -3005 264026 -2959 264038
rect -2909 264026 -2863 264038
rect -2795 264026 -2749 264038
rect -2699 264026 -2653 264038
rect -2585 264026 -2539 264038
rect -2489 264026 -2443 264038
rect -2375 264026 -2329 264038
rect -2279 264026 -2233 264038
rect -2165 264026 -2119 264038
rect -2069 264026 -2023 264038
rect -1955 264026 -1909 264038
rect -1859 264026 -1813 264038
rect -1745 264026 -1699 264038
rect -1649 264026 -1603 264038
rect -1535 264026 -1489 264038
rect -1439 264026 -1393 264038
rect -1325 264026 -1279 264038
rect -1229 264026 -1183 264038
rect -1115 264026 -1069 264038
rect -1019 264026 -973 264038
rect -905 264026 -859 264038
rect -809 264026 -763 264038
rect -695 264026 -649 264038
rect -599 264026 -553 264038
rect -485 264026 -439 264038
rect -389 264026 -343 264038
rect -275 264026 -229 264038
rect -179 264026 -133 264038
rect -65 264026 -19 264038
rect 31 264026 77 264038
rect 145 264026 191 264038
rect 241 264026 287 264038
rect 355 264026 401 264038
rect 451 264026 497 264038
rect 565 264026 611 264038
rect 661 264026 707 264038
rect 775 264026 821 264038
rect 871 264026 917 264038
rect 985 264026 1031 264038
rect 1081 264026 1127 264038
rect 1195 264026 1241 264038
rect 1291 264026 1337 264038
rect 1405 264026 1451 264038
rect 1501 264026 1547 264038
rect 1615 264026 1661 264038
rect 1711 264026 1757 264038
rect 1825 264026 1871 264038
rect 1921 264026 1967 264038
rect 2035 264026 2081 264038
rect 2131 264026 2177 264038
rect 2245 264026 2291 264038
rect 2341 264026 2387 264038
rect 2455 264026 2501 264038
rect 2551 264026 2597 264038
rect 2665 264026 2711 264038
rect 2761 264026 2807 264038
rect 2875 264026 2921 264038
rect 2971 264026 3017 264038
rect 3085 264026 3131 264038
rect 3181 264026 3227 264038
rect 3295 264026 3341 264038
rect 3391 264026 3437 264038
rect 3505 264026 3551 264038
rect 3601 264026 3647 264038
rect 3715 264026 3761 264038
rect 3811 264026 3857 264038
rect 3925 264026 3971 264038
rect 4021 264026 4067 264038
rect 4135 264026 4181 264038
rect 4231 264026 4277 264038
rect 4345 264026 4391 264038
rect 4441 264026 4487 264038
rect 4555 264026 4601 264038
rect 4651 264026 4697 264038
rect 4765 264026 4811 264038
rect 4861 264026 4907 264038
rect 4975 264026 5021 264038
rect 5071 264026 5117 264038
rect 5185 264026 5231 264038
rect 5281 264026 5327 264038
rect 5395 264026 5441 264038
rect 5491 264026 5537 264038
rect 5605 264026 5651 264038
rect 5701 264026 5747 264038
rect 5815 264026 5861 264038
rect 5911 264026 5957 264038
rect 6025 264026 6071 264038
rect 6121 264026 6167 264038
rect 6235 264026 6281 264038
rect 6331 264026 6377 264038
rect 6445 264026 6491 264038
rect 6541 264026 6587 264038
rect 6655 264026 6701 264038
rect 6751 264026 6797 264038
rect 6865 264026 6911 264038
rect 6961 264026 7007 264038
rect 7075 264026 7121 264038
rect 7171 264026 7217 264038
rect 7285 264026 7331 264038
rect 7381 264026 7427 264038
rect 7495 264026 7541 264038
rect 7591 264026 7637 264038
rect 7705 264026 7751 264038
rect 7801 264026 7847 264038
rect 7915 264026 7961 264038
rect 8011 264026 8057 264038
rect 8125 264026 8171 264038
rect 8221 264026 8267 264038
rect 8335 264026 8381 264038
rect 8431 264026 8477 264038
rect 8545 264026 8591 264038
rect 8641 264026 8687 264038
rect 8755 264026 8801 264038
rect 8851 264026 8897 264038
rect 8965 264026 9011 264038
rect 9061 264026 9107 264038
rect 9175 264026 9221 264038
rect 9271 264026 9317 264038
rect 9385 264026 9431 264038
rect 9481 264026 9527 264038
rect 9595 264026 9641 264038
rect 9691 264026 9737 264038
rect 9805 264026 9851 264038
rect 9901 264026 9947 264038
rect 10015 264026 10061 264038
rect 10111 264026 10157 264038
rect 10225 264026 10271 264038
rect 10321 264026 10367 264038
rect 10435 264026 10481 264038
rect 10531 264026 10577 264038
rect 10645 264026 10691 264038
rect 10741 264026 10787 264038
rect 10855 264026 10901 264038
rect 10951 264026 10997 264038
rect 11065 264026 11111 264038
rect 11161 264026 11207 264038
rect 11275 264026 11321 264038
rect 11371 264026 11417 264038
rect 11485 264026 11531 264038
rect 11581 264026 11627 264038
rect 11695 264026 11741 264038
rect 11791 264026 11837 264038
rect 11905 264026 11951 264038
rect 12001 264026 12047 264038
rect 12115 264026 12161 264038
rect 12211 264026 12257 264038
rect 12325 264026 12371 264038
rect 12421 264026 12467 264038
rect 12535 264026 12581 264038
rect 12631 264026 12677 264038
rect 12745 264026 12791 264038
rect 12841 264026 12887 264038
rect 12955 264026 13001 264038
rect 13051 264026 13097 264038
rect 13165 264026 13211 264038
rect 13261 264026 13307 264038
rect 13375 264026 13421 264038
rect 13471 264026 13517 264038
rect 13585 264026 13631 264038
rect 13681 264026 13727 264038
rect 13795 264026 13841 264038
rect 13891 264026 13937 264038
rect 14005 264026 14051 264038
rect 14101 264026 14147 264038
rect 14215 264026 14261 264038
rect 14311 264026 14357 264038
rect 14425 264026 14471 264038
rect 14521 264026 14567 264038
rect 14635 264026 14681 264038
rect 14731 264026 14777 264038
rect 14845 264026 14891 264038
rect 14941 264026 14987 264038
rect 15055 264026 15101 264038
rect 15151 264026 15197 264038
rect 15265 264026 15311 264038
rect 15361 264026 15407 264038
rect 15475 264026 15521 264038
rect 15571 264026 15617 264038
rect 15685 264026 15731 264038
rect 15781 264026 15827 264038
rect 15895 264026 15941 264038
rect 15991 264026 16037 264038
rect 16105 264026 16151 264038
rect 16201 264026 16247 264038
rect 16315 264026 16361 264038
rect 16411 264026 16457 264038
rect 16525 264026 16571 264038
rect 16621 264026 16667 264038
rect 16735 264026 16781 264038
rect 16831 264026 16877 264038
rect 16945 264026 16991 264038
rect 17041 264026 17087 264038
rect 17155 264026 17201 264038
rect 17251 264026 17297 264038
rect 17365 264026 17411 264038
rect 17461 264026 17507 264038
rect 17575 264026 17621 264038
rect 17671 264026 17717 264038
rect 17785 264026 17831 264038
rect 17881 264026 17927 264038
rect 17995 264026 18041 264038
rect 18091 264026 18137 264038
rect 18205 264026 18251 264038
rect 18301 264026 18347 264038
rect 18415 264026 18461 264038
rect 18511 264026 18557 264038
rect 18625 264026 18671 264038
rect 18721 264026 18767 264038
rect 18835 264026 18881 264038
rect 18931 264026 18977 264038
rect 19045 264026 19091 264038
rect 19141 264026 19187 264038
rect 19255 264026 19301 264038
rect 19351 264026 19397 264038
rect 19465 264026 19511 264038
rect 19561 264026 19607 264038
rect 19675 264026 19721 264038
rect 19771 264026 19817 264038
rect 19885 264026 19931 264038
rect 19981 264026 20027 264038
rect 20095 264026 20141 264038
rect 20191 264026 20237 264038
rect 20305 264026 20351 264038
rect 20401 264026 20447 264038
rect 20515 264026 20561 264038
rect 20611 264026 20657 264038
rect 20725 264026 20771 264038
rect 20821 264026 20867 264038
rect 20935 264026 20981 264038
rect 21031 264026 21077 264038
rect 21145 264026 21191 264038
rect 21241 264026 21287 264038
rect 21355 264026 21401 264038
rect 21451 264026 21497 264038
rect 21565 264026 21611 264038
rect 21661 264026 21707 264038
rect 21775 264026 21821 264038
rect 21871 264026 21917 264038
rect 21985 264026 22031 264038
rect 22081 264026 22127 264038
rect 22195 264026 22241 264038
rect 22291 264026 22337 264038
rect 22405 264026 22451 264038
rect 22501 264026 22547 264038
rect 22615 264026 22661 264038
rect 22711 264026 22757 264038
rect 22825 264026 22871 264038
rect 22921 264026 22967 264038
rect 23035 264026 23081 264038
rect 23131 264026 23177 264038
rect 23245 264026 23291 264038
rect 23341 264026 23387 264038
rect 23455 264026 23501 264038
rect 23551 264026 23597 264038
rect 23665 264026 23711 264038
rect 23761 264026 23807 264038
rect 23875 264026 23921 264038
rect 23971 264026 24017 264038
rect 24085 264026 24131 264038
rect 24181 264026 24227 264038
rect 24295 264026 24341 264038
rect 24391 264026 24437 264038
rect 24505 264026 24551 264038
rect 24601 264026 24647 264038
rect 24715 264026 24761 264038
rect 24811 264026 24857 264038
rect 24925 264026 24971 264038
rect 25021 264026 25067 264038
rect 25135 264026 25181 264038
rect 25231 264026 25277 264038
rect 25345 264026 25391 264038
rect 25441 264026 25487 264038
rect 25555 264026 25601 264038
rect 25651 264026 25697 264038
rect 25765 264026 25811 264038
rect 25861 264026 25907 264038
rect 25975 264026 26021 264038
rect 26071 264026 26117 264038
rect 26185 264026 26231 264038
rect 26281 264026 26327 264038
rect 26395 264026 26441 264038
rect 26491 264026 26537 264038
rect 26605 264026 26651 264038
rect 26701 264026 26747 264038
rect 26815 264026 26861 264038
rect 26911 264026 26957 264038
rect 27025 264026 27071 264038
rect 27121 264026 27167 264038
rect 27235 264026 27281 264038
rect 27331 264026 27423 264038
rect -4015 263250 -4005 264026
rect -3963 263250 -3953 264026
rect -3805 263250 -3795 264026
rect -3753 263250 -3743 264026
rect -3595 263250 -3585 264026
rect -3543 263250 -3533 264026
rect -3385 263250 -3375 264026
rect -3333 263250 -3323 264026
rect -3175 263250 -3165 264026
rect -3123 263250 -3113 264026
rect -2965 263250 -2955 264026
rect -2913 263250 -2903 264026
rect -2755 263250 -2745 264026
rect -2703 263250 -2693 264026
rect -2545 263250 -2535 264026
rect -2493 263250 -2483 264026
rect -2335 263250 -2325 264026
rect -2283 263250 -2273 264026
rect -2125 263250 -2115 264026
rect -2073 263250 -2063 264026
rect -1915 263250 -1905 264026
rect -1863 263250 -1853 264026
rect -1705 263250 -1695 264026
rect -1653 263250 -1643 264026
rect -1495 263250 -1485 264026
rect -1443 263250 -1433 264026
rect -1285 263250 -1275 264026
rect -1233 263250 -1223 264026
rect -1075 263250 -1065 264026
rect -1023 263250 -1013 264026
rect -865 263250 -855 264026
rect -813 263250 -803 264026
rect -655 263250 -645 264026
rect -603 263250 -593 264026
rect -445 263250 -435 264026
rect -393 263250 -383 264026
rect -235 263250 -225 264026
rect -183 263250 -173 264026
rect -25 263250 -15 264026
rect 27 263250 37 264026
rect 185 263250 195 264026
rect 237 263250 247 264026
rect 395 263250 405 264026
rect 447 263250 457 264026
rect 605 263250 615 264026
rect 657 263250 667 264026
rect 815 263250 825 264026
rect 867 263250 877 264026
rect 1025 263250 1035 264026
rect 1077 263250 1087 264026
rect 1235 263250 1245 264026
rect 1287 263250 1297 264026
rect 1445 263250 1455 264026
rect 1497 263250 1507 264026
rect 1655 263250 1665 264026
rect 1707 263250 1717 264026
rect 1865 263250 1875 264026
rect 1917 263250 1927 264026
rect 2075 263250 2085 264026
rect 2127 263250 2137 264026
rect 2285 263250 2295 264026
rect 2337 263250 2347 264026
rect 2495 263250 2505 264026
rect 2547 263250 2557 264026
rect 2705 263250 2715 264026
rect 2757 263250 2767 264026
rect 2915 263250 2925 264026
rect 2967 263250 2977 264026
rect 3125 263250 3135 264026
rect 3177 263250 3187 264026
rect 3335 263250 3345 264026
rect 3387 263250 3397 264026
rect 3545 263250 3555 264026
rect 3597 263250 3607 264026
rect 3755 263250 3765 264026
rect 3807 263250 3817 264026
rect 3965 263250 3975 264026
rect 4017 263250 4027 264026
rect 4175 263250 4185 264026
rect 4227 263250 4237 264026
rect 4385 263250 4395 264026
rect 4437 263250 4447 264026
rect 4595 263250 4605 264026
rect 4647 263250 4657 264026
rect 4805 263250 4815 264026
rect 4857 263250 4867 264026
rect 5015 263250 5025 264026
rect 5067 263250 5077 264026
rect 5225 263250 5235 264026
rect 5277 263250 5287 264026
rect 5435 263250 5445 264026
rect 5487 263250 5497 264026
rect 5645 263250 5655 264026
rect 5697 263250 5707 264026
rect 5855 263250 5865 264026
rect 5907 263250 5917 264026
rect 6065 263250 6075 264026
rect 6117 263250 6127 264026
rect 6275 263250 6285 264026
rect 6327 263250 6337 264026
rect 6485 263250 6495 264026
rect 6537 263250 6547 264026
rect 6695 263250 6705 264026
rect 6747 263250 6757 264026
rect 6905 263250 6915 264026
rect 6957 263250 6967 264026
rect 7115 263250 7125 264026
rect 7167 263250 7177 264026
rect 7325 263250 7335 264026
rect 7377 263250 7387 264026
rect 7535 263250 7545 264026
rect 7587 263250 7597 264026
rect 7745 263250 7755 264026
rect 7797 263250 7807 264026
rect 7955 263250 7965 264026
rect 8007 263250 8017 264026
rect 8165 263250 8175 264026
rect 8217 263250 8227 264026
rect 8375 263250 8385 264026
rect 8427 263250 8437 264026
rect 8585 263250 8595 264026
rect 8637 263250 8647 264026
rect 8795 263250 8805 264026
rect 8847 263250 8857 264026
rect 9005 263250 9015 264026
rect 9057 263250 9067 264026
rect 9215 263250 9225 264026
rect 9267 263250 9277 264026
rect 9425 263250 9435 264026
rect 9477 263250 9487 264026
rect 9635 263250 9645 264026
rect 9687 263250 9697 264026
rect 9845 263250 9855 264026
rect 9897 263250 9907 264026
rect 10055 263250 10065 264026
rect 10107 263250 10117 264026
rect 10265 263250 10275 264026
rect 10317 263250 10327 264026
rect 10475 263250 10485 264026
rect 10527 263250 10537 264026
rect 10685 263250 10695 264026
rect 10737 263250 10747 264026
rect 10895 263250 10905 264026
rect 10947 263250 10957 264026
rect 11105 263250 11115 264026
rect 11157 263250 11167 264026
rect 11315 263250 11325 264026
rect 11367 263250 11377 264026
rect 11525 263250 11535 264026
rect 11577 263250 11587 264026
rect 11735 263250 11745 264026
rect 11787 263250 11797 264026
rect 11945 263250 11955 264026
rect 11997 263250 12007 264026
rect 12155 263250 12165 264026
rect 12207 263250 12217 264026
rect 12365 263250 12375 264026
rect 12417 263250 12427 264026
rect 12575 263250 12585 264026
rect 12627 263250 12637 264026
rect 12785 263250 12795 264026
rect 12837 263250 12847 264026
rect 12995 263250 13005 264026
rect 13047 263250 13057 264026
rect 13205 263250 13215 264026
rect 13257 263250 13267 264026
rect 13415 263250 13425 264026
rect 13467 263250 13477 264026
rect 13625 263250 13635 264026
rect 13677 263250 13687 264026
rect 13835 263250 13845 264026
rect 13887 263250 13897 264026
rect 14045 263250 14055 264026
rect 14097 263250 14107 264026
rect 14255 263250 14265 264026
rect 14307 263250 14317 264026
rect 14465 263250 14475 264026
rect 14517 263250 14527 264026
rect 14675 263250 14685 264026
rect 14727 263250 14737 264026
rect 14885 263250 14895 264026
rect 14937 263250 14947 264026
rect 15095 263250 15105 264026
rect 15147 263250 15157 264026
rect 15305 263250 15315 264026
rect 15357 263250 15367 264026
rect 15515 263250 15525 264026
rect 15567 263250 15577 264026
rect 15725 263250 15735 264026
rect 15777 263250 15787 264026
rect 15935 263250 15945 264026
rect 15987 263250 15997 264026
rect 16145 263250 16155 264026
rect 16197 263250 16207 264026
rect 16355 263250 16365 264026
rect 16407 263250 16417 264026
rect 16565 263250 16575 264026
rect 16617 263250 16627 264026
rect 16775 263250 16785 264026
rect 16827 263250 16837 264026
rect 16985 263250 16995 264026
rect 17037 263250 17047 264026
rect 17195 263250 17205 264026
rect 17247 263250 17257 264026
rect 17405 263250 17415 264026
rect 17457 263250 17467 264026
rect 17615 263250 17625 264026
rect 17667 263250 17677 264026
rect 17825 263250 17835 264026
rect 17877 263250 17887 264026
rect 18035 263250 18045 264026
rect 18087 263250 18097 264026
rect 18245 263250 18255 264026
rect 18297 263250 18307 264026
rect 18455 263250 18465 264026
rect 18507 263250 18517 264026
rect 18665 263250 18675 264026
rect 18717 263250 18727 264026
rect 18875 263250 18885 264026
rect 18927 263250 18937 264026
rect 19085 263250 19095 264026
rect 19137 263250 19147 264026
rect 19295 263250 19305 264026
rect 19347 263250 19357 264026
rect 19505 263250 19515 264026
rect 19557 263250 19567 264026
rect 19715 263250 19725 264026
rect 19767 263250 19777 264026
rect 19925 263250 19935 264026
rect 19977 263250 19987 264026
rect 20135 263250 20145 264026
rect 20187 263250 20197 264026
rect 20345 263250 20355 264026
rect 20397 263250 20407 264026
rect 20555 263250 20565 264026
rect 20607 263250 20617 264026
rect 20765 263250 20775 264026
rect 20817 263250 20827 264026
rect 20975 263250 20985 264026
rect 21027 263250 21037 264026
rect 21185 263250 21195 264026
rect 21237 263250 21247 264026
rect 21395 263250 21405 264026
rect 21447 263250 21457 264026
rect 21605 263250 21615 264026
rect 21657 263250 21667 264026
rect 21815 263250 21825 264026
rect 21867 263250 21877 264026
rect 22025 263250 22035 264026
rect 22077 263250 22087 264026
rect 22235 263250 22245 264026
rect 22287 263250 22297 264026
rect 22445 263250 22455 264026
rect 22497 263250 22507 264026
rect 22655 263250 22665 264026
rect 22707 263250 22717 264026
rect 22865 263250 22875 264026
rect 22917 263250 22927 264026
rect 23075 263250 23085 264026
rect 23127 263250 23137 264026
rect 23285 263250 23295 264026
rect 23337 263250 23347 264026
rect 23495 263250 23505 264026
rect 23547 263250 23557 264026
rect 23705 263250 23715 264026
rect 23757 263250 23767 264026
rect 23915 263250 23925 264026
rect 23967 263250 23977 264026
rect 24125 263250 24135 264026
rect 24177 263250 24187 264026
rect 24335 263250 24345 264026
rect 24387 263250 24397 264026
rect 24545 263250 24555 264026
rect 24597 263250 24607 264026
rect 24755 263250 24765 264026
rect 24807 263250 24817 264026
rect 24965 263250 24975 264026
rect 25017 263250 25027 264026
rect 25175 263250 25185 264026
rect 25227 263250 25237 264026
rect 25385 263250 25395 264026
rect 25437 263250 25447 264026
rect 25595 263250 25605 264026
rect 25647 263250 25657 264026
rect 25805 263250 25815 264026
rect 25857 263250 25867 264026
rect 26015 263250 26025 264026
rect 26067 263250 26077 264026
rect 26225 263250 26235 264026
rect 26277 263250 26287 264026
rect 26435 263250 26445 264026
rect 26487 263250 26497 264026
rect 26645 263250 26655 264026
rect 26697 263250 26707 264026
rect 26855 263250 26865 264026
rect 26907 263250 26917 264026
rect 27065 263250 27075 264026
rect 27117 263250 27127 264026
rect 27275 263250 27285 264026
rect 27331 263250 27337 264026
rect 27371 263250 27423 264026
rect -4070 263238 -4009 263250
rect -3959 263238 -3913 263250
rect -3845 263238 -3799 263250
rect -3749 263238 -3703 263250
rect -3635 263238 -3589 263250
rect -3539 263238 -3493 263250
rect -3425 263238 -3379 263250
rect -3329 263238 -3283 263250
rect -3215 263238 -3169 263250
rect -3119 263238 -3073 263250
rect -3005 263238 -2959 263250
rect -2909 263238 -2863 263250
rect -2795 263238 -2749 263250
rect -2699 263238 -2653 263250
rect -2585 263238 -2539 263250
rect -2489 263238 -2443 263250
rect -2375 263238 -2329 263250
rect -2279 263238 -2233 263250
rect -2165 263238 -2119 263250
rect -2069 263238 -2023 263250
rect -1955 263238 -1909 263250
rect -1859 263238 -1813 263250
rect -1745 263238 -1699 263250
rect -1649 263238 -1603 263250
rect -1535 263238 -1489 263250
rect -1439 263238 -1393 263250
rect -1325 263238 -1279 263250
rect -1229 263238 -1183 263250
rect -1115 263238 -1069 263250
rect -1019 263238 -973 263250
rect -905 263238 -859 263250
rect -809 263238 -763 263250
rect -695 263238 -649 263250
rect -599 263238 -553 263250
rect -485 263238 -439 263250
rect -389 263238 -343 263250
rect -275 263238 -229 263250
rect -179 263238 -133 263250
rect -65 263238 -19 263250
rect 31 263238 77 263250
rect 145 263238 191 263250
rect 241 263238 287 263250
rect 355 263238 401 263250
rect 451 263238 497 263250
rect 565 263238 611 263250
rect 661 263238 707 263250
rect 775 263238 821 263250
rect 871 263238 917 263250
rect 985 263238 1031 263250
rect 1081 263238 1127 263250
rect 1195 263238 1241 263250
rect 1291 263238 1337 263250
rect 1405 263238 1451 263250
rect 1501 263238 1547 263250
rect 1615 263238 1661 263250
rect 1711 263238 1757 263250
rect 1825 263238 1871 263250
rect 1921 263238 1967 263250
rect 2035 263238 2081 263250
rect 2131 263238 2177 263250
rect 2245 263238 2291 263250
rect 2341 263238 2387 263250
rect 2455 263238 2501 263250
rect 2551 263238 2597 263250
rect 2665 263238 2711 263250
rect 2761 263238 2807 263250
rect 2875 263238 2921 263250
rect 2971 263238 3017 263250
rect 3085 263238 3131 263250
rect 3181 263238 3227 263250
rect 3295 263238 3341 263250
rect 3391 263238 3437 263250
rect 3505 263238 3551 263250
rect 3601 263238 3647 263250
rect 3715 263238 3761 263250
rect 3811 263238 3857 263250
rect 3925 263238 3971 263250
rect 4021 263238 4067 263250
rect 4135 263238 4181 263250
rect 4231 263238 4277 263250
rect 4345 263238 4391 263250
rect 4441 263238 4487 263250
rect 4555 263238 4601 263250
rect 4651 263238 4697 263250
rect 4765 263238 4811 263250
rect 4861 263238 4907 263250
rect 4975 263238 5021 263250
rect 5071 263238 5117 263250
rect 5185 263238 5231 263250
rect 5281 263238 5327 263250
rect 5395 263238 5441 263250
rect 5491 263238 5537 263250
rect 5605 263238 5651 263250
rect 5701 263238 5747 263250
rect 5815 263238 5861 263250
rect 5911 263238 5957 263250
rect 6025 263238 6071 263250
rect 6121 263238 6167 263250
rect 6235 263238 6281 263250
rect 6331 263238 6377 263250
rect 6445 263238 6491 263250
rect 6541 263238 6587 263250
rect 6655 263238 6701 263250
rect 6751 263238 6797 263250
rect 6865 263238 6911 263250
rect 6961 263238 7007 263250
rect 7075 263238 7121 263250
rect 7171 263238 7217 263250
rect 7285 263238 7331 263250
rect 7381 263238 7427 263250
rect 7495 263238 7541 263250
rect 7591 263238 7637 263250
rect 7705 263238 7751 263250
rect 7801 263238 7847 263250
rect 7915 263238 7961 263250
rect 8011 263238 8057 263250
rect 8125 263238 8171 263250
rect 8221 263238 8267 263250
rect 8335 263238 8381 263250
rect 8431 263238 8477 263250
rect 8545 263238 8591 263250
rect 8641 263238 8687 263250
rect 8755 263238 8801 263250
rect 8851 263238 8897 263250
rect 8965 263238 9011 263250
rect 9061 263238 9107 263250
rect 9175 263238 9221 263250
rect 9271 263238 9317 263250
rect 9385 263238 9431 263250
rect 9481 263238 9527 263250
rect 9595 263238 9641 263250
rect 9691 263238 9737 263250
rect 9805 263238 9851 263250
rect 9901 263238 9947 263250
rect 10015 263238 10061 263250
rect 10111 263238 10157 263250
rect 10225 263238 10271 263250
rect 10321 263238 10367 263250
rect 10435 263238 10481 263250
rect 10531 263238 10577 263250
rect 10645 263238 10691 263250
rect 10741 263238 10787 263250
rect 10855 263238 10901 263250
rect 10951 263238 10997 263250
rect 11065 263238 11111 263250
rect 11161 263238 11207 263250
rect 11275 263238 11321 263250
rect 11371 263238 11417 263250
rect 11485 263238 11531 263250
rect 11581 263238 11627 263250
rect 11695 263238 11741 263250
rect 11791 263238 11837 263250
rect 11905 263238 11951 263250
rect 12001 263238 12047 263250
rect 12115 263238 12161 263250
rect 12211 263238 12257 263250
rect 12325 263238 12371 263250
rect 12421 263238 12467 263250
rect 12535 263238 12581 263250
rect 12631 263238 12677 263250
rect 12745 263238 12791 263250
rect 12841 263238 12887 263250
rect 12955 263238 13001 263250
rect 13051 263238 13097 263250
rect 13165 263238 13211 263250
rect 13261 263238 13307 263250
rect 13375 263238 13421 263250
rect 13471 263238 13517 263250
rect 13585 263238 13631 263250
rect 13681 263238 13727 263250
rect 13795 263238 13841 263250
rect 13891 263238 13937 263250
rect 14005 263238 14051 263250
rect 14101 263238 14147 263250
rect 14215 263238 14261 263250
rect 14311 263238 14357 263250
rect 14425 263238 14471 263250
rect 14521 263238 14567 263250
rect 14635 263238 14681 263250
rect 14731 263238 14777 263250
rect 14845 263238 14891 263250
rect 14941 263238 14987 263250
rect 15055 263238 15101 263250
rect 15151 263238 15197 263250
rect 15265 263238 15311 263250
rect 15361 263238 15407 263250
rect 15475 263238 15521 263250
rect 15571 263238 15617 263250
rect 15685 263238 15731 263250
rect 15781 263238 15827 263250
rect 15895 263238 15941 263250
rect 15991 263238 16037 263250
rect 16105 263238 16151 263250
rect 16201 263238 16247 263250
rect 16315 263238 16361 263250
rect 16411 263238 16457 263250
rect 16525 263238 16571 263250
rect 16621 263238 16667 263250
rect 16735 263238 16781 263250
rect 16831 263238 16877 263250
rect 16945 263238 16991 263250
rect 17041 263238 17087 263250
rect 17155 263238 17201 263250
rect 17251 263238 17297 263250
rect 17365 263238 17411 263250
rect 17461 263238 17507 263250
rect 17575 263238 17621 263250
rect 17671 263238 17717 263250
rect 17785 263238 17831 263250
rect 17881 263238 17927 263250
rect 17995 263238 18041 263250
rect 18091 263238 18137 263250
rect 18205 263238 18251 263250
rect 18301 263238 18347 263250
rect 18415 263238 18461 263250
rect 18511 263238 18557 263250
rect 18625 263238 18671 263250
rect 18721 263238 18767 263250
rect 18835 263238 18881 263250
rect 18931 263238 18977 263250
rect 19045 263238 19091 263250
rect 19141 263238 19187 263250
rect 19255 263238 19301 263250
rect 19351 263238 19397 263250
rect 19465 263238 19511 263250
rect 19561 263238 19607 263250
rect 19675 263238 19721 263250
rect 19771 263238 19817 263250
rect 19885 263238 19931 263250
rect 19981 263238 20027 263250
rect 20095 263238 20141 263250
rect 20191 263238 20237 263250
rect 20305 263238 20351 263250
rect 20401 263238 20447 263250
rect 20515 263238 20561 263250
rect 20611 263238 20657 263250
rect 20725 263238 20771 263250
rect 20821 263238 20867 263250
rect 20935 263238 20981 263250
rect 21031 263238 21077 263250
rect 21145 263238 21191 263250
rect 21241 263238 21287 263250
rect 21355 263238 21401 263250
rect 21451 263238 21497 263250
rect 21565 263238 21611 263250
rect 21661 263238 21707 263250
rect 21775 263238 21821 263250
rect 21871 263238 21917 263250
rect 21985 263238 22031 263250
rect 22081 263238 22127 263250
rect 22195 263238 22241 263250
rect 22291 263238 22337 263250
rect 22405 263238 22451 263250
rect 22501 263238 22547 263250
rect 22615 263238 22661 263250
rect 22711 263238 22757 263250
rect 22825 263238 22871 263250
rect 22921 263238 22967 263250
rect 23035 263238 23081 263250
rect 23131 263238 23177 263250
rect 23245 263238 23291 263250
rect 23341 263238 23387 263250
rect 23455 263238 23501 263250
rect 23551 263238 23597 263250
rect 23665 263238 23711 263250
rect 23761 263238 23807 263250
rect 23875 263238 23921 263250
rect 23971 263238 24017 263250
rect 24085 263238 24131 263250
rect 24181 263238 24227 263250
rect 24295 263238 24341 263250
rect 24391 263238 24437 263250
rect 24505 263238 24551 263250
rect 24601 263238 24647 263250
rect 24715 263238 24761 263250
rect 24811 263238 24857 263250
rect 24925 263238 24971 263250
rect 25021 263238 25067 263250
rect 25135 263238 25181 263250
rect 25231 263238 25277 263250
rect 25345 263238 25391 263250
rect 25441 263238 25487 263250
rect 25555 263238 25601 263250
rect 25651 263238 25697 263250
rect 25765 263238 25811 263250
rect 25861 263238 25907 263250
rect 25975 263238 26021 263250
rect 26071 263238 26117 263250
rect 26185 263238 26231 263250
rect 26281 263238 26327 263250
rect 26395 263238 26441 263250
rect 26491 263238 26537 263250
rect 26605 263238 26651 263250
rect 26701 263238 26747 263250
rect 26815 263238 26861 263250
rect 26911 263238 26957 263250
rect 27025 263238 27071 263250
rect 27121 263238 27167 263250
rect 27235 263238 27281 263250
rect 27331 263238 27423 263250
rect -3797 263204 -3751 263210
rect -3377 263204 -3331 263210
rect -2957 263204 -2911 263210
rect -2537 263204 -2491 263210
rect -2117 263204 -2071 263210
rect -1697 263204 -1651 263210
rect -1277 263204 -1231 263210
rect -857 263204 -811 263210
rect -437 263204 -391 263210
rect -17 263204 29 263210
rect 403 263204 449 263210
rect 823 263204 869 263210
rect 1243 263204 1289 263210
rect 1663 263204 1709 263210
rect 2083 263204 2129 263210
rect 2503 263204 2549 263210
rect 2923 263204 2969 263210
rect 3343 263204 3389 263210
rect 3763 263204 3809 263210
rect 4183 263204 4229 263210
rect 4603 263204 4649 263210
rect 5023 263204 5069 263210
rect 5443 263204 5489 263210
rect 5863 263204 5909 263210
rect 6283 263204 6329 263210
rect 6703 263204 6749 263210
rect 7123 263204 7169 263210
rect 7543 263204 7589 263210
rect 7963 263204 8009 263210
rect 8383 263204 8429 263210
rect 8803 263204 8849 263210
rect 9223 263204 9269 263210
rect 9643 263204 9689 263210
rect 10063 263204 10109 263210
rect 10483 263204 10529 263210
rect 10903 263204 10949 263210
rect 11323 263204 11369 263210
rect 11743 263204 11789 263210
rect 12163 263204 12209 263210
rect 12583 263204 12629 263210
rect 13003 263204 13049 263210
rect 13423 263204 13469 263210
rect 13843 263204 13889 263210
rect 14263 263204 14309 263210
rect 14683 263204 14729 263210
rect 15103 263204 15149 263210
rect 15523 263204 15569 263210
rect 15943 263204 15989 263210
rect 16363 263204 16409 263210
rect 16783 263204 16829 263210
rect 17203 263204 17249 263210
rect 17623 263204 17669 263210
rect 18043 263204 18089 263210
rect 18463 263204 18509 263210
rect 18883 263204 18929 263210
rect 19303 263204 19349 263210
rect 19723 263204 19769 263210
rect 20143 263204 20189 263210
rect 20563 263204 20609 263210
rect 20983 263204 21029 263210
rect 21403 263204 21449 263210
rect 21823 263204 21869 263210
rect 22243 263204 22289 263210
rect 22663 263204 22709 263210
rect 23083 263204 23129 263210
rect 23503 263204 23549 263210
rect 23923 263204 23969 263210
rect 24343 263204 24389 263210
rect 24763 263204 24809 263210
rect 25183 263204 25229 263210
rect 25603 263204 25649 263210
rect 26023 263204 26069 263210
rect 26443 263204 26489 263210
rect 26863 263204 26909 263210
rect 27283 263204 27329 263210
rect -3803 263198 -3745 263204
rect -3383 263198 -3325 263204
rect -2963 263198 -2905 263204
rect -2543 263198 -2485 263204
rect -2123 263198 -2065 263204
rect -1703 263198 -1645 263204
rect -1283 263198 -1225 263204
rect -863 263198 -805 263204
rect -443 263198 -385 263204
rect -23 263198 35 263204
rect 397 263198 455 263204
rect 817 263198 875 263204
rect 1237 263198 1295 263204
rect 1657 263198 1715 263204
rect 2077 263198 2135 263204
rect 2497 263198 2555 263204
rect 2917 263198 2975 263204
rect 3337 263198 3395 263204
rect 3757 263198 3815 263204
rect 4177 263198 4235 263204
rect 4597 263198 4655 263204
rect 5017 263198 5075 263204
rect 5437 263198 5495 263204
rect 5857 263198 5915 263204
rect 6277 263198 6335 263204
rect 6697 263198 6755 263204
rect 7117 263198 7175 263204
rect 7537 263198 7595 263204
rect 7957 263198 8015 263204
rect 8377 263198 8435 263204
rect 8797 263198 8855 263204
rect 9217 263198 9275 263204
rect 9637 263198 9695 263204
rect 10057 263198 10115 263204
rect 10477 263198 10535 263204
rect 10897 263198 10955 263204
rect 11317 263198 11375 263204
rect 11737 263198 11795 263204
rect 12157 263198 12215 263204
rect 12577 263198 12635 263204
rect 12997 263198 13055 263204
rect 13417 263198 13475 263204
rect 13837 263198 13895 263204
rect 14257 263198 14315 263204
rect 14677 263198 14735 263204
rect 15097 263198 15155 263204
rect 15517 263198 15575 263204
rect 15937 263198 15995 263204
rect 16357 263198 16415 263204
rect 16777 263198 16835 263204
rect 17197 263198 17255 263204
rect 17617 263198 17675 263204
rect 18037 263198 18095 263204
rect 18457 263198 18515 263204
rect 18877 263198 18935 263204
rect 19297 263198 19355 263204
rect 19717 263198 19775 263204
rect 20137 263198 20195 263204
rect 20557 263198 20615 263204
rect 20977 263198 21035 263204
rect 21397 263198 21455 263204
rect 21817 263198 21875 263204
rect 22237 263198 22295 263204
rect 22657 263198 22715 263204
rect 23077 263198 23135 263204
rect 23497 263198 23555 263204
rect 23917 263198 23975 263204
rect 24337 263198 24395 263204
rect 24757 263198 24815 263204
rect 25177 263198 25235 263204
rect 25597 263198 25655 263204
rect 26017 263198 26075 263204
rect 26437 263198 26495 263204
rect 26857 263198 26915 263204
rect 27277 263198 27335 263204
rect -5008 263056 -3791 263198
rect -3757 263056 -3371 263198
rect -3337 263056 -2951 263198
rect -2917 263056 -2531 263198
rect -2497 263056 -2111 263198
rect -2077 263056 -1691 263198
rect -1657 263056 -1271 263198
rect -1237 263056 -851 263198
rect -817 263056 -431 263198
rect -397 263056 -11 263198
rect 23 263056 409 263198
rect 443 263056 829 263198
rect 863 263056 1249 263198
rect 1283 263056 1669 263198
rect 1703 263056 2089 263198
rect 2123 263056 2509 263198
rect 2543 263056 2929 263198
rect 2963 263056 3349 263198
rect 3383 263056 3769 263198
rect 3803 263056 4189 263198
rect 4223 263056 4609 263198
rect 4643 263056 5029 263198
rect 5063 263056 5449 263198
rect 5483 263056 5869 263198
rect 5903 263056 6289 263198
rect 6323 263056 6709 263198
rect 6743 263056 7129 263198
rect 7163 263056 7549 263198
rect 7583 263056 7969 263198
rect 8003 263056 8389 263198
rect 8423 263056 8809 263198
rect 8843 263056 9229 263198
rect 9263 263056 9649 263198
rect 9683 263056 10069 263198
rect 10103 263056 10489 263198
rect 10523 263056 10909 263198
rect 10943 263056 11329 263198
rect 11363 263056 11749 263198
rect 11783 263056 12169 263198
rect 12203 263056 12589 263198
rect 12623 263056 13009 263198
rect 13043 263056 13429 263198
rect 13463 263056 13849 263198
rect 13883 263056 14269 263198
rect 14303 263056 14689 263198
rect 14723 263056 15109 263198
rect 15143 263056 15529 263198
rect 15563 263056 15949 263198
rect 15983 263056 16369 263198
rect 16403 263056 16789 263198
rect 16823 263056 17209 263198
rect 17243 263056 17629 263198
rect 17663 263056 18049 263198
rect 18083 263056 18469 263198
rect 18503 263056 18889 263198
rect 18923 263056 19309 263198
rect 19343 263056 19729 263198
rect 19763 263056 20149 263198
rect 20183 263056 20569 263198
rect 20603 263056 20989 263198
rect 21023 263056 21409 263198
rect 21443 263056 21829 263198
rect 21863 263056 22249 263198
rect 22283 263056 22669 263198
rect 22703 263056 23089 263198
rect 23123 263056 23509 263198
rect 23543 263056 23929 263198
rect 23963 263056 24349 263198
rect 24383 263056 24769 263198
rect 24803 263056 25189 263198
rect 25223 263056 25609 263198
rect 25643 263056 26029 263198
rect 26063 263056 26449 263198
rect 26483 263056 26869 263198
rect 26903 263056 27289 263198
rect 27323 263158 27335 263198
rect 27323 263096 27329 263158
rect 27323 263056 27335 263096
rect -5008 262184 -4244 263056
rect -3803 263050 -3745 263056
rect -3383 263050 -3325 263056
rect -2963 263050 -2905 263056
rect -2543 263050 -2485 263056
rect -2123 263050 -2065 263056
rect -1703 263050 -1645 263056
rect -1283 263050 -1225 263056
rect -863 263050 -805 263056
rect -443 263050 -385 263056
rect -23 263050 35 263056
rect 397 263050 455 263056
rect 817 263050 875 263056
rect 1237 263050 1295 263056
rect 1657 263050 1715 263056
rect 2077 263050 2135 263056
rect 2497 263050 2555 263056
rect 2917 263050 2975 263056
rect 3337 263050 3395 263056
rect 3757 263050 3815 263056
rect 4177 263050 4235 263056
rect 4597 263050 4655 263056
rect 5017 263050 5075 263056
rect 5437 263050 5495 263056
rect 5857 263050 5915 263056
rect 6277 263050 6335 263056
rect 6697 263050 6755 263056
rect 7117 263050 7175 263056
rect 7537 263050 7595 263056
rect 7957 263050 8015 263056
rect 8377 263050 8435 263056
rect 8797 263050 8855 263056
rect 9217 263050 9275 263056
rect 9637 263050 9695 263056
rect 10057 263050 10115 263056
rect 10477 263050 10535 263056
rect 10897 263050 10955 263056
rect 11317 263050 11375 263056
rect 11737 263050 11795 263056
rect 12157 263050 12215 263056
rect 12577 263050 12635 263056
rect 12997 263050 13055 263056
rect 13417 263050 13475 263056
rect 13837 263050 13895 263056
rect 14257 263050 14315 263056
rect 14677 263050 14735 263056
rect 15097 263050 15155 263056
rect 15517 263050 15575 263056
rect 15937 263050 15995 263056
rect 16357 263050 16415 263056
rect 16777 263050 16835 263056
rect 17197 263050 17255 263056
rect 17617 263050 17675 263056
rect 18037 263050 18095 263056
rect 18457 263050 18515 263056
rect 18877 263050 18935 263056
rect 19297 263050 19355 263056
rect 19717 263050 19775 263056
rect 20137 263050 20195 263056
rect 20557 263050 20615 263056
rect 20977 263050 21035 263056
rect 21397 263050 21455 263056
rect 21817 263050 21875 263056
rect 22237 263050 22295 263056
rect 22657 263050 22715 263056
rect 23077 263050 23135 263056
rect 23497 263050 23555 263056
rect 23917 263050 23975 263056
rect 24337 263050 24395 263056
rect 24757 263050 24815 263056
rect 25177 263050 25235 263056
rect 25597 263050 25655 263056
rect 26017 263050 26075 263056
rect 26437 263050 26495 263056
rect 26857 263050 26915 263056
rect 27277 263050 27335 263056
rect -3797 263044 -3751 263050
rect -3377 263044 -3331 263050
rect -2957 263044 -2911 263050
rect -2537 263044 -2491 263050
rect -2117 263044 -2071 263050
rect -1697 263044 -1651 263050
rect -1277 263044 -1231 263050
rect -857 263044 -811 263050
rect -437 263044 -391 263050
rect -17 263044 29 263050
rect 403 263044 449 263050
rect 823 263044 869 263050
rect 1243 263044 1289 263050
rect 1663 263044 1709 263050
rect 2083 263044 2129 263050
rect 2503 263044 2549 263050
rect 2923 263044 2969 263050
rect 3343 263044 3389 263050
rect 3763 263044 3809 263050
rect 4183 263044 4229 263050
rect 4603 263044 4649 263050
rect 5023 263044 5069 263050
rect 5443 263044 5489 263050
rect 5863 263044 5909 263050
rect 6283 263044 6329 263050
rect 6703 263044 6749 263050
rect 7123 263044 7169 263050
rect 7543 263044 7589 263050
rect 7963 263044 8009 263050
rect 8383 263044 8429 263050
rect 8803 263044 8849 263050
rect 9223 263044 9269 263050
rect 9643 263044 9689 263050
rect 10063 263044 10109 263050
rect 10483 263044 10529 263050
rect 10903 263044 10949 263050
rect 11323 263044 11369 263050
rect 11743 263044 11789 263050
rect 12163 263044 12209 263050
rect 12583 263044 12629 263050
rect 13003 263044 13049 263050
rect 13423 263044 13469 263050
rect 13843 263044 13889 263050
rect 14263 263044 14309 263050
rect 14683 263044 14729 263050
rect 15103 263044 15149 263050
rect 15523 263044 15569 263050
rect 15943 263044 15989 263050
rect 16363 263044 16409 263050
rect 16783 263044 16829 263050
rect 17203 263044 17249 263050
rect 17623 263044 17669 263050
rect 18043 263044 18089 263050
rect 18463 263044 18509 263050
rect 18883 263044 18929 263050
rect 19303 263044 19349 263050
rect 19723 263044 19769 263050
rect 20143 263044 20189 263050
rect 20563 263044 20609 263050
rect 20983 263044 21029 263050
rect 21403 263044 21449 263050
rect 21823 263044 21869 263050
rect 22243 263044 22289 263050
rect 22663 263044 22709 263050
rect 23083 263044 23129 263050
rect 23503 263044 23549 263050
rect 23923 263044 23969 263050
rect 24343 263044 24389 263050
rect 24763 263044 24809 263050
rect 25183 263044 25229 263050
rect 25603 263044 25649 263050
rect 26023 263044 26069 263050
rect 26443 263044 26489 263050
rect 26863 263044 26909 263050
rect 27283 263044 27329 263050
rect 27375 263016 27423 263238
rect -4070 263004 -4009 263016
rect -3959 263004 -3913 263016
rect -3845 263004 -3799 263016
rect -3749 263004 -3703 263016
rect -3635 263004 -3589 263016
rect -3539 263004 -3493 263016
rect -3425 263004 -3379 263016
rect -3329 263004 -3283 263016
rect -3215 263004 -3169 263016
rect -3119 263004 -3073 263016
rect -3005 263004 -2959 263016
rect -2909 263004 -2863 263016
rect -2795 263004 -2749 263016
rect -2699 263004 -2653 263016
rect -2585 263004 -2539 263016
rect -2489 263004 -2443 263016
rect -2375 263004 -2329 263016
rect -2279 263004 -2233 263016
rect -2165 263004 -2119 263016
rect -2069 263004 -2023 263016
rect -1955 263004 -1909 263016
rect -1859 263004 -1813 263016
rect -1745 263004 -1699 263016
rect -1649 263004 -1603 263016
rect -1535 263004 -1489 263016
rect -1439 263004 -1393 263016
rect -1325 263004 -1279 263016
rect -1229 263004 -1183 263016
rect -1115 263004 -1069 263016
rect -1019 263004 -973 263016
rect -905 263004 -859 263016
rect -809 263004 -763 263016
rect -695 263004 -649 263016
rect -599 263004 -553 263016
rect -485 263004 -439 263016
rect -389 263004 -343 263016
rect -275 263004 -229 263016
rect -179 263004 -133 263016
rect -65 263004 -19 263016
rect 31 263004 77 263016
rect 145 263004 191 263016
rect 241 263004 287 263016
rect 355 263004 401 263016
rect 451 263004 497 263016
rect 565 263004 611 263016
rect 661 263004 707 263016
rect 775 263004 821 263016
rect 871 263004 917 263016
rect 985 263004 1031 263016
rect 1081 263004 1127 263016
rect 1195 263004 1241 263016
rect 1291 263004 1337 263016
rect 1405 263004 1451 263016
rect 1501 263004 1547 263016
rect 1615 263004 1661 263016
rect 1711 263004 1757 263016
rect 1825 263004 1871 263016
rect 1921 263004 1967 263016
rect 2035 263004 2081 263016
rect 2131 263004 2177 263016
rect 2245 263004 2291 263016
rect 2341 263004 2387 263016
rect 2455 263004 2501 263016
rect 2551 263004 2597 263016
rect 2665 263004 2711 263016
rect 2761 263004 2807 263016
rect 2875 263004 2921 263016
rect 2971 263004 3017 263016
rect 3085 263004 3131 263016
rect 3181 263004 3227 263016
rect 3295 263004 3341 263016
rect 3391 263004 3437 263016
rect 3505 263004 3551 263016
rect 3601 263004 3647 263016
rect 3715 263004 3761 263016
rect 3811 263004 3857 263016
rect 3925 263004 3971 263016
rect 4021 263004 4067 263016
rect 4135 263004 4181 263016
rect 4231 263004 4277 263016
rect 4345 263004 4391 263016
rect 4441 263004 4487 263016
rect 4555 263004 4601 263016
rect 4651 263004 4697 263016
rect 4765 263004 4811 263016
rect 4861 263004 4907 263016
rect 4975 263004 5021 263016
rect 5071 263004 5117 263016
rect 5185 263004 5231 263016
rect 5281 263004 5327 263016
rect 5395 263004 5441 263016
rect 5491 263004 5537 263016
rect 5605 263004 5651 263016
rect 5701 263004 5747 263016
rect 5815 263004 5861 263016
rect 5911 263004 5957 263016
rect 6025 263004 6071 263016
rect 6121 263004 6167 263016
rect 6235 263004 6281 263016
rect 6331 263004 6377 263016
rect 6445 263004 6491 263016
rect 6541 263004 6587 263016
rect 6655 263004 6701 263016
rect 6751 263004 6797 263016
rect 6865 263004 6911 263016
rect 6961 263004 7007 263016
rect 7075 263004 7121 263016
rect 7171 263004 7217 263016
rect 7285 263004 7331 263016
rect 7381 263004 7427 263016
rect 7495 263004 7541 263016
rect 7591 263004 7637 263016
rect 7705 263004 7751 263016
rect 7801 263004 7847 263016
rect 7915 263004 7961 263016
rect 8011 263004 8057 263016
rect 8125 263004 8171 263016
rect 8221 263004 8267 263016
rect 8335 263004 8381 263016
rect 8431 263004 8477 263016
rect 8545 263004 8591 263016
rect 8641 263004 8687 263016
rect 8755 263004 8801 263016
rect 8851 263004 8897 263016
rect 8965 263004 9011 263016
rect 9061 263004 9107 263016
rect 9175 263004 9221 263016
rect 9271 263004 9317 263016
rect 9385 263004 9431 263016
rect 9481 263004 9527 263016
rect 9595 263004 9641 263016
rect 9691 263004 9737 263016
rect 9805 263004 9851 263016
rect 9901 263004 9947 263016
rect 10015 263004 10061 263016
rect 10111 263004 10157 263016
rect 10225 263004 10271 263016
rect 10321 263004 10367 263016
rect 10435 263004 10481 263016
rect 10531 263004 10577 263016
rect 10645 263004 10691 263016
rect 10741 263004 10787 263016
rect 10855 263004 10901 263016
rect 10951 263004 10997 263016
rect 11065 263004 11111 263016
rect 11161 263004 11207 263016
rect 11275 263004 11321 263016
rect 11371 263004 11417 263016
rect 11485 263004 11531 263016
rect 11581 263004 11627 263016
rect 11695 263004 11741 263016
rect 11791 263004 11837 263016
rect 11905 263004 11951 263016
rect 12001 263004 12047 263016
rect 12115 263004 12161 263016
rect 12211 263004 12257 263016
rect 12325 263004 12371 263016
rect 12421 263004 12467 263016
rect 12535 263004 12581 263016
rect 12631 263004 12677 263016
rect 12745 263004 12791 263016
rect 12841 263004 12887 263016
rect 12955 263004 13001 263016
rect 13051 263004 13097 263016
rect 13165 263004 13211 263016
rect 13261 263004 13307 263016
rect 13375 263004 13421 263016
rect 13471 263004 13517 263016
rect 13585 263004 13631 263016
rect 13681 263004 13727 263016
rect 13795 263004 13841 263016
rect 13891 263004 13937 263016
rect 14005 263004 14051 263016
rect 14101 263004 14147 263016
rect 14215 263004 14261 263016
rect 14311 263004 14357 263016
rect 14425 263004 14471 263016
rect 14521 263004 14567 263016
rect 14635 263004 14681 263016
rect 14731 263004 14777 263016
rect 14845 263004 14891 263016
rect 14941 263004 14987 263016
rect 15055 263004 15101 263016
rect 15151 263004 15197 263016
rect 15265 263004 15311 263016
rect 15361 263004 15407 263016
rect 15475 263004 15521 263016
rect 15571 263004 15617 263016
rect 15685 263004 15731 263016
rect 15781 263004 15827 263016
rect 15895 263004 15941 263016
rect 15991 263004 16037 263016
rect 16105 263004 16151 263016
rect 16201 263004 16247 263016
rect 16315 263004 16361 263016
rect 16411 263004 16457 263016
rect 16525 263004 16571 263016
rect 16621 263004 16667 263016
rect 16735 263004 16781 263016
rect 16831 263004 16877 263016
rect 16945 263004 16991 263016
rect 17041 263004 17087 263016
rect 17155 263004 17201 263016
rect 17251 263004 17297 263016
rect 17365 263004 17411 263016
rect 17461 263004 17507 263016
rect 17575 263004 17621 263016
rect 17671 263004 17717 263016
rect 17785 263004 17831 263016
rect 17881 263004 17927 263016
rect 17995 263004 18041 263016
rect 18091 263004 18137 263016
rect 18205 263004 18251 263016
rect 18301 263004 18347 263016
rect 18415 263004 18461 263016
rect 18511 263004 18557 263016
rect 18625 263004 18671 263016
rect 18721 263004 18767 263016
rect 18835 263004 18881 263016
rect 18931 263004 18977 263016
rect 19045 263004 19091 263016
rect 19141 263004 19187 263016
rect 19255 263004 19301 263016
rect 19351 263004 19397 263016
rect 19465 263004 19511 263016
rect 19561 263004 19607 263016
rect 19675 263004 19721 263016
rect 19771 263004 19817 263016
rect 19885 263004 19931 263016
rect 19981 263004 20027 263016
rect 20095 263004 20141 263016
rect 20191 263004 20237 263016
rect 20305 263004 20351 263016
rect 20401 263004 20447 263016
rect 20515 263004 20561 263016
rect 20611 263004 20657 263016
rect 20725 263004 20771 263016
rect 20821 263004 20867 263016
rect 20935 263004 20981 263016
rect 21031 263004 21077 263016
rect 21145 263004 21191 263016
rect 21241 263004 21287 263016
rect 21355 263004 21401 263016
rect 21451 263004 21497 263016
rect 21565 263004 21611 263016
rect 21661 263004 21707 263016
rect 21775 263004 21821 263016
rect 21871 263004 21917 263016
rect 21985 263004 22031 263016
rect 22081 263004 22127 263016
rect 22195 263004 22241 263016
rect 22291 263004 22337 263016
rect 22405 263004 22451 263016
rect 22501 263004 22547 263016
rect 22615 263004 22661 263016
rect 22711 263004 22757 263016
rect 22825 263004 22871 263016
rect 22921 263004 22967 263016
rect 23035 263004 23081 263016
rect 23131 263004 23177 263016
rect 23245 263004 23291 263016
rect 23341 263004 23387 263016
rect 23455 263004 23501 263016
rect 23551 263004 23597 263016
rect 23665 263004 23711 263016
rect 23761 263004 23807 263016
rect 23875 263004 23921 263016
rect 23971 263004 24017 263016
rect 24085 263004 24131 263016
rect 24181 263004 24227 263016
rect 24295 263004 24341 263016
rect 24391 263004 24437 263016
rect 24505 263004 24551 263016
rect 24601 263004 24647 263016
rect 24715 263004 24761 263016
rect 24811 263004 24857 263016
rect 24925 263004 24971 263016
rect 25021 263004 25067 263016
rect 25135 263004 25181 263016
rect 25231 263004 25277 263016
rect 25345 263004 25391 263016
rect 25441 263004 25487 263016
rect 25555 263004 25601 263016
rect 25651 263004 25697 263016
rect 25765 263004 25811 263016
rect 25861 263004 25907 263016
rect 25975 263004 26021 263016
rect 26071 263004 26117 263016
rect 26185 263004 26231 263016
rect 26281 263004 26327 263016
rect 26395 263004 26441 263016
rect 26491 263004 26537 263016
rect 26605 263004 26651 263016
rect 26701 263004 26747 263016
rect 26815 263004 26861 263016
rect 26911 263004 26957 263016
rect 27025 263004 27071 263016
rect 27121 263004 27167 263016
rect 27235 263004 27281 263016
rect 27331 263004 27423 263016
rect -4015 262228 -4005 263004
rect -3963 262228 -3953 263004
rect -3805 262228 -3795 263004
rect -3753 262228 -3743 263004
rect -3595 262228 -3585 263004
rect -3543 262228 -3533 263004
rect -3385 262228 -3375 263004
rect -3333 262228 -3323 263004
rect -3175 262228 -3165 263004
rect -3123 262228 -3113 263004
rect -2965 262228 -2955 263004
rect -2913 262228 -2903 263004
rect -2755 262228 -2745 263004
rect -2703 262228 -2693 263004
rect -2545 262228 -2535 263004
rect -2493 262228 -2483 263004
rect -2335 262228 -2325 263004
rect -2283 262228 -2273 263004
rect -2125 262228 -2115 263004
rect -2073 262228 -2063 263004
rect -1915 262228 -1905 263004
rect -1863 262228 -1853 263004
rect -1705 262228 -1695 263004
rect -1653 262228 -1643 263004
rect -1495 262228 -1485 263004
rect -1443 262228 -1433 263004
rect -1285 262228 -1275 263004
rect -1233 262228 -1223 263004
rect -1075 262228 -1065 263004
rect -1023 262228 -1013 263004
rect -865 262228 -855 263004
rect -813 262228 -803 263004
rect -655 262228 -645 263004
rect -603 262228 -593 263004
rect -445 262228 -435 263004
rect -393 262228 -383 263004
rect -235 262228 -225 263004
rect -183 262228 -173 263004
rect -25 262228 -15 263004
rect 27 262228 37 263004
rect 185 262228 195 263004
rect 237 262228 247 263004
rect 395 262228 405 263004
rect 447 262228 457 263004
rect 605 262228 615 263004
rect 657 262228 667 263004
rect 815 262228 825 263004
rect 867 262228 877 263004
rect 1025 262228 1035 263004
rect 1077 262228 1087 263004
rect 1235 262228 1245 263004
rect 1287 262228 1297 263004
rect 1445 262228 1455 263004
rect 1497 262228 1507 263004
rect 1655 262228 1665 263004
rect 1707 262228 1717 263004
rect 1865 262228 1875 263004
rect 1917 262228 1927 263004
rect 2075 262228 2085 263004
rect 2127 262228 2137 263004
rect 2285 262228 2295 263004
rect 2337 262228 2347 263004
rect 2495 262228 2505 263004
rect 2547 262228 2557 263004
rect 2705 262228 2715 263004
rect 2757 262228 2767 263004
rect 2915 262228 2925 263004
rect 2967 262228 2977 263004
rect 3125 262228 3135 263004
rect 3177 262228 3187 263004
rect 3335 262228 3345 263004
rect 3387 262228 3397 263004
rect 3545 262228 3555 263004
rect 3597 262228 3607 263004
rect 3755 262228 3765 263004
rect 3807 262228 3817 263004
rect 3965 262228 3975 263004
rect 4017 262228 4027 263004
rect 4175 262228 4185 263004
rect 4227 262228 4237 263004
rect 4385 262228 4395 263004
rect 4437 262228 4447 263004
rect 4595 262228 4605 263004
rect 4647 262228 4657 263004
rect 4805 262228 4815 263004
rect 4857 262228 4867 263004
rect 5015 262228 5025 263004
rect 5067 262228 5077 263004
rect 5225 262228 5235 263004
rect 5277 262228 5287 263004
rect 5435 262228 5445 263004
rect 5487 262228 5497 263004
rect 5645 262228 5655 263004
rect 5697 262228 5707 263004
rect 5855 262228 5865 263004
rect 5907 262228 5917 263004
rect 6065 262228 6075 263004
rect 6117 262228 6127 263004
rect 6275 262228 6285 263004
rect 6327 262228 6337 263004
rect 6485 262228 6495 263004
rect 6537 262228 6547 263004
rect 6695 262228 6705 263004
rect 6747 262228 6757 263004
rect 6905 262228 6915 263004
rect 6957 262228 6967 263004
rect 7115 262228 7125 263004
rect 7167 262228 7177 263004
rect 7325 262228 7335 263004
rect 7377 262228 7387 263004
rect 7535 262228 7545 263004
rect 7587 262228 7597 263004
rect 7745 262228 7755 263004
rect 7797 262228 7807 263004
rect 7955 262228 7965 263004
rect 8007 262228 8017 263004
rect 8165 262228 8175 263004
rect 8217 262228 8227 263004
rect 8375 262228 8385 263004
rect 8427 262228 8437 263004
rect 8585 262228 8595 263004
rect 8637 262228 8647 263004
rect 8795 262228 8805 263004
rect 8847 262228 8857 263004
rect 9005 262228 9015 263004
rect 9057 262228 9067 263004
rect 9215 262228 9225 263004
rect 9267 262228 9277 263004
rect 9425 262228 9435 263004
rect 9477 262228 9487 263004
rect 9635 262228 9645 263004
rect 9687 262228 9697 263004
rect 9845 262228 9855 263004
rect 9897 262228 9907 263004
rect 10055 262228 10065 263004
rect 10107 262228 10117 263004
rect 10265 262228 10275 263004
rect 10317 262228 10327 263004
rect 10475 262228 10485 263004
rect 10527 262228 10537 263004
rect 10685 262228 10695 263004
rect 10737 262228 10747 263004
rect 10895 262228 10905 263004
rect 10947 262228 10957 263004
rect 11105 262228 11115 263004
rect 11157 262228 11167 263004
rect 11315 262228 11325 263004
rect 11367 262228 11377 263004
rect 11525 262228 11535 263004
rect 11577 262228 11587 263004
rect 11735 262228 11745 263004
rect 11787 262228 11797 263004
rect 11945 262228 11955 263004
rect 11997 262228 12007 263004
rect 12155 262228 12165 263004
rect 12207 262228 12217 263004
rect 12365 262228 12375 263004
rect 12417 262228 12427 263004
rect 12575 262228 12585 263004
rect 12627 262228 12637 263004
rect 12785 262228 12795 263004
rect 12837 262228 12847 263004
rect 12995 262228 13005 263004
rect 13047 262228 13057 263004
rect 13205 262228 13215 263004
rect 13257 262228 13267 263004
rect 13415 262228 13425 263004
rect 13467 262228 13477 263004
rect 13625 262228 13635 263004
rect 13677 262228 13687 263004
rect 13835 262228 13845 263004
rect 13887 262228 13897 263004
rect 14045 262228 14055 263004
rect 14097 262228 14107 263004
rect 14255 262228 14265 263004
rect 14307 262228 14317 263004
rect 14465 262228 14475 263004
rect 14517 262228 14527 263004
rect 14675 262228 14685 263004
rect 14727 262228 14737 263004
rect 14885 262228 14895 263004
rect 14937 262228 14947 263004
rect 15095 262228 15105 263004
rect 15147 262228 15157 263004
rect 15305 262228 15315 263004
rect 15357 262228 15367 263004
rect 15515 262228 15525 263004
rect 15567 262228 15577 263004
rect 15725 262228 15735 263004
rect 15777 262228 15787 263004
rect 15935 262228 15945 263004
rect 15987 262228 15997 263004
rect 16145 262228 16155 263004
rect 16197 262228 16207 263004
rect 16355 262228 16365 263004
rect 16407 262228 16417 263004
rect 16565 262228 16575 263004
rect 16617 262228 16627 263004
rect 16775 262228 16785 263004
rect 16827 262228 16837 263004
rect 16985 262228 16995 263004
rect 17037 262228 17047 263004
rect 17195 262228 17205 263004
rect 17247 262228 17257 263004
rect 17405 262228 17415 263004
rect 17457 262228 17467 263004
rect 17615 262228 17625 263004
rect 17667 262228 17677 263004
rect 17825 262228 17835 263004
rect 17877 262228 17887 263004
rect 18035 262228 18045 263004
rect 18087 262228 18097 263004
rect 18245 262228 18255 263004
rect 18297 262228 18307 263004
rect 18455 262228 18465 263004
rect 18507 262228 18517 263004
rect 18665 262228 18675 263004
rect 18717 262228 18727 263004
rect 18875 262228 18885 263004
rect 18927 262228 18937 263004
rect 19085 262228 19095 263004
rect 19137 262228 19147 263004
rect 19295 262228 19305 263004
rect 19347 262228 19357 263004
rect 19505 262228 19515 263004
rect 19557 262228 19567 263004
rect 19715 262228 19725 263004
rect 19767 262228 19777 263004
rect 19925 262228 19935 263004
rect 19977 262228 19987 263004
rect 20135 262228 20145 263004
rect 20187 262228 20197 263004
rect 20345 262228 20355 263004
rect 20397 262228 20407 263004
rect 20555 262228 20565 263004
rect 20607 262228 20617 263004
rect 20765 262228 20775 263004
rect 20817 262228 20827 263004
rect 20975 262228 20985 263004
rect 21027 262228 21037 263004
rect 21185 262228 21195 263004
rect 21237 262228 21247 263004
rect 21395 262228 21405 263004
rect 21447 262228 21457 263004
rect 21605 262228 21615 263004
rect 21657 262228 21667 263004
rect 21815 262228 21825 263004
rect 21867 262228 21877 263004
rect 22025 262228 22035 263004
rect 22077 262228 22087 263004
rect 22235 262228 22245 263004
rect 22287 262228 22297 263004
rect 22445 262228 22455 263004
rect 22497 262228 22507 263004
rect 22655 262228 22665 263004
rect 22707 262228 22717 263004
rect 22865 262228 22875 263004
rect 22917 262228 22927 263004
rect 23075 262228 23085 263004
rect 23127 262228 23137 263004
rect 23285 262228 23295 263004
rect 23337 262228 23347 263004
rect 23495 262228 23505 263004
rect 23547 262228 23557 263004
rect 23705 262228 23715 263004
rect 23757 262228 23767 263004
rect 23915 262228 23925 263004
rect 23967 262228 23977 263004
rect 24125 262228 24135 263004
rect 24177 262228 24187 263004
rect 24335 262228 24345 263004
rect 24387 262228 24397 263004
rect 24545 262228 24555 263004
rect 24597 262228 24607 263004
rect 24755 262228 24765 263004
rect 24807 262228 24817 263004
rect 24965 262228 24975 263004
rect 25017 262228 25027 263004
rect 25175 262228 25185 263004
rect 25227 262228 25237 263004
rect 25385 262228 25395 263004
rect 25437 262228 25447 263004
rect 25595 262228 25605 263004
rect 25647 262228 25657 263004
rect 25805 262228 25815 263004
rect 25857 262228 25867 263004
rect 26015 262228 26025 263004
rect 26067 262228 26077 263004
rect 26225 262228 26235 263004
rect 26277 262228 26287 263004
rect 26435 262228 26445 263004
rect 26487 262228 26497 263004
rect 26645 262228 26655 263004
rect 26697 262228 26707 263004
rect 26855 262228 26865 263004
rect 26907 262228 26917 263004
rect 27065 262228 27075 263004
rect 27117 262228 27127 263004
rect 27275 262228 27285 263004
rect 27331 262228 27337 263004
rect 27371 262228 27423 263004
rect -4070 262216 -4009 262228
rect -3959 262216 -3913 262228
rect -3845 262216 -3799 262228
rect -3749 262216 -3703 262228
rect -3635 262216 -3589 262228
rect -3539 262216 -3493 262228
rect -3425 262216 -3379 262228
rect -3329 262216 -3283 262228
rect -3215 262216 -3169 262228
rect -3119 262216 -3073 262228
rect -3005 262216 -2959 262228
rect -2909 262216 -2863 262228
rect -2795 262216 -2749 262228
rect -2699 262216 -2653 262228
rect -2585 262216 -2539 262228
rect -2489 262216 -2443 262228
rect -2375 262216 -2329 262228
rect -2279 262216 -2233 262228
rect -2165 262216 -2119 262228
rect -2069 262216 -2023 262228
rect -1955 262216 -1909 262228
rect -1859 262216 -1813 262228
rect -1745 262216 -1699 262228
rect -1649 262216 -1603 262228
rect -1535 262216 -1489 262228
rect -1439 262216 -1393 262228
rect -1325 262216 -1279 262228
rect -1229 262216 -1183 262228
rect -1115 262216 -1069 262228
rect -1019 262216 -973 262228
rect -905 262216 -859 262228
rect -809 262216 -763 262228
rect -695 262216 -649 262228
rect -599 262216 -553 262228
rect -485 262216 -439 262228
rect -389 262216 -343 262228
rect -275 262216 -229 262228
rect -179 262216 -133 262228
rect -65 262216 -19 262228
rect 31 262216 77 262228
rect 145 262216 191 262228
rect 241 262216 287 262228
rect 355 262216 401 262228
rect 451 262216 497 262228
rect 565 262216 611 262228
rect 661 262216 707 262228
rect 775 262216 821 262228
rect 871 262216 917 262228
rect 985 262216 1031 262228
rect 1081 262216 1127 262228
rect 1195 262216 1241 262228
rect 1291 262216 1337 262228
rect 1405 262216 1451 262228
rect 1501 262216 1547 262228
rect 1615 262216 1661 262228
rect 1711 262216 1757 262228
rect 1825 262216 1871 262228
rect 1921 262216 1967 262228
rect 2035 262216 2081 262228
rect 2131 262216 2177 262228
rect 2245 262216 2291 262228
rect 2341 262216 2387 262228
rect 2455 262216 2501 262228
rect 2551 262216 2597 262228
rect 2665 262216 2711 262228
rect 2761 262216 2807 262228
rect 2875 262216 2921 262228
rect 2971 262216 3017 262228
rect 3085 262216 3131 262228
rect 3181 262216 3227 262228
rect 3295 262216 3341 262228
rect 3391 262216 3437 262228
rect 3505 262216 3551 262228
rect 3601 262216 3647 262228
rect 3715 262216 3761 262228
rect 3811 262216 3857 262228
rect 3925 262216 3971 262228
rect 4021 262216 4067 262228
rect 4135 262216 4181 262228
rect 4231 262216 4277 262228
rect 4345 262216 4391 262228
rect 4441 262216 4487 262228
rect 4555 262216 4601 262228
rect 4651 262216 4697 262228
rect 4765 262216 4811 262228
rect 4861 262216 4907 262228
rect 4975 262216 5021 262228
rect 5071 262216 5117 262228
rect 5185 262216 5231 262228
rect 5281 262216 5327 262228
rect 5395 262216 5441 262228
rect 5491 262216 5537 262228
rect 5605 262216 5651 262228
rect 5701 262216 5747 262228
rect 5815 262216 5861 262228
rect 5911 262216 5957 262228
rect 6025 262216 6071 262228
rect 6121 262216 6167 262228
rect 6235 262216 6281 262228
rect 6331 262216 6377 262228
rect 6445 262216 6491 262228
rect 6541 262216 6587 262228
rect 6655 262216 6701 262228
rect 6751 262216 6797 262228
rect 6865 262216 6911 262228
rect 6961 262216 7007 262228
rect 7075 262216 7121 262228
rect 7171 262216 7217 262228
rect 7285 262216 7331 262228
rect 7381 262216 7427 262228
rect 7495 262216 7541 262228
rect 7591 262216 7637 262228
rect 7705 262216 7751 262228
rect 7801 262216 7847 262228
rect 7915 262216 7961 262228
rect 8011 262216 8057 262228
rect 8125 262216 8171 262228
rect 8221 262216 8267 262228
rect 8335 262216 8381 262228
rect 8431 262216 8477 262228
rect 8545 262216 8591 262228
rect 8641 262216 8687 262228
rect 8755 262216 8801 262228
rect 8851 262216 8897 262228
rect 8965 262216 9011 262228
rect 9061 262216 9107 262228
rect 9175 262216 9221 262228
rect 9271 262216 9317 262228
rect 9385 262216 9431 262228
rect 9481 262216 9527 262228
rect 9595 262216 9641 262228
rect 9691 262216 9737 262228
rect 9805 262216 9851 262228
rect 9901 262216 9947 262228
rect 10015 262216 10061 262228
rect 10111 262216 10157 262228
rect 10225 262216 10271 262228
rect 10321 262216 10367 262228
rect 10435 262216 10481 262228
rect 10531 262216 10577 262228
rect 10645 262216 10691 262228
rect 10741 262216 10787 262228
rect 10855 262216 10901 262228
rect 10951 262216 10997 262228
rect 11065 262216 11111 262228
rect 11161 262216 11207 262228
rect 11275 262216 11321 262228
rect 11371 262216 11417 262228
rect 11485 262216 11531 262228
rect 11581 262216 11627 262228
rect 11695 262216 11741 262228
rect 11791 262216 11837 262228
rect 11905 262216 11951 262228
rect 12001 262216 12047 262228
rect 12115 262216 12161 262228
rect 12211 262216 12257 262228
rect 12325 262216 12371 262228
rect 12421 262216 12467 262228
rect 12535 262216 12581 262228
rect 12631 262216 12677 262228
rect 12745 262216 12791 262228
rect 12841 262216 12887 262228
rect 12955 262216 13001 262228
rect 13051 262216 13097 262228
rect 13165 262216 13211 262228
rect 13261 262216 13307 262228
rect 13375 262216 13421 262228
rect 13471 262216 13517 262228
rect 13585 262216 13631 262228
rect 13681 262216 13727 262228
rect 13795 262216 13841 262228
rect 13891 262216 13937 262228
rect 14005 262216 14051 262228
rect 14101 262216 14147 262228
rect 14215 262216 14261 262228
rect 14311 262216 14357 262228
rect 14425 262216 14471 262228
rect 14521 262216 14567 262228
rect 14635 262216 14681 262228
rect 14731 262216 14777 262228
rect 14845 262216 14891 262228
rect 14941 262216 14987 262228
rect 15055 262216 15101 262228
rect 15151 262216 15197 262228
rect 15265 262216 15311 262228
rect 15361 262216 15407 262228
rect 15475 262216 15521 262228
rect 15571 262216 15617 262228
rect 15685 262216 15731 262228
rect 15781 262216 15827 262228
rect 15895 262216 15941 262228
rect 15991 262216 16037 262228
rect 16105 262216 16151 262228
rect 16201 262216 16247 262228
rect 16315 262216 16361 262228
rect 16411 262216 16457 262228
rect 16525 262216 16571 262228
rect 16621 262216 16667 262228
rect 16735 262216 16781 262228
rect 16831 262216 16877 262228
rect 16945 262216 16991 262228
rect 17041 262216 17087 262228
rect 17155 262216 17201 262228
rect 17251 262216 17297 262228
rect 17365 262216 17411 262228
rect 17461 262216 17507 262228
rect 17575 262216 17621 262228
rect 17671 262216 17717 262228
rect 17785 262216 17831 262228
rect 17881 262216 17927 262228
rect 17995 262216 18041 262228
rect 18091 262216 18137 262228
rect 18205 262216 18251 262228
rect 18301 262216 18347 262228
rect 18415 262216 18461 262228
rect 18511 262216 18557 262228
rect 18625 262216 18671 262228
rect 18721 262216 18767 262228
rect 18835 262216 18881 262228
rect 18931 262216 18977 262228
rect 19045 262216 19091 262228
rect 19141 262216 19187 262228
rect 19255 262216 19301 262228
rect 19351 262216 19397 262228
rect 19465 262216 19511 262228
rect 19561 262216 19607 262228
rect 19675 262216 19721 262228
rect 19771 262216 19817 262228
rect 19885 262216 19931 262228
rect 19981 262216 20027 262228
rect 20095 262216 20141 262228
rect 20191 262216 20237 262228
rect 20305 262216 20351 262228
rect 20401 262216 20447 262228
rect 20515 262216 20561 262228
rect 20611 262216 20657 262228
rect 20725 262216 20771 262228
rect 20821 262216 20867 262228
rect 20935 262216 20981 262228
rect 21031 262216 21077 262228
rect 21145 262216 21191 262228
rect 21241 262216 21287 262228
rect 21355 262216 21401 262228
rect 21451 262216 21497 262228
rect 21565 262216 21611 262228
rect 21661 262216 21707 262228
rect 21775 262216 21821 262228
rect 21871 262216 21917 262228
rect 21985 262216 22031 262228
rect 22081 262216 22127 262228
rect 22195 262216 22241 262228
rect 22291 262216 22337 262228
rect 22405 262216 22451 262228
rect 22501 262216 22547 262228
rect 22615 262216 22661 262228
rect 22711 262216 22757 262228
rect 22825 262216 22871 262228
rect 22921 262216 22967 262228
rect 23035 262216 23081 262228
rect 23131 262216 23177 262228
rect 23245 262216 23291 262228
rect 23341 262216 23387 262228
rect 23455 262216 23501 262228
rect 23551 262216 23597 262228
rect 23665 262216 23711 262228
rect 23761 262216 23807 262228
rect 23875 262216 23921 262228
rect 23971 262216 24017 262228
rect 24085 262216 24131 262228
rect 24181 262216 24227 262228
rect 24295 262216 24341 262228
rect 24391 262216 24437 262228
rect 24505 262216 24551 262228
rect 24601 262216 24647 262228
rect 24715 262216 24761 262228
rect 24811 262216 24857 262228
rect 24925 262216 24971 262228
rect 25021 262216 25067 262228
rect 25135 262216 25181 262228
rect 25231 262216 25277 262228
rect 25345 262216 25391 262228
rect 25441 262216 25487 262228
rect 25555 262216 25601 262228
rect 25651 262216 25697 262228
rect 25765 262216 25811 262228
rect 25861 262216 25907 262228
rect 25975 262216 26021 262228
rect 26071 262216 26117 262228
rect 26185 262216 26231 262228
rect 26281 262216 26327 262228
rect 26395 262216 26441 262228
rect 26491 262216 26537 262228
rect 26605 262216 26651 262228
rect 26701 262216 26747 262228
rect 26815 262216 26861 262228
rect 26911 262216 26957 262228
rect 27025 262216 27071 262228
rect 27121 262216 27167 262228
rect 27235 262216 27281 262228
rect 27331 262216 27423 262228
rect -5008 262178 27285 262184
rect -5008 262144 -4001 262178
rect -3905 262144 -3581 262178
rect -3485 262144 -3161 262178
rect -3065 262144 -2741 262178
rect -2645 262144 -2321 262178
rect -2225 262144 -1901 262178
rect -1805 262144 -1481 262178
rect -1385 262144 -1061 262178
rect -965 262144 -641 262178
rect -545 262144 -221 262178
rect -125 262144 199 262178
rect 295 262144 619 262178
rect 715 262144 1039 262178
rect 1135 262144 1459 262178
rect 1555 262144 1879 262178
rect 1975 262144 2299 262178
rect 2395 262144 2719 262178
rect 2815 262144 3139 262178
rect 3235 262144 3559 262178
rect 3655 262144 3979 262178
rect 4075 262144 4399 262178
rect 4495 262144 4819 262178
rect 4915 262144 5239 262178
rect 5335 262144 5659 262178
rect 5755 262144 6079 262178
rect 6175 262144 6499 262178
rect 6595 262144 6919 262178
rect 7015 262144 7339 262178
rect 7435 262144 7759 262178
rect 7855 262144 8179 262178
rect 8275 262144 8599 262178
rect 8695 262144 9019 262178
rect 9115 262144 9439 262178
rect 9535 262144 9859 262178
rect 9955 262144 10279 262178
rect 10375 262144 10699 262178
rect 10795 262144 11119 262178
rect 11215 262144 11539 262178
rect 11635 262144 11959 262178
rect 12055 262144 12379 262178
rect 12475 262144 12799 262178
rect 12895 262144 13219 262178
rect 13315 262144 13639 262178
rect 13735 262144 14059 262178
rect 14155 262144 14479 262178
rect 14575 262144 14899 262178
rect 14995 262144 15319 262178
rect 15415 262144 15739 262178
rect 15835 262144 16159 262178
rect 16255 262144 16579 262178
rect 16675 262144 16999 262178
rect 17095 262144 17419 262178
rect 17515 262144 17839 262178
rect 17935 262144 18259 262178
rect 18355 262144 18679 262178
rect 18775 262144 19099 262178
rect 19195 262144 19519 262178
rect 19615 262144 19939 262178
rect 20035 262144 20359 262178
rect 20455 262144 20779 262178
rect 20875 262144 21199 262178
rect 21295 262144 21619 262178
rect 21715 262144 22039 262178
rect 22135 262144 22459 262178
rect 22555 262144 22879 262178
rect 22975 262144 23299 262178
rect 23395 262144 23719 262178
rect 23815 262144 24139 262178
rect 24235 262144 24559 262178
rect 24655 262144 24979 262178
rect 25075 262144 25399 262178
rect 25495 262144 25819 262178
rect 25915 262144 26239 262178
rect 26335 262144 26659 262178
rect 26755 262144 27079 262178
rect 27175 262144 27285 262178
rect -5008 262138 27285 262144
rect -5008 254582 27285 254588
rect -5008 254548 -4001 254582
rect -3905 254548 -3581 254582
rect -3485 254548 -3161 254582
rect -3065 254548 -2741 254582
rect -2645 254548 -2321 254582
rect -2225 254548 -1901 254582
rect -1805 254548 -1481 254582
rect -1385 254548 -1061 254582
rect -965 254548 -641 254582
rect -545 254548 -221 254582
rect -125 254548 199 254582
rect 295 254548 619 254582
rect 715 254548 1039 254582
rect 1135 254548 1459 254582
rect 1555 254548 1879 254582
rect 1975 254548 2299 254582
rect 2395 254548 2719 254582
rect 2815 254548 3139 254582
rect 3235 254548 3559 254582
rect 3655 254548 3979 254582
rect 4075 254548 4399 254582
rect 4495 254548 4819 254582
rect 4915 254548 5239 254582
rect 5335 254548 5659 254582
rect 5755 254548 6079 254582
rect 6175 254548 6499 254582
rect 6595 254548 6919 254582
rect 7015 254548 7339 254582
rect 7435 254548 7759 254582
rect 7855 254548 8179 254582
rect 8275 254548 8599 254582
rect 8695 254548 9019 254582
rect 9115 254548 9439 254582
rect 9535 254548 9859 254582
rect 9955 254548 10279 254582
rect 10375 254548 10699 254582
rect 10795 254548 11119 254582
rect 11215 254548 11539 254582
rect 11635 254548 11959 254582
rect 12055 254548 12379 254582
rect 12475 254548 12799 254582
rect 12895 254548 13219 254582
rect 13315 254548 13639 254582
rect 13735 254548 14059 254582
rect 14155 254548 14479 254582
rect 14575 254548 14899 254582
rect 14995 254548 15319 254582
rect 15415 254548 15739 254582
rect 15835 254548 16159 254582
rect 16255 254548 16579 254582
rect 16675 254548 16999 254582
rect 17095 254548 17419 254582
rect 17515 254548 17839 254582
rect 17935 254548 18259 254582
rect 18355 254548 18679 254582
rect 18775 254548 19099 254582
rect 19195 254548 19519 254582
rect 19615 254548 19939 254582
rect 20035 254548 20359 254582
rect 20455 254548 20779 254582
rect 20875 254548 21199 254582
rect 21295 254548 21619 254582
rect 21715 254548 22039 254582
rect 22135 254548 22459 254582
rect 22555 254548 22879 254582
rect 22975 254548 23299 254582
rect 23395 254548 23719 254582
rect 23815 254548 24139 254582
rect 24235 254548 24559 254582
rect 24655 254548 24979 254582
rect 25075 254548 25399 254582
rect 25495 254548 25819 254582
rect 25915 254548 26239 254582
rect 26335 254548 26659 254582
rect 26755 254548 27079 254582
rect 27175 254548 27285 254582
rect -5008 254542 27285 254548
rect -5008 253654 -4142 254542
rect -4055 254489 -4009 254501
rect -3959 254489 -3913 254501
rect -3845 254489 -3799 254501
rect -3749 254489 -3703 254501
rect -3635 254489 -3589 254501
rect -3539 254490 -3493 254501
rect -3425 254490 -3379 254501
rect -3329 254490 -3283 254501
rect -3215 254490 -3169 254501
rect -3119 254490 -3073 254501
rect -3005 254490 -2959 254501
rect -2909 254490 -2863 254501
rect -2795 254490 -2749 254501
rect -2699 254490 -2653 254501
rect -2585 254490 -2539 254501
rect -2489 254490 -2443 254501
rect -2375 254490 -2329 254501
rect -2279 254490 -2233 254501
rect -2165 254490 -2119 254501
rect -2069 254490 -2023 254501
rect -1955 254490 -1909 254501
rect -1859 254490 -1813 254501
rect -1745 254490 -1699 254501
rect -1649 254490 -1603 254501
rect -1535 254490 -1489 254501
rect -1439 254490 -1393 254501
rect -1325 254490 -1279 254501
rect -1229 254490 -1183 254501
rect -1115 254490 -1069 254501
rect -1019 254490 -973 254501
rect -905 254490 -859 254501
rect -809 254490 -763 254501
rect -695 254490 -649 254501
rect -599 254490 -553 254501
rect -485 254490 -439 254501
rect -389 254490 -343 254501
rect -275 254490 -229 254501
rect -179 254490 -133 254501
rect -65 254490 -19 254501
rect 31 254490 77 254501
rect 145 254490 191 254501
rect 241 254490 287 254501
rect 355 254490 401 254501
rect 451 254490 497 254501
rect 565 254490 611 254501
rect 661 254490 707 254501
rect 775 254490 821 254501
rect 871 254490 917 254501
rect 985 254490 1031 254501
rect 1081 254490 1127 254501
rect 1195 254490 1241 254501
rect 1291 254490 1337 254501
rect 1405 254490 1451 254501
rect 1501 254490 1547 254501
rect 1615 254490 1661 254501
rect 1711 254490 1757 254501
rect 1825 254490 1871 254501
rect 1921 254490 1967 254501
rect 2035 254490 2081 254501
rect 2131 254490 2177 254501
rect 2245 254490 2291 254501
rect 2341 254490 2387 254501
rect 2455 254490 2501 254501
rect 2551 254490 2597 254501
rect 2665 254490 2711 254501
rect 2761 254490 2807 254501
rect 2875 254490 2921 254501
rect 2971 254490 3017 254501
rect 3085 254490 3131 254501
rect 3181 254490 3227 254501
rect 3295 254490 3341 254501
rect 3391 254490 3437 254501
rect 3505 254490 3551 254501
rect 3601 254490 3647 254501
rect 3715 254490 3761 254501
rect 3811 254490 3857 254501
rect 3925 254490 3971 254501
rect 4021 254490 4067 254501
rect 4135 254490 4181 254501
rect 4231 254490 4277 254501
rect 4345 254490 4391 254501
rect 4441 254490 4487 254501
rect 4555 254490 4601 254501
rect 4651 254490 4697 254501
rect 4765 254490 4811 254501
rect 4861 254490 4907 254501
rect 4975 254490 5021 254501
rect 5071 254490 5117 254501
rect 5185 254490 5231 254501
rect 5281 254490 5327 254501
rect 5395 254490 5441 254501
rect 5491 254490 5537 254501
rect 5605 254490 5651 254501
rect 5701 254490 5747 254501
rect 5815 254490 5861 254501
rect 5911 254490 5957 254501
rect 6025 254490 6071 254501
rect 6121 254490 6167 254501
rect 6235 254490 6281 254501
rect 6331 254490 6377 254501
rect 6445 254490 6491 254501
rect 6541 254490 6587 254501
rect 6655 254490 6701 254501
rect 6751 254490 6797 254501
rect 6865 254490 6911 254501
rect 6961 254490 7007 254501
rect 7075 254490 7121 254501
rect 7171 254490 7217 254501
rect 7285 254490 7331 254501
rect 7381 254490 7427 254501
rect 7495 254490 7541 254501
rect 7591 254490 7637 254501
rect 7705 254490 7751 254501
rect 7801 254490 7847 254501
rect 7915 254490 7961 254501
rect 8011 254490 8057 254501
rect 8125 254490 8171 254501
rect 8221 254490 8267 254501
rect 8335 254490 8381 254501
rect 8431 254490 8477 254501
rect 8545 254490 8591 254501
rect 8641 254490 8687 254501
rect 8755 254490 8801 254501
rect 8851 254490 8897 254501
rect 8965 254490 9011 254501
rect 9061 254490 9107 254501
rect 9175 254490 9221 254501
rect 9271 254490 9317 254501
rect 9385 254490 9431 254501
rect 9481 254490 9527 254501
rect 9595 254490 9641 254501
rect 9691 254490 9737 254501
rect 9805 254490 9851 254501
rect 9901 254490 9947 254501
rect 10015 254490 10061 254501
rect 10111 254490 10157 254501
rect 10225 254490 10271 254501
rect 10321 254490 10367 254501
rect 10435 254490 10481 254501
rect 10531 254490 10577 254501
rect 10645 254490 10691 254501
rect 10741 254490 10787 254501
rect 10855 254490 10901 254501
rect 10951 254490 10997 254501
rect 11065 254490 11111 254501
rect 11161 254490 11207 254501
rect 11275 254490 11321 254501
rect 11371 254490 11417 254501
rect 11485 254490 11531 254501
rect 11581 254490 11627 254501
rect 11695 254490 11741 254501
rect 11791 254490 11837 254501
rect 11905 254490 11951 254501
rect 12001 254490 12047 254501
rect 12115 254490 12161 254501
rect 12211 254490 12257 254501
rect 12325 254490 12371 254501
rect 12421 254490 12467 254501
rect 12535 254490 12581 254501
rect 12631 254490 12677 254501
rect 12745 254490 12791 254501
rect 12841 254490 12887 254501
rect 12955 254490 13001 254501
rect 13051 254490 13097 254501
rect 13165 254490 13211 254501
rect 13261 254490 13307 254501
rect 13375 254490 13421 254501
rect 13471 254490 13517 254501
rect 13585 254490 13631 254501
rect 13681 254490 13727 254501
rect 13795 254490 13841 254501
rect 13891 254490 13937 254501
rect 14005 254490 14051 254501
rect 14101 254490 14147 254501
rect 14215 254490 14261 254501
rect 14311 254490 14357 254501
rect 14425 254490 14471 254501
rect 14521 254490 14567 254501
rect 14635 254490 14681 254501
rect 14731 254490 14777 254501
rect 14845 254490 14891 254501
rect 14941 254490 14987 254501
rect 15055 254490 15101 254501
rect 15151 254490 15197 254501
rect 15265 254490 15311 254501
rect 15361 254490 15407 254501
rect 15475 254490 15521 254501
rect 15571 254490 15617 254501
rect 15685 254490 15731 254501
rect 15781 254490 15827 254501
rect 15895 254490 15941 254501
rect 15991 254490 16037 254501
rect 16105 254490 16151 254501
rect 16201 254490 16247 254501
rect 16315 254490 16361 254501
rect 16411 254490 16457 254501
rect 16525 254490 16571 254501
rect 16621 254490 16667 254501
rect 16735 254490 16781 254501
rect 16831 254490 16877 254501
rect 16945 254490 16991 254501
rect 17041 254490 17087 254501
rect 17155 254490 17201 254501
rect 17251 254490 17297 254501
rect 17365 254490 17411 254501
rect 17461 254490 17507 254501
rect 17575 254490 17621 254501
rect 17671 254490 17717 254501
rect 17785 254490 17831 254501
rect 17881 254490 17927 254501
rect 17995 254490 18041 254501
rect 18091 254490 18137 254501
rect 18205 254490 18251 254501
rect 18301 254490 18347 254501
rect 18415 254490 18461 254501
rect 18511 254490 18557 254501
rect 18625 254490 18671 254501
rect 18721 254490 18767 254501
rect 18835 254490 18881 254501
rect 18931 254490 18977 254501
rect 19045 254490 19091 254501
rect 19141 254490 19187 254501
rect 19255 254490 19301 254501
rect 19351 254490 19397 254501
rect 19465 254490 19511 254501
rect 19561 254490 19607 254501
rect 19675 254490 19721 254501
rect 19771 254490 19817 254501
rect 19885 254490 19931 254501
rect 19981 254490 20027 254501
rect 20095 254490 20141 254501
rect 20191 254490 20237 254501
rect 20305 254490 20351 254501
rect 20401 254490 20447 254501
rect 20515 254490 20561 254501
rect 20611 254490 20657 254501
rect 20725 254490 20771 254501
rect 20821 254490 20867 254501
rect 20935 254490 20981 254501
rect 21031 254490 21077 254501
rect 21145 254490 21191 254501
rect 21241 254490 21287 254501
rect 21355 254490 21401 254501
rect 21451 254490 21497 254501
rect 21565 254490 21611 254501
rect 21661 254490 21707 254501
rect 21775 254490 21821 254501
rect 21871 254490 21917 254501
rect 21985 254490 22031 254501
rect 22081 254490 22127 254501
rect 22195 254490 22241 254501
rect 22291 254490 22337 254501
rect 22405 254490 22451 254501
rect 22501 254490 22547 254501
rect 22615 254490 22661 254501
rect 22711 254490 22757 254501
rect 22825 254490 22871 254501
rect 22921 254490 22967 254501
rect 23035 254490 23081 254501
rect 23131 254490 23177 254501
rect 23245 254490 23291 254501
rect 23341 254490 23387 254501
rect 23455 254490 23501 254501
rect 23551 254490 23597 254501
rect 23665 254490 23711 254501
rect 23761 254490 23807 254501
rect 23875 254490 23921 254501
rect 23971 254490 24017 254501
rect 24085 254490 24131 254501
rect 24181 254490 24227 254501
rect 24295 254490 24341 254501
rect 24391 254490 24437 254501
rect 24505 254490 24551 254501
rect 24601 254490 24647 254501
rect 24715 254490 24761 254501
rect 24811 254490 24857 254501
rect 24925 254490 24971 254501
rect 25021 254490 25067 254501
rect 25135 254490 25181 254501
rect 25231 254490 25277 254501
rect 25345 254490 25391 254501
rect 25441 254490 25487 254501
rect 25555 254490 25601 254501
rect 25651 254490 25697 254501
rect 25765 254490 25811 254501
rect 25861 254490 25907 254501
rect 25975 254490 26021 254501
rect 26071 254490 26117 254501
rect 26185 254490 26231 254501
rect 26281 254490 26327 254501
rect 26395 254490 26441 254501
rect 26491 254490 26537 254501
rect 26605 254490 26651 254501
rect 26701 254490 26747 254501
rect 26815 254490 26861 254501
rect 26911 254490 26957 254501
rect 27025 254490 27071 254501
rect 27121 254490 27167 254501
rect 27235 254490 27281 254501
rect -4079 253713 -4069 254489
rect -4015 253713 -4005 254489
rect -3963 253713 -3953 254489
rect -3805 253713 -3795 254489
rect -3753 253713 -3743 254489
rect -3595 253713 -3585 254489
rect -3543 253713 -3533 254490
rect -3385 253713 -3375 254490
rect -3333 253713 -3323 254490
rect -3175 253713 -3165 254490
rect -3123 253713 -3113 254490
rect -2965 253713 -2955 254490
rect -2913 253713 -2903 254490
rect -2755 253713 -2745 254490
rect -2703 253713 -2693 254490
rect -2545 253713 -2535 254490
rect -2493 253713 -2483 254490
rect -2335 253713 -2325 254490
rect -2283 253713 -2273 254490
rect -2125 253713 -2115 254490
rect -2073 253713 -2063 254490
rect -1915 253713 -1905 254490
rect -1863 253713 -1853 254490
rect -1705 253713 -1695 254490
rect -1653 253713 -1643 254490
rect -1495 253713 -1485 254490
rect -1443 253713 -1433 254490
rect -1285 253713 -1275 254490
rect -1233 253713 -1223 254490
rect -1075 253713 -1065 254490
rect -1023 253713 -1013 254490
rect -865 253713 -855 254490
rect -813 253713 -803 254490
rect -655 253713 -645 254490
rect -603 253713 -593 254490
rect -445 253713 -435 254490
rect -393 253713 -383 254490
rect -235 253713 -225 254490
rect -183 253713 -173 254490
rect -25 253713 -15 254490
rect 27 253713 37 254490
rect 185 253713 195 254490
rect 237 253713 247 254490
rect 395 253713 405 254490
rect 447 253713 457 254490
rect 605 253713 615 254490
rect 657 253713 667 254490
rect 815 253713 825 254490
rect 867 253713 877 254490
rect 1025 253713 1035 254490
rect 1077 253713 1087 254490
rect 1235 253713 1245 254490
rect 1287 253713 1297 254490
rect 1445 253713 1455 254490
rect 1497 253713 1507 254490
rect 1655 253713 1665 254490
rect 1707 253713 1717 254490
rect 1865 253713 1875 254490
rect 1917 253713 1927 254490
rect 2075 253713 2085 254490
rect 2127 253713 2137 254490
rect 2285 253713 2295 254490
rect 2337 253713 2347 254490
rect 2495 253713 2505 254490
rect 2547 253713 2557 254490
rect 2705 253713 2715 254490
rect 2757 253713 2767 254490
rect 2915 253713 2925 254490
rect 2967 253713 2977 254490
rect 3125 253713 3135 254490
rect 3177 253713 3187 254490
rect 3335 253713 3345 254490
rect 3387 253713 3397 254490
rect 3545 253713 3555 254490
rect 3597 253713 3607 254490
rect 3755 253713 3765 254490
rect 3807 253713 3817 254490
rect 3965 253713 3975 254490
rect 4017 253713 4027 254490
rect 4175 253713 4185 254490
rect 4227 253713 4237 254490
rect 4385 253713 4395 254490
rect 4437 253713 4447 254490
rect 4595 253713 4605 254490
rect 4647 253713 4657 254490
rect 4805 253713 4815 254490
rect 4857 253713 4867 254490
rect 5015 253713 5025 254490
rect 5067 253713 5077 254490
rect 5225 253713 5235 254490
rect 5277 253713 5287 254490
rect 5435 253713 5445 254490
rect 5487 253713 5497 254490
rect 5645 253713 5655 254490
rect 5697 253713 5707 254490
rect 5855 253713 5865 254490
rect 5907 253713 5917 254490
rect 6065 253713 6075 254490
rect 6117 253713 6127 254490
rect 6275 253713 6285 254490
rect 6327 253713 6337 254490
rect 6485 253713 6495 254490
rect 6537 253713 6547 254490
rect 6695 253713 6705 254490
rect 6747 253713 6757 254490
rect 6905 253713 6915 254490
rect 6957 253713 6967 254490
rect 7115 253713 7125 254490
rect 7167 253713 7177 254490
rect 7325 253713 7335 254490
rect 7377 253713 7387 254490
rect 7535 253713 7545 254490
rect 7587 253713 7597 254490
rect 7745 253713 7755 254490
rect 7797 253713 7807 254490
rect 7955 253713 7965 254490
rect 8007 253713 8017 254490
rect 8165 253713 8175 254490
rect 8217 253713 8227 254490
rect 8375 253713 8385 254490
rect 8427 253713 8437 254490
rect 8585 253713 8595 254490
rect 8637 253713 8647 254490
rect 8795 253713 8805 254490
rect 8847 253713 8857 254490
rect 9005 253713 9015 254490
rect 9057 253713 9067 254490
rect 9215 253713 9225 254490
rect 9267 253713 9277 254490
rect 9425 253713 9435 254490
rect 9477 253713 9487 254490
rect 9635 253713 9645 254490
rect 9687 253713 9697 254490
rect 9845 253713 9855 254490
rect 9897 253713 9907 254490
rect 10055 253713 10065 254490
rect 10107 253713 10117 254490
rect 10265 253713 10275 254490
rect 10317 253713 10327 254490
rect 10475 253713 10485 254490
rect 10527 253713 10537 254490
rect 10685 253713 10695 254490
rect 10737 253713 10747 254490
rect 10895 253713 10905 254490
rect 10947 253713 10957 254490
rect 11105 253713 11115 254490
rect 11157 253713 11167 254490
rect 11315 253713 11325 254490
rect 11367 253713 11377 254490
rect 11525 253713 11535 254490
rect 11577 253713 11587 254490
rect 11735 253713 11745 254490
rect 11787 253713 11797 254490
rect 11945 253713 11955 254490
rect 11997 253713 12007 254490
rect 12155 253713 12165 254490
rect 12207 253713 12217 254490
rect 12365 253713 12375 254490
rect 12417 253713 12427 254490
rect 12575 253713 12585 254490
rect 12627 253713 12637 254490
rect 12785 253713 12795 254490
rect 12837 253713 12847 254490
rect 12995 253713 13005 254490
rect 13047 253713 13057 254490
rect 13205 253713 13215 254490
rect 13257 253713 13267 254490
rect 13415 253713 13425 254490
rect 13467 253713 13477 254490
rect 13625 253713 13635 254490
rect 13677 253713 13687 254490
rect 13835 253713 13845 254490
rect 13887 253713 13897 254490
rect 14045 253713 14055 254490
rect 14097 253713 14107 254490
rect 14255 253713 14265 254490
rect 14307 253713 14317 254490
rect 14465 253713 14475 254490
rect 14517 253713 14527 254490
rect 14675 253713 14685 254490
rect 14727 253713 14737 254490
rect 14885 253713 14895 254490
rect 14937 253713 14947 254490
rect 15095 253713 15105 254490
rect 15147 253713 15157 254490
rect 15305 253713 15315 254490
rect 15357 253713 15367 254490
rect 15515 253713 15525 254490
rect 15567 253713 15577 254490
rect 15725 253713 15735 254490
rect 15777 253713 15787 254490
rect 15935 253713 15945 254490
rect 15987 253713 15997 254490
rect 16145 253713 16155 254490
rect 16197 253713 16207 254490
rect 16355 253713 16365 254490
rect 16407 253713 16417 254490
rect 16565 253713 16575 254490
rect 16617 253713 16627 254490
rect 16775 253713 16785 254490
rect 16827 253713 16837 254490
rect 16985 253713 16995 254490
rect 17037 253713 17047 254490
rect 17195 253713 17205 254490
rect 17247 253713 17257 254490
rect 17405 253713 17415 254490
rect 17457 253713 17467 254490
rect 17615 253713 17625 254490
rect 17667 253713 17677 254490
rect 17825 253713 17835 254490
rect 17877 253713 17887 254490
rect 18035 253713 18045 254490
rect 18087 253713 18097 254490
rect 18245 253713 18255 254490
rect 18297 253713 18307 254490
rect 18455 253713 18465 254490
rect 18507 253713 18517 254490
rect 18665 253713 18675 254490
rect 18717 253713 18727 254490
rect 18875 253713 18885 254490
rect 18927 253713 18937 254490
rect 19085 253713 19095 254490
rect 19137 253713 19147 254490
rect 19295 253713 19305 254490
rect 19347 253713 19357 254490
rect 19505 253713 19515 254490
rect 19557 253713 19567 254490
rect 19715 253713 19725 254490
rect 19767 253713 19777 254490
rect 19925 253713 19935 254490
rect 19977 253713 19987 254490
rect 20135 253713 20145 254490
rect 20187 253713 20197 254490
rect 20345 253713 20355 254490
rect 20397 253713 20407 254490
rect 20555 253713 20565 254490
rect 20607 253713 20617 254490
rect 20765 253713 20775 254490
rect 20817 253713 20827 254490
rect 20975 253713 20985 254490
rect 21027 253713 21037 254490
rect 21185 253713 21195 254490
rect 21237 253713 21247 254490
rect 21395 253713 21405 254490
rect 21447 253713 21457 254490
rect 21605 253713 21615 254490
rect 21657 253713 21667 254490
rect 21815 253713 21825 254490
rect 21867 253713 21877 254490
rect 22025 253713 22035 254490
rect 22077 253713 22087 254490
rect 22235 253713 22245 254490
rect 22287 253713 22297 254490
rect 22445 253713 22455 254490
rect 22497 253713 22507 254490
rect 22655 253713 22665 254490
rect 22707 253713 22717 254490
rect 22865 253713 22875 254490
rect 22917 253713 22927 254490
rect 23075 253713 23085 254490
rect 23127 253713 23137 254490
rect 23285 253713 23295 254490
rect 23337 253713 23347 254490
rect 23495 253713 23505 254490
rect 23547 253713 23557 254490
rect 23705 253713 23715 254490
rect 23757 253713 23767 254490
rect 23915 253713 23925 254490
rect 23967 253713 23977 254490
rect 24125 253713 24135 254490
rect 24177 253713 24187 254490
rect 24335 253713 24345 254490
rect 24387 253713 24397 254490
rect 24545 253713 24555 254490
rect 24597 253713 24607 254490
rect 24755 253713 24765 254490
rect 24807 253713 24817 254490
rect 24965 253713 24975 254490
rect 25017 253713 25027 254490
rect 25175 253713 25185 254490
rect 25227 253713 25237 254490
rect 25385 253713 25395 254490
rect 25437 253713 25447 254490
rect 25595 253713 25605 254490
rect 25647 253713 25657 254490
rect 25805 253713 25815 254490
rect 25857 253713 25867 254490
rect 26015 253713 26025 254490
rect 26067 253713 26077 254490
rect 26225 253713 26235 254490
rect 26277 253713 26287 254490
rect 26435 253713 26445 254490
rect 26487 253713 26497 254490
rect 26645 253713 26655 254490
rect 26697 253713 26707 254490
rect 26855 253713 26865 254490
rect 26907 253713 26917 254490
rect 27065 253713 27075 254490
rect 27117 253713 27127 254490
rect 27275 253713 27285 254490
rect 27331 254489 27566 254501
rect 27331 253713 27337 254489
rect 27371 253713 27566 254489
rect -4055 253701 -4009 253713
rect -3959 253701 -3913 253713
rect -3845 253701 -3799 253713
rect -3749 253701 -3703 253713
rect -3635 253701 -3589 253713
rect -3539 253701 -3493 253713
rect -3425 253701 -3379 253713
rect -3329 253701 -3283 253713
rect -3215 253701 -3169 253713
rect -3119 253701 -3073 253713
rect -3005 253701 -2959 253713
rect -2909 253701 -2863 253713
rect -2795 253701 -2749 253713
rect -2699 253701 -2653 253713
rect -2585 253701 -2539 253713
rect -2489 253701 -2443 253713
rect -2375 253701 -2329 253713
rect -2279 253701 -2233 253713
rect -2165 253701 -2119 253713
rect -2069 253701 -2023 253713
rect -1955 253701 -1909 253713
rect -1859 253701 -1813 253713
rect -1745 253701 -1699 253713
rect -1649 253701 -1603 253713
rect -1535 253701 -1489 253713
rect -1439 253701 -1393 253713
rect -1325 253701 -1279 253713
rect -1229 253701 -1183 253713
rect -1115 253701 -1069 253713
rect -1019 253701 -973 253713
rect -905 253701 -859 253713
rect -809 253701 -763 253713
rect -695 253701 -649 253713
rect -599 253701 -553 253713
rect -485 253701 -439 253713
rect -389 253701 -343 253713
rect -275 253701 -229 253713
rect -179 253701 -133 253713
rect -65 253701 -19 253713
rect 31 253701 77 253713
rect 145 253701 191 253713
rect 241 253701 287 253713
rect 355 253701 401 253713
rect 451 253701 497 253713
rect 565 253701 611 253713
rect 661 253701 707 253713
rect 775 253701 821 253713
rect 871 253701 917 253713
rect 985 253701 1031 253713
rect 1081 253701 1127 253713
rect 1195 253701 1241 253713
rect 1291 253701 1337 253713
rect 1405 253701 1451 253713
rect 1501 253701 1547 253713
rect 1615 253701 1661 253713
rect 1711 253701 1757 253713
rect 1825 253701 1871 253713
rect 1921 253701 1967 253713
rect 2035 253701 2081 253713
rect 2131 253701 2177 253713
rect 2245 253701 2291 253713
rect 2341 253701 2387 253713
rect 2455 253701 2501 253713
rect 2551 253701 2597 253713
rect 2665 253701 2711 253713
rect 2761 253701 2807 253713
rect 2875 253701 2921 253713
rect 2971 253701 3017 253713
rect 3085 253701 3131 253713
rect 3181 253701 3227 253713
rect 3295 253701 3341 253713
rect 3391 253701 3437 253713
rect 3505 253701 3551 253713
rect 3601 253701 3647 253713
rect 3715 253701 3761 253713
rect 3811 253701 3857 253713
rect 3925 253701 3971 253713
rect 4021 253701 4067 253713
rect 4135 253701 4181 253713
rect 4231 253701 4277 253713
rect 4345 253701 4391 253713
rect 4441 253701 4487 253713
rect 4555 253701 4601 253713
rect 4651 253701 4697 253713
rect 4765 253701 4811 253713
rect 4861 253701 4907 253713
rect 4975 253701 5021 253713
rect 5071 253701 5117 253713
rect 5185 253701 5231 253713
rect 5281 253701 5327 253713
rect 5395 253701 5441 253713
rect 5491 253701 5537 253713
rect 5605 253701 5651 253713
rect 5701 253701 5747 253713
rect 5815 253701 5861 253713
rect 5911 253701 5957 253713
rect 6025 253701 6071 253713
rect 6121 253701 6167 253713
rect 6235 253701 6281 253713
rect 6331 253701 6377 253713
rect 6445 253701 6491 253713
rect 6541 253701 6587 253713
rect 6655 253701 6701 253713
rect 6751 253701 6797 253713
rect 6865 253701 6911 253713
rect 6961 253701 7007 253713
rect 7075 253701 7121 253713
rect 7171 253701 7217 253713
rect 7285 253701 7331 253713
rect 7381 253701 7427 253713
rect 7495 253701 7541 253713
rect 7591 253701 7637 253713
rect 7705 253701 7751 253713
rect 7801 253701 7847 253713
rect 7915 253701 7961 253713
rect 8011 253701 8057 253713
rect 8125 253701 8171 253713
rect 8221 253701 8267 253713
rect 8335 253701 8381 253713
rect 8431 253701 8477 253713
rect 8545 253701 8591 253713
rect 8641 253701 8687 253713
rect 8755 253701 8801 253713
rect 8851 253701 8897 253713
rect 8965 253701 9011 253713
rect 9061 253701 9107 253713
rect 9175 253701 9221 253713
rect 9271 253701 9317 253713
rect 9385 253701 9431 253713
rect 9481 253701 9527 253713
rect 9595 253701 9641 253713
rect 9691 253701 9737 253713
rect 9805 253701 9851 253713
rect 9901 253701 9947 253713
rect 10015 253701 10061 253713
rect 10111 253701 10157 253713
rect 10225 253701 10271 253713
rect 10321 253701 10367 253713
rect 10435 253701 10481 253713
rect 10531 253701 10577 253713
rect 10645 253701 10691 253713
rect 10741 253701 10787 253713
rect 10855 253701 10901 253713
rect 10951 253701 10997 253713
rect 11065 253701 11111 253713
rect 11161 253701 11207 253713
rect 11275 253701 11321 253713
rect 11371 253701 11417 253713
rect 11485 253701 11531 253713
rect 11581 253701 11627 253713
rect 11695 253701 11741 253713
rect 11791 253701 11837 253713
rect 11905 253701 11951 253713
rect 12001 253701 12047 253713
rect 12115 253701 12161 253713
rect 12211 253701 12257 253713
rect 12325 253701 12371 253713
rect 12421 253701 12467 253713
rect 12535 253701 12581 253713
rect 12631 253701 12677 253713
rect 12745 253701 12791 253713
rect 12841 253701 12887 253713
rect 12955 253701 13001 253713
rect 13051 253701 13097 253713
rect 13165 253701 13211 253713
rect 13261 253701 13307 253713
rect 13375 253701 13421 253713
rect 13471 253701 13517 253713
rect 13585 253701 13631 253713
rect 13681 253701 13727 253713
rect 13795 253701 13841 253713
rect 13891 253701 13937 253713
rect 14005 253701 14051 253713
rect 14101 253701 14147 253713
rect 14215 253701 14261 253713
rect 14311 253701 14357 253713
rect 14425 253701 14471 253713
rect 14521 253701 14567 253713
rect 14635 253701 14681 253713
rect 14731 253701 14777 253713
rect 14845 253701 14891 253713
rect 14941 253701 14987 253713
rect 15055 253701 15101 253713
rect 15151 253701 15197 253713
rect 15265 253701 15311 253713
rect 15361 253701 15407 253713
rect 15475 253701 15521 253713
rect 15571 253701 15617 253713
rect 15685 253701 15731 253713
rect 15781 253701 15827 253713
rect 15895 253701 15941 253713
rect 15991 253701 16037 253713
rect 16105 253701 16151 253713
rect 16201 253701 16247 253713
rect 16315 253701 16361 253713
rect 16411 253701 16457 253713
rect 16525 253701 16571 253713
rect 16621 253701 16667 253713
rect 16735 253701 16781 253713
rect 16831 253701 16877 253713
rect 16945 253701 16991 253713
rect 17041 253701 17087 253713
rect 17155 253701 17201 253713
rect 17251 253701 17297 253713
rect 17365 253701 17411 253713
rect 17461 253701 17507 253713
rect 17575 253701 17621 253713
rect 17671 253701 17717 253713
rect 17785 253701 17831 253713
rect 17881 253701 17927 253713
rect 17995 253701 18041 253713
rect 18091 253701 18137 253713
rect 18205 253701 18251 253713
rect 18301 253701 18347 253713
rect 18415 253701 18461 253713
rect 18511 253701 18557 253713
rect 18625 253701 18671 253713
rect 18721 253701 18767 253713
rect 18835 253701 18881 253713
rect 18931 253701 18977 253713
rect 19045 253701 19091 253713
rect 19141 253701 19187 253713
rect 19255 253701 19301 253713
rect 19351 253701 19397 253713
rect 19465 253701 19511 253713
rect 19561 253701 19607 253713
rect 19675 253701 19721 253713
rect 19771 253701 19817 253713
rect 19885 253701 19931 253713
rect 19981 253701 20027 253713
rect 20095 253701 20141 253713
rect 20191 253701 20237 253713
rect 20305 253701 20351 253713
rect 20401 253701 20447 253713
rect 20515 253701 20561 253713
rect 20611 253701 20657 253713
rect 20725 253701 20771 253713
rect 20821 253701 20867 253713
rect 20935 253701 20981 253713
rect 21031 253701 21077 253713
rect 21145 253701 21191 253713
rect 21241 253701 21287 253713
rect 21355 253701 21401 253713
rect 21451 253701 21497 253713
rect 21565 253701 21611 253713
rect 21661 253701 21707 253713
rect 21775 253701 21821 253713
rect 21871 253701 21917 253713
rect 21985 253701 22031 253713
rect 22081 253701 22127 253713
rect 22195 253701 22241 253713
rect 22291 253701 22337 253713
rect 22405 253701 22451 253713
rect 22501 253701 22547 253713
rect 22615 253701 22661 253713
rect 22711 253701 22757 253713
rect 22825 253701 22871 253713
rect 22921 253701 22967 253713
rect 23035 253701 23081 253713
rect 23131 253701 23177 253713
rect 23245 253701 23291 253713
rect 23341 253701 23387 253713
rect 23455 253701 23501 253713
rect 23551 253701 23597 253713
rect 23665 253701 23711 253713
rect 23761 253701 23807 253713
rect 23875 253701 23921 253713
rect 23971 253701 24017 253713
rect 24085 253701 24131 253713
rect 24181 253701 24227 253713
rect 24295 253701 24341 253713
rect 24391 253701 24437 253713
rect 24505 253701 24551 253713
rect 24601 253701 24647 253713
rect 24715 253701 24761 253713
rect 24811 253701 24857 253713
rect 24925 253701 24971 253713
rect 25021 253701 25067 253713
rect 25135 253701 25181 253713
rect 25231 253701 25277 253713
rect 25345 253701 25391 253713
rect 25441 253701 25487 253713
rect 25555 253701 25601 253713
rect 25651 253701 25697 253713
rect 25765 253701 25811 253713
rect 25861 253701 25907 253713
rect 25975 253701 26021 253713
rect 26071 253701 26117 253713
rect 26185 253701 26231 253713
rect 26281 253701 26327 253713
rect 26395 253701 26441 253713
rect 26491 253701 26537 253713
rect 26605 253701 26651 253713
rect 26701 253701 26747 253713
rect 26815 253701 26861 253713
rect 26911 253701 26957 253713
rect 27025 253701 27071 253713
rect 27121 253701 27167 253713
rect 27235 253701 27281 253713
rect 27331 253701 27566 253713
rect -3803 253654 27335 253666
rect -5008 253512 -3791 253654
rect -3757 253512 -3371 253654
rect -3337 253512 -2951 253654
rect -2917 253512 -2531 253654
rect -2497 253512 -2111 253654
rect -2077 253512 -1691 253654
rect -1657 253512 -1271 253654
rect -1237 253512 -851 253654
rect -817 253512 -431 253654
rect -397 253512 -11 253654
rect 23 253512 409 253654
rect 443 253512 829 253654
rect 863 253512 1249 253654
rect 1283 253512 1669 253654
rect 1703 253512 2089 253654
rect 2123 253512 2509 253654
rect 2543 253512 2929 253654
rect 2963 253512 3349 253654
rect 3383 253512 3769 253654
rect 3803 253512 4189 253654
rect 4223 253512 4609 253654
rect 4643 253512 5029 253654
rect 5063 253512 5449 253654
rect 5483 253512 5869 253654
rect 5903 253512 6289 253654
rect 6323 253512 6709 253654
rect 6743 253512 7129 253654
rect 7163 253512 7549 253654
rect 7583 253512 7969 253654
rect 8003 253512 8389 253654
rect 8423 253512 8809 253654
rect 8843 253512 9229 253654
rect 9263 253512 9649 253654
rect 9683 253512 10069 253654
rect 10103 253512 10489 253654
rect 10523 253512 10909 253654
rect 10943 253512 11329 253654
rect 11363 253512 11749 253654
rect 11783 253512 12169 253654
rect 12203 253512 12589 253654
rect 12623 253512 13009 253654
rect 13043 253512 13429 253654
rect 13463 253512 13849 253654
rect 13883 253512 14269 253654
rect 14303 253512 14689 253654
rect 14723 253512 15109 253654
rect 15143 253512 15529 253654
rect 15563 253512 15949 253654
rect 15983 253512 16369 253654
rect 16403 253512 16789 253654
rect 16823 253512 17209 253654
rect 17243 253512 17629 253654
rect 17663 253512 18049 253654
rect 18083 253512 18469 253654
rect 18503 253512 18889 253654
rect 18923 253512 19309 253654
rect 19343 253512 19729 253654
rect 19763 253512 20149 253654
rect 20183 253512 20569 253654
rect 20603 253512 20989 253654
rect 21023 253512 21409 253654
rect 21443 253512 21829 253654
rect 21863 253512 22249 253654
rect 22283 253512 22669 253654
rect 22703 253512 23089 253654
rect 23123 253512 23509 253654
rect 23543 253512 23929 253654
rect 23963 253512 24349 253654
rect 24383 253512 24769 253654
rect 24803 253512 25189 253654
rect 25223 253512 25609 253654
rect 25643 253512 26029 253654
rect 26063 253512 26449 253654
rect 26483 253512 26869 253654
rect 26903 253512 27289 253654
rect 27323 253512 27335 253654
rect -5008 252618 -4142 253512
rect -3803 253500 27335 253512
rect 27377 253465 27566 253701
rect -4055 253453 -4009 253465
rect -3959 253453 -3913 253465
rect -3845 253453 -3799 253465
rect -3749 253453 -3703 253465
rect -3635 253453 -3589 253465
rect -3539 253454 -3493 253465
rect -3425 253454 -3379 253465
rect -3329 253454 -3283 253465
rect -3215 253454 -3169 253465
rect -3119 253454 -3073 253465
rect -3005 253454 -2959 253465
rect -2909 253454 -2863 253465
rect -2795 253454 -2749 253465
rect -2699 253454 -2653 253465
rect -2585 253454 -2539 253465
rect -2489 253454 -2443 253465
rect -2375 253454 -2329 253465
rect -2279 253454 -2233 253465
rect -2165 253454 -2119 253465
rect -2069 253454 -2023 253465
rect -1955 253454 -1909 253465
rect -1859 253454 -1813 253465
rect -1745 253454 -1699 253465
rect -1649 253454 -1603 253465
rect -1535 253454 -1489 253465
rect -1439 253454 -1393 253465
rect -1325 253454 -1279 253465
rect -1229 253454 -1183 253465
rect -1115 253454 -1069 253465
rect -1019 253454 -973 253465
rect -905 253454 -859 253465
rect -809 253454 -763 253465
rect -695 253454 -649 253465
rect -599 253454 -553 253465
rect -485 253454 -439 253465
rect -389 253454 -343 253465
rect -275 253454 -229 253465
rect -179 253454 -133 253465
rect -65 253454 -19 253465
rect 31 253454 77 253465
rect 145 253454 191 253465
rect 241 253454 287 253465
rect 355 253454 401 253465
rect 451 253454 497 253465
rect 565 253454 611 253465
rect 661 253454 707 253465
rect 775 253454 821 253465
rect 871 253454 917 253465
rect 985 253454 1031 253465
rect 1081 253454 1127 253465
rect 1195 253454 1241 253465
rect 1291 253454 1337 253465
rect 1405 253454 1451 253465
rect 1501 253454 1547 253465
rect 1615 253454 1661 253465
rect 1711 253454 1757 253465
rect 1825 253454 1871 253465
rect 1921 253454 1967 253465
rect 2035 253454 2081 253465
rect 2131 253454 2177 253465
rect 2245 253454 2291 253465
rect 2341 253454 2387 253465
rect 2455 253454 2501 253465
rect 2551 253454 2597 253465
rect 2665 253454 2711 253465
rect 2761 253454 2807 253465
rect 2875 253454 2921 253465
rect 2971 253454 3017 253465
rect 3085 253454 3131 253465
rect 3181 253454 3227 253465
rect 3295 253454 3341 253465
rect 3391 253454 3437 253465
rect 3505 253454 3551 253465
rect 3601 253454 3647 253465
rect 3715 253454 3761 253465
rect 3811 253454 3857 253465
rect 3925 253454 3971 253465
rect 4021 253454 4067 253465
rect 4135 253454 4181 253465
rect 4231 253454 4277 253465
rect 4345 253454 4391 253465
rect 4441 253454 4487 253465
rect 4555 253454 4601 253465
rect 4651 253454 4697 253465
rect 4765 253454 4811 253465
rect 4861 253454 4907 253465
rect 4975 253454 5021 253465
rect 5071 253454 5117 253465
rect 5185 253454 5231 253465
rect 5281 253454 5327 253465
rect 5395 253454 5441 253465
rect 5491 253454 5537 253465
rect 5605 253454 5651 253465
rect 5701 253454 5747 253465
rect 5815 253454 5861 253465
rect 5911 253454 5957 253465
rect 6025 253454 6071 253465
rect 6121 253454 6167 253465
rect 6235 253454 6281 253465
rect 6331 253454 6377 253465
rect 6445 253454 6491 253465
rect 6541 253454 6587 253465
rect 6655 253454 6701 253465
rect 6751 253454 6797 253465
rect 6865 253454 6911 253465
rect 6961 253454 7007 253465
rect 7075 253454 7121 253465
rect 7171 253454 7217 253465
rect 7285 253454 7331 253465
rect 7381 253454 7427 253465
rect 7495 253454 7541 253465
rect 7591 253454 7637 253465
rect 7705 253454 7751 253465
rect 7801 253454 7847 253465
rect 7915 253454 7961 253465
rect 8011 253454 8057 253465
rect 8125 253454 8171 253465
rect 8221 253454 8267 253465
rect 8335 253454 8381 253465
rect 8431 253454 8477 253465
rect 8545 253454 8591 253465
rect 8641 253454 8687 253465
rect 8755 253454 8801 253465
rect 8851 253454 8897 253465
rect 8965 253454 9011 253465
rect 9061 253454 9107 253465
rect 9175 253454 9221 253465
rect 9271 253454 9317 253465
rect 9385 253454 9431 253465
rect 9481 253454 9527 253465
rect 9595 253454 9641 253465
rect 9691 253454 9737 253465
rect 9805 253454 9851 253465
rect 9901 253454 9947 253465
rect 10015 253454 10061 253465
rect 10111 253454 10157 253465
rect 10225 253454 10271 253465
rect 10321 253454 10367 253465
rect 10435 253454 10481 253465
rect 10531 253454 10577 253465
rect 10645 253454 10691 253465
rect 10741 253454 10787 253465
rect 10855 253454 10901 253465
rect 10951 253454 10997 253465
rect 11065 253454 11111 253465
rect 11161 253454 11207 253465
rect 11275 253454 11321 253465
rect 11371 253454 11417 253465
rect 11485 253454 11531 253465
rect 11581 253454 11627 253465
rect 11695 253454 11741 253465
rect 11791 253454 11837 253465
rect 11905 253454 11951 253465
rect 12001 253454 12047 253465
rect 12115 253454 12161 253465
rect 12211 253454 12257 253465
rect 12325 253454 12371 253465
rect 12421 253454 12467 253465
rect 12535 253454 12581 253465
rect 12631 253454 12677 253465
rect 12745 253454 12791 253465
rect 12841 253454 12887 253465
rect 12955 253454 13001 253465
rect 13051 253454 13097 253465
rect 13165 253454 13211 253465
rect 13261 253454 13307 253465
rect 13375 253454 13421 253465
rect 13471 253454 13517 253465
rect 13585 253454 13631 253465
rect 13681 253454 13727 253465
rect 13795 253454 13841 253465
rect 13891 253454 13937 253465
rect 14005 253454 14051 253465
rect 14101 253454 14147 253465
rect 14215 253454 14261 253465
rect 14311 253454 14357 253465
rect 14425 253454 14471 253465
rect 14521 253454 14567 253465
rect 14635 253454 14681 253465
rect 14731 253454 14777 253465
rect 14845 253454 14891 253465
rect 14941 253454 14987 253465
rect 15055 253454 15101 253465
rect 15151 253454 15197 253465
rect 15265 253454 15311 253465
rect 15361 253454 15407 253465
rect 15475 253454 15521 253465
rect 15571 253454 15617 253465
rect 15685 253454 15731 253465
rect 15781 253454 15827 253465
rect 15895 253454 15941 253465
rect 15991 253454 16037 253465
rect 16105 253454 16151 253465
rect 16201 253454 16247 253465
rect 16315 253454 16361 253465
rect 16411 253454 16457 253465
rect 16525 253454 16571 253465
rect 16621 253454 16667 253465
rect 16735 253454 16781 253465
rect 16831 253454 16877 253465
rect 16945 253454 16991 253465
rect 17041 253454 17087 253465
rect 17155 253454 17201 253465
rect 17251 253454 17297 253465
rect 17365 253454 17411 253465
rect 17461 253454 17507 253465
rect 17575 253454 17621 253465
rect 17671 253454 17717 253465
rect 17785 253454 17831 253465
rect 17881 253454 17927 253465
rect 17995 253454 18041 253465
rect 18091 253454 18137 253465
rect 18205 253454 18251 253465
rect 18301 253454 18347 253465
rect 18415 253454 18461 253465
rect 18511 253454 18557 253465
rect 18625 253454 18671 253465
rect 18721 253454 18767 253465
rect 18835 253454 18881 253465
rect 18931 253454 18977 253465
rect 19045 253454 19091 253465
rect 19141 253454 19187 253465
rect 19255 253454 19301 253465
rect 19351 253454 19397 253465
rect 19465 253454 19511 253465
rect 19561 253454 19607 253465
rect 19675 253454 19721 253465
rect 19771 253454 19817 253465
rect 19885 253454 19931 253465
rect 19981 253454 20027 253465
rect 20095 253454 20141 253465
rect 20191 253454 20237 253465
rect 20305 253454 20351 253465
rect 20401 253454 20447 253465
rect 20515 253454 20561 253465
rect 20611 253454 20657 253465
rect 20725 253454 20771 253465
rect 20821 253454 20867 253465
rect 20935 253454 20981 253465
rect 21031 253454 21077 253465
rect 21145 253454 21191 253465
rect 21241 253454 21287 253465
rect 21355 253454 21401 253465
rect 21451 253454 21497 253465
rect 21565 253454 21611 253465
rect 21661 253454 21707 253465
rect 21775 253454 21821 253465
rect 21871 253454 21917 253465
rect 21985 253454 22031 253465
rect 22081 253454 22127 253465
rect 22195 253454 22241 253465
rect 22291 253454 22337 253465
rect 22405 253454 22451 253465
rect 22501 253454 22547 253465
rect 22615 253454 22661 253465
rect 22711 253454 22757 253465
rect 22825 253454 22871 253465
rect 22921 253454 22967 253465
rect 23035 253454 23081 253465
rect 23131 253454 23177 253465
rect 23245 253454 23291 253465
rect 23341 253454 23387 253465
rect 23455 253454 23501 253465
rect 23551 253454 23597 253465
rect 23665 253454 23711 253465
rect 23761 253454 23807 253465
rect 23875 253454 23921 253465
rect 23971 253454 24017 253465
rect 24085 253454 24131 253465
rect 24181 253454 24227 253465
rect 24295 253454 24341 253465
rect 24391 253454 24437 253465
rect 24505 253454 24551 253465
rect 24601 253454 24647 253465
rect 24715 253454 24761 253465
rect 24811 253454 24857 253465
rect 24925 253454 24971 253465
rect 25021 253454 25067 253465
rect 25135 253454 25181 253465
rect 25231 253454 25277 253465
rect 25345 253454 25391 253465
rect 25441 253454 25487 253465
rect 25555 253454 25601 253465
rect 25651 253454 25697 253465
rect 25765 253454 25811 253465
rect 25861 253454 25907 253465
rect 25975 253454 26021 253465
rect 26071 253454 26117 253465
rect 26185 253454 26231 253465
rect 26281 253454 26327 253465
rect 26395 253454 26441 253465
rect 26491 253454 26537 253465
rect 26605 253454 26651 253465
rect 26701 253454 26747 253465
rect 26815 253454 26861 253465
rect 26911 253454 26957 253465
rect 27025 253454 27071 253465
rect 27121 253454 27167 253465
rect 27235 253454 27281 253465
rect -4079 252677 -4069 253453
rect -4015 252677 -4005 253453
rect -3963 252677 -3953 253453
rect -3805 252677 -3795 253453
rect -3753 252677 -3743 253453
rect -3595 252677 -3585 253453
rect -3543 252677 -3533 253454
rect -3385 252677 -3375 253454
rect -3333 252677 -3323 253454
rect -3175 252677 -3165 253454
rect -3123 252677 -3113 253454
rect -2965 252677 -2955 253454
rect -2913 252677 -2903 253454
rect -2755 252677 -2745 253454
rect -2703 252677 -2693 253454
rect -2545 252677 -2535 253454
rect -2493 252677 -2483 253454
rect -2335 252677 -2325 253454
rect -2283 252677 -2273 253454
rect -2125 252677 -2115 253454
rect -2073 252677 -2063 253454
rect -1915 252677 -1905 253454
rect -1863 252677 -1853 253454
rect -1705 252677 -1695 253454
rect -1653 252677 -1643 253454
rect -1495 252677 -1485 253454
rect -1443 252677 -1433 253454
rect -1285 252677 -1275 253454
rect -1233 252677 -1223 253454
rect -1075 252677 -1065 253454
rect -1023 252677 -1013 253454
rect -865 252677 -855 253454
rect -813 252677 -803 253454
rect -655 252677 -645 253454
rect -603 252677 -593 253454
rect -445 252677 -435 253454
rect -393 252677 -383 253454
rect -235 252677 -225 253454
rect -183 252677 -173 253454
rect -25 252677 -15 253454
rect 27 252677 37 253454
rect 185 252677 195 253454
rect 237 252677 247 253454
rect 395 252677 405 253454
rect 447 252677 457 253454
rect 605 252677 615 253454
rect 657 252677 667 253454
rect 815 252677 825 253454
rect 867 252677 877 253454
rect 1025 252677 1035 253454
rect 1077 252677 1087 253454
rect 1235 252677 1245 253454
rect 1287 252677 1297 253454
rect 1445 252677 1455 253454
rect 1497 252677 1507 253454
rect 1655 252677 1665 253454
rect 1707 252677 1717 253454
rect 1865 252677 1875 253454
rect 1917 252677 1927 253454
rect 2075 252677 2085 253454
rect 2127 252677 2137 253454
rect 2285 252677 2295 253454
rect 2337 252677 2347 253454
rect 2495 252677 2505 253454
rect 2547 252677 2557 253454
rect 2705 252677 2715 253454
rect 2757 252677 2767 253454
rect 2915 252677 2925 253454
rect 2967 252677 2977 253454
rect 3125 252677 3135 253454
rect 3177 252677 3187 253454
rect 3335 252677 3345 253454
rect 3387 252677 3397 253454
rect 3545 252677 3555 253454
rect 3597 252677 3607 253454
rect 3755 252677 3765 253454
rect 3807 252677 3817 253454
rect 3965 252677 3975 253454
rect 4017 252677 4027 253454
rect 4175 252677 4185 253454
rect 4227 252677 4237 253454
rect 4385 252677 4395 253454
rect 4437 252677 4447 253454
rect 4595 252677 4605 253454
rect 4647 252677 4657 253454
rect 4805 252677 4815 253454
rect 4857 252677 4867 253454
rect 5015 252677 5025 253454
rect 5067 252677 5077 253454
rect 5225 252677 5235 253454
rect 5277 252677 5287 253454
rect 5435 252677 5445 253454
rect 5487 252677 5497 253454
rect 5645 252677 5655 253454
rect 5697 252677 5707 253454
rect 5855 252677 5865 253454
rect 5907 252677 5917 253454
rect 6065 252677 6075 253454
rect 6117 252677 6127 253454
rect 6275 252677 6285 253454
rect 6327 252677 6337 253454
rect 6485 252677 6495 253454
rect 6537 252677 6547 253454
rect 6695 252677 6705 253454
rect 6747 252677 6757 253454
rect 6905 252677 6915 253454
rect 6957 252677 6967 253454
rect 7115 252677 7125 253454
rect 7167 252677 7177 253454
rect 7325 252677 7335 253454
rect 7377 252677 7387 253454
rect 7535 252677 7545 253454
rect 7587 252677 7597 253454
rect 7745 252677 7755 253454
rect 7797 252677 7807 253454
rect 7955 252677 7965 253454
rect 8007 252677 8017 253454
rect 8165 252677 8175 253454
rect 8217 252677 8227 253454
rect 8375 252677 8385 253454
rect 8427 252677 8437 253454
rect 8585 252677 8595 253454
rect 8637 252677 8647 253454
rect 8795 252677 8805 253454
rect 8847 252677 8857 253454
rect 9005 252677 9015 253454
rect 9057 252677 9067 253454
rect 9215 252677 9225 253454
rect 9267 252677 9277 253454
rect 9425 252677 9435 253454
rect 9477 252677 9487 253454
rect 9635 252677 9645 253454
rect 9687 252677 9697 253454
rect 9845 252677 9855 253454
rect 9897 252677 9907 253454
rect 10055 252677 10065 253454
rect 10107 252677 10117 253454
rect 10265 252677 10275 253454
rect 10317 252677 10327 253454
rect 10475 252677 10485 253454
rect 10527 252677 10537 253454
rect 10685 252677 10695 253454
rect 10737 252677 10747 253454
rect 10895 252677 10905 253454
rect 10947 252677 10957 253454
rect 11105 252677 11115 253454
rect 11157 252677 11167 253454
rect 11315 252677 11325 253454
rect 11367 252677 11377 253454
rect 11525 252677 11535 253454
rect 11577 252677 11587 253454
rect 11735 252677 11745 253454
rect 11787 252677 11797 253454
rect 11945 252677 11955 253454
rect 11997 252677 12007 253454
rect 12155 252677 12165 253454
rect 12207 252677 12217 253454
rect 12365 252677 12375 253454
rect 12417 252677 12427 253454
rect 12575 252677 12585 253454
rect 12627 252677 12637 253454
rect 12785 252677 12795 253454
rect 12837 252677 12847 253454
rect 12995 252677 13005 253454
rect 13047 252677 13057 253454
rect 13205 252677 13215 253454
rect 13257 252677 13267 253454
rect 13415 252677 13425 253454
rect 13467 252677 13477 253454
rect 13625 252677 13635 253454
rect 13677 252677 13687 253454
rect 13835 252677 13845 253454
rect 13887 252677 13897 253454
rect 14045 252677 14055 253454
rect 14097 252677 14107 253454
rect 14255 252677 14265 253454
rect 14307 252677 14317 253454
rect 14465 252677 14475 253454
rect 14517 252677 14527 253454
rect 14675 252677 14685 253454
rect 14727 252677 14737 253454
rect 14885 252677 14895 253454
rect 14937 252677 14947 253454
rect 15095 252677 15105 253454
rect 15147 252677 15157 253454
rect 15305 252677 15315 253454
rect 15357 252677 15367 253454
rect 15515 252677 15525 253454
rect 15567 252677 15577 253454
rect 15725 252677 15735 253454
rect 15777 252677 15787 253454
rect 15935 252677 15945 253454
rect 15987 252677 15997 253454
rect 16145 252677 16155 253454
rect 16197 252677 16207 253454
rect 16355 252677 16365 253454
rect 16407 252677 16417 253454
rect 16565 252677 16575 253454
rect 16617 252677 16627 253454
rect 16775 252677 16785 253454
rect 16827 252677 16837 253454
rect 16985 252677 16995 253454
rect 17037 252677 17047 253454
rect 17195 252677 17205 253454
rect 17247 252677 17257 253454
rect 17405 252677 17415 253454
rect 17457 252677 17467 253454
rect 17615 252677 17625 253454
rect 17667 252677 17677 253454
rect 17825 252677 17835 253454
rect 17877 252677 17887 253454
rect 18035 252677 18045 253454
rect 18087 252677 18097 253454
rect 18245 252677 18255 253454
rect 18297 252677 18307 253454
rect 18455 252677 18465 253454
rect 18507 252677 18517 253454
rect 18665 252677 18675 253454
rect 18717 252677 18727 253454
rect 18875 252677 18885 253454
rect 18927 252677 18937 253454
rect 19085 252677 19095 253454
rect 19137 252677 19147 253454
rect 19295 252677 19305 253454
rect 19347 252677 19357 253454
rect 19505 252677 19515 253454
rect 19557 252677 19567 253454
rect 19715 252677 19725 253454
rect 19767 252677 19777 253454
rect 19925 252677 19935 253454
rect 19977 252677 19987 253454
rect 20135 252677 20145 253454
rect 20187 252677 20197 253454
rect 20345 252677 20355 253454
rect 20397 252677 20407 253454
rect 20555 252677 20565 253454
rect 20607 252677 20617 253454
rect 20765 252677 20775 253454
rect 20817 252677 20827 253454
rect 20975 252677 20985 253454
rect 21027 252677 21037 253454
rect 21185 252677 21195 253454
rect 21237 252677 21247 253454
rect 21395 252677 21405 253454
rect 21447 252677 21457 253454
rect 21605 252677 21615 253454
rect 21657 252677 21667 253454
rect 21815 252677 21825 253454
rect 21867 252677 21877 253454
rect 22025 252677 22035 253454
rect 22077 252677 22087 253454
rect 22235 252677 22245 253454
rect 22287 252677 22297 253454
rect 22445 252677 22455 253454
rect 22497 252677 22507 253454
rect 22655 252677 22665 253454
rect 22707 252677 22717 253454
rect 22865 252677 22875 253454
rect 22917 252677 22927 253454
rect 23075 252677 23085 253454
rect 23127 252677 23137 253454
rect 23285 252677 23295 253454
rect 23337 252677 23347 253454
rect 23495 252677 23505 253454
rect 23547 252677 23557 253454
rect 23705 252677 23715 253454
rect 23757 252677 23767 253454
rect 23915 252677 23925 253454
rect 23967 252677 23977 253454
rect 24125 252677 24135 253454
rect 24177 252677 24187 253454
rect 24335 252677 24345 253454
rect 24387 252677 24397 253454
rect 24545 252677 24555 253454
rect 24597 252677 24607 253454
rect 24755 252677 24765 253454
rect 24807 252677 24817 253454
rect 24965 252677 24975 253454
rect 25017 252677 25027 253454
rect 25175 252677 25185 253454
rect 25227 252677 25237 253454
rect 25385 252677 25395 253454
rect 25437 252677 25447 253454
rect 25595 252677 25605 253454
rect 25647 252677 25657 253454
rect 25805 252677 25815 253454
rect 25857 252677 25867 253454
rect 26015 252677 26025 253454
rect 26067 252677 26077 253454
rect 26225 252677 26235 253454
rect 26277 252677 26287 253454
rect 26435 252677 26445 253454
rect 26487 252677 26497 253454
rect 26645 252677 26655 253454
rect 26697 252677 26707 253454
rect 26855 252677 26865 253454
rect 26907 252677 26917 253454
rect 27065 252677 27075 253454
rect 27117 252677 27127 253454
rect 27275 252677 27285 253454
rect 27331 253453 27566 253465
rect 27331 252677 27337 253453
rect 27371 252677 27566 253453
rect -4055 252665 -4009 252677
rect -3959 252665 -3913 252677
rect -3845 252665 -3799 252677
rect -3749 252665 -3703 252677
rect -3635 252665 -3589 252677
rect -3539 252665 -3493 252677
rect -3425 252665 -3379 252677
rect -3329 252665 -3283 252677
rect -3215 252665 -3169 252677
rect -3119 252665 -3073 252677
rect -3005 252665 -2959 252677
rect -2909 252665 -2863 252677
rect -2795 252665 -2749 252677
rect -2699 252665 -2653 252677
rect -2585 252665 -2539 252677
rect -2489 252665 -2443 252677
rect -2375 252665 -2329 252677
rect -2279 252665 -2233 252677
rect -2165 252665 -2119 252677
rect -2069 252665 -2023 252677
rect -1955 252665 -1909 252677
rect -1859 252665 -1813 252677
rect -1745 252665 -1699 252677
rect -1649 252665 -1603 252677
rect -1535 252665 -1489 252677
rect -1439 252665 -1393 252677
rect -1325 252665 -1279 252677
rect -1229 252665 -1183 252677
rect -1115 252665 -1069 252677
rect -1019 252665 -973 252677
rect -905 252665 -859 252677
rect -809 252665 -763 252677
rect -695 252665 -649 252677
rect -599 252665 -553 252677
rect -485 252665 -439 252677
rect -389 252665 -343 252677
rect -275 252665 -229 252677
rect -179 252665 -133 252677
rect -65 252665 -19 252677
rect 31 252665 77 252677
rect 145 252665 191 252677
rect 241 252665 287 252677
rect 355 252665 401 252677
rect 451 252665 497 252677
rect 565 252665 611 252677
rect 661 252665 707 252677
rect 775 252665 821 252677
rect 871 252665 917 252677
rect 985 252665 1031 252677
rect 1081 252665 1127 252677
rect 1195 252665 1241 252677
rect 1291 252665 1337 252677
rect 1405 252665 1451 252677
rect 1501 252665 1547 252677
rect 1615 252665 1661 252677
rect 1711 252665 1757 252677
rect 1825 252665 1871 252677
rect 1921 252665 1967 252677
rect 2035 252665 2081 252677
rect 2131 252665 2177 252677
rect 2245 252665 2291 252677
rect 2341 252665 2387 252677
rect 2455 252665 2501 252677
rect 2551 252665 2597 252677
rect 2665 252665 2711 252677
rect 2761 252665 2807 252677
rect 2875 252665 2921 252677
rect 2971 252665 3017 252677
rect 3085 252665 3131 252677
rect 3181 252665 3227 252677
rect 3295 252665 3341 252677
rect 3391 252665 3437 252677
rect 3505 252665 3551 252677
rect 3601 252665 3647 252677
rect 3715 252665 3761 252677
rect 3811 252665 3857 252677
rect 3925 252665 3971 252677
rect 4021 252665 4067 252677
rect 4135 252665 4181 252677
rect 4231 252665 4277 252677
rect 4345 252665 4391 252677
rect 4441 252665 4487 252677
rect 4555 252665 4601 252677
rect 4651 252665 4697 252677
rect 4765 252665 4811 252677
rect 4861 252665 4907 252677
rect 4975 252665 5021 252677
rect 5071 252665 5117 252677
rect 5185 252665 5231 252677
rect 5281 252665 5327 252677
rect 5395 252665 5441 252677
rect 5491 252665 5537 252677
rect 5605 252665 5651 252677
rect 5701 252665 5747 252677
rect 5815 252665 5861 252677
rect 5911 252665 5957 252677
rect 6025 252665 6071 252677
rect 6121 252665 6167 252677
rect 6235 252665 6281 252677
rect 6331 252665 6377 252677
rect 6445 252665 6491 252677
rect 6541 252665 6587 252677
rect 6655 252665 6701 252677
rect 6751 252665 6797 252677
rect 6865 252665 6911 252677
rect 6961 252665 7007 252677
rect 7075 252665 7121 252677
rect 7171 252665 7217 252677
rect 7285 252665 7331 252677
rect 7381 252665 7427 252677
rect 7495 252665 7541 252677
rect 7591 252665 7637 252677
rect 7705 252665 7751 252677
rect 7801 252665 7847 252677
rect 7915 252665 7961 252677
rect 8011 252665 8057 252677
rect 8125 252665 8171 252677
rect 8221 252665 8267 252677
rect 8335 252665 8381 252677
rect 8431 252665 8477 252677
rect 8545 252665 8591 252677
rect 8641 252665 8687 252677
rect 8755 252665 8801 252677
rect 8851 252665 8897 252677
rect 8965 252665 9011 252677
rect 9061 252665 9107 252677
rect 9175 252665 9221 252677
rect 9271 252665 9317 252677
rect 9385 252665 9431 252677
rect 9481 252665 9527 252677
rect 9595 252665 9641 252677
rect 9691 252665 9737 252677
rect 9805 252665 9851 252677
rect 9901 252665 9947 252677
rect 10015 252665 10061 252677
rect 10111 252665 10157 252677
rect 10225 252665 10271 252677
rect 10321 252665 10367 252677
rect 10435 252665 10481 252677
rect 10531 252665 10577 252677
rect 10645 252665 10691 252677
rect 10741 252665 10787 252677
rect 10855 252665 10901 252677
rect 10951 252665 10997 252677
rect 11065 252665 11111 252677
rect 11161 252665 11207 252677
rect 11275 252665 11321 252677
rect 11371 252665 11417 252677
rect 11485 252665 11531 252677
rect 11581 252665 11627 252677
rect 11695 252665 11741 252677
rect 11791 252665 11837 252677
rect 11905 252665 11951 252677
rect 12001 252665 12047 252677
rect 12115 252665 12161 252677
rect 12211 252665 12257 252677
rect 12325 252665 12371 252677
rect 12421 252665 12467 252677
rect 12535 252665 12581 252677
rect 12631 252665 12677 252677
rect 12745 252665 12791 252677
rect 12841 252665 12887 252677
rect 12955 252665 13001 252677
rect 13051 252665 13097 252677
rect 13165 252665 13211 252677
rect 13261 252665 13307 252677
rect 13375 252665 13421 252677
rect 13471 252665 13517 252677
rect 13585 252665 13631 252677
rect 13681 252665 13727 252677
rect 13795 252665 13841 252677
rect 13891 252665 13937 252677
rect 14005 252665 14051 252677
rect 14101 252665 14147 252677
rect 14215 252665 14261 252677
rect 14311 252665 14357 252677
rect 14425 252665 14471 252677
rect 14521 252665 14567 252677
rect 14635 252665 14681 252677
rect 14731 252665 14777 252677
rect 14845 252665 14891 252677
rect 14941 252665 14987 252677
rect 15055 252665 15101 252677
rect 15151 252665 15197 252677
rect 15265 252665 15311 252677
rect 15361 252665 15407 252677
rect 15475 252665 15521 252677
rect 15571 252665 15617 252677
rect 15685 252665 15731 252677
rect 15781 252665 15827 252677
rect 15895 252665 15941 252677
rect 15991 252665 16037 252677
rect 16105 252665 16151 252677
rect 16201 252665 16247 252677
rect 16315 252665 16361 252677
rect 16411 252665 16457 252677
rect 16525 252665 16571 252677
rect 16621 252665 16667 252677
rect 16735 252665 16781 252677
rect 16831 252665 16877 252677
rect 16945 252665 16991 252677
rect 17041 252665 17087 252677
rect 17155 252665 17201 252677
rect 17251 252665 17297 252677
rect 17365 252665 17411 252677
rect 17461 252665 17507 252677
rect 17575 252665 17621 252677
rect 17671 252665 17717 252677
rect 17785 252665 17831 252677
rect 17881 252665 17927 252677
rect 17995 252665 18041 252677
rect 18091 252665 18137 252677
rect 18205 252665 18251 252677
rect 18301 252665 18347 252677
rect 18415 252665 18461 252677
rect 18511 252665 18557 252677
rect 18625 252665 18671 252677
rect 18721 252665 18767 252677
rect 18835 252665 18881 252677
rect 18931 252665 18977 252677
rect 19045 252665 19091 252677
rect 19141 252665 19187 252677
rect 19255 252665 19301 252677
rect 19351 252665 19397 252677
rect 19465 252665 19511 252677
rect 19561 252665 19607 252677
rect 19675 252665 19721 252677
rect 19771 252665 19817 252677
rect 19885 252665 19931 252677
rect 19981 252665 20027 252677
rect 20095 252665 20141 252677
rect 20191 252665 20237 252677
rect 20305 252665 20351 252677
rect 20401 252665 20447 252677
rect 20515 252665 20561 252677
rect 20611 252665 20657 252677
rect 20725 252665 20771 252677
rect 20821 252665 20867 252677
rect 20935 252665 20981 252677
rect 21031 252665 21077 252677
rect 21145 252665 21191 252677
rect 21241 252665 21287 252677
rect 21355 252665 21401 252677
rect 21451 252665 21497 252677
rect 21565 252665 21611 252677
rect 21661 252665 21707 252677
rect 21775 252665 21821 252677
rect 21871 252665 21917 252677
rect 21985 252665 22031 252677
rect 22081 252665 22127 252677
rect 22195 252665 22241 252677
rect 22291 252665 22337 252677
rect 22405 252665 22451 252677
rect 22501 252665 22547 252677
rect 22615 252665 22661 252677
rect 22711 252665 22757 252677
rect 22825 252665 22871 252677
rect 22921 252665 22967 252677
rect 23035 252665 23081 252677
rect 23131 252665 23177 252677
rect 23245 252665 23291 252677
rect 23341 252665 23387 252677
rect 23455 252665 23501 252677
rect 23551 252665 23597 252677
rect 23665 252665 23711 252677
rect 23761 252665 23807 252677
rect 23875 252665 23921 252677
rect 23971 252665 24017 252677
rect 24085 252665 24131 252677
rect 24181 252665 24227 252677
rect 24295 252665 24341 252677
rect 24391 252665 24437 252677
rect 24505 252665 24551 252677
rect 24601 252665 24647 252677
rect 24715 252665 24761 252677
rect 24811 252665 24857 252677
rect 24925 252665 24971 252677
rect 25021 252665 25067 252677
rect 25135 252665 25181 252677
rect 25231 252665 25277 252677
rect 25345 252665 25391 252677
rect 25441 252665 25487 252677
rect 25555 252665 25601 252677
rect 25651 252665 25697 252677
rect 25765 252665 25811 252677
rect 25861 252665 25907 252677
rect 25975 252665 26021 252677
rect 26071 252665 26117 252677
rect 26185 252665 26231 252677
rect 26281 252665 26327 252677
rect 26395 252665 26441 252677
rect 26491 252665 26537 252677
rect 26605 252665 26651 252677
rect 26701 252665 26747 252677
rect 26815 252665 26861 252677
rect 26911 252665 26957 252677
rect 27025 252665 27071 252677
rect 27121 252665 27167 252677
rect 27235 252665 27281 252677
rect 27331 252665 27566 252677
rect -4013 252618 27125 252630
rect -5008 252476 -4001 252618
rect -3967 252476 -3581 252618
rect -3547 252476 -3161 252618
rect -3127 252476 -2741 252618
rect -2707 252476 -2321 252618
rect -2287 252476 -1901 252618
rect -1867 252476 -1481 252618
rect -1447 252476 -1061 252618
rect -1027 252476 -641 252618
rect -607 252476 -221 252618
rect -187 252476 199 252618
rect 233 252476 619 252618
rect 653 252476 1039 252618
rect 1073 252476 1459 252618
rect 1493 252476 1879 252618
rect 1913 252476 2299 252618
rect 2333 252476 2719 252618
rect 2753 252476 3139 252618
rect 3173 252476 3559 252618
rect 3593 252476 3979 252618
rect 4013 252476 4399 252618
rect 4433 252476 4819 252618
rect 4853 252476 5239 252618
rect 5273 252476 5659 252618
rect 5693 252476 6079 252618
rect 6113 252476 6499 252618
rect 6533 252476 6919 252618
rect 6953 252476 7339 252618
rect 7373 252476 7759 252618
rect 7793 252476 8179 252618
rect 8213 252476 8599 252618
rect 8633 252476 9019 252618
rect 9053 252476 9439 252618
rect 9473 252476 9859 252618
rect 9893 252476 10279 252618
rect 10313 252476 10699 252618
rect 10733 252476 11119 252618
rect 11153 252476 11539 252618
rect 11573 252476 11959 252618
rect 11993 252476 12379 252618
rect 12413 252476 12799 252618
rect 12833 252476 13219 252618
rect 13253 252476 13639 252618
rect 13673 252476 14059 252618
rect 14093 252476 14479 252618
rect 14513 252476 14899 252618
rect 14933 252476 15319 252618
rect 15353 252476 15739 252618
rect 15773 252476 16159 252618
rect 16193 252476 16579 252618
rect 16613 252476 16999 252618
rect 17033 252476 17419 252618
rect 17453 252476 17839 252618
rect 17873 252476 18259 252618
rect 18293 252476 18679 252618
rect 18713 252476 19099 252618
rect 19133 252476 19519 252618
rect 19553 252476 19939 252618
rect 19973 252476 20359 252618
rect 20393 252476 20779 252618
rect 20813 252476 21199 252618
rect 21233 252476 21619 252618
rect 21653 252476 22039 252618
rect 22073 252476 22459 252618
rect 22493 252476 22879 252618
rect 22913 252476 23299 252618
rect 23333 252476 23719 252618
rect 23753 252476 24139 252618
rect 24173 252476 24559 252618
rect 24593 252476 24979 252618
rect 25013 252476 25399 252618
rect 25433 252476 25819 252618
rect 25853 252476 26239 252618
rect 26273 252476 26659 252618
rect 26693 252476 27079 252618
rect 27113 252476 27125 252618
rect -5008 251582 -4142 252476
rect -4013 252464 27125 252476
rect 27377 252429 27566 252665
rect -4055 252417 -4009 252429
rect -3959 252417 -3913 252429
rect -3845 252417 -3799 252429
rect -3749 252417 -3703 252429
rect -3635 252417 -3589 252429
rect -3539 252418 -3493 252429
rect -3425 252418 -3379 252429
rect -3329 252418 -3283 252429
rect -3215 252418 -3169 252429
rect -3119 252418 -3073 252429
rect -3005 252418 -2959 252429
rect -2909 252418 -2863 252429
rect -2795 252418 -2749 252429
rect -2699 252418 -2653 252429
rect -2585 252418 -2539 252429
rect -2489 252418 -2443 252429
rect -2375 252418 -2329 252429
rect -2279 252418 -2233 252429
rect -2165 252418 -2119 252429
rect -2069 252418 -2023 252429
rect -1955 252418 -1909 252429
rect -1859 252418 -1813 252429
rect -1745 252418 -1699 252429
rect -1649 252418 -1603 252429
rect -1535 252418 -1489 252429
rect -1439 252418 -1393 252429
rect -1325 252418 -1279 252429
rect -1229 252418 -1183 252429
rect -1115 252418 -1069 252429
rect -1019 252418 -973 252429
rect -905 252418 -859 252429
rect -809 252418 -763 252429
rect -695 252418 -649 252429
rect -599 252418 -553 252429
rect -485 252418 -439 252429
rect -389 252418 -343 252429
rect -275 252418 -229 252429
rect -179 252418 -133 252429
rect -65 252418 -19 252429
rect 31 252418 77 252429
rect 145 252418 191 252429
rect 241 252418 287 252429
rect 355 252418 401 252429
rect 451 252418 497 252429
rect 565 252418 611 252429
rect 661 252418 707 252429
rect 775 252418 821 252429
rect 871 252418 917 252429
rect 985 252418 1031 252429
rect 1081 252418 1127 252429
rect 1195 252418 1241 252429
rect 1291 252418 1337 252429
rect 1405 252418 1451 252429
rect 1501 252418 1547 252429
rect 1615 252418 1661 252429
rect 1711 252418 1757 252429
rect 1825 252418 1871 252429
rect 1921 252418 1967 252429
rect 2035 252418 2081 252429
rect 2131 252418 2177 252429
rect 2245 252418 2291 252429
rect 2341 252418 2387 252429
rect 2455 252418 2501 252429
rect 2551 252418 2597 252429
rect 2665 252418 2711 252429
rect 2761 252418 2807 252429
rect 2875 252418 2921 252429
rect 2971 252418 3017 252429
rect 3085 252418 3131 252429
rect 3181 252418 3227 252429
rect 3295 252418 3341 252429
rect 3391 252418 3437 252429
rect 3505 252418 3551 252429
rect 3601 252418 3647 252429
rect 3715 252418 3761 252429
rect 3811 252418 3857 252429
rect 3925 252418 3971 252429
rect 4021 252418 4067 252429
rect 4135 252418 4181 252429
rect 4231 252418 4277 252429
rect 4345 252418 4391 252429
rect 4441 252418 4487 252429
rect 4555 252418 4601 252429
rect 4651 252418 4697 252429
rect 4765 252418 4811 252429
rect 4861 252418 4907 252429
rect 4975 252418 5021 252429
rect 5071 252418 5117 252429
rect 5185 252418 5231 252429
rect 5281 252418 5327 252429
rect 5395 252418 5441 252429
rect 5491 252418 5537 252429
rect 5605 252418 5651 252429
rect 5701 252418 5747 252429
rect 5815 252418 5861 252429
rect 5911 252418 5957 252429
rect 6025 252418 6071 252429
rect 6121 252418 6167 252429
rect 6235 252418 6281 252429
rect 6331 252418 6377 252429
rect 6445 252418 6491 252429
rect 6541 252418 6587 252429
rect 6655 252418 6701 252429
rect 6751 252418 6797 252429
rect 6865 252418 6911 252429
rect 6961 252418 7007 252429
rect 7075 252418 7121 252429
rect 7171 252418 7217 252429
rect 7285 252418 7331 252429
rect 7381 252418 7427 252429
rect 7495 252418 7541 252429
rect 7591 252418 7637 252429
rect 7705 252418 7751 252429
rect 7801 252418 7847 252429
rect 7915 252418 7961 252429
rect 8011 252418 8057 252429
rect 8125 252418 8171 252429
rect 8221 252418 8267 252429
rect 8335 252418 8381 252429
rect 8431 252418 8477 252429
rect 8545 252418 8591 252429
rect 8641 252418 8687 252429
rect 8755 252418 8801 252429
rect 8851 252418 8897 252429
rect 8965 252418 9011 252429
rect 9061 252418 9107 252429
rect 9175 252418 9221 252429
rect 9271 252418 9317 252429
rect 9385 252418 9431 252429
rect 9481 252418 9527 252429
rect 9595 252418 9641 252429
rect 9691 252418 9737 252429
rect 9805 252418 9851 252429
rect 9901 252418 9947 252429
rect 10015 252418 10061 252429
rect 10111 252418 10157 252429
rect 10225 252418 10271 252429
rect 10321 252418 10367 252429
rect 10435 252418 10481 252429
rect 10531 252418 10577 252429
rect 10645 252418 10691 252429
rect 10741 252418 10787 252429
rect 10855 252418 10901 252429
rect 10951 252418 10997 252429
rect 11065 252418 11111 252429
rect 11161 252418 11207 252429
rect 11275 252418 11321 252429
rect 11371 252418 11417 252429
rect 11485 252418 11531 252429
rect 11581 252418 11627 252429
rect 11695 252418 11741 252429
rect 11791 252418 11837 252429
rect 11905 252418 11951 252429
rect 12001 252418 12047 252429
rect 12115 252418 12161 252429
rect 12211 252418 12257 252429
rect 12325 252418 12371 252429
rect 12421 252418 12467 252429
rect 12535 252418 12581 252429
rect 12631 252418 12677 252429
rect 12745 252418 12791 252429
rect 12841 252418 12887 252429
rect 12955 252418 13001 252429
rect 13051 252418 13097 252429
rect 13165 252418 13211 252429
rect 13261 252418 13307 252429
rect 13375 252418 13421 252429
rect 13471 252418 13517 252429
rect 13585 252418 13631 252429
rect 13681 252418 13727 252429
rect 13795 252418 13841 252429
rect 13891 252418 13937 252429
rect 14005 252418 14051 252429
rect 14101 252418 14147 252429
rect 14215 252418 14261 252429
rect 14311 252418 14357 252429
rect 14425 252418 14471 252429
rect 14521 252418 14567 252429
rect 14635 252418 14681 252429
rect 14731 252418 14777 252429
rect 14845 252418 14891 252429
rect 14941 252418 14987 252429
rect 15055 252418 15101 252429
rect 15151 252418 15197 252429
rect 15265 252418 15311 252429
rect 15361 252418 15407 252429
rect 15475 252418 15521 252429
rect 15571 252418 15617 252429
rect 15685 252418 15731 252429
rect 15781 252418 15827 252429
rect 15895 252418 15941 252429
rect 15991 252418 16037 252429
rect 16105 252418 16151 252429
rect 16201 252418 16247 252429
rect 16315 252418 16361 252429
rect 16411 252418 16457 252429
rect 16525 252418 16571 252429
rect 16621 252418 16667 252429
rect 16735 252418 16781 252429
rect 16831 252418 16877 252429
rect 16945 252418 16991 252429
rect 17041 252418 17087 252429
rect 17155 252418 17201 252429
rect 17251 252418 17297 252429
rect 17365 252418 17411 252429
rect 17461 252418 17507 252429
rect 17575 252418 17621 252429
rect 17671 252418 17717 252429
rect 17785 252418 17831 252429
rect 17881 252418 17927 252429
rect 17995 252418 18041 252429
rect 18091 252418 18137 252429
rect 18205 252418 18251 252429
rect 18301 252418 18347 252429
rect 18415 252418 18461 252429
rect 18511 252418 18557 252429
rect 18625 252418 18671 252429
rect 18721 252418 18767 252429
rect 18835 252418 18881 252429
rect 18931 252418 18977 252429
rect 19045 252418 19091 252429
rect 19141 252418 19187 252429
rect 19255 252418 19301 252429
rect 19351 252418 19397 252429
rect 19465 252418 19511 252429
rect 19561 252418 19607 252429
rect 19675 252418 19721 252429
rect 19771 252418 19817 252429
rect 19885 252418 19931 252429
rect 19981 252418 20027 252429
rect 20095 252418 20141 252429
rect 20191 252418 20237 252429
rect 20305 252418 20351 252429
rect 20401 252418 20447 252429
rect 20515 252418 20561 252429
rect 20611 252418 20657 252429
rect 20725 252418 20771 252429
rect 20821 252418 20867 252429
rect 20935 252418 20981 252429
rect 21031 252418 21077 252429
rect 21145 252418 21191 252429
rect 21241 252418 21287 252429
rect 21355 252418 21401 252429
rect 21451 252418 21497 252429
rect 21565 252418 21611 252429
rect 21661 252418 21707 252429
rect 21775 252418 21821 252429
rect 21871 252418 21917 252429
rect 21985 252418 22031 252429
rect 22081 252418 22127 252429
rect 22195 252418 22241 252429
rect 22291 252418 22337 252429
rect 22405 252418 22451 252429
rect 22501 252418 22547 252429
rect 22615 252418 22661 252429
rect 22711 252418 22757 252429
rect 22825 252418 22871 252429
rect 22921 252418 22967 252429
rect 23035 252418 23081 252429
rect 23131 252418 23177 252429
rect 23245 252418 23291 252429
rect 23341 252418 23387 252429
rect 23455 252418 23501 252429
rect 23551 252418 23597 252429
rect 23665 252418 23711 252429
rect 23761 252418 23807 252429
rect 23875 252418 23921 252429
rect 23971 252418 24017 252429
rect 24085 252418 24131 252429
rect 24181 252418 24227 252429
rect 24295 252418 24341 252429
rect 24391 252418 24437 252429
rect 24505 252418 24551 252429
rect 24601 252418 24647 252429
rect 24715 252418 24761 252429
rect 24811 252418 24857 252429
rect 24925 252418 24971 252429
rect 25021 252418 25067 252429
rect 25135 252418 25181 252429
rect 25231 252418 25277 252429
rect 25345 252418 25391 252429
rect 25441 252418 25487 252429
rect 25555 252418 25601 252429
rect 25651 252418 25697 252429
rect 25765 252418 25811 252429
rect 25861 252418 25907 252429
rect 25975 252418 26021 252429
rect 26071 252418 26117 252429
rect 26185 252418 26231 252429
rect 26281 252418 26327 252429
rect 26395 252418 26441 252429
rect 26491 252418 26537 252429
rect 26605 252418 26651 252429
rect 26701 252418 26747 252429
rect 26815 252418 26861 252429
rect 26911 252418 26957 252429
rect 27025 252418 27071 252429
rect 27121 252418 27167 252429
rect 27235 252418 27281 252429
rect -4079 251641 -4069 252417
rect -4015 251641 -4005 252417
rect -3963 251641 -3953 252417
rect -3805 251641 -3795 252417
rect -3753 251641 -3743 252417
rect -3595 251641 -3585 252417
rect -3543 251641 -3533 252418
rect -3385 251641 -3375 252418
rect -3333 251641 -3323 252418
rect -3175 251641 -3165 252418
rect -3123 251641 -3113 252418
rect -2965 251641 -2955 252418
rect -2913 251641 -2903 252418
rect -2755 251641 -2745 252418
rect -2703 251641 -2693 252418
rect -2545 251641 -2535 252418
rect -2493 251641 -2483 252418
rect -2335 251641 -2325 252418
rect -2283 251641 -2273 252418
rect -2125 251641 -2115 252418
rect -2073 251641 -2063 252418
rect -1915 251641 -1905 252418
rect -1863 251641 -1853 252418
rect -1705 251641 -1695 252418
rect -1653 251641 -1643 252418
rect -1495 251641 -1485 252418
rect -1443 251641 -1433 252418
rect -1285 251641 -1275 252418
rect -1233 251641 -1223 252418
rect -1075 251641 -1065 252418
rect -1023 251641 -1013 252418
rect -865 251641 -855 252418
rect -813 251641 -803 252418
rect -655 251641 -645 252418
rect -603 251641 -593 252418
rect -445 251641 -435 252418
rect -393 251641 -383 252418
rect -235 251641 -225 252418
rect -183 251641 -173 252418
rect -25 251641 -15 252418
rect 27 251641 37 252418
rect 185 251641 195 252418
rect 237 251641 247 252418
rect 395 251641 405 252418
rect 447 251641 457 252418
rect 605 251641 615 252418
rect 657 251641 667 252418
rect 815 251641 825 252418
rect 867 251641 877 252418
rect 1025 251641 1035 252418
rect 1077 251641 1087 252418
rect 1235 251641 1245 252418
rect 1287 251641 1297 252418
rect 1445 251641 1455 252418
rect 1497 251641 1507 252418
rect 1655 251641 1665 252418
rect 1707 251641 1717 252418
rect 1865 251641 1875 252418
rect 1917 251641 1927 252418
rect 2075 251641 2085 252418
rect 2127 251641 2137 252418
rect 2285 251641 2295 252418
rect 2337 251641 2347 252418
rect 2495 251641 2505 252418
rect 2547 251641 2557 252418
rect 2705 251641 2715 252418
rect 2757 251641 2767 252418
rect 2915 251641 2925 252418
rect 2967 251641 2977 252418
rect 3125 251641 3135 252418
rect 3177 251641 3187 252418
rect 3335 251641 3345 252418
rect 3387 251641 3397 252418
rect 3545 251641 3555 252418
rect 3597 251641 3607 252418
rect 3755 251641 3765 252418
rect 3807 251641 3817 252418
rect 3965 251641 3975 252418
rect 4017 251641 4027 252418
rect 4175 251641 4185 252418
rect 4227 251641 4237 252418
rect 4385 251641 4395 252418
rect 4437 251641 4447 252418
rect 4595 251641 4605 252418
rect 4647 251641 4657 252418
rect 4805 251641 4815 252418
rect 4857 251641 4867 252418
rect 5015 251641 5025 252418
rect 5067 251641 5077 252418
rect 5225 251641 5235 252418
rect 5277 251641 5287 252418
rect 5435 251641 5445 252418
rect 5487 251641 5497 252418
rect 5645 251641 5655 252418
rect 5697 251641 5707 252418
rect 5855 251641 5865 252418
rect 5907 251641 5917 252418
rect 6065 251641 6075 252418
rect 6117 251641 6127 252418
rect 6275 251641 6285 252418
rect 6327 251641 6337 252418
rect 6485 251641 6495 252418
rect 6537 251641 6547 252418
rect 6695 251641 6705 252418
rect 6747 251641 6757 252418
rect 6905 251641 6915 252418
rect 6957 251641 6967 252418
rect 7115 251641 7125 252418
rect 7167 251641 7177 252418
rect 7325 251641 7335 252418
rect 7377 251641 7387 252418
rect 7535 251641 7545 252418
rect 7587 251641 7597 252418
rect 7745 251641 7755 252418
rect 7797 251641 7807 252418
rect 7955 251641 7965 252418
rect 8007 251641 8017 252418
rect 8165 251641 8175 252418
rect 8217 251641 8227 252418
rect 8375 251641 8385 252418
rect 8427 251641 8437 252418
rect 8585 251641 8595 252418
rect 8637 251641 8647 252418
rect 8795 251641 8805 252418
rect 8847 251641 8857 252418
rect 9005 251641 9015 252418
rect 9057 251641 9067 252418
rect 9215 251641 9225 252418
rect 9267 251641 9277 252418
rect 9425 251641 9435 252418
rect 9477 251641 9487 252418
rect 9635 251641 9645 252418
rect 9687 251641 9697 252418
rect 9845 251641 9855 252418
rect 9897 251641 9907 252418
rect 10055 251641 10065 252418
rect 10107 251641 10117 252418
rect 10265 251641 10275 252418
rect 10317 251641 10327 252418
rect 10475 251641 10485 252418
rect 10527 251641 10537 252418
rect 10685 251641 10695 252418
rect 10737 251641 10747 252418
rect 10895 251641 10905 252418
rect 10947 251641 10957 252418
rect 11105 251641 11115 252418
rect 11157 251641 11167 252418
rect 11315 251641 11325 252418
rect 11367 251641 11377 252418
rect 11525 251641 11535 252418
rect 11577 251641 11587 252418
rect 11735 251641 11745 252418
rect 11787 251641 11797 252418
rect 11945 251641 11955 252418
rect 11997 251641 12007 252418
rect 12155 251641 12165 252418
rect 12207 251641 12217 252418
rect 12365 251641 12375 252418
rect 12417 251641 12427 252418
rect 12575 251641 12585 252418
rect 12627 251641 12637 252418
rect 12785 251641 12795 252418
rect 12837 251641 12847 252418
rect 12995 251641 13005 252418
rect 13047 251641 13057 252418
rect 13205 251641 13215 252418
rect 13257 251641 13267 252418
rect 13415 251641 13425 252418
rect 13467 251641 13477 252418
rect 13625 251641 13635 252418
rect 13677 251641 13687 252418
rect 13835 251641 13845 252418
rect 13887 251641 13897 252418
rect 14045 251641 14055 252418
rect 14097 251641 14107 252418
rect 14255 251641 14265 252418
rect 14307 251641 14317 252418
rect 14465 251641 14475 252418
rect 14517 251641 14527 252418
rect 14675 251641 14685 252418
rect 14727 251641 14737 252418
rect 14885 251641 14895 252418
rect 14937 251641 14947 252418
rect 15095 251641 15105 252418
rect 15147 251641 15157 252418
rect 15305 251641 15315 252418
rect 15357 251641 15367 252418
rect 15515 251641 15525 252418
rect 15567 251641 15577 252418
rect 15725 251641 15735 252418
rect 15777 251641 15787 252418
rect 15935 251641 15945 252418
rect 15987 251641 15997 252418
rect 16145 251641 16155 252418
rect 16197 251641 16207 252418
rect 16355 251641 16365 252418
rect 16407 251641 16417 252418
rect 16565 251641 16575 252418
rect 16617 251641 16627 252418
rect 16775 251641 16785 252418
rect 16827 251641 16837 252418
rect 16985 251641 16995 252418
rect 17037 251641 17047 252418
rect 17195 251641 17205 252418
rect 17247 251641 17257 252418
rect 17405 251641 17415 252418
rect 17457 251641 17467 252418
rect 17615 251641 17625 252418
rect 17667 251641 17677 252418
rect 17825 251641 17835 252418
rect 17877 251641 17887 252418
rect 18035 251641 18045 252418
rect 18087 251641 18097 252418
rect 18245 251641 18255 252418
rect 18297 251641 18307 252418
rect 18455 251641 18465 252418
rect 18507 251641 18517 252418
rect 18665 251641 18675 252418
rect 18717 251641 18727 252418
rect 18875 251641 18885 252418
rect 18927 251641 18937 252418
rect 19085 251641 19095 252418
rect 19137 251641 19147 252418
rect 19295 251641 19305 252418
rect 19347 251641 19357 252418
rect 19505 251641 19515 252418
rect 19557 251641 19567 252418
rect 19715 251641 19725 252418
rect 19767 251641 19777 252418
rect 19925 251641 19935 252418
rect 19977 251641 19987 252418
rect 20135 251641 20145 252418
rect 20187 251641 20197 252418
rect 20345 251641 20355 252418
rect 20397 251641 20407 252418
rect 20555 251641 20565 252418
rect 20607 251641 20617 252418
rect 20765 251641 20775 252418
rect 20817 251641 20827 252418
rect 20975 251641 20985 252418
rect 21027 251641 21037 252418
rect 21185 251641 21195 252418
rect 21237 251641 21247 252418
rect 21395 251641 21405 252418
rect 21447 251641 21457 252418
rect 21605 251641 21615 252418
rect 21657 251641 21667 252418
rect 21815 251641 21825 252418
rect 21867 251641 21877 252418
rect 22025 251641 22035 252418
rect 22077 251641 22087 252418
rect 22235 251641 22245 252418
rect 22287 251641 22297 252418
rect 22445 251641 22455 252418
rect 22497 251641 22507 252418
rect 22655 251641 22665 252418
rect 22707 251641 22717 252418
rect 22865 251641 22875 252418
rect 22917 251641 22927 252418
rect 23075 251641 23085 252418
rect 23127 251641 23137 252418
rect 23285 251641 23295 252418
rect 23337 251641 23347 252418
rect 23495 251641 23505 252418
rect 23547 251641 23557 252418
rect 23705 251641 23715 252418
rect 23757 251641 23767 252418
rect 23915 251641 23925 252418
rect 23967 251641 23977 252418
rect 24125 251641 24135 252418
rect 24177 251641 24187 252418
rect 24335 251641 24345 252418
rect 24387 251641 24397 252418
rect 24545 251641 24555 252418
rect 24597 251641 24607 252418
rect 24755 251641 24765 252418
rect 24807 251641 24817 252418
rect 24965 251641 24975 252418
rect 25017 251641 25027 252418
rect 25175 251641 25185 252418
rect 25227 251641 25237 252418
rect 25385 251641 25395 252418
rect 25437 251641 25447 252418
rect 25595 251641 25605 252418
rect 25647 251641 25657 252418
rect 25805 251641 25815 252418
rect 25857 251641 25867 252418
rect 26015 251641 26025 252418
rect 26067 251641 26077 252418
rect 26225 251641 26235 252418
rect 26277 251641 26287 252418
rect 26435 251641 26445 252418
rect 26487 251641 26497 252418
rect 26645 251641 26655 252418
rect 26697 251641 26707 252418
rect 26855 251641 26865 252418
rect 26907 251641 26917 252418
rect 27065 251641 27075 252418
rect 27117 251641 27127 252418
rect 27275 251641 27285 252418
rect 27331 252417 27566 252429
rect 27331 251641 27337 252417
rect 27371 251641 27566 252417
rect -4055 251629 -4009 251641
rect -3959 251629 -3913 251641
rect -3845 251629 -3799 251641
rect -3749 251629 -3703 251641
rect -3635 251629 -3589 251641
rect -3539 251629 -3493 251641
rect -3425 251629 -3379 251641
rect -3329 251629 -3283 251641
rect -3215 251629 -3169 251641
rect -3119 251629 -3073 251641
rect -3005 251629 -2959 251641
rect -2909 251629 -2863 251641
rect -2795 251629 -2749 251641
rect -2699 251629 -2653 251641
rect -2585 251629 -2539 251641
rect -2489 251629 -2443 251641
rect -2375 251629 -2329 251641
rect -2279 251629 -2233 251641
rect -2165 251629 -2119 251641
rect -2069 251629 -2023 251641
rect -1955 251629 -1909 251641
rect -1859 251629 -1813 251641
rect -1745 251629 -1699 251641
rect -1649 251629 -1603 251641
rect -1535 251629 -1489 251641
rect -1439 251629 -1393 251641
rect -1325 251629 -1279 251641
rect -1229 251629 -1183 251641
rect -1115 251629 -1069 251641
rect -1019 251629 -973 251641
rect -905 251629 -859 251641
rect -809 251629 -763 251641
rect -695 251629 -649 251641
rect -599 251629 -553 251641
rect -485 251629 -439 251641
rect -389 251629 -343 251641
rect -275 251629 -229 251641
rect -179 251629 -133 251641
rect -65 251629 -19 251641
rect 31 251629 77 251641
rect 145 251629 191 251641
rect 241 251629 287 251641
rect 355 251629 401 251641
rect 451 251629 497 251641
rect 565 251629 611 251641
rect 661 251629 707 251641
rect 775 251629 821 251641
rect 871 251629 917 251641
rect 985 251629 1031 251641
rect 1081 251629 1127 251641
rect 1195 251629 1241 251641
rect 1291 251629 1337 251641
rect 1405 251629 1451 251641
rect 1501 251629 1547 251641
rect 1615 251629 1661 251641
rect 1711 251629 1757 251641
rect 1825 251629 1871 251641
rect 1921 251629 1967 251641
rect 2035 251629 2081 251641
rect 2131 251629 2177 251641
rect 2245 251629 2291 251641
rect 2341 251629 2387 251641
rect 2455 251629 2501 251641
rect 2551 251629 2597 251641
rect 2665 251629 2711 251641
rect 2761 251629 2807 251641
rect 2875 251629 2921 251641
rect 2971 251629 3017 251641
rect 3085 251629 3131 251641
rect 3181 251629 3227 251641
rect 3295 251629 3341 251641
rect 3391 251629 3437 251641
rect 3505 251629 3551 251641
rect 3601 251629 3647 251641
rect 3715 251629 3761 251641
rect 3811 251629 3857 251641
rect 3925 251629 3971 251641
rect 4021 251629 4067 251641
rect 4135 251629 4181 251641
rect 4231 251629 4277 251641
rect 4345 251629 4391 251641
rect 4441 251629 4487 251641
rect 4555 251629 4601 251641
rect 4651 251629 4697 251641
rect 4765 251629 4811 251641
rect 4861 251629 4907 251641
rect 4975 251629 5021 251641
rect 5071 251629 5117 251641
rect 5185 251629 5231 251641
rect 5281 251629 5327 251641
rect 5395 251629 5441 251641
rect 5491 251629 5537 251641
rect 5605 251629 5651 251641
rect 5701 251629 5747 251641
rect 5815 251629 5861 251641
rect 5911 251629 5957 251641
rect 6025 251629 6071 251641
rect 6121 251629 6167 251641
rect 6235 251629 6281 251641
rect 6331 251629 6377 251641
rect 6445 251629 6491 251641
rect 6541 251629 6587 251641
rect 6655 251629 6701 251641
rect 6751 251629 6797 251641
rect 6865 251629 6911 251641
rect 6961 251629 7007 251641
rect 7075 251629 7121 251641
rect 7171 251629 7217 251641
rect 7285 251629 7331 251641
rect 7381 251629 7427 251641
rect 7495 251629 7541 251641
rect 7591 251629 7637 251641
rect 7705 251629 7751 251641
rect 7801 251629 7847 251641
rect 7915 251629 7961 251641
rect 8011 251629 8057 251641
rect 8125 251629 8171 251641
rect 8221 251629 8267 251641
rect 8335 251629 8381 251641
rect 8431 251629 8477 251641
rect 8545 251629 8591 251641
rect 8641 251629 8687 251641
rect 8755 251629 8801 251641
rect 8851 251629 8897 251641
rect 8965 251629 9011 251641
rect 9061 251629 9107 251641
rect 9175 251629 9221 251641
rect 9271 251629 9317 251641
rect 9385 251629 9431 251641
rect 9481 251629 9527 251641
rect 9595 251629 9641 251641
rect 9691 251629 9737 251641
rect 9805 251629 9851 251641
rect 9901 251629 9947 251641
rect 10015 251629 10061 251641
rect 10111 251629 10157 251641
rect 10225 251629 10271 251641
rect 10321 251629 10367 251641
rect 10435 251629 10481 251641
rect 10531 251629 10577 251641
rect 10645 251629 10691 251641
rect 10741 251629 10787 251641
rect 10855 251629 10901 251641
rect 10951 251629 10997 251641
rect 11065 251629 11111 251641
rect 11161 251629 11207 251641
rect 11275 251629 11321 251641
rect 11371 251629 11417 251641
rect 11485 251629 11531 251641
rect 11581 251629 11627 251641
rect 11695 251629 11741 251641
rect 11791 251629 11837 251641
rect 11905 251629 11951 251641
rect 12001 251629 12047 251641
rect 12115 251629 12161 251641
rect 12211 251629 12257 251641
rect 12325 251629 12371 251641
rect 12421 251629 12467 251641
rect 12535 251629 12581 251641
rect 12631 251629 12677 251641
rect 12745 251629 12791 251641
rect 12841 251629 12887 251641
rect 12955 251629 13001 251641
rect 13051 251629 13097 251641
rect 13165 251629 13211 251641
rect 13261 251629 13307 251641
rect 13375 251629 13421 251641
rect 13471 251629 13517 251641
rect 13585 251629 13631 251641
rect 13681 251629 13727 251641
rect 13795 251629 13841 251641
rect 13891 251629 13937 251641
rect 14005 251629 14051 251641
rect 14101 251629 14147 251641
rect 14215 251629 14261 251641
rect 14311 251629 14357 251641
rect 14425 251629 14471 251641
rect 14521 251629 14567 251641
rect 14635 251629 14681 251641
rect 14731 251629 14777 251641
rect 14845 251629 14891 251641
rect 14941 251629 14987 251641
rect 15055 251629 15101 251641
rect 15151 251629 15197 251641
rect 15265 251629 15311 251641
rect 15361 251629 15407 251641
rect 15475 251629 15521 251641
rect 15571 251629 15617 251641
rect 15685 251629 15731 251641
rect 15781 251629 15827 251641
rect 15895 251629 15941 251641
rect 15991 251629 16037 251641
rect 16105 251629 16151 251641
rect 16201 251629 16247 251641
rect 16315 251629 16361 251641
rect 16411 251629 16457 251641
rect 16525 251629 16571 251641
rect 16621 251629 16667 251641
rect 16735 251629 16781 251641
rect 16831 251629 16877 251641
rect 16945 251629 16991 251641
rect 17041 251629 17087 251641
rect 17155 251629 17201 251641
rect 17251 251629 17297 251641
rect 17365 251629 17411 251641
rect 17461 251629 17507 251641
rect 17575 251629 17621 251641
rect 17671 251629 17717 251641
rect 17785 251629 17831 251641
rect 17881 251629 17927 251641
rect 17995 251629 18041 251641
rect 18091 251629 18137 251641
rect 18205 251629 18251 251641
rect 18301 251629 18347 251641
rect 18415 251629 18461 251641
rect 18511 251629 18557 251641
rect 18625 251629 18671 251641
rect 18721 251629 18767 251641
rect 18835 251629 18881 251641
rect 18931 251629 18977 251641
rect 19045 251629 19091 251641
rect 19141 251629 19187 251641
rect 19255 251629 19301 251641
rect 19351 251629 19397 251641
rect 19465 251629 19511 251641
rect 19561 251629 19607 251641
rect 19675 251629 19721 251641
rect 19771 251629 19817 251641
rect 19885 251629 19931 251641
rect 19981 251629 20027 251641
rect 20095 251629 20141 251641
rect 20191 251629 20237 251641
rect 20305 251629 20351 251641
rect 20401 251629 20447 251641
rect 20515 251629 20561 251641
rect 20611 251629 20657 251641
rect 20725 251629 20771 251641
rect 20821 251629 20867 251641
rect 20935 251629 20981 251641
rect 21031 251629 21077 251641
rect 21145 251629 21191 251641
rect 21241 251629 21287 251641
rect 21355 251629 21401 251641
rect 21451 251629 21497 251641
rect 21565 251629 21611 251641
rect 21661 251629 21707 251641
rect 21775 251629 21821 251641
rect 21871 251629 21917 251641
rect 21985 251629 22031 251641
rect 22081 251629 22127 251641
rect 22195 251629 22241 251641
rect 22291 251629 22337 251641
rect 22405 251629 22451 251641
rect 22501 251629 22547 251641
rect 22615 251629 22661 251641
rect 22711 251629 22757 251641
rect 22825 251629 22871 251641
rect 22921 251629 22967 251641
rect 23035 251629 23081 251641
rect 23131 251629 23177 251641
rect 23245 251629 23291 251641
rect 23341 251629 23387 251641
rect 23455 251629 23501 251641
rect 23551 251629 23597 251641
rect 23665 251629 23711 251641
rect 23761 251629 23807 251641
rect 23875 251629 23921 251641
rect 23971 251629 24017 251641
rect 24085 251629 24131 251641
rect 24181 251629 24227 251641
rect 24295 251629 24341 251641
rect 24391 251629 24437 251641
rect 24505 251629 24551 251641
rect 24601 251629 24647 251641
rect 24715 251629 24761 251641
rect 24811 251629 24857 251641
rect 24925 251629 24971 251641
rect 25021 251629 25067 251641
rect 25135 251629 25181 251641
rect 25231 251629 25277 251641
rect 25345 251629 25391 251641
rect 25441 251629 25487 251641
rect 25555 251629 25601 251641
rect 25651 251629 25697 251641
rect 25765 251629 25811 251641
rect 25861 251629 25907 251641
rect 25975 251629 26021 251641
rect 26071 251629 26117 251641
rect 26185 251629 26231 251641
rect 26281 251629 26327 251641
rect 26395 251629 26441 251641
rect 26491 251629 26537 251641
rect 26605 251629 26651 251641
rect 26701 251629 26747 251641
rect 26815 251629 26861 251641
rect 26911 251629 26957 251641
rect 27025 251629 27071 251641
rect 27121 251629 27167 251641
rect 27235 251629 27281 251641
rect 27331 251629 27566 251641
rect -3803 251582 27335 251594
rect -5008 251440 -3791 251582
rect -3757 251440 -3371 251582
rect -3337 251440 -2951 251582
rect -2917 251440 -2531 251582
rect -2497 251440 -2111 251582
rect -2077 251440 -1691 251582
rect -1657 251440 -1271 251582
rect -1237 251440 -851 251582
rect -817 251440 -431 251582
rect -397 251440 -11 251582
rect 23 251440 409 251582
rect 443 251440 829 251582
rect 863 251440 1249 251582
rect 1283 251440 1669 251582
rect 1703 251440 2089 251582
rect 2123 251440 2509 251582
rect 2543 251440 2929 251582
rect 2963 251440 3349 251582
rect 3383 251440 3769 251582
rect 3803 251440 4189 251582
rect 4223 251440 4609 251582
rect 4643 251440 5029 251582
rect 5063 251440 5449 251582
rect 5483 251440 5869 251582
rect 5903 251440 6289 251582
rect 6323 251440 6709 251582
rect 6743 251440 7129 251582
rect 7163 251440 7549 251582
rect 7583 251440 7969 251582
rect 8003 251440 8389 251582
rect 8423 251440 8809 251582
rect 8843 251440 9229 251582
rect 9263 251440 9649 251582
rect 9683 251440 10069 251582
rect 10103 251440 10489 251582
rect 10523 251440 10909 251582
rect 10943 251440 11329 251582
rect 11363 251440 11749 251582
rect 11783 251440 12169 251582
rect 12203 251440 12589 251582
rect 12623 251440 13009 251582
rect 13043 251440 13429 251582
rect 13463 251440 13849 251582
rect 13883 251440 14269 251582
rect 14303 251440 14689 251582
rect 14723 251440 15109 251582
rect 15143 251440 15529 251582
rect 15563 251440 15949 251582
rect 15983 251440 16369 251582
rect 16403 251440 16789 251582
rect 16823 251440 17209 251582
rect 17243 251440 17629 251582
rect 17663 251440 18049 251582
rect 18083 251440 18469 251582
rect 18503 251440 18889 251582
rect 18923 251440 19309 251582
rect 19343 251440 19729 251582
rect 19763 251440 20149 251582
rect 20183 251440 20569 251582
rect 20603 251440 20989 251582
rect 21023 251440 21409 251582
rect 21443 251440 21829 251582
rect 21863 251440 22249 251582
rect 22283 251440 22669 251582
rect 22703 251440 23089 251582
rect 23123 251440 23509 251582
rect 23543 251440 23929 251582
rect 23963 251440 24349 251582
rect 24383 251440 24769 251582
rect 24803 251440 25189 251582
rect 25223 251440 25609 251582
rect 25643 251440 26029 251582
rect 26063 251440 26449 251582
rect 26483 251440 26869 251582
rect 26903 251440 27289 251582
rect 27323 251440 27335 251582
rect -5008 250546 -4142 251440
rect -3803 251428 27335 251440
rect 27377 251393 27566 251629
rect -4055 251381 -4009 251393
rect -3959 251381 -3913 251393
rect -3845 251381 -3799 251393
rect -3749 251381 -3703 251393
rect -3635 251381 -3589 251393
rect -3539 251382 -3493 251393
rect -3425 251382 -3379 251393
rect -3329 251382 -3283 251393
rect -3215 251382 -3169 251393
rect -3119 251382 -3073 251393
rect -3005 251382 -2959 251393
rect -2909 251382 -2863 251393
rect -2795 251382 -2749 251393
rect -2699 251382 -2653 251393
rect -2585 251382 -2539 251393
rect -2489 251382 -2443 251393
rect -2375 251382 -2329 251393
rect -2279 251382 -2233 251393
rect -2165 251382 -2119 251393
rect -2069 251382 -2023 251393
rect -1955 251382 -1909 251393
rect -1859 251382 -1813 251393
rect -1745 251382 -1699 251393
rect -1649 251382 -1603 251393
rect -1535 251382 -1489 251393
rect -1439 251382 -1393 251393
rect -1325 251382 -1279 251393
rect -1229 251382 -1183 251393
rect -1115 251382 -1069 251393
rect -1019 251382 -973 251393
rect -905 251382 -859 251393
rect -809 251382 -763 251393
rect -695 251382 -649 251393
rect -599 251382 -553 251393
rect -485 251382 -439 251393
rect -389 251382 -343 251393
rect -275 251382 -229 251393
rect -179 251382 -133 251393
rect -65 251382 -19 251393
rect 31 251382 77 251393
rect 145 251382 191 251393
rect 241 251382 287 251393
rect 355 251382 401 251393
rect 451 251382 497 251393
rect 565 251382 611 251393
rect 661 251382 707 251393
rect 775 251382 821 251393
rect 871 251382 917 251393
rect 985 251382 1031 251393
rect 1081 251382 1127 251393
rect 1195 251382 1241 251393
rect 1291 251382 1337 251393
rect 1405 251382 1451 251393
rect 1501 251382 1547 251393
rect 1615 251382 1661 251393
rect 1711 251382 1757 251393
rect 1825 251382 1871 251393
rect 1921 251382 1967 251393
rect 2035 251382 2081 251393
rect 2131 251382 2177 251393
rect 2245 251382 2291 251393
rect 2341 251382 2387 251393
rect 2455 251382 2501 251393
rect 2551 251382 2597 251393
rect 2665 251382 2711 251393
rect 2761 251382 2807 251393
rect 2875 251382 2921 251393
rect 2971 251382 3017 251393
rect 3085 251382 3131 251393
rect 3181 251382 3227 251393
rect 3295 251382 3341 251393
rect 3391 251382 3437 251393
rect 3505 251382 3551 251393
rect 3601 251382 3647 251393
rect 3715 251382 3761 251393
rect 3811 251382 3857 251393
rect 3925 251382 3971 251393
rect 4021 251382 4067 251393
rect 4135 251382 4181 251393
rect 4231 251382 4277 251393
rect 4345 251382 4391 251393
rect 4441 251382 4487 251393
rect 4555 251382 4601 251393
rect 4651 251382 4697 251393
rect 4765 251382 4811 251393
rect 4861 251382 4907 251393
rect 4975 251382 5021 251393
rect 5071 251382 5117 251393
rect 5185 251382 5231 251393
rect 5281 251382 5327 251393
rect 5395 251382 5441 251393
rect 5491 251382 5537 251393
rect 5605 251382 5651 251393
rect 5701 251382 5747 251393
rect 5815 251382 5861 251393
rect 5911 251382 5957 251393
rect 6025 251382 6071 251393
rect 6121 251382 6167 251393
rect 6235 251382 6281 251393
rect 6331 251382 6377 251393
rect 6445 251382 6491 251393
rect 6541 251382 6587 251393
rect 6655 251382 6701 251393
rect 6751 251382 6797 251393
rect 6865 251382 6911 251393
rect 6961 251382 7007 251393
rect 7075 251382 7121 251393
rect 7171 251382 7217 251393
rect 7285 251382 7331 251393
rect 7381 251382 7427 251393
rect 7495 251382 7541 251393
rect 7591 251382 7637 251393
rect 7705 251382 7751 251393
rect 7801 251382 7847 251393
rect 7915 251382 7961 251393
rect 8011 251382 8057 251393
rect 8125 251382 8171 251393
rect 8221 251382 8267 251393
rect 8335 251382 8381 251393
rect 8431 251382 8477 251393
rect 8545 251382 8591 251393
rect 8641 251382 8687 251393
rect 8755 251382 8801 251393
rect 8851 251382 8897 251393
rect 8965 251382 9011 251393
rect 9061 251382 9107 251393
rect 9175 251382 9221 251393
rect 9271 251382 9317 251393
rect 9385 251382 9431 251393
rect 9481 251382 9527 251393
rect 9595 251382 9641 251393
rect 9691 251382 9737 251393
rect 9805 251382 9851 251393
rect 9901 251382 9947 251393
rect 10015 251382 10061 251393
rect 10111 251382 10157 251393
rect 10225 251382 10271 251393
rect 10321 251382 10367 251393
rect 10435 251382 10481 251393
rect 10531 251382 10577 251393
rect 10645 251382 10691 251393
rect 10741 251382 10787 251393
rect 10855 251382 10901 251393
rect 10951 251382 10997 251393
rect 11065 251382 11111 251393
rect 11161 251382 11207 251393
rect 11275 251382 11321 251393
rect 11371 251382 11417 251393
rect 11485 251382 11531 251393
rect 11581 251382 11627 251393
rect 11695 251382 11741 251393
rect 11791 251382 11837 251393
rect 11905 251382 11951 251393
rect 12001 251382 12047 251393
rect 12115 251382 12161 251393
rect 12211 251382 12257 251393
rect 12325 251382 12371 251393
rect 12421 251382 12467 251393
rect 12535 251382 12581 251393
rect 12631 251382 12677 251393
rect 12745 251382 12791 251393
rect 12841 251382 12887 251393
rect 12955 251382 13001 251393
rect 13051 251382 13097 251393
rect 13165 251382 13211 251393
rect 13261 251382 13307 251393
rect 13375 251382 13421 251393
rect 13471 251382 13517 251393
rect 13585 251382 13631 251393
rect 13681 251382 13727 251393
rect 13795 251382 13841 251393
rect 13891 251382 13937 251393
rect 14005 251382 14051 251393
rect 14101 251382 14147 251393
rect 14215 251382 14261 251393
rect 14311 251382 14357 251393
rect 14425 251382 14471 251393
rect 14521 251382 14567 251393
rect 14635 251382 14681 251393
rect 14731 251382 14777 251393
rect 14845 251382 14891 251393
rect 14941 251382 14987 251393
rect 15055 251382 15101 251393
rect 15151 251382 15197 251393
rect 15265 251382 15311 251393
rect 15361 251382 15407 251393
rect 15475 251382 15521 251393
rect 15571 251382 15617 251393
rect 15685 251382 15731 251393
rect 15781 251382 15827 251393
rect 15895 251382 15941 251393
rect 15991 251382 16037 251393
rect 16105 251382 16151 251393
rect 16201 251382 16247 251393
rect 16315 251382 16361 251393
rect 16411 251382 16457 251393
rect 16525 251382 16571 251393
rect 16621 251382 16667 251393
rect 16735 251382 16781 251393
rect 16831 251382 16877 251393
rect 16945 251382 16991 251393
rect 17041 251382 17087 251393
rect 17155 251382 17201 251393
rect 17251 251382 17297 251393
rect 17365 251382 17411 251393
rect 17461 251382 17507 251393
rect 17575 251382 17621 251393
rect 17671 251382 17717 251393
rect 17785 251382 17831 251393
rect 17881 251382 17927 251393
rect 17995 251382 18041 251393
rect 18091 251382 18137 251393
rect 18205 251382 18251 251393
rect 18301 251382 18347 251393
rect 18415 251382 18461 251393
rect 18511 251382 18557 251393
rect 18625 251382 18671 251393
rect 18721 251382 18767 251393
rect 18835 251382 18881 251393
rect 18931 251382 18977 251393
rect 19045 251382 19091 251393
rect 19141 251382 19187 251393
rect 19255 251382 19301 251393
rect 19351 251382 19397 251393
rect 19465 251382 19511 251393
rect 19561 251382 19607 251393
rect 19675 251382 19721 251393
rect 19771 251382 19817 251393
rect 19885 251382 19931 251393
rect 19981 251382 20027 251393
rect 20095 251382 20141 251393
rect 20191 251382 20237 251393
rect 20305 251382 20351 251393
rect 20401 251382 20447 251393
rect 20515 251382 20561 251393
rect 20611 251382 20657 251393
rect 20725 251382 20771 251393
rect 20821 251382 20867 251393
rect 20935 251382 20981 251393
rect 21031 251382 21077 251393
rect 21145 251382 21191 251393
rect 21241 251382 21287 251393
rect 21355 251382 21401 251393
rect 21451 251382 21497 251393
rect 21565 251382 21611 251393
rect 21661 251382 21707 251393
rect 21775 251382 21821 251393
rect 21871 251382 21917 251393
rect 21985 251382 22031 251393
rect 22081 251382 22127 251393
rect 22195 251382 22241 251393
rect 22291 251382 22337 251393
rect 22405 251382 22451 251393
rect 22501 251382 22547 251393
rect 22615 251382 22661 251393
rect 22711 251382 22757 251393
rect 22825 251382 22871 251393
rect 22921 251382 22967 251393
rect 23035 251382 23081 251393
rect 23131 251382 23177 251393
rect 23245 251382 23291 251393
rect 23341 251382 23387 251393
rect 23455 251382 23501 251393
rect 23551 251382 23597 251393
rect 23665 251382 23711 251393
rect 23761 251382 23807 251393
rect 23875 251382 23921 251393
rect 23971 251382 24017 251393
rect 24085 251382 24131 251393
rect 24181 251382 24227 251393
rect 24295 251382 24341 251393
rect 24391 251382 24437 251393
rect 24505 251382 24551 251393
rect 24601 251382 24647 251393
rect 24715 251382 24761 251393
rect 24811 251382 24857 251393
rect 24925 251382 24971 251393
rect 25021 251382 25067 251393
rect 25135 251382 25181 251393
rect 25231 251382 25277 251393
rect 25345 251382 25391 251393
rect 25441 251382 25487 251393
rect 25555 251382 25601 251393
rect 25651 251382 25697 251393
rect 25765 251382 25811 251393
rect 25861 251382 25907 251393
rect 25975 251382 26021 251393
rect 26071 251382 26117 251393
rect 26185 251382 26231 251393
rect 26281 251382 26327 251393
rect 26395 251382 26441 251393
rect 26491 251382 26537 251393
rect 26605 251382 26651 251393
rect 26701 251382 26747 251393
rect 26815 251382 26861 251393
rect 26911 251382 26957 251393
rect 27025 251382 27071 251393
rect 27121 251382 27167 251393
rect 27235 251382 27281 251393
rect -4079 250605 -4069 251381
rect -4015 250605 -4005 251381
rect -3963 250605 -3953 251381
rect -3805 250605 -3795 251381
rect -3753 250605 -3743 251381
rect -3595 250605 -3585 251381
rect -3543 250605 -3533 251382
rect -3385 250605 -3375 251382
rect -3333 250605 -3323 251382
rect -3175 250605 -3165 251382
rect -3123 250605 -3113 251382
rect -2965 250605 -2955 251382
rect -2913 250605 -2903 251382
rect -2755 250605 -2745 251382
rect -2703 250605 -2693 251382
rect -2545 250605 -2535 251382
rect -2493 250605 -2483 251382
rect -2335 250605 -2325 251382
rect -2283 250605 -2273 251382
rect -2125 250605 -2115 251382
rect -2073 250605 -2063 251382
rect -1915 250605 -1905 251382
rect -1863 250605 -1853 251382
rect -1705 250605 -1695 251382
rect -1653 250605 -1643 251382
rect -1495 250605 -1485 251382
rect -1443 250605 -1433 251382
rect -1285 250605 -1275 251382
rect -1233 250605 -1223 251382
rect -1075 250605 -1065 251382
rect -1023 250605 -1013 251382
rect -865 250605 -855 251382
rect -813 250605 -803 251382
rect -655 250605 -645 251382
rect -603 250605 -593 251382
rect -445 250605 -435 251382
rect -393 250605 -383 251382
rect -235 250605 -225 251382
rect -183 250605 -173 251382
rect -25 250605 -15 251382
rect 27 250605 37 251382
rect 185 250605 195 251382
rect 237 250605 247 251382
rect 395 250605 405 251382
rect 447 250605 457 251382
rect 605 250605 615 251382
rect 657 250605 667 251382
rect 815 250605 825 251382
rect 867 250605 877 251382
rect 1025 250605 1035 251382
rect 1077 250605 1087 251382
rect 1235 250605 1245 251382
rect 1287 250605 1297 251382
rect 1445 250605 1455 251382
rect 1497 250605 1507 251382
rect 1655 250605 1665 251382
rect 1707 250605 1717 251382
rect 1865 250605 1875 251382
rect 1917 250605 1927 251382
rect 2075 250605 2085 251382
rect 2127 250605 2137 251382
rect 2285 250605 2295 251382
rect 2337 250605 2347 251382
rect 2495 250605 2505 251382
rect 2547 250605 2557 251382
rect 2705 250605 2715 251382
rect 2757 250605 2767 251382
rect 2915 250605 2925 251382
rect 2967 250605 2977 251382
rect 3125 250605 3135 251382
rect 3177 250605 3187 251382
rect 3335 250605 3345 251382
rect 3387 250605 3397 251382
rect 3545 250605 3555 251382
rect 3597 250605 3607 251382
rect 3755 250605 3765 251382
rect 3807 250605 3817 251382
rect 3965 250605 3975 251382
rect 4017 250605 4027 251382
rect 4175 250605 4185 251382
rect 4227 250605 4237 251382
rect 4385 250605 4395 251382
rect 4437 250605 4447 251382
rect 4595 250605 4605 251382
rect 4647 250605 4657 251382
rect 4805 250605 4815 251382
rect 4857 250605 4867 251382
rect 5015 250605 5025 251382
rect 5067 250605 5077 251382
rect 5225 250605 5235 251382
rect 5277 250605 5287 251382
rect 5435 250605 5445 251382
rect 5487 250605 5497 251382
rect 5645 250605 5655 251382
rect 5697 250605 5707 251382
rect 5855 250605 5865 251382
rect 5907 250605 5917 251382
rect 6065 250605 6075 251382
rect 6117 250605 6127 251382
rect 6275 250605 6285 251382
rect 6327 250605 6337 251382
rect 6485 250605 6495 251382
rect 6537 250605 6547 251382
rect 6695 250605 6705 251382
rect 6747 250605 6757 251382
rect 6905 250605 6915 251382
rect 6957 250605 6967 251382
rect 7115 250605 7125 251382
rect 7167 250605 7177 251382
rect 7325 250605 7335 251382
rect 7377 250605 7387 251382
rect 7535 250605 7545 251382
rect 7587 250605 7597 251382
rect 7745 250605 7755 251382
rect 7797 250605 7807 251382
rect 7955 250605 7965 251382
rect 8007 250605 8017 251382
rect 8165 250605 8175 251382
rect 8217 250605 8227 251382
rect 8375 250605 8385 251382
rect 8427 250605 8437 251382
rect 8585 250605 8595 251382
rect 8637 250605 8647 251382
rect 8795 250605 8805 251382
rect 8847 250605 8857 251382
rect 9005 250605 9015 251382
rect 9057 250605 9067 251382
rect 9215 250605 9225 251382
rect 9267 250605 9277 251382
rect 9425 250605 9435 251382
rect 9477 250605 9487 251382
rect 9635 250605 9645 251382
rect 9687 250605 9697 251382
rect 9845 250605 9855 251382
rect 9897 250605 9907 251382
rect 10055 250605 10065 251382
rect 10107 250605 10117 251382
rect 10265 250605 10275 251382
rect 10317 250605 10327 251382
rect 10475 250605 10485 251382
rect 10527 250605 10537 251382
rect 10685 250605 10695 251382
rect 10737 250605 10747 251382
rect 10895 250605 10905 251382
rect 10947 250605 10957 251382
rect 11105 250605 11115 251382
rect 11157 250605 11167 251382
rect 11315 250605 11325 251382
rect 11367 250605 11377 251382
rect 11525 250605 11535 251382
rect 11577 250605 11587 251382
rect 11735 250605 11745 251382
rect 11787 250605 11797 251382
rect 11945 250605 11955 251382
rect 11997 250605 12007 251382
rect 12155 250605 12165 251382
rect 12207 250605 12217 251382
rect 12365 250605 12375 251382
rect 12417 250605 12427 251382
rect 12575 250605 12585 251382
rect 12627 250605 12637 251382
rect 12785 250605 12795 251382
rect 12837 250605 12847 251382
rect 12995 250605 13005 251382
rect 13047 250605 13057 251382
rect 13205 250605 13215 251382
rect 13257 250605 13267 251382
rect 13415 250605 13425 251382
rect 13467 250605 13477 251382
rect 13625 250605 13635 251382
rect 13677 250605 13687 251382
rect 13835 250605 13845 251382
rect 13887 250605 13897 251382
rect 14045 250605 14055 251382
rect 14097 250605 14107 251382
rect 14255 250605 14265 251382
rect 14307 250605 14317 251382
rect 14465 250605 14475 251382
rect 14517 250605 14527 251382
rect 14675 250605 14685 251382
rect 14727 250605 14737 251382
rect 14885 250605 14895 251382
rect 14937 250605 14947 251382
rect 15095 250605 15105 251382
rect 15147 250605 15157 251382
rect 15305 250605 15315 251382
rect 15357 250605 15367 251382
rect 15515 250605 15525 251382
rect 15567 250605 15577 251382
rect 15725 250605 15735 251382
rect 15777 250605 15787 251382
rect 15935 250605 15945 251382
rect 15987 250605 15997 251382
rect 16145 250605 16155 251382
rect 16197 250605 16207 251382
rect 16355 250605 16365 251382
rect 16407 250605 16417 251382
rect 16565 250605 16575 251382
rect 16617 250605 16627 251382
rect 16775 250605 16785 251382
rect 16827 250605 16837 251382
rect 16985 250605 16995 251382
rect 17037 250605 17047 251382
rect 17195 250605 17205 251382
rect 17247 250605 17257 251382
rect 17405 250605 17415 251382
rect 17457 250605 17467 251382
rect 17615 250605 17625 251382
rect 17667 250605 17677 251382
rect 17825 250605 17835 251382
rect 17877 250605 17887 251382
rect 18035 250605 18045 251382
rect 18087 250605 18097 251382
rect 18245 250605 18255 251382
rect 18297 250605 18307 251382
rect 18455 250605 18465 251382
rect 18507 250605 18517 251382
rect 18665 250605 18675 251382
rect 18717 250605 18727 251382
rect 18875 250605 18885 251382
rect 18927 250605 18937 251382
rect 19085 250605 19095 251382
rect 19137 250605 19147 251382
rect 19295 250605 19305 251382
rect 19347 250605 19357 251382
rect 19505 250605 19515 251382
rect 19557 250605 19567 251382
rect 19715 250605 19725 251382
rect 19767 250605 19777 251382
rect 19925 250605 19935 251382
rect 19977 250605 19987 251382
rect 20135 250605 20145 251382
rect 20187 250605 20197 251382
rect 20345 250605 20355 251382
rect 20397 250605 20407 251382
rect 20555 250605 20565 251382
rect 20607 250605 20617 251382
rect 20765 250605 20775 251382
rect 20817 250605 20827 251382
rect 20975 250605 20985 251382
rect 21027 250605 21037 251382
rect 21185 250605 21195 251382
rect 21237 250605 21247 251382
rect 21395 250605 21405 251382
rect 21447 250605 21457 251382
rect 21605 250605 21615 251382
rect 21657 250605 21667 251382
rect 21815 250605 21825 251382
rect 21867 250605 21877 251382
rect 22025 250605 22035 251382
rect 22077 250605 22087 251382
rect 22235 250605 22245 251382
rect 22287 250605 22297 251382
rect 22445 250605 22455 251382
rect 22497 250605 22507 251382
rect 22655 250605 22665 251382
rect 22707 250605 22717 251382
rect 22865 250605 22875 251382
rect 22917 250605 22927 251382
rect 23075 250605 23085 251382
rect 23127 250605 23137 251382
rect 23285 250605 23295 251382
rect 23337 250605 23347 251382
rect 23495 250605 23505 251382
rect 23547 250605 23557 251382
rect 23705 250605 23715 251382
rect 23757 250605 23767 251382
rect 23915 250605 23925 251382
rect 23967 250605 23977 251382
rect 24125 250605 24135 251382
rect 24177 250605 24187 251382
rect 24335 250605 24345 251382
rect 24387 250605 24397 251382
rect 24545 250605 24555 251382
rect 24597 250605 24607 251382
rect 24755 250605 24765 251382
rect 24807 250605 24817 251382
rect 24965 250605 24975 251382
rect 25017 250605 25027 251382
rect 25175 250605 25185 251382
rect 25227 250605 25237 251382
rect 25385 250605 25395 251382
rect 25437 250605 25447 251382
rect 25595 250605 25605 251382
rect 25647 250605 25657 251382
rect 25805 250605 25815 251382
rect 25857 250605 25867 251382
rect 26015 250605 26025 251382
rect 26067 250605 26077 251382
rect 26225 250605 26235 251382
rect 26277 250605 26287 251382
rect 26435 250605 26445 251382
rect 26487 250605 26497 251382
rect 26645 250605 26655 251382
rect 26697 250605 26707 251382
rect 26855 250605 26865 251382
rect 26907 250605 26917 251382
rect 27065 250605 27075 251382
rect 27117 250605 27127 251382
rect 27275 250605 27285 251382
rect 27331 251381 27566 251393
rect 27331 250605 27337 251381
rect 27371 250605 27566 251381
rect -4055 250593 -4009 250605
rect -3959 250593 -3913 250605
rect -3845 250593 -3799 250605
rect -3749 250593 -3703 250605
rect -3635 250593 -3589 250605
rect -3539 250593 -3493 250605
rect -3425 250593 -3379 250605
rect -3329 250593 -3283 250605
rect -3215 250593 -3169 250605
rect -3119 250593 -3073 250605
rect -3005 250593 -2959 250605
rect -2909 250593 -2863 250605
rect -2795 250593 -2749 250605
rect -2699 250593 -2653 250605
rect -2585 250593 -2539 250605
rect -2489 250593 -2443 250605
rect -2375 250593 -2329 250605
rect -2279 250593 -2233 250605
rect -2165 250593 -2119 250605
rect -2069 250593 -2023 250605
rect -1955 250593 -1909 250605
rect -1859 250593 -1813 250605
rect -1745 250593 -1699 250605
rect -1649 250593 -1603 250605
rect -1535 250593 -1489 250605
rect -1439 250593 -1393 250605
rect -1325 250593 -1279 250605
rect -1229 250593 -1183 250605
rect -1115 250593 -1069 250605
rect -1019 250593 -973 250605
rect -905 250593 -859 250605
rect -809 250593 -763 250605
rect -695 250593 -649 250605
rect -599 250593 -553 250605
rect -485 250593 -439 250605
rect -389 250593 -343 250605
rect -275 250593 -229 250605
rect -179 250593 -133 250605
rect -65 250593 -19 250605
rect 31 250593 77 250605
rect 145 250593 191 250605
rect 241 250593 287 250605
rect 355 250593 401 250605
rect 451 250593 497 250605
rect 565 250593 611 250605
rect 661 250593 707 250605
rect 775 250593 821 250605
rect 871 250593 917 250605
rect 985 250593 1031 250605
rect 1081 250593 1127 250605
rect 1195 250593 1241 250605
rect 1291 250593 1337 250605
rect 1405 250593 1451 250605
rect 1501 250593 1547 250605
rect 1615 250593 1661 250605
rect 1711 250593 1757 250605
rect 1825 250593 1871 250605
rect 1921 250593 1967 250605
rect 2035 250593 2081 250605
rect 2131 250593 2177 250605
rect 2245 250593 2291 250605
rect 2341 250593 2387 250605
rect 2455 250593 2501 250605
rect 2551 250593 2597 250605
rect 2665 250593 2711 250605
rect 2761 250593 2807 250605
rect 2875 250593 2921 250605
rect 2971 250593 3017 250605
rect 3085 250593 3131 250605
rect 3181 250593 3227 250605
rect 3295 250593 3341 250605
rect 3391 250593 3437 250605
rect 3505 250593 3551 250605
rect 3601 250593 3647 250605
rect 3715 250593 3761 250605
rect 3811 250593 3857 250605
rect 3925 250593 3971 250605
rect 4021 250593 4067 250605
rect 4135 250593 4181 250605
rect 4231 250593 4277 250605
rect 4345 250593 4391 250605
rect 4441 250593 4487 250605
rect 4555 250593 4601 250605
rect 4651 250593 4697 250605
rect 4765 250593 4811 250605
rect 4861 250593 4907 250605
rect 4975 250593 5021 250605
rect 5071 250593 5117 250605
rect 5185 250593 5231 250605
rect 5281 250593 5327 250605
rect 5395 250593 5441 250605
rect 5491 250593 5537 250605
rect 5605 250593 5651 250605
rect 5701 250593 5747 250605
rect 5815 250593 5861 250605
rect 5911 250593 5957 250605
rect 6025 250593 6071 250605
rect 6121 250593 6167 250605
rect 6235 250593 6281 250605
rect 6331 250593 6377 250605
rect 6445 250593 6491 250605
rect 6541 250593 6587 250605
rect 6655 250593 6701 250605
rect 6751 250593 6797 250605
rect 6865 250593 6911 250605
rect 6961 250593 7007 250605
rect 7075 250593 7121 250605
rect 7171 250593 7217 250605
rect 7285 250593 7331 250605
rect 7381 250593 7427 250605
rect 7495 250593 7541 250605
rect 7591 250593 7637 250605
rect 7705 250593 7751 250605
rect 7801 250593 7847 250605
rect 7915 250593 7961 250605
rect 8011 250593 8057 250605
rect 8125 250593 8171 250605
rect 8221 250593 8267 250605
rect 8335 250593 8381 250605
rect 8431 250593 8477 250605
rect 8545 250593 8591 250605
rect 8641 250593 8687 250605
rect 8755 250593 8801 250605
rect 8851 250593 8897 250605
rect 8965 250593 9011 250605
rect 9061 250593 9107 250605
rect 9175 250593 9221 250605
rect 9271 250593 9317 250605
rect 9385 250593 9431 250605
rect 9481 250593 9527 250605
rect 9595 250593 9641 250605
rect 9691 250593 9737 250605
rect 9805 250593 9851 250605
rect 9901 250593 9947 250605
rect 10015 250593 10061 250605
rect 10111 250593 10157 250605
rect 10225 250593 10271 250605
rect 10321 250593 10367 250605
rect 10435 250593 10481 250605
rect 10531 250593 10577 250605
rect 10645 250593 10691 250605
rect 10741 250593 10787 250605
rect 10855 250593 10901 250605
rect 10951 250593 10997 250605
rect 11065 250593 11111 250605
rect 11161 250593 11207 250605
rect 11275 250593 11321 250605
rect 11371 250593 11417 250605
rect 11485 250593 11531 250605
rect 11581 250593 11627 250605
rect 11695 250593 11741 250605
rect 11791 250593 11837 250605
rect 11905 250593 11951 250605
rect 12001 250593 12047 250605
rect 12115 250593 12161 250605
rect 12211 250593 12257 250605
rect 12325 250593 12371 250605
rect 12421 250593 12467 250605
rect 12535 250593 12581 250605
rect 12631 250593 12677 250605
rect 12745 250593 12791 250605
rect 12841 250593 12887 250605
rect 12955 250593 13001 250605
rect 13051 250593 13097 250605
rect 13165 250593 13211 250605
rect 13261 250593 13307 250605
rect 13375 250593 13421 250605
rect 13471 250593 13517 250605
rect 13585 250593 13631 250605
rect 13681 250593 13727 250605
rect 13795 250593 13841 250605
rect 13891 250593 13937 250605
rect 14005 250593 14051 250605
rect 14101 250593 14147 250605
rect 14215 250593 14261 250605
rect 14311 250593 14357 250605
rect 14425 250593 14471 250605
rect 14521 250593 14567 250605
rect 14635 250593 14681 250605
rect 14731 250593 14777 250605
rect 14845 250593 14891 250605
rect 14941 250593 14987 250605
rect 15055 250593 15101 250605
rect 15151 250593 15197 250605
rect 15265 250593 15311 250605
rect 15361 250593 15407 250605
rect 15475 250593 15521 250605
rect 15571 250593 15617 250605
rect 15685 250593 15731 250605
rect 15781 250593 15827 250605
rect 15895 250593 15941 250605
rect 15991 250593 16037 250605
rect 16105 250593 16151 250605
rect 16201 250593 16247 250605
rect 16315 250593 16361 250605
rect 16411 250593 16457 250605
rect 16525 250593 16571 250605
rect 16621 250593 16667 250605
rect 16735 250593 16781 250605
rect 16831 250593 16877 250605
rect 16945 250593 16991 250605
rect 17041 250593 17087 250605
rect 17155 250593 17201 250605
rect 17251 250593 17297 250605
rect 17365 250593 17411 250605
rect 17461 250593 17507 250605
rect 17575 250593 17621 250605
rect 17671 250593 17717 250605
rect 17785 250593 17831 250605
rect 17881 250593 17927 250605
rect 17995 250593 18041 250605
rect 18091 250593 18137 250605
rect 18205 250593 18251 250605
rect 18301 250593 18347 250605
rect 18415 250593 18461 250605
rect 18511 250593 18557 250605
rect 18625 250593 18671 250605
rect 18721 250593 18767 250605
rect 18835 250593 18881 250605
rect 18931 250593 18977 250605
rect 19045 250593 19091 250605
rect 19141 250593 19187 250605
rect 19255 250593 19301 250605
rect 19351 250593 19397 250605
rect 19465 250593 19511 250605
rect 19561 250593 19607 250605
rect 19675 250593 19721 250605
rect 19771 250593 19817 250605
rect 19885 250593 19931 250605
rect 19981 250593 20027 250605
rect 20095 250593 20141 250605
rect 20191 250593 20237 250605
rect 20305 250593 20351 250605
rect 20401 250593 20447 250605
rect 20515 250593 20561 250605
rect 20611 250593 20657 250605
rect 20725 250593 20771 250605
rect 20821 250593 20867 250605
rect 20935 250593 20981 250605
rect 21031 250593 21077 250605
rect 21145 250593 21191 250605
rect 21241 250593 21287 250605
rect 21355 250593 21401 250605
rect 21451 250593 21497 250605
rect 21565 250593 21611 250605
rect 21661 250593 21707 250605
rect 21775 250593 21821 250605
rect 21871 250593 21917 250605
rect 21985 250593 22031 250605
rect 22081 250593 22127 250605
rect 22195 250593 22241 250605
rect 22291 250593 22337 250605
rect 22405 250593 22451 250605
rect 22501 250593 22547 250605
rect 22615 250593 22661 250605
rect 22711 250593 22757 250605
rect 22825 250593 22871 250605
rect 22921 250593 22967 250605
rect 23035 250593 23081 250605
rect 23131 250593 23177 250605
rect 23245 250593 23291 250605
rect 23341 250593 23387 250605
rect 23455 250593 23501 250605
rect 23551 250593 23597 250605
rect 23665 250593 23711 250605
rect 23761 250593 23807 250605
rect 23875 250593 23921 250605
rect 23971 250593 24017 250605
rect 24085 250593 24131 250605
rect 24181 250593 24227 250605
rect 24295 250593 24341 250605
rect 24391 250593 24437 250605
rect 24505 250593 24551 250605
rect 24601 250593 24647 250605
rect 24715 250593 24761 250605
rect 24811 250593 24857 250605
rect 24925 250593 24971 250605
rect 25021 250593 25067 250605
rect 25135 250593 25181 250605
rect 25231 250593 25277 250605
rect 25345 250593 25391 250605
rect 25441 250593 25487 250605
rect 25555 250593 25601 250605
rect 25651 250593 25697 250605
rect 25765 250593 25811 250605
rect 25861 250593 25907 250605
rect 25975 250593 26021 250605
rect 26071 250593 26117 250605
rect 26185 250593 26231 250605
rect 26281 250593 26327 250605
rect 26395 250593 26441 250605
rect 26491 250593 26537 250605
rect 26605 250593 26651 250605
rect 26701 250593 26747 250605
rect 26815 250593 26861 250605
rect 26911 250593 26957 250605
rect 27025 250593 27071 250605
rect 27121 250593 27167 250605
rect 27235 250593 27281 250605
rect 27331 250593 27566 250605
rect -4013 250546 27125 250558
rect -5008 250404 -4001 250546
rect -3967 250404 -3581 250546
rect -3547 250404 -3161 250546
rect -3127 250404 -2741 250546
rect -2707 250404 -2321 250546
rect -2287 250404 -1901 250546
rect -1867 250404 -1481 250546
rect -1447 250404 -1061 250546
rect -1027 250404 -641 250546
rect -607 250404 -221 250546
rect -187 250404 199 250546
rect 233 250404 619 250546
rect 653 250404 1039 250546
rect 1073 250404 1459 250546
rect 1493 250404 1879 250546
rect 1913 250404 2299 250546
rect 2333 250404 2719 250546
rect 2753 250404 3139 250546
rect 3173 250404 3559 250546
rect 3593 250404 3979 250546
rect 4013 250404 4399 250546
rect 4433 250404 4819 250546
rect 4853 250404 5239 250546
rect 5273 250404 5659 250546
rect 5693 250404 6079 250546
rect 6113 250404 6499 250546
rect 6533 250404 6919 250546
rect 6953 250404 7339 250546
rect 7373 250404 7759 250546
rect 7793 250404 8179 250546
rect 8213 250404 8599 250546
rect 8633 250404 9019 250546
rect 9053 250404 9439 250546
rect 9473 250404 9859 250546
rect 9893 250404 10279 250546
rect 10313 250404 10699 250546
rect 10733 250404 11119 250546
rect 11153 250404 11539 250546
rect 11573 250404 11959 250546
rect 11993 250404 12379 250546
rect 12413 250404 12799 250546
rect 12833 250404 13219 250546
rect 13253 250404 13639 250546
rect 13673 250404 14059 250546
rect 14093 250404 14479 250546
rect 14513 250404 14899 250546
rect 14933 250404 15319 250546
rect 15353 250404 15739 250546
rect 15773 250404 16159 250546
rect 16193 250404 16579 250546
rect 16613 250404 16999 250546
rect 17033 250404 17419 250546
rect 17453 250404 17839 250546
rect 17873 250404 18259 250546
rect 18293 250404 18679 250546
rect 18713 250404 19099 250546
rect 19133 250404 19519 250546
rect 19553 250404 19939 250546
rect 19973 250404 20359 250546
rect 20393 250404 20779 250546
rect 20813 250404 21199 250546
rect 21233 250404 21619 250546
rect 21653 250404 22039 250546
rect 22073 250404 22459 250546
rect 22493 250404 22879 250546
rect 22913 250404 23299 250546
rect 23333 250404 23719 250546
rect 23753 250404 24139 250546
rect 24173 250404 24559 250546
rect 24593 250404 24979 250546
rect 25013 250404 25399 250546
rect 25433 250404 25819 250546
rect 25853 250404 26239 250546
rect 26273 250404 26659 250546
rect 26693 250404 27079 250546
rect 27113 250404 27125 250546
rect -5008 249516 -4142 250404
rect -4013 250392 27125 250404
rect 27377 250357 27566 250593
rect -4055 250345 -4009 250357
rect -3959 250345 -3913 250357
rect -3845 250345 -3799 250357
rect -3749 250345 -3703 250357
rect -3635 250345 -3589 250357
rect -3539 250346 -3493 250357
rect -3425 250346 -3379 250357
rect -3329 250346 -3283 250357
rect -3215 250346 -3169 250357
rect -3119 250346 -3073 250357
rect -3005 250346 -2959 250357
rect -2909 250346 -2863 250357
rect -2795 250346 -2749 250357
rect -2699 250346 -2653 250357
rect -2585 250346 -2539 250357
rect -2489 250346 -2443 250357
rect -2375 250346 -2329 250357
rect -2279 250346 -2233 250357
rect -2165 250346 -2119 250357
rect -2069 250346 -2023 250357
rect -1955 250346 -1909 250357
rect -1859 250346 -1813 250357
rect -1745 250346 -1699 250357
rect -1649 250346 -1603 250357
rect -1535 250346 -1489 250357
rect -1439 250346 -1393 250357
rect -1325 250346 -1279 250357
rect -1229 250346 -1183 250357
rect -1115 250346 -1069 250357
rect -1019 250346 -973 250357
rect -905 250346 -859 250357
rect -809 250346 -763 250357
rect -695 250346 -649 250357
rect -599 250346 -553 250357
rect -485 250346 -439 250357
rect -389 250346 -343 250357
rect -275 250346 -229 250357
rect -179 250346 -133 250357
rect -65 250346 -19 250357
rect 31 250346 77 250357
rect 145 250346 191 250357
rect 241 250346 287 250357
rect 355 250346 401 250357
rect 451 250346 497 250357
rect 565 250346 611 250357
rect 661 250346 707 250357
rect 775 250346 821 250357
rect 871 250346 917 250357
rect 985 250346 1031 250357
rect 1081 250346 1127 250357
rect 1195 250346 1241 250357
rect 1291 250346 1337 250357
rect 1405 250346 1451 250357
rect 1501 250346 1547 250357
rect 1615 250346 1661 250357
rect 1711 250346 1757 250357
rect 1825 250346 1871 250357
rect 1921 250346 1967 250357
rect 2035 250346 2081 250357
rect 2131 250346 2177 250357
rect 2245 250346 2291 250357
rect 2341 250346 2387 250357
rect 2455 250346 2501 250357
rect 2551 250346 2597 250357
rect 2665 250346 2711 250357
rect 2761 250346 2807 250357
rect 2875 250346 2921 250357
rect 2971 250346 3017 250357
rect 3085 250346 3131 250357
rect 3181 250346 3227 250357
rect 3295 250346 3341 250357
rect 3391 250346 3437 250357
rect 3505 250346 3551 250357
rect 3601 250346 3647 250357
rect 3715 250346 3761 250357
rect 3811 250346 3857 250357
rect 3925 250346 3971 250357
rect 4021 250346 4067 250357
rect 4135 250346 4181 250357
rect 4231 250346 4277 250357
rect 4345 250346 4391 250357
rect 4441 250346 4487 250357
rect 4555 250346 4601 250357
rect 4651 250346 4697 250357
rect 4765 250346 4811 250357
rect 4861 250346 4907 250357
rect 4975 250346 5021 250357
rect 5071 250346 5117 250357
rect 5185 250346 5231 250357
rect 5281 250346 5327 250357
rect 5395 250346 5441 250357
rect 5491 250346 5537 250357
rect 5605 250346 5651 250357
rect 5701 250346 5747 250357
rect 5815 250346 5861 250357
rect 5911 250346 5957 250357
rect 6025 250346 6071 250357
rect 6121 250346 6167 250357
rect 6235 250346 6281 250357
rect 6331 250346 6377 250357
rect 6445 250346 6491 250357
rect 6541 250346 6587 250357
rect 6655 250346 6701 250357
rect 6751 250346 6797 250357
rect 6865 250346 6911 250357
rect 6961 250346 7007 250357
rect 7075 250346 7121 250357
rect 7171 250346 7217 250357
rect 7285 250346 7331 250357
rect 7381 250346 7427 250357
rect 7495 250346 7541 250357
rect 7591 250346 7637 250357
rect 7705 250346 7751 250357
rect 7801 250346 7847 250357
rect 7915 250346 7961 250357
rect 8011 250346 8057 250357
rect 8125 250346 8171 250357
rect 8221 250346 8267 250357
rect 8335 250346 8381 250357
rect 8431 250346 8477 250357
rect 8545 250346 8591 250357
rect 8641 250346 8687 250357
rect 8755 250346 8801 250357
rect 8851 250346 8897 250357
rect 8965 250346 9011 250357
rect 9061 250346 9107 250357
rect 9175 250346 9221 250357
rect 9271 250346 9317 250357
rect 9385 250346 9431 250357
rect 9481 250346 9527 250357
rect 9595 250346 9641 250357
rect 9691 250346 9737 250357
rect 9805 250346 9851 250357
rect 9901 250346 9947 250357
rect 10015 250346 10061 250357
rect 10111 250346 10157 250357
rect 10225 250346 10271 250357
rect 10321 250346 10367 250357
rect 10435 250346 10481 250357
rect 10531 250346 10577 250357
rect 10645 250346 10691 250357
rect 10741 250346 10787 250357
rect 10855 250346 10901 250357
rect 10951 250346 10997 250357
rect 11065 250346 11111 250357
rect 11161 250346 11207 250357
rect 11275 250346 11321 250357
rect 11371 250346 11417 250357
rect 11485 250346 11531 250357
rect 11581 250346 11627 250357
rect 11695 250346 11741 250357
rect 11791 250346 11837 250357
rect 11905 250346 11951 250357
rect 12001 250346 12047 250357
rect 12115 250346 12161 250357
rect 12211 250346 12257 250357
rect 12325 250346 12371 250357
rect 12421 250346 12467 250357
rect 12535 250346 12581 250357
rect 12631 250346 12677 250357
rect 12745 250346 12791 250357
rect 12841 250346 12887 250357
rect 12955 250346 13001 250357
rect 13051 250346 13097 250357
rect 13165 250346 13211 250357
rect 13261 250346 13307 250357
rect 13375 250346 13421 250357
rect 13471 250346 13517 250357
rect 13585 250346 13631 250357
rect 13681 250346 13727 250357
rect 13795 250346 13841 250357
rect 13891 250346 13937 250357
rect 14005 250346 14051 250357
rect 14101 250346 14147 250357
rect 14215 250346 14261 250357
rect 14311 250346 14357 250357
rect 14425 250346 14471 250357
rect 14521 250346 14567 250357
rect 14635 250346 14681 250357
rect 14731 250346 14777 250357
rect 14845 250346 14891 250357
rect 14941 250346 14987 250357
rect 15055 250346 15101 250357
rect 15151 250346 15197 250357
rect 15265 250346 15311 250357
rect 15361 250346 15407 250357
rect 15475 250346 15521 250357
rect 15571 250346 15617 250357
rect 15685 250346 15731 250357
rect 15781 250346 15827 250357
rect 15895 250346 15941 250357
rect 15991 250346 16037 250357
rect 16105 250346 16151 250357
rect 16201 250346 16247 250357
rect 16315 250346 16361 250357
rect 16411 250346 16457 250357
rect 16525 250346 16571 250357
rect 16621 250346 16667 250357
rect 16735 250346 16781 250357
rect 16831 250346 16877 250357
rect 16945 250346 16991 250357
rect 17041 250346 17087 250357
rect 17155 250346 17201 250357
rect 17251 250346 17297 250357
rect 17365 250346 17411 250357
rect 17461 250346 17507 250357
rect 17575 250346 17621 250357
rect 17671 250346 17717 250357
rect 17785 250346 17831 250357
rect 17881 250346 17927 250357
rect 17995 250346 18041 250357
rect 18091 250346 18137 250357
rect 18205 250346 18251 250357
rect 18301 250346 18347 250357
rect 18415 250346 18461 250357
rect 18511 250346 18557 250357
rect 18625 250346 18671 250357
rect 18721 250346 18767 250357
rect 18835 250346 18881 250357
rect 18931 250346 18977 250357
rect 19045 250346 19091 250357
rect 19141 250346 19187 250357
rect 19255 250346 19301 250357
rect 19351 250346 19397 250357
rect 19465 250346 19511 250357
rect 19561 250346 19607 250357
rect 19675 250346 19721 250357
rect 19771 250346 19817 250357
rect 19885 250346 19931 250357
rect 19981 250346 20027 250357
rect 20095 250346 20141 250357
rect 20191 250346 20237 250357
rect 20305 250346 20351 250357
rect 20401 250346 20447 250357
rect 20515 250346 20561 250357
rect 20611 250346 20657 250357
rect 20725 250346 20771 250357
rect 20821 250346 20867 250357
rect 20935 250346 20981 250357
rect 21031 250346 21077 250357
rect 21145 250346 21191 250357
rect 21241 250346 21287 250357
rect 21355 250346 21401 250357
rect 21451 250346 21497 250357
rect 21565 250346 21611 250357
rect 21661 250346 21707 250357
rect 21775 250346 21821 250357
rect 21871 250346 21917 250357
rect 21985 250346 22031 250357
rect 22081 250346 22127 250357
rect 22195 250346 22241 250357
rect 22291 250346 22337 250357
rect 22405 250346 22451 250357
rect 22501 250346 22547 250357
rect 22615 250346 22661 250357
rect 22711 250346 22757 250357
rect 22825 250346 22871 250357
rect 22921 250346 22967 250357
rect 23035 250346 23081 250357
rect 23131 250346 23177 250357
rect 23245 250346 23291 250357
rect 23341 250346 23387 250357
rect 23455 250346 23501 250357
rect 23551 250346 23597 250357
rect 23665 250346 23711 250357
rect 23761 250346 23807 250357
rect 23875 250346 23921 250357
rect 23971 250346 24017 250357
rect 24085 250346 24131 250357
rect 24181 250346 24227 250357
rect 24295 250346 24341 250357
rect 24391 250346 24437 250357
rect 24505 250346 24551 250357
rect 24601 250346 24647 250357
rect 24715 250346 24761 250357
rect 24811 250346 24857 250357
rect 24925 250346 24971 250357
rect 25021 250346 25067 250357
rect 25135 250346 25181 250357
rect 25231 250346 25277 250357
rect 25345 250346 25391 250357
rect 25441 250346 25487 250357
rect 25555 250346 25601 250357
rect 25651 250346 25697 250357
rect 25765 250346 25811 250357
rect 25861 250346 25907 250357
rect 25975 250346 26021 250357
rect 26071 250346 26117 250357
rect 26185 250346 26231 250357
rect 26281 250346 26327 250357
rect 26395 250346 26441 250357
rect 26491 250346 26537 250357
rect 26605 250346 26651 250357
rect 26701 250346 26747 250357
rect 26815 250346 26861 250357
rect 26911 250346 26957 250357
rect 27025 250346 27071 250357
rect 27121 250346 27167 250357
rect 27235 250346 27281 250357
rect -4079 249569 -4069 250345
rect -4015 249569 -4005 250345
rect -3963 249569 -3953 250345
rect -3805 249569 -3795 250345
rect -3753 249569 -3743 250345
rect -3595 249569 -3585 250345
rect -3543 249569 -3533 250346
rect -3385 249569 -3375 250346
rect -3333 249569 -3323 250346
rect -3175 249569 -3165 250346
rect -3123 249569 -3113 250346
rect -2965 249569 -2955 250346
rect -2913 249569 -2903 250346
rect -2755 249569 -2745 250346
rect -2703 249569 -2693 250346
rect -2545 249569 -2535 250346
rect -2493 249569 -2483 250346
rect -2335 249569 -2325 250346
rect -2283 249569 -2273 250346
rect -2125 249569 -2115 250346
rect -2073 249569 -2063 250346
rect -1915 249569 -1905 250346
rect -1863 249569 -1853 250346
rect -1705 249569 -1695 250346
rect -1653 249569 -1643 250346
rect -1495 249569 -1485 250346
rect -1443 249569 -1433 250346
rect -1285 249569 -1275 250346
rect -1233 249569 -1223 250346
rect -1075 249569 -1065 250346
rect -1023 249569 -1013 250346
rect -865 249569 -855 250346
rect -813 249569 -803 250346
rect -655 249569 -645 250346
rect -603 249569 -593 250346
rect -445 249569 -435 250346
rect -393 249569 -383 250346
rect -235 249569 -225 250346
rect -183 249569 -173 250346
rect -25 249569 -15 250346
rect 27 249569 37 250346
rect 185 249569 195 250346
rect 237 249569 247 250346
rect 395 249569 405 250346
rect 447 249569 457 250346
rect 605 249569 615 250346
rect 657 249569 667 250346
rect 815 249569 825 250346
rect 867 249569 877 250346
rect 1025 249569 1035 250346
rect 1077 249569 1087 250346
rect 1235 249569 1245 250346
rect 1287 249569 1297 250346
rect 1445 249569 1455 250346
rect 1497 249569 1507 250346
rect 1655 249569 1665 250346
rect 1707 249569 1717 250346
rect 1865 249569 1875 250346
rect 1917 249569 1927 250346
rect 2075 249569 2085 250346
rect 2127 249569 2137 250346
rect 2285 249569 2295 250346
rect 2337 249569 2347 250346
rect 2495 249569 2505 250346
rect 2547 249569 2557 250346
rect 2705 249569 2715 250346
rect 2757 249569 2767 250346
rect 2915 249569 2925 250346
rect 2967 249569 2977 250346
rect 3125 249569 3135 250346
rect 3177 249569 3187 250346
rect 3335 249569 3345 250346
rect 3387 249569 3397 250346
rect 3545 249569 3555 250346
rect 3597 249569 3607 250346
rect 3755 249569 3765 250346
rect 3807 249569 3817 250346
rect 3965 249569 3975 250346
rect 4017 249569 4027 250346
rect 4175 249569 4185 250346
rect 4227 249569 4237 250346
rect 4385 249569 4395 250346
rect 4437 249569 4447 250346
rect 4595 249569 4605 250346
rect 4647 249569 4657 250346
rect 4805 249569 4815 250346
rect 4857 249569 4867 250346
rect 5015 249569 5025 250346
rect 5067 249569 5077 250346
rect 5225 249569 5235 250346
rect 5277 249569 5287 250346
rect 5435 249569 5445 250346
rect 5487 249569 5497 250346
rect 5645 249569 5655 250346
rect 5697 249569 5707 250346
rect 5855 249569 5865 250346
rect 5907 249569 5917 250346
rect 6065 249569 6075 250346
rect 6117 249569 6127 250346
rect 6275 249569 6285 250346
rect 6327 249569 6337 250346
rect 6485 249569 6495 250346
rect 6537 249569 6547 250346
rect 6695 249569 6705 250346
rect 6747 249569 6757 250346
rect 6905 249569 6915 250346
rect 6957 249569 6967 250346
rect 7115 249569 7125 250346
rect 7167 249569 7177 250346
rect 7325 249569 7335 250346
rect 7377 249569 7387 250346
rect 7535 249569 7545 250346
rect 7587 249569 7597 250346
rect 7745 249569 7755 250346
rect 7797 249569 7807 250346
rect 7955 249569 7965 250346
rect 8007 249569 8017 250346
rect 8165 249569 8175 250346
rect 8217 249569 8227 250346
rect 8375 249569 8385 250346
rect 8427 249569 8437 250346
rect 8585 249569 8595 250346
rect 8637 249569 8647 250346
rect 8795 249569 8805 250346
rect 8847 249569 8857 250346
rect 9005 249569 9015 250346
rect 9057 249569 9067 250346
rect 9215 249569 9225 250346
rect 9267 249569 9277 250346
rect 9425 249569 9435 250346
rect 9477 249569 9487 250346
rect 9635 249569 9645 250346
rect 9687 249569 9697 250346
rect 9845 249569 9855 250346
rect 9897 249569 9907 250346
rect 10055 249569 10065 250346
rect 10107 249569 10117 250346
rect 10265 249569 10275 250346
rect 10317 249569 10327 250346
rect 10475 249569 10485 250346
rect 10527 249569 10537 250346
rect 10685 249569 10695 250346
rect 10737 249569 10747 250346
rect 10895 249569 10905 250346
rect 10947 249569 10957 250346
rect 11105 249569 11115 250346
rect 11157 249569 11167 250346
rect 11315 249569 11325 250346
rect 11367 249569 11377 250346
rect 11525 249569 11535 250346
rect 11577 249569 11587 250346
rect 11735 249569 11745 250346
rect 11787 249569 11797 250346
rect 11945 249569 11955 250346
rect 11997 249569 12007 250346
rect 12155 249569 12165 250346
rect 12207 249569 12217 250346
rect 12365 249569 12375 250346
rect 12417 249569 12427 250346
rect 12575 249569 12585 250346
rect 12627 249569 12637 250346
rect 12785 249569 12795 250346
rect 12837 249569 12847 250346
rect 12995 249569 13005 250346
rect 13047 249569 13057 250346
rect 13205 249569 13215 250346
rect 13257 249569 13267 250346
rect 13415 249569 13425 250346
rect 13467 249569 13477 250346
rect 13625 249569 13635 250346
rect 13677 249569 13687 250346
rect 13835 249569 13845 250346
rect 13887 249569 13897 250346
rect 14045 249569 14055 250346
rect 14097 249569 14107 250346
rect 14255 249569 14265 250346
rect 14307 249569 14317 250346
rect 14465 249569 14475 250346
rect 14517 249569 14527 250346
rect 14675 249569 14685 250346
rect 14727 249569 14737 250346
rect 14885 249569 14895 250346
rect 14937 249569 14947 250346
rect 15095 249569 15105 250346
rect 15147 249569 15157 250346
rect 15305 249569 15315 250346
rect 15357 249569 15367 250346
rect 15515 249569 15525 250346
rect 15567 249569 15577 250346
rect 15725 249569 15735 250346
rect 15777 249569 15787 250346
rect 15935 249569 15945 250346
rect 15987 249569 15997 250346
rect 16145 249569 16155 250346
rect 16197 249569 16207 250346
rect 16355 249569 16365 250346
rect 16407 249569 16417 250346
rect 16565 249569 16575 250346
rect 16617 249569 16627 250346
rect 16775 249569 16785 250346
rect 16827 249569 16837 250346
rect 16985 249569 16995 250346
rect 17037 249569 17047 250346
rect 17195 249569 17205 250346
rect 17247 249569 17257 250346
rect 17405 249569 17415 250346
rect 17457 249569 17467 250346
rect 17615 249569 17625 250346
rect 17667 249569 17677 250346
rect 17825 249569 17835 250346
rect 17877 249569 17887 250346
rect 18035 249569 18045 250346
rect 18087 249569 18097 250346
rect 18245 249569 18255 250346
rect 18297 249569 18307 250346
rect 18455 249569 18465 250346
rect 18507 249569 18517 250346
rect 18665 249569 18675 250346
rect 18717 249569 18727 250346
rect 18875 249569 18885 250346
rect 18927 249569 18937 250346
rect 19085 249569 19095 250346
rect 19137 249569 19147 250346
rect 19295 249569 19305 250346
rect 19347 249569 19357 250346
rect 19505 249569 19515 250346
rect 19557 249569 19567 250346
rect 19715 249569 19725 250346
rect 19767 249569 19777 250346
rect 19925 249569 19935 250346
rect 19977 249569 19987 250346
rect 20135 249569 20145 250346
rect 20187 249569 20197 250346
rect 20345 249569 20355 250346
rect 20397 249569 20407 250346
rect 20555 249569 20565 250346
rect 20607 249569 20617 250346
rect 20765 249569 20775 250346
rect 20817 249569 20827 250346
rect 20975 249569 20985 250346
rect 21027 249569 21037 250346
rect 21185 249569 21195 250346
rect 21237 249569 21247 250346
rect 21395 249569 21405 250346
rect 21447 249569 21457 250346
rect 21605 249569 21615 250346
rect 21657 249569 21667 250346
rect 21815 249569 21825 250346
rect 21867 249569 21877 250346
rect 22025 249569 22035 250346
rect 22077 249569 22087 250346
rect 22235 249569 22245 250346
rect 22287 249569 22297 250346
rect 22445 249569 22455 250346
rect 22497 249569 22507 250346
rect 22655 249569 22665 250346
rect 22707 249569 22717 250346
rect 22865 249569 22875 250346
rect 22917 249569 22927 250346
rect 23075 249569 23085 250346
rect 23127 249569 23137 250346
rect 23285 249569 23295 250346
rect 23337 249569 23347 250346
rect 23495 249569 23505 250346
rect 23547 249569 23557 250346
rect 23705 249569 23715 250346
rect 23757 249569 23767 250346
rect 23915 249569 23925 250346
rect 23967 249569 23977 250346
rect 24125 249569 24135 250346
rect 24177 249569 24187 250346
rect 24335 249569 24345 250346
rect 24387 249569 24397 250346
rect 24545 249569 24555 250346
rect 24597 249569 24607 250346
rect 24755 249569 24765 250346
rect 24807 249569 24817 250346
rect 24965 249569 24975 250346
rect 25017 249569 25027 250346
rect 25175 249569 25185 250346
rect 25227 249569 25237 250346
rect 25385 249569 25395 250346
rect 25437 249569 25447 250346
rect 25595 249569 25605 250346
rect 25647 249569 25657 250346
rect 25805 249569 25815 250346
rect 25857 249569 25867 250346
rect 26015 249569 26025 250346
rect 26067 249569 26077 250346
rect 26225 249569 26235 250346
rect 26277 249569 26287 250346
rect 26435 249569 26445 250346
rect 26487 249569 26497 250346
rect 26645 249569 26655 250346
rect 26697 249569 26707 250346
rect 26855 249569 26865 250346
rect 26907 249569 26917 250346
rect 27065 249569 27075 250346
rect 27117 249569 27127 250346
rect 27275 249569 27285 250346
rect 27331 250345 27566 250357
rect 27331 249569 27337 250345
rect 27371 249569 27566 250345
rect -4055 249557 -4009 249569
rect -3959 249557 -3913 249569
rect -3845 249557 -3799 249569
rect -3749 249557 -3703 249569
rect -3635 249557 -3589 249569
rect -3539 249557 -3493 249569
rect -3425 249557 -3379 249569
rect -3329 249557 -3283 249569
rect -3215 249557 -3169 249569
rect -3119 249557 -3073 249569
rect -3005 249557 -2959 249569
rect -2909 249557 -2863 249569
rect -2795 249557 -2749 249569
rect -2699 249557 -2653 249569
rect -2585 249557 -2539 249569
rect -2489 249557 -2443 249569
rect -2375 249557 -2329 249569
rect -2279 249557 -2233 249569
rect -2165 249557 -2119 249569
rect -2069 249557 -2023 249569
rect -1955 249557 -1909 249569
rect -1859 249557 -1813 249569
rect -1745 249557 -1699 249569
rect -1649 249557 -1603 249569
rect -1535 249557 -1489 249569
rect -1439 249557 -1393 249569
rect -1325 249557 -1279 249569
rect -1229 249557 -1183 249569
rect -1115 249557 -1069 249569
rect -1019 249557 -973 249569
rect -905 249557 -859 249569
rect -809 249557 -763 249569
rect -695 249557 -649 249569
rect -599 249557 -553 249569
rect -485 249557 -439 249569
rect -389 249557 -343 249569
rect -275 249557 -229 249569
rect -179 249557 -133 249569
rect -65 249557 -19 249569
rect 31 249557 77 249569
rect 145 249557 191 249569
rect 241 249557 287 249569
rect 355 249557 401 249569
rect 451 249557 497 249569
rect 565 249557 611 249569
rect 661 249557 707 249569
rect 775 249557 821 249569
rect 871 249557 917 249569
rect 985 249557 1031 249569
rect 1081 249557 1127 249569
rect 1195 249557 1241 249569
rect 1291 249557 1337 249569
rect 1405 249557 1451 249569
rect 1501 249557 1547 249569
rect 1615 249557 1661 249569
rect 1711 249557 1757 249569
rect 1825 249557 1871 249569
rect 1921 249557 1967 249569
rect 2035 249557 2081 249569
rect 2131 249557 2177 249569
rect 2245 249557 2291 249569
rect 2341 249557 2387 249569
rect 2455 249557 2501 249569
rect 2551 249557 2597 249569
rect 2665 249557 2711 249569
rect 2761 249557 2807 249569
rect 2875 249557 2921 249569
rect 2971 249557 3017 249569
rect 3085 249557 3131 249569
rect 3181 249557 3227 249569
rect 3295 249557 3341 249569
rect 3391 249557 3437 249569
rect 3505 249557 3551 249569
rect 3601 249557 3647 249569
rect 3715 249557 3761 249569
rect 3811 249557 3857 249569
rect 3925 249557 3971 249569
rect 4021 249557 4067 249569
rect 4135 249557 4181 249569
rect 4231 249557 4277 249569
rect 4345 249557 4391 249569
rect 4441 249557 4487 249569
rect 4555 249557 4601 249569
rect 4651 249557 4697 249569
rect 4765 249557 4811 249569
rect 4861 249557 4907 249569
rect 4975 249557 5021 249569
rect 5071 249557 5117 249569
rect 5185 249557 5231 249569
rect 5281 249557 5327 249569
rect 5395 249557 5441 249569
rect 5491 249557 5537 249569
rect 5605 249557 5651 249569
rect 5701 249557 5747 249569
rect 5815 249557 5861 249569
rect 5911 249557 5957 249569
rect 6025 249557 6071 249569
rect 6121 249557 6167 249569
rect 6235 249557 6281 249569
rect 6331 249557 6377 249569
rect 6445 249557 6491 249569
rect 6541 249557 6587 249569
rect 6655 249557 6701 249569
rect 6751 249557 6797 249569
rect 6865 249557 6911 249569
rect 6961 249557 7007 249569
rect 7075 249557 7121 249569
rect 7171 249557 7217 249569
rect 7285 249557 7331 249569
rect 7381 249557 7427 249569
rect 7495 249557 7541 249569
rect 7591 249557 7637 249569
rect 7705 249557 7751 249569
rect 7801 249557 7847 249569
rect 7915 249557 7961 249569
rect 8011 249557 8057 249569
rect 8125 249557 8171 249569
rect 8221 249557 8267 249569
rect 8335 249557 8381 249569
rect 8431 249557 8477 249569
rect 8545 249557 8591 249569
rect 8641 249557 8687 249569
rect 8755 249557 8801 249569
rect 8851 249557 8897 249569
rect 8965 249557 9011 249569
rect 9061 249557 9107 249569
rect 9175 249557 9221 249569
rect 9271 249557 9317 249569
rect 9385 249557 9431 249569
rect 9481 249557 9527 249569
rect 9595 249557 9641 249569
rect 9691 249557 9737 249569
rect 9805 249557 9851 249569
rect 9901 249557 9947 249569
rect 10015 249557 10061 249569
rect 10111 249557 10157 249569
rect 10225 249557 10271 249569
rect 10321 249557 10367 249569
rect 10435 249557 10481 249569
rect 10531 249557 10577 249569
rect 10645 249557 10691 249569
rect 10741 249557 10787 249569
rect 10855 249557 10901 249569
rect 10951 249557 10997 249569
rect 11065 249557 11111 249569
rect 11161 249557 11207 249569
rect 11275 249557 11321 249569
rect 11371 249557 11417 249569
rect 11485 249557 11531 249569
rect 11581 249557 11627 249569
rect 11695 249557 11741 249569
rect 11791 249557 11837 249569
rect 11905 249557 11951 249569
rect 12001 249557 12047 249569
rect 12115 249557 12161 249569
rect 12211 249557 12257 249569
rect 12325 249557 12371 249569
rect 12421 249557 12467 249569
rect 12535 249557 12581 249569
rect 12631 249557 12677 249569
rect 12745 249557 12791 249569
rect 12841 249557 12887 249569
rect 12955 249557 13001 249569
rect 13051 249557 13097 249569
rect 13165 249557 13211 249569
rect 13261 249557 13307 249569
rect 13375 249557 13421 249569
rect 13471 249557 13517 249569
rect 13585 249557 13631 249569
rect 13681 249557 13727 249569
rect 13795 249557 13841 249569
rect 13891 249557 13937 249569
rect 14005 249557 14051 249569
rect 14101 249557 14147 249569
rect 14215 249557 14261 249569
rect 14311 249557 14357 249569
rect 14425 249557 14471 249569
rect 14521 249557 14567 249569
rect 14635 249557 14681 249569
rect 14731 249557 14777 249569
rect 14845 249557 14891 249569
rect 14941 249557 14987 249569
rect 15055 249557 15101 249569
rect 15151 249557 15197 249569
rect 15265 249557 15311 249569
rect 15361 249557 15407 249569
rect 15475 249557 15521 249569
rect 15571 249557 15617 249569
rect 15685 249557 15731 249569
rect 15781 249557 15827 249569
rect 15895 249557 15941 249569
rect 15991 249557 16037 249569
rect 16105 249557 16151 249569
rect 16201 249557 16247 249569
rect 16315 249557 16361 249569
rect 16411 249557 16457 249569
rect 16525 249557 16571 249569
rect 16621 249557 16667 249569
rect 16735 249557 16781 249569
rect 16831 249557 16877 249569
rect 16945 249557 16991 249569
rect 17041 249557 17087 249569
rect 17155 249557 17201 249569
rect 17251 249557 17297 249569
rect 17365 249557 17411 249569
rect 17461 249557 17507 249569
rect 17575 249557 17621 249569
rect 17671 249557 17717 249569
rect 17785 249557 17831 249569
rect 17881 249557 17927 249569
rect 17995 249557 18041 249569
rect 18091 249557 18137 249569
rect 18205 249557 18251 249569
rect 18301 249557 18347 249569
rect 18415 249557 18461 249569
rect 18511 249557 18557 249569
rect 18625 249557 18671 249569
rect 18721 249557 18767 249569
rect 18835 249557 18881 249569
rect 18931 249557 18977 249569
rect 19045 249557 19091 249569
rect 19141 249557 19187 249569
rect 19255 249557 19301 249569
rect 19351 249557 19397 249569
rect 19465 249557 19511 249569
rect 19561 249557 19607 249569
rect 19675 249557 19721 249569
rect 19771 249557 19817 249569
rect 19885 249557 19931 249569
rect 19981 249557 20027 249569
rect 20095 249557 20141 249569
rect 20191 249557 20237 249569
rect 20305 249557 20351 249569
rect 20401 249557 20447 249569
rect 20515 249557 20561 249569
rect 20611 249557 20657 249569
rect 20725 249557 20771 249569
rect 20821 249557 20867 249569
rect 20935 249557 20981 249569
rect 21031 249557 21077 249569
rect 21145 249557 21191 249569
rect 21241 249557 21287 249569
rect 21355 249557 21401 249569
rect 21451 249557 21497 249569
rect 21565 249557 21611 249569
rect 21661 249557 21707 249569
rect 21775 249557 21821 249569
rect 21871 249557 21917 249569
rect 21985 249557 22031 249569
rect 22081 249557 22127 249569
rect 22195 249557 22241 249569
rect 22291 249557 22337 249569
rect 22405 249557 22451 249569
rect 22501 249557 22547 249569
rect 22615 249557 22661 249569
rect 22711 249557 22757 249569
rect 22825 249557 22871 249569
rect 22921 249557 22967 249569
rect 23035 249557 23081 249569
rect 23131 249557 23177 249569
rect 23245 249557 23291 249569
rect 23341 249557 23387 249569
rect 23455 249557 23501 249569
rect 23551 249557 23597 249569
rect 23665 249557 23711 249569
rect 23761 249557 23807 249569
rect 23875 249557 23921 249569
rect 23971 249557 24017 249569
rect 24085 249557 24131 249569
rect 24181 249557 24227 249569
rect 24295 249557 24341 249569
rect 24391 249557 24437 249569
rect 24505 249557 24551 249569
rect 24601 249557 24647 249569
rect 24715 249557 24761 249569
rect 24811 249557 24857 249569
rect 24925 249557 24971 249569
rect 25021 249557 25067 249569
rect 25135 249557 25181 249569
rect 25231 249557 25277 249569
rect 25345 249557 25391 249569
rect 25441 249557 25487 249569
rect 25555 249557 25601 249569
rect 25651 249557 25697 249569
rect 25765 249557 25811 249569
rect 25861 249557 25907 249569
rect 25975 249557 26021 249569
rect 26071 249557 26117 249569
rect 26185 249557 26231 249569
rect 26281 249557 26327 249569
rect 26395 249557 26441 249569
rect 26491 249557 26537 249569
rect 26605 249557 26651 249569
rect 26701 249557 26747 249569
rect 26815 249557 26861 249569
rect 26911 249557 26957 249569
rect 27025 249557 27071 249569
rect 27121 249557 27167 249569
rect 27235 249557 27281 249569
rect 27331 249557 27566 249569
rect -5008 249510 27397 249516
rect -5008 249476 -3791 249510
rect -3695 249476 -3371 249510
rect -3275 249476 -2951 249510
rect -2855 249476 -2531 249510
rect -2435 249476 -2111 249510
rect -2015 249476 -1691 249510
rect -1595 249476 -1271 249510
rect -1175 249476 -851 249510
rect -755 249476 -431 249510
rect -335 249476 -11 249510
rect 85 249476 409 249510
rect 505 249476 829 249510
rect 925 249476 1249 249510
rect 1345 249476 1669 249510
rect 1765 249476 2089 249510
rect 2185 249476 2509 249510
rect 2605 249476 2929 249510
rect 3025 249476 3349 249510
rect 3445 249476 3769 249510
rect 3865 249476 4189 249510
rect 4285 249476 4609 249510
rect 4705 249476 5029 249510
rect 5125 249476 5449 249510
rect 5545 249476 5869 249510
rect 5965 249476 6289 249510
rect 6385 249476 6709 249510
rect 6805 249476 7129 249510
rect 7225 249476 7549 249510
rect 7645 249476 7969 249510
rect 8065 249476 8389 249510
rect 8485 249476 8809 249510
rect 8905 249476 9229 249510
rect 9325 249476 9649 249510
rect 9745 249476 10069 249510
rect 10165 249476 10489 249510
rect 10585 249476 10909 249510
rect 11005 249476 11329 249510
rect 11425 249476 11749 249510
rect 11845 249476 12169 249510
rect 12265 249476 12589 249510
rect 12685 249476 13009 249510
rect 13105 249476 13429 249510
rect 13525 249476 13849 249510
rect 13945 249476 14269 249510
rect 14365 249476 14689 249510
rect 14785 249476 15109 249510
rect 15205 249476 15529 249510
rect 15625 249476 15949 249510
rect 16045 249476 16369 249510
rect 16465 249476 16789 249510
rect 16885 249476 17209 249510
rect 17305 249476 17629 249510
rect 17725 249476 18049 249510
rect 18145 249476 18469 249510
rect 18565 249476 18889 249510
rect 18985 249476 19309 249510
rect 19405 249476 19729 249510
rect 19825 249476 20149 249510
rect 20245 249476 20569 249510
rect 20665 249476 20989 249510
rect 21085 249476 21409 249510
rect 21505 249476 21829 249510
rect 21925 249476 22249 249510
rect 22345 249476 22669 249510
rect 22765 249476 23089 249510
rect 23185 249476 23509 249510
rect 23605 249476 23929 249510
rect 24025 249476 24349 249510
rect 24445 249476 24769 249510
rect 24865 249476 25189 249510
rect 25285 249476 25609 249510
rect 25705 249476 26029 249510
rect 26125 249476 26449 249510
rect 26545 249476 26869 249510
rect 26965 249476 27289 249510
rect 27385 249476 27397 249510
rect -5008 249470 27397 249476
rect -5008 249278 -4142 249470
rect 27450 249408 27566 249557
rect -4013 249278 27196 249279
rect -5008 249273 27197 249278
rect -5008 249239 -4001 249273
rect -3905 249239 -3581 249273
rect -3485 249239 -3161 249273
rect -3065 249239 -2741 249273
rect -2645 249239 -2321 249273
rect -2225 249239 -1901 249273
rect -1805 249239 -1481 249273
rect -1385 249239 -1061 249273
rect -965 249239 -641 249273
rect -545 249239 -221 249273
rect -125 249239 199 249273
rect 295 249239 619 249273
rect 715 249239 1039 249273
rect 1135 249239 1459 249273
rect 1555 249239 1879 249273
rect 1975 249239 2299 249273
rect 2395 249239 2719 249273
rect 2815 249239 3139 249273
rect 3235 249239 3559 249273
rect 3655 249239 3979 249273
rect 4075 249239 4399 249273
rect 4495 249239 4819 249273
rect 4915 249239 5239 249273
rect 5335 249239 5659 249273
rect 5755 249239 6079 249273
rect 6175 249239 6499 249273
rect 6595 249239 6919 249273
rect 7015 249239 7339 249273
rect 7435 249239 7759 249273
rect 7855 249239 8179 249273
rect 8275 249239 8599 249273
rect 8695 249239 9019 249273
rect 9115 249239 9439 249273
rect 9535 249239 9859 249273
rect 9955 249239 10279 249273
rect 10375 249239 10699 249273
rect 10795 249239 11119 249273
rect 11215 249239 11539 249273
rect 11635 249239 11959 249273
rect 12055 249239 12379 249273
rect 12475 249239 12799 249273
rect 12895 249239 13219 249273
rect 13315 249239 13639 249273
rect 13735 249239 14059 249273
rect 14155 249239 14479 249273
rect 14575 249239 14899 249273
rect 14995 249239 15319 249273
rect 15415 249239 15739 249273
rect 15835 249239 16159 249273
rect 16255 249239 16579 249273
rect 16675 249239 16999 249273
rect 17095 249239 17419 249273
rect 17515 249239 17839 249273
rect 17935 249239 18259 249273
rect 18355 249239 18679 249273
rect 18775 249239 19099 249273
rect 19195 249239 19519 249273
rect 19615 249239 19939 249273
rect 20035 249239 20359 249273
rect 20455 249239 20779 249273
rect 20875 249239 21199 249273
rect 21295 249239 21619 249273
rect 21715 249239 22039 249273
rect 22135 249239 22459 249273
rect 22555 249239 22879 249273
rect 22975 249239 23299 249273
rect 23395 249239 23719 249273
rect 23815 249239 24139 249273
rect 24235 249239 24559 249273
rect 24655 249239 24979 249273
rect 25075 249239 25399 249273
rect 25495 249239 25819 249273
rect 25915 249239 26239 249273
rect 26335 249239 26659 249273
rect 26755 249239 27079 249273
rect 27175 249239 27197 249273
rect -5008 249232 27197 249239
rect -5008 248345 -4142 249232
rect 27377 249192 27566 249408
rect -4055 249180 -4009 249192
rect -3959 249180 -3913 249192
rect -3845 249180 -3799 249192
rect -3749 249180 -3703 249192
rect -3635 249180 -3589 249192
rect -3539 249181 -3493 249192
rect -3425 249181 -3379 249192
rect -3329 249181 -3283 249192
rect -3215 249181 -3169 249192
rect -3119 249181 -3073 249192
rect -3005 249181 -2959 249192
rect -2909 249181 -2863 249192
rect -2795 249181 -2749 249192
rect -2699 249181 -2653 249192
rect -2585 249181 -2539 249192
rect -2489 249181 -2443 249192
rect -2375 249181 -2329 249192
rect -2279 249181 -2233 249192
rect -2165 249181 -2119 249192
rect -2069 249181 -2023 249192
rect -1955 249181 -1909 249192
rect -1859 249181 -1813 249192
rect -1745 249181 -1699 249192
rect -1649 249181 -1603 249192
rect -1535 249181 -1489 249192
rect -1439 249181 -1393 249192
rect -1325 249181 -1279 249192
rect -1229 249181 -1183 249192
rect -1115 249181 -1069 249192
rect -1019 249181 -973 249192
rect -905 249181 -859 249192
rect -809 249181 -763 249192
rect -695 249181 -649 249192
rect -599 249181 -553 249192
rect -485 249181 -439 249192
rect -389 249181 -343 249192
rect -275 249181 -229 249192
rect -179 249181 -133 249192
rect -65 249181 -19 249192
rect 31 249181 77 249192
rect 145 249181 191 249192
rect 241 249181 287 249192
rect 355 249181 401 249192
rect 451 249181 497 249192
rect 565 249181 611 249192
rect 661 249181 707 249192
rect 775 249181 821 249192
rect 871 249181 917 249192
rect 985 249181 1031 249192
rect 1081 249181 1127 249192
rect 1195 249181 1241 249192
rect 1291 249181 1337 249192
rect 1405 249181 1451 249192
rect 1501 249181 1547 249192
rect 1615 249181 1661 249192
rect 1711 249181 1757 249192
rect 1825 249181 1871 249192
rect 1921 249181 1967 249192
rect 2035 249181 2081 249192
rect 2131 249181 2177 249192
rect 2245 249181 2291 249192
rect 2341 249181 2387 249192
rect 2455 249181 2501 249192
rect 2551 249181 2597 249192
rect 2665 249181 2711 249192
rect 2761 249181 2807 249192
rect 2875 249181 2921 249192
rect 2971 249181 3017 249192
rect 3085 249181 3131 249192
rect 3181 249181 3227 249192
rect 3295 249181 3341 249192
rect 3391 249181 3437 249192
rect 3505 249181 3551 249192
rect 3601 249181 3647 249192
rect 3715 249181 3761 249192
rect 3811 249181 3857 249192
rect 3925 249181 3971 249192
rect 4021 249181 4067 249192
rect 4135 249181 4181 249192
rect 4231 249181 4277 249192
rect 4345 249181 4391 249192
rect 4441 249181 4487 249192
rect 4555 249181 4601 249192
rect 4651 249181 4697 249192
rect 4765 249181 4811 249192
rect 4861 249181 4907 249192
rect 4975 249181 5021 249192
rect 5071 249181 5117 249192
rect 5185 249181 5231 249192
rect 5281 249181 5327 249192
rect 5395 249181 5441 249192
rect 5491 249181 5537 249192
rect 5605 249181 5651 249192
rect 5701 249181 5747 249192
rect 5815 249181 5861 249192
rect 5911 249181 5957 249192
rect 6025 249181 6071 249192
rect 6121 249181 6167 249192
rect 6235 249181 6281 249192
rect 6331 249181 6377 249192
rect 6445 249181 6491 249192
rect 6541 249181 6587 249192
rect 6655 249181 6701 249192
rect 6751 249181 6797 249192
rect 6865 249181 6911 249192
rect 6961 249181 7007 249192
rect 7075 249181 7121 249192
rect 7171 249181 7217 249192
rect 7285 249181 7331 249192
rect 7381 249181 7427 249192
rect 7495 249181 7541 249192
rect 7591 249181 7637 249192
rect 7705 249181 7751 249192
rect 7801 249181 7847 249192
rect 7915 249181 7961 249192
rect 8011 249181 8057 249192
rect 8125 249181 8171 249192
rect 8221 249181 8267 249192
rect 8335 249181 8381 249192
rect 8431 249181 8477 249192
rect 8545 249181 8591 249192
rect 8641 249181 8687 249192
rect 8755 249181 8801 249192
rect 8851 249181 8897 249192
rect 8965 249181 9011 249192
rect 9061 249181 9107 249192
rect 9175 249181 9221 249192
rect 9271 249181 9317 249192
rect 9385 249181 9431 249192
rect 9481 249181 9527 249192
rect 9595 249181 9641 249192
rect 9691 249181 9737 249192
rect 9805 249181 9851 249192
rect 9901 249181 9947 249192
rect 10015 249181 10061 249192
rect 10111 249181 10157 249192
rect 10225 249181 10271 249192
rect 10321 249181 10367 249192
rect 10435 249181 10481 249192
rect 10531 249181 10577 249192
rect 10645 249181 10691 249192
rect 10741 249181 10787 249192
rect 10855 249181 10901 249192
rect 10951 249181 10997 249192
rect 11065 249181 11111 249192
rect 11161 249181 11207 249192
rect 11275 249181 11321 249192
rect 11371 249181 11417 249192
rect 11485 249181 11531 249192
rect 11581 249181 11627 249192
rect 11695 249181 11741 249192
rect 11791 249181 11837 249192
rect 11905 249181 11951 249192
rect 12001 249181 12047 249192
rect 12115 249181 12161 249192
rect 12211 249181 12257 249192
rect 12325 249181 12371 249192
rect 12421 249181 12467 249192
rect 12535 249181 12581 249192
rect 12631 249181 12677 249192
rect 12745 249181 12791 249192
rect 12841 249181 12887 249192
rect 12955 249181 13001 249192
rect 13051 249181 13097 249192
rect 13165 249181 13211 249192
rect 13261 249181 13307 249192
rect 13375 249181 13421 249192
rect 13471 249181 13517 249192
rect 13585 249181 13631 249192
rect 13681 249181 13727 249192
rect 13795 249181 13841 249192
rect 13891 249181 13937 249192
rect 14005 249181 14051 249192
rect 14101 249181 14147 249192
rect 14215 249181 14261 249192
rect 14311 249181 14357 249192
rect 14425 249181 14471 249192
rect 14521 249181 14567 249192
rect 14635 249181 14681 249192
rect 14731 249181 14777 249192
rect 14845 249181 14891 249192
rect 14941 249181 14987 249192
rect 15055 249181 15101 249192
rect 15151 249181 15197 249192
rect 15265 249181 15311 249192
rect 15361 249181 15407 249192
rect 15475 249181 15521 249192
rect 15571 249181 15617 249192
rect 15685 249181 15731 249192
rect 15781 249181 15827 249192
rect 15895 249181 15941 249192
rect 15991 249181 16037 249192
rect 16105 249181 16151 249192
rect 16201 249181 16247 249192
rect 16315 249181 16361 249192
rect 16411 249181 16457 249192
rect 16525 249181 16571 249192
rect 16621 249181 16667 249192
rect 16735 249181 16781 249192
rect 16831 249181 16877 249192
rect 16945 249181 16991 249192
rect 17041 249181 17087 249192
rect 17155 249181 17201 249192
rect 17251 249181 17297 249192
rect 17365 249181 17411 249192
rect 17461 249181 17507 249192
rect 17575 249181 17621 249192
rect 17671 249181 17717 249192
rect 17785 249181 17831 249192
rect 17881 249181 17927 249192
rect 17995 249181 18041 249192
rect 18091 249181 18137 249192
rect 18205 249181 18251 249192
rect 18301 249181 18347 249192
rect 18415 249181 18461 249192
rect 18511 249181 18557 249192
rect 18625 249181 18671 249192
rect 18721 249181 18767 249192
rect 18835 249181 18881 249192
rect 18931 249181 18977 249192
rect 19045 249181 19091 249192
rect 19141 249181 19187 249192
rect 19255 249181 19301 249192
rect 19351 249181 19397 249192
rect 19465 249181 19511 249192
rect 19561 249181 19607 249192
rect 19675 249181 19721 249192
rect 19771 249181 19817 249192
rect 19885 249181 19931 249192
rect 19981 249181 20027 249192
rect 20095 249181 20141 249192
rect 20191 249181 20237 249192
rect 20305 249181 20351 249192
rect 20401 249181 20447 249192
rect 20515 249181 20561 249192
rect 20611 249181 20657 249192
rect 20725 249181 20771 249192
rect 20821 249181 20867 249192
rect 20935 249181 20981 249192
rect 21031 249181 21077 249192
rect 21145 249181 21191 249192
rect 21241 249181 21287 249192
rect 21355 249181 21401 249192
rect 21451 249181 21497 249192
rect 21565 249181 21611 249192
rect 21661 249181 21707 249192
rect 21775 249181 21821 249192
rect 21871 249181 21917 249192
rect 21985 249181 22031 249192
rect 22081 249181 22127 249192
rect 22195 249181 22241 249192
rect 22291 249181 22337 249192
rect 22405 249181 22451 249192
rect 22501 249181 22547 249192
rect 22615 249181 22661 249192
rect 22711 249181 22757 249192
rect 22825 249181 22871 249192
rect 22921 249181 22967 249192
rect 23035 249181 23081 249192
rect 23131 249181 23177 249192
rect 23245 249181 23291 249192
rect 23341 249181 23387 249192
rect 23455 249181 23501 249192
rect 23551 249181 23597 249192
rect 23665 249181 23711 249192
rect 23761 249181 23807 249192
rect 23875 249181 23921 249192
rect 23971 249181 24017 249192
rect 24085 249181 24131 249192
rect 24181 249181 24227 249192
rect 24295 249181 24341 249192
rect 24391 249181 24437 249192
rect 24505 249181 24551 249192
rect 24601 249181 24647 249192
rect 24715 249181 24761 249192
rect 24811 249181 24857 249192
rect 24925 249181 24971 249192
rect 25021 249181 25067 249192
rect 25135 249181 25181 249192
rect 25231 249181 25277 249192
rect 25345 249181 25391 249192
rect 25441 249181 25487 249192
rect 25555 249181 25601 249192
rect 25651 249181 25697 249192
rect 25765 249181 25811 249192
rect 25861 249181 25907 249192
rect 25975 249181 26021 249192
rect 26071 249181 26117 249192
rect 26185 249181 26231 249192
rect 26281 249181 26327 249192
rect 26395 249181 26441 249192
rect 26491 249181 26537 249192
rect 26605 249181 26651 249192
rect 26701 249181 26747 249192
rect 26815 249181 26861 249192
rect 26911 249181 26957 249192
rect 27025 249181 27071 249192
rect 27121 249181 27167 249192
rect 27235 249181 27281 249192
rect -4085 248404 -4075 249180
rect -4015 248404 -4005 249180
rect -3963 248404 -3953 249180
rect -3805 248404 -3795 249180
rect -3753 248404 -3743 249180
rect -3595 248404 -3585 249180
rect -3543 248404 -3533 249181
rect -3385 248404 -3375 249181
rect -3333 248404 -3323 249181
rect -3175 248404 -3165 249181
rect -3123 248404 -3113 249181
rect -2965 248404 -2955 249181
rect -2913 248404 -2903 249181
rect -2755 248404 -2745 249181
rect -2703 248404 -2693 249181
rect -2545 248404 -2535 249181
rect -2493 248404 -2483 249181
rect -2335 248404 -2325 249181
rect -2283 248404 -2273 249181
rect -2125 248404 -2115 249181
rect -2073 248404 -2063 249181
rect -1915 248404 -1905 249181
rect -1863 248404 -1853 249181
rect -1705 248404 -1695 249181
rect -1653 248404 -1643 249181
rect -1495 248404 -1485 249181
rect -1443 248404 -1433 249181
rect -1285 248404 -1275 249181
rect -1233 248404 -1223 249181
rect -1075 248404 -1065 249181
rect -1023 248404 -1013 249181
rect -865 248404 -855 249181
rect -813 248404 -803 249181
rect -655 248404 -645 249181
rect -603 248404 -593 249181
rect -445 248404 -435 249181
rect -393 248404 -383 249181
rect -235 248404 -225 249181
rect -183 248404 -173 249181
rect -25 248404 -15 249181
rect 27 248404 37 249181
rect 185 248404 195 249181
rect 237 248404 247 249181
rect 395 248404 405 249181
rect 447 248404 457 249181
rect 605 248404 615 249181
rect 657 248404 667 249181
rect 815 248404 825 249181
rect 867 248404 877 249181
rect 1025 248404 1035 249181
rect 1077 248404 1087 249181
rect 1235 248404 1245 249181
rect 1287 248404 1297 249181
rect 1445 248404 1455 249181
rect 1497 248404 1507 249181
rect 1655 248404 1665 249181
rect 1707 248404 1717 249181
rect 1865 248404 1875 249181
rect 1917 248404 1927 249181
rect 2075 248404 2085 249181
rect 2127 248404 2137 249181
rect 2285 248404 2295 249181
rect 2337 248404 2347 249181
rect 2495 248404 2505 249181
rect 2547 248404 2557 249181
rect 2705 248404 2715 249181
rect 2757 248404 2767 249181
rect 2915 248404 2925 249181
rect 2967 248404 2977 249181
rect 3125 248404 3135 249181
rect 3177 248404 3187 249181
rect 3335 248404 3345 249181
rect 3387 248404 3397 249181
rect 3545 248404 3555 249181
rect 3597 248404 3607 249181
rect 3755 248404 3765 249181
rect 3807 248404 3817 249181
rect 3965 248404 3975 249181
rect 4017 248404 4027 249181
rect 4175 248404 4185 249181
rect 4227 248404 4237 249181
rect 4385 248404 4395 249181
rect 4437 248404 4447 249181
rect 4595 248404 4605 249181
rect 4647 248404 4657 249181
rect 4805 248404 4815 249181
rect 4857 248404 4867 249181
rect 5015 248404 5025 249181
rect 5067 248404 5077 249181
rect 5225 248404 5235 249181
rect 5277 248404 5287 249181
rect 5435 248404 5445 249181
rect 5487 248404 5497 249181
rect 5645 248404 5655 249181
rect 5697 248404 5707 249181
rect 5855 248404 5865 249181
rect 5907 248404 5917 249181
rect 6065 248404 6075 249181
rect 6117 248404 6127 249181
rect 6275 248404 6285 249181
rect 6327 248404 6337 249181
rect 6485 248404 6495 249181
rect 6537 248404 6547 249181
rect 6695 248404 6705 249181
rect 6747 248404 6757 249181
rect 6905 248404 6915 249181
rect 6957 248404 6967 249181
rect 7115 248404 7125 249181
rect 7167 248404 7177 249181
rect 7325 248404 7335 249181
rect 7377 248404 7387 249181
rect 7535 248404 7545 249181
rect 7587 248404 7597 249181
rect 7745 248404 7755 249181
rect 7797 248404 7807 249181
rect 7955 248404 7965 249181
rect 8007 248404 8017 249181
rect 8165 248404 8175 249181
rect 8217 248404 8227 249181
rect 8375 248404 8385 249181
rect 8427 248404 8437 249181
rect 8585 248404 8595 249181
rect 8637 248404 8647 249181
rect 8795 248404 8805 249181
rect 8847 248404 8857 249181
rect 9005 248404 9015 249181
rect 9057 248404 9067 249181
rect 9215 248404 9225 249181
rect 9267 248404 9277 249181
rect 9425 248404 9435 249181
rect 9477 248404 9487 249181
rect 9635 248404 9645 249181
rect 9687 248404 9697 249181
rect 9845 248404 9855 249181
rect 9897 248404 9907 249181
rect 10055 248404 10065 249181
rect 10107 248404 10117 249181
rect 10265 248404 10275 249181
rect 10317 248404 10327 249181
rect 10475 248404 10485 249181
rect 10527 248404 10537 249181
rect 10685 248404 10695 249181
rect 10737 248404 10747 249181
rect 10895 248404 10905 249181
rect 10947 248404 10957 249181
rect 11105 248404 11115 249181
rect 11157 248404 11167 249181
rect 11315 248404 11325 249181
rect 11367 248404 11377 249181
rect 11525 248404 11535 249181
rect 11577 248404 11587 249181
rect 11735 248404 11745 249181
rect 11787 248404 11797 249181
rect 11945 248404 11955 249181
rect 11997 248404 12007 249181
rect 12155 248404 12165 249181
rect 12207 248404 12217 249181
rect 12365 248404 12375 249181
rect 12417 248404 12427 249181
rect 12575 248404 12585 249181
rect 12627 248404 12637 249181
rect 12785 248404 12795 249181
rect 12837 248404 12847 249181
rect 12995 248404 13005 249181
rect 13047 248404 13057 249181
rect 13205 248404 13215 249181
rect 13257 248404 13267 249181
rect 13415 248404 13425 249181
rect 13467 248404 13477 249181
rect 13625 248404 13635 249181
rect 13677 248404 13687 249181
rect 13835 248404 13845 249181
rect 13887 248404 13897 249181
rect 14045 248404 14055 249181
rect 14097 248404 14107 249181
rect 14255 248404 14265 249181
rect 14307 248404 14317 249181
rect 14465 248404 14475 249181
rect 14517 248404 14527 249181
rect 14675 248404 14685 249181
rect 14727 248404 14737 249181
rect 14885 248404 14895 249181
rect 14937 248404 14947 249181
rect 15095 248404 15105 249181
rect 15147 248404 15157 249181
rect 15305 248404 15315 249181
rect 15357 248404 15367 249181
rect 15515 248404 15525 249181
rect 15567 248404 15577 249181
rect 15725 248404 15735 249181
rect 15777 248404 15787 249181
rect 15935 248404 15945 249181
rect 15987 248404 15997 249181
rect 16145 248404 16155 249181
rect 16197 248404 16207 249181
rect 16355 248404 16365 249181
rect 16407 248404 16417 249181
rect 16565 248404 16575 249181
rect 16617 248404 16627 249181
rect 16775 248404 16785 249181
rect 16827 248404 16837 249181
rect 16985 248404 16995 249181
rect 17037 248404 17047 249181
rect 17195 248404 17205 249181
rect 17247 248404 17257 249181
rect 17405 248404 17415 249181
rect 17457 248404 17467 249181
rect 17615 248404 17625 249181
rect 17667 248404 17677 249181
rect 17825 248404 17835 249181
rect 17877 248404 17887 249181
rect 18035 248404 18045 249181
rect 18087 248404 18097 249181
rect 18245 248404 18255 249181
rect 18297 248404 18307 249181
rect 18455 248404 18465 249181
rect 18507 248404 18517 249181
rect 18665 248404 18675 249181
rect 18717 248404 18727 249181
rect 18875 248404 18885 249181
rect 18927 248404 18937 249181
rect 19085 248404 19095 249181
rect 19137 248404 19147 249181
rect 19295 248404 19305 249181
rect 19347 248404 19357 249181
rect 19505 248404 19515 249181
rect 19557 248404 19567 249181
rect 19715 248404 19725 249181
rect 19767 248404 19777 249181
rect 19925 248404 19935 249181
rect 19977 248404 19987 249181
rect 20135 248404 20145 249181
rect 20187 248404 20197 249181
rect 20345 248404 20355 249181
rect 20397 248404 20407 249181
rect 20555 248404 20565 249181
rect 20607 248404 20617 249181
rect 20765 248404 20775 249181
rect 20817 248404 20827 249181
rect 20975 248404 20985 249181
rect 21027 248404 21037 249181
rect 21185 248404 21195 249181
rect 21237 248404 21247 249181
rect 21395 248404 21405 249181
rect 21447 248404 21457 249181
rect 21605 248404 21615 249181
rect 21657 248404 21667 249181
rect 21815 248404 21825 249181
rect 21867 248404 21877 249181
rect 22025 248404 22035 249181
rect 22077 248404 22087 249181
rect 22235 248404 22245 249181
rect 22287 248404 22297 249181
rect 22445 248404 22455 249181
rect 22497 248404 22507 249181
rect 22655 248404 22665 249181
rect 22707 248404 22717 249181
rect 22865 248404 22875 249181
rect 22917 248404 22927 249181
rect 23075 248404 23085 249181
rect 23127 248404 23137 249181
rect 23285 248404 23295 249181
rect 23337 248404 23347 249181
rect 23495 248404 23505 249181
rect 23547 248404 23557 249181
rect 23705 248404 23715 249181
rect 23757 248404 23767 249181
rect 23915 248404 23925 249181
rect 23967 248404 23977 249181
rect 24125 248404 24135 249181
rect 24177 248404 24187 249181
rect 24335 248404 24345 249181
rect 24387 248404 24397 249181
rect 24545 248404 24555 249181
rect 24597 248404 24607 249181
rect 24755 248404 24765 249181
rect 24807 248404 24817 249181
rect 24965 248404 24975 249181
rect 25017 248404 25027 249181
rect 25175 248404 25185 249181
rect 25227 248404 25237 249181
rect 25385 248404 25395 249181
rect 25437 248404 25447 249181
rect 25595 248404 25605 249181
rect 25647 248404 25657 249181
rect 25805 248404 25815 249181
rect 25857 248404 25867 249181
rect 26015 248404 26025 249181
rect 26067 248404 26077 249181
rect 26225 248404 26235 249181
rect 26277 248404 26287 249181
rect 26435 248404 26445 249181
rect 26487 248404 26497 249181
rect 26645 248404 26655 249181
rect 26697 248404 26707 249181
rect 26855 248404 26865 249181
rect 26907 248404 26917 249181
rect 27065 248404 27075 249181
rect 27117 248404 27127 249181
rect 27275 248404 27285 249181
rect 27331 249180 27566 249192
rect 27331 248404 27337 249180
rect 27371 248404 27566 249180
rect -4055 248392 -4009 248404
rect -3959 248392 -3913 248404
rect -3845 248392 -3799 248404
rect -3749 248392 -3703 248404
rect -3635 248392 -3589 248404
rect -3539 248392 -3493 248404
rect -3425 248392 -3379 248404
rect -3329 248392 -3283 248404
rect -3215 248392 -3169 248404
rect -3119 248392 -3073 248404
rect -3005 248392 -2959 248404
rect -2909 248392 -2863 248404
rect -2795 248392 -2749 248404
rect -2699 248392 -2653 248404
rect -2585 248392 -2539 248404
rect -2489 248392 -2443 248404
rect -2375 248392 -2329 248404
rect -2279 248392 -2233 248404
rect -2165 248392 -2119 248404
rect -2069 248392 -2023 248404
rect -1955 248392 -1909 248404
rect -1859 248392 -1813 248404
rect -1745 248392 -1699 248404
rect -1649 248392 -1603 248404
rect -1535 248392 -1489 248404
rect -1439 248392 -1393 248404
rect -1325 248392 -1279 248404
rect -1229 248392 -1183 248404
rect -1115 248392 -1069 248404
rect -1019 248392 -973 248404
rect -905 248392 -859 248404
rect -809 248392 -763 248404
rect -695 248392 -649 248404
rect -599 248392 -553 248404
rect -485 248392 -439 248404
rect -389 248392 -343 248404
rect -275 248392 -229 248404
rect -179 248392 -133 248404
rect -65 248392 -19 248404
rect 31 248392 77 248404
rect 145 248392 191 248404
rect 241 248392 287 248404
rect 355 248392 401 248404
rect 451 248392 497 248404
rect 565 248392 611 248404
rect 661 248392 707 248404
rect 775 248392 821 248404
rect 871 248392 917 248404
rect 985 248392 1031 248404
rect 1081 248392 1127 248404
rect 1195 248392 1241 248404
rect 1291 248392 1337 248404
rect 1405 248392 1451 248404
rect 1501 248392 1547 248404
rect 1615 248392 1661 248404
rect 1711 248392 1757 248404
rect 1825 248392 1871 248404
rect 1921 248392 1967 248404
rect 2035 248392 2081 248404
rect 2131 248392 2177 248404
rect 2245 248392 2291 248404
rect 2341 248392 2387 248404
rect 2455 248392 2501 248404
rect 2551 248392 2597 248404
rect 2665 248392 2711 248404
rect 2761 248392 2807 248404
rect 2875 248392 2921 248404
rect 2971 248392 3017 248404
rect 3085 248392 3131 248404
rect 3181 248392 3227 248404
rect 3295 248392 3341 248404
rect 3391 248392 3437 248404
rect 3505 248392 3551 248404
rect 3601 248392 3647 248404
rect 3715 248392 3761 248404
rect 3811 248392 3857 248404
rect 3925 248392 3971 248404
rect 4021 248392 4067 248404
rect 4135 248392 4181 248404
rect 4231 248392 4277 248404
rect 4345 248392 4391 248404
rect 4441 248392 4487 248404
rect 4555 248392 4601 248404
rect 4651 248392 4697 248404
rect 4765 248392 4811 248404
rect 4861 248392 4907 248404
rect 4975 248392 5021 248404
rect 5071 248392 5117 248404
rect 5185 248392 5231 248404
rect 5281 248392 5327 248404
rect 5395 248392 5441 248404
rect 5491 248392 5537 248404
rect 5605 248392 5651 248404
rect 5701 248392 5747 248404
rect 5815 248392 5861 248404
rect 5911 248392 5957 248404
rect 6025 248392 6071 248404
rect 6121 248392 6167 248404
rect 6235 248392 6281 248404
rect 6331 248392 6377 248404
rect 6445 248392 6491 248404
rect 6541 248392 6587 248404
rect 6655 248392 6701 248404
rect 6751 248392 6797 248404
rect 6865 248392 6911 248404
rect 6961 248392 7007 248404
rect 7075 248392 7121 248404
rect 7171 248392 7217 248404
rect 7285 248392 7331 248404
rect 7381 248392 7427 248404
rect 7495 248392 7541 248404
rect 7591 248392 7637 248404
rect 7705 248392 7751 248404
rect 7801 248392 7847 248404
rect 7915 248392 7961 248404
rect 8011 248392 8057 248404
rect 8125 248392 8171 248404
rect 8221 248392 8267 248404
rect 8335 248392 8381 248404
rect 8431 248392 8477 248404
rect 8545 248392 8591 248404
rect 8641 248392 8687 248404
rect 8755 248392 8801 248404
rect 8851 248392 8897 248404
rect 8965 248392 9011 248404
rect 9061 248392 9107 248404
rect 9175 248392 9221 248404
rect 9271 248392 9317 248404
rect 9385 248392 9431 248404
rect 9481 248392 9527 248404
rect 9595 248392 9641 248404
rect 9691 248392 9737 248404
rect 9805 248392 9851 248404
rect 9901 248392 9947 248404
rect 10015 248392 10061 248404
rect 10111 248392 10157 248404
rect 10225 248392 10271 248404
rect 10321 248392 10367 248404
rect 10435 248392 10481 248404
rect 10531 248392 10577 248404
rect 10645 248392 10691 248404
rect 10741 248392 10787 248404
rect 10855 248392 10901 248404
rect 10951 248392 10997 248404
rect 11065 248392 11111 248404
rect 11161 248392 11207 248404
rect 11275 248392 11321 248404
rect 11371 248392 11417 248404
rect 11485 248392 11531 248404
rect 11581 248392 11627 248404
rect 11695 248392 11741 248404
rect 11791 248392 11837 248404
rect 11905 248392 11951 248404
rect 12001 248392 12047 248404
rect 12115 248392 12161 248404
rect 12211 248392 12257 248404
rect 12325 248392 12371 248404
rect 12421 248392 12467 248404
rect 12535 248392 12581 248404
rect 12631 248392 12677 248404
rect 12745 248392 12791 248404
rect 12841 248392 12887 248404
rect 12955 248392 13001 248404
rect 13051 248392 13097 248404
rect 13165 248392 13211 248404
rect 13261 248392 13307 248404
rect 13375 248392 13421 248404
rect 13471 248392 13517 248404
rect 13585 248392 13631 248404
rect 13681 248392 13727 248404
rect 13795 248392 13841 248404
rect 13891 248392 13937 248404
rect 14005 248392 14051 248404
rect 14101 248392 14147 248404
rect 14215 248392 14261 248404
rect 14311 248392 14357 248404
rect 14425 248392 14471 248404
rect 14521 248392 14567 248404
rect 14635 248392 14681 248404
rect 14731 248392 14777 248404
rect 14845 248392 14891 248404
rect 14941 248392 14987 248404
rect 15055 248392 15101 248404
rect 15151 248392 15197 248404
rect 15265 248392 15311 248404
rect 15361 248392 15407 248404
rect 15475 248392 15521 248404
rect 15571 248392 15617 248404
rect 15685 248392 15731 248404
rect 15781 248392 15827 248404
rect 15895 248392 15941 248404
rect 15991 248392 16037 248404
rect 16105 248392 16151 248404
rect 16201 248392 16247 248404
rect 16315 248392 16361 248404
rect 16411 248392 16457 248404
rect 16525 248392 16571 248404
rect 16621 248392 16667 248404
rect 16735 248392 16781 248404
rect 16831 248392 16877 248404
rect 16945 248392 16991 248404
rect 17041 248392 17087 248404
rect 17155 248392 17201 248404
rect 17251 248392 17297 248404
rect 17365 248392 17411 248404
rect 17461 248392 17507 248404
rect 17575 248392 17621 248404
rect 17671 248392 17717 248404
rect 17785 248392 17831 248404
rect 17881 248392 17927 248404
rect 17995 248392 18041 248404
rect 18091 248392 18137 248404
rect 18205 248392 18251 248404
rect 18301 248392 18347 248404
rect 18415 248392 18461 248404
rect 18511 248392 18557 248404
rect 18625 248392 18671 248404
rect 18721 248392 18767 248404
rect 18835 248392 18881 248404
rect 18931 248392 18977 248404
rect 19045 248392 19091 248404
rect 19141 248392 19187 248404
rect 19255 248392 19301 248404
rect 19351 248392 19397 248404
rect 19465 248392 19511 248404
rect 19561 248392 19607 248404
rect 19675 248392 19721 248404
rect 19771 248392 19817 248404
rect 19885 248392 19931 248404
rect 19981 248392 20027 248404
rect 20095 248392 20141 248404
rect 20191 248392 20237 248404
rect 20305 248392 20351 248404
rect 20401 248392 20447 248404
rect 20515 248392 20561 248404
rect 20611 248392 20657 248404
rect 20725 248392 20771 248404
rect 20821 248392 20867 248404
rect 20935 248392 20981 248404
rect 21031 248392 21077 248404
rect 21145 248392 21191 248404
rect 21241 248392 21287 248404
rect 21355 248392 21401 248404
rect 21451 248392 21497 248404
rect 21565 248392 21611 248404
rect 21661 248392 21707 248404
rect 21775 248392 21821 248404
rect 21871 248392 21917 248404
rect 21985 248392 22031 248404
rect 22081 248392 22127 248404
rect 22195 248392 22241 248404
rect 22291 248392 22337 248404
rect 22405 248392 22451 248404
rect 22501 248392 22547 248404
rect 22615 248392 22661 248404
rect 22711 248392 22757 248404
rect 22825 248392 22871 248404
rect 22921 248392 22967 248404
rect 23035 248392 23081 248404
rect 23131 248392 23177 248404
rect 23245 248392 23291 248404
rect 23341 248392 23387 248404
rect 23455 248392 23501 248404
rect 23551 248392 23597 248404
rect 23665 248392 23711 248404
rect 23761 248392 23807 248404
rect 23875 248392 23921 248404
rect 23971 248392 24017 248404
rect 24085 248392 24131 248404
rect 24181 248392 24227 248404
rect 24295 248392 24341 248404
rect 24391 248392 24437 248404
rect 24505 248392 24551 248404
rect 24601 248392 24647 248404
rect 24715 248392 24761 248404
rect 24811 248392 24857 248404
rect 24925 248392 24971 248404
rect 25021 248392 25067 248404
rect 25135 248392 25181 248404
rect 25231 248392 25277 248404
rect 25345 248392 25391 248404
rect 25441 248392 25487 248404
rect 25555 248392 25601 248404
rect 25651 248392 25697 248404
rect 25765 248392 25811 248404
rect 25861 248392 25907 248404
rect 25975 248392 26021 248404
rect 26071 248392 26117 248404
rect 26185 248392 26231 248404
rect 26281 248392 26327 248404
rect 26395 248392 26441 248404
rect 26491 248392 26537 248404
rect 26605 248392 26651 248404
rect 26701 248392 26747 248404
rect 26815 248392 26861 248404
rect 26911 248392 26957 248404
rect 27025 248392 27071 248404
rect 27121 248392 27167 248404
rect 27235 248392 27281 248404
rect 27331 248392 27566 248404
rect -3803 248345 27335 248357
rect -5008 248203 -3791 248345
rect -3757 248203 -3371 248345
rect -3337 248203 -2951 248345
rect -2917 248203 -2531 248345
rect -2497 248203 -2111 248345
rect -2077 248203 -1691 248345
rect -1657 248203 -1271 248345
rect -1237 248203 -851 248345
rect -817 248203 -431 248345
rect -397 248203 -11 248345
rect 23 248203 409 248345
rect 443 248203 829 248345
rect 863 248203 1249 248345
rect 1283 248203 1669 248345
rect 1703 248203 2089 248345
rect 2123 248203 2509 248345
rect 2543 248203 2929 248345
rect 2963 248203 3349 248345
rect 3383 248203 3769 248345
rect 3803 248203 4189 248345
rect 4223 248203 4609 248345
rect 4643 248203 5029 248345
rect 5063 248203 5449 248345
rect 5483 248203 5869 248345
rect 5903 248203 6289 248345
rect 6323 248203 6709 248345
rect 6743 248203 7129 248345
rect 7163 248203 7549 248345
rect 7583 248203 7969 248345
rect 8003 248203 8389 248345
rect 8423 248203 8809 248345
rect 8843 248203 9229 248345
rect 9263 248203 9649 248345
rect 9683 248203 10069 248345
rect 10103 248203 10489 248345
rect 10523 248203 10909 248345
rect 10943 248203 11329 248345
rect 11363 248203 11749 248345
rect 11783 248203 12169 248345
rect 12203 248203 12589 248345
rect 12623 248203 13009 248345
rect 13043 248203 13429 248345
rect 13463 248203 13849 248345
rect 13883 248203 14269 248345
rect 14303 248203 14689 248345
rect 14723 248203 15109 248345
rect 15143 248203 15529 248345
rect 15563 248203 15949 248345
rect 15983 248203 16369 248345
rect 16403 248203 16789 248345
rect 16823 248203 17209 248345
rect 17243 248203 17629 248345
rect 17663 248203 18049 248345
rect 18083 248203 18469 248345
rect 18503 248203 18889 248345
rect 18923 248203 19309 248345
rect 19343 248203 19729 248345
rect 19763 248203 20149 248345
rect 20183 248203 20569 248345
rect 20603 248203 20989 248345
rect 21023 248203 21409 248345
rect 21443 248203 21829 248345
rect 21863 248203 22249 248345
rect 22283 248203 22669 248345
rect 22703 248203 23089 248345
rect 23123 248203 23509 248345
rect 23543 248203 23929 248345
rect 23963 248203 24349 248345
rect 24383 248203 24769 248345
rect 24803 248203 25189 248345
rect 25223 248203 25609 248345
rect 25643 248203 26029 248345
rect 26063 248203 26449 248345
rect 26483 248203 26869 248345
rect 26903 248203 27289 248345
rect 27323 248203 27335 248345
rect -5008 247309 -4142 248203
rect -3803 248191 27335 248203
rect 27377 248156 27566 248392
rect -4055 248144 -4009 248156
rect -3959 248144 -3913 248156
rect -3845 248144 -3799 248156
rect -3749 248144 -3703 248156
rect -3635 248144 -3589 248156
rect -3539 248145 -3493 248156
rect -3425 248145 -3379 248156
rect -3329 248145 -3283 248156
rect -3215 248145 -3169 248156
rect -3119 248145 -3073 248156
rect -3005 248145 -2959 248156
rect -2909 248145 -2863 248156
rect -2795 248145 -2749 248156
rect -2699 248145 -2653 248156
rect -2585 248145 -2539 248156
rect -2489 248145 -2443 248156
rect -2375 248145 -2329 248156
rect -2279 248145 -2233 248156
rect -2165 248145 -2119 248156
rect -2069 248145 -2023 248156
rect -1955 248145 -1909 248156
rect -1859 248145 -1813 248156
rect -1745 248145 -1699 248156
rect -1649 248145 -1603 248156
rect -1535 248145 -1489 248156
rect -1439 248145 -1393 248156
rect -1325 248145 -1279 248156
rect -1229 248145 -1183 248156
rect -1115 248145 -1069 248156
rect -1019 248145 -973 248156
rect -905 248145 -859 248156
rect -809 248145 -763 248156
rect -695 248145 -649 248156
rect -599 248145 -553 248156
rect -485 248145 -439 248156
rect -389 248145 -343 248156
rect -275 248145 -229 248156
rect -179 248145 -133 248156
rect -65 248145 -19 248156
rect 31 248145 77 248156
rect 145 248145 191 248156
rect 241 248145 287 248156
rect 355 248145 401 248156
rect 451 248145 497 248156
rect 565 248145 611 248156
rect 661 248145 707 248156
rect 775 248145 821 248156
rect 871 248145 917 248156
rect 985 248145 1031 248156
rect 1081 248145 1127 248156
rect 1195 248145 1241 248156
rect 1291 248145 1337 248156
rect 1405 248145 1451 248156
rect 1501 248145 1547 248156
rect 1615 248145 1661 248156
rect 1711 248145 1757 248156
rect 1825 248145 1871 248156
rect 1921 248145 1967 248156
rect 2035 248145 2081 248156
rect 2131 248145 2177 248156
rect 2245 248145 2291 248156
rect 2341 248145 2387 248156
rect 2455 248145 2501 248156
rect 2551 248145 2597 248156
rect 2665 248145 2711 248156
rect 2761 248145 2807 248156
rect 2875 248145 2921 248156
rect 2971 248145 3017 248156
rect 3085 248145 3131 248156
rect 3181 248145 3227 248156
rect 3295 248145 3341 248156
rect 3391 248145 3437 248156
rect 3505 248145 3551 248156
rect 3601 248145 3647 248156
rect 3715 248145 3761 248156
rect 3811 248145 3857 248156
rect 3925 248145 3971 248156
rect 4021 248145 4067 248156
rect 4135 248145 4181 248156
rect 4231 248145 4277 248156
rect 4345 248145 4391 248156
rect 4441 248145 4487 248156
rect 4555 248145 4601 248156
rect 4651 248145 4697 248156
rect 4765 248145 4811 248156
rect 4861 248145 4907 248156
rect 4975 248145 5021 248156
rect 5071 248145 5117 248156
rect 5185 248145 5231 248156
rect 5281 248145 5327 248156
rect 5395 248145 5441 248156
rect 5491 248145 5537 248156
rect 5605 248145 5651 248156
rect 5701 248145 5747 248156
rect 5815 248145 5861 248156
rect 5911 248145 5957 248156
rect 6025 248145 6071 248156
rect 6121 248145 6167 248156
rect 6235 248145 6281 248156
rect 6331 248145 6377 248156
rect 6445 248145 6491 248156
rect 6541 248145 6587 248156
rect 6655 248145 6701 248156
rect 6751 248145 6797 248156
rect 6865 248145 6911 248156
rect 6961 248145 7007 248156
rect 7075 248145 7121 248156
rect 7171 248145 7217 248156
rect 7285 248145 7331 248156
rect 7381 248145 7427 248156
rect 7495 248145 7541 248156
rect 7591 248145 7637 248156
rect 7705 248145 7751 248156
rect 7801 248145 7847 248156
rect 7915 248145 7961 248156
rect 8011 248145 8057 248156
rect 8125 248145 8171 248156
rect 8221 248145 8267 248156
rect 8335 248145 8381 248156
rect 8431 248145 8477 248156
rect 8545 248145 8591 248156
rect 8641 248145 8687 248156
rect 8755 248145 8801 248156
rect 8851 248145 8897 248156
rect 8965 248145 9011 248156
rect 9061 248145 9107 248156
rect 9175 248145 9221 248156
rect 9271 248145 9317 248156
rect 9385 248145 9431 248156
rect 9481 248145 9527 248156
rect 9595 248145 9641 248156
rect 9691 248145 9737 248156
rect 9805 248145 9851 248156
rect 9901 248145 9947 248156
rect 10015 248145 10061 248156
rect 10111 248145 10157 248156
rect 10225 248145 10271 248156
rect 10321 248145 10367 248156
rect 10435 248145 10481 248156
rect 10531 248145 10577 248156
rect 10645 248145 10691 248156
rect 10741 248145 10787 248156
rect 10855 248145 10901 248156
rect 10951 248145 10997 248156
rect 11065 248145 11111 248156
rect 11161 248145 11207 248156
rect 11275 248145 11321 248156
rect 11371 248145 11417 248156
rect 11485 248145 11531 248156
rect 11581 248145 11627 248156
rect 11695 248145 11741 248156
rect 11791 248145 11837 248156
rect 11905 248145 11951 248156
rect 12001 248145 12047 248156
rect 12115 248145 12161 248156
rect 12211 248145 12257 248156
rect 12325 248145 12371 248156
rect 12421 248145 12467 248156
rect 12535 248145 12581 248156
rect 12631 248145 12677 248156
rect 12745 248145 12791 248156
rect 12841 248145 12887 248156
rect 12955 248145 13001 248156
rect 13051 248145 13097 248156
rect 13165 248145 13211 248156
rect 13261 248145 13307 248156
rect 13375 248145 13421 248156
rect 13471 248145 13517 248156
rect 13585 248145 13631 248156
rect 13681 248145 13727 248156
rect 13795 248145 13841 248156
rect 13891 248145 13937 248156
rect 14005 248145 14051 248156
rect 14101 248145 14147 248156
rect 14215 248145 14261 248156
rect 14311 248145 14357 248156
rect 14425 248145 14471 248156
rect 14521 248145 14567 248156
rect 14635 248145 14681 248156
rect 14731 248145 14777 248156
rect 14845 248145 14891 248156
rect 14941 248145 14987 248156
rect 15055 248145 15101 248156
rect 15151 248145 15197 248156
rect 15265 248145 15311 248156
rect 15361 248145 15407 248156
rect 15475 248145 15521 248156
rect 15571 248145 15617 248156
rect 15685 248145 15731 248156
rect 15781 248145 15827 248156
rect 15895 248145 15941 248156
rect 15991 248145 16037 248156
rect 16105 248145 16151 248156
rect 16201 248145 16247 248156
rect 16315 248145 16361 248156
rect 16411 248145 16457 248156
rect 16525 248145 16571 248156
rect 16621 248145 16667 248156
rect 16735 248145 16781 248156
rect 16831 248145 16877 248156
rect 16945 248145 16991 248156
rect 17041 248145 17087 248156
rect 17155 248145 17201 248156
rect 17251 248145 17297 248156
rect 17365 248145 17411 248156
rect 17461 248145 17507 248156
rect 17575 248145 17621 248156
rect 17671 248145 17717 248156
rect 17785 248145 17831 248156
rect 17881 248145 17927 248156
rect 17995 248145 18041 248156
rect 18091 248145 18137 248156
rect 18205 248145 18251 248156
rect 18301 248145 18347 248156
rect 18415 248145 18461 248156
rect 18511 248145 18557 248156
rect 18625 248145 18671 248156
rect 18721 248145 18767 248156
rect 18835 248145 18881 248156
rect 18931 248145 18977 248156
rect 19045 248145 19091 248156
rect 19141 248145 19187 248156
rect 19255 248145 19301 248156
rect 19351 248145 19397 248156
rect 19465 248145 19511 248156
rect 19561 248145 19607 248156
rect 19675 248145 19721 248156
rect 19771 248145 19817 248156
rect 19885 248145 19931 248156
rect 19981 248145 20027 248156
rect 20095 248145 20141 248156
rect 20191 248145 20237 248156
rect 20305 248145 20351 248156
rect 20401 248145 20447 248156
rect 20515 248145 20561 248156
rect 20611 248145 20657 248156
rect 20725 248145 20771 248156
rect 20821 248145 20867 248156
rect 20935 248145 20981 248156
rect 21031 248145 21077 248156
rect 21145 248145 21191 248156
rect 21241 248145 21287 248156
rect 21355 248145 21401 248156
rect 21451 248145 21497 248156
rect 21565 248145 21611 248156
rect 21661 248145 21707 248156
rect 21775 248145 21821 248156
rect 21871 248145 21917 248156
rect 21985 248145 22031 248156
rect 22081 248145 22127 248156
rect 22195 248145 22241 248156
rect 22291 248145 22337 248156
rect 22405 248145 22451 248156
rect 22501 248145 22547 248156
rect 22615 248145 22661 248156
rect 22711 248145 22757 248156
rect 22825 248145 22871 248156
rect 22921 248145 22967 248156
rect 23035 248145 23081 248156
rect 23131 248145 23177 248156
rect 23245 248145 23291 248156
rect 23341 248145 23387 248156
rect 23455 248145 23501 248156
rect 23551 248145 23597 248156
rect 23665 248145 23711 248156
rect 23761 248145 23807 248156
rect 23875 248145 23921 248156
rect 23971 248145 24017 248156
rect 24085 248145 24131 248156
rect 24181 248145 24227 248156
rect 24295 248145 24341 248156
rect 24391 248145 24437 248156
rect 24505 248145 24551 248156
rect 24601 248145 24647 248156
rect 24715 248145 24761 248156
rect 24811 248145 24857 248156
rect 24925 248145 24971 248156
rect 25021 248145 25067 248156
rect 25135 248145 25181 248156
rect 25231 248145 25277 248156
rect 25345 248145 25391 248156
rect 25441 248145 25487 248156
rect 25555 248145 25601 248156
rect 25651 248145 25697 248156
rect 25765 248145 25811 248156
rect 25861 248145 25907 248156
rect 25975 248145 26021 248156
rect 26071 248145 26117 248156
rect 26185 248145 26231 248156
rect 26281 248145 26327 248156
rect 26395 248145 26441 248156
rect 26491 248145 26537 248156
rect 26605 248145 26651 248156
rect 26701 248145 26747 248156
rect 26815 248145 26861 248156
rect 26911 248145 26957 248156
rect 27025 248145 27071 248156
rect 27121 248145 27167 248156
rect 27235 248145 27281 248156
rect -4085 247368 -4075 248144
rect -4015 247368 -4005 248144
rect -3963 247368 -3953 248144
rect -3805 247368 -3795 248144
rect -3753 247368 -3743 248144
rect -3595 247368 -3585 248144
rect -3543 247368 -3533 248145
rect -3385 247368 -3375 248145
rect -3333 247368 -3323 248145
rect -3175 247368 -3165 248145
rect -3123 247368 -3113 248145
rect -2965 247368 -2955 248145
rect -2913 247368 -2903 248145
rect -2755 247368 -2745 248145
rect -2703 247368 -2693 248145
rect -2545 247368 -2535 248145
rect -2493 247368 -2483 248145
rect -2335 247368 -2325 248145
rect -2283 247368 -2273 248145
rect -2125 247368 -2115 248145
rect -2073 247368 -2063 248145
rect -1915 247368 -1905 248145
rect -1863 247368 -1853 248145
rect -1705 247368 -1695 248145
rect -1653 247368 -1643 248145
rect -1495 247368 -1485 248145
rect -1443 247368 -1433 248145
rect -1285 247368 -1275 248145
rect -1233 247368 -1223 248145
rect -1075 247368 -1065 248145
rect -1023 247368 -1013 248145
rect -865 247368 -855 248145
rect -813 247368 -803 248145
rect -655 247368 -645 248145
rect -603 247368 -593 248145
rect -445 247368 -435 248145
rect -393 247368 -383 248145
rect -235 247368 -225 248145
rect -183 247368 -173 248145
rect -25 247368 -15 248145
rect 27 247368 37 248145
rect 185 247368 195 248145
rect 237 247368 247 248145
rect 395 247368 405 248145
rect 447 247368 457 248145
rect 605 247368 615 248145
rect 657 247368 667 248145
rect 815 247368 825 248145
rect 867 247368 877 248145
rect 1025 247368 1035 248145
rect 1077 247368 1087 248145
rect 1235 247368 1245 248145
rect 1287 247368 1297 248145
rect 1445 247368 1455 248145
rect 1497 247368 1507 248145
rect 1655 247368 1665 248145
rect 1707 247368 1717 248145
rect 1865 247368 1875 248145
rect 1917 247368 1927 248145
rect 2075 247368 2085 248145
rect 2127 247368 2137 248145
rect 2285 247368 2295 248145
rect 2337 247368 2347 248145
rect 2495 247368 2505 248145
rect 2547 247368 2557 248145
rect 2705 247368 2715 248145
rect 2757 247368 2767 248145
rect 2915 247368 2925 248145
rect 2967 247368 2977 248145
rect 3125 247368 3135 248145
rect 3177 247368 3187 248145
rect 3335 247368 3345 248145
rect 3387 247368 3397 248145
rect 3545 247368 3555 248145
rect 3597 247368 3607 248145
rect 3755 247368 3765 248145
rect 3807 247368 3817 248145
rect 3965 247368 3975 248145
rect 4017 247368 4027 248145
rect 4175 247368 4185 248145
rect 4227 247368 4237 248145
rect 4385 247368 4395 248145
rect 4437 247368 4447 248145
rect 4595 247368 4605 248145
rect 4647 247368 4657 248145
rect 4805 247368 4815 248145
rect 4857 247368 4867 248145
rect 5015 247368 5025 248145
rect 5067 247368 5077 248145
rect 5225 247368 5235 248145
rect 5277 247368 5287 248145
rect 5435 247368 5445 248145
rect 5487 247368 5497 248145
rect 5645 247368 5655 248145
rect 5697 247368 5707 248145
rect 5855 247368 5865 248145
rect 5907 247368 5917 248145
rect 6065 247368 6075 248145
rect 6117 247368 6127 248145
rect 6275 247368 6285 248145
rect 6327 247368 6337 248145
rect 6485 247368 6495 248145
rect 6537 247368 6547 248145
rect 6695 247368 6705 248145
rect 6747 247368 6757 248145
rect 6905 247368 6915 248145
rect 6957 247368 6967 248145
rect 7115 247368 7125 248145
rect 7167 247368 7177 248145
rect 7325 247368 7335 248145
rect 7377 247368 7387 248145
rect 7535 247368 7545 248145
rect 7587 247368 7597 248145
rect 7745 247368 7755 248145
rect 7797 247368 7807 248145
rect 7955 247368 7965 248145
rect 8007 247368 8017 248145
rect 8165 247368 8175 248145
rect 8217 247368 8227 248145
rect 8375 247368 8385 248145
rect 8427 247368 8437 248145
rect 8585 247368 8595 248145
rect 8637 247368 8647 248145
rect 8795 247368 8805 248145
rect 8847 247368 8857 248145
rect 9005 247368 9015 248145
rect 9057 247368 9067 248145
rect 9215 247368 9225 248145
rect 9267 247368 9277 248145
rect 9425 247368 9435 248145
rect 9477 247368 9487 248145
rect 9635 247368 9645 248145
rect 9687 247368 9697 248145
rect 9845 247368 9855 248145
rect 9897 247368 9907 248145
rect 10055 247368 10065 248145
rect 10107 247368 10117 248145
rect 10265 247368 10275 248145
rect 10317 247368 10327 248145
rect 10475 247368 10485 248145
rect 10527 247368 10537 248145
rect 10685 247368 10695 248145
rect 10737 247368 10747 248145
rect 10895 247368 10905 248145
rect 10947 247368 10957 248145
rect 11105 247368 11115 248145
rect 11157 247368 11167 248145
rect 11315 247368 11325 248145
rect 11367 247368 11377 248145
rect 11525 247368 11535 248145
rect 11577 247368 11587 248145
rect 11735 247368 11745 248145
rect 11787 247368 11797 248145
rect 11945 247368 11955 248145
rect 11997 247368 12007 248145
rect 12155 247368 12165 248145
rect 12207 247368 12217 248145
rect 12365 247368 12375 248145
rect 12417 247368 12427 248145
rect 12575 247368 12585 248145
rect 12627 247368 12637 248145
rect 12785 247368 12795 248145
rect 12837 247368 12847 248145
rect 12995 247368 13005 248145
rect 13047 247368 13057 248145
rect 13205 247368 13215 248145
rect 13257 247368 13267 248145
rect 13415 247368 13425 248145
rect 13467 247368 13477 248145
rect 13625 247368 13635 248145
rect 13677 247368 13687 248145
rect 13835 247368 13845 248145
rect 13887 247368 13897 248145
rect 14045 247368 14055 248145
rect 14097 247368 14107 248145
rect 14255 247368 14265 248145
rect 14307 247368 14317 248145
rect 14465 247368 14475 248145
rect 14517 247368 14527 248145
rect 14675 247368 14685 248145
rect 14727 247368 14737 248145
rect 14885 247368 14895 248145
rect 14937 247368 14947 248145
rect 15095 247368 15105 248145
rect 15147 247368 15157 248145
rect 15305 247368 15315 248145
rect 15357 247368 15367 248145
rect 15515 247368 15525 248145
rect 15567 247368 15577 248145
rect 15725 247368 15735 248145
rect 15777 247368 15787 248145
rect 15935 247368 15945 248145
rect 15987 247368 15997 248145
rect 16145 247368 16155 248145
rect 16197 247368 16207 248145
rect 16355 247368 16365 248145
rect 16407 247368 16417 248145
rect 16565 247368 16575 248145
rect 16617 247368 16627 248145
rect 16775 247368 16785 248145
rect 16827 247368 16837 248145
rect 16985 247368 16995 248145
rect 17037 247368 17047 248145
rect 17195 247368 17205 248145
rect 17247 247368 17257 248145
rect 17405 247368 17415 248145
rect 17457 247368 17467 248145
rect 17615 247368 17625 248145
rect 17667 247368 17677 248145
rect 17825 247368 17835 248145
rect 17877 247368 17887 248145
rect 18035 247368 18045 248145
rect 18087 247368 18097 248145
rect 18245 247368 18255 248145
rect 18297 247368 18307 248145
rect 18455 247368 18465 248145
rect 18507 247368 18517 248145
rect 18665 247368 18675 248145
rect 18717 247368 18727 248145
rect 18875 247368 18885 248145
rect 18927 247368 18937 248145
rect 19085 247368 19095 248145
rect 19137 247368 19147 248145
rect 19295 247368 19305 248145
rect 19347 247368 19357 248145
rect 19505 247368 19515 248145
rect 19557 247368 19567 248145
rect 19715 247368 19725 248145
rect 19767 247368 19777 248145
rect 19925 247368 19935 248145
rect 19977 247368 19987 248145
rect 20135 247368 20145 248145
rect 20187 247368 20197 248145
rect 20345 247368 20355 248145
rect 20397 247368 20407 248145
rect 20555 247368 20565 248145
rect 20607 247368 20617 248145
rect 20765 247368 20775 248145
rect 20817 247368 20827 248145
rect 20975 247368 20985 248145
rect 21027 247368 21037 248145
rect 21185 247368 21195 248145
rect 21237 247368 21247 248145
rect 21395 247368 21405 248145
rect 21447 247368 21457 248145
rect 21605 247368 21615 248145
rect 21657 247368 21667 248145
rect 21815 247368 21825 248145
rect 21867 247368 21877 248145
rect 22025 247368 22035 248145
rect 22077 247368 22087 248145
rect 22235 247368 22245 248145
rect 22287 247368 22297 248145
rect 22445 247368 22455 248145
rect 22497 247368 22507 248145
rect 22655 247368 22665 248145
rect 22707 247368 22717 248145
rect 22865 247368 22875 248145
rect 22917 247368 22927 248145
rect 23075 247368 23085 248145
rect 23127 247368 23137 248145
rect 23285 247368 23295 248145
rect 23337 247368 23347 248145
rect 23495 247368 23505 248145
rect 23547 247368 23557 248145
rect 23705 247368 23715 248145
rect 23757 247368 23767 248145
rect 23915 247368 23925 248145
rect 23967 247368 23977 248145
rect 24125 247368 24135 248145
rect 24177 247368 24187 248145
rect 24335 247368 24345 248145
rect 24387 247368 24397 248145
rect 24545 247368 24555 248145
rect 24597 247368 24607 248145
rect 24755 247368 24765 248145
rect 24807 247368 24817 248145
rect 24965 247368 24975 248145
rect 25017 247368 25027 248145
rect 25175 247368 25185 248145
rect 25227 247368 25237 248145
rect 25385 247368 25395 248145
rect 25437 247368 25447 248145
rect 25595 247368 25605 248145
rect 25647 247368 25657 248145
rect 25805 247368 25815 248145
rect 25857 247368 25867 248145
rect 26015 247368 26025 248145
rect 26067 247368 26077 248145
rect 26225 247368 26235 248145
rect 26277 247368 26287 248145
rect 26435 247368 26445 248145
rect 26487 247368 26497 248145
rect 26645 247368 26655 248145
rect 26697 247368 26707 248145
rect 26855 247368 26865 248145
rect 26907 247368 26917 248145
rect 27065 247368 27075 248145
rect 27117 247368 27127 248145
rect 27275 247368 27285 248145
rect 27331 248144 27566 248156
rect 27331 247368 27337 248144
rect 27371 247368 27566 248144
rect -4055 247356 -4009 247368
rect -3959 247356 -3913 247368
rect -3845 247356 -3799 247368
rect -3749 247356 -3703 247368
rect -3635 247356 -3589 247368
rect -3539 247356 -3493 247368
rect -3425 247356 -3379 247368
rect -3329 247356 -3283 247368
rect -3215 247356 -3169 247368
rect -3119 247356 -3073 247368
rect -3005 247356 -2959 247368
rect -2909 247356 -2863 247368
rect -2795 247356 -2749 247368
rect -2699 247356 -2653 247368
rect -2585 247356 -2539 247368
rect -2489 247356 -2443 247368
rect -2375 247356 -2329 247368
rect -2279 247356 -2233 247368
rect -2165 247356 -2119 247368
rect -2069 247356 -2023 247368
rect -1955 247356 -1909 247368
rect -1859 247356 -1813 247368
rect -1745 247356 -1699 247368
rect -1649 247356 -1603 247368
rect -1535 247356 -1489 247368
rect -1439 247356 -1393 247368
rect -1325 247356 -1279 247368
rect -1229 247356 -1183 247368
rect -1115 247356 -1069 247368
rect -1019 247356 -973 247368
rect -905 247356 -859 247368
rect -809 247356 -763 247368
rect -695 247356 -649 247368
rect -599 247356 -553 247368
rect -485 247356 -439 247368
rect -389 247356 -343 247368
rect -275 247356 -229 247368
rect -179 247356 -133 247368
rect -65 247356 -19 247368
rect 31 247356 77 247368
rect 145 247356 191 247368
rect 241 247356 287 247368
rect 355 247356 401 247368
rect 451 247356 497 247368
rect 565 247356 611 247368
rect 661 247356 707 247368
rect 775 247356 821 247368
rect 871 247356 917 247368
rect 985 247356 1031 247368
rect 1081 247356 1127 247368
rect 1195 247356 1241 247368
rect 1291 247356 1337 247368
rect 1405 247356 1451 247368
rect 1501 247356 1547 247368
rect 1615 247356 1661 247368
rect 1711 247356 1757 247368
rect 1825 247356 1871 247368
rect 1921 247356 1967 247368
rect 2035 247356 2081 247368
rect 2131 247356 2177 247368
rect 2245 247356 2291 247368
rect 2341 247356 2387 247368
rect 2455 247356 2501 247368
rect 2551 247356 2597 247368
rect 2665 247356 2711 247368
rect 2761 247356 2807 247368
rect 2875 247356 2921 247368
rect 2971 247356 3017 247368
rect 3085 247356 3131 247368
rect 3181 247356 3227 247368
rect 3295 247356 3341 247368
rect 3391 247356 3437 247368
rect 3505 247356 3551 247368
rect 3601 247356 3647 247368
rect 3715 247356 3761 247368
rect 3811 247356 3857 247368
rect 3925 247356 3971 247368
rect 4021 247356 4067 247368
rect 4135 247356 4181 247368
rect 4231 247356 4277 247368
rect 4345 247356 4391 247368
rect 4441 247356 4487 247368
rect 4555 247356 4601 247368
rect 4651 247356 4697 247368
rect 4765 247356 4811 247368
rect 4861 247356 4907 247368
rect 4975 247356 5021 247368
rect 5071 247356 5117 247368
rect 5185 247356 5231 247368
rect 5281 247356 5327 247368
rect 5395 247356 5441 247368
rect 5491 247356 5537 247368
rect 5605 247356 5651 247368
rect 5701 247356 5747 247368
rect 5815 247356 5861 247368
rect 5911 247356 5957 247368
rect 6025 247356 6071 247368
rect 6121 247356 6167 247368
rect 6235 247356 6281 247368
rect 6331 247356 6377 247368
rect 6445 247356 6491 247368
rect 6541 247356 6587 247368
rect 6655 247356 6701 247368
rect 6751 247356 6797 247368
rect 6865 247356 6911 247368
rect 6961 247356 7007 247368
rect 7075 247356 7121 247368
rect 7171 247356 7217 247368
rect 7285 247356 7331 247368
rect 7381 247356 7427 247368
rect 7495 247356 7541 247368
rect 7591 247356 7637 247368
rect 7705 247356 7751 247368
rect 7801 247356 7847 247368
rect 7915 247356 7961 247368
rect 8011 247356 8057 247368
rect 8125 247356 8171 247368
rect 8221 247356 8267 247368
rect 8335 247356 8381 247368
rect 8431 247356 8477 247368
rect 8545 247356 8591 247368
rect 8641 247356 8687 247368
rect 8755 247356 8801 247368
rect 8851 247356 8897 247368
rect 8965 247356 9011 247368
rect 9061 247356 9107 247368
rect 9175 247356 9221 247368
rect 9271 247356 9317 247368
rect 9385 247356 9431 247368
rect 9481 247356 9527 247368
rect 9595 247356 9641 247368
rect 9691 247356 9737 247368
rect 9805 247356 9851 247368
rect 9901 247356 9947 247368
rect 10015 247356 10061 247368
rect 10111 247356 10157 247368
rect 10225 247356 10271 247368
rect 10321 247356 10367 247368
rect 10435 247356 10481 247368
rect 10531 247356 10577 247368
rect 10645 247356 10691 247368
rect 10741 247356 10787 247368
rect 10855 247356 10901 247368
rect 10951 247356 10997 247368
rect 11065 247356 11111 247368
rect 11161 247356 11207 247368
rect 11275 247356 11321 247368
rect 11371 247356 11417 247368
rect 11485 247356 11531 247368
rect 11581 247356 11627 247368
rect 11695 247356 11741 247368
rect 11791 247356 11837 247368
rect 11905 247356 11951 247368
rect 12001 247356 12047 247368
rect 12115 247356 12161 247368
rect 12211 247356 12257 247368
rect 12325 247356 12371 247368
rect 12421 247356 12467 247368
rect 12535 247356 12581 247368
rect 12631 247356 12677 247368
rect 12745 247356 12791 247368
rect 12841 247356 12887 247368
rect 12955 247356 13001 247368
rect 13051 247356 13097 247368
rect 13165 247356 13211 247368
rect 13261 247356 13307 247368
rect 13375 247356 13421 247368
rect 13471 247356 13517 247368
rect 13585 247356 13631 247368
rect 13681 247356 13727 247368
rect 13795 247356 13841 247368
rect 13891 247356 13937 247368
rect 14005 247356 14051 247368
rect 14101 247356 14147 247368
rect 14215 247356 14261 247368
rect 14311 247356 14357 247368
rect 14425 247356 14471 247368
rect 14521 247356 14567 247368
rect 14635 247356 14681 247368
rect 14731 247356 14777 247368
rect 14845 247356 14891 247368
rect 14941 247356 14987 247368
rect 15055 247356 15101 247368
rect 15151 247356 15197 247368
rect 15265 247356 15311 247368
rect 15361 247356 15407 247368
rect 15475 247356 15521 247368
rect 15571 247356 15617 247368
rect 15685 247356 15731 247368
rect 15781 247356 15827 247368
rect 15895 247356 15941 247368
rect 15991 247356 16037 247368
rect 16105 247356 16151 247368
rect 16201 247356 16247 247368
rect 16315 247356 16361 247368
rect 16411 247356 16457 247368
rect 16525 247356 16571 247368
rect 16621 247356 16667 247368
rect 16735 247356 16781 247368
rect 16831 247356 16877 247368
rect 16945 247356 16991 247368
rect 17041 247356 17087 247368
rect 17155 247356 17201 247368
rect 17251 247356 17297 247368
rect 17365 247356 17411 247368
rect 17461 247356 17507 247368
rect 17575 247356 17621 247368
rect 17671 247356 17717 247368
rect 17785 247356 17831 247368
rect 17881 247356 17927 247368
rect 17995 247356 18041 247368
rect 18091 247356 18137 247368
rect 18205 247356 18251 247368
rect 18301 247356 18347 247368
rect 18415 247356 18461 247368
rect 18511 247356 18557 247368
rect 18625 247356 18671 247368
rect 18721 247356 18767 247368
rect 18835 247356 18881 247368
rect 18931 247356 18977 247368
rect 19045 247356 19091 247368
rect 19141 247356 19187 247368
rect 19255 247356 19301 247368
rect 19351 247356 19397 247368
rect 19465 247356 19511 247368
rect 19561 247356 19607 247368
rect 19675 247356 19721 247368
rect 19771 247356 19817 247368
rect 19885 247356 19931 247368
rect 19981 247356 20027 247368
rect 20095 247356 20141 247368
rect 20191 247356 20237 247368
rect 20305 247356 20351 247368
rect 20401 247356 20447 247368
rect 20515 247356 20561 247368
rect 20611 247356 20657 247368
rect 20725 247356 20771 247368
rect 20821 247356 20867 247368
rect 20935 247356 20981 247368
rect 21031 247356 21077 247368
rect 21145 247356 21191 247368
rect 21241 247356 21287 247368
rect 21355 247356 21401 247368
rect 21451 247356 21497 247368
rect 21565 247356 21611 247368
rect 21661 247356 21707 247368
rect 21775 247356 21821 247368
rect 21871 247356 21917 247368
rect 21985 247356 22031 247368
rect 22081 247356 22127 247368
rect 22195 247356 22241 247368
rect 22291 247356 22337 247368
rect 22405 247356 22451 247368
rect 22501 247356 22547 247368
rect 22615 247356 22661 247368
rect 22711 247356 22757 247368
rect 22825 247356 22871 247368
rect 22921 247356 22967 247368
rect 23035 247356 23081 247368
rect 23131 247356 23177 247368
rect 23245 247356 23291 247368
rect 23341 247356 23387 247368
rect 23455 247356 23501 247368
rect 23551 247356 23597 247368
rect 23665 247356 23711 247368
rect 23761 247356 23807 247368
rect 23875 247356 23921 247368
rect 23971 247356 24017 247368
rect 24085 247356 24131 247368
rect 24181 247356 24227 247368
rect 24295 247356 24341 247368
rect 24391 247356 24437 247368
rect 24505 247356 24551 247368
rect 24601 247356 24647 247368
rect 24715 247356 24761 247368
rect 24811 247356 24857 247368
rect 24925 247356 24971 247368
rect 25021 247356 25067 247368
rect 25135 247356 25181 247368
rect 25231 247356 25277 247368
rect 25345 247356 25391 247368
rect 25441 247356 25487 247368
rect 25555 247356 25601 247368
rect 25651 247356 25697 247368
rect 25765 247356 25811 247368
rect 25861 247356 25907 247368
rect 25975 247356 26021 247368
rect 26071 247356 26117 247368
rect 26185 247356 26231 247368
rect 26281 247356 26327 247368
rect 26395 247356 26441 247368
rect 26491 247356 26537 247368
rect 26605 247356 26651 247368
rect 26701 247356 26747 247368
rect 26815 247356 26861 247368
rect 26911 247356 26957 247368
rect 27025 247356 27071 247368
rect 27121 247356 27167 247368
rect 27235 247356 27281 247368
rect 27331 247356 27566 247368
rect -4013 247309 27125 247321
rect -5008 247167 -4001 247309
rect -3967 247167 -3581 247309
rect -3547 247167 -3161 247309
rect -3127 247167 -2741 247309
rect -2707 247167 -2321 247309
rect -2287 247167 -1901 247309
rect -1867 247167 -1481 247309
rect -1447 247167 -1061 247309
rect -1027 247167 -641 247309
rect -607 247167 -221 247309
rect -187 247167 199 247309
rect 233 247167 619 247309
rect 653 247167 1039 247309
rect 1073 247167 1459 247309
rect 1493 247167 1879 247309
rect 1913 247167 2299 247309
rect 2333 247167 2719 247309
rect 2753 247167 3139 247309
rect 3173 247167 3559 247309
rect 3593 247167 3979 247309
rect 4013 247167 4399 247309
rect 4433 247167 4819 247309
rect 4853 247167 5239 247309
rect 5273 247167 5659 247309
rect 5693 247167 6079 247309
rect 6113 247167 6499 247309
rect 6533 247167 6919 247309
rect 6953 247167 7339 247309
rect 7373 247167 7759 247309
rect 7793 247167 8179 247309
rect 8213 247167 8599 247309
rect 8633 247167 9019 247309
rect 9053 247167 9439 247309
rect 9473 247167 9859 247309
rect 9893 247167 10279 247309
rect 10313 247167 10699 247309
rect 10733 247167 11119 247309
rect 11153 247167 11539 247309
rect 11573 247167 11959 247309
rect 11993 247167 12379 247309
rect 12413 247167 12799 247309
rect 12833 247167 13219 247309
rect 13253 247167 13639 247309
rect 13673 247167 14059 247309
rect 14093 247167 14479 247309
rect 14513 247167 14899 247309
rect 14933 247167 15319 247309
rect 15353 247167 15739 247309
rect 15773 247167 16159 247309
rect 16193 247167 16579 247309
rect 16613 247167 16999 247309
rect 17033 247167 17419 247309
rect 17453 247167 17839 247309
rect 17873 247167 18259 247309
rect 18293 247167 18679 247309
rect 18713 247167 19099 247309
rect 19133 247167 19519 247309
rect 19553 247167 19939 247309
rect 19973 247167 20359 247309
rect 20393 247167 20779 247309
rect 20813 247167 21199 247309
rect 21233 247167 21619 247309
rect 21653 247167 22039 247309
rect 22073 247167 22459 247309
rect 22493 247167 22879 247309
rect 22913 247167 23299 247309
rect 23333 247167 23719 247309
rect 23753 247167 24139 247309
rect 24173 247167 24559 247309
rect 24593 247167 24979 247309
rect 25013 247167 25399 247309
rect 25433 247167 25819 247309
rect 25853 247167 26239 247309
rect 26273 247167 26659 247309
rect 26693 247167 27079 247309
rect 27113 247167 27125 247309
rect -5008 246273 -4142 247167
rect -4013 247155 27125 247167
rect 27377 247120 27566 247356
rect -4055 247108 -4009 247120
rect -3959 247108 -3913 247120
rect -3845 247108 -3799 247120
rect -3749 247108 -3703 247120
rect -3635 247108 -3589 247120
rect -3539 247109 -3493 247120
rect -3425 247109 -3379 247120
rect -3329 247109 -3283 247120
rect -3215 247109 -3169 247120
rect -3119 247109 -3073 247120
rect -3005 247109 -2959 247120
rect -2909 247109 -2863 247120
rect -2795 247109 -2749 247120
rect -2699 247109 -2653 247120
rect -2585 247109 -2539 247120
rect -2489 247109 -2443 247120
rect -2375 247109 -2329 247120
rect -2279 247109 -2233 247120
rect -2165 247109 -2119 247120
rect -2069 247109 -2023 247120
rect -1955 247109 -1909 247120
rect -1859 247109 -1813 247120
rect -1745 247109 -1699 247120
rect -1649 247109 -1603 247120
rect -1535 247109 -1489 247120
rect -1439 247109 -1393 247120
rect -1325 247109 -1279 247120
rect -1229 247109 -1183 247120
rect -1115 247109 -1069 247120
rect -1019 247109 -973 247120
rect -905 247109 -859 247120
rect -809 247109 -763 247120
rect -695 247109 -649 247120
rect -599 247109 -553 247120
rect -485 247109 -439 247120
rect -389 247109 -343 247120
rect -275 247109 -229 247120
rect -179 247109 -133 247120
rect -65 247109 -19 247120
rect 31 247109 77 247120
rect 145 247109 191 247120
rect 241 247109 287 247120
rect 355 247109 401 247120
rect 451 247109 497 247120
rect 565 247109 611 247120
rect 661 247109 707 247120
rect 775 247109 821 247120
rect 871 247109 917 247120
rect 985 247109 1031 247120
rect 1081 247109 1127 247120
rect 1195 247109 1241 247120
rect 1291 247109 1337 247120
rect 1405 247109 1451 247120
rect 1501 247109 1547 247120
rect 1615 247109 1661 247120
rect 1711 247109 1757 247120
rect 1825 247109 1871 247120
rect 1921 247109 1967 247120
rect 2035 247109 2081 247120
rect 2131 247109 2177 247120
rect 2245 247109 2291 247120
rect 2341 247109 2387 247120
rect 2455 247109 2501 247120
rect 2551 247109 2597 247120
rect 2665 247109 2711 247120
rect 2761 247109 2807 247120
rect 2875 247109 2921 247120
rect 2971 247109 3017 247120
rect 3085 247109 3131 247120
rect 3181 247109 3227 247120
rect 3295 247109 3341 247120
rect 3391 247109 3437 247120
rect 3505 247109 3551 247120
rect 3601 247109 3647 247120
rect 3715 247109 3761 247120
rect 3811 247109 3857 247120
rect 3925 247109 3971 247120
rect 4021 247109 4067 247120
rect 4135 247109 4181 247120
rect 4231 247109 4277 247120
rect 4345 247109 4391 247120
rect 4441 247109 4487 247120
rect 4555 247109 4601 247120
rect 4651 247109 4697 247120
rect 4765 247109 4811 247120
rect 4861 247109 4907 247120
rect 4975 247109 5021 247120
rect 5071 247109 5117 247120
rect 5185 247109 5231 247120
rect 5281 247109 5327 247120
rect 5395 247109 5441 247120
rect 5491 247109 5537 247120
rect 5605 247109 5651 247120
rect 5701 247109 5747 247120
rect 5815 247109 5861 247120
rect 5911 247109 5957 247120
rect 6025 247109 6071 247120
rect 6121 247109 6167 247120
rect 6235 247109 6281 247120
rect 6331 247109 6377 247120
rect 6445 247109 6491 247120
rect 6541 247109 6587 247120
rect 6655 247109 6701 247120
rect 6751 247109 6797 247120
rect 6865 247109 6911 247120
rect 6961 247109 7007 247120
rect 7075 247109 7121 247120
rect 7171 247109 7217 247120
rect 7285 247109 7331 247120
rect 7381 247109 7427 247120
rect 7495 247109 7541 247120
rect 7591 247109 7637 247120
rect 7705 247109 7751 247120
rect 7801 247109 7847 247120
rect 7915 247109 7961 247120
rect 8011 247109 8057 247120
rect 8125 247109 8171 247120
rect 8221 247109 8267 247120
rect 8335 247109 8381 247120
rect 8431 247109 8477 247120
rect 8545 247109 8591 247120
rect 8641 247109 8687 247120
rect 8755 247109 8801 247120
rect 8851 247109 8897 247120
rect 8965 247109 9011 247120
rect 9061 247109 9107 247120
rect 9175 247109 9221 247120
rect 9271 247109 9317 247120
rect 9385 247109 9431 247120
rect 9481 247109 9527 247120
rect 9595 247109 9641 247120
rect 9691 247109 9737 247120
rect 9805 247109 9851 247120
rect 9901 247109 9947 247120
rect 10015 247109 10061 247120
rect 10111 247109 10157 247120
rect 10225 247109 10271 247120
rect 10321 247109 10367 247120
rect 10435 247109 10481 247120
rect 10531 247109 10577 247120
rect 10645 247109 10691 247120
rect 10741 247109 10787 247120
rect 10855 247109 10901 247120
rect 10951 247109 10997 247120
rect 11065 247109 11111 247120
rect 11161 247109 11207 247120
rect 11275 247109 11321 247120
rect 11371 247109 11417 247120
rect 11485 247109 11531 247120
rect 11581 247109 11627 247120
rect 11695 247109 11741 247120
rect 11791 247109 11837 247120
rect 11905 247109 11951 247120
rect 12001 247109 12047 247120
rect 12115 247109 12161 247120
rect 12211 247109 12257 247120
rect 12325 247109 12371 247120
rect 12421 247109 12467 247120
rect 12535 247109 12581 247120
rect 12631 247109 12677 247120
rect 12745 247109 12791 247120
rect 12841 247109 12887 247120
rect 12955 247109 13001 247120
rect 13051 247109 13097 247120
rect 13165 247109 13211 247120
rect 13261 247109 13307 247120
rect 13375 247109 13421 247120
rect 13471 247109 13517 247120
rect 13585 247109 13631 247120
rect 13681 247109 13727 247120
rect 13795 247109 13841 247120
rect 13891 247109 13937 247120
rect 14005 247109 14051 247120
rect 14101 247109 14147 247120
rect 14215 247109 14261 247120
rect 14311 247109 14357 247120
rect 14425 247109 14471 247120
rect 14521 247109 14567 247120
rect 14635 247109 14681 247120
rect 14731 247109 14777 247120
rect 14845 247109 14891 247120
rect 14941 247109 14987 247120
rect 15055 247109 15101 247120
rect 15151 247109 15197 247120
rect 15265 247109 15311 247120
rect 15361 247109 15407 247120
rect 15475 247109 15521 247120
rect 15571 247109 15617 247120
rect 15685 247109 15731 247120
rect 15781 247109 15827 247120
rect 15895 247109 15941 247120
rect 15991 247109 16037 247120
rect 16105 247109 16151 247120
rect 16201 247109 16247 247120
rect 16315 247109 16361 247120
rect 16411 247109 16457 247120
rect 16525 247109 16571 247120
rect 16621 247109 16667 247120
rect 16735 247109 16781 247120
rect 16831 247109 16877 247120
rect 16945 247109 16991 247120
rect 17041 247109 17087 247120
rect 17155 247109 17201 247120
rect 17251 247109 17297 247120
rect 17365 247109 17411 247120
rect 17461 247109 17507 247120
rect 17575 247109 17621 247120
rect 17671 247109 17717 247120
rect 17785 247109 17831 247120
rect 17881 247109 17927 247120
rect 17995 247109 18041 247120
rect 18091 247109 18137 247120
rect 18205 247109 18251 247120
rect 18301 247109 18347 247120
rect 18415 247109 18461 247120
rect 18511 247109 18557 247120
rect 18625 247109 18671 247120
rect 18721 247109 18767 247120
rect 18835 247109 18881 247120
rect 18931 247109 18977 247120
rect 19045 247109 19091 247120
rect 19141 247109 19187 247120
rect 19255 247109 19301 247120
rect 19351 247109 19397 247120
rect 19465 247109 19511 247120
rect 19561 247109 19607 247120
rect 19675 247109 19721 247120
rect 19771 247109 19817 247120
rect 19885 247109 19931 247120
rect 19981 247109 20027 247120
rect 20095 247109 20141 247120
rect 20191 247109 20237 247120
rect 20305 247109 20351 247120
rect 20401 247109 20447 247120
rect 20515 247109 20561 247120
rect 20611 247109 20657 247120
rect 20725 247109 20771 247120
rect 20821 247109 20867 247120
rect 20935 247109 20981 247120
rect 21031 247109 21077 247120
rect 21145 247109 21191 247120
rect 21241 247109 21287 247120
rect 21355 247109 21401 247120
rect 21451 247109 21497 247120
rect 21565 247109 21611 247120
rect 21661 247109 21707 247120
rect 21775 247109 21821 247120
rect 21871 247109 21917 247120
rect 21985 247109 22031 247120
rect 22081 247109 22127 247120
rect 22195 247109 22241 247120
rect 22291 247109 22337 247120
rect 22405 247109 22451 247120
rect 22501 247109 22547 247120
rect 22615 247109 22661 247120
rect 22711 247109 22757 247120
rect 22825 247109 22871 247120
rect 22921 247109 22967 247120
rect 23035 247109 23081 247120
rect 23131 247109 23177 247120
rect 23245 247109 23291 247120
rect 23341 247109 23387 247120
rect 23455 247109 23501 247120
rect 23551 247109 23597 247120
rect 23665 247109 23711 247120
rect 23761 247109 23807 247120
rect 23875 247109 23921 247120
rect 23971 247109 24017 247120
rect 24085 247109 24131 247120
rect 24181 247109 24227 247120
rect 24295 247109 24341 247120
rect 24391 247109 24437 247120
rect 24505 247109 24551 247120
rect 24601 247109 24647 247120
rect 24715 247109 24761 247120
rect 24811 247109 24857 247120
rect 24925 247109 24971 247120
rect 25021 247109 25067 247120
rect 25135 247109 25181 247120
rect 25231 247109 25277 247120
rect 25345 247109 25391 247120
rect 25441 247109 25487 247120
rect 25555 247109 25601 247120
rect 25651 247109 25697 247120
rect 25765 247109 25811 247120
rect 25861 247109 25907 247120
rect 25975 247109 26021 247120
rect 26071 247109 26117 247120
rect 26185 247109 26231 247120
rect 26281 247109 26327 247120
rect 26395 247109 26441 247120
rect 26491 247109 26537 247120
rect 26605 247109 26651 247120
rect 26701 247109 26747 247120
rect 26815 247109 26861 247120
rect 26911 247109 26957 247120
rect 27025 247109 27071 247120
rect 27121 247109 27167 247120
rect 27235 247109 27281 247120
rect -4085 246332 -4075 247108
rect -4015 246332 -4005 247108
rect -3963 246332 -3953 247108
rect -3805 246332 -3795 247108
rect -3753 246332 -3743 247108
rect -3595 246332 -3585 247108
rect -3543 246332 -3533 247109
rect -3385 246332 -3375 247109
rect -3333 246332 -3323 247109
rect -3175 246332 -3165 247109
rect -3123 246332 -3113 247109
rect -2965 246332 -2955 247109
rect -2913 246332 -2903 247109
rect -2755 246332 -2745 247109
rect -2703 246332 -2693 247109
rect -2545 246332 -2535 247109
rect -2493 246332 -2483 247109
rect -2335 246332 -2325 247109
rect -2283 246332 -2273 247109
rect -2125 246332 -2115 247109
rect -2073 246332 -2063 247109
rect -1915 246332 -1905 247109
rect -1863 246332 -1853 247109
rect -1705 246332 -1695 247109
rect -1653 246332 -1643 247109
rect -1495 246332 -1485 247109
rect -1443 246332 -1433 247109
rect -1285 246332 -1275 247109
rect -1233 246332 -1223 247109
rect -1075 246332 -1065 247109
rect -1023 246332 -1013 247109
rect -865 246332 -855 247109
rect -813 246332 -803 247109
rect -655 246332 -645 247109
rect -603 246332 -593 247109
rect -445 246332 -435 247109
rect -393 246332 -383 247109
rect -235 246332 -225 247109
rect -183 246332 -173 247109
rect -25 246332 -15 247109
rect 27 246332 37 247109
rect 185 246332 195 247109
rect 237 246332 247 247109
rect 395 246332 405 247109
rect 447 246332 457 247109
rect 605 246332 615 247109
rect 657 246332 667 247109
rect 815 246332 825 247109
rect 867 246332 877 247109
rect 1025 246332 1035 247109
rect 1077 246332 1087 247109
rect 1235 246332 1245 247109
rect 1287 246332 1297 247109
rect 1445 246332 1455 247109
rect 1497 246332 1507 247109
rect 1655 246332 1665 247109
rect 1707 246332 1717 247109
rect 1865 246332 1875 247109
rect 1917 246332 1927 247109
rect 2075 246332 2085 247109
rect 2127 246332 2137 247109
rect 2285 246332 2295 247109
rect 2337 246332 2347 247109
rect 2495 246332 2505 247109
rect 2547 246332 2557 247109
rect 2705 246332 2715 247109
rect 2757 246332 2767 247109
rect 2915 246332 2925 247109
rect 2967 246332 2977 247109
rect 3125 246332 3135 247109
rect 3177 246332 3187 247109
rect 3335 246332 3345 247109
rect 3387 246332 3397 247109
rect 3545 246332 3555 247109
rect 3597 246332 3607 247109
rect 3755 246332 3765 247109
rect 3807 246332 3817 247109
rect 3965 246332 3975 247109
rect 4017 246332 4027 247109
rect 4175 246332 4185 247109
rect 4227 246332 4237 247109
rect 4385 246332 4395 247109
rect 4437 246332 4447 247109
rect 4595 246332 4605 247109
rect 4647 246332 4657 247109
rect 4805 246332 4815 247109
rect 4857 246332 4867 247109
rect 5015 246332 5025 247109
rect 5067 246332 5077 247109
rect 5225 246332 5235 247109
rect 5277 246332 5287 247109
rect 5435 246332 5445 247109
rect 5487 246332 5497 247109
rect 5645 246332 5655 247109
rect 5697 246332 5707 247109
rect 5855 246332 5865 247109
rect 5907 246332 5917 247109
rect 6065 246332 6075 247109
rect 6117 246332 6127 247109
rect 6275 246332 6285 247109
rect 6327 246332 6337 247109
rect 6485 246332 6495 247109
rect 6537 246332 6547 247109
rect 6695 246332 6705 247109
rect 6747 246332 6757 247109
rect 6905 246332 6915 247109
rect 6957 246332 6967 247109
rect 7115 246332 7125 247109
rect 7167 246332 7177 247109
rect 7325 246332 7335 247109
rect 7377 246332 7387 247109
rect 7535 246332 7545 247109
rect 7587 246332 7597 247109
rect 7745 246332 7755 247109
rect 7797 246332 7807 247109
rect 7955 246332 7965 247109
rect 8007 246332 8017 247109
rect 8165 246332 8175 247109
rect 8217 246332 8227 247109
rect 8375 246332 8385 247109
rect 8427 246332 8437 247109
rect 8585 246332 8595 247109
rect 8637 246332 8647 247109
rect 8795 246332 8805 247109
rect 8847 246332 8857 247109
rect 9005 246332 9015 247109
rect 9057 246332 9067 247109
rect 9215 246332 9225 247109
rect 9267 246332 9277 247109
rect 9425 246332 9435 247109
rect 9477 246332 9487 247109
rect 9635 246332 9645 247109
rect 9687 246332 9697 247109
rect 9845 246332 9855 247109
rect 9897 246332 9907 247109
rect 10055 246332 10065 247109
rect 10107 246332 10117 247109
rect 10265 246332 10275 247109
rect 10317 246332 10327 247109
rect 10475 246332 10485 247109
rect 10527 246332 10537 247109
rect 10685 246332 10695 247109
rect 10737 246332 10747 247109
rect 10895 246332 10905 247109
rect 10947 246332 10957 247109
rect 11105 246332 11115 247109
rect 11157 246332 11167 247109
rect 11315 246332 11325 247109
rect 11367 246332 11377 247109
rect 11525 246332 11535 247109
rect 11577 246332 11587 247109
rect 11735 246332 11745 247109
rect 11787 246332 11797 247109
rect 11945 246332 11955 247109
rect 11997 246332 12007 247109
rect 12155 246332 12165 247109
rect 12207 246332 12217 247109
rect 12365 246332 12375 247109
rect 12417 246332 12427 247109
rect 12575 246332 12585 247109
rect 12627 246332 12637 247109
rect 12785 246332 12795 247109
rect 12837 246332 12847 247109
rect 12995 246332 13005 247109
rect 13047 246332 13057 247109
rect 13205 246332 13215 247109
rect 13257 246332 13267 247109
rect 13415 246332 13425 247109
rect 13467 246332 13477 247109
rect 13625 246332 13635 247109
rect 13677 246332 13687 247109
rect 13835 246332 13845 247109
rect 13887 246332 13897 247109
rect 14045 246332 14055 247109
rect 14097 246332 14107 247109
rect 14255 246332 14265 247109
rect 14307 246332 14317 247109
rect 14465 246332 14475 247109
rect 14517 246332 14527 247109
rect 14675 246332 14685 247109
rect 14727 246332 14737 247109
rect 14885 246332 14895 247109
rect 14937 246332 14947 247109
rect 15095 246332 15105 247109
rect 15147 246332 15157 247109
rect 15305 246332 15315 247109
rect 15357 246332 15367 247109
rect 15515 246332 15525 247109
rect 15567 246332 15577 247109
rect 15725 246332 15735 247109
rect 15777 246332 15787 247109
rect 15935 246332 15945 247109
rect 15987 246332 15997 247109
rect 16145 246332 16155 247109
rect 16197 246332 16207 247109
rect 16355 246332 16365 247109
rect 16407 246332 16417 247109
rect 16565 246332 16575 247109
rect 16617 246332 16627 247109
rect 16775 246332 16785 247109
rect 16827 246332 16837 247109
rect 16985 246332 16995 247109
rect 17037 246332 17047 247109
rect 17195 246332 17205 247109
rect 17247 246332 17257 247109
rect 17405 246332 17415 247109
rect 17457 246332 17467 247109
rect 17615 246332 17625 247109
rect 17667 246332 17677 247109
rect 17825 246332 17835 247109
rect 17877 246332 17887 247109
rect 18035 246332 18045 247109
rect 18087 246332 18097 247109
rect 18245 246332 18255 247109
rect 18297 246332 18307 247109
rect 18455 246332 18465 247109
rect 18507 246332 18517 247109
rect 18665 246332 18675 247109
rect 18717 246332 18727 247109
rect 18875 246332 18885 247109
rect 18927 246332 18937 247109
rect 19085 246332 19095 247109
rect 19137 246332 19147 247109
rect 19295 246332 19305 247109
rect 19347 246332 19357 247109
rect 19505 246332 19515 247109
rect 19557 246332 19567 247109
rect 19715 246332 19725 247109
rect 19767 246332 19777 247109
rect 19925 246332 19935 247109
rect 19977 246332 19987 247109
rect 20135 246332 20145 247109
rect 20187 246332 20197 247109
rect 20345 246332 20355 247109
rect 20397 246332 20407 247109
rect 20555 246332 20565 247109
rect 20607 246332 20617 247109
rect 20765 246332 20775 247109
rect 20817 246332 20827 247109
rect 20975 246332 20985 247109
rect 21027 246332 21037 247109
rect 21185 246332 21195 247109
rect 21237 246332 21247 247109
rect 21395 246332 21405 247109
rect 21447 246332 21457 247109
rect 21605 246332 21615 247109
rect 21657 246332 21667 247109
rect 21815 246332 21825 247109
rect 21867 246332 21877 247109
rect 22025 246332 22035 247109
rect 22077 246332 22087 247109
rect 22235 246332 22245 247109
rect 22287 246332 22297 247109
rect 22445 246332 22455 247109
rect 22497 246332 22507 247109
rect 22655 246332 22665 247109
rect 22707 246332 22717 247109
rect 22865 246332 22875 247109
rect 22917 246332 22927 247109
rect 23075 246332 23085 247109
rect 23127 246332 23137 247109
rect 23285 246332 23295 247109
rect 23337 246332 23347 247109
rect 23495 246332 23505 247109
rect 23547 246332 23557 247109
rect 23705 246332 23715 247109
rect 23757 246332 23767 247109
rect 23915 246332 23925 247109
rect 23967 246332 23977 247109
rect 24125 246332 24135 247109
rect 24177 246332 24187 247109
rect 24335 246332 24345 247109
rect 24387 246332 24397 247109
rect 24545 246332 24555 247109
rect 24597 246332 24607 247109
rect 24755 246332 24765 247109
rect 24807 246332 24817 247109
rect 24965 246332 24975 247109
rect 25017 246332 25027 247109
rect 25175 246332 25185 247109
rect 25227 246332 25237 247109
rect 25385 246332 25395 247109
rect 25437 246332 25447 247109
rect 25595 246332 25605 247109
rect 25647 246332 25657 247109
rect 25805 246332 25815 247109
rect 25857 246332 25867 247109
rect 26015 246332 26025 247109
rect 26067 246332 26077 247109
rect 26225 246332 26235 247109
rect 26277 246332 26287 247109
rect 26435 246332 26445 247109
rect 26487 246332 26497 247109
rect 26645 246332 26655 247109
rect 26697 246332 26707 247109
rect 26855 246332 26865 247109
rect 26907 246332 26917 247109
rect 27065 246332 27075 247109
rect 27117 246332 27127 247109
rect 27275 246332 27285 247109
rect 27331 247108 27566 247120
rect 27331 246332 27337 247108
rect 27371 246332 27566 247108
rect -4055 246320 -4009 246332
rect -3959 246320 -3913 246332
rect -3845 246320 -3799 246332
rect -3749 246320 -3703 246332
rect -3635 246320 -3589 246332
rect -3539 246320 -3493 246332
rect -3425 246320 -3379 246332
rect -3329 246320 -3283 246332
rect -3215 246320 -3169 246332
rect -3119 246320 -3073 246332
rect -3005 246320 -2959 246332
rect -2909 246320 -2863 246332
rect -2795 246320 -2749 246332
rect -2699 246320 -2653 246332
rect -2585 246320 -2539 246332
rect -2489 246320 -2443 246332
rect -2375 246320 -2329 246332
rect -2279 246320 -2233 246332
rect -2165 246320 -2119 246332
rect -2069 246320 -2023 246332
rect -1955 246320 -1909 246332
rect -1859 246320 -1813 246332
rect -1745 246320 -1699 246332
rect -1649 246320 -1603 246332
rect -1535 246320 -1489 246332
rect -1439 246320 -1393 246332
rect -1325 246320 -1279 246332
rect -1229 246320 -1183 246332
rect -1115 246320 -1069 246332
rect -1019 246320 -973 246332
rect -905 246320 -859 246332
rect -809 246320 -763 246332
rect -695 246320 -649 246332
rect -599 246320 -553 246332
rect -485 246320 -439 246332
rect -389 246320 -343 246332
rect -275 246320 -229 246332
rect -179 246320 -133 246332
rect -65 246320 -19 246332
rect 31 246320 77 246332
rect 145 246320 191 246332
rect 241 246320 287 246332
rect 355 246320 401 246332
rect 451 246320 497 246332
rect 565 246320 611 246332
rect 661 246320 707 246332
rect 775 246320 821 246332
rect 871 246320 917 246332
rect 985 246320 1031 246332
rect 1081 246320 1127 246332
rect 1195 246320 1241 246332
rect 1291 246320 1337 246332
rect 1405 246320 1451 246332
rect 1501 246320 1547 246332
rect 1615 246320 1661 246332
rect 1711 246320 1757 246332
rect 1825 246320 1871 246332
rect 1921 246320 1967 246332
rect 2035 246320 2081 246332
rect 2131 246320 2177 246332
rect 2245 246320 2291 246332
rect 2341 246320 2387 246332
rect 2455 246320 2501 246332
rect 2551 246320 2597 246332
rect 2665 246320 2711 246332
rect 2761 246320 2807 246332
rect 2875 246320 2921 246332
rect 2971 246320 3017 246332
rect 3085 246320 3131 246332
rect 3181 246320 3227 246332
rect 3295 246320 3341 246332
rect 3391 246320 3437 246332
rect 3505 246320 3551 246332
rect 3601 246320 3647 246332
rect 3715 246320 3761 246332
rect 3811 246320 3857 246332
rect 3925 246320 3971 246332
rect 4021 246320 4067 246332
rect 4135 246320 4181 246332
rect 4231 246320 4277 246332
rect 4345 246320 4391 246332
rect 4441 246320 4487 246332
rect 4555 246320 4601 246332
rect 4651 246320 4697 246332
rect 4765 246320 4811 246332
rect 4861 246320 4907 246332
rect 4975 246320 5021 246332
rect 5071 246320 5117 246332
rect 5185 246320 5231 246332
rect 5281 246320 5327 246332
rect 5395 246320 5441 246332
rect 5491 246320 5537 246332
rect 5605 246320 5651 246332
rect 5701 246320 5747 246332
rect 5815 246320 5861 246332
rect 5911 246320 5957 246332
rect 6025 246320 6071 246332
rect 6121 246320 6167 246332
rect 6235 246320 6281 246332
rect 6331 246320 6377 246332
rect 6445 246320 6491 246332
rect 6541 246320 6587 246332
rect 6655 246320 6701 246332
rect 6751 246320 6797 246332
rect 6865 246320 6911 246332
rect 6961 246320 7007 246332
rect 7075 246320 7121 246332
rect 7171 246320 7217 246332
rect 7285 246320 7331 246332
rect 7381 246320 7427 246332
rect 7495 246320 7541 246332
rect 7591 246320 7637 246332
rect 7705 246320 7751 246332
rect 7801 246320 7847 246332
rect 7915 246320 7961 246332
rect 8011 246320 8057 246332
rect 8125 246320 8171 246332
rect 8221 246320 8267 246332
rect 8335 246320 8381 246332
rect 8431 246320 8477 246332
rect 8545 246320 8591 246332
rect 8641 246320 8687 246332
rect 8755 246320 8801 246332
rect 8851 246320 8897 246332
rect 8965 246320 9011 246332
rect 9061 246320 9107 246332
rect 9175 246320 9221 246332
rect 9271 246320 9317 246332
rect 9385 246320 9431 246332
rect 9481 246320 9527 246332
rect 9595 246320 9641 246332
rect 9691 246320 9737 246332
rect 9805 246320 9851 246332
rect 9901 246320 9947 246332
rect 10015 246320 10061 246332
rect 10111 246320 10157 246332
rect 10225 246320 10271 246332
rect 10321 246320 10367 246332
rect 10435 246320 10481 246332
rect 10531 246320 10577 246332
rect 10645 246320 10691 246332
rect 10741 246320 10787 246332
rect 10855 246320 10901 246332
rect 10951 246320 10997 246332
rect 11065 246320 11111 246332
rect 11161 246320 11207 246332
rect 11275 246320 11321 246332
rect 11371 246320 11417 246332
rect 11485 246320 11531 246332
rect 11581 246320 11627 246332
rect 11695 246320 11741 246332
rect 11791 246320 11837 246332
rect 11905 246320 11951 246332
rect 12001 246320 12047 246332
rect 12115 246320 12161 246332
rect 12211 246320 12257 246332
rect 12325 246320 12371 246332
rect 12421 246320 12467 246332
rect 12535 246320 12581 246332
rect 12631 246320 12677 246332
rect 12745 246320 12791 246332
rect 12841 246320 12887 246332
rect 12955 246320 13001 246332
rect 13051 246320 13097 246332
rect 13165 246320 13211 246332
rect 13261 246320 13307 246332
rect 13375 246320 13421 246332
rect 13471 246320 13517 246332
rect 13585 246320 13631 246332
rect 13681 246320 13727 246332
rect 13795 246320 13841 246332
rect 13891 246320 13937 246332
rect 14005 246320 14051 246332
rect 14101 246320 14147 246332
rect 14215 246320 14261 246332
rect 14311 246320 14357 246332
rect 14425 246320 14471 246332
rect 14521 246320 14567 246332
rect 14635 246320 14681 246332
rect 14731 246320 14777 246332
rect 14845 246320 14891 246332
rect 14941 246320 14987 246332
rect 15055 246320 15101 246332
rect 15151 246320 15197 246332
rect 15265 246320 15311 246332
rect 15361 246320 15407 246332
rect 15475 246320 15521 246332
rect 15571 246320 15617 246332
rect 15685 246320 15731 246332
rect 15781 246320 15827 246332
rect 15895 246320 15941 246332
rect 15991 246320 16037 246332
rect 16105 246320 16151 246332
rect 16201 246320 16247 246332
rect 16315 246320 16361 246332
rect 16411 246320 16457 246332
rect 16525 246320 16571 246332
rect 16621 246320 16667 246332
rect 16735 246320 16781 246332
rect 16831 246320 16877 246332
rect 16945 246320 16991 246332
rect 17041 246320 17087 246332
rect 17155 246320 17201 246332
rect 17251 246320 17297 246332
rect 17365 246320 17411 246332
rect 17461 246320 17507 246332
rect 17575 246320 17621 246332
rect 17671 246320 17717 246332
rect 17785 246320 17831 246332
rect 17881 246320 17927 246332
rect 17995 246320 18041 246332
rect 18091 246320 18137 246332
rect 18205 246320 18251 246332
rect 18301 246320 18347 246332
rect 18415 246320 18461 246332
rect 18511 246320 18557 246332
rect 18625 246320 18671 246332
rect 18721 246320 18767 246332
rect 18835 246320 18881 246332
rect 18931 246320 18977 246332
rect 19045 246320 19091 246332
rect 19141 246320 19187 246332
rect 19255 246320 19301 246332
rect 19351 246320 19397 246332
rect 19465 246320 19511 246332
rect 19561 246320 19607 246332
rect 19675 246320 19721 246332
rect 19771 246320 19817 246332
rect 19885 246320 19931 246332
rect 19981 246320 20027 246332
rect 20095 246320 20141 246332
rect 20191 246320 20237 246332
rect 20305 246320 20351 246332
rect 20401 246320 20447 246332
rect 20515 246320 20561 246332
rect 20611 246320 20657 246332
rect 20725 246320 20771 246332
rect 20821 246320 20867 246332
rect 20935 246320 20981 246332
rect 21031 246320 21077 246332
rect 21145 246320 21191 246332
rect 21241 246320 21287 246332
rect 21355 246320 21401 246332
rect 21451 246320 21497 246332
rect 21565 246320 21611 246332
rect 21661 246320 21707 246332
rect 21775 246320 21821 246332
rect 21871 246320 21917 246332
rect 21985 246320 22031 246332
rect 22081 246320 22127 246332
rect 22195 246320 22241 246332
rect 22291 246320 22337 246332
rect 22405 246320 22451 246332
rect 22501 246320 22547 246332
rect 22615 246320 22661 246332
rect 22711 246320 22757 246332
rect 22825 246320 22871 246332
rect 22921 246320 22967 246332
rect 23035 246320 23081 246332
rect 23131 246320 23177 246332
rect 23245 246320 23291 246332
rect 23341 246320 23387 246332
rect 23455 246320 23501 246332
rect 23551 246320 23597 246332
rect 23665 246320 23711 246332
rect 23761 246320 23807 246332
rect 23875 246320 23921 246332
rect 23971 246320 24017 246332
rect 24085 246320 24131 246332
rect 24181 246320 24227 246332
rect 24295 246320 24341 246332
rect 24391 246320 24437 246332
rect 24505 246320 24551 246332
rect 24601 246320 24647 246332
rect 24715 246320 24761 246332
rect 24811 246320 24857 246332
rect 24925 246320 24971 246332
rect 25021 246320 25067 246332
rect 25135 246320 25181 246332
rect 25231 246320 25277 246332
rect 25345 246320 25391 246332
rect 25441 246320 25487 246332
rect 25555 246320 25601 246332
rect 25651 246320 25697 246332
rect 25765 246320 25811 246332
rect 25861 246320 25907 246332
rect 25975 246320 26021 246332
rect 26071 246320 26117 246332
rect 26185 246320 26231 246332
rect 26281 246320 26327 246332
rect 26395 246320 26441 246332
rect 26491 246320 26537 246332
rect 26605 246320 26651 246332
rect 26701 246320 26747 246332
rect 26815 246320 26861 246332
rect 26911 246320 26957 246332
rect 27025 246320 27071 246332
rect 27121 246320 27167 246332
rect 27235 246320 27281 246332
rect 27331 246320 27566 246332
rect -3803 246273 27335 246285
rect -5008 246131 -3791 246273
rect -3757 246131 -3371 246273
rect -3337 246131 -2951 246273
rect -2917 246131 -2531 246273
rect -2497 246131 -2111 246273
rect -2077 246131 -1691 246273
rect -1657 246131 -1271 246273
rect -1237 246131 -851 246273
rect -817 246131 -431 246273
rect -397 246131 -11 246273
rect 23 246131 409 246273
rect 443 246131 829 246273
rect 863 246131 1249 246273
rect 1283 246131 1669 246273
rect 1703 246131 2089 246273
rect 2123 246131 2509 246273
rect 2543 246131 2929 246273
rect 2963 246131 3349 246273
rect 3383 246131 3769 246273
rect 3803 246131 4189 246273
rect 4223 246131 4609 246273
rect 4643 246131 5029 246273
rect 5063 246131 5449 246273
rect 5483 246131 5869 246273
rect 5903 246131 6289 246273
rect 6323 246131 6709 246273
rect 6743 246131 7129 246273
rect 7163 246131 7549 246273
rect 7583 246131 7969 246273
rect 8003 246131 8389 246273
rect 8423 246131 8809 246273
rect 8843 246131 9229 246273
rect 9263 246131 9649 246273
rect 9683 246131 10069 246273
rect 10103 246131 10489 246273
rect 10523 246131 10909 246273
rect 10943 246131 11329 246273
rect 11363 246131 11749 246273
rect 11783 246131 12169 246273
rect 12203 246131 12589 246273
rect 12623 246131 13009 246273
rect 13043 246131 13429 246273
rect 13463 246131 13849 246273
rect 13883 246131 14269 246273
rect 14303 246131 14689 246273
rect 14723 246131 15109 246273
rect 15143 246131 15529 246273
rect 15563 246131 15949 246273
rect 15983 246131 16369 246273
rect 16403 246131 16789 246273
rect 16823 246131 17209 246273
rect 17243 246131 17629 246273
rect 17663 246131 18049 246273
rect 18083 246131 18469 246273
rect 18503 246131 18889 246273
rect 18923 246131 19309 246273
rect 19343 246131 19729 246273
rect 19763 246131 20149 246273
rect 20183 246131 20569 246273
rect 20603 246131 20989 246273
rect 21023 246131 21409 246273
rect 21443 246131 21829 246273
rect 21863 246131 22249 246273
rect 22283 246131 22669 246273
rect 22703 246131 23089 246273
rect 23123 246131 23509 246273
rect 23543 246131 23929 246273
rect 23963 246131 24349 246273
rect 24383 246131 24769 246273
rect 24803 246131 25189 246273
rect 25223 246131 25609 246273
rect 25643 246131 26029 246273
rect 26063 246131 26449 246273
rect 26483 246131 26869 246273
rect 26903 246131 27289 246273
rect 27323 246131 27335 246273
rect -5008 245237 -4142 246131
rect -3803 246119 27335 246131
rect 27377 246084 27566 246320
rect -4055 246072 -4009 246084
rect -3959 246072 -3913 246084
rect -3845 246072 -3799 246084
rect -3749 246072 -3703 246084
rect -3635 246072 -3589 246084
rect -3539 246073 -3493 246084
rect -3425 246073 -3379 246084
rect -3329 246073 -3283 246084
rect -3215 246073 -3169 246084
rect -3119 246073 -3073 246084
rect -3005 246073 -2959 246084
rect -2909 246073 -2863 246084
rect -2795 246073 -2749 246084
rect -2699 246073 -2653 246084
rect -2585 246073 -2539 246084
rect -2489 246073 -2443 246084
rect -2375 246073 -2329 246084
rect -2279 246073 -2233 246084
rect -2165 246073 -2119 246084
rect -2069 246073 -2023 246084
rect -1955 246073 -1909 246084
rect -1859 246073 -1813 246084
rect -1745 246073 -1699 246084
rect -1649 246073 -1603 246084
rect -1535 246073 -1489 246084
rect -1439 246073 -1393 246084
rect -1325 246073 -1279 246084
rect -1229 246073 -1183 246084
rect -1115 246073 -1069 246084
rect -1019 246073 -973 246084
rect -905 246073 -859 246084
rect -809 246073 -763 246084
rect -695 246073 -649 246084
rect -599 246073 -553 246084
rect -485 246073 -439 246084
rect -389 246073 -343 246084
rect -275 246073 -229 246084
rect -179 246073 -133 246084
rect -65 246073 -19 246084
rect 31 246073 77 246084
rect 145 246073 191 246084
rect 241 246073 287 246084
rect 355 246073 401 246084
rect 451 246073 497 246084
rect 565 246073 611 246084
rect 661 246073 707 246084
rect 775 246073 821 246084
rect 871 246073 917 246084
rect 985 246073 1031 246084
rect 1081 246073 1127 246084
rect 1195 246073 1241 246084
rect 1291 246073 1337 246084
rect 1405 246073 1451 246084
rect 1501 246073 1547 246084
rect 1615 246073 1661 246084
rect 1711 246073 1757 246084
rect 1825 246073 1871 246084
rect 1921 246073 1967 246084
rect 2035 246073 2081 246084
rect 2131 246073 2177 246084
rect 2245 246073 2291 246084
rect 2341 246073 2387 246084
rect 2455 246073 2501 246084
rect 2551 246073 2597 246084
rect 2665 246073 2711 246084
rect 2761 246073 2807 246084
rect 2875 246073 2921 246084
rect 2971 246073 3017 246084
rect 3085 246073 3131 246084
rect 3181 246073 3227 246084
rect 3295 246073 3341 246084
rect 3391 246073 3437 246084
rect 3505 246073 3551 246084
rect 3601 246073 3647 246084
rect 3715 246073 3761 246084
rect 3811 246073 3857 246084
rect 3925 246073 3971 246084
rect 4021 246073 4067 246084
rect 4135 246073 4181 246084
rect 4231 246073 4277 246084
rect 4345 246073 4391 246084
rect 4441 246073 4487 246084
rect 4555 246073 4601 246084
rect 4651 246073 4697 246084
rect 4765 246073 4811 246084
rect 4861 246073 4907 246084
rect 4975 246073 5021 246084
rect 5071 246073 5117 246084
rect 5185 246073 5231 246084
rect 5281 246073 5327 246084
rect 5395 246073 5441 246084
rect 5491 246073 5537 246084
rect 5605 246073 5651 246084
rect 5701 246073 5747 246084
rect 5815 246073 5861 246084
rect 5911 246073 5957 246084
rect 6025 246073 6071 246084
rect 6121 246073 6167 246084
rect 6235 246073 6281 246084
rect 6331 246073 6377 246084
rect 6445 246073 6491 246084
rect 6541 246073 6587 246084
rect 6655 246073 6701 246084
rect 6751 246073 6797 246084
rect 6865 246073 6911 246084
rect 6961 246073 7007 246084
rect 7075 246073 7121 246084
rect 7171 246073 7217 246084
rect 7285 246073 7331 246084
rect 7381 246073 7427 246084
rect 7495 246073 7541 246084
rect 7591 246073 7637 246084
rect 7705 246073 7751 246084
rect 7801 246073 7847 246084
rect 7915 246073 7961 246084
rect 8011 246073 8057 246084
rect 8125 246073 8171 246084
rect 8221 246073 8267 246084
rect 8335 246073 8381 246084
rect 8431 246073 8477 246084
rect 8545 246073 8591 246084
rect 8641 246073 8687 246084
rect 8755 246073 8801 246084
rect 8851 246073 8897 246084
rect 8965 246073 9011 246084
rect 9061 246073 9107 246084
rect 9175 246073 9221 246084
rect 9271 246073 9317 246084
rect 9385 246073 9431 246084
rect 9481 246073 9527 246084
rect 9595 246073 9641 246084
rect 9691 246073 9737 246084
rect 9805 246073 9851 246084
rect 9901 246073 9947 246084
rect 10015 246073 10061 246084
rect 10111 246073 10157 246084
rect 10225 246073 10271 246084
rect 10321 246073 10367 246084
rect 10435 246073 10481 246084
rect 10531 246073 10577 246084
rect 10645 246073 10691 246084
rect 10741 246073 10787 246084
rect 10855 246073 10901 246084
rect 10951 246073 10997 246084
rect 11065 246073 11111 246084
rect 11161 246073 11207 246084
rect 11275 246073 11321 246084
rect 11371 246073 11417 246084
rect 11485 246073 11531 246084
rect 11581 246073 11627 246084
rect 11695 246073 11741 246084
rect 11791 246073 11837 246084
rect 11905 246073 11951 246084
rect 12001 246073 12047 246084
rect 12115 246073 12161 246084
rect 12211 246073 12257 246084
rect 12325 246073 12371 246084
rect 12421 246073 12467 246084
rect 12535 246073 12581 246084
rect 12631 246073 12677 246084
rect 12745 246073 12791 246084
rect 12841 246073 12887 246084
rect 12955 246073 13001 246084
rect 13051 246073 13097 246084
rect 13165 246073 13211 246084
rect 13261 246073 13307 246084
rect 13375 246073 13421 246084
rect 13471 246073 13517 246084
rect 13585 246073 13631 246084
rect 13681 246073 13727 246084
rect 13795 246073 13841 246084
rect 13891 246073 13937 246084
rect 14005 246073 14051 246084
rect 14101 246073 14147 246084
rect 14215 246073 14261 246084
rect 14311 246073 14357 246084
rect 14425 246073 14471 246084
rect 14521 246073 14567 246084
rect 14635 246073 14681 246084
rect 14731 246073 14777 246084
rect 14845 246073 14891 246084
rect 14941 246073 14987 246084
rect 15055 246073 15101 246084
rect 15151 246073 15197 246084
rect 15265 246073 15311 246084
rect 15361 246073 15407 246084
rect 15475 246073 15521 246084
rect 15571 246073 15617 246084
rect 15685 246073 15731 246084
rect 15781 246073 15827 246084
rect 15895 246073 15941 246084
rect 15991 246073 16037 246084
rect 16105 246073 16151 246084
rect 16201 246073 16247 246084
rect 16315 246073 16361 246084
rect 16411 246073 16457 246084
rect 16525 246073 16571 246084
rect 16621 246073 16667 246084
rect 16735 246073 16781 246084
rect 16831 246073 16877 246084
rect 16945 246073 16991 246084
rect 17041 246073 17087 246084
rect 17155 246073 17201 246084
rect 17251 246073 17297 246084
rect 17365 246073 17411 246084
rect 17461 246073 17507 246084
rect 17575 246073 17621 246084
rect 17671 246073 17717 246084
rect 17785 246073 17831 246084
rect 17881 246073 17927 246084
rect 17995 246073 18041 246084
rect 18091 246073 18137 246084
rect 18205 246073 18251 246084
rect 18301 246073 18347 246084
rect 18415 246073 18461 246084
rect 18511 246073 18557 246084
rect 18625 246073 18671 246084
rect 18721 246073 18767 246084
rect 18835 246073 18881 246084
rect 18931 246073 18977 246084
rect 19045 246073 19091 246084
rect 19141 246073 19187 246084
rect 19255 246073 19301 246084
rect 19351 246073 19397 246084
rect 19465 246073 19511 246084
rect 19561 246073 19607 246084
rect 19675 246073 19721 246084
rect 19771 246073 19817 246084
rect 19885 246073 19931 246084
rect 19981 246073 20027 246084
rect 20095 246073 20141 246084
rect 20191 246073 20237 246084
rect 20305 246073 20351 246084
rect 20401 246073 20447 246084
rect 20515 246073 20561 246084
rect 20611 246073 20657 246084
rect 20725 246073 20771 246084
rect 20821 246073 20867 246084
rect 20935 246073 20981 246084
rect 21031 246073 21077 246084
rect 21145 246073 21191 246084
rect 21241 246073 21287 246084
rect 21355 246073 21401 246084
rect 21451 246073 21497 246084
rect 21565 246073 21611 246084
rect 21661 246073 21707 246084
rect 21775 246073 21821 246084
rect 21871 246073 21917 246084
rect 21985 246073 22031 246084
rect 22081 246073 22127 246084
rect 22195 246073 22241 246084
rect 22291 246073 22337 246084
rect 22405 246073 22451 246084
rect 22501 246073 22547 246084
rect 22615 246073 22661 246084
rect 22711 246073 22757 246084
rect 22825 246073 22871 246084
rect 22921 246073 22967 246084
rect 23035 246073 23081 246084
rect 23131 246073 23177 246084
rect 23245 246073 23291 246084
rect 23341 246073 23387 246084
rect 23455 246073 23501 246084
rect 23551 246073 23597 246084
rect 23665 246073 23711 246084
rect 23761 246073 23807 246084
rect 23875 246073 23921 246084
rect 23971 246073 24017 246084
rect 24085 246073 24131 246084
rect 24181 246073 24227 246084
rect 24295 246073 24341 246084
rect 24391 246073 24437 246084
rect 24505 246073 24551 246084
rect 24601 246073 24647 246084
rect 24715 246073 24761 246084
rect 24811 246073 24857 246084
rect 24925 246073 24971 246084
rect 25021 246073 25067 246084
rect 25135 246073 25181 246084
rect 25231 246073 25277 246084
rect 25345 246073 25391 246084
rect 25441 246073 25487 246084
rect 25555 246073 25601 246084
rect 25651 246073 25697 246084
rect 25765 246073 25811 246084
rect 25861 246073 25907 246084
rect 25975 246073 26021 246084
rect 26071 246073 26117 246084
rect 26185 246073 26231 246084
rect 26281 246073 26327 246084
rect 26395 246073 26441 246084
rect 26491 246073 26537 246084
rect 26605 246073 26651 246084
rect 26701 246073 26747 246084
rect 26815 246073 26861 246084
rect 26911 246073 26957 246084
rect 27025 246073 27071 246084
rect 27121 246073 27167 246084
rect 27235 246073 27281 246084
rect -4085 245296 -4075 246072
rect -4015 245296 -4005 246072
rect -3963 245296 -3953 246072
rect -3805 245296 -3795 246072
rect -3753 245296 -3743 246072
rect -3595 245296 -3585 246072
rect -3543 245296 -3533 246073
rect -3385 245296 -3375 246073
rect -3333 245296 -3323 246073
rect -3175 245296 -3165 246073
rect -3123 245296 -3113 246073
rect -2965 245296 -2955 246073
rect -2913 245296 -2903 246073
rect -2755 245296 -2745 246073
rect -2703 245296 -2693 246073
rect -2545 245296 -2535 246073
rect -2493 245296 -2483 246073
rect -2335 245296 -2325 246073
rect -2283 245296 -2273 246073
rect -2125 245296 -2115 246073
rect -2073 245296 -2063 246073
rect -1915 245296 -1905 246073
rect -1863 245296 -1853 246073
rect -1705 245296 -1695 246073
rect -1653 245296 -1643 246073
rect -1495 245296 -1485 246073
rect -1443 245296 -1433 246073
rect -1285 245296 -1275 246073
rect -1233 245296 -1223 246073
rect -1075 245296 -1065 246073
rect -1023 245296 -1013 246073
rect -865 245296 -855 246073
rect -813 245296 -803 246073
rect -655 245296 -645 246073
rect -603 245296 -593 246073
rect -445 245296 -435 246073
rect -393 245296 -383 246073
rect -235 245296 -225 246073
rect -183 245296 -173 246073
rect -25 245296 -15 246073
rect 27 245296 37 246073
rect 185 245296 195 246073
rect 237 245296 247 246073
rect 395 245296 405 246073
rect 447 245296 457 246073
rect 605 245296 615 246073
rect 657 245296 667 246073
rect 815 245296 825 246073
rect 867 245296 877 246073
rect 1025 245296 1035 246073
rect 1077 245296 1087 246073
rect 1235 245296 1245 246073
rect 1287 245296 1297 246073
rect 1445 245296 1455 246073
rect 1497 245296 1507 246073
rect 1655 245296 1665 246073
rect 1707 245296 1717 246073
rect 1865 245296 1875 246073
rect 1917 245296 1927 246073
rect 2075 245296 2085 246073
rect 2127 245296 2137 246073
rect 2285 245296 2295 246073
rect 2337 245296 2347 246073
rect 2495 245296 2505 246073
rect 2547 245296 2557 246073
rect 2705 245296 2715 246073
rect 2757 245296 2767 246073
rect 2915 245296 2925 246073
rect 2967 245296 2977 246073
rect 3125 245296 3135 246073
rect 3177 245296 3187 246073
rect 3335 245296 3345 246073
rect 3387 245296 3397 246073
rect 3545 245296 3555 246073
rect 3597 245296 3607 246073
rect 3755 245296 3765 246073
rect 3807 245296 3817 246073
rect 3965 245296 3975 246073
rect 4017 245296 4027 246073
rect 4175 245296 4185 246073
rect 4227 245296 4237 246073
rect 4385 245296 4395 246073
rect 4437 245296 4447 246073
rect 4595 245296 4605 246073
rect 4647 245296 4657 246073
rect 4805 245296 4815 246073
rect 4857 245296 4867 246073
rect 5015 245296 5025 246073
rect 5067 245296 5077 246073
rect 5225 245296 5235 246073
rect 5277 245296 5287 246073
rect 5435 245296 5445 246073
rect 5487 245296 5497 246073
rect 5645 245296 5655 246073
rect 5697 245296 5707 246073
rect 5855 245296 5865 246073
rect 5907 245296 5917 246073
rect 6065 245296 6075 246073
rect 6117 245296 6127 246073
rect 6275 245296 6285 246073
rect 6327 245296 6337 246073
rect 6485 245296 6495 246073
rect 6537 245296 6547 246073
rect 6695 245296 6705 246073
rect 6747 245296 6757 246073
rect 6905 245296 6915 246073
rect 6957 245296 6967 246073
rect 7115 245296 7125 246073
rect 7167 245296 7177 246073
rect 7325 245296 7335 246073
rect 7377 245296 7387 246073
rect 7535 245296 7545 246073
rect 7587 245296 7597 246073
rect 7745 245296 7755 246073
rect 7797 245296 7807 246073
rect 7955 245296 7965 246073
rect 8007 245296 8017 246073
rect 8165 245296 8175 246073
rect 8217 245296 8227 246073
rect 8375 245296 8385 246073
rect 8427 245296 8437 246073
rect 8585 245296 8595 246073
rect 8637 245296 8647 246073
rect 8795 245296 8805 246073
rect 8847 245296 8857 246073
rect 9005 245296 9015 246073
rect 9057 245296 9067 246073
rect 9215 245296 9225 246073
rect 9267 245296 9277 246073
rect 9425 245296 9435 246073
rect 9477 245296 9487 246073
rect 9635 245296 9645 246073
rect 9687 245296 9697 246073
rect 9845 245296 9855 246073
rect 9897 245296 9907 246073
rect 10055 245296 10065 246073
rect 10107 245296 10117 246073
rect 10265 245296 10275 246073
rect 10317 245296 10327 246073
rect 10475 245296 10485 246073
rect 10527 245296 10537 246073
rect 10685 245296 10695 246073
rect 10737 245296 10747 246073
rect 10895 245296 10905 246073
rect 10947 245296 10957 246073
rect 11105 245296 11115 246073
rect 11157 245296 11167 246073
rect 11315 245296 11325 246073
rect 11367 245296 11377 246073
rect 11525 245296 11535 246073
rect 11577 245296 11587 246073
rect 11735 245296 11745 246073
rect 11787 245296 11797 246073
rect 11945 245296 11955 246073
rect 11997 245296 12007 246073
rect 12155 245296 12165 246073
rect 12207 245296 12217 246073
rect 12365 245296 12375 246073
rect 12417 245296 12427 246073
rect 12575 245296 12585 246073
rect 12627 245296 12637 246073
rect 12785 245296 12795 246073
rect 12837 245296 12847 246073
rect 12995 245296 13005 246073
rect 13047 245296 13057 246073
rect 13205 245296 13215 246073
rect 13257 245296 13267 246073
rect 13415 245296 13425 246073
rect 13467 245296 13477 246073
rect 13625 245296 13635 246073
rect 13677 245296 13687 246073
rect 13835 245296 13845 246073
rect 13887 245296 13897 246073
rect 14045 245296 14055 246073
rect 14097 245296 14107 246073
rect 14255 245296 14265 246073
rect 14307 245296 14317 246073
rect 14465 245296 14475 246073
rect 14517 245296 14527 246073
rect 14675 245296 14685 246073
rect 14727 245296 14737 246073
rect 14885 245296 14895 246073
rect 14937 245296 14947 246073
rect 15095 245296 15105 246073
rect 15147 245296 15157 246073
rect 15305 245296 15315 246073
rect 15357 245296 15367 246073
rect 15515 245296 15525 246073
rect 15567 245296 15577 246073
rect 15725 245296 15735 246073
rect 15777 245296 15787 246073
rect 15935 245296 15945 246073
rect 15987 245296 15997 246073
rect 16145 245296 16155 246073
rect 16197 245296 16207 246073
rect 16355 245296 16365 246073
rect 16407 245296 16417 246073
rect 16565 245296 16575 246073
rect 16617 245296 16627 246073
rect 16775 245296 16785 246073
rect 16827 245296 16837 246073
rect 16985 245296 16995 246073
rect 17037 245296 17047 246073
rect 17195 245296 17205 246073
rect 17247 245296 17257 246073
rect 17405 245296 17415 246073
rect 17457 245296 17467 246073
rect 17615 245296 17625 246073
rect 17667 245296 17677 246073
rect 17825 245296 17835 246073
rect 17877 245296 17887 246073
rect 18035 245296 18045 246073
rect 18087 245296 18097 246073
rect 18245 245296 18255 246073
rect 18297 245296 18307 246073
rect 18455 245296 18465 246073
rect 18507 245296 18517 246073
rect 18665 245296 18675 246073
rect 18717 245296 18727 246073
rect 18875 245296 18885 246073
rect 18927 245296 18937 246073
rect 19085 245296 19095 246073
rect 19137 245296 19147 246073
rect 19295 245296 19305 246073
rect 19347 245296 19357 246073
rect 19505 245296 19515 246073
rect 19557 245296 19567 246073
rect 19715 245296 19725 246073
rect 19767 245296 19777 246073
rect 19925 245296 19935 246073
rect 19977 245296 19987 246073
rect 20135 245296 20145 246073
rect 20187 245296 20197 246073
rect 20345 245296 20355 246073
rect 20397 245296 20407 246073
rect 20555 245296 20565 246073
rect 20607 245296 20617 246073
rect 20765 245296 20775 246073
rect 20817 245296 20827 246073
rect 20975 245296 20985 246073
rect 21027 245296 21037 246073
rect 21185 245296 21195 246073
rect 21237 245296 21247 246073
rect 21395 245296 21405 246073
rect 21447 245296 21457 246073
rect 21605 245296 21615 246073
rect 21657 245296 21667 246073
rect 21815 245296 21825 246073
rect 21867 245296 21877 246073
rect 22025 245296 22035 246073
rect 22077 245296 22087 246073
rect 22235 245296 22245 246073
rect 22287 245296 22297 246073
rect 22445 245296 22455 246073
rect 22497 245296 22507 246073
rect 22655 245296 22665 246073
rect 22707 245296 22717 246073
rect 22865 245296 22875 246073
rect 22917 245296 22927 246073
rect 23075 245296 23085 246073
rect 23127 245296 23137 246073
rect 23285 245296 23295 246073
rect 23337 245296 23347 246073
rect 23495 245296 23505 246073
rect 23547 245296 23557 246073
rect 23705 245296 23715 246073
rect 23757 245296 23767 246073
rect 23915 245296 23925 246073
rect 23967 245296 23977 246073
rect 24125 245296 24135 246073
rect 24177 245296 24187 246073
rect 24335 245296 24345 246073
rect 24387 245296 24397 246073
rect 24545 245296 24555 246073
rect 24597 245296 24607 246073
rect 24755 245296 24765 246073
rect 24807 245296 24817 246073
rect 24965 245296 24975 246073
rect 25017 245296 25027 246073
rect 25175 245296 25185 246073
rect 25227 245296 25237 246073
rect 25385 245296 25395 246073
rect 25437 245296 25447 246073
rect 25595 245296 25605 246073
rect 25647 245296 25657 246073
rect 25805 245296 25815 246073
rect 25857 245296 25867 246073
rect 26015 245296 26025 246073
rect 26067 245296 26077 246073
rect 26225 245296 26235 246073
rect 26277 245296 26287 246073
rect 26435 245296 26445 246073
rect 26487 245296 26497 246073
rect 26645 245296 26655 246073
rect 26697 245296 26707 246073
rect 26855 245296 26865 246073
rect 26907 245296 26917 246073
rect 27065 245296 27075 246073
rect 27117 245296 27127 246073
rect 27275 245296 27285 246073
rect 27331 246072 27566 246084
rect 27331 245296 27337 246072
rect 27371 245296 27566 246072
rect -4055 245284 -4009 245296
rect -3959 245284 -3913 245296
rect -3845 245284 -3799 245296
rect -3749 245284 -3703 245296
rect -3635 245284 -3589 245296
rect -3539 245284 -3493 245296
rect -3425 245284 -3379 245296
rect -3329 245284 -3283 245296
rect -3215 245284 -3169 245296
rect -3119 245284 -3073 245296
rect -3005 245284 -2959 245296
rect -2909 245284 -2863 245296
rect -2795 245284 -2749 245296
rect -2699 245284 -2653 245296
rect -2585 245284 -2539 245296
rect -2489 245284 -2443 245296
rect -2375 245284 -2329 245296
rect -2279 245284 -2233 245296
rect -2165 245284 -2119 245296
rect -2069 245284 -2023 245296
rect -1955 245284 -1909 245296
rect -1859 245284 -1813 245296
rect -1745 245284 -1699 245296
rect -1649 245284 -1603 245296
rect -1535 245284 -1489 245296
rect -1439 245284 -1393 245296
rect -1325 245284 -1279 245296
rect -1229 245284 -1183 245296
rect -1115 245284 -1069 245296
rect -1019 245284 -973 245296
rect -905 245284 -859 245296
rect -809 245284 -763 245296
rect -695 245284 -649 245296
rect -599 245284 -553 245296
rect -485 245284 -439 245296
rect -389 245284 -343 245296
rect -275 245284 -229 245296
rect -179 245284 -133 245296
rect -65 245284 -19 245296
rect 31 245284 77 245296
rect 145 245284 191 245296
rect 241 245284 287 245296
rect 355 245284 401 245296
rect 451 245284 497 245296
rect 565 245284 611 245296
rect 661 245284 707 245296
rect 775 245284 821 245296
rect 871 245284 917 245296
rect 985 245284 1031 245296
rect 1081 245284 1127 245296
rect 1195 245284 1241 245296
rect 1291 245284 1337 245296
rect 1405 245284 1451 245296
rect 1501 245284 1547 245296
rect 1615 245284 1661 245296
rect 1711 245284 1757 245296
rect 1825 245284 1871 245296
rect 1921 245284 1967 245296
rect 2035 245284 2081 245296
rect 2131 245284 2177 245296
rect 2245 245284 2291 245296
rect 2341 245284 2387 245296
rect 2455 245284 2501 245296
rect 2551 245284 2597 245296
rect 2665 245284 2711 245296
rect 2761 245284 2807 245296
rect 2875 245284 2921 245296
rect 2971 245284 3017 245296
rect 3085 245284 3131 245296
rect 3181 245284 3227 245296
rect 3295 245284 3341 245296
rect 3391 245284 3437 245296
rect 3505 245284 3551 245296
rect 3601 245284 3647 245296
rect 3715 245284 3761 245296
rect 3811 245284 3857 245296
rect 3925 245284 3971 245296
rect 4021 245284 4067 245296
rect 4135 245284 4181 245296
rect 4231 245284 4277 245296
rect 4345 245284 4391 245296
rect 4441 245284 4487 245296
rect 4555 245284 4601 245296
rect 4651 245284 4697 245296
rect 4765 245284 4811 245296
rect 4861 245284 4907 245296
rect 4975 245284 5021 245296
rect 5071 245284 5117 245296
rect 5185 245284 5231 245296
rect 5281 245284 5327 245296
rect 5395 245284 5441 245296
rect 5491 245284 5537 245296
rect 5605 245284 5651 245296
rect 5701 245284 5747 245296
rect 5815 245284 5861 245296
rect 5911 245284 5957 245296
rect 6025 245284 6071 245296
rect 6121 245284 6167 245296
rect 6235 245284 6281 245296
rect 6331 245284 6377 245296
rect 6445 245284 6491 245296
rect 6541 245284 6587 245296
rect 6655 245284 6701 245296
rect 6751 245284 6797 245296
rect 6865 245284 6911 245296
rect 6961 245284 7007 245296
rect 7075 245284 7121 245296
rect 7171 245284 7217 245296
rect 7285 245284 7331 245296
rect 7381 245284 7427 245296
rect 7495 245284 7541 245296
rect 7591 245284 7637 245296
rect 7705 245284 7751 245296
rect 7801 245284 7847 245296
rect 7915 245284 7961 245296
rect 8011 245284 8057 245296
rect 8125 245284 8171 245296
rect 8221 245284 8267 245296
rect 8335 245284 8381 245296
rect 8431 245284 8477 245296
rect 8545 245284 8591 245296
rect 8641 245284 8687 245296
rect 8755 245284 8801 245296
rect 8851 245284 8897 245296
rect 8965 245284 9011 245296
rect 9061 245284 9107 245296
rect 9175 245284 9221 245296
rect 9271 245284 9317 245296
rect 9385 245284 9431 245296
rect 9481 245284 9527 245296
rect 9595 245284 9641 245296
rect 9691 245284 9737 245296
rect 9805 245284 9851 245296
rect 9901 245284 9947 245296
rect 10015 245284 10061 245296
rect 10111 245284 10157 245296
rect 10225 245284 10271 245296
rect 10321 245284 10367 245296
rect 10435 245284 10481 245296
rect 10531 245284 10577 245296
rect 10645 245284 10691 245296
rect 10741 245284 10787 245296
rect 10855 245284 10901 245296
rect 10951 245284 10997 245296
rect 11065 245284 11111 245296
rect 11161 245284 11207 245296
rect 11275 245284 11321 245296
rect 11371 245284 11417 245296
rect 11485 245284 11531 245296
rect 11581 245284 11627 245296
rect 11695 245284 11741 245296
rect 11791 245284 11837 245296
rect 11905 245284 11951 245296
rect 12001 245284 12047 245296
rect 12115 245284 12161 245296
rect 12211 245284 12257 245296
rect 12325 245284 12371 245296
rect 12421 245284 12467 245296
rect 12535 245284 12581 245296
rect 12631 245284 12677 245296
rect 12745 245284 12791 245296
rect 12841 245284 12887 245296
rect 12955 245284 13001 245296
rect 13051 245284 13097 245296
rect 13165 245284 13211 245296
rect 13261 245284 13307 245296
rect 13375 245284 13421 245296
rect 13471 245284 13517 245296
rect 13585 245284 13631 245296
rect 13681 245284 13727 245296
rect 13795 245284 13841 245296
rect 13891 245284 13937 245296
rect 14005 245284 14051 245296
rect 14101 245284 14147 245296
rect 14215 245284 14261 245296
rect 14311 245284 14357 245296
rect 14425 245284 14471 245296
rect 14521 245284 14567 245296
rect 14635 245284 14681 245296
rect 14731 245284 14777 245296
rect 14845 245284 14891 245296
rect 14941 245284 14987 245296
rect 15055 245284 15101 245296
rect 15151 245284 15197 245296
rect 15265 245284 15311 245296
rect 15361 245284 15407 245296
rect 15475 245284 15521 245296
rect 15571 245284 15617 245296
rect 15685 245284 15731 245296
rect 15781 245284 15827 245296
rect 15895 245284 15941 245296
rect 15991 245284 16037 245296
rect 16105 245284 16151 245296
rect 16201 245284 16247 245296
rect 16315 245284 16361 245296
rect 16411 245284 16457 245296
rect 16525 245284 16571 245296
rect 16621 245284 16667 245296
rect 16735 245284 16781 245296
rect 16831 245284 16877 245296
rect 16945 245284 16991 245296
rect 17041 245284 17087 245296
rect 17155 245284 17201 245296
rect 17251 245284 17297 245296
rect 17365 245284 17411 245296
rect 17461 245284 17507 245296
rect 17575 245284 17621 245296
rect 17671 245284 17717 245296
rect 17785 245284 17831 245296
rect 17881 245284 17927 245296
rect 17995 245284 18041 245296
rect 18091 245284 18137 245296
rect 18205 245284 18251 245296
rect 18301 245284 18347 245296
rect 18415 245284 18461 245296
rect 18511 245284 18557 245296
rect 18625 245284 18671 245296
rect 18721 245284 18767 245296
rect 18835 245284 18881 245296
rect 18931 245284 18977 245296
rect 19045 245284 19091 245296
rect 19141 245284 19187 245296
rect 19255 245284 19301 245296
rect 19351 245284 19397 245296
rect 19465 245284 19511 245296
rect 19561 245284 19607 245296
rect 19675 245284 19721 245296
rect 19771 245284 19817 245296
rect 19885 245284 19931 245296
rect 19981 245284 20027 245296
rect 20095 245284 20141 245296
rect 20191 245284 20237 245296
rect 20305 245284 20351 245296
rect 20401 245284 20447 245296
rect 20515 245284 20561 245296
rect 20611 245284 20657 245296
rect 20725 245284 20771 245296
rect 20821 245284 20867 245296
rect 20935 245284 20981 245296
rect 21031 245284 21077 245296
rect 21145 245284 21191 245296
rect 21241 245284 21287 245296
rect 21355 245284 21401 245296
rect 21451 245284 21497 245296
rect 21565 245284 21611 245296
rect 21661 245284 21707 245296
rect 21775 245284 21821 245296
rect 21871 245284 21917 245296
rect 21985 245284 22031 245296
rect 22081 245284 22127 245296
rect 22195 245284 22241 245296
rect 22291 245284 22337 245296
rect 22405 245284 22451 245296
rect 22501 245284 22547 245296
rect 22615 245284 22661 245296
rect 22711 245284 22757 245296
rect 22825 245284 22871 245296
rect 22921 245284 22967 245296
rect 23035 245284 23081 245296
rect 23131 245284 23177 245296
rect 23245 245284 23291 245296
rect 23341 245284 23387 245296
rect 23455 245284 23501 245296
rect 23551 245284 23597 245296
rect 23665 245284 23711 245296
rect 23761 245284 23807 245296
rect 23875 245284 23921 245296
rect 23971 245284 24017 245296
rect 24085 245284 24131 245296
rect 24181 245284 24227 245296
rect 24295 245284 24341 245296
rect 24391 245284 24437 245296
rect 24505 245284 24551 245296
rect 24601 245284 24647 245296
rect 24715 245284 24761 245296
rect 24811 245284 24857 245296
rect 24925 245284 24971 245296
rect 25021 245284 25067 245296
rect 25135 245284 25181 245296
rect 25231 245284 25277 245296
rect 25345 245284 25391 245296
rect 25441 245284 25487 245296
rect 25555 245284 25601 245296
rect 25651 245284 25697 245296
rect 25765 245284 25811 245296
rect 25861 245284 25907 245296
rect 25975 245284 26021 245296
rect 26071 245284 26117 245296
rect 26185 245284 26231 245296
rect 26281 245284 26327 245296
rect 26395 245284 26441 245296
rect 26491 245284 26537 245296
rect 26605 245284 26651 245296
rect 26701 245284 26747 245296
rect 26815 245284 26861 245296
rect 26911 245284 26957 245296
rect 27025 245284 27071 245296
rect 27121 245284 27167 245296
rect 27235 245284 27281 245296
rect 27331 245284 27566 245296
rect -4013 245237 27125 245249
rect -5008 245095 -4001 245237
rect -3967 245095 -3581 245237
rect -3547 245095 -3161 245237
rect -3127 245095 -2741 245237
rect -2707 245095 -2321 245237
rect -2287 245095 -1901 245237
rect -1867 245095 -1481 245237
rect -1447 245095 -1061 245237
rect -1027 245095 -641 245237
rect -607 245095 -221 245237
rect -187 245095 199 245237
rect 233 245095 619 245237
rect 653 245095 1039 245237
rect 1073 245095 1459 245237
rect 1493 245095 1879 245237
rect 1913 245095 2299 245237
rect 2333 245095 2719 245237
rect 2753 245095 3139 245237
rect 3173 245095 3559 245237
rect 3593 245095 3979 245237
rect 4013 245095 4399 245237
rect 4433 245095 4819 245237
rect 4853 245095 5239 245237
rect 5273 245095 5659 245237
rect 5693 245095 6079 245237
rect 6113 245095 6499 245237
rect 6533 245095 6919 245237
rect 6953 245095 7339 245237
rect 7373 245095 7759 245237
rect 7793 245095 8179 245237
rect 8213 245095 8599 245237
rect 8633 245095 9019 245237
rect 9053 245095 9439 245237
rect 9473 245095 9859 245237
rect 9893 245095 10279 245237
rect 10313 245095 10699 245237
rect 10733 245095 11119 245237
rect 11153 245095 11539 245237
rect 11573 245095 11959 245237
rect 11993 245095 12379 245237
rect 12413 245095 12799 245237
rect 12833 245095 13219 245237
rect 13253 245095 13639 245237
rect 13673 245095 14059 245237
rect 14093 245095 14479 245237
rect 14513 245095 14899 245237
rect 14933 245095 15319 245237
rect 15353 245095 15739 245237
rect 15773 245095 16159 245237
rect 16193 245095 16579 245237
rect 16613 245095 16999 245237
rect 17033 245095 17419 245237
rect 17453 245095 17839 245237
rect 17873 245095 18259 245237
rect 18293 245095 18679 245237
rect 18713 245095 19099 245237
rect 19133 245095 19519 245237
rect 19553 245095 19939 245237
rect 19973 245095 20359 245237
rect 20393 245095 20779 245237
rect 20813 245095 21199 245237
rect 21233 245095 21619 245237
rect 21653 245095 22039 245237
rect 22073 245095 22459 245237
rect 22493 245095 22879 245237
rect 22913 245095 23299 245237
rect 23333 245095 23719 245237
rect 23753 245095 24139 245237
rect 24173 245095 24559 245237
rect 24593 245095 24979 245237
rect 25013 245095 25399 245237
rect 25433 245095 25819 245237
rect 25853 245095 26239 245237
rect 26273 245095 26659 245237
rect 26693 245095 27079 245237
rect 27113 245095 27125 245237
rect -5008 244207 -4142 245095
rect -4013 245083 27125 245095
rect 27377 245048 27566 245284
rect -4056 245036 -4009 245048
rect -3959 245036 -3913 245048
rect -3845 245036 -3799 245048
rect -3749 245036 -3703 245048
rect -3635 245036 -3589 245048
rect -3539 245037 -3493 245048
rect -3425 245037 -3379 245048
rect -3329 245037 -3283 245048
rect -3215 245037 -3169 245048
rect -3119 245037 -3073 245048
rect -3005 245037 -2959 245048
rect -2909 245037 -2863 245048
rect -2795 245037 -2749 245048
rect -2699 245037 -2653 245048
rect -2585 245037 -2539 245048
rect -2489 245037 -2443 245048
rect -2375 245037 -2329 245048
rect -2279 245037 -2233 245048
rect -2165 245037 -2119 245048
rect -2069 245037 -2023 245048
rect -1955 245037 -1909 245048
rect -1859 245037 -1813 245048
rect -1745 245037 -1699 245048
rect -1649 245037 -1603 245048
rect -1535 245037 -1489 245048
rect -1439 245037 -1393 245048
rect -1325 245037 -1279 245048
rect -1229 245037 -1183 245048
rect -1115 245037 -1069 245048
rect -1019 245037 -973 245048
rect -905 245037 -859 245048
rect -809 245037 -763 245048
rect -695 245037 -649 245048
rect -599 245037 -553 245048
rect -485 245037 -439 245048
rect -389 245037 -343 245048
rect -275 245037 -229 245048
rect -179 245037 -133 245048
rect -65 245037 -19 245048
rect 31 245037 77 245048
rect 145 245037 191 245048
rect 241 245037 287 245048
rect 355 245037 401 245048
rect 451 245037 497 245048
rect 565 245037 611 245048
rect 661 245037 707 245048
rect 775 245037 821 245048
rect 871 245037 917 245048
rect 985 245037 1031 245048
rect 1081 245037 1127 245048
rect 1195 245037 1241 245048
rect 1291 245037 1337 245048
rect 1405 245037 1451 245048
rect 1501 245037 1547 245048
rect 1615 245037 1661 245048
rect 1711 245037 1757 245048
rect 1825 245037 1871 245048
rect 1921 245037 1967 245048
rect 2035 245037 2081 245048
rect 2131 245037 2177 245048
rect 2245 245037 2291 245048
rect 2341 245037 2387 245048
rect 2455 245037 2501 245048
rect 2551 245037 2597 245048
rect 2665 245037 2711 245048
rect 2761 245037 2807 245048
rect 2875 245037 2921 245048
rect 2971 245037 3017 245048
rect 3085 245037 3131 245048
rect 3181 245037 3227 245048
rect 3295 245037 3341 245048
rect 3391 245037 3437 245048
rect 3505 245037 3551 245048
rect 3601 245037 3647 245048
rect 3715 245037 3761 245048
rect 3811 245037 3857 245048
rect 3925 245037 3971 245048
rect 4021 245037 4067 245048
rect 4135 245037 4181 245048
rect 4231 245037 4277 245048
rect 4345 245037 4391 245048
rect 4441 245037 4487 245048
rect 4555 245037 4601 245048
rect 4651 245037 4697 245048
rect 4765 245037 4811 245048
rect 4861 245037 4907 245048
rect 4975 245037 5021 245048
rect 5071 245037 5117 245048
rect 5185 245037 5231 245048
rect 5281 245037 5327 245048
rect 5395 245037 5441 245048
rect 5491 245037 5537 245048
rect 5605 245037 5651 245048
rect 5701 245037 5747 245048
rect 5815 245037 5861 245048
rect 5911 245037 5957 245048
rect 6025 245037 6071 245048
rect 6121 245037 6167 245048
rect 6235 245037 6281 245048
rect 6331 245037 6377 245048
rect 6445 245037 6491 245048
rect 6541 245037 6587 245048
rect 6655 245037 6701 245048
rect 6751 245037 6797 245048
rect 6865 245037 6911 245048
rect 6961 245037 7007 245048
rect 7075 245037 7121 245048
rect 7171 245037 7217 245048
rect 7285 245037 7331 245048
rect 7381 245037 7427 245048
rect 7495 245037 7541 245048
rect 7591 245037 7637 245048
rect 7705 245037 7751 245048
rect 7801 245037 7847 245048
rect 7915 245037 7961 245048
rect 8011 245037 8057 245048
rect 8125 245037 8171 245048
rect 8221 245037 8267 245048
rect 8335 245037 8381 245048
rect 8431 245037 8477 245048
rect 8545 245037 8591 245048
rect 8641 245037 8687 245048
rect 8755 245037 8801 245048
rect 8851 245037 8897 245048
rect 8965 245037 9011 245048
rect 9061 245037 9107 245048
rect 9175 245037 9221 245048
rect 9271 245037 9317 245048
rect 9385 245037 9431 245048
rect 9481 245037 9527 245048
rect 9595 245037 9641 245048
rect 9691 245037 9737 245048
rect 9805 245037 9851 245048
rect 9901 245037 9947 245048
rect 10015 245037 10061 245048
rect 10111 245037 10157 245048
rect 10225 245037 10271 245048
rect 10321 245037 10367 245048
rect 10435 245037 10481 245048
rect 10531 245037 10577 245048
rect 10645 245037 10691 245048
rect 10741 245037 10787 245048
rect 10855 245037 10901 245048
rect 10951 245037 10997 245048
rect 11065 245037 11111 245048
rect 11161 245037 11207 245048
rect 11275 245037 11321 245048
rect 11371 245037 11417 245048
rect 11485 245037 11531 245048
rect 11581 245037 11627 245048
rect 11695 245037 11741 245048
rect 11791 245037 11837 245048
rect 11905 245037 11951 245048
rect 12001 245037 12047 245048
rect 12115 245037 12161 245048
rect 12211 245037 12257 245048
rect 12325 245037 12371 245048
rect 12421 245037 12467 245048
rect 12535 245037 12581 245048
rect 12631 245037 12677 245048
rect 12745 245037 12791 245048
rect 12841 245037 12887 245048
rect 12955 245037 13001 245048
rect 13051 245037 13097 245048
rect 13165 245037 13211 245048
rect 13261 245037 13307 245048
rect 13375 245037 13421 245048
rect 13471 245037 13517 245048
rect 13585 245037 13631 245048
rect 13681 245037 13727 245048
rect 13795 245037 13841 245048
rect 13891 245037 13937 245048
rect 14005 245037 14051 245048
rect 14101 245037 14147 245048
rect 14215 245037 14261 245048
rect 14311 245037 14357 245048
rect 14425 245037 14471 245048
rect 14521 245037 14567 245048
rect 14635 245037 14681 245048
rect 14731 245037 14777 245048
rect 14845 245037 14891 245048
rect 14941 245037 14987 245048
rect 15055 245037 15101 245048
rect 15151 245037 15197 245048
rect 15265 245037 15311 245048
rect 15361 245037 15407 245048
rect 15475 245037 15521 245048
rect 15571 245037 15617 245048
rect 15685 245037 15731 245048
rect 15781 245037 15827 245048
rect 15895 245037 15941 245048
rect 15991 245037 16037 245048
rect 16105 245037 16151 245048
rect 16201 245037 16247 245048
rect 16315 245037 16361 245048
rect 16411 245037 16457 245048
rect 16525 245037 16571 245048
rect 16621 245037 16667 245048
rect 16735 245037 16781 245048
rect 16831 245037 16877 245048
rect 16945 245037 16991 245048
rect 17041 245037 17087 245048
rect 17155 245037 17201 245048
rect 17251 245037 17297 245048
rect 17365 245037 17411 245048
rect 17461 245037 17507 245048
rect 17575 245037 17621 245048
rect 17671 245037 17717 245048
rect 17785 245037 17831 245048
rect 17881 245037 17927 245048
rect 17995 245037 18041 245048
rect 18091 245037 18137 245048
rect 18205 245037 18251 245048
rect 18301 245037 18347 245048
rect 18415 245037 18461 245048
rect 18511 245037 18557 245048
rect 18625 245037 18671 245048
rect 18721 245037 18767 245048
rect 18835 245037 18881 245048
rect 18931 245037 18977 245048
rect 19045 245037 19091 245048
rect 19141 245037 19187 245048
rect 19255 245037 19301 245048
rect 19351 245037 19397 245048
rect 19465 245037 19511 245048
rect 19561 245037 19607 245048
rect 19675 245037 19721 245048
rect 19771 245037 19817 245048
rect 19885 245037 19931 245048
rect 19981 245037 20027 245048
rect 20095 245037 20141 245048
rect 20191 245037 20237 245048
rect 20305 245037 20351 245048
rect 20401 245037 20447 245048
rect 20515 245037 20561 245048
rect 20611 245037 20657 245048
rect 20725 245037 20771 245048
rect 20821 245037 20867 245048
rect 20935 245037 20981 245048
rect 21031 245037 21077 245048
rect 21145 245037 21191 245048
rect 21241 245037 21287 245048
rect 21355 245037 21401 245048
rect 21451 245037 21497 245048
rect 21565 245037 21611 245048
rect 21661 245037 21707 245048
rect 21775 245037 21821 245048
rect 21871 245037 21917 245048
rect 21985 245037 22031 245048
rect 22081 245037 22127 245048
rect 22195 245037 22241 245048
rect 22291 245037 22337 245048
rect 22405 245037 22451 245048
rect 22501 245037 22547 245048
rect 22615 245037 22661 245048
rect 22711 245037 22757 245048
rect 22825 245037 22871 245048
rect 22921 245037 22967 245048
rect 23035 245037 23081 245048
rect 23131 245037 23177 245048
rect 23245 245037 23291 245048
rect 23341 245037 23387 245048
rect 23455 245037 23501 245048
rect 23551 245037 23597 245048
rect 23665 245037 23711 245048
rect 23761 245037 23807 245048
rect 23875 245037 23921 245048
rect 23971 245037 24017 245048
rect 24085 245037 24131 245048
rect 24181 245037 24227 245048
rect 24295 245037 24341 245048
rect 24391 245037 24437 245048
rect 24505 245037 24551 245048
rect 24601 245037 24647 245048
rect 24715 245037 24761 245048
rect 24811 245037 24857 245048
rect 24925 245037 24971 245048
rect 25021 245037 25067 245048
rect 25135 245037 25181 245048
rect 25231 245037 25277 245048
rect 25345 245037 25391 245048
rect 25441 245037 25487 245048
rect 25555 245037 25601 245048
rect 25651 245037 25697 245048
rect 25765 245037 25811 245048
rect 25861 245037 25907 245048
rect 25975 245037 26021 245048
rect 26071 245037 26117 245048
rect 26185 245037 26231 245048
rect 26281 245037 26327 245048
rect 26395 245037 26441 245048
rect 26491 245037 26537 245048
rect 26605 245037 26651 245048
rect 26701 245037 26747 245048
rect 26815 245037 26861 245048
rect 26911 245037 26957 245048
rect 27025 245037 27071 245048
rect 27121 245037 27167 245048
rect 27235 245037 27281 245048
rect -4085 244260 -4075 245036
rect -4015 244260 -4005 245036
rect -3963 244260 -3953 245036
rect -3805 244260 -3795 245036
rect -3753 244260 -3743 245036
rect -3595 244260 -3585 245036
rect -3543 244260 -3533 245037
rect -3385 244260 -3375 245037
rect -3333 244260 -3323 245037
rect -3175 244260 -3165 245037
rect -3123 244260 -3113 245037
rect -2965 244260 -2955 245037
rect -2913 244260 -2903 245037
rect -2755 244260 -2745 245037
rect -2703 244260 -2693 245037
rect -2545 244260 -2535 245037
rect -2493 244260 -2483 245037
rect -2335 244260 -2325 245037
rect -2283 244260 -2273 245037
rect -2125 244260 -2115 245037
rect -2073 244260 -2063 245037
rect -1915 244260 -1905 245037
rect -1863 244260 -1853 245037
rect -1705 244260 -1695 245037
rect -1653 244260 -1643 245037
rect -1495 244260 -1485 245037
rect -1443 244260 -1433 245037
rect -1285 244260 -1275 245037
rect -1233 244260 -1223 245037
rect -1075 244260 -1065 245037
rect -1023 244260 -1013 245037
rect -865 244260 -855 245037
rect -813 244260 -803 245037
rect -655 244260 -645 245037
rect -603 244260 -593 245037
rect -445 244260 -435 245037
rect -393 244260 -383 245037
rect -235 244260 -225 245037
rect -183 244260 -173 245037
rect -25 244260 -15 245037
rect 27 244260 37 245037
rect 185 244260 195 245037
rect 237 244260 247 245037
rect 395 244260 405 245037
rect 447 244260 457 245037
rect 605 244260 615 245037
rect 657 244260 667 245037
rect 815 244260 825 245037
rect 867 244260 877 245037
rect 1025 244260 1035 245037
rect 1077 244260 1087 245037
rect 1235 244260 1245 245037
rect 1287 244260 1297 245037
rect 1445 244260 1455 245037
rect 1497 244260 1507 245037
rect 1655 244260 1665 245037
rect 1707 244260 1717 245037
rect 1865 244260 1875 245037
rect 1917 244260 1927 245037
rect 2075 244260 2085 245037
rect 2127 244260 2137 245037
rect 2285 244260 2295 245037
rect 2337 244260 2347 245037
rect 2495 244260 2505 245037
rect 2547 244260 2557 245037
rect 2705 244260 2715 245037
rect 2757 244260 2767 245037
rect 2915 244260 2925 245037
rect 2967 244260 2977 245037
rect 3125 244260 3135 245037
rect 3177 244260 3187 245037
rect 3335 244260 3345 245037
rect 3387 244260 3397 245037
rect 3545 244260 3555 245037
rect 3597 244260 3607 245037
rect 3755 244260 3765 245037
rect 3807 244260 3817 245037
rect 3965 244260 3975 245037
rect 4017 244260 4027 245037
rect 4175 244260 4185 245037
rect 4227 244260 4237 245037
rect 4385 244260 4395 245037
rect 4437 244260 4447 245037
rect 4595 244260 4605 245037
rect 4647 244260 4657 245037
rect 4805 244260 4815 245037
rect 4857 244260 4867 245037
rect 5015 244260 5025 245037
rect 5067 244260 5077 245037
rect 5225 244260 5235 245037
rect 5277 244260 5287 245037
rect 5435 244260 5445 245037
rect 5487 244260 5497 245037
rect 5645 244260 5655 245037
rect 5697 244260 5707 245037
rect 5855 244260 5865 245037
rect 5907 244260 5917 245037
rect 6065 244260 6075 245037
rect 6117 244260 6127 245037
rect 6275 244260 6285 245037
rect 6327 244260 6337 245037
rect 6485 244260 6495 245037
rect 6537 244260 6547 245037
rect 6695 244260 6705 245037
rect 6747 244260 6757 245037
rect 6905 244260 6915 245037
rect 6957 244260 6967 245037
rect 7115 244260 7125 245037
rect 7167 244260 7177 245037
rect 7325 244260 7335 245037
rect 7377 244260 7387 245037
rect 7535 244260 7545 245037
rect 7587 244260 7597 245037
rect 7745 244260 7755 245037
rect 7797 244260 7807 245037
rect 7955 244260 7965 245037
rect 8007 244260 8017 245037
rect 8165 244260 8175 245037
rect 8217 244260 8227 245037
rect 8375 244260 8385 245037
rect 8427 244260 8437 245037
rect 8585 244260 8595 245037
rect 8637 244260 8647 245037
rect 8795 244260 8805 245037
rect 8847 244260 8857 245037
rect 9005 244260 9015 245037
rect 9057 244260 9067 245037
rect 9215 244260 9225 245037
rect 9267 244260 9277 245037
rect 9425 244260 9435 245037
rect 9477 244260 9487 245037
rect 9635 244260 9645 245037
rect 9687 244260 9697 245037
rect 9845 244260 9855 245037
rect 9897 244260 9907 245037
rect 10055 244260 10065 245037
rect 10107 244260 10117 245037
rect 10265 244260 10275 245037
rect 10317 244260 10327 245037
rect 10475 244260 10485 245037
rect 10527 244260 10537 245037
rect 10685 244260 10695 245037
rect 10737 244260 10747 245037
rect 10895 244260 10905 245037
rect 10947 244260 10957 245037
rect 11105 244260 11115 245037
rect 11157 244260 11167 245037
rect 11315 244260 11325 245037
rect 11367 244260 11377 245037
rect 11525 244260 11535 245037
rect 11577 244260 11587 245037
rect 11735 244260 11745 245037
rect 11787 244260 11797 245037
rect 11945 244260 11955 245037
rect 11997 244260 12007 245037
rect 12155 244260 12165 245037
rect 12207 244260 12217 245037
rect 12365 244260 12375 245037
rect 12417 244260 12427 245037
rect 12575 244260 12585 245037
rect 12627 244260 12637 245037
rect 12785 244260 12795 245037
rect 12837 244260 12847 245037
rect 12995 244260 13005 245037
rect 13047 244260 13057 245037
rect 13205 244260 13215 245037
rect 13257 244260 13267 245037
rect 13415 244260 13425 245037
rect 13467 244260 13477 245037
rect 13625 244260 13635 245037
rect 13677 244260 13687 245037
rect 13835 244260 13845 245037
rect 13887 244260 13897 245037
rect 14045 244260 14055 245037
rect 14097 244260 14107 245037
rect 14255 244260 14265 245037
rect 14307 244260 14317 245037
rect 14465 244260 14475 245037
rect 14517 244260 14527 245037
rect 14675 244260 14685 245037
rect 14727 244260 14737 245037
rect 14885 244260 14895 245037
rect 14937 244260 14947 245037
rect 15095 244260 15105 245037
rect 15147 244260 15157 245037
rect 15305 244260 15315 245037
rect 15357 244260 15367 245037
rect 15515 244260 15525 245037
rect 15567 244260 15577 245037
rect 15725 244260 15735 245037
rect 15777 244260 15787 245037
rect 15935 244260 15945 245037
rect 15987 244260 15997 245037
rect 16145 244260 16155 245037
rect 16197 244260 16207 245037
rect 16355 244260 16365 245037
rect 16407 244260 16417 245037
rect 16565 244260 16575 245037
rect 16617 244260 16627 245037
rect 16775 244260 16785 245037
rect 16827 244260 16837 245037
rect 16985 244260 16995 245037
rect 17037 244260 17047 245037
rect 17195 244260 17205 245037
rect 17247 244260 17257 245037
rect 17405 244260 17415 245037
rect 17457 244260 17467 245037
rect 17615 244260 17625 245037
rect 17667 244260 17677 245037
rect 17825 244260 17835 245037
rect 17877 244260 17887 245037
rect 18035 244260 18045 245037
rect 18087 244260 18097 245037
rect 18245 244260 18255 245037
rect 18297 244260 18307 245037
rect 18455 244260 18465 245037
rect 18507 244260 18517 245037
rect 18665 244260 18675 245037
rect 18717 244260 18727 245037
rect 18875 244260 18885 245037
rect 18927 244260 18937 245037
rect 19085 244260 19095 245037
rect 19137 244260 19147 245037
rect 19295 244260 19305 245037
rect 19347 244260 19357 245037
rect 19505 244260 19515 245037
rect 19557 244260 19567 245037
rect 19715 244260 19725 245037
rect 19767 244260 19777 245037
rect 19925 244260 19935 245037
rect 19977 244260 19987 245037
rect 20135 244260 20145 245037
rect 20187 244260 20197 245037
rect 20345 244260 20355 245037
rect 20397 244260 20407 245037
rect 20555 244260 20565 245037
rect 20607 244260 20617 245037
rect 20765 244260 20775 245037
rect 20817 244260 20827 245037
rect 20975 244260 20985 245037
rect 21027 244260 21037 245037
rect 21185 244260 21195 245037
rect 21237 244260 21247 245037
rect 21395 244260 21405 245037
rect 21447 244260 21457 245037
rect 21605 244260 21615 245037
rect 21657 244260 21667 245037
rect 21815 244260 21825 245037
rect 21867 244260 21877 245037
rect 22025 244260 22035 245037
rect 22077 244260 22087 245037
rect 22235 244260 22245 245037
rect 22287 244260 22297 245037
rect 22445 244260 22455 245037
rect 22497 244260 22507 245037
rect 22655 244260 22665 245037
rect 22707 244260 22717 245037
rect 22865 244260 22875 245037
rect 22917 244260 22927 245037
rect 23075 244260 23085 245037
rect 23127 244260 23137 245037
rect 23285 244260 23295 245037
rect 23337 244260 23347 245037
rect 23495 244260 23505 245037
rect 23547 244260 23557 245037
rect 23705 244260 23715 245037
rect 23757 244260 23767 245037
rect 23915 244260 23925 245037
rect 23967 244260 23977 245037
rect 24125 244260 24135 245037
rect 24177 244260 24187 245037
rect 24335 244260 24345 245037
rect 24387 244260 24397 245037
rect 24545 244260 24555 245037
rect 24597 244260 24607 245037
rect 24755 244260 24765 245037
rect 24807 244260 24817 245037
rect 24965 244260 24975 245037
rect 25017 244260 25027 245037
rect 25175 244260 25185 245037
rect 25227 244260 25237 245037
rect 25385 244260 25395 245037
rect 25437 244260 25447 245037
rect 25595 244260 25605 245037
rect 25647 244260 25657 245037
rect 25805 244260 25815 245037
rect 25857 244260 25867 245037
rect 26015 244260 26025 245037
rect 26067 244260 26077 245037
rect 26225 244260 26235 245037
rect 26277 244260 26287 245037
rect 26435 244260 26445 245037
rect 26487 244260 26497 245037
rect 26645 244260 26655 245037
rect 26697 244260 26707 245037
rect 26855 244260 26865 245037
rect 26907 244260 26917 245037
rect 27065 244260 27075 245037
rect 27117 244260 27127 245037
rect 27275 244260 27285 245037
rect 27331 245036 27566 245048
rect 27331 244260 27337 245036
rect 27371 244260 27566 245036
rect -4056 244248 -4009 244260
rect -3959 244248 -3913 244260
rect -3845 244248 -3799 244260
rect -3749 244248 -3703 244260
rect -3635 244248 -3589 244260
rect -3539 244248 -3493 244260
rect -3425 244248 -3379 244260
rect -3329 244248 -3283 244260
rect -3215 244248 -3169 244260
rect -3119 244248 -3073 244260
rect -3005 244248 -2959 244260
rect -2909 244248 -2863 244260
rect -2795 244248 -2749 244260
rect -2699 244248 -2653 244260
rect -2585 244248 -2539 244260
rect -2489 244248 -2443 244260
rect -2375 244248 -2329 244260
rect -2279 244248 -2233 244260
rect -2165 244248 -2119 244260
rect -2069 244248 -2023 244260
rect -1955 244248 -1909 244260
rect -1859 244248 -1813 244260
rect -1745 244248 -1699 244260
rect -1649 244248 -1603 244260
rect -1535 244248 -1489 244260
rect -1439 244248 -1393 244260
rect -1325 244248 -1279 244260
rect -1229 244248 -1183 244260
rect -1115 244248 -1069 244260
rect -1019 244248 -973 244260
rect -905 244248 -859 244260
rect -809 244248 -763 244260
rect -695 244248 -649 244260
rect -599 244248 -553 244260
rect -485 244248 -439 244260
rect -389 244248 -343 244260
rect -275 244248 -229 244260
rect -179 244248 -133 244260
rect -65 244248 -19 244260
rect 31 244248 77 244260
rect 145 244248 191 244260
rect 241 244248 287 244260
rect 355 244248 401 244260
rect 451 244248 497 244260
rect 565 244248 611 244260
rect 661 244248 707 244260
rect 775 244248 821 244260
rect 871 244248 917 244260
rect 985 244248 1031 244260
rect 1081 244248 1127 244260
rect 1195 244248 1241 244260
rect 1291 244248 1337 244260
rect 1405 244248 1451 244260
rect 1501 244248 1547 244260
rect 1615 244248 1661 244260
rect 1711 244248 1757 244260
rect 1825 244248 1871 244260
rect 1921 244248 1967 244260
rect 2035 244248 2081 244260
rect 2131 244248 2177 244260
rect 2245 244248 2291 244260
rect 2341 244248 2387 244260
rect 2455 244248 2501 244260
rect 2551 244248 2597 244260
rect 2665 244248 2711 244260
rect 2761 244248 2807 244260
rect 2875 244248 2921 244260
rect 2971 244248 3017 244260
rect 3085 244248 3131 244260
rect 3181 244248 3227 244260
rect 3295 244248 3341 244260
rect 3391 244248 3437 244260
rect 3505 244248 3551 244260
rect 3601 244248 3647 244260
rect 3715 244248 3761 244260
rect 3811 244248 3857 244260
rect 3925 244248 3971 244260
rect 4021 244248 4067 244260
rect 4135 244248 4181 244260
rect 4231 244248 4277 244260
rect 4345 244248 4391 244260
rect 4441 244248 4487 244260
rect 4555 244248 4601 244260
rect 4651 244248 4697 244260
rect 4765 244248 4811 244260
rect 4861 244248 4907 244260
rect 4975 244248 5021 244260
rect 5071 244248 5117 244260
rect 5185 244248 5231 244260
rect 5281 244248 5327 244260
rect 5395 244248 5441 244260
rect 5491 244248 5537 244260
rect 5605 244248 5651 244260
rect 5701 244248 5747 244260
rect 5815 244248 5861 244260
rect 5911 244248 5957 244260
rect 6025 244248 6071 244260
rect 6121 244248 6167 244260
rect 6235 244248 6281 244260
rect 6331 244248 6377 244260
rect 6445 244248 6491 244260
rect 6541 244248 6587 244260
rect 6655 244248 6701 244260
rect 6751 244248 6797 244260
rect 6865 244248 6911 244260
rect 6961 244248 7007 244260
rect 7075 244248 7121 244260
rect 7171 244248 7217 244260
rect 7285 244248 7331 244260
rect 7381 244248 7427 244260
rect 7495 244248 7541 244260
rect 7591 244248 7637 244260
rect 7705 244248 7751 244260
rect 7801 244248 7847 244260
rect 7915 244248 7961 244260
rect 8011 244248 8057 244260
rect 8125 244248 8171 244260
rect 8221 244248 8267 244260
rect 8335 244248 8381 244260
rect 8431 244248 8477 244260
rect 8545 244248 8591 244260
rect 8641 244248 8687 244260
rect 8755 244248 8801 244260
rect 8851 244248 8897 244260
rect 8965 244248 9011 244260
rect 9061 244248 9107 244260
rect 9175 244248 9221 244260
rect 9271 244248 9317 244260
rect 9385 244248 9431 244260
rect 9481 244248 9527 244260
rect 9595 244248 9641 244260
rect 9691 244248 9737 244260
rect 9805 244248 9851 244260
rect 9901 244248 9947 244260
rect 10015 244248 10061 244260
rect 10111 244248 10157 244260
rect 10225 244248 10271 244260
rect 10321 244248 10367 244260
rect 10435 244248 10481 244260
rect 10531 244248 10577 244260
rect 10645 244248 10691 244260
rect 10741 244248 10787 244260
rect 10855 244248 10901 244260
rect 10951 244248 10997 244260
rect 11065 244248 11111 244260
rect 11161 244248 11207 244260
rect 11275 244248 11321 244260
rect 11371 244248 11417 244260
rect 11485 244248 11531 244260
rect 11581 244248 11627 244260
rect 11695 244248 11741 244260
rect 11791 244248 11837 244260
rect 11905 244248 11951 244260
rect 12001 244248 12047 244260
rect 12115 244248 12161 244260
rect 12211 244248 12257 244260
rect 12325 244248 12371 244260
rect 12421 244248 12467 244260
rect 12535 244248 12581 244260
rect 12631 244248 12677 244260
rect 12745 244248 12791 244260
rect 12841 244248 12887 244260
rect 12955 244248 13001 244260
rect 13051 244248 13097 244260
rect 13165 244248 13211 244260
rect 13261 244248 13307 244260
rect 13375 244248 13421 244260
rect 13471 244248 13517 244260
rect 13585 244248 13631 244260
rect 13681 244248 13727 244260
rect 13795 244248 13841 244260
rect 13891 244248 13937 244260
rect 14005 244248 14051 244260
rect 14101 244248 14147 244260
rect 14215 244248 14261 244260
rect 14311 244248 14357 244260
rect 14425 244248 14471 244260
rect 14521 244248 14567 244260
rect 14635 244248 14681 244260
rect 14731 244248 14777 244260
rect 14845 244248 14891 244260
rect 14941 244248 14987 244260
rect 15055 244248 15101 244260
rect 15151 244248 15197 244260
rect 15265 244248 15311 244260
rect 15361 244248 15407 244260
rect 15475 244248 15521 244260
rect 15571 244248 15617 244260
rect 15685 244248 15731 244260
rect 15781 244248 15827 244260
rect 15895 244248 15941 244260
rect 15991 244248 16037 244260
rect 16105 244248 16151 244260
rect 16201 244248 16247 244260
rect 16315 244248 16361 244260
rect 16411 244248 16457 244260
rect 16525 244248 16571 244260
rect 16621 244248 16667 244260
rect 16735 244248 16781 244260
rect 16831 244248 16877 244260
rect 16945 244248 16991 244260
rect 17041 244248 17087 244260
rect 17155 244248 17201 244260
rect 17251 244248 17297 244260
rect 17365 244248 17411 244260
rect 17461 244248 17507 244260
rect 17575 244248 17621 244260
rect 17671 244248 17717 244260
rect 17785 244248 17831 244260
rect 17881 244248 17927 244260
rect 17995 244248 18041 244260
rect 18091 244248 18137 244260
rect 18205 244248 18251 244260
rect 18301 244248 18347 244260
rect 18415 244248 18461 244260
rect 18511 244248 18557 244260
rect 18625 244248 18671 244260
rect 18721 244248 18767 244260
rect 18835 244248 18881 244260
rect 18931 244248 18977 244260
rect 19045 244248 19091 244260
rect 19141 244248 19187 244260
rect 19255 244248 19301 244260
rect 19351 244248 19397 244260
rect 19465 244248 19511 244260
rect 19561 244248 19607 244260
rect 19675 244248 19721 244260
rect 19771 244248 19817 244260
rect 19885 244248 19931 244260
rect 19981 244248 20027 244260
rect 20095 244248 20141 244260
rect 20191 244248 20237 244260
rect 20305 244248 20351 244260
rect 20401 244248 20447 244260
rect 20515 244248 20561 244260
rect 20611 244248 20657 244260
rect 20725 244248 20771 244260
rect 20821 244248 20867 244260
rect 20935 244248 20981 244260
rect 21031 244248 21077 244260
rect 21145 244248 21191 244260
rect 21241 244248 21287 244260
rect 21355 244248 21401 244260
rect 21451 244248 21497 244260
rect 21565 244248 21611 244260
rect 21661 244248 21707 244260
rect 21775 244248 21821 244260
rect 21871 244248 21917 244260
rect 21985 244248 22031 244260
rect 22081 244248 22127 244260
rect 22195 244248 22241 244260
rect 22291 244248 22337 244260
rect 22405 244248 22451 244260
rect 22501 244248 22547 244260
rect 22615 244248 22661 244260
rect 22711 244248 22757 244260
rect 22825 244248 22871 244260
rect 22921 244248 22967 244260
rect 23035 244248 23081 244260
rect 23131 244248 23177 244260
rect 23245 244248 23291 244260
rect 23341 244248 23387 244260
rect 23455 244248 23501 244260
rect 23551 244248 23597 244260
rect 23665 244248 23711 244260
rect 23761 244248 23807 244260
rect 23875 244248 23921 244260
rect 23971 244248 24017 244260
rect 24085 244248 24131 244260
rect 24181 244248 24227 244260
rect 24295 244248 24341 244260
rect 24391 244248 24437 244260
rect 24505 244248 24551 244260
rect 24601 244248 24647 244260
rect 24715 244248 24761 244260
rect 24811 244248 24857 244260
rect 24925 244248 24971 244260
rect 25021 244248 25067 244260
rect 25135 244248 25181 244260
rect 25231 244248 25277 244260
rect 25345 244248 25391 244260
rect 25441 244248 25487 244260
rect 25555 244248 25601 244260
rect 25651 244248 25697 244260
rect 25765 244248 25811 244260
rect 25861 244248 25907 244260
rect 25975 244248 26021 244260
rect 26071 244248 26117 244260
rect 26185 244248 26231 244260
rect 26281 244248 26327 244260
rect 26395 244248 26441 244260
rect 26491 244248 26537 244260
rect 26605 244248 26651 244260
rect 26701 244248 26747 244260
rect 26815 244248 26861 244260
rect 26911 244248 26957 244260
rect 27025 244248 27071 244260
rect 27121 244248 27167 244260
rect 27235 244248 27281 244260
rect 27331 244248 27566 244260
rect -5008 244201 27406 244207
rect -5008 244167 -3791 244201
rect -3695 244167 -3371 244201
rect -3275 244167 -2951 244201
rect -2855 244167 -2531 244201
rect -2435 244167 -2111 244201
rect -2015 244167 -1691 244201
rect -1595 244167 -1271 244201
rect -1175 244167 -851 244201
rect -755 244167 -431 244201
rect -335 244167 -11 244201
rect 85 244167 409 244201
rect 505 244167 829 244201
rect 925 244167 1249 244201
rect 1345 244167 1669 244201
rect 1765 244167 2089 244201
rect 2185 244167 2509 244201
rect 2605 244167 2929 244201
rect 3025 244167 3349 244201
rect 3445 244167 3769 244201
rect 3865 244167 4189 244201
rect 4285 244167 4609 244201
rect 4705 244167 5029 244201
rect 5125 244167 5449 244201
rect 5545 244167 5869 244201
rect 5965 244167 6289 244201
rect 6385 244167 6709 244201
rect 6805 244167 7129 244201
rect 7225 244167 7549 244201
rect 7645 244167 7969 244201
rect 8065 244167 8389 244201
rect 8485 244167 8809 244201
rect 8905 244167 9229 244201
rect 9325 244167 9649 244201
rect 9745 244167 10069 244201
rect 10165 244167 10489 244201
rect 10585 244167 10909 244201
rect 11005 244167 11329 244201
rect 11425 244167 11749 244201
rect 11845 244167 12169 244201
rect 12265 244167 12589 244201
rect 12685 244167 13009 244201
rect 13105 244167 13429 244201
rect 13525 244167 13849 244201
rect 13945 244167 14269 244201
rect 14365 244167 14689 244201
rect 14785 244167 15109 244201
rect 15205 244167 15529 244201
rect 15625 244167 15949 244201
rect 16045 244167 16369 244201
rect 16465 244167 16789 244201
rect 16885 244167 17209 244201
rect 17305 244167 17629 244201
rect 17725 244167 18049 244201
rect 18145 244167 18469 244201
rect 18565 244167 18889 244201
rect 18985 244167 19309 244201
rect 19405 244167 19729 244201
rect 19825 244167 20149 244201
rect 20245 244167 20569 244201
rect 20665 244167 20989 244201
rect 21085 244167 21409 244201
rect 21505 244167 21829 244201
rect 21925 244167 22249 244201
rect 22345 244167 22669 244201
rect 22765 244167 23089 244201
rect 23185 244167 23509 244201
rect 23605 244167 23929 244201
rect 24025 244167 24349 244201
rect 24445 244167 24769 244201
rect 24865 244167 25189 244201
rect 25285 244167 25609 244201
rect 25705 244167 26029 244201
rect 26125 244167 26449 244201
rect 26545 244167 26869 244201
rect 26965 244167 27289 244201
rect 27385 244167 27406 244201
rect -5008 244161 27406 244167
rect 27467 244071 27566 244248
rect -4175 244065 27566 244071
rect -4175 243960 -4163 244065
rect 27485 244041 27566 244065
rect -4175 243954 27414 243960
rect 27404 243841 27414 243954
rect 27614 243841 27624 244041
<< via1 >>
rect 27310 264317 27510 264430
rect -4163 264212 27486 264317
rect 27486 264230 27510 264317
rect -4070 263250 -4049 264026
rect -4049 263250 -4015 264026
rect -3953 263250 -3919 264026
rect -3919 263250 -3839 264026
rect -3839 263250 -3805 264026
rect -3743 263250 -3709 264026
rect -3709 263250 -3629 264026
rect -3629 263250 -3595 264026
rect -3533 263250 -3499 264026
rect -3499 263250 -3419 264026
rect -3419 263250 -3385 264026
rect -3323 263250 -3289 264026
rect -3289 263250 -3209 264026
rect -3209 263250 -3175 264026
rect -3113 263250 -3079 264026
rect -3079 263250 -2999 264026
rect -2999 263250 -2965 264026
rect -2903 263250 -2869 264026
rect -2869 263250 -2789 264026
rect -2789 263250 -2755 264026
rect -2693 263250 -2659 264026
rect -2659 263250 -2579 264026
rect -2579 263250 -2545 264026
rect -2483 263250 -2449 264026
rect -2449 263250 -2369 264026
rect -2369 263250 -2335 264026
rect -2273 263250 -2239 264026
rect -2239 263250 -2159 264026
rect -2159 263250 -2125 264026
rect -2063 263250 -2029 264026
rect -2029 263250 -1949 264026
rect -1949 263250 -1915 264026
rect -1853 263250 -1819 264026
rect -1819 263250 -1739 264026
rect -1739 263250 -1705 264026
rect -1643 263250 -1609 264026
rect -1609 263250 -1529 264026
rect -1529 263250 -1495 264026
rect -1433 263250 -1399 264026
rect -1399 263250 -1319 264026
rect -1319 263250 -1285 264026
rect -1223 263250 -1189 264026
rect -1189 263250 -1109 264026
rect -1109 263250 -1075 264026
rect -1013 263250 -979 264026
rect -979 263250 -899 264026
rect -899 263250 -865 264026
rect -803 263250 -769 264026
rect -769 263250 -689 264026
rect -689 263250 -655 264026
rect -593 263250 -559 264026
rect -559 263250 -479 264026
rect -479 263250 -445 264026
rect -383 263250 -349 264026
rect -349 263250 -269 264026
rect -269 263250 -235 264026
rect -173 263250 -139 264026
rect -139 263250 -59 264026
rect -59 263250 -25 264026
rect 37 263250 71 264026
rect 71 263250 151 264026
rect 151 263250 185 264026
rect 247 263250 281 264026
rect 281 263250 361 264026
rect 361 263250 395 264026
rect 457 263250 491 264026
rect 491 263250 571 264026
rect 571 263250 605 264026
rect 667 263250 701 264026
rect 701 263250 781 264026
rect 781 263250 815 264026
rect 877 263250 911 264026
rect 911 263250 991 264026
rect 991 263250 1025 264026
rect 1087 263250 1121 264026
rect 1121 263250 1201 264026
rect 1201 263250 1235 264026
rect 1297 263250 1331 264026
rect 1331 263250 1411 264026
rect 1411 263250 1445 264026
rect 1507 263250 1541 264026
rect 1541 263250 1621 264026
rect 1621 263250 1655 264026
rect 1717 263250 1751 264026
rect 1751 263250 1831 264026
rect 1831 263250 1865 264026
rect 1927 263250 1961 264026
rect 1961 263250 2041 264026
rect 2041 263250 2075 264026
rect 2137 263250 2171 264026
rect 2171 263250 2251 264026
rect 2251 263250 2285 264026
rect 2347 263250 2381 264026
rect 2381 263250 2461 264026
rect 2461 263250 2495 264026
rect 2557 263250 2591 264026
rect 2591 263250 2671 264026
rect 2671 263250 2705 264026
rect 2767 263250 2801 264026
rect 2801 263250 2881 264026
rect 2881 263250 2915 264026
rect 2977 263250 3011 264026
rect 3011 263250 3091 264026
rect 3091 263250 3125 264026
rect 3187 263250 3221 264026
rect 3221 263250 3301 264026
rect 3301 263250 3335 264026
rect 3397 263250 3431 264026
rect 3431 263250 3511 264026
rect 3511 263250 3545 264026
rect 3607 263250 3641 264026
rect 3641 263250 3721 264026
rect 3721 263250 3755 264026
rect 3817 263250 3851 264026
rect 3851 263250 3931 264026
rect 3931 263250 3965 264026
rect 4027 263250 4061 264026
rect 4061 263250 4141 264026
rect 4141 263250 4175 264026
rect 4237 263250 4271 264026
rect 4271 263250 4351 264026
rect 4351 263250 4385 264026
rect 4447 263250 4481 264026
rect 4481 263250 4561 264026
rect 4561 263250 4595 264026
rect 4657 263250 4691 264026
rect 4691 263250 4771 264026
rect 4771 263250 4805 264026
rect 4867 263250 4901 264026
rect 4901 263250 4981 264026
rect 4981 263250 5015 264026
rect 5077 263250 5111 264026
rect 5111 263250 5191 264026
rect 5191 263250 5225 264026
rect 5287 263250 5321 264026
rect 5321 263250 5401 264026
rect 5401 263250 5435 264026
rect 5497 263250 5531 264026
rect 5531 263250 5611 264026
rect 5611 263250 5645 264026
rect 5707 263250 5741 264026
rect 5741 263250 5821 264026
rect 5821 263250 5855 264026
rect 5917 263250 5951 264026
rect 5951 263250 6031 264026
rect 6031 263250 6065 264026
rect 6127 263250 6161 264026
rect 6161 263250 6241 264026
rect 6241 263250 6275 264026
rect 6337 263250 6371 264026
rect 6371 263250 6451 264026
rect 6451 263250 6485 264026
rect 6547 263250 6581 264026
rect 6581 263250 6661 264026
rect 6661 263250 6695 264026
rect 6757 263250 6791 264026
rect 6791 263250 6871 264026
rect 6871 263250 6905 264026
rect 6967 263250 7001 264026
rect 7001 263250 7081 264026
rect 7081 263250 7115 264026
rect 7177 263250 7211 264026
rect 7211 263250 7291 264026
rect 7291 263250 7325 264026
rect 7387 263250 7421 264026
rect 7421 263250 7501 264026
rect 7501 263250 7535 264026
rect 7597 263250 7631 264026
rect 7631 263250 7711 264026
rect 7711 263250 7745 264026
rect 7807 263250 7841 264026
rect 7841 263250 7921 264026
rect 7921 263250 7955 264026
rect 8017 263250 8051 264026
rect 8051 263250 8131 264026
rect 8131 263250 8165 264026
rect 8227 263250 8261 264026
rect 8261 263250 8341 264026
rect 8341 263250 8375 264026
rect 8437 263250 8471 264026
rect 8471 263250 8551 264026
rect 8551 263250 8585 264026
rect 8647 263250 8681 264026
rect 8681 263250 8761 264026
rect 8761 263250 8795 264026
rect 8857 263250 8891 264026
rect 8891 263250 8971 264026
rect 8971 263250 9005 264026
rect 9067 263250 9101 264026
rect 9101 263250 9181 264026
rect 9181 263250 9215 264026
rect 9277 263250 9311 264026
rect 9311 263250 9391 264026
rect 9391 263250 9425 264026
rect 9487 263250 9521 264026
rect 9521 263250 9601 264026
rect 9601 263250 9635 264026
rect 9697 263250 9731 264026
rect 9731 263250 9811 264026
rect 9811 263250 9845 264026
rect 9907 263250 9941 264026
rect 9941 263250 10021 264026
rect 10021 263250 10055 264026
rect 10117 263250 10151 264026
rect 10151 263250 10231 264026
rect 10231 263250 10265 264026
rect 10327 263250 10361 264026
rect 10361 263250 10441 264026
rect 10441 263250 10475 264026
rect 10537 263250 10571 264026
rect 10571 263250 10651 264026
rect 10651 263250 10685 264026
rect 10747 263250 10781 264026
rect 10781 263250 10861 264026
rect 10861 263250 10895 264026
rect 10957 263250 10991 264026
rect 10991 263250 11071 264026
rect 11071 263250 11105 264026
rect 11167 263250 11201 264026
rect 11201 263250 11281 264026
rect 11281 263250 11315 264026
rect 11377 263250 11411 264026
rect 11411 263250 11491 264026
rect 11491 263250 11525 264026
rect 11587 263250 11621 264026
rect 11621 263250 11701 264026
rect 11701 263250 11735 264026
rect 11797 263250 11831 264026
rect 11831 263250 11911 264026
rect 11911 263250 11945 264026
rect 12007 263250 12041 264026
rect 12041 263250 12121 264026
rect 12121 263250 12155 264026
rect 12217 263250 12251 264026
rect 12251 263250 12331 264026
rect 12331 263250 12365 264026
rect 12427 263250 12461 264026
rect 12461 263250 12541 264026
rect 12541 263250 12575 264026
rect 12637 263250 12671 264026
rect 12671 263250 12751 264026
rect 12751 263250 12785 264026
rect 12847 263250 12881 264026
rect 12881 263250 12961 264026
rect 12961 263250 12995 264026
rect 13057 263250 13091 264026
rect 13091 263250 13171 264026
rect 13171 263250 13205 264026
rect 13267 263250 13301 264026
rect 13301 263250 13381 264026
rect 13381 263250 13415 264026
rect 13477 263250 13511 264026
rect 13511 263250 13591 264026
rect 13591 263250 13625 264026
rect 13687 263250 13721 264026
rect 13721 263250 13801 264026
rect 13801 263250 13835 264026
rect 13897 263250 13931 264026
rect 13931 263250 14011 264026
rect 14011 263250 14045 264026
rect 14107 263250 14141 264026
rect 14141 263250 14221 264026
rect 14221 263250 14255 264026
rect 14317 263250 14351 264026
rect 14351 263250 14431 264026
rect 14431 263250 14465 264026
rect 14527 263250 14561 264026
rect 14561 263250 14641 264026
rect 14641 263250 14675 264026
rect 14737 263250 14771 264026
rect 14771 263250 14851 264026
rect 14851 263250 14885 264026
rect 14947 263250 14981 264026
rect 14981 263250 15061 264026
rect 15061 263250 15095 264026
rect 15157 263250 15191 264026
rect 15191 263250 15271 264026
rect 15271 263250 15305 264026
rect 15367 263250 15401 264026
rect 15401 263250 15481 264026
rect 15481 263250 15515 264026
rect 15577 263250 15611 264026
rect 15611 263250 15691 264026
rect 15691 263250 15725 264026
rect 15787 263250 15821 264026
rect 15821 263250 15901 264026
rect 15901 263250 15935 264026
rect 15997 263250 16031 264026
rect 16031 263250 16111 264026
rect 16111 263250 16145 264026
rect 16207 263250 16241 264026
rect 16241 263250 16321 264026
rect 16321 263250 16355 264026
rect 16417 263250 16451 264026
rect 16451 263250 16531 264026
rect 16531 263250 16565 264026
rect 16627 263250 16661 264026
rect 16661 263250 16741 264026
rect 16741 263250 16775 264026
rect 16837 263250 16871 264026
rect 16871 263250 16951 264026
rect 16951 263250 16985 264026
rect 17047 263250 17081 264026
rect 17081 263250 17161 264026
rect 17161 263250 17195 264026
rect 17257 263250 17291 264026
rect 17291 263250 17371 264026
rect 17371 263250 17405 264026
rect 17467 263250 17501 264026
rect 17501 263250 17581 264026
rect 17581 263250 17615 264026
rect 17677 263250 17711 264026
rect 17711 263250 17791 264026
rect 17791 263250 17825 264026
rect 17887 263250 17921 264026
rect 17921 263250 18001 264026
rect 18001 263250 18035 264026
rect 18097 263250 18131 264026
rect 18131 263250 18211 264026
rect 18211 263250 18245 264026
rect 18307 263250 18341 264026
rect 18341 263250 18421 264026
rect 18421 263250 18455 264026
rect 18517 263250 18551 264026
rect 18551 263250 18631 264026
rect 18631 263250 18665 264026
rect 18727 263250 18761 264026
rect 18761 263250 18841 264026
rect 18841 263250 18875 264026
rect 18937 263250 18971 264026
rect 18971 263250 19051 264026
rect 19051 263250 19085 264026
rect 19147 263250 19181 264026
rect 19181 263250 19261 264026
rect 19261 263250 19295 264026
rect 19357 263250 19391 264026
rect 19391 263250 19471 264026
rect 19471 263250 19505 264026
rect 19567 263250 19601 264026
rect 19601 263250 19681 264026
rect 19681 263250 19715 264026
rect 19777 263250 19811 264026
rect 19811 263250 19891 264026
rect 19891 263250 19925 264026
rect 19987 263250 20021 264026
rect 20021 263250 20101 264026
rect 20101 263250 20135 264026
rect 20197 263250 20231 264026
rect 20231 263250 20311 264026
rect 20311 263250 20345 264026
rect 20407 263250 20441 264026
rect 20441 263250 20521 264026
rect 20521 263250 20555 264026
rect 20617 263250 20651 264026
rect 20651 263250 20731 264026
rect 20731 263250 20765 264026
rect 20827 263250 20861 264026
rect 20861 263250 20941 264026
rect 20941 263250 20975 264026
rect 21037 263250 21071 264026
rect 21071 263250 21151 264026
rect 21151 263250 21185 264026
rect 21247 263250 21281 264026
rect 21281 263250 21361 264026
rect 21361 263250 21395 264026
rect 21457 263250 21491 264026
rect 21491 263250 21571 264026
rect 21571 263250 21605 264026
rect 21667 263250 21701 264026
rect 21701 263250 21781 264026
rect 21781 263250 21815 264026
rect 21877 263250 21911 264026
rect 21911 263250 21991 264026
rect 21991 263250 22025 264026
rect 22087 263250 22121 264026
rect 22121 263250 22201 264026
rect 22201 263250 22235 264026
rect 22297 263250 22331 264026
rect 22331 263250 22411 264026
rect 22411 263250 22445 264026
rect 22507 263250 22541 264026
rect 22541 263250 22621 264026
rect 22621 263250 22655 264026
rect 22717 263250 22751 264026
rect 22751 263250 22831 264026
rect 22831 263250 22865 264026
rect 22927 263250 22961 264026
rect 22961 263250 23041 264026
rect 23041 263250 23075 264026
rect 23137 263250 23171 264026
rect 23171 263250 23251 264026
rect 23251 263250 23285 264026
rect 23347 263250 23381 264026
rect 23381 263250 23461 264026
rect 23461 263250 23495 264026
rect 23557 263250 23591 264026
rect 23591 263250 23671 264026
rect 23671 263250 23705 264026
rect 23767 263250 23801 264026
rect 23801 263250 23881 264026
rect 23881 263250 23915 264026
rect 23977 263250 24011 264026
rect 24011 263250 24091 264026
rect 24091 263250 24125 264026
rect 24187 263250 24221 264026
rect 24221 263250 24301 264026
rect 24301 263250 24335 264026
rect 24397 263250 24431 264026
rect 24431 263250 24511 264026
rect 24511 263250 24545 264026
rect 24607 263250 24641 264026
rect 24641 263250 24721 264026
rect 24721 263250 24755 264026
rect 24817 263250 24851 264026
rect 24851 263250 24931 264026
rect 24931 263250 24965 264026
rect 25027 263250 25061 264026
rect 25061 263250 25141 264026
rect 25141 263250 25175 264026
rect 25237 263250 25271 264026
rect 25271 263250 25351 264026
rect 25351 263250 25385 264026
rect 25447 263250 25481 264026
rect 25481 263250 25561 264026
rect 25561 263250 25595 264026
rect 25657 263250 25691 264026
rect 25691 263250 25771 264026
rect 25771 263250 25805 264026
rect 25867 263250 25901 264026
rect 25901 263250 25981 264026
rect 25981 263250 26015 264026
rect 26077 263250 26111 264026
rect 26111 263250 26191 264026
rect 26191 263250 26225 264026
rect 26287 263250 26321 264026
rect 26321 263250 26401 264026
rect 26401 263250 26435 264026
rect 26497 263250 26531 264026
rect 26531 263250 26611 264026
rect 26611 263250 26645 264026
rect 26707 263250 26741 264026
rect 26741 263250 26821 264026
rect 26821 263250 26855 264026
rect 26917 263250 26951 264026
rect 26951 263250 27031 264026
rect 27031 263250 27065 264026
rect 27127 263250 27161 264026
rect 27161 263250 27241 264026
rect 27241 263250 27275 264026
rect -4070 262228 -4049 263004
rect -4049 262228 -4015 263004
rect -3953 262228 -3919 263004
rect -3919 262228 -3839 263004
rect -3839 262228 -3805 263004
rect -3743 262228 -3709 263004
rect -3709 262228 -3629 263004
rect -3629 262228 -3595 263004
rect -3533 262228 -3499 263004
rect -3499 262228 -3419 263004
rect -3419 262228 -3385 263004
rect -3323 262228 -3289 263004
rect -3289 262228 -3209 263004
rect -3209 262228 -3175 263004
rect -3113 262228 -3079 263004
rect -3079 262228 -2999 263004
rect -2999 262228 -2965 263004
rect -2903 262228 -2869 263004
rect -2869 262228 -2789 263004
rect -2789 262228 -2755 263004
rect -2693 262228 -2659 263004
rect -2659 262228 -2579 263004
rect -2579 262228 -2545 263004
rect -2483 262228 -2449 263004
rect -2449 262228 -2369 263004
rect -2369 262228 -2335 263004
rect -2273 262228 -2239 263004
rect -2239 262228 -2159 263004
rect -2159 262228 -2125 263004
rect -2063 262228 -2029 263004
rect -2029 262228 -1949 263004
rect -1949 262228 -1915 263004
rect -1853 262228 -1819 263004
rect -1819 262228 -1739 263004
rect -1739 262228 -1705 263004
rect -1643 262228 -1609 263004
rect -1609 262228 -1529 263004
rect -1529 262228 -1495 263004
rect -1433 262228 -1399 263004
rect -1399 262228 -1319 263004
rect -1319 262228 -1285 263004
rect -1223 262228 -1189 263004
rect -1189 262228 -1109 263004
rect -1109 262228 -1075 263004
rect -1013 262228 -979 263004
rect -979 262228 -899 263004
rect -899 262228 -865 263004
rect -803 262228 -769 263004
rect -769 262228 -689 263004
rect -689 262228 -655 263004
rect -593 262228 -559 263004
rect -559 262228 -479 263004
rect -479 262228 -445 263004
rect -383 262228 -349 263004
rect -349 262228 -269 263004
rect -269 262228 -235 263004
rect -173 262228 -139 263004
rect -139 262228 -59 263004
rect -59 262228 -25 263004
rect 37 262228 71 263004
rect 71 262228 151 263004
rect 151 262228 185 263004
rect 247 262228 281 263004
rect 281 262228 361 263004
rect 361 262228 395 263004
rect 457 262228 491 263004
rect 491 262228 571 263004
rect 571 262228 605 263004
rect 667 262228 701 263004
rect 701 262228 781 263004
rect 781 262228 815 263004
rect 877 262228 911 263004
rect 911 262228 991 263004
rect 991 262228 1025 263004
rect 1087 262228 1121 263004
rect 1121 262228 1201 263004
rect 1201 262228 1235 263004
rect 1297 262228 1331 263004
rect 1331 262228 1411 263004
rect 1411 262228 1445 263004
rect 1507 262228 1541 263004
rect 1541 262228 1621 263004
rect 1621 262228 1655 263004
rect 1717 262228 1751 263004
rect 1751 262228 1831 263004
rect 1831 262228 1865 263004
rect 1927 262228 1961 263004
rect 1961 262228 2041 263004
rect 2041 262228 2075 263004
rect 2137 262228 2171 263004
rect 2171 262228 2251 263004
rect 2251 262228 2285 263004
rect 2347 262228 2381 263004
rect 2381 262228 2461 263004
rect 2461 262228 2495 263004
rect 2557 262228 2591 263004
rect 2591 262228 2671 263004
rect 2671 262228 2705 263004
rect 2767 262228 2801 263004
rect 2801 262228 2881 263004
rect 2881 262228 2915 263004
rect 2977 262228 3011 263004
rect 3011 262228 3091 263004
rect 3091 262228 3125 263004
rect 3187 262228 3221 263004
rect 3221 262228 3301 263004
rect 3301 262228 3335 263004
rect 3397 262228 3431 263004
rect 3431 262228 3511 263004
rect 3511 262228 3545 263004
rect 3607 262228 3641 263004
rect 3641 262228 3721 263004
rect 3721 262228 3755 263004
rect 3817 262228 3851 263004
rect 3851 262228 3931 263004
rect 3931 262228 3965 263004
rect 4027 262228 4061 263004
rect 4061 262228 4141 263004
rect 4141 262228 4175 263004
rect 4237 262228 4271 263004
rect 4271 262228 4351 263004
rect 4351 262228 4385 263004
rect 4447 262228 4481 263004
rect 4481 262228 4561 263004
rect 4561 262228 4595 263004
rect 4657 262228 4691 263004
rect 4691 262228 4771 263004
rect 4771 262228 4805 263004
rect 4867 262228 4901 263004
rect 4901 262228 4981 263004
rect 4981 262228 5015 263004
rect 5077 262228 5111 263004
rect 5111 262228 5191 263004
rect 5191 262228 5225 263004
rect 5287 262228 5321 263004
rect 5321 262228 5401 263004
rect 5401 262228 5435 263004
rect 5497 262228 5531 263004
rect 5531 262228 5611 263004
rect 5611 262228 5645 263004
rect 5707 262228 5741 263004
rect 5741 262228 5821 263004
rect 5821 262228 5855 263004
rect 5917 262228 5951 263004
rect 5951 262228 6031 263004
rect 6031 262228 6065 263004
rect 6127 262228 6161 263004
rect 6161 262228 6241 263004
rect 6241 262228 6275 263004
rect 6337 262228 6371 263004
rect 6371 262228 6451 263004
rect 6451 262228 6485 263004
rect 6547 262228 6581 263004
rect 6581 262228 6661 263004
rect 6661 262228 6695 263004
rect 6757 262228 6791 263004
rect 6791 262228 6871 263004
rect 6871 262228 6905 263004
rect 6967 262228 7001 263004
rect 7001 262228 7081 263004
rect 7081 262228 7115 263004
rect 7177 262228 7211 263004
rect 7211 262228 7291 263004
rect 7291 262228 7325 263004
rect 7387 262228 7421 263004
rect 7421 262228 7501 263004
rect 7501 262228 7535 263004
rect 7597 262228 7631 263004
rect 7631 262228 7711 263004
rect 7711 262228 7745 263004
rect 7807 262228 7841 263004
rect 7841 262228 7921 263004
rect 7921 262228 7955 263004
rect 8017 262228 8051 263004
rect 8051 262228 8131 263004
rect 8131 262228 8165 263004
rect 8227 262228 8261 263004
rect 8261 262228 8341 263004
rect 8341 262228 8375 263004
rect 8437 262228 8471 263004
rect 8471 262228 8551 263004
rect 8551 262228 8585 263004
rect 8647 262228 8681 263004
rect 8681 262228 8761 263004
rect 8761 262228 8795 263004
rect 8857 262228 8891 263004
rect 8891 262228 8971 263004
rect 8971 262228 9005 263004
rect 9067 262228 9101 263004
rect 9101 262228 9181 263004
rect 9181 262228 9215 263004
rect 9277 262228 9311 263004
rect 9311 262228 9391 263004
rect 9391 262228 9425 263004
rect 9487 262228 9521 263004
rect 9521 262228 9601 263004
rect 9601 262228 9635 263004
rect 9697 262228 9731 263004
rect 9731 262228 9811 263004
rect 9811 262228 9845 263004
rect 9907 262228 9941 263004
rect 9941 262228 10021 263004
rect 10021 262228 10055 263004
rect 10117 262228 10151 263004
rect 10151 262228 10231 263004
rect 10231 262228 10265 263004
rect 10327 262228 10361 263004
rect 10361 262228 10441 263004
rect 10441 262228 10475 263004
rect 10537 262228 10571 263004
rect 10571 262228 10651 263004
rect 10651 262228 10685 263004
rect 10747 262228 10781 263004
rect 10781 262228 10861 263004
rect 10861 262228 10895 263004
rect 10957 262228 10991 263004
rect 10991 262228 11071 263004
rect 11071 262228 11105 263004
rect 11167 262228 11201 263004
rect 11201 262228 11281 263004
rect 11281 262228 11315 263004
rect 11377 262228 11411 263004
rect 11411 262228 11491 263004
rect 11491 262228 11525 263004
rect 11587 262228 11621 263004
rect 11621 262228 11701 263004
rect 11701 262228 11735 263004
rect 11797 262228 11831 263004
rect 11831 262228 11911 263004
rect 11911 262228 11945 263004
rect 12007 262228 12041 263004
rect 12041 262228 12121 263004
rect 12121 262228 12155 263004
rect 12217 262228 12251 263004
rect 12251 262228 12331 263004
rect 12331 262228 12365 263004
rect 12427 262228 12461 263004
rect 12461 262228 12541 263004
rect 12541 262228 12575 263004
rect 12637 262228 12671 263004
rect 12671 262228 12751 263004
rect 12751 262228 12785 263004
rect 12847 262228 12881 263004
rect 12881 262228 12961 263004
rect 12961 262228 12995 263004
rect 13057 262228 13091 263004
rect 13091 262228 13171 263004
rect 13171 262228 13205 263004
rect 13267 262228 13301 263004
rect 13301 262228 13381 263004
rect 13381 262228 13415 263004
rect 13477 262228 13511 263004
rect 13511 262228 13591 263004
rect 13591 262228 13625 263004
rect 13687 262228 13721 263004
rect 13721 262228 13801 263004
rect 13801 262228 13835 263004
rect 13897 262228 13931 263004
rect 13931 262228 14011 263004
rect 14011 262228 14045 263004
rect 14107 262228 14141 263004
rect 14141 262228 14221 263004
rect 14221 262228 14255 263004
rect 14317 262228 14351 263004
rect 14351 262228 14431 263004
rect 14431 262228 14465 263004
rect 14527 262228 14561 263004
rect 14561 262228 14641 263004
rect 14641 262228 14675 263004
rect 14737 262228 14771 263004
rect 14771 262228 14851 263004
rect 14851 262228 14885 263004
rect 14947 262228 14981 263004
rect 14981 262228 15061 263004
rect 15061 262228 15095 263004
rect 15157 262228 15191 263004
rect 15191 262228 15271 263004
rect 15271 262228 15305 263004
rect 15367 262228 15401 263004
rect 15401 262228 15481 263004
rect 15481 262228 15515 263004
rect 15577 262228 15611 263004
rect 15611 262228 15691 263004
rect 15691 262228 15725 263004
rect 15787 262228 15821 263004
rect 15821 262228 15901 263004
rect 15901 262228 15935 263004
rect 15997 262228 16031 263004
rect 16031 262228 16111 263004
rect 16111 262228 16145 263004
rect 16207 262228 16241 263004
rect 16241 262228 16321 263004
rect 16321 262228 16355 263004
rect 16417 262228 16451 263004
rect 16451 262228 16531 263004
rect 16531 262228 16565 263004
rect 16627 262228 16661 263004
rect 16661 262228 16741 263004
rect 16741 262228 16775 263004
rect 16837 262228 16871 263004
rect 16871 262228 16951 263004
rect 16951 262228 16985 263004
rect 17047 262228 17081 263004
rect 17081 262228 17161 263004
rect 17161 262228 17195 263004
rect 17257 262228 17291 263004
rect 17291 262228 17371 263004
rect 17371 262228 17405 263004
rect 17467 262228 17501 263004
rect 17501 262228 17581 263004
rect 17581 262228 17615 263004
rect 17677 262228 17711 263004
rect 17711 262228 17791 263004
rect 17791 262228 17825 263004
rect 17887 262228 17921 263004
rect 17921 262228 18001 263004
rect 18001 262228 18035 263004
rect 18097 262228 18131 263004
rect 18131 262228 18211 263004
rect 18211 262228 18245 263004
rect 18307 262228 18341 263004
rect 18341 262228 18421 263004
rect 18421 262228 18455 263004
rect 18517 262228 18551 263004
rect 18551 262228 18631 263004
rect 18631 262228 18665 263004
rect 18727 262228 18761 263004
rect 18761 262228 18841 263004
rect 18841 262228 18875 263004
rect 18937 262228 18971 263004
rect 18971 262228 19051 263004
rect 19051 262228 19085 263004
rect 19147 262228 19181 263004
rect 19181 262228 19261 263004
rect 19261 262228 19295 263004
rect 19357 262228 19391 263004
rect 19391 262228 19471 263004
rect 19471 262228 19505 263004
rect 19567 262228 19601 263004
rect 19601 262228 19681 263004
rect 19681 262228 19715 263004
rect 19777 262228 19811 263004
rect 19811 262228 19891 263004
rect 19891 262228 19925 263004
rect 19987 262228 20021 263004
rect 20021 262228 20101 263004
rect 20101 262228 20135 263004
rect 20197 262228 20231 263004
rect 20231 262228 20311 263004
rect 20311 262228 20345 263004
rect 20407 262228 20441 263004
rect 20441 262228 20521 263004
rect 20521 262228 20555 263004
rect 20617 262228 20651 263004
rect 20651 262228 20731 263004
rect 20731 262228 20765 263004
rect 20827 262228 20861 263004
rect 20861 262228 20941 263004
rect 20941 262228 20975 263004
rect 21037 262228 21071 263004
rect 21071 262228 21151 263004
rect 21151 262228 21185 263004
rect 21247 262228 21281 263004
rect 21281 262228 21361 263004
rect 21361 262228 21395 263004
rect 21457 262228 21491 263004
rect 21491 262228 21571 263004
rect 21571 262228 21605 263004
rect 21667 262228 21701 263004
rect 21701 262228 21781 263004
rect 21781 262228 21815 263004
rect 21877 262228 21911 263004
rect 21911 262228 21991 263004
rect 21991 262228 22025 263004
rect 22087 262228 22121 263004
rect 22121 262228 22201 263004
rect 22201 262228 22235 263004
rect 22297 262228 22331 263004
rect 22331 262228 22411 263004
rect 22411 262228 22445 263004
rect 22507 262228 22541 263004
rect 22541 262228 22621 263004
rect 22621 262228 22655 263004
rect 22717 262228 22751 263004
rect 22751 262228 22831 263004
rect 22831 262228 22865 263004
rect 22927 262228 22961 263004
rect 22961 262228 23041 263004
rect 23041 262228 23075 263004
rect 23137 262228 23171 263004
rect 23171 262228 23251 263004
rect 23251 262228 23285 263004
rect 23347 262228 23381 263004
rect 23381 262228 23461 263004
rect 23461 262228 23495 263004
rect 23557 262228 23591 263004
rect 23591 262228 23671 263004
rect 23671 262228 23705 263004
rect 23767 262228 23801 263004
rect 23801 262228 23881 263004
rect 23881 262228 23915 263004
rect 23977 262228 24011 263004
rect 24011 262228 24091 263004
rect 24091 262228 24125 263004
rect 24187 262228 24221 263004
rect 24221 262228 24301 263004
rect 24301 262228 24335 263004
rect 24397 262228 24431 263004
rect 24431 262228 24511 263004
rect 24511 262228 24545 263004
rect 24607 262228 24641 263004
rect 24641 262228 24721 263004
rect 24721 262228 24755 263004
rect 24817 262228 24851 263004
rect 24851 262228 24931 263004
rect 24931 262228 24965 263004
rect 25027 262228 25061 263004
rect 25061 262228 25141 263004
rect 25141 262228 25175 263004
rect 25237 262228 25271 263004
rect 25271 262228 25351 263004
rect 25351 262228 25385 263004
rect 25447 262228 25481 263004
rect 25481 262228 25561 263004
rect 25561 262228 25595 263004
rect 25657 262228 25691 263004
rect 25691 262228 25771 263004
rect 25771 262228 25805 263004
rect 25867 262228 25901 263004
rect 25901 262228 25981 263004
rect 25981 262228 26015 263004
rect 26077 262228 26111 263004
rect 26111 262228 26191 263004
rect 26191 262228 26225 263004
rect 26287 262228 26321 263004
rect 26321 262228 26401 263004
rect 26401 262228 26435 263004
rect 26497 262228 26531 263004
rect 26531 262228 26611 263004
rect 26611 262228 26645 263004
rect 26707 262228 26741 263004
rect 26741 262228 26821 263004
rect 26821 262228 26855 263004
rect 26917 262228 26951 263004
rect 26951 262228 27031 263004
rect 27031 262228 27065 263004
rect 27127 262228 27161 263004
rect 27161 262228 27241 263004
rect 27241 262228 27275 263004
rect -4069 253713 -4049 254489
rect -4049 253713 -4015 254489
rect -3953 253713 -3919 254489
rect -3919 253713 -3839 254489
rect -3839 253713 -3805 254489
rect -3743 253713 -3709 254489
rect -3709 253713 -3629 254489
rect -3629 253713 -3595 254489
rect -3533 254489 -3385 254490
rect -3533 253713 -3499 254489
rect -3499 253713 -3419 254489
rect -3419 253713 -3385 254489
rect -3323 254489 -3175 254490
rect -3323 253713 -3289 254489
rect -3289 253713 -3209 254489
rect -3209 253713 -3175 254489
rect -3113 254489 -2965 254490
rect -3113 253713 -3079 254489
rect -3079 253713 -2999 254489
rect -2999 253713 -2965 254489
rect -2903 254489 -2755 254490
rect -2903 253713 -2869 254489
rect -2869 253713 -2789 254489
rect -2789 253713 -2755 254489
rect -2693 254489 -2545 254490
rect -2693 253713 -2659 254489
rect -2659 253713 -2579 254489
rect -2579 253713 -2545 254489
rect -2483 254489 -2335 254490
rect -2483 253713 -2449 254489
rect -2449 253713 -2369 254489
rect -2369 253713 -2335 254489
rect -2273 254489 -2125 254490
rect -2273 253713 -2239 254489
rect -2239 253713 -2159 254489
rect -2159 253713 -2125 254489
rect -2063 254489 -1915 254490
rect -2063 253713 -2029 254489
rect -2029 253713 -1949 254489
rect -1949 253713 -1915 254489
rect -1853 254489 -1705 254490
rect -1853 253713 -1819 254489
rect -1819 253713 -1739 254489
rect -1739 253713 -1705 254489
rect -1643 254489 -1495 254490
rect -1643 253713 -1609 254489
rect -1609 253713 -1529 254489
rect -1529 253713 -1495 254489
rect -1433 254489 -1285 254490
rect -1433 253713 -1399 254489
rect -1399 253713 -1319 254489
rect -1319 253713 -1285 254489
rect -1223 254489 -1075 254490
rect -1223 253713 -1189 254489
rect -1189 253713 -1109 254489
rect -1109 253713 -1075 254489
rect -1013 254489 -865 254490
rect -1013 253713 -979 254489
rect -979 253713 -899 254489
rect -899 253713 -865 254489
rect -803 254489 -655 254490
rect -803 253713 -769 254489
rect -769 253713 -689 254489
rect -689 253713 -655 254489
rect -593 254489 -445 254490
rect -593 253713 -559 254489
rect -559 253713 -479 254489
rect -479 253713 -445 254489
rect -383 254489 -235 254490
rect -383 253713 -349 254489
rect -349 253713 -269 254489
rect -269 253713 -235 254489
rect -173 254489 -25 254490
rect -173 253713 -139 254489
rect -139 253713 -59 254489
rect -59 253713 -25 254489
rect 37 254489 185 254490
rect 37 253713 71 254489
rect 71 253713 151 254489
rect 151 253713 185 254489
rect 247 254489 395 254490
rect 247 253713 281 254489
rect 281 253713 361 254489
rect 361 253713 395 254489
rect 457 254489 605 254490
rect 457 253713 491 254489
rect 491 253713 571 254489
rect 571 253713 605 254489
rect 667 254489 815 254490
rect 667 253713 701 254489
rect 701 253713 781 254489
rect 781 253713 815 254489
rect 877 254489 1025 254490
rect 877 253713 911 254489
rect 911 253713 991 254489
rect 991 253713 1025 254489
rect 1087 254489 1235 254490
rect 1087 253713 1121 254489
rect 1121 253713 1201 254489
rect 1201 253713 1235 254489
rect 1297 254489 1445 254490
rect 1297 253713 1331 254489
rect 1331 253713 1411 254489
rect 1411 253713 1445 254489
rect 1507 254489 1655 254490
rect 1507 253713 1541 254489
rect 1541 253713 1621 254489
rect 1621 253713 1655 254489
rect 1717 254489 1865 254490
rect 1717 253713 1751 254489
rect 1751 253713 1831 254489
rect 1831 253713 1865 254489
rect 1927 254489 2075 254490
rect 1927 253713 1961 254489
rect 1961 253713 2041 254489
rect 2041 253713 2075 254489
rect 2137 254489 2285 254490
rect 2137 253713 2171 254489
rect 2171 253713 2251 254489
rect 2251 253713 2285 254489
rect 2347 254489 2495 254490
rect 2347 253713 2381 254489
rect 2381 253713 2461 254489
rect 2461 253713 2495 254489
rect 2557 254489 2705 254490
rect 2557 253713 2591 254489
rect 2591 253713 2671 254489
rect 2671 253713 2705 254489
rect 2767 254489 2915 254490
rect 2767 253713 2801 254489
rect 2801 253713 2881 254489
rect 2881 253713 2915 254489
rect 2977 254489 3125 254490
rect 2977 253713 3011 254489
rect 3011 253713 3091 254489
rect 3091 253713 3125 254489
rect 3187 254489 3335 254490
rect 3187 253713 3221 254489
rect 3221 253713 3301 254489
rect 3301 253713 3335 254489
rect 3397 254489 3545 254490
rect 3397 253713 3431 254489
rect 3431 253713 3511 254489
rect 3511 253713 3545 254489
rect 3607 254489 3755 254490
rect 3607 253713 3641 254489
rect 3641 253713 3721 254489
rect 3721 253713 3755 254489
rect 3817 254489 3965 254490
rect 3817 253713 3851 254489
rect 3851 253713 3931 254489
rect 3931 253713 3965 254489
rect 4027 254489 4175 254490
rect 4027 253713 4061 254489
rect 4061 253713 4141 254489
rect 4141 253713 4175 254489
rect 4237 254489 4385 254490
rect 4237 253713 4271 254489
rect 4271 253713 4351 254489
rect 4351 253713 4385 254489
rect 4447 254489 4595 254490
rect 4447 253713 4481 254489
rect 4481 253713 4561 254489
rect 4561 253713 4595 254489
rect 4657 254489 4805 254490
rect 4657 253713 4691 254489
rect 4691 253713 4771 254489
rect 4771 253713 4805 254489
rect 4867 254489 5015 254490
rect 4867 253713 4901 254489
rect 4901 253713 4981 254489
rect 4981 253713 5015 254489
rect 5077 254489 5225 254490
rect 5077 253713 5111 254489
rect 5111 253713 5191 254489
rect 5191 253713 5225 254489
rect 5287 254489 5435 254490
rect 5287 253713 5321 254489
rect 5321 253713 5401 254489
rect 5401 253713 5435 254489
rect 5497 254489 5645 254490
rect 5497 253713 5531 254489
rect 5531 253713 5611 254489
rect 5611 253713 5645 254489
rect 5707 254489 5855 254490
rect 5707 253713 5741 254489
rect 5741 253713 5821 254489
rect 5821 253713 5855 254489
rect 5917 254489 6065 254490
rect 5917 253713 5951 254489
rect 5951 253713 6031 254489
rect 6031 253713 6065 254489
rect 6127 254489 6275 254490
rect 6127 253713 6161 254489
rect 6161 253713 6241 254489
rect 6241 253713 6275 254489
rect 6337 254489 6485 254490
rect 6337 253713 6371 254489
rect 6371 253713 6451 254489
rect 6451 253713 6485 254489
rect 6547 254489 6695 254490
rect 6547 253713 6581 254489
rect 6581 253713 6661 254489
rect 6661 253713 6695 254489
rect 6757 254489 6905 254490
rect 6757 253713 6791 254489
rect 6791 253713 6871 254489
rect 6871 253713 6905 254489
rect 6967 254489 7115 254490
rect 6967 253713 7001 254489
rect 7001 253713 7081 254489
rect 7081 253713 7115 254489
rect 7177 254489 7325 254490
rect 7177 253713 7211 254489
rect 7211 253713 7291 254489
rect 7291 253713 7325 254489
rect 7387 254489 7535 254490
rect 7387 253713 7421 254489
rect 7421 253713 7501 254489
rect 7501 253713 7535 254489
rect 7597 254489 7745 254490
rect 7597 253713 7631 254489
rect 7631 253713 7711 254489
rect 7711 253713 7745 254489
rect 7807 254489 7955 254490
rect 7807 253713 7841 254489
rect 7841 253713 7921 254489
rect 7921 253713 7955 254489
rect 8017 254489 8165 254490
rect 8017 253713 8051 254489
rect 8051 253713 8131 254489
rect 8131 253713 8165 254489
rect 8227 254489 8375 254490
rect 8227 253713 8261 254489
rect 8261 253713 8341 254489
rect 8341 253713 8375 254489
rect 8437 254489 8585 254490
rect 8437 253713 8471 254489
rect 8471 253713 8551 254489
rect 8551 253713 8585 254489
rect 8647 254489 8795 254490
rect 8647 253713 8681 254489
rect 8681 253713 8761 254489
rect 8761 253713 8795 254489
rect 8857 254489 9005 254490
rect 8857 253713 8891 254489
rect 8891 253713 8971 254489
rect 8971 253713 9005 254489
rect 9067 254489 9215 254490
rect 9067 253713 9101 254489
rect 9101 253713 9181 254489
rect 9181 253713 9215 254489
rect 9277 254489 9425 254490
rect 9277 253713 9311 254489
rect 9311 253713 9391 254489
rect 9391 253713 9425 254489
rect 9487 254489 9635 254490
rect 9487 253713 9521 254489
rect 9521 253713 9601 254489
rect 9601 253713 9635 254489
rect 9697 254489 9845 254490
rect 9697 253713 9731 254489
rect 9731 253713 9811 254489
rect 9811 253713 9845 254489
rect 9907 254489 10055 254490
rect 9907 253713 9941 254489
rect 9941 253713 10021 254489
rect 10021 253713 10055 254489
rect 10117 254489 10265 254490
rect 10117 253713 10151 254489
rect 10151 253713 10231 254489
rect 10231 253713 10265 254489
rect 10327 254489 10475 254490
rect 10327 253713 10361 254489
rect 10361 253713 10441 254489
rect 10441 253713 10475 254489
rect 10537 254489 10685 254490
rect 10537 253713 10571 254489
rect 10571 253713 10651 254489
rect 10651 253713 10685 254489
rect 10747 254489 10895 254490
rect 10747 253713 10781 254489
rect 10781 253713 10861 254489
rect 10861 253713 10895 254489
rect 10957 254489 11105 254490
rect 10957 253713 10991 254489
rect 10991 253713 11071 254489
rect 11071 253713 11105 254489
rect 11167 254489 11315 254490
rect 11167 253713 11201 254489
rect 11201 253713 11281 254489
rect 11281 253713 11315 254489
rect 11377 254489 11525 254490
rect 11377 253713 11411 254489
rect 11411 253713 11491 254489
rect 11491 253713 11525 254489
rect 11587 254489 11735 254490
rect 11587 253713 11621 254489
rect 11621 253713 11701 254489
rect 11701 253713 11735 254489
rect 11797 254489 11945 254490
rect 11797 253713 11831 254489
rect 11831 253713 11911 254489
rect 11911 253713 11945 254489
rect 12007 254489 12155 254490
rect 12007 253713 12041 254489
rect 12041 253713 12121 254489
rect 12121 253713 12155 254489
rect 12217 254489 12365 254490
rect 12217 253713 12251 254489
rect 12251 253713 12331 254489
rect 12331 253713 12365 254489
rect 12427 254489 12575 254490
rect 12427 253713 12461 254489
rect 12461 253713 12541 254489
rect 12541 253713 12575 254489
rect 12637 254489 12785 254490
rect 12637 253713 12671 254489
rect 12671 253713 12751 254489
rect 12751 253713 12785 254489
rect 12847 254489 12995 254490
rect 12847 253713 12881 254489
rect 12881 253713 12961 254489
rect 12961 253713 12995 254489
rect 13057 254489 13205 254490
rect 13057 253713 13091 254489
rect 13091 253713 13171 254489
rect 13171 253713 13205 254489
rect 13267 254489 13415 254490
rect 13267 253713 13301 254489
rect 13301 253713 13381 254489
rect 13381 253713 13415 254489
rect 13477 254489 13625 254490
rect 13477 253713 13511 254489
rect 13511 253713 13591 254489
rect 13591 253713 13625 254489
rect 13687 254489 13835 254490
rect 13687 253713 13721 254489
rect 13721 253713 13801 254489
rect 13801 253713 13835 254489
rect 13897 254489 14045 254490
rect 13897 253713 13931 254489
rect 13931 253713 14011 254489
rect 14011 253713 14045 254489
rect 14107 254489 14255 254490
rect 14107 253713 14141 254489
rect 14141 253713 14221 254489
rect 14221 253713 14255 254489
rect 14317 254489 14465 254490
rect 14317 253713 14351 254489
rect 14351 253713 14431 254489
rect 14431 253713 14465 254489
rect 14527 254489 14675 254490
rect 14527 253713 14561 254489
rect 14561 253713 14641 254489
rect 14641 253713 14675 254489
rect 14737 254489 14885 254490
rect 14737 253713 14771 254489
rect 14771 253713 14851 254489
rect 14851 253713 14885 254489
rect 14947 254489 15095 254490
rect 14947 253713 14981 254489
rect 14981 253713 15061 254489
rect 15061 253713 15095 254489
rect 15157 254489 15305 254490
rect 15157 253713 15191 254489
rect 15191 253713 15271 254489
rect 15271 253713 15305 254489
rect 15367 254489 15515 254490
rect 15367 253713 15401 254489
rect 15401 253713 15481 254489
rect 15481 253713 15515 254489
rect 15577 254489 15725 254490
rect 15577 253713 15611 254489
rect 15611 253713 15691 254489
rect 15691 253713 15725 254489
rect 15787 254489 15935 254490
rect 15787 253713 15821 254489
rect 15821 253713 15901 254489
rect 15901 253713 15935 254489
rect 15997 254489 16145 254490
rect 15997 253713 16031 254489
rect 16031 253713 16111 254489
rect 16111 253713 16145 254489
rect 16207 254489 16355 254490
rect 16207 253713 16241 254489
rect 16241 253713 16321 254489
rect 16321 253713 16355 254489
rect 16417 254489 16565 254490
rect 16417 253713 16451 254489
rect 16451 253713 16531 254489
rect 16531 253713 16565 254489
rect 16627 254489 16775 254490
rect 16627 253713 16661 254489
rect 16661 253713 16741 254489
rect 16741 253713 16775 254489
rect 16837 254489 16985 254490
rect 16837 253713 16871 254489
rect 16871 253713 16951 254489
rect 16951 253713 16985 254489
rect 17047 254489 17195 254490
rect 17047 253713 17081 254489
rect 17081 253713 17161 254489
rect 17161 253713 17195 254489
rect 17257 254489 17405 254490
rect 17257 253713 17291 254489
rect 17291 253713 17371 254489
rect 17371 253713 17405 254489
rect 17467 254489 17615 254490
rect 17467 253713 17501 254489
rect 17501 253713 17581 254489
rect 17581 253713 17615 254489
rect 17677 254489 17825 254490
rect 17677 253713 17711 254489
rect 17711 253713 17791 254489
rect 17791 253713 17825 254489
rect 17887 254489 18035 254490
rect 17887 253713 17921 254489
rect 17921 253713 18001 254489
rect 18001 253713 18035 254489
rect 18097 254489 18245 254490
rect 18097 253713 18131 254489
rect 18131 253713 18211 254489
rect 18211 253713 18245 254489
rect 18307 254489 18455 254490
rect 18307 253713 18341 254489
rect 18341 253713 18421 254489
rect 18421 253713 18455 254489
rect 18517 254489 18665 254490
rect 18517 253713 18551 254489
rect 18551 253713 18631 254489
rect 18631 253713 18665 254489
rect 18727 254489 18875 254490
rect 18727 253713 18761 254489
rect 18761 253713 18841 254489
rect 18841 253713 18875 254489
rect 18937 254489 19085 254490
rect 18937 253713 18971 254489
rect 18971 253713 19051 254489
rect 19051 253713 19085 254489
rect 19147 254489 19295 254490
rect 19147 253713 19181 254489
rect 19181 253713 19261 254489
rect 19261 253713 19295 254489
rect 19357 254489 19505 254490
rect 19357 253713 19391 254489
rect 19391 253713 19471 254489
rect 19471 253713 19505 254489
rect 19567 254489 19715 254490
rect 19567 253713 19601 254489
rect 19601 253713 19681 254489
rect 19681 253713 19715 254489
rect 19777 254489 19925 254490
rect 19777 253713 19811 254489
rect 19811 253713 19891 254489
rect 19891 253713 19925 254489
rect 19987 254489 20135 254490
rect 19987 253713 20021 254489
rect 20021 253713 20101 254489
rect 20101 253713 20135 254489
rect 20197 254489 20345 254490
rect 20197 253713 20231 254489
rect 20231 253713 20311 254489
rect 20311 253713 20345 254489
rect 20407 254489 20555 254490
rect 20407 253713 20441 254489
rect 20441 253713 20521 254489
rect 20521 253713 20555 254489
rect 20617 254489 20765 254490
rect 20617 253713 20651 254489
rect 20651 253713 20731 254489
rect 20731 253713 20765 254489
rect 20827 254489 20975 254490
rect 20827 253713 20861 254489
rect 20861 253713 20941 254489
rect 20941 253713 20975 254489
rect 21037 254489 21185 254490
rect 21037 253713 21071 254489
rect 21071 253713 21151 254489
rect 21151 253713 21185 254489
rect 21247 254489 21395 254490
rect 21247 253713 21281 254489
rect 21281 253713 21361 254489
rect 21361 253713 21395 254489
rect 21457 254489 21605 254490
rect 21457 253713 21491 254489
rect 21491 253713 21571 254489
rect 21571 253713 21605 254489
rect 21667 254489 21815 254490
rect 21667 253713 21701 254489
rect 21701 253713 21781 254489
rect 21781 253713 21815 254489
rect 21877 254489 22025 254490
rect 21877 253713 21911 254489
rect 21911 253713 21991 254489
rect 21991 253713 22025 254489
rect 22087 254489 22235 254490
rect 22087 253713 22121 254489
rect 22121 253713 22201 254489
rect 22201 253713 22235 254489
rect 22297 254489 22445 254490
rect 22297 253713 22331 254489
rect 22331 253713 22411 254489
rect 22411 253713 22445 254489
rect 22507 254489 22655 254490
rect 22507 253713 22541 254489
rect 22541 253713 22621 254489
rect 22621 253713 22655 254489
rect 22717 254489 22865 254490
rect 22717 253713 22751 254489
rect 22751 253713 22831 254489
rect 22831 253713 22865 254489
rect 22927 254489 23075 254490
rect 22927 253713 22961 254489
rect 22961 253713 23041 254489
rect 23041 253713 23075 254489
rect 23137 254489 23285 254490
rect 23137 253713 23171 254489
rect 23171 253713 23251 254489
rect 23251 253713 23285 254489
rect 23347 254489 23495 254490
rect 23347 253713 23381 254489
rect 23381 253713 23461 254489
rect 23461 253713 23495 254489
rect 23557 254489 23705 254490
rect 23557 253713 23591 254489
rect 23591 253713 23671 254489
rect 23671 253713 23705 254489
rect 23767 254489 23915 254490
rect 23767 253713 23801 254489
rect 23801 253713 23881 254489
rect 23881 253713 23915 254489
rect 23977 254489 24125 254490
rect 23977 253713 24011 254489
rect 24011 253713 24091 254489
rect 24091 253713 24125 254489
rect 24187 254489 24335 254490
rect 24187 253713 24221 254489
rect 24221 253713 24301 254489
rect 24301 253713 24335 254489
rect 24397 254489 24545 254490
rect 24397 253713 24431 254489
rect 24431 253713 24511 254489
rect 24511 253713 24545 254489
rect 24607 254489 24755 254490
rect 24607 253713 24641 254489
rect 24641 253713 24721 254489
rect 24721 253713 24755 254489
rect 24817 254489 24965 254490
rect 24817 253713 24851 254489
rect 24851 253713 24931 254489
rect 24931 253713 24965 254489
rect 25027 254489 25175 254490
rect 25027 253713 25061 254489
rect 25061 253713 25141 254489
rect 25141 253713 25175 254489
rect 25237 254489 25385 254490
rect 25237 253713 25271 254489
rect 25271 253713 25351 254489
rect 25351 253713 25385 254489
rect 25447 254489 25595 254490
rect 25447 253713 25481 254489
rect 25481 253713 25561 254489
rect 25561 253713 25595 254489
rect 25657 254489 25805 254490
rect 25657 253713 25691 254489
rect 25691 253713 25771 254489
rect 25771 253713 25805 254489
rect 25867 254489 26015 254490
rect 25867 253713 25901 254489
rect 25901 253713 25981 254489
rect 25981 253713 26015 254489
rect 26077 254489 26225 254490
rect 26077 253713 26111 254489
rect 26111 253713 26191 254489
rect 26191 253713 26225 254489
rect 26287 254489 26435 254490
rect 26287 253713 26321 254489
rect 26321 253713 26401 254489
rect 26401 253713 26435 254489
rect 26497 254489 26645 254490
rect 26497 253713 26531 254489
rect 26531 253713 26611 254489
rect 26611 253713 26645 254489
rect 26707 254489 26855 254490
rect 26707 253713 26741 254489
rect 26741 253713 26821 254489
rect 26821 253713 26855 254489
rect 26917 254489 27065 254490
rect 26917 253713 26951 254489
rect 26951 253713 27031 254489
rect 27031 253713 27065 254489
rect 27127 254489 27275 254490
rect 27127 253713 27161 254489
rect 27161 253713 27241 254489
rect 27241 253713 27275 254489
rect -4069 252677 -4049 253453
rect -4049 252677 -4015 253453
rect -3953 252677 -3919 253453
rect -3919 252677 -3839 253453
rect -3839 252677 -3805 253453
rect -3743 252677 -3709 253453
rect -3709 252677 -3629 253453
rect -3629 252677 -3595 253453
rect -3533 253453 -3385 253454
rect -3533 252677 -3499 253453
rect -3499 252677 -3419 253453
rect -3419 252677 -3385 253453
rect -3323 253453 -3175 253454
rect -3323 252677 -3289 253453
rect -3289 252677 -3209 253453
rect -3209 252677 -3175 253453
rect -3113 253453 -2965 253454
rect -3113 252677 -3079 253453
rect -3079 252677 -2999 253453
rect -2999 252677 -2965 253453
rect -2903 253453 -2755 253454
rect -2903 252677 -2869 253453
rect -2869 252677 -2789 253453
rect -2789 252677 -2755 253453
rect -2693 253453 -2545 253454
rect -2693 252677 -2659 253453
rect -2659 252677 -2579 253453
rect -2579 252677 -2545 253453
rect -2483 253453 -2335 253454
rect -2483 252677 -2449 253453
rect -2449 252677 -2369 253453
rect -2369 252677 -2335 253453
rect -2273 253453 -2125 253454
rect -2273 252677 -2239 253453
rect -2239 252677 -2159 253453
rect -2159 252677 -2125 253453
rect -2063 253453 -1915 253454
rect -2063 252677 -2029 253453
rect -2029 252677 -1949 253453
rect -1949 252677 -1915 253453
rect -1853 253453 -1705 253454
rect -1853 252677 -1819 253453
rect -1819 252677 -1739 253453
rect -1739 252677 -1705 253453
rect -1643 253453 -1495 253454
rect -1643 252677 -1609 253453
rect -1609 252677 -1529 253453
rect -1529 252677 -1495 253453
rect -1433 253453 -1285 253454
rect -1433 252677 -1399 253453
rect -1399 252677 -1319 253453
rect -1319 252677 -1285 253453
rect -1223 253453 -1075 253454
rect -1223 252677 -1189 253453
rect -1189 252677 -1109 253453
rect -1109 252677 -1075 253453
rect -1013 253453 -865 253454
rect -1013 252677 -979 253453
rect -979 252677 -899 253453
rect -899 252677 -865 253453
rect -803 253453 -655 253454
rect -803 252677 -769 253453
rect -769 252677 -689 253453
rect -689 252677 -655 253453
rect -593 253453 -445 253454
rect -593 252677 -559 253453
rect -559 252677 -479 253453
rect -479 252677 -445 253453
rect -383 253453 -235 253454
rect -383 252677 -349 253453
rect -349 252677 -269 253453
rect -269 252677 -235 253453
rect -173 253453 -25 253454
rect -173 252677 -139 253453
rect -139 252677 -59 253453
rect -59 252677 -25 253453
rect 37 253453 185 253454
rect 37 252677 71 253453
rect 71 252677 151 253453
rect 151 252677 185 253453
rect 247 253453 395 253454
rect 247 252677 281 253453
rect 281 252677 361 253453
rect 361 252677 395 253453
rect 457 253453 605 253454
rect 457 252677 491 253453
rect 491 252677 571 253453
rect 571 252677 605 253453
rect 667 253453 815 253454
rect 667 252677 701 253453
rect 701 252677 781 253453
rect 781 252677 815 253453
rect 877 253453 1025 253454
rect 877 252677 911 253453
rect 911 252677 991 253453
rect 991 252677 1025 253453
rect 1087 253453 1235 253454
rect 1087 252677 1121 253453
rect 1121 252677 1201 253453
rect 1201 252677 1235 253453
rect 1297 253453 1445 253454
rect 1297 252677 1331 253453
rect 1331 252677 1411 253453
rect 1411 252677 1445 253453
rect 1507 253453 1655 253454
rect 1507 252677 1541 253453
rect 1541 252677 1621 253453
rect 1621 252677 1655 253453
rect 1717 253453 1865 253454
rect 1717 252677 1751 253453
rect 1751 252677 1831 253453
rect 1831 252677 1865 253453
rect 1927 253453 2075 253454
rect 1927 252677 1961 253453
rect 1961 252677 2041 253453
rect 2041 252677 2075 253453
rect 2137 253453 2285 253454
rect 2137 252677 2171 253453
rect 2171 252677 2251 253453
rect 2251 252677 2285 253453
rect 2347 253453 2495 253454
rect 2347 252677 2381 253453
rect 2381 252677 2461 253453
rect 2461 252677 2495 253453
rect 2557 253453 2705 253454
rect 2557 252677 2591 253453
rect 2591 252677 2671 253453
rect 2671 252677 2705 253453
rect 2767 253453 2915 253454
rect 2767 252677 2801 253453
rect 2801 252677 2881 253453
rect 2881 252677 2915 253453
rect 2977 253453 3125 253454
rect 2977 252677 3011 253453
rect 3011 252677 3091 253453
rect 3091 252677 3125 253453
rect 3187 253453 3335 253454
rect 3187 252677 3221 253453
rect 3221 252677 3301 253453
rect 3301 252677 3335 253453
rect 3397 253453 3545 253454
rect 3397 252677 3431 253453
rect 3431 252677 3511 253453
rect 3511 252677 3545 253453
rect 3607 253453 3755 253454
rect 3607 252677 3641 253453
rect 3641 252677 3721 253453
rect 3721 252677 3755 253453
rect 3817 253453 3965 253454
rect 3817 252677 3851 253453
rect 3851 252677 3931 253453
rect 3931 252677 3965 253453
rect 4027 253453 4175 253454
rect 4027 252677 4061 253453
rect 4061 252677 4141 253453
rect 4141 252677 4175 253453
rect 4237 253453 4385 253454
rect 4237 252677 4271 253453
rect 4271 252677 4351 253453
rect 4351 252677 4385 253453
rect 4447 253453 4595 253454
rect 4447 252677 4481 253453
rect 4481 252677 4561 253453
rect 4561 252677 4595 253453
rect 4657 253453 4805 253454
rect 4657 252677 4691 253453
rect 4691 252677 4771 253453
rect 4771 252677 4805 253453
rect 4867 253453 5015 253454
rect 4867 252677 4901 253453
rect 4901 252677 4981 253453
rect 4981 252677 5015 253453
rect 5077 253453 5225 253454
rect 5077 252677 5111 253453
rect 5111 252677 5191 253453
rect 5191 252677 5225 253453
rect 5287 253453 5435 253454
rect 5287 252677 5321 253453
rect 5321 252677 5401 253453
rect 5401 252677 5435 253453
rect 5497 253453 5645 253454
rect 5497 252677 5531 253453
rect 5531 252677 5611 253453
rect 5611 252677 5645 253453
rect 5707 253453 5855 253454
rect 5707 252677 5741 253453
rect 5741 252677 5821 253453
rect 5821 252677 5855 253453
rect 5917 253453 6065 253454
rect 5917 252677 5951 253453
rect 5951 252677 6031 253453
rect 6031 252677 6065 253453
rect 6127 253453 6275 253454
rect 6127 252677 6161 253453
rect 6161 252677 6241 253453
rect 6241 252677 6275 253453
rect 6337 253453 6485 253454
rect 6337 252677 6371 253453
rect 6371 252677 6451 253453
rect 6451 252677 6485 253453
rect 6547 253453 6695 253454
rect 6547 252677 6581 253453
rect 6581 252677 6661 253453
rect 6661 252677 6695 253453
rect 6757 253453 6905 253454
rect 6757 252677 6791 253453
rect 6791 252677 6871 253453
rect 6871 252677 6905 253453
rect 6967 253453 7115 253454
rect 6967 252677 7001 253453
rect 7001 252677 7081 253453
rect 7081 252677 7115 253453
rect 7177 253453 7325 253454
rect 7177 252677 7211 253453
rect 7211 252677 7291 253453
rect 7291 252677 7325 253453
rect 7387 253453 7535 253454
rect 7387 252677 7421 253453
rect 7421 252677 7501 253453
rect 7501 252677 7535 253453
rect 7597 253453 7745 253454
rect 7597 252677 7631 253453
rect 7631 252677 7711 253453
rect 7711 252677 7745 253453
rect 7807 253453 7955 253454
rect 7807 252677 7841 253453
rect 7841 252677 7921 253453
rect 7921 252677 7955 253453
rect 8017 253453 8165 253454
rect 8017 252677 8051 253453
rect 8051 252677 8131 253453
rect 8131 252677 8165 253453
rect 8227 253453 8375 253454
rect 8227 252677 8261 253453
rect 8261 252677 8341 253453
rect 8341 252677 8375 253453
rect 8437 253453 8585 253454
rect 8437 252677 8471 253453
rect 8471 252677 8551 253453
rect 8551 252677 8585 253453
rect 8647 253453 8795 253454
rect 8647 252677 8681 253453
rect 8681 252677 8761 253453
rect 8761 252677 8795 253453
rect 8857 253453 9005 253454
rect 8857 252677 8891 253453
rect 8891 252677 8971 253453
rect 8971 252677 9005 253453
rect 9067 253453 9215 253454
rect 9067 252677 9101 253453
rect 9101 252677 9181 253453
rect 9181 252677 9215 253453
rect 9277 253453 9425 253454
rect 9277 252677 9311 253453
rect 9311 252677 9391 253453
rect 9391 252677 9425 253453
rect 9487 253453 9635 253454
rect 9487 252677 9521 253453
rect 9521 252677 9601 253453
rect 9601 252677 9635 253453
rect 9697 253453 9845 253454
rect 9697 252677 9731 253453
rect 9731 252677 9811 253453
rect 9811 252677 9845 253453
rect 9907 253453 10055 253454
rect 9907 252677 9941 253453
rect 9941 252677 10021 253453
rect 10021 252677 10055 253453
rect 10117 253453 10265 253454
rect 10117 252677 10151 253453
rect 10151 252677 10231 253453
rect 10231 252677 10265 253453
rect 10327 253453 10475 253454
rect 10327 252677 10361 253453
rect 10361 252677 10441 253453
rect 10441 252677 10475 253453
rect 10537 253453 10685 253454
rect 10537 252677 10571 253453
rect 10571 252677 10651 253453
rect 10651 252677 10685 253453
rect 10747 253453 10895 253454
rect 10747 252677 10781 253453
rect 10781 252677 10861 253453
rect 10861 252677 10895 253453
rect 10957 253453 11105 253454
rect 10957 252677 10991 253453
rect 10991 252677 11071 253453
rect 11071 252677 11105 253453
rect 11167 253453 11315 253454
rect 11167 252677 11201 253453
rect 11201 252677 11281 253453
rect 11281 252677 11315 253453
rect 11377 253453 11525 253454
rect 11377 252677 11411 253453
rect 11411 252677 11491 253453
rect 11491 252677 11525 253453
rect 11587 253453 11735 253454
rect 11587 252677 11621 253453
rect 11621 252677 11701 253453
rect 11701 252677 11735 253453
rect 11797 253453 11945 253454
rect 11797 252677 11831 253453
rect 11831 252677 11911 253453
rect 11911 252677 11945 253453
rect 12007 253453 12155 253454
rect 12007 252677 12041 253453
rect 12041 252677 12121 253453
rect 12121 252677 12155 253453
rect 12217 253453 12365 253454
rect 12217 252677 12251 253453
rect 12251 252677 12331 253453
rect 12331 252677 12365 253453
rect 12427 253453 12575 253454
rect 12427 252677 12461 253453
rect 12461 252677 12541 253453
rect 12541 252677 12575 253453
rect 12637 253453 12785 253454
rect 12637 252677 12671 253453
rect 12671 252677 12751 253453
rect 12751 252677 12785 253453
rect 12847 253453 12995 253454
rect 12847 252677 12881 253453
rect 12881 252677 12961 253453
rect 12961 252677 12995 253453
rect 13057 253453 13205 253454
rect 13057 252677 13091 253453
rect 13091 252677 13171 253453
rect 13171 252677 13205 253453
rect 13267 253453 13415 253454
rect 13267 252677 13301 253453
rect 13301 252677 13381 253453
rect 13381 252677 13415 253453
rect 13477 253453 13625 253454
rect 13477 252677 13511 253453
rect 13511 252677 13591 253453
rect 13591 252677 13625 253453
rect 13687 253453 13835 253454
rect 13687 252677 13721 253453
rect 13721 252677 13801 253453
rect 13801 252677 13835 253453
rect 13897 253453 14045 253454
rect 13897 252677 13931 253453
rect 13931 252677 14011 253453
rect 14011 252677 14045 253453
rect 14107 253453 14255 253454
rect 14107 252677 14141 253453
rect 14141 252677 14221 253453
rect 14221 252677 14255 253453
rect 14317 253453 14465 253454
rect 14317 252677 14351 253453
rect 14351 252677 14431 253453
rect 14431 252677 14465 253453
rect 14527 253453 14675 253454
rect 14527 252677 14561 253453
rect 14561 252677 14641 253453
rect 14641 252677 14675 253453
rect 14737 253453 14885 253454
rect 14737 252677 14771 253453
rect 14771 252677 14851 253453
rect 14851 252677 14885 253453
rect 14947 253453 15095 253454
rect 14947 252677 14981 253453
rect 14981 252677 15061 253453
rect 15061 252677 15095 253453
rect 15157 253453 15305 253454
rect 15157 252677 15191 253453
rect 15191 252677 15271 253453
rect 15271 252677 15305 253453
rect 15367 253453 15515 253454
rect 15367 252677 15401 253453
rect 15401 252677 15481 253453
rect 15481 252677 15515 253453
rect 15577 253453 15725 253454
rect 15577 252677 15611 253453
rect 15611 252677 15691 253453
rect 15691 252677 15725 253453
rect 15787 253453 15935 253454
rect 15787 252677 15821 253453
rect 15821 252677 15901 253453
rect 15901 252677 15935 253453
rect 15997 253453 16145 253454
rect 15997 252677 16031 253453
rect 16031 252677 16111 253453
rect 16111 252677 16145 253453
rect 16207 253453 16355 253454
rect 16207 252677 16241 253453
rect 16241 252677 16321 253453
rect 16321 252677 16355 253453
rect 16417 253453 16565 253454
rect 16417 252677 16451 253453
rect 16451 252677 16531 253453
rect 16531 252677 16565 253453
rect 16627 253453 16775 253454
rect 16627 252677 16661 253453
rect 16661 252677 16741 253453
rect 16741 252677 16775 253453
rect 16837 253453 16985 253454
rect 16837 252677 16871 253453
rect 16871 252677 16951 253453
rect 16951 252677 16985 253453
rect 17047 253453 17195 253454
rect 17047 252677 17081 253453
rect 17081 252677 17161 253453
rect 17161 252677 17195 253453
rect 17257 253453 17405 253454
rect 17257 252677 17291 253453
rect 17291 252677 17371 253453
rect 17371 252677 17405 253453
rect 17467 253453 17615 253454
rect 17467 252677 17501 253453
rect 17501 252677 17581 253453
rect 17581 252677 17615 253453
rect 17677 253453 17825 253454
rect 17677 252677 17711 253453
rect 17711 252677 17791 253453
rect 17791 252677 17825 253453
rect 17887 253453 18035 253454
rect 17887 252677 17921 253453
rect 17921 252677 18001 253453
rect 18001 252677 18035 253453
rect 18097 253453 18245 253454
rect 18097 252677 18131 253453
rect 18131 252677 18211 253453
rect 18211 252677 18245 253453
rect 18307 253453 18455 253454
rect 18307 252677 18341 253453
rect 18341 252677 18421 253453
rect 18421 252677 18455 253453
rect 18517 253453 18665 253454
rect 18517 252677 18551 253453
rect 18551 252677 18631 253453
rect 18631 252677 18665 253453
rect 18727 253453 18875 253454
rect 18727 252677 18761 253453
rect 18761 252677 18841 253453
rect 18841 252677 18875 253453
rect 18937 253453 19085 253454
rect 18937 252677 18971 253453
rect 18971 252677 19051 253453
rect 19051 252677 19085 253453
rect 19147 253453 19295 253454
rect 19147 252677 19181 253453
rect 19181 252677 19261 253453
rect 19261 252677 19295 253453
rect 19357 253453 19505 253454
rect 19357 252677 19391 253453
rect 19391 252677 19471 253453
rect 19471 252677 19505 253453
rect 19567 253453 19715 253454
rect 19567 252677 19601 253453
rect 19601 252677 19681 253453
rect 19681 252677 19715 253453
rect 19777 253453 19925 253454
rect 19777 252677 19811 253453
rect 19811 252677 19891 253453
rect 19891 252677 19925 253453
rect 19987 253453 20135 253454
rect 19987 252677 20021 253453
rect 20021 252677 20101 253453
rect 20101 252677 20135 253453
rect 20197 253453 20345 253454
rect 20197 252677 20231 253453
rect 20231 252677 20311 253453
rect 20311 252677 20345 253453
rect 20407 253453 20555 253454
rect 20407 252677 20441 253453
rect 20441 252677 20521 253453
rect 20521 252677 20555 253453
rect 20617 253453 20765 253454
rect 20617 252677 20651 253453
rect 20651 252677 20731 253453
rect 20731 252677 20765 253453
rect 20827 253453 20975 253454
rect 20827 252677 20861 253453
rect 20861 252677 20941 253453
rect 20941 252677 20975 253453
rect 21037 253453 21185 253454
rect 21037 252677 21071 253453
rect 21071 252677 21151 253453
rect 21151 252677 21185 253453
rect 21247 253453 21395 253454
rect 21247 252677 21281 253453
rect 21281 252677 21361 253453
rect 21361 252677 21395 253453
rect 21457 253453 21605 253454
rect 21457 252677 21491 253453
rect 21491 252677 21571 253453
rect 21571 252677 21605 253453
rect 21667 253453 21815 253454
rect 21667 252677 21701 253453
rect 21701 252677 21781 253453
rect 21781 252677 21815 253453
rect 21877 253453 22025 253454
rect 21877 252677 21911 253453
rect 21911 252677 21991 253453
rect 21991 252677 22025 253453
rect 22087 253453 22235 253454
rect 22087 252677 22121 253453
rect 22121 252677 22201 253453
rect 22201 252677 22235 253453
rect 22297 253453 22445 253454
rect 22297 252677 22331 253453
rect 22331 252677 22411 253453
rect 22411 252677 22445 253453
rect 22507 253453 22655 253454
rect 22507 252677 22541 253453
rect 22541 252677 22621 253453
rect 22621 252677 22655 253453
rect 22717 253453 22865 253454
rect 22717 252677 22751 253453
rect 22751 252677 22831 253453
rect 22831 252677 22865 253453
rect 22927 253453 23075 253454
rect 22927 252677 22961 253453
rect 22961 252677 23041 253453
rect 23041 252677 23075 253453
rect 23137 253453 23285 253454
rect 23137 252677 23171 253453
rect 23171 252677 23251 253453
rect 23251 252677 23285 253453
rect 23347 253453 23495 253454
rect 23347 252677 23381 253453
rect 23381 252677 23461 253453
rect 23461 252677 23495 253453
rect 23557 253453 23705 253454
rect 23557 252677 23591 253453
rect 23591 252677 23671 253453
rect 23671 252677 23705 253453
rect 23767 253453 23915 253454
rect 23767 252677 23801 253453
rect 23801 252677 23881 253453
rect 23881 252677 23915 253453
rect 23977 253453 24125 253454
rect 23977 252677 24011 253453
rect 24011 252677 24091 253453
rect 24091 252677 24125 253453
rect 24187 253453 24335 253454
rect 24187 252677 24221 253453
rect 24221 252677 24301 253453
rect 24301 252677 24335 253453
rect 24397 253453 24545 253454
rect 24397 252677 24431 253453
rect 24431 252677 24511 253453
rect 24511 252677 24545 253453
rect 24607 253453 24755 253454
rect 24607 252677 24641 253453
rect 24641 252677 24721 253453
rect 24721 252677 24755 253453
rect 24817 253453 24965 253454
rect 24817 252677 24851 253453
rect 24851 252677 24931 253453
rect 24931 252677 24965 253453
rect 25027 253453 25175 253454
rect 25027 252677 25061 253453
rect 25061 252677 25141 253453
rect 25141 252677 25175 253453
rect 25237 253453 25385 253454
rect 25237 252677 25271 253453
rect 25271 252677 25351 253453
rect 25351 252677 25385 253453
rect 25447 253453 25595 253454
rect 25447 252677 25481 253453
rect 25481 252677 25561 253453
rect 25561 252677 25595 253453
rect 25657 253453 25805 253454
rect 25657 252677 25691 253453
rect 25691 252677 25771 253453
rect 25771 252677 25805 253453
rect 25867 253453 26015 253454
rect 25867 252677 25901 253453
rect 25901 252677 25981 253453
rect 25981 252677 26015 253453
rect 26077 253453 26225 253454
rect 26077 252677 26111 253453
rect 26111 252677 26191 253453
rect 26191 252677 26225 253453
rect 26287 253453 26435 253454
rect 26287 252677 26321 253453
rect 26321 252677 26401 253453
rect 26401 252677 26435 253453
rect 26497 253453 26645 253454
rect 26497 252677 26531 253453
rect 26531 252677 26611 253453
rect 26611 252677 26645 253453
rect 26707 253453 26855 253454
rect 26707 252677 26741 253453
rect 26741 252677 26821 253453
rect 26821 252677 26855 253453
rect 26917 253453 27065 253454
rect 26917 252677 26951 253453
rect 26951 252677 27031 253453
rect 27031 252677 27065 253453
rect 27127 253453 27275 253454
rect 27127 252677 27161 253453
rect 27161 252677 27241 253453
rect 27241 252677 27275 253453
rect -4069 251641 -4049 252417
rect -4049 251641 -4015 252417
rect -3953 251641 -3919 252417
rect -3919 251641 -3839 252417
rect -3839 251641 -3805 252417
rect -3743 251641 -3709 252417
rect -3709 251641 -3629 252417
rect -3629 251641 -3595 252417
rect -3533 252417 -3385 252418
rect -3533 251641 -3499 252417
rect -3499 251641 -3419 252417
rect -3419 251641 -3385 252417
rect -3323 252417 -3175 252418
rect -3323 251641 -3289 252417
rect -3289 251641 -3209 252417
rect -3209 251641 -3175 252417
rect -3113 252417 -2965 252418
rect -3113 251641 -3079 252417
rect -3079 251641 -2999 252417
rect -2999 251641 -2965 252417
rect -2903 252417 -2755 252418
rect -2903 251641 -2869 252417
rect -2869 251641 -2789 252417
rect -2789 251641 -2755 252417
rect -2693 252417 -2545 252418
rect -2693 251641 -2659 252417
rect -2659 251641 -2579 252417
rect -2579 251641 -2545 252417
rect -2483 252417 -2335 252418
rect -2483 251641 -2449 252417
rect -2449 251641 -2369 252417
rect -2369 251641 -2335 252417
rect -2273 252417 -2125 252418
rect -2273 251641 -2239 252417
rect -2239 251641 -2159 252417
rect -2159 251641 -2125 252417
rect -2063 252417 -1915 252418
rect -2063 251641 -2029 252417
rect -2029 251641 -1949 252417
rect -1949 251641 -1915 252417
rect -1853 252417 -1705 252418
rect -1853 251641 -1819 252417
rect -1819 251641 -1739 252417
rect -1739 251641 -1705 252417
rect -1643 252417 -1495 252418
rect -1643 251641 -1609 252417
rect -1609 251641 -1529 252417
rect -1529 251641 -1495 252417
rect -1433 252417 -1285 252418
rect -1433 251641 -1399 252417
rect -1399 251641 -1319 252417
rect -1319 251641 -1285 252417
rect -1223 252417 -1075 252418
rect -1223 251641 -1189 252417
rect -1189 251641 -1109 252417
rect -1109 251641 -1075 252417
rect -1013 252417 -865 252418
rect -1013 251641 -979 252417
rect -979 251641 -899 252417
rect -899 251641 -865 252417
rect -803 252417 -655 252418
rect -803 251641 -769 252417
rect -769 251641 -689 252417
rect -689 251641 -655 252417
rect -593 252417 -445 252418
rect -593 251641 -559 252417
rect -559 251641 -479 252417
rect -479 251641 -445 252417
rect -383 252417 -235 252418
rect -383 251641 -349 252417
rect -349 251641 -269 252417
rect -269 251641 -235 252417
rect -173 252417 -25 252418
rect -173 251641 -139 252417
rect -139 251641 -59 252417
rect -59 251641 -25 252417
rect 37 252417 185 252418
rect 37 251641 71 252417
rect 71 251641 151 252417
rect 151 251641 185 252417
rect 247 252417 395 252418
rect 247 251641 281 252417
rect 281 251641 361 252417
rect 361 251641 395 252417
rect 457 252417 605 252418
rect 457 251641 491 252417
rect 491 251641 571 252417
rect 571 251641 605 252417
rect 667 252417 815 252418
rect 667 251641 701 252417
rect 701 251641 781 252417
rect 781 251641 815 252417
rect 877 252417 1025 252418
rect 877 251641 911 252417
rect 911 251641 991 252417
rect 991 251641 1025 252417
rect 1087 252417 1235 252418
rect 1087 251641 1121 252417
rect 1121 251641 1201 252417
rect 1201 251641 1235 252417
rect 1297 252417 1445 252418
rect 1297 251641 1331 252417
rect 1331 251641 1411 252417
rect 1411 251641 1445 252417
rect 1507 252417 1655 252418
rect 1507 251641 1541 252417
rect 1541 251641 1621 252417
rect 1621 251641 1655 252417
rect 1717 252417 1865 252418
rect 1717 251641 1751 252417
rect 1751 251641 1831 252417
rect 1831 251641 1865 252417
rect 1927 252417 2075 252418
rect 1927 251641 1961 252417
rect 1961 251641 2041 252417
rect 2041 251641 2075 252417
rect 2137 252417 2285 252418
rect 2137 251641 2171 252417
rect 2171 251641 2251 252417
rect 2251 251641 2285 252417
rect 2347 252417 2495 252418
rect 2347 251641 2381 252417
rect 2381 251641 2461 252417
rect 2461 251641 2495 252417
rect 2557 252417 2705 252418
rect 2557 251641 2591 252417
rect 2591 251641 2671 252417
rect 2671 251641 2705 252417
rect 2767 252417 2915 252418
rect 2767 251641 2801 252417
rect 2801 251641 2881 252417
rect 2881 251641 2915 252417
rect 2977 252417 3125 252418
rect 2977 251641 3011 252417
rect 3011 251641 3091 252417
rect 3091 251641 3125 252417
rect 3187 252417 3335 252418
rect 3187 251641 3221 252417
rect 3221 251641 3301 252417
rect 3301 251641 3335 252417
rect 3397 252417 3545 252418
rect 3397 251641 3431 252417
rect 3431 251641 3511 252417
rect 3511 251641 3545 252417
rect 3607 252417 3755 252418
rect 3607 251641 3641 252417
rect 3641 251641 3721 252417
rect 3721 251641 3755 252417
rect 3817 252417 3965 252418
rect 3817 251641 3851 252417
rect 3851 251641 3931 252417
rect 3931 251641 3965 252417
rect 4027 252417 4175 252418
rect 4027 251641 4061 252417
rect 4061 251641 4141 252417
rect 4141 251641 4175 252417
rect 4237 252417 4385 252418
rect 4237 251641 4271 252417
rect 4271 251641 4351 252417
rect 4351 251641 4385 252417
rect 4447 252417 4595 252418
rect 4447 251641 4481 252417
rect 4481 251641 4561 252417
rect 4561 251641 4595 252417
rect 4657 252417 4805 252418
rect 4657 251641 4691 252417
rect 4691 251641 4771 252417
rect 4771 251641 4805 252417
rect 4867 252417 5015 252418
rect 4867 251641 4901 252417
rect 4901 251641 4981 252417
rect 4981 251641 5015 252417
rect 5077 252417 5225 252418
rect 5077 251641 5111 252417
rect 5111 251641 5191 252417
rect 5191 251641 5225 252417
rect 5287 252417 5435 252418
rect 5287 251641 5321 252417
rect 5321 251641 5401 252417
rect 5401 251641 5435 252417
rect 5497 252417 5645 252418
rect 5497 251641 5531 252417
rect 5531 251641 5611 252417
rect 5611 251641 5645 252417
rect 5707 252417 5855 252418
rect 5707 251641 5741 252417
rect 5741 251641 5821 252417
rect 5821 251641 5855 252417
rect 5917 252417 6065 252418
rect 5917 251641 5951 252417
rect 5951 251641 6031 252417
rect 6031 251641 6065 252417
rect 6127 252417 6275 252418
rect 6127 251641 6161 252417
rect 6161 251641 6241 252417
rect 6241 251641 6275 252417
rect 6337 252417 6485 252418
rect 6337 251641 6371 252417
rect 6371 251641 6451 252417
rect 6451 251641 6485 252417
rect 6547 252417 6695 252418
rect 6547 251641 6581 252417
rect 6581 251641 6661 252417
rect 6661 251641 6695 252417
rect 6757 252417 6905 252418
rect 6757 251641 6791 252417
rect 6791 251641 6871 252417
rect 6871 251641 6905 252417
rect 6967 252417 7115 252418
rect 6967 251641 7001 252417
rect 7001 251641 7081 252417
rect 7081 251641 7115 252417
rect 7177 252417 7325 252418
rect 7177 251641 7211 252417
rect 7211 251641 7291 252417
rect 7291 251641 7325 252417
rect 7387 252417 7535 252418
rect 7387 251641 7421 252417
rect 7421 251641 7501 252417
rect 7501 251641 7535 252417
rect 7597 252417 7745 252418
rect 7597 251641 7631 252417
rect 7631 251641 7711 252417
rect 7711 251641 7745 252417
rect 7807 252417 7955 252418
rect 7807 251641 7841 252417
rect 7841 251641 7921 252417
rect 7921 251641 7955 252417
rect 8017 252417 8165 252418
rect 8017 251641 8051 252417
rect 8051 251641 8131 252417
rect 8131 251641 8165 252417
rect 8227 252417 8375 252418
rect 8227 251641 8261 252417
rect 8261 251641 8341 252417
rect 8341 251641 8375 252417
rect 8437 252417 8585 252418
rect 8437 251641 8471 252417
rect 8471 251641 8551 252417
rect 8551 251641 8585 252417
rect 8647 252417 8795 252418
rect 8647 251641 8681 252417
rect 8681 251641 8761 252417
rect 8761 251641 8795 252417
rect 8857 252417 9005 252418
rect 8857 251641 8891 252417
rect 8891 251641 8971 252417
rect 8971 251641 9005 252417
rect 9067 252417 9215 252418
rect 9067 251641 9101 252417
rect 9101 251641 9181 252417
rect 9181 251641 9215 252417
rect 9277 252417 9425 252418
rect 9277 251641 9311 252417
rect 9311 251641 9391 252417
rect 9391 251641 9425 252417
rect 9487 252417 9635 252418
rect 9487 251641 9521 252417
rect 9521 251641 9601 252417
rect 9601 251641 9635 252417
rect 9697 252417 9845 252418
rect 9697 251641 9731 252417
rect 9731 251641 9811 252417
rect 9811 251641 9845 252417
rect 9907 252417 10055 252418
rect 9907 251641 9941 252417
rect 9941 251641 10021 252417
rect 10021 251641 10055 252417
rect 10117 252417 10265 252418
rect 10117 251641 10151 252417
rect 10151 251641 10231 252417
rect 10231 251641 10265 252417
rect 10327 252417 10475 252418
rect 10327 251641 10361 252417
rect 10361 251641 10441 252417
rect 10441 251641 10475 252417
rect 10537 252417 10685 252418
rect 10537 251641 10571 252417
rect 10571 251641 10651 252417
rect 10651 251641 10685 252417
rect 10747 252417 10895 252418
rect 10747 251641 10781 252417
rect 10781 251641 10861 252417
rect 10861 251641 10895 252417
rect 10957 252417 11105 252418
rect 10957 251641 10991 252417
rect 10991 251641 11071 252417
rect 11071 251641 11105 252417
rect 11167 252417 11315 252418
rect 11167 251641 11201 252417
rect 11201 251641 11281 252417
rect 11281 251641 11315 252417
rect 11377 252417 11525 252418
rect 11377 251641 11411 252417
rect 11411 251641 11491 252417
rect 11491 251641 11525 252417
rect 11587 252417 11735 252418
rect 11587 251641 11621 252417
rect 11621 251641 11701 252417
rect 11701 251641 11735 252417
rect 11797 252417 11945 252418
rect 11797 251641 11831 252417
rect 11831 251641 11911 252417
rect 11911 251641 11945 252417
rect 12007 252417 12155 252418
rect 12007 251641 12041 252417
rect 12041 251641 12121 252417
rect 12121 251641 12155 252417
rect 12217 252417 12365 252418
rect 12217 251641 12251 252417
rect 12251 251641 12331 252417
rect 12331 251641 12365 252417
rect 12427 252417 12575 252418
rect 12427 251641 12461 252417
rect 12461 251641 12541 252417
rect 12541 251641 12575 252417
rect 12637 252417 12785 252418
rect 12637 251641 12671 252417
rect 12671 251641 12751 252417
rect 12751 251641 12785 252417
rect 12847 252417 12995 252418
rect 12847 251641 12881 252417
rect 12881 251641 12961 252417
rect 12961 251641 12995 252417
rect 13057 252417 13205 252418
rect 13057 251641 13091 252417
rect 13091 251641 13171 252417
rect 13171 251641 13205 252417
rect 13267 252417 13415 252418
rect 13267 251641 13301 252417
rect 13301 251641 13381 252417
rect 13381 251641 13415 252417
rect 13477 252417 13625 252418
rect 13477 251641 13511 252417
rect 13511 251641 13591 252417
rect 13591 251641 13625 252417
rect 13687 252417 13835 252418
rect 13687 251641 13721 252417
rect 13721 251641 13801 252417
rect 13801 251641 13835 252417
rect 13897 252417 14045 252418
rect 13897 251641 13931 252417
rect 13931 251641 14011 252417
rect 14011 251641 14045 252417
rect 14107 252417 14255 252418
rect 14107 251641 14141 252417
rect 14141 251641 14221 252417
rect 14221 251641 14255 252417
rect 14317 252417 14465 252418
rect 14317 251641 14351 252417
rect 14351 251641 14431 252417
rect 14431 251641 14465 252417
rect 14527 252417 14675 252418
rect 14527 251641 14561 252417
rect 14561 251641 14641 252417
rect 14641 251641 14675 252417
rect 14737 252417 14885 252418
rect 14737 251641 14771 252417
rect 14771 251641 14851 252417
rect 14851 251641 14885 252417
rect 14947 252417 15095 252418
rect 14947 251641 14981 252417
rect 14981 251641 15061 252417
rect 15061 251641 15095 252417
rect 15157 252417 15305 252418
rect 15157 251641 15191 252417
rect 15191 251641 15271 252417
rect 15271 251641 15305 252417
rect 15367 252417 15515 252418
rect 15367 251641 15401 252417
rect 15401 251641 15481 252417
rect 15481 251641 15515 252417
rect 15577 252417 15725 252418
rect 15577 251641 15611 252417
rect 15611 251641 15691 252417
rect 15691 251641 15725 252417
rect 15787 252417 15935 252418
rect 15787 251641 15821 252417
rect 15821 251641 15901 252417
rect 15901 251641 15935 252417
rect 15997 252417 16145 252418
rect 15997 251641 16031 252417
rect 16031 251641 16111 252417
rect 16111 251641 16145 252417
rect 16207 252417 16355 252418
rect 16207 251641 16241 252417
rect 16241 251641 16321 252417
rect 16321 251641 16355 252417
rect 16417 252417 16565 252418
rect 16417 251641 16451 252417
rect 16451 251641 16531 252417
rect 16531 251641 16565 252417
rect 16627 252417 16775 252418
rect 16627 251641 16661 252417
rect 16661 251641 16741 252417
rect 16741 251641 16775 252417
rect 16837 252417 16985 252418
rect 16837 251641 16871 252417
rect 16871 251641 16951 252417
rect 16951 251641 16985 252417
rect 17047 252417 17195 252418
rect 17047 251641 17081 252417
rect 17081 251641 17161 252417
rect 17161 251641 17195 252417
rect 17257 252417 17405 252418
rect 17257 251641 17291 252417
rect 17291 251641 17371 252417
rect 17371 251641 17405 252417
rect 17467 252417 17615 252418
rect 17467 251641 17501 252417
rect 17501 251641 17581 252417
rect 17581 251641 17615 252417
rect 17677 252417 17825 252418
rect 17677 251641 17711 252417
rect 17711 251641 17791 252417
rect 17791 251641 17825 252417
rect 17887 252417 18035 252418
rect 17887 251641 17921 252417
rect 17921 251641 18001 252417
rect 18001 251641 18035 252417
rect 18097 252417 18245 252418
rect 18097 251641 18131 252417
rect 18131 251641 18211 252417
rect 18211 251641 18245 252417
rect 18307 252417 18455 252418
rect 18307 251641 18341 252417
rect 18341 251641 18421 252417
rect 18421 251641 18455 252417
rect 18517 252417 18665 252418
rect 18517 251641 18551 252417
rect 18551 251641 18631 252417
rect 18631 251641 18665 252417
rect 18727 252417 18875 252418
rect 18727 251641 18761 252417
rect 18761 251641 18841 252417
rect 18841 251641 18875 252417
rect 18937 252417 19085 252418
rect 18937 251641 18971 252417
rect 18971 251641 19051 252417
rect 19051 251641 19085 252417
rect 19147 252417 19295 252418
rect 19147 251641 19181 252417
rect 19181 251641 19261 252417
rect 19261 251641 19295 252417
rect 19357 252417 19505 252418
rect 19357 251641 19391 252417
rect 19391 251641 19471 252417
rect 19471 251641 19505 252417
rect 19567 252417 19715 252418
rect 19567 251641 19601 252417
rect 19601 251641 19681 252417
rect 19681 251641 19715 252417
rect 19777 252417 19925 252418
rect 19777 251641 19811 252417
rect 19811 251641 19891 252417
rect 19891 251641 19925 252417
rect 19987 252417 20135 252418
rect 19987 251641 20021 252417
rect 20021 251641 20101 252417
rect 20101 251641 20135 252417
rect 20197 252417 20345 252418
rect 20197 251641 20231 252417
rect 20231 251641 20311 252417
rect 20311 251641 20345 252417
rect 20407 252417 20555 252418
rect 20407 251641 20441 252417
rect 20441 251641 20521 252417
rect 20521 251641 20555 252417
rect 20617 252417 20765 252418
rect 20617 251641 20651 252417
rect 20651 251641 20731 252417
rect 20731 251641 20765 252417
rect 20827 252417 20975 252418
rect 20827 251641 20861 252417
rect 20861 251641 20941 252417
rect 20941 251641 20975 252417
rect 21037 252417 21185 252418
rect 21037 251641 21071 252417
rect 21071 251641 21151 252417
rect 21151 251641 21185 252417
rect 21247 252417 21395 252418
rect 21247 251641 21281 252417
rect 21281 251641 21361 252417
rect 21361 251641 21395 252417
rect 21457 252417 21605 252418
rect 21457 251641 21491 252417
rect 21491 251641 21571 252417
rect 21571 251641 21605 252417
rect 21667 252417 21815 252418
rect 21667 251641 21701 252417
rect 21701 251641 21781 252417
rect 21781 251641 21815 252417
rect 21877 252417 22025 252418
rect 21877 251641 21911 252417
rect 21911 251641 21991 252417
rect 21991 251641 22025 252417
rect 22087 252417 22235 252418
rect 22087 251641 22121 252417
rect 22121 251641 22201 252417
rect 22201 251641 22235 252417
rect 22297 252417 22445 252418
rect 22297 251641 22331 252417
rect 22331 251641 22411 252417
rect 22411 251641 22445 252417
rect 22507 252417 22655 252418
rect 22507 251641 22541 252417
rect 22541 251641 22621 252417
rect 22621 251641 22655 252417
rect 22717 252417 22865 252418
rect 22717 251641 22751 252417
rect 22751 251641 22831 252417
rect 22831 251641 22865 252417
rect 22927 252417 23075 252418
rect 22927 251641 22961 252417
rect 22961 251641 23041 252417
rect 23041 251641 23075 252417
rect 23137 252417 23285 252418
rect 23137 251641 23171 252417
rect 23171 251641 23251 252417
rect 23251 251641 23285 252417
rect 23347 252417 23495 252418
rect 23347 251641 23381 252417
rect 23381 251641 23461 252417
rect 23461 251641 23495 252417
rect 23557 252417 23705 252418
rect 23557 251641 23591 252417
rect 23591 251641 23671 252417
rect 23671 251641 23705 252417
rect 23767 252417 23915 252418
rect 23767 251641 23801 252417
rect 23801 251641 23881 252417
rect 23881 251641 23915 252417
rect 23977 252417 24125 252418
rect 23977 251641 24011 252417
rect 24011 251641 24091 252417
rect 24091 251641 24125 252417
rect 24187 252417 24335 252418
rect 24187 251641 24221 252417
rect 24221 251641 24301 252417
rect 24301 251641 24335 252417
rect 24397 252417 24545 252418
rect 24397 251641 24431 252417
rect 24431 251641 24511 252417
rect 24511 251641 24545 252417
rect 24607 252417 24755 252418
rect 24607 251641 24641 252417
rect 24641 251641 24721 252417
rect 24721 251641 24755 252417
rect 24817 252417 24965 252418
rect 24817 251641 24851 252417
rect 24851 251641 24931 252417
rect 24931 251641 24965 252417
rect 25027 252417 25175 252418
rect 25027 251641 25061 252417
rect 25061 251641 25141 252417
rect 25141 251641 25175 252417
rect 25237 252417 25385 252418
rect 25237 251641 25271 252417
rect 25271 251641 25351 252417
rect 25351 251641 25385 252417
rect 25447 252417 25595 252418
rect 25447 251641 25481 252417
rect 25481 251641 25561 252417
rect 25561 251641 25595 252417
rect 25657 252417 25805 252418
rect 25657 251641 25691 252417
rect 25691 251641 25771 252417
rect 25771 251641 25805 252417
rect 25867 252417 26015 252418
rect 25867 251641 25901 252417
rect 25901 251641 25981 252417
rect 25981 251641 26015 252417
rect 26077 252417 26225 252418
rect 26077 251641 26111 252417
rect 26111 251641 26191 252417
rect 26191 251641 26225 252417
rect 26287 252417 26435 252418
rect 26287 251641 26321 252417
rect 26321 251641 26401 252417
rect 26401 251641 26435 252417
rect 26497 252417 26645 252418
rect 26497 251641 26531 252417
rect 26531 251641 26611 252417
rect 26611 251641 26645 252417
rect 26707 252417 26855 252418
rect 26707 251641 26741 252417
rect 26741 251641 26821 252417
rect 26821 251641 26855 252417
rect 26917 252417 27065 252418
rect 26917 251641 26951 252417
rect 26951 251641 27031 252417
rect 27031 251641 27065 252417
rect 27127 252417 27275 252418
rect 27127 251641 27161 252417
rect 27161 251641 27241 252417
rect 27241 251641 27275 252417
rect -4069 250605 -4049 251381
rect -4049 250605 -4015 251381
rect -3953 250605 -3919 251381
rect -3919 250605 -3839 251381
rect -3839 250605 -3805 251381
rect -3743 250605 -3709 251381
rect -3709 250605 -3629 251381
rect -3629 250605 -3595 251381
rect -3533 251381 -3385 251382
rect -3533 250605 -3499 251381
rect -3499 250605 -3419 251381
rect -3419 250605 -3385 251381
rect -3323 251381 -3175 251382
rect -3323 250605 -3289 251381
rect -3289 250605 -3209 251381
rect -3209 250605 -3175 251381
rect -3113 251381 -2965 251382
rect -3113 250605 -3079 251381
rect -3079 250605 -2999 251381
rect -2999 250605 -2965 251381
rect -2903 251381 -2755 251382
rect -2903 250605 -2869 251381
rect -2869 250605 -2789 251381
rect -2789 250605 -2755 251381
rect -2693 251381 -2545 251382
rect -2693 250605 -2659 251381
rect -2659 250605 -2579 251381
rect -2579 250605 -2545 251381
rect -2483 251381 -2335 251382
rect -2483 250605 -2449 251381
rect -2449 250605 -2369 251381
rect -2369 250605 -2335 251381
rect -2273 251381 -2125 251382
rect -2273 250605 -2239 251381
rect -2239 250605 -2159 251381
rect -2159 250605 -2125 251381
rect -2063 251381 -1915 251382
rect -2063 250605 -2029 251381
rect -2029 250605 -1949 251381
rect -1949 250605 -1915 251381
rect -1853 251381 -1705 251382
rect -1853 250605 -1819 251381
rect -1819 250605 -1739 251381
rect -1739 250605 -1705 251381
rect -1643 251381 -1495 251382
rect -1643 250605 -1609 251381
rect -1609 250605 -1529 251381
rect -1529 250605 -1495 251381
rect -1433 251381 -1285 251382
rect -1433 250605 -1399 251381
rect -1399 250605 -1319 251381
rect -1319 250605 -1285 251381
rect -1223 251381 -1075 251382
rect -1223 250605 -1189 251381
rect -1189 250605 -1109 251381
rect -1109 250605 -1075 251381
rect -1013 251381 -865 251382
rect -1013 250605 -979 251381
rect -979 250605 -899 251381
rect -899 250605 -865 251381
rect -803 251381 -655 251382
rect -803 250605 -769 251381
rect -769 250605 -689 251381
rect -689 250605 -655 251381
rect -593 251381 -445 251382
rect -593 250605 -559 251381
rect -559 250605 -479 251381
rect -479 250605 -445 251381
rect -383 251381 -235 251382
rect -383 250605 -349 251381
rect -349 250605 -269 251381
rect -269 250605 -235 251381
rect -173 251381 -25 251382
rect -173 250605 -139 251381
rect -139 250605 -59 251381
rect -59 250605 -25 251381
rect 37 251381 185 251382
rect 37 250605 71 251381
rect 71 250605 151 251381
rect 151 250605 185 251381
rect 247 251381 395 251382
rect 247 250605 281 251381
rect 281 250605 361 251381
rect 361 250605 395 251381
rect 457 251381 605 251382
rect 457 250605 491 251381
rect 491 250605 571 251381
rect 571 250605 605 251381
rect 667 251381 815 251382
rect 667 250605 701 251381
rect 701 250605 781 251381
rect 781 250605 815 251381
rect 877 251381 1025 251382
rect 877 250605 911 251381
rect 911 250605 991 251381
rect 991 250605 1025 251381
rect 1087 251381 1235 251382
rect 1087 250605 1121 251381
rect 1121 250605 1201 251381
rect 1201 250605 1235 251381
rect 1297 251381 1445 251382
rect 1297 250605 1331 251381
rect 1331 250605 1411 251381
rect 1411 250605 1445 251381
rect 1507 251381 1655 251382
rect 1507 250605 1541 251381
rect 1541 250605 1621 251381
rect 1621 250605 1655 251381
rect 1717 251381 1865 251382
rect 1717 250605 1751 251381
rect 1751 250605 1831 251381
rect 1831 250605 1865 251381
rect 1927 251381 2075 251382
rect 1927 250605 1961 251381
rect 1961 250605 2041 251381
rect 2041 250605 2075 251381
rect 2137 251381 2285 251382
rect 2137 250605 2171 251381
rect 2171 250605 2251 251381
rect 2251 250605 2285 251381
rect 2347 251381 2495 251382
rect 2347 250605 2381 251381
rect 2381 250605 2461 251381
rect 2461 250605 2495 251381
rect 2557 251381 2705 251382
rect 2557 250605 2591 251381
rect 2591 250605 2671 251381
rect 2671 250605 2705 251381
rect 2767 251381 2915 251382
rect 2767 250605 2801 251381
rect 2801 250605 2881 251381
rect 2881 250605 2915 251381
rect 2977 251381 3125 251382
rect 2977 250605 3011 251381
rect 3011 250605 3091 251381
rect 3091 250605 3125 251381
rect 3187 251381 3335 251382
rect 3187 250605 3221 251381
rect 3221 250605 3301 251381
rect 3301 250605 3335 251381
rect 3397 251381 3545 251382
rect 3397 250605 3431 251381
rect 3431 250605 3511 251381
rect 3511 250605 3545 251381
rect 3607 251381 3755 251382
rect 3607 250605 3641 251381
rect 3641 250605 3721 251381
rect 3721 250605 3755 251381
rect 3817 251381 3965 251382
rect 3817 250605 3851 251381
rect 3851 250605 3931 251381
rect 3931 250605 3965 251381
rect 4027 251381 4175 251382
rect 4027 250605 4061 251381
rect 4061 250605 4141 251381
rect 4141 250605 4175 251381
rect 4237 251381 4385 251382
rect 4237 250605 4271 251381
rect 4271 250605 4351 251381
rect 4351 250605 4385 251381
rect 4447 251381 4595 251382
rect 4447 250605 4481 251381
rect 4481 250605 4561 251381
rect 4561 250605 4595 251381
rect 4657 251381 4805 251382
rect 4657 250605 4691 251381
rect 4691 250605 4771 251381
rect 4771 250605 4805 251381
rect 4867 251381 5015 251382
rect 4867 250605 4901 251381
rect 4901 250605 4981 251381
rect 4981 250605 5015 251381
rect 5077 251381 5225 251382
rect 5077 250605 5111 251381
rect 5111 250605 5191 251381
rect 5191 250605 5225 251381
rect 5287 251381 5435 251382
rect 5287 250605 5321 251381
rect 5321 250605 5401 251381
rect 5401 250605 5435 251381
rect 5497 251381 5645 251382
rect 5497 250605 5531 251381
rect 5531 250605 5611 251381
rect 5611 250605 5645 251381
rect 5707 251381 5855 251382
rect 5707 250605 5741 251381
rect 5741 250605 5821 251381
rect 5821 250605 5855 251381
rect 5917 251381 6065 251382
rect 5917 250605 5951 251381
rect 5951 250605 6031 251381
rect 6031 250605 6065 251381
rect 6127 251381 6275 251382
rect 6127 250605 6161 251381
rect 6161 250605 6241 251381
rect 6241 250605 6275 251381
rect 6337 251381 6485 251382
rect 6337 250605 6371 251381
rect 6371 250605 6451 251381
rect 6451 250605 6485 251381
rect 6547 251381 6695 251382
rect 6547 250605 6581 251381
rect 6581 250605 6661 251381
rect 6661 250605 6695 251381
rect 6757 251381 6905 251382
rect 6757 250605 6791 251381
rect 6791 250605 6871 251381
rect 6871 250605 6905 251381
rect 6967 251381 7115 251382
rect 6967 250605 7001 251381
rect 7001 250605 7081 251381
rect 7081 250605 7115 251381
rect 7177 251381 7325 251382
rect 7177 250605 7211 251381
rect 7211 250605 7291 251381
rect 7291 250605 7325 251381
rect 7387 251381 7535 251382
rect 7387 250605 7421 251381
rect 7421 250605 7501 251381
rect 7501 250605 7535 251381
rect 7597 251381 7745 251382
rect 7597 250605 7631 251381
rect 7631 250605 7711 251381
rect 7711 250605 7745 251381
rect 7807 251381 7955 251382
rect 7807 250605 7841 251381
rect 7841 250605 7921 251381
rect 7921 250605 7955 251381
rect 8017 251381 8165 251382
rect 8017 250605 8051 251381
rect 8051 250605 8131 251381
rect 8131 250605 8165 251381
rect 8227 251381 8375 251382
rect 8227 250605 8261 251381
rect 8261 250605 8341 251381
rect 8341 250605 8375 251381
rect 8437 251381 8585 251382
rect 8437 250605 8471 251381
rect 8471 250605 8551 251381
rect 8551 250605 8585 251381
rect 8647 251381 8795 251382
rect 8647 250605 8681 251381
rect 8681 250605 8761 251381
rect 8761 250605 8795 251381
rect 8857 251381 9005 251382
rect 8857 250605 8891 251381
rect 8891 250605 8971 251381
rect 8971 250605 9005 251381
rect 9067 251381 9215 251382
rect 9067 250605 9101 251381
rect 9101 250605 9181 251381
rect 9181 250605 9215 251381
rect 9277 251381 9425 251382
rect 9277 250605 9311 251381
rect 9311 250605 9391 251381
rect 9391 250605 9425 251381
rect 9487 251381 9635 251382
rect 9487 250605 9521 251381
rect 9521 250605 9601 251381
rect 9601 250605 9635 251381
rect 9697 251381 9845 251382
rect 9697 250605 9731 251381
rect 9731 250605 9811 251381
rect 9811 250605 9845 251381
rect 9907 251381 10055 251382
rect 9907 250605 9941 251381
rect 9941 250605 10021 251381
rect 10021 250605 10055 251381
rect 10117 251381 10265 251382
rect 10117 250605 10151 251381
rect 10151 250605 10231 251381
rect 10231 250605 10265 251381
rect 10327 251381 10475 251382
rect 10327 250605 10361 251381
rect 10361 250605 10441 251381
rect 10441 250605 10475 251381
rect 10537 251381 10685 251382
rect 10537 250605 10571 251381
rect 10571 250605 10651 251381
rect 10651 250605 10685 251381
rect 10747 251381 10895 251382
rect 10747 250605 10781 251381
rect 10781 250605 10861 251381
rect 10861 250605 10895 251381
rect 10957 251381 11105 251382
rect 10957 250605 10991 251381
rect 10991 250605 11071 251381
rect 11071 250605 11105 251381
rect 11167 251381 11315 251382
rect 11167 250605 11201 251381
rect 11201 250605 11281 251381
rect 11281 250605 11315 251381
rect 11377 251381 11525 251382
rect 11377 250605 11411 251381
rect 11411 250605 11491 251381
rect 11491 250605 11525 251381
rect 11587 251381 11735 251382
rect 11587 250605 11621 251381
rect 11621 250605 11701 251381
rect 11701 250605 11735 251381
rect 11797 251381 11945 251382
rect 11797 250605 11831 251381
rect 11831 250605 11911 251381
rect 11911 250605 11945 251381
rect 12007 251381 12155 251382
rect 12007 250605 12041 251381
rect 12041 250605 12121 251381
rect 12121 250605 12155 251381
rect 12217 251381 12365 251382
rect 12217 250605 12251 251381
rect 12251 250605 12331 251381
rect 12331 250605 12365 251381
rect 12427 251381 12575 251382
rect 12427 250605 12461 251381
rect 12461 250605 12541 251381
rect 12541 250605 12575 251381
rect 12637 251381 12785 251382
rect 12637 250605 12671 251381
rect 12671 250605 12751 251381
rect 12751 250605 12785 251381
rect 12847 251381 12995 251382
rect 12847 250605 12881 251381
rect 12881 250605 12961 251381
rect 12961 250605 12995 251381
rect 13057 251381 13205 251382
rect 13057 250605 13091 251381
rect 13091 250605 13171 251381
rect 13171 250605 13205 251381
rect 13267 251381 13415 251382
rect 13267 250605 13301 251381
rect 13301 250605 13381 251381
rect 13381 250605 13415 251381
rect 13477 251381 13625 251382
rect 13477 250605 13511 251381
rect 13511 250605 13591 251381
rect 13591 250605 13625 251381
rect 13687 251381 13835 251382
rect 13687 250605 13721 251381
rect 13721 250605 13801 251381
rect 13801 250605 13835 251381
rect 13897 251381 14045 251382
rect 13897 250605 13931 251381
rect 13931 250605 14011 251381
rect 14011 250605 14045 251381
rect 14107 251381 14255 251382
rect 14107 250605 14141 251381
rect 14141 250605 14221 251381
rect 14221 250605 14255 251381
rect 14317 251381 14465 251382
rect 14317 250605 14351 251381
rect 14351 250605 14431 251381
rect 14431 250605 14465 251381
rect 14527 251381 14675 251382
rect 14527 250605 14561 251381
rect 14561 250605 14641 251381
rect 14641 250605 14675 251381
rect 14737 251381 14885 251382
rect 14737 250605 14771 251381
rect 14771 250605 14851 251381
rect 14851 250605 14885 251381
rect 14947 251381 15095 251382
rect 14947 250605 14981 251381
rect 14981 250605 15061 251381
rect 15061 250605 15095 251381
rect 15157 251381 15305 251382
rect 15157 250605 15191 251381
rect 15191 250605 15271 251381
rect 15271 250605 15305 251381
rect 15367 251381 15515 251382
rect 15367 250605 15401 251381
rect 15401 250605 15481 251381
rect 15481 250605 15515 251381
rect 15577 251381 15725 251382
rect 15577 250605 15611 251381
rect 15611 250605 15691 251381
rect 15691 250605 15725 251381
rect 15787 251381 15935 251382
rect 15787 250605 15821 251381
rect 15821 250605 15901 251381
rect 15901 250605 15935 251381
rect 15997 251381 16145 251382
rect 15997 250605 16031 251381
rect 16031 250605 16111 251381
rect 16111 250605 16145 251381
rect 16207 251381 16355 251382
rect 16207 250605 16241 251381
rect 16241 250605 16321 251381
rect 16321 250605 16355 251381
rect 16417 251381 16565 251382
rect 16417 250605 16451 251381
rect 16451 250605 16531 251381
rect 16531 250605 16565 251381
rect 16627 251381 16775 251382
rect 16627 250605 16661 251381
rect 16661 250605 16741 251381
rect 16741 250605 16775 251381
rect 16837 251381 16985 251382
rect 16837 250605 16871 251381
rect 16871 250605 16951 251381
rect 16951 250605 16985 251381
rect 17047 251381 17195 251382
rect 17047 250605 17081 251381
rect 17081 250605 17161 251381
rect 17161 250605 17195 251381
rect 17257 251381 17405 251382
rect 17257 250605 17291 251381
rect 17291 250605 17371 251381
rect 17371 250605 17405 251381
rect 17467 251381 17615 251382
rect 17467 250605 17501 251381
rect 17501 250605 17581 251381
rect 17581 250605 17615 251381
rect 17677 251381 17825 251382
rect 17677 250605 17711 251381
rect 17711 250605 17791 251381
rect 17791 250605 17825 251381
rect 17887 251381 18035 251382
rect 17887 250605 17921 251381
rect 17921 250605 18001 251381
rect 18001 250605 18035 251381
rect 18097 251381 18245 251382
rect 18097 250605 18131 251381
rect 18131 250605 18211 251381
rect 18211 250605 18245 251381
rect 18307 251381 18455 251382
rect 18307 250605 18341 251381
rect 18341 250605 18421 251381
rect 18421 250605 18455 251381
rect 18517 251381 18665 251382
rect 18517 250605 18551 251381
rect 18551 250605 18631 251381
rect 18631 250605 18665 251381
rect 18727 251381 18875 251382
rect 18727 250605 18761 251381
rect 18761 250605 18841 251381
rect 18841 250605 18875 251381
rect 18937 251381 19085 251382
rect 18937 250605 18971 251381
rect 18971 250605 19051 251381
rect 19051 250605 19085 251381
rect 19147 251381 19295 251382
rect 19147 250605 19181 251381
rect 19181 250605 19261 251381
rect 19261 250605 19295 251381
rect 19357 251381 19505 251382
rect 19357 250605 19391 251381
rect 19391 250605 19471 251381
rect 19471 250605 19505 251381
rect 19567 251381 19715 251382
rect 19567 250605 19601 251381
rect 19601 250605 19681 251381
rect 19681 250605 19715 251381
rect 19777 251381 19925 251382
rect 19777 250605 19811 251381
rect 19811 250605 19891 251381
rect 19891 250605 19925 251381
rect 19987 251381 20135 251382
rect 19987 250605 20021 251381
rect 20021 250605 20101 251381
rect 20101 250605 20135 251381
rect 20197 251381 20345 251382
rect 20197 250605 20231 251381
rect 20231 250605 20311 251381
rect 20311 250605 20345 251381
rect 20407 251381 20555 251382
rect 20407 250605 20441 251381
rect 20441 250605 20521 251381
rect 20521 250605 20555 251381
rect 20617 251381 20765 251382
rect 20617 250605 20651 251381
rect 20651 250605 20731 251381
rect 20731 250605 20765 251381
rect 20827 251381 20975 251382
rect 20827 250605 20861 251381
rect 20861 250605 20941 251381
rect 20941 250605 20975 251381
rect 21037 251381 21185 251382
rect 21037 250605 21071 251381
rect 21071 250605 21151 251381
rect 21151 250605 21185 251381
rect 21247 251381 21395 251382
rect 21247 250605 21281 251381
rect 21281 250605 21361 251381
rect 21361 250605 21395 251381
rect 21457 251381 21605 251382
rect 21457 250605 21491 251381
rect 21491 250605 21571 251381
rect 21571 250605 21605 251381
rect 21667 251381 21815 251382
rect 21667 250605 21701 251381
rect 21701 250605 21781 251381
rect 21781 250605 21815 251381
rect 21877 251381 22025 251382
rect 21877 250605 21911 251381
rect 21911 250605 21991 251381
rect 21991 250605 22025 251381
rect 22087 251381 22235 251382
rect 22087 250605 22121 251381
rect 22121 250605 22201 251381
rect 22201 250605 22235 251381
rect 22297 251381 22445 251382
rect 22297 250605 22331 251381
rect 22331 250605 22411 251381
rect 22411 250605 22445 251381
rect 22507 251381 22655 251382
rect 22507 250605 22541 251381
rect 22541 250605 22621 251381
rect 22621 250605 22655 251381
rect 22717 251381 22865 251382
rect 22717 250605 22751 251381
rect 22751 250605 22831 251381
rect 22831 250605 22865 251381
rect 22927 251381 23075 251382
rect 22927 250605 22961 251381
rect 22961 250605 23041 251381
rect 23041 250605 23075 251381
rect 23137 251381 23285 251382
rect 23137 250605 23171 251381
rect 23171 250605 23251 251381
rect 23251 250605 23285 251381
rect 23347 251381 23495 251382
rect 23347 250605 23381 251381
rect 23381 250605 23461 251381
rect 23461 250605 23495 251381
rect 23557 251381 23705 251382
rect 23557 250605 23591 251381
rect 23591 250605 23671 251381
rect 23671 250605 23705 251381
rect 23767 251381 23915 251382
rect 23767 250605 23801 251381
rect 23801 250605 23881 251381
rect 23881 250605 23915 251381
rect 23977 251381 24125 251382
rect 23977 250605 24011 251381
rect 24011 250605 24091 251381
rect 24091 250605 24125 251381
rect 24187 251381 24335 251382
rect 24187 250605 24221 251381
rect 24221 250605 24301 251381
rect 24301 250605 24335 251381
rect 24397 251381 24545 251382
rect 24397 250605 24431 251381
rect 24431 250605 24511 251381
rect 24511 250605 24545 251381
rect 24607 251381 24755 251382
rect 24607 250605 24641 251381
rect 24641 250605 24721 251381
rect 24721 250605 24755 251381
rect 24817 251381 24965 251382
rect 24817 250605 24851 251381
rect 24851 250605 24931 251381
rect 24931 250605 24965 251381
rect 25027 251381 25175 251382
rect 25027 250605 25061 251381
rect 25061 250605 25141 251381
rect 25141 250605 25175 251381
rect 25237 251381 25385 251382
rect 25237 250605 25271 251381
rect 25271 250605 25351 251381
rect 25351 250605 25385 251381
rect 25447 251381 25595 251382
rect 25447 250605 25481 251381
rect 25481 250605 25561 251381
rect 25561 250605 25595 251381
rect 25657 251381 25805 251382
rect 25657 250605 25691 251381
rect 25691 250605 25771 251381
rect 25771 250605 25805 251381
rect 25867 251381 26015 251382
rect 25867 250605 25901 251381
rect 25901 250605 25981 251381
rect 25981 250605 26015 251381
rect 26077 251381 26225 251382
rect 26077 250605 26111 251381
rect 26111 250605 26191 251381
rect 26191 250605 26225 251381
rect 26287 251381 26435 251382
rect 26287 250605 26321 251381
rect 26321 250605 26401 251381
rect 26401 250605 26435 251381
rect 26497 251381 26645 251382
rect 26497 250605 26531 251381
rect 26531 250605 26611 251381
rect 26611 250605 26645 251381
rect 26707 251381 26855 251382
rect 26707 250605 26741 251381
rect 26741 250605 26821 251381
rect 26821 250605 26855 251381
rect 26917 251381 27065 251382
rect 26917 250605 26951 251381
rect 26951 250605 27031 251381
rect 27031 250605 27065 251381
rect 27127 251381 27275 251382
rect 27127 250605 27161 251381
rect 27161 250605 27241 251381
rect 27241 250605 27275 251381
rect -4069 249569 -4049 250345
rect -4049 249569 -4015 250345
rect -3953 249569 -3919 250345
rect -3919 249569 -3839 250345
rect -3839 249569 -3805 250345
rect -3743 249569 -3709 250345
rect -3709 249569 -3629 250345
rect -3629 249569 -3595 250345
rect -3533 250345 -3385 250346
rect -3533 249569 -3499 250345
rect -3499 249569 -3419 250345
rect -3419 249569 -3385 250345
rect -3323 250345 -3175 250346
rect -3323 249569 -3289 250345
rect -3289 249569 -3209 250345
rect -3209 249569 -3175 250345
rect -3113 250345 -2965 250346
rect -3113 249569 -3079 250345
rect -3079 249569 -2999 250345
rect -2999 249569 -2965 250345
rect -2903 250345 -2755 250346
rect -2903 249569 -2869 250345
rect -2869 249569 -2789 250345
rect -2789 249569 -2755 250345
rect -2693 250345 -2545 250346
rect -2693 249569 -2659 250345
rect -2659 249569 -2579 250345
rect -2579 249569 -2545 250345
rect -2483 250345 -2335 250346
rect -2483 249569 -2449 250345
rect -2449 249569 -2369 250345
rect -2369 249569 -2335 250345
rect -2273 250345 -2125 250346
rect -2273 249569 -2239 250345
rect -2239 249569 -2159 250345
rect -2159 249569 -2125 250345
rect -2063 250345 -1915 250346
rect -2063 249569 -2029 250345
rect -2029 249569 -1949 250345
rect -1949 249569 -1915 250345
rect -1853 250345 -1705 250346
rect -1853 249569 -1819 250345
rect -1819 249569 -1739 250345
rect -1739 249569 -1705 250345
rect -1643 250345 -1495 250346
rect -1643 249569 -1609 250345
rect -1609 249569 -1529 250345
rect -1529 249569 -1495 250345
rect -1433 250345 -1285 250346
rect -1433 249569 -1399 250345
rect -1399 249569 -1319 250345
rect -1319 249569 -1285 250345
rect -1223 250345 -1075 250346
rect -1223 249569 -1189 250345
rect -1189 249569 -1109 250345
rect -1109 249569 -1075 250345
rect -1013 250345 -865 250346
rect -1013 249569 -979 250345
rect -979 249569 -899 250345
rect -899 249569 -865 250345
rect -803 250345 -655 250346
rect -803 249569 -769 250345
rect -769 249569 -689 250345
rect -689 249569 -655 250345
rect -593 250345 -445 250346
rect -593 249569 -559 250345
rect -559 249569 -479 250345
rect -479 249569 -445 250345
rect -383 250345 -235 250346
rect -383 249569 -349 250345
rect -349 249569 -269 250345
rect -269 249569 -235 250345
rect -173 250345 -25 250346
rect -173 249569 -139 250345
rect -139 249569 -59 250345
rect -59 249569 -25 250345
rect 37 250345 185 250346
rect 37 249569 71 250345
rect 71 249569 151 250345
rect 151 249569 185 250345
rect 247 250345 395 250346
rect 247 249569 281 250345
rect 281 249569 361 250345
rect 361 249569 395 250345
rect 457 250345 605 250346
rect 457 249569 491 250345
rect 491 249569 571 250345
rect 571 249569 605 250345
rect 667 250345 815 250346
rect 667 249569 701 250345
rect 701 249569 781 250345
rect 781 249569 815 250345
rect 877 250345 1025 250346
rect 877 249569 911 250345
rect 911 249569 991 250345
rect 991 249569 1025 250345
rect 1087 250345 1235 250346
rect 1087 249569 1121 250345
rect 1121 249569 1201 250345
rect 1201 249569 1235 250345
rect 1297 250345 1445 250346
rect 1297 249569 1331 250345
rect 1331 249569 1411 250345
rect 1411 249569 1445 250345
rect 1507 250345 1655 250346
rect 1507 249569 1541 250345
rect 1541 249569 1621 250345
rect 1621 249569 1655 250345
rect 1717 250345 1865 250346
rect 1717 249569 1751 250345
rect 1751 249569 1831 250345
rect 1831 249569 1865 250345
rect 1927 250345 2075 250346
rect 1927 249569 1961 250345
rect 1961 249569 2041 250345
rect 2041 249569 2075 250345
rect 2137 250345 2285 250346
rect 2137 249569 2171 250345
rect 2171 249569 2251 250345
rect 2251 249569 2285 250345
rect 2347 250345 2495 250346
rect 2347 249569 2381 250345
rect 2381 249569 2461 250345
rect 2461 249569 2495 250345
rect 2557 250345 2705 250346
rect 2557 249569 2591 250345
rect 2591 249569 2671 250345
rect 2671 249569 2705 250345
rect 2767 250345 2915 250346
rect 2767 249569 2801 250345
rect 2801 249569 2881 250345
rect 2881 249569 2915 250345
rect 2977 250345 3125 250346
rect 2977 249569 3011 250345
rect 3011 249569 3091 250345
rect 3091 249569 3125 250345
rect 3187 250345 3335 250346
rect 3187 249569 3221 250345
rect 3221 249569 3301 250345
rect 3301 249569 3335 250345
rect 3397 250345 3545 250346
rect 3397 249569 3431 250345
rect 3431 249569 3511 250345
rect 3511 249569 3545 250345
rect 3607 250345 3755 250346
rect 3607 249569 3641 250345
rect 3641 249569 3721 250345
rect 3721 249569 3755 250345
rect 3817 250345 3965 250346
rect 3817 249569 3851 250345
rect 3851 249569 3931 250345
rect 3931 249569 3965 250345
rect 4027 250345 4175 250346
rect 4027 249569 4061 250345
rect 4061 249569 4141 250345
rect 4141 249569 4175 250345
rect 4237 250345 4385 250346
rect 4237 249569 4271 250345
rect 4271 249569 4351 250345
rect 4351 249569 4385 250345
rect 4447 250345 4595 250346
rect 4447 249569 4481 250345
rect 4481 249569 4561 250345
rect 4561 249569 4595 250345
rect 4657 250345 4805 250346
rect 4657 249569 4691 250345
rect 4691 249569 4771 250345
rect 4771 249569 4805 250345
rect 4867 250345 5015 250346
rect 4867 249569 4901 250345
rect 4901 249569 4981 250345
rect 4981 249569 5015 250345
rect 5077 250345 5225 250346
rect 5077 249569 5111 250345
rect 5111 249569 5191 250345
rect 5191 249569 5225 250345
rect 5287 250345 5435 250346
rect 5287 249569 5321 250345
rect 5321 249569 5401 250345
rect 5401 249569 5435 250345
rect 5497 250345 5645 250346
rect 5497 249569 5531 250345
rect 5531 249569 5611 250345
rect 5611 249569 5645 250345
rect 5707 250345 5855 250346
rect 5707 249569 5741 250345
rect 5741 249569 5821 250345
rect 5821 249569 5855 250345
rect 5917 250345 6065 250346
rect 5917 249569 5951 250345
rect 5951 249569 6031 250345
rect 6031 249569 6065 250345
rect 6127 250345 6275 250346
rect 6127 249569 6161 250345
rect 6161 249569 6241 250345
rect 6241 249569 6275 250345
rect 6337 250345 6485 250346
rect 6337 249569 6371 250345
rect 6371 249569 6451 250345
rect 6451 249569 6485 250345
rect 6547 250345 6695 250346
rect 6547 249569 6581 250345
rect 6581 249569 6661 250345
rect 6661 249569 6695 250345
rect 6757 250345 6905 250346
rect 6757 249569 6791 250345
rect 6791 249569 6871 250345
rect 6871 249569 6905 250345
rect 6967 250345 7115 250346
rect 6967 249569 7001 250345
rect 7001 249569 7081 250345
rect 7081 249569 7115 250345
rect 7177 250345 7325 250346
rect 7177 249569 7211 250345
rect 7211 249569 7291 250345
rect 7291 249569 7325 250345
rect 7387 250345 7535 250346
rect 7387 249569 7421 250345
rect 7421 249569 7501 250345
rect 7501 249569 7535 250345
rect 7597 250345 7745 250346
rect 7597 249569 7631 250345
rect 7631 249569 7711 250345
rect 7711 249569 7745 250345
rect 7807 250345 7955 250346
rect 7807 249569 7841 250345
rect 7841 249569 7921 250345
rect 7921 249569 7955 250345
rect 8017 250345 8165 250346
rect 8017 249569 8051 250345
rect 8051 249569 8131 250345
rect 8131 249569 8165 250345
rect 8227 250345 8375 250346
rect 8227 249569 8261 250345
rect 8261 249569 8341 250345
rect 8341 249569 8375 250345
rect 8437 250345 8585 250346
rect 8437 249569 8471 250345
rect 8471 249569 8551 250345
rect 8551 249569 8585 250345
rect 8647 250345 8795 250346
rect 8647 249569 8681 250345
rect 8681 249569 8761 250345
rect 8761 249569 8795 250345
rect 8857 250345 9005 250346
rect 8857 249569 8891 250345
rect 8891 249569 8971 250345
rect 8971 249569 9005 250345
rect 9067 250345 9215 250346
rect 9067 249569 9101 250345
rect 9101 249569 9181 250345
rect 9181 249569 9215 250345
rect 9277 250345 9425 250346
rect 9277 249569 9311 250345
rect 9311 249569 9391 250345
rect 9391 249569 9425 250345
rect 9487 250345 9635 250346
rect 9487 249569 9521 250345
rect 9521 249569 9601 250345
rect 9601 249569 9635 250345
rect 9697 250345 9845 250346
rect 9697 249569 9731 250345
rect 9731 249569 9811 250345
rect 9811 249569 9845 250345
rect 9907 250345 10055 250346
rect 9907 249569 9941 250345
rect 9941 249569 10021 250345
rect 10021 249569 10055 250345
rect 10117 250345 10265 250346
rect 10117 249569 10151 250345
rect 10151 249569 10231 250345
rect 10231 249569 10265 250345
rect 10327 250345 10475 250346
rect 10327 249569 10361 250345
rect 10361 249569 10441 250345
rect 10441 249569 10475 250345
rect 10537 250345 10685 250346
rect 10537 249569 10571 250345
rect 10571 249569 10651 250345
rect 10651 249569 10685 250345
rect 10747 250345 10895 250346
rect 10747 249569 10781 250345
rect 10781 249569 10861 250345
rect 10861 249569 10895 250345
rect 10957 250345 11105 250346
rect 10957 249569 10991 250345
rect 10991 249569 11071 250345
rect 11071 249569 11105 250345
rect 11167 250345 11315 250346
rect 11167 249569 11201 250345
rect 11201 249569 11281 250345
rect 11281 249569 11315 250345
rect 11377 250345 11525 250346
rect 11377 249569 11411 250345
rect 11411 249569 11491 250345
rect 11491 249569 11525 250345
rect 11587 250345 11735 250346
rect 11587 249569 11621 250345
rect 11621 249569 11701 250345
rect 11701 249569 11735 250345
rect 11797 250345 11945 250346
rect 11797 249569 11831 250345
rect 11831 249569 11911 250345
rect 11911 249569 11945 250345
rect 12007 250345 12155 250346
rect 12007 249569 12041 250345
rect 12041 249569 12121 250345
rect 12121 249569 12155 250345
rect 12217 250345 12365 250346
rect 12217 249569 12251 250345
rect 12251 249569 12331 250345
rect 12331 249569 12365 250345
rect 12427 250345 12575 250346
rect 12427 249569 12461 250345
rect 12461 249569 12541 250345
rect 12541 249569 12575 250345
rect 12637 250345 12785 250346
rect 12637 249569 12671 250345
rect 12671 249569 12751 250345
rect 12751 249569 12785 250345
rect 12847 250345 12995 250346
rect 12847 249569 12881 250345
rect 12881 249569 12961 250345
rect 12961 249569 12995 250345
rect 13057 250345 13205 250346
rect 13057 249569 13091 250345
rect 13091 249569 13171 250345
rect 13171 249569 13205 250345
rect 13267 250345 13415 250346
rect 13267 249569 13301 250345
rect 13301 249569 13381 250345
rect 13381 249569 13415 250345
rect 13477 250345 13625 250346
rect 13477 249569 13511 250345
rect 13511 249569 13591 250345
rect 13591 249569 13625 250345
rect 13687 250345 13835 250346
rect 13687 249569 13721 250345
rect 13721 249569 13801 250345
rect 13801 249569 13835 250345
rect 13897 250345 14045 250346
rect 13897 249569 13931 250345
rect 13931 249569 14011 250345
rect 14011 249569 14045 250345
rect 14107 250345 14255 250346
rect 14107 249569 14141 250345
rect 14141 249569 14221 250345
rect 14221 249569 14255 250345
rect 14317 250345 14465 250346
rect 14317 249569 14351 250345
rect 14351 249569 14431 250345
rect 14431 249569 14465 250345
rect 14527 250345 14675 250346
rect 14527 249569 14561 250345
rect 14561 249569 14641 250345
rect 14641 249569 14675 250345
rect 14737 250345 14885 250346
rect 14737 249569 14771 250345
rect 14771 249569 14851 250345
rect 14851 249569 14885 250345
rect 14947 250345 15095 250346
rect 14947 249569 14981 250345
rect 14981 249569 15061 250345
rect 15061 249569 15095 250345
rect 15157 250345 15305 250346
rect 15157 249569 15191 250345
rect 15191 249569 15271 250345
rect 15271 249569 15305 250345
rect 15367 250345 15515 250346
rect 15367 249569 15401 250345
rect 15401 249569 15481 250345
rect 15481 249569 15515 250345
rect 15577 250345 15725 250346
rect 15577 249569 15611 250345
rect 15611 249569 15691 250345
rect 15691 249569 15725 250345
rect 15787 250345 15935 250346
rect 15787 249569 15821 250345
rect 15821 249569 15901 250345
rect 15901 249569 15935 250345
rect 15997 250345 16145 250346
rect 15997 249569 16031 250345
rect 16031 249569 16111 250345
rect 16111 249569 16145 250345
rect 16207 250345 16355 250346
rect 16207 249569 16241 250345
rect 16241 249569 16321 250345
rect 16321 249569 16355 250345
rect 16417 250345 16565 250346
rect 16417 249569 16451 250345
rect 16451 249569 16531 250345
rect 16531 249569 16565 250345
rect 16627 250345 16775 250346
rect 16627 249569 16661 250345
rect 16661 249569 16741 250345
rect 16741 249569 16775 250345
rect 16837 250345 16985 250346
rect 16837 249569 16871 250345
rect 16871 249569 16951 250345
rect 16951 249569 16985 250345
rect 17047 250345 17195 250346
rect 17047 249569 17081 250345
rect 17081 249569 17161 250345
rect 17161 249569 17195 250345
rect 17257 250345 17405 250346
rect 17257 249569 17291 250345
rect 17291 249569 17371 250345
rect 17371 249569 17405 250345
rect 17467 250345 17615 250346
rect 17467 249569 17501 250345
rect 17501 249569 17581 250345
rect 17581 249569 17615 250345
rect 17677 250345 17825 250346
rect 17677 249569 17711 250345
rect 17711 249569 17791 250345
rect 17791 249569 17825 250345
rect 17887 250345 18035 250346
rect 17887 249569 17921 250345
rect 17921 249569 18001 250345
rect 18001 249569 18035 250345
rect 18097 250345 18245 250346
rect 18097 249569 18131 250345
rect 18131 249569 18211 250345
rect 18211 249569 18245 250345
rect 18307 250345 18455 250346
rect 18307 249569 18341 250345
rect 18341 249569 18421 250345
rect 18421 249569 18455 250345
rect 18517 250345 18665 250346
rect 18517 249569 18551 250345
rect 18551 249569 18631 250345
rect 18631 249569 18665 250345
rect 18727 250345 18875 250346
rect 18727 249569 18761 250345
rect 18761 249569 18841 250345
rect 18841 249569 18875 250345
rect 18937 250345 19085 250346
rect 18937 249569 18971 250345
rect 18971 249569 19051 250345
rect 19051 249569 19085 250345
rect 19147 250345 19295 250346
rect 19147 249569 19181 250345
rect 19181 249569 19261 250345
rect 19261 249569 19295 250345
rect 19357 250345 19505 250346
rect 19357 249569 19391 250345
rect 19391 249569 19471 250345
rect 19471 249569 19505 250345
rect 19567 250345 19715 250346
rect 19567 249569 19601 250345
rect 19601 249569 19681 250345
rect 19681 249569 19715 250345
rect 19777 250345 19925 250346
rect 19777 249569 19811 250345
rect 19811 249569 19891 250345
rect 19891 249569 19925 250345
rect 19987 250345 20135 250346
rect 19987 249569 20021 250345
rect 20021 249569 20101 250345
rect 20101 249569 20135 250345
rect 20197 250345 20345 250346
rect 20197 249569 20231 250345
rect 20231 249569 20311 250345
rect 20311 249569 20345 250345
rect 20407 250345 20555 250346
rect 20407 249569 20441 250345
rect 20441 249569 20521 250345
rect 20521 249569 20555 250345
rect 20617 250345 20765 250346
rect 20617 249569 20651 250345
rect 20651 249569 20731 250345
rect 20731 249569 20765 250345
rect 20827 250345 20975 250346
rect 20827 249569 20861 250345
rect 20861 249569 20941 250345
rect 20941 249569 20975 250345
rect 21037 250345 21185 250346
rect 21037 249569 21071 250345
rect 21071 249569 21151 250345
rect 21151 249569 21185 250345
rect 21247 250345 21395 250346
rect 21247 249569 21281 250345
rect 21281 249569 21361 250345
rect 21361 249569 21395 250345
rect 21457 250345 21605 250346
rect 21457 249569 21491 250345
rect 21491 249569 21571 250345
rect 21571 249569 21605 250345
rect 21667 250345 21815 250346
rect 21667 249569 21701 250345
rect 21701 249569 21781 250345
rect 21781 249569 21815 250345
rect 21877 250345 22025 250346
rect 21877 249569 21911 250345
rect 21911 249569 21991 250345
rect 21991 249569 22025 250345
rect 22087 250345 22235 250346
rect 22087 249569 22121 250345
rect 22121 249569 22201 250345
rect 22201 249569 22235 250345
rect 22297 250345 22445 250346
rect 22297 249569 22331 250345
rect 22331 249569 22411 250345
rect 22411 249569 22445 250345
rect 22507 250345 22655 250346
rect 22507 249569 22541 250345
rect 22541 249569 22621 250345
rect 22621 249569 22655 250345
rect 22717 250345 22865 250346
rect 22717 249569 22751 250345
rect 22751 249569 22831 250345
rect 22831 249569 22865 250345
rect 22927 250345 23075 250346
rect 22927 249569 22961 250345
rect 22961 249569 23041 250345
rect 23041 249569 23075 250345
rect 23137 250345 23285 250346
rect 23137 249569 23171 250345
rect 23171 249569 23251 250345
rect 23251 249569 23285 250345
rect 23347 250345 23495 250346
rect 23347 249569 23381 250345
rect 23381 249569 23461 250345
rect 23461 249569 23495 250345
rect 23557 250345 23705 250346
rect 23557 249569 23591 250345
rect 23591 249569 23671 250345
rect 23671 249569 23705 250345
rect 23767 250345 23915 250346
rect 23767 249569 23801 250345
rect 23801 249569 23881 250345
rect 23881 249569 23915 250345
rect 23977 250345 24125 250346
rect 23977 249569 24011 250345
rect 24011 249569 24091 250345
rect 24091 249569 24125 250345
rect 24187 250345 24335 250346
rect 24187 249569 24221 250345
rect 24221 249569 24301 250345
rect 24301 249569 24335 250345
rect 24397 250345 24545 250346
rect 24397 249569 24431 250345
rect 24431 249569 24511 250345
rect 24511 249569 24545 250345
rect 24607 250345 24755 250346
rect 24607 249569 24641 250345
rect 24641 249569 24721 250345
rect 24721 249569 24755 250345
rect 24817 250345 24965 250346
rect 24817 249569 24851 250345
rect 24851 249569 24931 250345
rect 24931 249569 24965 250345
rect 25027 250345 25175 250346
rect 25027 249569 25061 250345
rect 25061 249569 25141 250345
rect 25141 249569 25175 250345
rect 25237 250345 25385 250346
rect 25237 249569 25271 250345
rect 25271 249569 25351 250345
rect 25351 249569 25385 250345
rect 25447 250345 25595 250346
rect 25447 249569 25481 250345
rect 25481 249569 25561 250345
rect 25561 249569 25595 250345
rect 25657 250345 25805 250346
rect 25657 249569 25691 250345
rect 25691 249569 25771 250345
rect 25771 249569 25805 250345
rect 25867 250345 26015 250346
rect 25867 249569 25901 250345
rect 25901 249569 25981 250345
rect 25981 249569 26015 250345
rect 26077 250345 26225 250346
rect 26077 249569 26111 250345
rect 26111 249569 26191 250345
rect 26191 249569 26225 250345
rect 26287 250345 26435 250346
rect 26287 249569 26321 250345
rect 26321 249569 26401 250345
rect 26401 249569 26435 250345
rect 26497 250345 26645 250346
rect 26497 249569 26531 250345
rect 26531 249569 26611 250345
rect 26611 249569 26645 250345
rect 26707 250345 26855 250346
rect 26707 249569 26741 250345
rect 26741 249569 26821 250345
rect 26821 249569 26855 250345
rect 26917 250345 27065 250346
rect 26917 249569 26951 250345
rect 26951 249569 27031 250345
rect 27031 249569 27065 250345
rect 27127 250345 27275 250346
rect 27127 249569 27161 250345
rect 27161 249569 27241 250345
rect 27241 249569 27275 250345
rect -4075 248404 -4049 249180
rect -4049 248404 -4015 249180
rect -3953 248404 -3919 249180
rect -3919 248404 -3839 249180
rect -3839 248404 -3805 249180
rect -3743 248404 -3709 249180
rect -3709 248404 -3629 249180
rect -3629 248404 -3595 249180
rect -3533 249180 -3385 249181
rect -3533 248404 -3499 249180
rect -3499 248404 -3419 249180
rect -3419 248404 -3385 249180
rect -3323 249180 -3175 249181
rect -3323 248404 -3289 249180
rect -3289 248404 -3209 249180
rect -3209 248404 -3175 249180
rect -3113 249180 -2965 249181
rect -3113 248404 -3079 249180
rect -3079 248404 -2999 249180
rect -2999 248404 -2965 249180
rect -2903 249180 -2755 249181
rect -2903 248404 -2869 249180
rect -2869 248404 -2789 249180
rect -2789 248404 -2755 249180
rect -2693 249180 -2545 249181
rect -2693 248404 -2659 249180
rect -2659 248404 -2579 249180
rect -2579 248404 -2545 249180
rect -2483 249180 -2335 249181
rect -2483 248404 -2449 249180
rect -2449 248404 -2369 249180
rect -2369 248404 -2335 249180
rect -2273 249180 -2125 249181
rect -2273 248404 -2239 249180
rect -2239 248404 -2159 249180
rect -2159 248404 -2125 249180
rect -2063 249180 -1915 249181
rect -2063 248404 -2029 249180
rect -2029 248404 -1949 249180
rect -1949 248404 -1915 249180
rect -1853 249180 -1705 249181
rect -1853 248404 -1819 249180
rect -1819 248404 -1739 249180
rect -1739 248404 -1705 249180
rect -1643 249180 -1495 249181
rect -1643 248404 -1609 249180
rect -1609 248404 -1529 249180
rect -1529 248404 -1495 249180
rect -1433 249180 -1285 249181
rect -1433 248404 -1399 249180
rect -1399 248404 -1319 249180
rect -1319 248404 -1285 249180
rect -1223 249180 -1075 249181
rect -1223 248404 -1189 249180
rect -1189 248404 -1109 249180
rect -1109 248404 -1075 249180
rect -1013 249180 -865 249181
rect -1013 248404 -979 249180
rect -979 248404 -899 249180
rect -899 248404 -865 249180
rect -803 249180 -655 249181
rect -803 248404 -769 249180
rect -769 248404 -689 249180
rect -689 248404 -655 249180
rect -593 249180 -445 249181
rect -593 248404 -559 249180
rect -559 248404 -479 249180
rect -479 248404 -445 249180
rect -383 249180 -235 249181
rect -383 248404 -349 249180
rect -349 248404 -269 249180
rect -269 248404 -235 249180
rect -173 249180 -25 249181
rect -173 248404 -139 249180
rect -139 248404 -59 249180
rect -59 248404 -25 249180
rect 37 249180 185 249181
rect 37 248404 71 249180
rect 71 248404 151 249180
rect 151 248404 185 249180
rect 247 249180 395 249181
rect 247 248404 281 249180
rect 281 248404 361 249180
rect 361 248404 395 249180
rect 457 249180 605 249181
rect 457 248404 491 249180
rect 491 248404 571 249180
rect 571 248404 605 249180
rect 667 249180 815 249181
rect 667 248404 701 249180
rect 701 248404 781 249180
rect 781 248404 815 249180
rect 877 249180 1025 249181
rect 877 248404 911 249180
rect 911 248404 991 249180
rect 991 248404 1025 249180
rect 1087 249180 1235 249181
rect 1087 248404 1121 249180
rect 1121 248404 1201 249180
rect 1201 248404 1235 249180
rect 1297 249180 1445 249181
rect 1297 248404 1331 249180
rect 1331 248404 1411 249180
rect 1411 248404 1445 249180
rect 1507 249180 1655 249181
rect 1507 248404 1541 249180
rect 1541 248404 1621 249180
rect 1621 248404 1655 249180
rect 1717 249180 1865 249181
rect 1717 248404 1751 249180
rect 1751 248404 1831 249180
rect 1831 248404 1865 249180
rect 1927 249180 2075 249181
rect 1927 248404 1961 249180
rect 1961 248404 2041 249180
rect 2041 248404 2075 249180
rect 2137 249180 2285 249181
rect 2137 248404 2171 249180
rect 2171 248404 2251 249180
rect 2251 248404 2285 249180
rect 2347 249180 2495 249181
rect 2347 248404 2381 249180
rect 2381 248404 2461 249180
rect 2461 248404 2495 249180
rect 2557 249180 2705 249181
rect 2557 248404 2591 249180
rect 2591 248404 2671 249180
rect 2671 248404 2705 249180
rect 2767 249180 2915 249181
rect 2767 248404 2801 249180
rect 2801 248404 2881 249180
rect 2881 248404 2915 249180
rect 2977 249180 3125 249181
rect 2977 248404 3011 249180
rect 3011 248404 3091 249180
rect 3091 248404 3125 249180
rect 3187 249180 3335 249181
rect 3187 248404 3221 249180
rect 3221 248404 3301 249180
rect 3301 248404 3335 249180
rect 3397 249180 3545 249181
rect 3397 248404 3431 249180
rect 3431 248404 3511 249180
rect 3511 248404 3545 249180
rect 3607 249180 3755 249181
rect 3607 248404 3641 249180
rect 3641 248404 3721 249180
rect 3721 248404 3755 249180
rect 3817 249180 3965 249181
rect 3817 248404 3851 249180
rect 3851 248404 3931 249180
rect 3931 248404 3965 249180
rect 4027 249180 4175 249181
rect 4027 248404 4061 249180
rect 4061 248404 4141 249180
rect 4141 248404 4175 249180
rect 4237 249180 4385 249181
rect 4237 248404 4271 249180
rect 4271 248404 4351 249180
rect 4351 248404 4385 249180
rect 4447 249180 4595 249181
rect 4447 248404 4481 249180
rect 4481 248404 4561 249180
rect 4561 248404 4595 249180
rect 4657 249180 4805 249181
rect 4657 248404 4691 249180
rect 4691 248404 4771 249180
rect 4771 248404 4805 249180
rect 4867 249180 5015 249181
rect 4867 248404 4901 249180
rect 4901 248404 4981 249180
rect 4981 248404 5015 249180
rect 5077 249180 5225 249181
rect 5077 248404 5111 249180
rect 5111 248404 5191 249180
rect 5191 248404 5225 249180
rect 5287 249180 5435 249181
rect 5287 248404 5321 249180
rect 5321 248404 5401 249180
rect 5401 248404 5435 249180
rect 5497 249180 5645 249181
rect 5497 248404 5531 249180
rect 5531 248404 5611 249180
rect 5611 248404 5645 249180
rect 5707 249180 5855 249181
rect 5707 248404 5741 249180
rect 5741 248404 5821 249180
rect 5821 248404 5855 249180
rect 5917 249180 6065 249181
rect 5917 248404 5951 249180
rect 5951 248404 6031 249180
rect 6031 248404 6065 249180
rect 6127 249180 6275 249181
rect 6127 248404 6161 249180
rect 6161 248404 6241 249180
rect 6241 248404 6275 249180
rect 6337 249180 6485 249181
rect 6337 248404 6371 249180
rect 6371 248404 6451 249180
rect 6451 248404 6485 249180
rect 6547 249180 6695 249181
rect 6547 248404 6581 249180
rect 6581 248404 6661 249180
rect 6661 248404 6695 249180
rect 6757 249180 6905 249181
rect 6757 248404 6791 249180
rect 6791 248404 6871 249180
rect 6871 248404 6905 249180
rect 6967 249180 7115 249181
rect 6967 248404 7001 249180
rect 7001 248404 7081 249180
rect 7081 248404 7115 249180
rect 7177 249180 7325 249181
rect 7177 248404 7211 249180
rect 7211 248404 7291 249180
rect 7291 248404 7325 249180
rect 7387 249180 7535 249181
rect 7387 248404 7421 249180
rect 7421 248404 7501 249180
rect 7501 248404 7535 249180
rect 7597 249180 7745 249181
rect 7597 248404 7631 249180
rect 7631 248404 7711 249180
rect 7711 248404 7745 249180
rect 7807 249180 7955 249181
rect 7807 248404 7841 249180
rect 7841 248404 7921 249180
rect 7921 248404 7955 249180
rect 8017 249180 8165 249181
rect 8017 248404 8051 249180
rect 8051 248404 8131 249180
rect 8131 248404 8165 249180
rect 8227 249180 8375 249181
rect 8227 248404 8261 249180
rect 8261 248404 8341 249180
rect 8341 248404 8375 249180
rect 8437 249180 8585 249181
rect 8437 248404 8471 249180
rect 8471 248404 8551 249180
rect 8551 248404 8585 249180
rect 8647 249180 8795 249181
rect 8647 248404 8681 249180
rect 8681 248404 8761 249180
rect 8761 248404 8795 249180
rect 8857 249180 9005 249181
rect 8857 248404 8891 249180
rect 8891 248404 8971 249180
rect 8971 248404 9005 249180
rect 9067 249180 9215 249181
rect 9067 248404 9101 249180
rect 9101 248404 9181 249180
rect 9181 248404 9215 249180
rect 9277 249180 9425 249181
rect 9277 248404 9311 249180
rect 9311 248404 9391 249180
rect 9391 248404 9425 249180
rect 9487 249180 9635 249181
rect 9487 248404 9521 249180
rect 9521 248404 9601 249180
rect 9601 248404 9635 249180
rect 9697 249180 9845 249181
rect 9697 248404 9731 249180
rect 9731 248404 9811 249180
rect 9811 248404 9845 249180
rect 9907 249180 10055 249181
rect 9907 248404 9941 249180
rect 9941 248404 10021 249180
rect 10021 248404 10055 249180
rect 10117 249180 10265 249181
rect 10117 248404 10151 249180
rect 10151 248404 10231 249180
rect 10231 248404 10265 249180
rect 10327 249180 10475 249181
rect 10327 248404 10361 249180
rect 10361 248404 10441 249180
rect 10441 248404 10475 249180
rect 10537 249180 10685 249181
rect 10537 248404 10571 249180
rect 10571 248404 10651 249180
rect 10651 248404 10685 249180
rect 10747 249180 10895 249181
rect 10747 248404 10781 249180
rect 10781 248404 10861 249180
rect 10861 248404 10895 249180
rect 10957 249180 11105 249181
rect 10957 248404 10991 249180
rect 10991 248404 11071 249180
rect 11071 248404 11105 249180
rect 11167 249180 11315 249181
rect 11167 248404 11201 249180
rect 11201 248404 11281 249180
rect 11281 248404 11315 249180
rect 11377 249180 11525 249181
rect 11377 248404 11411 249180
rect 11411 248404 11491 249180
rect 11491 248404 11525 249180
rect 11587 249180 11735 249181
rect 11587 248404 11621 249180
rect 11621 248404 11701 249180
rect 11701 248404 11735 249180
rect 11797 249180 11945 249181
rect 11797 248404 11831 249180
rect 11831 248404 11911 249180
rect 11911 248404 11945 249180
rect 12007 249180 12155 249181
rect 12007 248404 12041 249180
rect 12041 248404 12121 249180
rect 12121 248404 12155 249180
rect 12217 249180 12365 249181
rect 12217 248404 12251 249180
rect 12251 248404 12331 249180
rect 12331 248404 12365 249180
rect 12427 249180 12575 249181
rect 12427 248404 12461 249180
rect 12461 248404 12541 249180
rect 12541 248404 12575 249180
rect 12637 249180 12785 249181
rect 12637 248404 12671 249180
rect 12671 248404 12751 249180
rect 12751 248404 12785 249180
rect 12847 249180 12995 249181
rect 12847 248404 12881 249180
rect 12881 248404 12961 249180
rect 12961 248404 12995 249180
rect 13057 249180 13205 249181
rect 13057 248404 13091 249180
rect 13091 248404 13171 249180
rect 13171 248404 13205 249180
rect 13267 249180 13415 249181
rect 13267 248404 13301 249180
rect 13301 248404 13381 249180
rect 13381 248404 13415 249180
rect 13477 249180 13625 249181
rect 13477 248404 13511 249180
rect 13511 248404 13591 249180
rect 13591 248404 13625 249180
rect 13687 249180 13835 249181
rect 13687 248404 13721 249180
rect 13721 248404 13801 249180
rect 13801 248404 13835 249180
rect 13897 249180 14045 249181
rect 13897 248404 13931 249180
rect 13931 248404 14011 249180
rect 14011 248404 14045 249180
rect 14107 249180 14255 249181
rect 14107 248404 14141 249180
rect 14141 248404 14221 249180
rect 14221 248404 14255 249180
rect 14317 249180 14465 249181
rect 14317 248404 14351 249180
rect 14351 248404 14431 249180
rect 14431 248404 14465 249180
rect 14527 249180 14675 249181
rect 14527 248404 14561 249180
rect 14561 248404 14641 249180
rect 14641 248404 14675 249180
rect 14737 249180 14885 249181
rect 14737 248404 14771 249180
rect 14771 248404 14851 249180
rect 14851 248404 14885 249180
rect 14947 249180 15095 249181
rect 14947 248404 14981 249180
rect 14981 248404 15061 249180
rect 15061 248404 15095 249180
rect 15157 249180 15305 249181
rect 15157 248404 15191 249180
rect 15191 248404 15271 249180
rect 15271 248404 15305 249180
rect 15367 249180 15515 249181
rect 15367 248404 15401 249180
rect 15401 248404 15481 249180
rect 15481 248404 15515 249180
rect 15577 249180 15725 249181
rect 15577 248404 15611 249180
rect 15611 248404 15691 249180
rect 15691 248404 15725 249180
rect 15787 249180 15935 249181
rect 15787 248404 15821 249180
rect 15821 248404 15901 249180
rect 15901 248404 15935 249180
rect 15997 249180 16145 249181
rect 15997 248404 16031 249180
rect 16031 248404 16111 249180
rect 16111 248404 16145 249180
rect 16207 249180 16355 249181
rect 16207 248404 16241 249180
rect 16241 248404 16321 249180
rect 16321 248404 16355 249180
rect 16417 249180 16565 249181
rect 16417 248404 16451 249180
rect 16451 248404 16531 249180
rect 16531 248404 16565 249180
rect 16627 249180 16775 249181
rect 16627 248404 16661 249180
rect 16661 248404 16741 249180
rect 16741 248404 16775 249180
rect 16837 249180 16985 249181
rect 16837 248404 16871 249180
rect 16871 248404 16951 249180
rect 16951 248404 16985 249180
rect 17047 249180 17195 249181
rect 17047 248404 17081 249180
rect 17081 248404 17161 249180
rect 17161 248404 17195 249180
rect 17257 249180 17405 249181
rect 17257 248404 17291 249180
rect 17291 248404 17371 249180
rect 17371 248404 17405 249180
rect 17467 249180 17615 249181
rect 17467 248404 17501 249180
rect 17501 248404 17581 249180
rect 17581 248404 17615 249180
rect 17677 249180 17825 249181
rect 17677 248404 17711 249180
rect 17711 248404 17791 249180
rect 17791 248404 17825 249180
rect 17887 249180 18035 249181
rect 17887 248404 17921 249180
rect 17921 248404 18001 249180
rect 18001 248404 18035 249180
rect 18097 249180 18245 249181
rect 18097 248404 18131 249180
rect 18131 248404 18211 249180
rect 18211 248404 18245 249180
rect 18307 249180 18455 249181
rect 18307 248404 18341 249180
rect 18341 248404 18421 249180
rect 18421 248404 18455 249180
rect 18517 249180 18665 249181
rect 18517 248404 18551 249180
rect 18551 248404 18631 249180
rect 18631 248404 18665 249180
rect 18727 249180 18875 249181
rect 18727 248404 18761 249180
rect 18761 248404 18841 249180
rect 18841 248404 18875 249180
rect 18937 249180 19085 249181
rect 18937 248404 18971 249180
rect 18971 248404 19051 249180
rect 19051 248404 19085 249180
rect 19147 249180 19295 249181
rect 19147 248404 19181 249180
rect 19181 248404 19261 249180
rect 19261 248404 19295 249180
rect 19357 249180 19505 249181
rect 19357 248404 19391 249180
rect 19391 248404 19471 249180
rect 19471 248404 19505 249180
rect 19567 249180 19715 249181
rect 19567 248404 19601 249180
rect 19601 248404 19681 249180
rect 19681 248404 19715 249180
rect 19777 249180 19925 249181
rect 19777 248404 19811 249180
rect 19811 248404 19891 249180
rect 19891 248404 19925 249180
rect 19987 249180 20135 249181
rect 19987 248404 20021 249180
rect 20021 248404 20101 249180
rect 20101 248404 20135 249180
rect 20197 249180 20345 249181
rect 20197 248404 20231 249180
rect 20231 248404 20311 249180
rect 20311 248404 20345 249180
rect 20407 249180 20555 249181
rect 20407 248404 20441 249180
rect 20441 248404 20521 249180
rect 20521 248404 20555 249180
rect 20617 249180 20765 249181
rect 20617 248404 20651 249180
rect 20651 248404 20731 249180
rect 20731 248404 20765 249180
rect 20827 249180 20975 249181
rect 20827 248404 20861 249180
rect 20861 248404 20941 249180
rect 20941 248404 20975 249180
rect 21037 249180 21185 249181
rect 21037 248404 21071 249180
rect 21071 248404 21151 249180
rect 21151 248404 21185 249180
rect 21247 249180 21395 249181
rect 21247 248404 21281 249180
rect 21281 248404 21361 249180
rect 21361 248404 21395 249180
rect 21457 249180 21605 249181
rect 21457 248404 21491 249180
rect 21491 248404 21571 249180
rect 21571 248404 21605 249180
rect 21667 249180 21815 249181
rect 21667 248404 21701 249180
rect 21701 248404 21781 249180
rect 21781 248404 21815 249180
rect 21877 249180 22025 249181
rect 21877 248404 21911 249180
rect 21911 248404 21991 249180
rect 21991 248404 22025 249180
rect 22087 249180 22235 249181
rect 22087 248404 22121 249180
rect 22121 248404 22201 249180
rect 22201 248404 22235 249180
rect 22297 249180 22445 249181
rect 22297 248404 22331 249180
rect 22331 248404 22411 249180
rect 22411 248404 22445 249180
rect 22507 249180 22655 249181
rect 22507 248404 22541 249180
rect 22541 248404 22621 249180
rect 22621 248404 22655 249180
rect 22717 249180 22865 249181
rect 22717 248404 22751 249180
rect 22751 248404 22831 249180
rect 22831 248404 22865 249180
rect 22927 249180 23075 249181
rect 22927 248404 22961 249180
rect 22961 248404 23041 249180
rect 23041 248404 23075 249180
rect 23137 249180 23285 249181
rect 23137 248404 23171 249180
rect 23171 248404 23251 249180
rect 23251 248404 23285 249180
rect 23347 249180 23495 249181
rect 23347 248404 23381 249180
rect 23381 248404 23461 249180
rect 23461 248404 23495 249180
rect 23557 249180 23705 249181
rect 23557 248404 23591 249180
rect 23591 248404 23671 249180
rect 23671 248404 23705 249180
rect 23767 249180 23915 249181
rect 23767 248404 23801 249180
rect 23801 248404 23881 249180
rect 23881 248404 23915 249180
rect 23977 249180 24125 249181
rect 23977 248404 24011 249180
rect 24011 248404 24091 249180
rect 24091 248404 24125 249180
rect 24187 249180 24335 249181
rect 24187 248404 24221 249180
rect 24221 248404 24301 249180
rect 24301 248404 24335 249180
rect 24397 249180 24545 249181
rect 24397 248404 24431 249180
rect 24431 248404 24511 249180
rect 24511 248404 24545 249180
rect 24607 249180 24755 249181
rect 24607 248404 24641 249180
rect 24641 248404 24721 249180
rect 24721 248404 24755 249180
rect 24817 249180 24965 249181
rect 24817 248404 24851 249180
rect 24851 248404 24931 249180
rect 24931 248404 24965 249180
rect 25027 249180 25175 249181
rect 25027 248404 25061 249180
rect 25061 248404 25141 249180
rect 25141 248404 25175 249180
rect 25237 249180 25385 249181
rect 25237 248404 25271 249180
rect 25271 248404 25351 249180
rect 25351 248404 25385 249180
rect 25447 249180 25595 249181
rect 25447 248404 25481 249180
rect 25481 248404 25561 249180
rect 25561 248404 25595 249180
rect 25657 249180 25805 249181
rect 25657 248404 25691 249180
rect 25691 248404 25771 249180
rect 25771 248404 25805 249180
rect 25867 249180 26015 249181
rect 25867 248404 25901 249180
rect 25901 248404 25981 249180
rect 25981 248404 26015 249180
rect 26077 249180 26225 249181
rect 26077 248404 26111 249180
rect 26111 248404 26191 249180
rect 26191 248404 26225 249180
rect 26287 249180 26435 249181
rect 26287 248404 26321 249180
rect 26321 248404 26401 249180
rect 26401 248404 26435 249180
rect 26497 249180 26645 249181
rect 26497 248404 26531 249180
rect 26531 248404 26611 249180
rect 26611 248404 26645 249180
rect 26707 249180 26855 249181
rect 26707 248404 26741 249180
rect 26741 248404 26821 249180
rect 26821 248404 26855 249180
rect 26917 249180 27065 249181
rect 26917 248404 26951 249180
rect 26951 248404 27031 249180
rect 27031 248404 27065 249180
rect 27127 249180 27275 249181
rect 27127 248404 27161 249180
rect 27161 248404 27241 249180
rect 27241 248404 27275 249180
rect -4075 247368 -4049 248144
rect -4049 247368 -4015 248144
rect -3953 247368 -3919 248144
rect -3919 247368 -3839 248144
rect -3839 247368 -3805 248144
rect -3743 247368 -3709 248144
rect -3709 247368 -3629 248144
rect -3629 247368 -3595 248144
rect -3533 248144 -3385 248145
rect -3533 247368 -3499 248144
rect -3499 247368 -3419 248144
rect -3419 247368 -3385 248144
rect -3323 248144 -3175 248145
rect -3323 247368 -3289 248144
rect -3289 247368 -3209 248144
rect -3209 247368 -3175 248144
rect -3113 248144 -2965 248145
rect -3113 247368 -3079 248144
rect -3079 247368 -2999 248144
rect -2999 247368 -2965 248144
rect -2903 248144 -2755 248145
rect -2903 247368 -2869 248144
rect -2869 247368 -2789 248144
rect -2789 247368 -2755 248144
rect -2693 248144 -2545 248145
rect -2693 247368 -2659 248144
rect -2659 247368 -2579 248144
rect -2579 247368 -2545 248144
rect -2483 248144 -2335 248145
rect -2483 247368 -2449 248144
rect -2449 247368 -2369 248144
rect -2369 247368 -2335 248144
rect -2273 248144 -2125 248145
rect -2273 247368 -2239 248144
rect -2239 247368 -2159 248144
rect -2159 247368 -2125 248144
rect -2063 248144 -1915 248145
rect -2063 247368 -2029 248144
rect -2029 247368 -1949 248144
rect -1949 247368 -1915 248144
rect -1853 248144 -1705 248145
rect -1853 247368 -1819 248144
rect -1819 247368 -1739 248144
rect -1739 247368 -1705 248144
rect -1643 248144 -1495 248145
rect -1643 247368 -1609 248144
rect -1609 247368 -1529 248144
rect -1529 247368 -1495 248144
rect -1433 248144 -1285 248145
rect -1433 247368 -1399 248144
rect -1399 247368 -1319 248144
rect -1319 247368 -1285 248144
rect -1223 248144 -1075 248145
rect -1223 247368 -1189 248144
rect -1189 247368 -1109 248144
rect -1109 247368 -1075 248144
rect -1013 248144 -865 248145
rect -1013 247368 -979 248144
rect -979 247368 -899 248144
rect -899 247368 -865 248144
rect -803 248144 -655 248145
rect -803 247368 -769 248144
rect -769 247368 -689 248144
rect -689 247368 -655 248144
rect -593 248144 -445 248145
rect -593 247368 -559 248144
rect -559 247368 -479 248144
rect -479 247368 -445 248144
rect -383 248144 -235 248145
rect -383 247368 -349 248144
rect -349 247368 -269 248144
rect -269 247368 -235 248144
rect -173 248144 -25 248145
rect -173 247368 -139 248144
rect -139 247368 -59 248144
rect -59 247368 -25 248144
rect 37 248144 185 248145
rect 37 247368 71 248144
rect 71 247368 151 248144
rect 151 247368 185 248144
rect 247 248144 395 248145
rect 247 247368 281 248144
rect 281 247368 361 248144
rect 361 247368 395 248144
rect 457 248144 605 248145
rect 457 247368 491 248144
rect 491 247368 571 248144
rect 571 247368 605 248144
rect 667 248144 815 248145
rect 667 247368 701 248144
rect 701 247368 781 248144
rect 781 247368 815 248144
rect 877 248144 1025 248145
rect 877 247368 911 248144
rect 911 247368 991 248144
rect 991 247368 1025 248144
rect 1087 248144 1235 248145
rect 1087 247368 1121 248144
rect 1121 247368 1201 248144
rect 1201 247368 1235 248144
rect 1297 248144 1445 248145
rect 1297 247368 1331 248144
rect 1331 247368 1411 248144
rect 1411 247368 1445 248144
rect 1507 248144 1655 248145
rect 1507 247368 1541 248144
rect 1541 247368 1621 248144
rect 1621 247368 1655 248144
rect 1717 248144 1865 248145
rect 1717 247368 1751 248144
rect 1751 247368 1831 248144
rect 1831 247368 1865 248144
rect 1927 248144 2075 248145
rect 1927 247368 1961 248144
rect 1961 247368 2041 248144
rect 2041 247368 2075 248144
rect 2137 248144 2285 248145
rect 2137 247368 2171 248144
rect 2171 247368 2251 248144
rect 2251 247368 2285 248144
rect 2347 248144 2495 248145
rect 2347 247368 2381 248144
rect 2381 247368 2461 248144
rect 2461 247368 2495 248144
rect 2557 248144 2705 248145
rect 2557 247368 2591 248144
rect 2591 247368 2671 248144
rect 2671 247368 2705 248144
rect 2767 248144 2915 248145
rect 2767 247368 2801 248144
rect 2801 247368 2881 248144
rect 2881 247368 2915 248144
rect 2977 248144 3125 248145
rect 2977 247368 3011 248144
rect 3011 247368 3091 248144
rect 3091 247368 3125 248144
rect 3187 248144 3335 248145
rect 3187 247368 3221 248144
rect 3221 247368 3301 248144
rect 3301 247368 3335 248144
rect 3397 248144 3545 248145
rect 3397 247368 3431 248144
rect 3431 247368 3511 248144
rect 3511 247368 3545 248144
rect 3607 248144 3755 248145
rect 3607 247368 3641 248144
rect 3641 247368 3721 248144
rect 3721 247368 3755 248144
rect 3817 248144 3965 248145
rect 3817 247368 3851 248144
rect 3851 247368 3931 248144
rect 3931 247368 3965 248144
rect 4027 248144 4175 248145
rect 4027 247368 4061 248144
rect 4061 247368 4141 248144
rect 4141 247368 4175 248144
rect 4237 248144 4385 248145
rect 4237 247368 4271 248144
rect 4271 247368 4351 248144
rect 4351 247368 4385 248144
rect 4447 248144 4595 248145
rect 4447 247368 4481 248144
rect 4481 247368 4561 248144
rect 4561 247368 4595 248144
rect 4657 248144 4805 248145
rect 4657 247368 4691 248144
rect 4691 247368 4771 248144
rect 4771 247368 4805 248144
rect 4867 248144 5015 248145
rect 4867 247368 4901 248144
rect 4901 247368 4981 248144
rect 4981 247368 5015 248144
rect 5077 248144 5225 248145
rect 5077 247368 5111 248144
rect 5111 247368 5191 248144
rect 5191 247368 5225 248144
rect 5287 248144 5435 248145
rect 5287 247368 5321 248144
rect 5321 247368 5401 248144
rect 5401 247368 5435 248144
rect 5497 248144 5645 248145
rect 5497 247368 5531 248144
rect 5531 247368 5611 248144
rect 5611 247368 5645 248144
rect 5707 248144 5855 248145
rect 5707 247368 5741 248144
rect 5741 247368 5821 248144
rect 5821 247368 5855 248144
rect 5917 248144 6065 248145
rect 5917 247368 5951 248144
rect 5951 247368 6031 248144
rect 6031 247368 6065 248144
rect 6127 248144 6275 248145
rect 6127 247368 6161 248144
rect 6161 247368 6241 248144
rect 6241 247368 6275 248144
rect 6337 248144 6485 248145
rect 6337 247368 6371 248144
rect 6371 247368 6451 248144
rect 6451 247368 6485 248144
rect 6547 248144 6695 248145
rect 6547 247368 6581 248144
rect 6581 247368 6661 248144
rect 6661 247368 6695 248144
rect 6757 248144 6905 248145
rect 6757 247368 6791 248144
rect 6791 247368 6871 248144
rect 6871 247368 6905 248144
rect 6967 248144 7115 248145
rect 6967 247368 7001 248144
rect 7001 247368 7081 248144
rect 7081 247368 7115 248144
rect 7177 248144 7325 248145
rect 7177 247368 7211 248144
rect 7211 247368 7291 248144
rect 7291 247368 7325 248144
rect 7387 248144 7535 248145
rect 7387 247368 7421 248144
rect 7421 247368 7501 248144
rect 7501 247368 7535 248144
rect 7597 248144 7745 248145
rect 7597 247368 7631 248144
rect 7631 247368 7711 248144
rect 7711 247368 7745 248144
rect 7807 248144 7955 248145
rect 7807 247368 7841 248144
rect 7841 247368 7921 248144
rect 7921 247368 7955 248144
rect 8017 248144 8165 248145
rect 8017 247368 8051 248144
rect 8051 247368 8131 248144
rect 8131 247368 8165 248144
rect 8227 248144 8375 248145
rect 8227 247368 8261 248144
rect 8261 247368 8341 248144
rect 8341 247368 8375 248144
rect 8437 248144 8585 248145
rect 8437 247368 8471 248144
rect 8471 247368 8551 248144
rect 8551 247368 8585 248144
rect 8647 248144 8795 248145
rect 8647 247368 8681 248144
rect 8681 247368 8761 248144
rect 8761 247368 8795 248144
rect 8857 248144 9005 248145
rect 8857 247368 8891 248144
rect 8891 247368 8971 248144
rect 8971 247368 9005 248144
rect 9067 248144 9215 248145
rect 9067 247368 9101 248144
rect 9101 247368 9181 248144
rect 9181 247368 9215 248144
rect 9277 248144 9425 248145
rect 9277 247368 9311 248144
rect 9311 247368 9391 248144
rect 9391 247368 9425 248144
rect 9487 248144 9635 248145
rect 9487 247368 9521 248144
rect 9521 247368 9601 248144
rect 9601 247368 9635 248144
rect 9697 248144 9845 248145
rect 9697 247368 9731 248144
rect 9731 247368 9811 248144
rect 9811 247368 9845 248144
rect 9907 248144 10055 248145
rect 9907 247368 9941 248144
rect 9941 247368 10021 248144
rect 10021 247368 10055 248144
rect 10117 248144 10265 248145
rect 10117 247368 10151 248144
rect 10151 247368 10231 248144
rect 10231 247368 10265 248144
rect 10327 248144 10475 248145
rect 10327 247368 10361 248144
rect 10361 247368 10441 248144
rect 10441 247368 10475 248144
rect 10537 248144 10685 248145
rect 10537 247368 10571 248144
rect 10571 247368 10651 248144
rect 10651 247368 10685 248144
rect 10747 248144 10895 248145
rect 10747 247368 10781 248144
rect 10781 247368 10861 248144
rect 10861 247368 10895 248144
rect 10957 248144 11105 248145
rect 10957 247368 10991 248144
rect 10991 247368 11071 248144
rect 11071 247368 11105 248144
rect 11167 248144 11315 248145
rect 11167 247368 11201 248144
rect 11201 247368 11281 248144
rect 11281 247368 11315 248144
rect 11377 248144 11525 248145
rect 11377 247368 11411 248144
rect 11411 247368 11491 248144
rect 11491 247368 11525 248144
rect 11587 248144 11735 248145
rect 11587 247368 11621 248144
rect 11621 247368 11701 248144
rect 11701 247368 11735 248144
rect 11797 248144 11945 248145
rect 11797 247368 11831 248144
rect 11831 247368 11911 248144
rect 11911 247368 11945 248144
rect 12007 248144 12155 248145
rect 12007 247368 12041 248144
rect 12041 247368 12121 248144
rect 12121 247368 12155 248144
rect 12217 248144 12365 248145
rect 12217 247368 12251 248144
rect 12251 247368 12331 248144
rect 12331 247368 12365 248144
rect 12427 248144 12575 248145
rect 12427 247368 12461 248144
rect 12461 247368 12541 248144
rect 12541 247368 12575 248144
rect 12637 248144 12785 248145
rect 12637 247368 12671 248144
rect 12671 247368 12751 248144
rect 12751 247368 12785 248144
rect 12847 248144 12995 248145
rect 12847 247368 12881 248144
rect 12881 247368 12961 248144
rect 12961 247368 12995 248144
rect 13057 248144 13205 248145
rect 13057 247368 13091 248144
rect 13091 247368 13171 248144
rect 13171 247368 13205 248144
rect 13267 248144 13415 248145
rect 13267 247368 13301 248144
rect 13301 247368 13381 248144
rect 13381 247368 13415 248144
rect 13477 248144 13625 248145
rect 13477 247368 13511 248144
rect 13511 247368 13591 248144
rect 13591 247368 13625 248144
rect 13687 248144 13835 248145
rect 13687 247368 13721 248144
rect 13721 247368 13801 248144
rect 13801 247368 13835 248144
rect 13897 248144 14045 248145
rect 13897 247368 13931 248144
rect 13931 247368 14011 248144
rect 14011 247368 14045 248144
rect 14107 248144 14255 248145
rect 14107 247368 14141 248144
rect 14141 247368 14221 248144
rect 14221 247368 14255 248144
rect 14317 248144 14465 248145
rect 14317 247368 14351 248144
rect 14351 247368 14431 248144
rect 14431 247368 14465 248144
rect 14527 248144 14675 248145
rect 14527 247368 14561 248144
rect 14561 247368 14641 248144
rect 14641 247368 14675 248144
rect 14737 248144 14885 248145
rect 14737 247368 14771 248144
rect 14771 247368 14851 248144
rect 14851 247368 14885 248144
rect 14947 248144 15095 248145
rect 14947 247368 14981 248144
rect 14981 247368 15061 248144
rect 15061 247368 15095 248144
rect 15157 248144 15305 248145
rect 15157 247368 15191 248144
rect 15191 247368 15271 248144
rect 15271 247368 15305 248144
rect 15367 248144 15515 248145
rect 15367 247368 15401 248144
rect 15401 247368 15481 248144
rect 15481 247368 15515 248144
rect 15577 248144 15725 248145
rect 15577 247368 15611 248144
rect 15611 247368 15691 248144
rect 15691 247368 15725 248144
rect 15787 248144 15935 248145
rect 15787 247368 15821 248144
rect 15821 247368 15901 248144
rect 15901 247368 15935 248144
rect 15997 248144 16145 248145
rect 15997 247368 16031 248144
rect 16031 247368 16111 248144
rect 16111 247368 16145 248144
rect 16207 248144 16355 248145
rect 16207 247368 16241 248144
rect 16241 247368 16321 248144
rect 16321 247368 16355 248144
rect 16417 248144 16565 248145
rect 16417 247368 16451 248144
rect 16451 247368 16531 248144
rect 16531 247368 16565 248144
rect 16627 248144 16775 248145
rect 16627 247368 16661 248144
rect 16661 247368 16741 248144
rect 16741 247368 16775 248144
rect 16837 248144 16985 248145
rect 16837 247368 16871 248144
rect 16871 247368 16951 248144
rect 16951 247368 16985 248144
rect 17047 248144 17195 248145
rect 17047 247368 17081 248144
rect 17081 247368 17161 248144
rect 17161 247368 17195 248144
rect 17257 248144 17405 248145
rect 17257 247368 17291 248144
rect 17291 247368 17371 248144
rect 17371 247368 17405 248144
rect 17467 248144 17615 248145
rect 17467 247368 17501 248144
rect 17501 247368 17581 248144
rect 17581 247368 17615 248144
rect 17677 248144 17825 248145
rect 17677 247368 17711 248144
rect 17711 247368 17791 248144
rect 17791 247368 17825 248144
rect 17887 248144 18035 248145
rect 17887 247368 17921 248144
rect 17921 247368 18001 248144
rect 18001 247368 18035 248144
rect 18097 248144 18245 248145
rect 18097 247368 18131 248144
rect 18131 247368 18211 248144
rect 18211 247368 18245 248144
rect 18307 248144 18455 248145
rect 18307 247368 18341 248144
rect 18341 247368 18421 248144
rect 18421 247368 18455 248144
rect 18517 248144 18665 248145
rect 18517 247368 18551 248144
rect 18551 247368 18631 248144
rect 18631 247368 18665 248144
rect 18727 248144 18875 248145
rect 18727 247368 18761 248144
rect 18761 247368 18841 248144
rect 18841 247368 18875 248144
rect 18937 248144 19085 248145
rect 18937 247368 18971 248144
rect 18971 247368 19051 248144
rect 19051 247368 19085 248144
rect 19147 248144 19295 248145
rect 19147 247368 19181 248144
rect 19181 247368 19261 248144
rect 19261 247368 19295 248144
rect 19357 248144 19505 248145
rect 19357 247368 19391 248144
rect 19391 247368 19471 248144
rect 19471 247368 19505 248144
rect 19567 248144 19715 248145
rect 19567 247368 19601 248144
rect 19601 247368 19681 248144
rect 19681 247368 19715 248144
rect 19777 248144 19925 248145
rect 19777 247368 19811 248144
rect 19811 247368 19891 248144
rect 19891 247368 19925 248144
rect 19987 248144 20135 248145
rect 19987 247368 20021 248144
rect 20021 247368 20101 248144
rect 20101 247368 20135 248144
rect 20197 248144 20345 248145
rect 20197 247368 20231 248144
rect 20231 247368 20311 248144
rect 20311 247368 20345 248144
rect 20407 248144 20555 248145
rect 20407 247368 20441 248144
rect 20441 247368 20521 248144
rect 20521 247368 20555 248144
rect 20617 248144 20765 248145
rect 20617 247368 20651 248144
rect 20651 247368 20731 248144
rect 20731 247368 20765 248144
rect 20827 248144 20975 248145
rect 20827 247368 20861 248144
rect 20861 247368 20941 248144
rect 20941 247368 20975 248144
rect 21037 248144 21185 248145
rect 21037 247368 21071 248144
rect 21071 247368 21151 248144
rect 21151 247368 21185 248144
rect 21247 248144 21395 248145
rect 21247 247368 21281 248144
rect 21281 247368 21361 248144
rect 21361 247368 21395 248144
rect 21457 248144 21605 248145
rect 21457 247368 21491 248144
rect 21491 247368 21571 248144
rect 21571 247368 21605 248144
rect 21667 248144 21815 248145
rect 21667 247368 21701 248144
rect 21701 247368 21781 248144
rect 21781 247368 21815 248144
rect 21877 248144 22025 248145
rect 21877 247368 21911 248144
rect 21911 247368 21991 248144
rect 21991 247368 22025 248144
rect 22087 248144 22235 248145
rect 22087 247368 22121 248144
rect 22121 247368 22201 248144
rect 22201 247368 22235 248144
rect 22297 248144 22445 248145
rect 22297 247368 22331 248144
rect 22331 247368 22411 248144
rect 22411 247368 22445 248144
rect 22507 248144 22655 248145
rect 22507 247368 22541 248144
rect 22541 247368 22621 248144
rect 22621 247368 22655 248144
rect 22717 248144 22865 248145
rect 22717 247368 22751 248144
rect 22751 247368 22831 248144
rect 22831 247368 22865 248144
rect 22927 248144 23075 248145
rect 22927 247368 22961 248144
rect 22961 247368 23041 248144
rect 23041 247368 23075 248144
rect 23137 248144 23285 248145
rect 23137 247368 23171 248144
rect 23171 247368 23251 248144
rect 23251 247368 23285 248144
rect 23347 248144 23495 248145
rect 23347 247368 23381 248144
rect 23381 247368 23461 248144
rect 23461 247368 23495 248144
rect 23557 248144 23705 248145
rect 23557 247368 23591 248144
rect 23591 247368 23671 248144
rect 23671 247368 23705 248144
rect 23767 248144 23915 248145
rect 23767 247368 23801 248144
rect 23801 247368 23881 248144
rect 23881 247368 23915 248144
rect 23977 248144 24125 248145
rect 23977 247368 24011 248144
rect 24011 247368 24091 248144
rect 24091 247368 24125 248144
rect 24187 248144 24335 248145
rect 24187 247368 24221 248144
rect 24221 247368 24301 248144
rect 24301 247368 24335 248144
rect 24397 248144 24545 248145
rect 24397 247368 24431 248144
rect 24431 247368 24511 248144
rect 24511 247368 24545 248144
rect 24607 248144 24755 248145
rect 24607 247368 24641 248144
rect 24641 247368 24721 248144
rect 24721 247368 24755 248144
rect 24817 248144 24965 248145
rect 24817 247368 24851 248144
rect 24851 247368 24931 248144
rect 24931 247368 24965 248144
rect 25027 248144 25175 248145
rect 25027 247368 25061 248144
rect 25061 247368 25141 248144
rect 25141 247368 25175 248144
rect 25237 248144 25385 248145
rect 25237 247368 25271 248144
rect 25271 247368 25351 248144
rect 25351 247368 25385 248144
rect 25447 248144 25595 248145
rect 25447 247368 25481 248144
rect 25481 247368 25561 248144
rect 25561 247368 25595 248144
rect 25657 248144 25805 248145
rect 25657 247368 25691 248144
rect 25691 247368 25771 248144
rect 25771 247368 25805 248144
rect 25867 248144 26015 248145
rect 25867 247368 25901 248144
rect 25901 247368 25981 248144
rect 25981 247368 26015 248144
rect 26077 248144 26225 248145
rect 26077 247368 26111 248144
rect 26111 247368 26191 248144
rect 26191 247368 26225 248144
rect 26287 248144 26435 248145
rect 26287 247368 26321 248144
rect 26321 247368 26401 248144
rect 26401 247368 26435 248144
rect 26497 248144 26645 248145
rect 26497 247368 26531 248144
rect 26531 247368 26611 248144
rect 26611 247368 26645 248144
rect 26707 248144 26855 248145
rect 26707 247368 26741 248144
rect 26741 247368 26821 248144
rect 26821 247368 26855 248144
rect 26917 248144 27065 248145
rect 26917 247368 26951 248144
rect 26951 247368 27031 248144
rect 27031 247368 27065 248144
rect 27127 248144 27275 248145
rect 27127 247368 27161 248144
rect 27161 247368 27241 248144
rect 27241 247368 27275 248144
rect -4075 246332 -4049 247108
rect -4049 246332 -4015 247108
rect -3953 246332 -3919 247108
rect -3919 246332 -3839 247108
rect -3839 246332 -3805 247108
rect -3743 246332 -3709 247108
rect -3709 246332 -3629 247108
rect -3629 246332 -3595 247108
rect -3533 247108 -3385 247109
rect -3533 246332 -3499 247108
rect -3499 246332 -3419 247108
rect -3419 246332 -3385 247108
rect -3323 247108 -3175 247109
rect -3323 246332 -3289 247108
rect -3289 246332 -3209 247108
rect -3209 246332 -3175 247108
rect -3113 247108 -2965 247109
rect -3113 246332 -3079 247108
rect -3079 246332 -2999 247108
rect -2999 246332 -2965 247108
rect -2903 247108 -2755 247109
rect -2903 246332 -2869 247108
rect -2869 246332 -2789 247108
rect -2789 246332 -2755 247108
rect -2693 247108 -2545 247109
rect -2693 246332 -2659 247108
rect -2659 246332 -2579 247108
rect -2579 246332 -2545 247108
rect -2483 247108 -2335 247109
rect -2483 246332 -2449 247108
rect -2449 246332 -2369 247108
rect -2369 246332 -2335 247108
rect -2273 247108 -2125 247109
rect -2273 246332 -2239 247108
rect -2239 246332 -2159 247108
rect -2159 246332 -2125 247108
rect -2063 247108 -1915 247109
rect -2063 246332 -2029 247108
rect -2029 246332 -1949 247108
rect -1949 246332 -1915 247108
rect -1853 247108 -1705 247109
rect -1853 246332 -1819 247108
rect -1819 246332 -1739 247108
rect -1739 246332 -1705 247108
rect -1643 247108 -1495 247109
rect -1643 246332 -1609 247108
rect -1609 246332 -1529 247108
rect -1529 246332 -1495 247108
rect -1433 247108 -1285 247109
rect -1433 246332 -1399 247108
rect -1399 246332 -1319 247108
rect -1319 246332 -1285 247108
rect -1223 247108 -1075 247109
rect -1223 246332 -1189 247108
rect -1189 246332 -1109 247108
rect -1109 246332 -1075 247108
rect -1013 247108 -865 247109
rect -1013 246332 -979 247108
rect -979 246332 -899 247108
rect -899 246332 -865 247108
rect -803 247108 -655 247109
rect -803 246332 -769 247108
rect -769 246332 -689 247108
rect -689 246332 -655 247108
rect -593 247108 -445 247109
rect -593 246332 -559 247108
rect -559 246332 -479 247108
rect -479 246332 -445 247108
rect -383 247108 -235 247109
rect -383 246332 -349 247108
rect -349 246332 -269 247108
rect -269 246332 -235 247108
rect -173 247108 -25 247109
rect -173 246332 -139 247108
rect -139 246332 -59 247108
rect -59 246332 -25 247108
rect 37 247108 185 247109
rect 37 246332 71 247108
rect 71 246332 151 247108
rect 151 246332 185 247108
rect 247 247108 395 247109
rect 247 246332 281 247108
rect 281 246332 361 247108
rect 361 246332 395 247108
rect 457 247108 605 247109
rect 457 246332 491 247108
rect 491 246332 571 247108
rect 571 246332 605 247108
rect 667 247108 815 247109
rect 667 246332 701 247108
rect 701 246332 781 247108
rect 781 246332 815 247108
rect 877 247108 1025 247109
rect 877 246332 911 247108
rect 911 246332 991 247108
rect 991 246332 1025 247108
rect 1087 247108 1235 247109
rect 1087 246332 1121 247108
rect 1121 246332 1201 247108
rect 1201 246332 1235 247108
rect 1297 247108 1445 247109
rect 1297 246332 1331 247108
rect 1331 246332 1411 247108
rect 1411 246332 1445 247108
rect 1507 247108 1655 247109
rect 1507 246332 1541 247108
rect 1541 246332 1621 247108
rect 1621 246332 1655 247108
rect 1717 247108 1865 247109
rect 1717 246332 1751 247108
rect 1751 246332 1831 247108
rect 1831 246332 1865 247108
rect 1927 247108 2075 247109
rect 1927 246332 1961 247108
rect 1961 246332 2041 247108
rect 2041 246332 2075 247108
rect 2137 247108 2285 247109
rect 2137 246332 2171 247108
rect 2171 246332 2251 247108
rect 2251 246332 2285 247108
rect 2347 247108 2495 247109
rect 2347 246332 2381 247108
rect 2381 246332 2461 247108
rect 2461 246332 2495 247108
rect 2557 247108 2705 247109
rect 2557 246332 2591 247108
rect 2591 246332 2671 247108
rect 2671 246332 2705 247108
rect 2767 247108 2915 247109
rect 2767 246332 2801 247108
rect 2801 246332 2881 247108
rect 2881 246332 2915 247108
rect 2977 247108 3125 247109
rect 2977 246332 3011 247108
rect 3011 246332 3091 247108
rect 3091 246332 3125 247108
rect 3187 247108 3335 247109
rect 3187 246332 3221 247108
rect 3221 246332 3301 247108
rect 3301 246332 3335 247108
rect 3397 247108 3545 247109
rect 3397 246332 3431 247108
rect 3431 246332 3511 247108
rect 3511 246332 3545 247108
rect 3607 247108 3755 247109
rect 3607 246332 3641 247108
rect 3641 246332 3721 247108
rect 3721 246332 3755 247108
rect 3817 247108 3965 247109
rect 3817 246332 3851 247108
rect 3851 246332 3931 247108
rect 3931 246332 3965 247108
rect 4027 247108 4175 247109
rect 4027 246332 4061 247108
rect 4061 246332 4141 247108
rect 4141 246332 4175 247108
rect 4237 247108 4385 247109
rect 4237 246332 4271 247108
rect 4271 246332 4351 247108
rect 4351 246332 4385 247108
rect 4447 247108 4595 247109
rect 4447 246332 4481 247108
rect 4481 246332 4561 247108
rect 4561 246332 4595 247108
rect 4657 247108 4805 247109
rect 4657 246332 4691 247108
rect 4691 246332 4771 247108
rect 4771 246332 4805 247108
rect 4867 247108 5015 247109
rect 4867 246332 4901 247108
rect 4901 246332 4981 247108
rect 4981 246332 5015 247108
rect 5077 247108 5225 247109
rect 5077 246332 5111 247108
rect 5111 246332 5191 247108
rect 5191 246332 5225 247108
rect 5287 247108 5435 247109
rect 5287 246332 5321 247108
rect 5321 246332 5401 247108
rect 5401 246332 5435 247108
rect 5497 247108 5645 247109
rect 5497 246332 5531 247108
rect 5531 246332 5611 247108
rect 5611 246332 5645 247108
rect 5707 247108 5855 247109
rect 5707 246332 5741 247108
rect 5741 246332 5821 247108
rect 5821 246332 5855 247108
rect 5917 247108 6065 247109
rect 5917 246332 5951 247108
rect 5951 246332 6031 247108
rect 6031 246332 6065 247108
rect 6127 247108 6275 247109
rect 6127 246332 6161 247108
rect 6161 246332 6241 247108
rect 6241 246332 6275 247108
rect 6337 247108 6485 247109
rect 6337 246332 6371 247108
rect 6371 246332 6451 247108
rect 6451 246332 6485 247108
rect 6547 247108 6695 247109
rect 6547 246332 6581 247108
rect 6581 246332 6661 247108
rect 6661 246332 6695 247108
rect 6757 247108 6905 247109
rect 6757 246332 6791 247108
rect 6791 246332 6871 247108
rect 6871 246332 6905 247108
rect 6967 247108 7115 247109
rect 6967 246332 7001 247108
rect 7001 246332 7081 247108
rect 7081 246332 7115 247108
rect 7177 247108 7325 247109
rect 7177 246332 7211 247108
rect 7211 246332 7291 247108
rect 7291 246332 7325 247108
rect 7387 247108 7535 247109
rect 7387 246332 7421 247108
rect 7421 246332 7501 247108
rect 7501 246332 7535 247108
rect 7597 247108 7745 247109
rect 7597 246332 7631 247108
rect 7631 246332 7711 247108
rect 7711 246332 7745 247108
rect 7807 247108 7955 247109
rect 7807 246332 7841 247108
rect 7841 246332 7921 247108
rect 7921 246332 7955 247108
rect 8017 247108 8165 247109
rect 8017 246332 8051 247108
rect 8051 246332 8131 247108
rect 8131 246332 8165 247108
rect 8227 247108 8375 247109
rect 8227 246332 8261 247108
rect 8261 246332 8341 247108
rect 8341 246332 8375 247108
rect 8437 247108 8585 247109
rect 8437 246332 8471 247108
rect 8471 246332 8551 247108
rect 8551 246332 8585 247108
rect 8647 247108 8795 247109
rect 8647 246332 8681 247108
rect 8681 246332 8761 247108
rect 8761 246332 8795 247108
rect 8857 247108 9005 247109
rect 8857 246332 8891 247108
rect 8891 246332 8971 247108
rect 8971 246332 9005 247108
rect 9067 247108 9215 247109
rect 9067 246332 9101 247108
rect 9101 246332 9181 247108
rect 9181 246332 9215 247108
rect 9277 247108 9425 247109
rect 9277 246332 9311 247108
rect 9311 246332 9391 247108
rect 9391 246332 9425 247108
rect 9487 247108 9635 247109
rect 9487 246332 9521 247108
rect 9521 246332 9601 247108
rect 9601 246332 9635 247108
rect 9697 247108 9845 247109
rect 9697 246332 9731 247108
rect 9731 246332 9811 247108
rect 9811 246332 9845 247108
rect 9907 247108 10055 247109
rect 9907 246332 9941 247108
rect 9941 246332 10021 247108
rect 10021 246332 10055 247108
rect 10117 247108 10265 247109
rect 10117 246332 10151 247108
rect 10151 246332 10231 247108
rect 10231 246332 10265 247108
rect 10327 247108 10475 247109
rect 10327 246332 10361 247108
rect 10361 246332 10441 247108
rect 10441 246332 10475 247108
rect 10537 247108 10685 247109
rect 10537 246332 10571 247108
rect 10571 246332 10651 247108
rect 10651 246332 10685 247108
rect 10747 247108 10895 247109
rect 10747 246332 10781 247108
rect 10781 246332 10861 247108
rect 10861 246332 10895 247108
rect 10957 247108 11105 247109
rect 10957 246332 10991 247108
rect 10991 246332 11071 247108
rect 11071 246332 11105 247108
rect 11167 247108 11315 247109
rect 11167 246332 11201 247108
rect 11201 246332 11281 247108
rect 11281 246332 11315 247108
rect 11377 247108 11525 247109
rect 11377 246332 11411 247108
rect 11411 246332 11491 247108
rect 11491 246332 11525 247108
rect 11587 247108 11735 247109
rect 11587 246332 11621 247108
rect 11621 246332 11701 247108
rect 11701 246332 11735 247108
rect 11797 247108 11945 247109
rect 11797 246332 11831 247108
rect 11831 246332 11911 247108
rect 11911 246332 11945 247108
rect 12007 247108 12155 247109
rect 12007 246332 12041 247108
rect 12041 246332 12121 247108
rect 12121 246332 12155 247108
rect 12217 247108 12365 247109
rect 12217 246332 12251 247108
rect 12251 246332 12331 247108
rect 12331 246332 12365 247108
rect 12427 247108 12575 247109
rect 12427 246332 12461 247108
rect 12461 246332 12541 247108
rect 12541 246332 12575 247108
rect 12637 247108 12785 247109
rect 12637 246332 12671 247108
rect 12671 246332 12751 247108
rect 12751 246332 12785 247108
rect 12847 247108 12995 247109
rect 12847 246332 12881 247108
rect 12881 246332 12961 247108
rect 12961 246332 12995 247108
rect 13057 247108 13205 247109
rect 13057 246332 13091 247108
rect 13091 246332 13171 247108
rect 13171 246332 13205 247108
rect 13267 247108 13415 247109
rect 13267 246332 13301 247108
rect 13301 246332 13381 247108
rect 13381 246332 13415 247108
rect 13477 247108 13625 247109
rect 13477 246332 13511 247108
rect 13511 246332 13591 247108
rect 13591 246332 13625 247108
rect 13687 247108 13835 247109
rect 13687 246332 13721 247108
rect 13721 246332 13801 247108
rect 13801 246332 13835 247108
rect 13897 247108 14045 247109
rect 13897 246332 13931 247108
rect 13931 246332 14011 247108
rect 14011 246332 14045 247108
rect 14107 247108 14255 247109
rect 14107 246332 14141 247108
rect 14141 246332 14221 247108
rect 14221 246332 14255 247108
rect 14317 247108 14465 247109
rect 14317 246332 14351 247108
rect 14351 246332 14431 247108
rect 14431 246332 14465 247108
rect 14527 247108 14675 247109
rect 14527 246332 14561 247108
rect 14561 246332 14641 247108
rect 14641 246332 14675 247108
rect 14737 247108 14885 247109
rect 14737 246332 14771 247108
rect 14771 246332 14851 247108
rect 14851 246332 14885 247108
rect 14947 247108 15095 247109
rect 14947 246332 14981 247108
rect 14981 246332 15061 247108
rect 15061 246332 15095 247108
rect 15157 247108 15305 247109
rect 15157 246332 15191 247108
rect 15191 246332 15271 247108
rect 15271 246332 15305 247108
rect 15367 247108 15515 247109
rect 15367 246332 15401 247108
rect 15401 246332 15481 247108
rect 15481 246332 15515 247108
rect 15577 247108 15725 247109
rect 15577 246332 15611 247108
rect 15611 246332 15691 247108
rect 15691 246332 15725 247108
rect 15787 247108 15935 247109
rect 15787 246332 15821 247108
rect 15821 246332 15901 247108
rect 15901 246332 15935 247108
rect 15997 247108 16145 247109
rect 15997 246332 16031 247108
rect 16031 246332 16111 247108
rect 16111 246332 16145 247108
rect 16207 247108 16355 247109
rect 16207 246332 16241 247108
rect 16241 246332 16321 247108
rect 16321 246332 16355 247108
rect 16417 247108 16565 247109
rect 16417 246332 16451 247108
rect 16451 246332 16531 247108
rect 16531 246332 16565 247108
rect 16627 247108 16775 247109
rect 16627 246332 16661 247108
rect 16661 246332 16741 247108
rect 16741 246332 16775 247108
rect 16837 247108 16985 247109
rect 16837 246332 16871 247108
rect 16871 246332 16951 247108
rect 16951 246332 16985 247108
rect 17047 247108 17195 247109
rect 17047 246332 17081 247108
rect 17081 246332 17161 247108
rect 17161 246332 17195 247108
rect 17257 247108 17405 247109
rect 17257 246332 17291 247108
rect 17291 246332 17371 247108
rect 17371 246332 17405 247108
rect 17467 247108 17615 247109
rect 17467 246332 17501 247108
rect 17501 246332 17581 247108
rect 17581 246332 17615 247108
rect 17677 247108 17825 247109
rect 17677 246332 17711 247108
rect 17711 246332 17791 247108
rect 17791 246332 17825 247108
rect 17887 247108 18035 247109
rect 17887 246332 17921 247108
rect 17921 246332 18001 247108
rect 18001 246332 18035 247108
rect 18097 247108 18245 247109
rect 18097 246332 18131 247108
rect 18131 246332 18211 247108
rect 18211 246332 18245 247108
rect 18307 247108 18455 247109
rect 18307 246332 18341 247108
rect 18341 246332 18421 247108
rect 18421 246332 18455 247108
rect 18517 247108 18665 247109
rect 18517 246332 18551 247108
rect 18551 246332 18631 247108
rect 18631 246332 18665 247108
rect 18727 247108 18875 247109
rect 18727 246332 18761 247108
rect 18761 246332 18841 247108
rect 18841 246332 18875 247108
rect 18937 247108 19085 247109
rect 18937 246332 18971 247108
rect 18971 246332 19051 247108
rect 19051 246332 19085 247108
rect 19147 247108 19295 247109
rect 19147 246332 19181 247108
rect 19181 246332 19261 247108
rect 19261 246332 19295 247108
rect 19357 247108 19505 247109
rect 19357 246332 19391 247108
rect 19391 246332 19471 247108
rect 19471 246332 19505 247108
rect 19567 247108 19715 247109
rect 19567 246332 19601 247108
rect 19601 246332 19681 247108
rect 19681 246332 19715 247108
rect 19777 247108 19925 247109
rect 19777 246332 19811 247108
rect 19811 246332 19891 247108
rect 19891 246332 19925 247108
rect 19987 247108 20135 247109
rect 19987 246332 20021 247108
rect 20021 246332 20101 247108
rect 20101 246332 20135 247108
rect 20197 247108 20345 247109
rect 20197 246332 20231 247108
rect 20231 246332 20311 247108
rect 20311 246332 20345 247108
rect 20407 247108 20555 247109
rect 20407 246332 20441 247108
rect 20441 246332 20521 247108
rect 20521 246332 20555 247108
rect 20617 247108 20765 247109
rect 20617 246332 20651 247108
rect 20651 246332 20731 247108
rect 20731 246332 20765 247108
rect 20827 247108 20975 247109
rect 20827 246332 20861 247108
rect 20861 246332 20941 247108
rect 20941 246332 20975 247108
rect 21037 247108 21185 247109
rect 21037 246332 21071 247108
rect 21071 246332 21151 247108
rect 21151 246332 21185 247108
rect 21247 247108 21395 247109
rect 21247 246332 21281 247108
rect 21281 246332 21361 247108
rect 21361 246332 21395 247108
rect 21457 247108 21605 247109
rect 21457 246332 21491 247108
rect 21491 246332 21571 247108
rect 21571 246332 21605 247108
rect 21667 247108 21815 247109
rect 21667 246332 21701 247108
rect 21701 246332 21781 247108
rect 21781 246332 21815 247108
rect 21877 247108 22025 247109
rect 21877 246332 21911 247108
rect 21911 246332 21991 247108
rect 21991 246332 22025 247108
rect 22087 247108 22235 247109
rect 22087 246332 22121 247108
rect 22121 246332 22201 247108
rect 22201 246332 22235 247108
rect 22297 247108 22445 247109
rect 22297 246332 22331 247108
rect 22331 246332 22411 247108
rect 22411 246332 22445 247108
rect 22507 247108 22655 247109
rect 22507 246332 22541 247108
rect 22541 246332 22621 247108
rect 22621 246332 22655 247108
rect 22717 247108 22865 247109
rect 22717 246332 22751 247108
rect 22751 246332 22831 247108
rect 22831 246332 22865 247108
rect 22927 247108 23075 247109
rect 22927 246332 22961 247108
rect 22961 246332 23041 247108
rect 23041 246332 23075 247108
rect 23137 247108 23285 247109
rect 23137 246332 23171 247108
rect 23171 246332 23251 247108
rect 23251 246332 23285 247108
rect 23347 247108 23495 247109
rect 23347 246332 23381 247108
rect 23381 246332 23461 247108
rect 23461 246332 23495 247108
rect 23557 247108 23705 247109
rect 23557 246332 23591 247108
rect 23591 246332 23671 247108
rect 23671 246332 23705 247108
rect 23767 247108 23915 247109
rect 23767 246332 23801 247108
rect 23801 246332 23881 247108
rect 23881 246332 23915 247108
rect 23977 247108 24125 247109
rect 23977 246332 24011 247108
rect 24011 246332 24091 247108
rect 24091 246332 24125 247108
rect 24187 247108 24335 247109
rect 24187 246332 24221 247108
rect 24221 246332 24301 247108
rect 24301 246332 24335 247108
rect 24397 247108 24545 247109
rect 24397 246332 24431 247108
rect 24431 246332 24511 247108
rect 24511 246332 24545 247108
rect 24607 247108 24755 247109
rect 24607 246332 24641 247108
rect 24641 246332 24721 247108
rect 24721 246332 24755 247108
rect 24817 247108 24965 247109
rect 24817 246332 24851 247108
rect 24851 246332 24931 247108
rect 24931 246332 24965 247108
rect 25027 247108 25175 247109
rect 25027 246332 25061 247108
rect 25061 246332 25141 247108
rect 25141 246332 25175 247108
rect 25237 247108 25385 247109
rect 25237 246332 25271 247108
rect 25271 246332 25351 247108
rect 25351 246332 25385 247108
rect 25447 247108 25595 247109
rect 25447 246332 25481 247108
rect 25481 246332 25561 247108
rect 25561 246332 25595 247108
rect 25657 247108 25805 247109
rect 25657 246332 25691 247108
rect 25691 246332 25771 247108
rect 25771 246332 25805 247108
rect 25867 247108 26015 247109
rect 25867 246332 25901 247108
rect 25901 246332 25981 247108
rect 25981 246332 26015 247108
rect 26077 247108 26225 247109
rect 26077 246332 26111 247108
rect 26111 246332 26191 247108
rect 26191 246332 26225 247108
rect 26287 247108 26435 247109
rect 26287 246332 26321 247108
rect 26321 246332 26401 247108
rect 26401 246332 26435 247108
rect 26497 247108 26645 247109
rect 26497 246332 26531 247108
rect 26531 246332 26611 247108
rect 26611 246332 26645 247108
rect 26707 247108 26855 247109
rect 26707 246332 26741 247108
rect 26741 246332 26821 247108
rect 26821 246332 26855 247108
rect 26917 247108 27065 247109
rect 26917 246332 26951 247108
rect 26951 246332 27031 247108
rect 27031 246332 27065 247108
rect 27127 247108 27275 247109
rect 27127 246332 27161 247108
rect 27161 246332 27241 247108
rect 27241 246332 27275 247108
rect -4075 245296 -4049 246072
rect -4049 245296 -4015 246072
rect -3953 245296 -3919 246072
rect -3919 245296 -3839 246072
rect -3839 245296 -3805 246072
rect -3743 245296 -3709 246072
rect -3709 245296 -3629 246072
rect -3629 245296 -3595 246072
rect -3533 246072 -3385 246073
rect -3533 245296 -3499 246072
rect -3499 245296 -3419 246072
rect -3419 245296 -3385 246072
rect -3323 246072 -3175 246073
rect -3323 245296 -3289 246072
rect -3289 245296 -3209 246072
rect -3209 245296 -3175 246072
rect -3113 246072 -2965 246073
rect -3113 245296 -3079 246072
rect -3079 245296 -2999 246072
rect -2999 245296 -2965 246072
rect -2903 246072 -2755 246073
rect -2903 245296 -2869 246072
rect -2869 245296 -2789 246072
rect -2789 245296 -2755 246072
rect -2693 246072 -2545 246073
rect -2693 245296 -2659 246072
rect -2659 245296 -2579 246072
rect -2579 245296 -2545 246072
rect -2483 246072 -2335 246073
rect -2483 245296 -2449 246072
rect -2449 245296 -2369 246072
rect -2369 245296 -2335 246072
rect -2273 246072 -2125 246073
rect -2273 245296 -2239 246072
rect -2239 245296 -2159 246072
rect -2159 245296 -2125 246072
rect -2063 246072 -1915 246073
rect -2063 245296 -2029 246072
rect -2029 245296 -1949 246072
rect -1949 245296 -1915 246072
rect -1853 246072 -1705 246073
rect -1853 245296 -1819 246072
rect -1819 245296 -1739 246072
rect -1739 245296 -1705 246072
rect -1643 246072 -1495 246073
rect -1643 245296 -1609 246072
rect -1609 245296 -1529 246072
rect -1529 245296 -1495 246072
rect -1433 246072 -1285 246073
rect -1433 245296 -1399 246072
rect -1399 245296 -1319 246072
rect -1319 245296 -1285 246072
rect -1223 246072 -1075 246073
rect -1223 245296 -1189 246072
rect -1189 245296 -1109 246072
rect -1109 245296 -1075 246072
rect -1013 246072 -865 246073
rect -1013 245296 -979 246072
rect -979 245296 -899 246072
rect -899 245296 -865 246072
rect -803 246072 -655 246073
rect -803 245296 -769 246072
rect -769 245296 -689 246072
rect -689 245296 -655 246072
rect -593 246072 -445 246073
rect -593 245296 -559 246072
rect -559 245296 -479 246072
rect -479 245296 -445 246072
rect -383 246072 -235 246073
rect -383 245296 -349 246072
rect -349 245296 -269 246072
rect -269 245296 -235 246072
rect -173 246072 -25 246073
rect -173 245296 -139 246072
rect -139 245296 -59 246072
rect -59 245296 -25 246072
rect 37 246072 185 246073
rect 37 245296 71 246072
rect 71 245296 151 246072
rect 151 245296 185 246072
rect 247 246072 395 246073
rect 247 245296 281 246072
rect 281 245296 361 246072
rect 361 245296 395 246072
rect 457 246072 605 246073
rect 457 245296 491 246072
rect 491 245296 571 246072
rect 571 245296 605 246072
rect 667 246072 815 246073
rect 667 245296 701 246072
rect 701 245296 781 246072
rect 781 245296 815 246072
rect 877 246072 1025 246073
rect 877 245296 911 246072
rect 911 245296 991 246072
rect 991 245296 1025 246072
rect 1087 246072 1235 246073
rect 1087 245296 1121 246072
rect 1121 245296 1201 246072
rect 1201 245296 1235 246072
rect 1297 246072 1445 246073
rect 1297 245296 1331 246072
rect 1331 245296 1411 246072
rect 1411 245296 1445 246072
rect 1507 246072 1655 246073
rect 1507 245296 1541 246072
rect 1541 245296 1621 246072
rect 1621 245296 1655 246072
rect 1717 246072 1865 246073
rect 1717 245296 1751 246072
rect 1751 245296 1831 246072
rect 1831 245296 1865 246072
rect 1927 246072 2075 246073
rect 1927 245296 1961 246072
rect 1961 245296 2041 246072
rect 2041 245296 2075 246072
rect 2137 246072 2285 246073
rect 2137 245296 2171 246072
rect 2171 245296 2251 246072
rect 2251 245296 2285 246072
rect 2347 246072 2495 246073
rect 2347 245296 2381 246072
rect 2381 245296 2461 246072
rect 2461 245296 2495 246072
rect 2557 246072 2705 246073
rect 2557 245296 2591 246072
rect 2591 245296 2671 246072
rect 2671 245296 2705 246072
rect 2767 246072 2915 246073
rect 2767 245296 2801 246072
rect 2801 245296 2881 246072
rect 2881 245296 2915 246072
rect 2977 246072 3125 246073
rect 2977 245296 3011 246072
rect 3011 245296 3091 246072
rect 3091 245296 3125 246072
rect 3187 246072 3335 246073
rect 3187 245296 3221 246072
rect 3221 245296 3301 246072
rect 3301 245296 3335 246072
rect 3397 246072 3545 246073
rect 3397 245296 3431 246072
rect 3431 245296 3511 246072
rect 3511 245296 3545 246072
rect 3607 246072 3755 246073
rect 3607 245296 3641 246072
rect 3641 245296 3721 246072
rect 3721 245296 3755 246072
rect 3817 246072 3965 246073
rect 3817 245296 3851 246072
rect 3851 245296 3931 246072
rect 3931 245296 3965 246072
rect 4027 246072 4175 246073
rect 4027 245296 4061 246072
rect 4061 245296 4141 246072
rect 4141 245296 4175 246072
rect 4237 246072 4385 246073
rect 4237 245296 4271 246072
rect 4271 245296 4351 246072
rect 4351 245296 4385 246072
rect 4447 246072 4595 246073
rect 4447 245296 4481 246072
rect 4481 245296 4561 246072
rect 4561 245296 4595 246072
rect 4657 246072 4805 246073
rect 4657 245296 4691 246072
rect 4691 245296 4771 246072
rect 4771 245296 4805 246072
rect 4867 246072 5015 246073
rect 4867 245296 4901 246072
rect 4901 245296 4981 246072
rect 4981 245296 5015 246072
rect 5077 246072 5225 246073
rect 5077 245296 5111 246072
rect 5111 245296 5191 246072
rect 5191 245296 5225 246072
rect 5287 246072 5435 246073
rect 5287 245296 5321 246072
rect 5321 245296 5401 246072
rect 5401 245296 5435 246072
rect 5497 246072 5645 246073
rect 5497 245296 5531 246072
rect 5531 245296 5611 246072
rect 5611 245296 5645 246072
rect 5707 246072 5855 246073
rect 5707 245296 5741 246072
rect 5741 245296 5821 246072
rect 5821 245296 5855 246072
rect 5917 246072 6065 246073
rect 5917 245296 5951 246072
rect 5951 245296 6031 246072
rect 6031 245296 6065 246072
rect 6127 246072 6275 246073
rect 6127 245296 6161 246072
rect 6161 245296 6241 246072
rect 6241 245296 6275 246072
rect 6337 246072 6485 246073
rect 6337 245296 6371 246072
rect 6371 245296 6451 246072
rect 6451 245296 6485 246072
rect 6547 246072 6695 246073
rect 6547 245296 6581 246072
rect 6581 245296 6661 246072
rect 6661 245296 6695 246072
rect 6757 246072 6905 246073
rect 6757 245296 6791 246072
rect 6791 245296 6871 246072
rect 6871 245296 6905 246072
rect 6967 246072 7115 246073
rect 6967 245296 7001 246072
rect 7001 245296 7081 246072
rect 7081 245296 7115 246072
rect 7177 246072 7325 246073
rect 7177 245296 7211 246072
rect 7211 245296 7291 246072
rect 7291 245296 7325 246072
rect 7387 246072 7535 246073
rect 7387 245296 7421 246072
rect 7421 245296 7501 246072
rect 7501 245296 7535 246072
rect 7597 246072 7745 246073
rect 7597 245296 7631 246072
rect 7631 245296 7711 246072
rect 7711 245296 7745 246072
rect 7807 246072 7955 246073
rect 7807 245296 7841 246072
rect 7841 245296 7921 246072
rect 7921 245296 7955 246072
rect 8017 246072 8165 246073
rect 8017 245296 8051 246072
rect 8051 245296 8131 246072
rect 8131 245296 8165 246072
rect 8227 246072 8375 246073
rect 8227 245296 8261 246072
rect 8261 245296 8341 246072
rect 8341 245296 8375 246072
rect 8437 246072 8585 246073
rect 8437 245296 8471 246072
rect 8471 245296 8551 246072
rect 8551 245296 8585 246072
rect 8647 246072 8795 246073
rect 8647 245296 8681 246072
rect 8681 245296 8761 246072
rect 8761 245296 8795 246072
rect 8857 246072 9005 246073
rect 8857 245296 8891 246072
rect 8891 245296 8971 246072
rect 8971 245296 9005 246072
rect 9067 246072 9215 246073
rect 9067 245296 9101 246072
rect 9101 245296 9181 246072
rect 9181 245296 9215 246072
rect 9277 246072 9425 246073
rect 9277 245296 9311 246072
rect 9311 245296 9391 246072
rect 9391 245296 9425 246072
rect 9487 246072 9635 246073
rect 9487 245296 9521 246072
rect 9521 245296 9601 246072
rect 9601 245296 9635 246072
rect 9697 246072 9845 246073
rect 9697 245296 9731 246072
rect 9731 245296 9811 246072
rect 9811 245296 9845 246072
rect 9907 246072 10055 246073
rect 9907 245296 9941 246072
rect 9941 245296 10021 246072
rect 10021 245296 10055 246072
rect 10117 246072 10265 246073
rect 10117 245296 10151 246072
rect 10151 245296 10231 246072
rect 10231 245296 10265 246072
rect 10327 246072 10475 246073
rect 10327 245296 10361 246072
rect 10361 245296 10441 246072
rect 10441 245296 10475 246072
rect 10537 246072 10685 246073
rect 10537 245296 10571 246072
rect 10571 245296 10651 246072
rect 10651 245296 10685 246072
rect 10747 246072 10895 246073
rect 10747 245296 10781 246072
rect 10781 245296 10861 246072
rect 10861 245296 10895 246072
rect 10957 246072 11105 246073
rect 10957 245296 10991 246072
rect 10991 245296 11071 246072
rect 11071 245296 11105 246072
rect 11167 246072 11315 246073
rect 11167 245296 11201 246072
rect 11201 245296 11281 246072
rect 11281 245296 11315 246072
rect 11377 246072 11525 246073
rect 11377 245296 11411 246072
rect 11411 245296 11491 246072
rect 11491 245296 11525 246072
rect 11587 246072 11735 246073
rect 11587 245296 11621 246072
rect 11621 245296 11701 246072
rect 11701 245296 11735 246072
rect 11797 246072 11945 246073
rect 11797 245296 11831 246072
rect 11831 245296 11911 246072
rect 11911 245296 11945 246072
rect 12007 246072 12155 246073
rect 12007 245296 12041 246072
rect 12041 245296 12121 246072
rect 12121 245296 12155 246072
rect 12217 246072 12365 246073
rect 12217 245296 12251 246072
rect 12251 245296 12331 246072
rect 12331 245296 12365 246072
rect 12427 246072 12575 246073
rect 12427 245296 12461 246072
rect 12461 245296 12541 246072
rect 12541 245296 12575 246072
rect 12637 246072 12785 246073
rect 12637 245296 12671 246072
rect 12671 245296 12751 246072
rect 12751 245296 12785 246072
rect 12847 246072 12995 246073
rect 12847 245296 12881 246072
rect 12881 245296 12961 246072
rect 12961 245296 12995 246072
rect 13057 246072 13205 246073
rect 13057 245296 13091 246072
rect 13091 245296 13171 246072
rect 13171 245296 13205 246072
rect 13267 246072 13415 246073
rect 13267 245296 13301 246072
rect 13301 245296 13381 246072
rect 13381 245296 13415 246072
rect 13477 246072 13625 246073
rect 13477 245296 13511 246072
rect 13511 245296 13591 246072
rect 13591 245296 13625 246072
rect 13687 246072 13835 246073
rect 13687 245296 13721 246072
rect 13721 245296 13801 246072
rect 13801 245296 13835 246072
rect 13897 246072 14045 246073
rect 13897 245296 13931 246072
rect 13931 245296 14011 246072
rect 14011 245296 14045 246072
rect 14107 246072 14255 246073
rect 14107 245296 14141 246072
rect 14141 245296 14221 246072
rect 14221 245296 14255 246072
rect 14317 246072 14465 246073
rect 14317 245296 14351 246072
rect 14351 245296 14431 246072
rect 14431 245296 14465 246072
rect 14527 246072 14675 246073
rect 14527 245296 14561 246072
rect 14561 245296 14641 246072
rect 14641 245296 14675 246072
rect 14737 246072 14885 246073
rect 14737 245296 14771 246072
rect 14771 245296 14851 246072
rect 14851 245296 14885 246072
rect 14947 246072 15095 246073
rect 14947 245296 14981 246072
rect 14981 245296 15061 246072
rect 15061 245296 15095 246072
rect 15157 246072 15305 246073
rect 15157 245296 15191 246072
rect 15191 245296 15271 246072
rect 15271 245296 15305 246072
rect 15367 246072 15515 246073
rect 15367 245296 15401 246072
rect 15401 245296 15481 246072
rect 15481 245296 15515 246072
rect 15577 246072 15725 246073
rect 15577 245296 15611 246072
rect 15611 245296 15691 246072
rect 15691 245296 15725 246072
rect 15787 246072 15935 246073
rect 15787 245296 15821 246072
rect 15821 245296 15901 246072
rect 15901 245296 15935 246072
rect 15997 246072 16145 246073
rect 15997 245296 16031 246072
rect 16031 245296 16111 246072
rect 16111 245296 16145 246072
rect 16207 246072 16355 246073
rect 16207 245296 16241 246072
rect 16241 245296 16321 246072
rect 16321 245296 16355 246072
rect 16417 246072 16565 246073
rect 16417 245296 16451 246072
rect 16451 245296 16531 246072
rect 16531 245296 16565 246072
rect 16627 246072 16775 246073
rect 16627 245296 16661 246072
rect 16661 245296 16741 246072
rect 16741 245296 16775 246072
rect 16837 246072 16985 246073
rect 16837 245296 16871 246072
rect 16871 245296 16951 246072
rect 16951 245296 16985 246072
rect 17047 246072 17195 246073
rect 17047 245296 17081 246072
rect 17081 245296 17161 246072
rect 17161 245296 17195 246072
rect 17257 246072 17405 246073
rect 17257 245296 17291 246072
rect 17291 245296 17371 246072
rect 17371 245296 17405 246072
rect 17467 246072 17615 246073
rect 17467 245296 17501 246072
rect 17501 245296 17581 246072
rect 17581 245296 17615 246072
rect 17677 246072 17825 246073
rect 17677 245296 17711 246072
rect 17711 245296 17791 246072
rect 17791 245296 17825 246072
rect 17887 246072 18035 246073
rect 17887 245296 17921 246072
rect 17921 245296 18001 246072
rect 18001 245296 18035 246072
rect 18097 246072 18245 246073
rect 18097 245296 18131 246072
rect 18131 245296 18211 246072
rect 18211 245296 18245 246072
rect 18307 246072 18455 246073
rect 18307 245296 18341 246072
rect 18341 245296 18421 246072
rect 18421 245296 18455 246072
rect 18517 246072 18665 246073
rect 18517 245296 18551 246072
rect 18551 245296 18631 246072
rect 18631 245296 18665 246072
rect 18727 246072 18875 246073
rect 18727 245296 18761 246072
rect 18761 245296 18841 246072
rect 18841 245296 18875 246072
rect 18937 246072 19085 246073
rect 18937 245296 18971 246072
rect 18971 245296 19051 246072
rect 19051 245296 19085 246072
rect 19147 246072 19295 246073
rect 19147 245296 19181 246072
rect 19181 245296 19261 246072
rect 19261 245296 19295 246072
rect 19357 246072 19505 246073
rect 19357 245296 19391 246072
rect 19391 245296 19471 246072
rect 19471 245296 19505 246072
rect 19567 246072 19715 246073
rect 19567 245296 19601 246072
rect 19601 245296 19681 246072
rect 19681 245296 19715 246072
rect 19777 246072 19925 246073
rect 19777 245296 19811 246072
rect 19811 245296 19891 246072
rect 19891 245296 19925 246072
rect 19987 246072 20135 246073
rect 19987 245296 20021 246072
rect 20021 245296 20101 246072
rect 20101 245296 20135 246072
rect 20197 246072 20345 246073
rect 20197 245296 20231 246072
rect 20231 245296 20311 246072
rect 20311 245296 20345 246072
rect 20407 246072 20555 246073
rect 20407 245296 20441 246072
rect 20441 245296 20521 246072
rect 20521 245296 20555 246072
rect 20617 246072 20765 246073
rect 20617 245296 20651 246072
rect 20651 245296 20731 246072
rect 20731 245296 20765 246072
rect 20827 246072 20975 246073
rect 20827 245296 20861 246072
rect 20861 245296 20941 246072
rect 20941 245296 20975 246072
rect 21037 246072 21185 246073
rect 21037 245296 21071 246072
rect 21071 245296 21151 246072
rect 21151 245296 21185 246072
rect 21247 246072 21395 246073
rect 21247 245296 21281 246072
rect 21281 245296 21361 246072
rect 21361 245296 21395 246072
rect 21457 246072 21605 246073
rect 21457 245296 21491 246072
rect 21491 245296 21571 246072
rect 21571 245296 21605 246072
rect 21667 246072 21815 246073
rect 21667 245296 21701 246072
rect 21701 245296 21781 246072
rect 21781 245296 21815 246072
rect 21877 246072 22025 246073
rect 21877 245296 21911 246072
rect 21911 245296 21991 246072
rect 21991 245296 22025 246072
rect 22087 246072 22235 246073
rect 22087 245296 22121 246072
rect 22121 245296 22201 246072
rect 22201 245296 22235 246072
rect 22297 246072 22445 246073
rect 22297 245296 22331 246072
rect 22331 245296 22411 246072
rect 22411 245296 22445 246072
rect 22507 246072 22655 246073
rect 22507 245296 22541 246072
rect 22541 245296 22621 246072
rect 22621 245296 22655 246072
rect 22717 246072 22865 246073
rect 22717 245296 22751 246072
rect 22751 245296 22831 246072
rect 22831 245296 22865 246072
rect 22927 246072 23075 246073
rect 22927 245296 22961 246072
rect 22961 245296 23041 246072
rect 23041 245296 23075 246072
rect 23137 246072 23285 246073
rect 23137 245296 23171 246072
rect 23171 245296 23251 246072
rect 23251 245296 23285 246072
rect 23347 246072 23495 246073
rect 23347 245296 23381 246072
rect 23381 245296 23461 246072
rect 23461 245296 23495 246072
rect 23557 246072 23705 246073
rect 23557 245296 23591 246072
rect 23591 245296 23671 246072
rect 23671 245296 23705 246072
rect 23767 246072 23915 246073
rect 23767 245296 23801 246072
rect 23801 245296 23881 246072
rect 23881 245296 23915 246072
rect 23977 246072 24125 246073
rect 23977 245296 24011 246072
rect 24011 245296 24091 246072
rect 24091 245296 24125 246072
rect 24187 246072 24335 246073
rect 24187 245296 24221 246072
rect 24221 245296 24301 246072
rect 24301 245296 24335 246072
rect 24397 246072 24545 246073
rect 24397 245296 24431 246072
rect 24431 245296 24511 246072
rect 24511 245296 24545 246072
rect 24607 246072 24755 246073
rect 24607 245296 24641 246072
rect 24641 245296 24721 246072
rect 24721 245296 24755 246072
rect 24817 246072 24965 246073
rect 24817 245296 24851 246072
rect 24851 245296 24931 246072
rect 24931 245296 24965 246072
rect 25027 246072 25175 246073
rect 25027 245296 25061 246072
rect 25061 245296 25141 246072
rect 25141 245296 25175 246072
rect 25237 246072 25385 246073
rect 25237 245296 25271 246072
rect 25271 245296 25351 246072
rect 25351 245296 25385 246072
rect 25447 246072 25595 246073
rect 25447 245296 25481 246072
rect 25481 245296 25561 246072
rect 25561 245296 25595 246072
rect 25657 246072 25805 246073
rect 25657 245296 25691 246072
rect 25691 245296 25771 246072
rect 25771 245296 25805 246072
rect 25867 246072 26015 246073
rect 25867 245296 25901 246072
rect 25901 245296 25981 246072
rect 25981 245296 26015 246072
rect 26077 246072 26225 246073
rect 26077 245296 26111 246072
rect 26111 245296 26191 246072
rect 26191 245296 26225 246072
rect 26287 246072 26435 246073
rect 26287 245296 26321 246072
rect 26321 245296 26401 246072
rect 26401 245296 26435 246072
rect 26497 246072 26645 246073
rect 26497 245296 26531 246072
rect 26531 245296 26611 246072
rect 26611 245296 26645 246072
rect 26707 246072 26855 246073
rect 26707 245296 26741 246072
rect 26741 245296 26821 246072
rect 26821 245296 26855 246072
rect 26917 246072 27065 246073
rect 26917 245296 26951 246072
rect 26951 245296 27031 246072
rect 27031 245296 27065 246072
rect 27127 246072 27275 246073
rect 27127 245296 27161 246072
rect 27161 245296 27241 246072
rect 27241 245296 27275 246072
rect -4075 244260 -4049 245036
rect -4049 244260 -4015 245036
rect -3953 244260 -3919 245036
rect -3919 244260 -3839 245036
rect -3839 244260 -3805 245036
rect -3743 244260 -3709 245036
rect -3709 244260 -3629 245036
rect -3629 244260 -3595 245036
rect -3533 245036 -3385 245037
rect -3533 244260 -3499 245036
rect -3499 244260 -3419 245036
rect -3419 244260 -3385 245036
rect -3323 245036 -3175 245037
rect -3323 244260 -3289 245036
rect -3289 244260 -3209 245036
rect -3209 244260 -3175 245036
rect -3113 245036 -2965 245037
rect -3113 244260 -3079 245036
rect -3079 244260 -2999 245036
rect -2999 244260 -2965 245036
rect -2903 245036 -2755 245037
rect -2903 244260 -2869 245036
rect -2869 244260 -2789 245036
rect -2789 244260 -2755 245036
rect -2693 245036 -2545 245037
rect -2693 244260 -2659 245036
rect -2659 244260 -2579 245036
rect -2579 244260 -2545 245036
rect -2483 245036 -2335 245037
rect -2483 244260 -2449 245036
rect -2449 244260 -2369 245036
rect -2369 244260 -2335 245036
rect -2273 245036 -2125 245037
rect -2273 244260 -2239 245036
rect -2239 244260 -2159 245036
rect -2159 244260 -2125 245036
rect -2063 245036 -1915 245037
rect -2063 244260 -2029 245036
rect -2029 244260 -1949 245036
rect -1949 244260 -1915 245036
rect -1853 245036 -1705 245037
rect -1853 244260 -1819 245036
rect -1819 244260 -1739 245036
rect -1739 244260 -1705 245036
rect -1643 245036 -1495 245037
rect -1643 244260 -1609 245036
rect -1609 244260 -1529 245036
rect -1529 244260 -1495 245036
rect -1433 245036 -1285 245037
rect -1433 244260 -1399 245036
rect -1399 244260 -1319 245036
rect -1319 244260 -1285 245036
rect -1223 245036 -1075 245037
rect -1223 244260 -1189 245036
rect -1189 244260 -1109 245036
rect -1109 244260 -1075 245036
rect -1013 245036 -865 245037
rect -1013 244260 -979 245036
rect -979 244260 -899 245036
rect -899 244260 -865 245036
rect -803 245036 -655 245037
rect -803 244260 -769 245036
rect -769 244260 -689 245036
rect -689 244260 -655 245036
rect -593 245036 -445 245037
rect -593 244260 -559 245036
rect -559 244260 -479 245036
rect -479 244260 -445 245036
rect -383 245036 -235 245037
rect -383 244260 -349 245036
rect -349 244260 -269 245036
rect -269 244260 -235 245036
rect -173 245036 -25 245037
rect -173 244260 -139 245036
rect -139 244260 -59 245036
rect -59 244260 -25 245036
rect 37 245036 185 245037
rect 37 244260 71 245036
rect 71 244260 151 245036
rect 151 244260 185 245036
rect 247 245036 395 245037
rect 247 244260 281 245036
rect 281 244260 361 245036
rect 361 244260 395 245036
rect 457 245036 605 245037
rect 457 244260 491 245036
rect 491 244260 571 245036
rect 571 244260 605 245036
rect 667 245036 815 245037
rect 667 244260 701 245036
rect 701 244260 781 245036
rect 781 244260 815 245036
rect 877 245036 1025 245037
rect 877 244260 911 245036
rect 911 244260 991 245036
rect 991 244260 1025 245036
rect 1087 245036 1235 245037
rect 1087 244260 1121 245036
rect 1121 244260 1201 245036
rect 1201 244260 1235 245036
rect 1297 245036 1445 245037
rect 1297 244260 1331 245036
rect 1331 244260 1411 245036
rect 1411 244260 1445 245036
rect 1507 245036 1655 245037
rect 1507 244260 1541 245036
rect 1541 244260 1621 245036
rect 1621 244260 1655 245036
rect 1717 245036 1865 245037
rect 1717 244260 1751 245036
rect 1751 244260 1831 245036
rect 1831 244260 1865 245036
rect 1927 245036 2075 245037
rect 1927 244260 1961 245036
rect 1961 244260 2041 245036
rect 2041 244260 2075 245036
rect 2137 245036 2285 245037
rect 2137 244260 2171 245036
rect 2171 244260 2251 245036
rect 2251 244260 2285 245036
rect 2347 245036 2495 245037
rect 2347 244260 2381 245036
rect 2381 244260 2461 245036
rect 2461 244260 2495 245036
rect 2557 245036 2705 245037
rect 2557 244260 2591 245036
rect 2591 244260 2671 245036
rect 2671 244260 2705 245036
rect 2767 245036 2915 245037
rect 2767 244260 2801 245036
rect 2801 244260 2881 245036
rect 2881 244260 2915 245036
rect 2977 245036 3125 245037
rect 2977 244260 3011 245036
rect 3011 244260 3091 245036
rect 3091 244260 3125 245036
rect 3187 245036 3335 245037
rect 3187 244260 3221 245036
rect 3221 244260 3301 245036
rect 3301 244260 3335 245036
rect 3397 245036 3545 245037
rect 3397 244260 3431 245036
rect 3431 244260 3511 245036
rect 3511 244260 3545 245036
rect 3607 245036 3755 245037
rect 3607 244260 3641 245036
rect 3641 244260 3721 245036
rect 3721 244260 3755 245036
rect 3817 245036 3965 245037
rect 3817 244260 3851 245036
rect 3851 244260 3931 245036
rect 3931 244260 3965 245036
rect 4027 245036 4175 245037
rect 4027 244260 4061 245036
rect 4061 244260 4141 245036
rect 4141 244260 4175 245036
rect 4237 245036 4385 245037
rect 4237 244260 4271 245036
rect 4271 244260 4351 245036
rect 4351 244260 4385 245036
rect 4447 245036 4595 245037
rect 4447 244260 4481 245036
rect 4481 244260 4561 245036
rect 4561 244260 4595 245036
rect 4657 245036 4805 245037
rect 4657 244260 4691 245036
rect 4691 244260 4771 245036
rect 4771 244260 4805 245036
rect 4867 245036 5015 245037
rect 4867 244260 4901 245036
rect 4901 244260 4981 245036
rect 4981 244260 5015 245036
rect 5077 245036 5225 245037
rect 5077 244260 5111 245036
rect 5111 244260 5191 245036
rect 5191 244260 5225 245036
rect 5287 245036 5435 245037
rect 5287 244260 5321 245036
rect 5321 244260 5401 245036
rect 5401 244260 5435 245036
rect 5497 245036 5645 245037
rect 5497 244260 5531 245036
rect 5531 244260 5611 245036
rect 5611 244260 5645 245036
rect 5707 245036 5855 245037
rect 5707 244260 5741 245036
rect 5741 244260 5821 245036
rect 5821 244260 5855 245036
rect 5917 245036 6065 245037
rect 5917 244260 5951 245036
rect 5951 244260 6031 245036
rect 6031 244260 6065 245036
rect 6127 245036 6275 245037
rect 6127 244260 6161 245036
rect 6161 244260 6241 245036
rect 6241 244260 6275 245036
rect 6337 245036 6485 245037
rect 6337 244260 6371 245036
rect 6371 244260 6451 245036
rect 6451 244260 6485 245036
rect 6547 245036 6695 245037
rect 6547 244260 6581 245036
rect 6581 244260 6661 245036
rect 6661 244260 6695 245036
rect 6757 245036 6905 245037
rect 6757 244260 6791 245036
rect 6791 244260 6871 245036
rect 6871 244260 6905 245036
rect 6967 245036 7115 245037
rect 6967 244260 7001 245036
rect 7001 244260 7081 245036
rect 7081 244260 7115 245036
rect 7177 245036 7325 245037
rect 7177 244260 7211 245036
rect 7211 244260 7291 245036
rect 7291 244260 7325 245036
rect 7387 245036 7535 245037
rect 7387 244260 7421 245036
rect 7421 244260 7501 245036
rect 7501 244260 7535 245036
rect 7597 245036 7745 245037
rect 7597 244260 7631 245036
rect 7631 244260 7711 245036
rect 7711 244260 7745 245036
rect 7807 245036 7955 245037
rect 7807 244260 7841 245036
rect 7841 244260 7921 245036
rect 7921 244260 7955 245036
rect 8017 245036 8165 245037
rect 8017 244260 8051 245036
rect 8051 244260 8131 245036
rect 8131 244260 8165 245036
rect 8227 245036 8375 245037
rect 8227 244260 8261 245036
rect 8261 244260 8341 245036
rect 8341 244260 8375 245036
rect 8437 245036 8585 245037
rect 8437 244260 8471 245036
rect 8471 244260 8551 245036
rect 8551 244260 8585 245036
rect 8647 245036 8795 245037
rect 8647 244260 8681 245036
rect 8681 244260 8761 245036
rect 8761 244260 8795 245036
rect 8857 245036 9005 245037
rect 8857 244260 8891 245036
rect 8891 244260 8971 245036
rect 8971 244260 9005 245036
rect 9067 245036 9215 245037
rect 9067 244260 9101 245036
rect 9101 244260 9181 245036
rect 9181 244260 9215 245036
rect 9277 245036 9425 245037
rect 9277 244260 9311 245036
rect 9311 244260 9391 245036
rect 9391 244260 9425 245036
rect 9487 245036 9635 245037
rect 9487 244260 9521 245036
rect 9521 244260 9601 245036
rect 9601 244260 9635 245036
rect 9697 245036 9845 245037
rect 9697 244260 9731 245036
rect 9731 244260 9811 245036
rect 9811 244260 9845 245036
rect 9907 245036 10055 245037
rect 9907 244260 9941 245036
rect 9941 244260 10021 245036
rect 10021 244260 10055 245036
rect 10117 245036 10265 245037
rect 10117 244260 10151 245036
rect 10151 244260 10231 245036
rect 10231 244260 10265 245036
rect 10327 245036 10475 245037
rect 10327 244260 10361 245036
rect 10361 244260 10441 245036
rect 10441 244260 10475 245036
rect 10537 245036 10685 245037
rect 10537 244260 10571 245036
rect 10571 244260 10651 245036
rect 10651 244260 10685 245036
rect 10747 245036 10895 245037
rect 10747 244260 10781 245036
rect 10781 244260 10861 245036
rect 10861 244260 10895 245036
rect 10957 245036 11105 245037
rect 10957 244260 10991 245036
rect 10991 244260 11071 245036
rect 11071 244260 11105 245036
rect 11167 245036 11315 245037
rect 11167 244260 11201 245036
rect 11201 244260 11281 245036
rect 11281 244260 11315 245036
rect 11377 245036 11525 245037
rect 11377 244260 11411 245036
rect 11411 244260 11491 245036
rect 11491 244260 11525 245036
rect 11587 245036 11735 245037
rect 11587 244260 11621 245036
rect 11621 244260 11701 245036
rect 11701 244260 11735 245036
rect 11797 245036 11945 245037
rect 11797 244260 11831 245036
rect 11831 244260 11911 245036
rect 11911 244260 11945 245036
rect 12007 245036 12155 245037
rect 12007 244260 12041 245036
rect 12041 244260 12121 245036
rect 12121 244260 12155 245036
rect 12217 245036 12365 245037
rect 12217 244260 12251 245036
rect 12251 244260 12331 245036
rect 12331 244260 12365 245036
rect 12427 245036 12575 245037
rect 12427 244260 12461 245036
rect 12461 244260 12541 245036
rect 12541 244260 12575 245036
rect 12637 245036 12785 245037
rect 12637 244260 12671 245036
rect 12671 244260 12751 245036
rect 12751 244260 12785 245036
rect 12847 245036 12995 245037
rect 12847 244260 12881 245036
rect 12881 244260 12961 245036
rect 12961 244260 12995 245036
rect 13057 245036 13205 245037
rect 13057 244260 13091 245036
rect 13091 244260 13171 245036
rect 13171 244260 13205 245036
rect 13267 245036 13415 245037
rect 13267 244260 13301 245036
rect 13301 244260 13381 245036
rect 13381 244260 13415 245036
rect 13477 245036 13625 245037
rect 13477 244260 13511 245036
rect 13511 244260 13591 245036
rect 13591 244260 13625 245036
rect 13687 245036 13835 245037
rect 13687 244260 13721 245036
rect 13721 244260 13801 245036
rect 13801 244260 13835 245036
rect 13897 245036 14045 245037
rect 13897 244260 13931 245036
rect 13931 244260 14011 245036
rect 14011 244260 14045 245036
rect 14107 245036 14255 245037
rect 14107 244260 14141 245036
rect 14141 244260 14221 245036
rect 14221 244260 14255 245036
rect 14317 245036 14465 245037
rect 14317 244260 14351 245036
rect 14351 244260 14431 245036
rect 14431 244260 14465 245036
rect 14527 245036 14675 245037
rect 14527 244260 14561 245036
rect 14561 244260 14641 245036
rect 14641 244260 14675 245036
rect 14737 245036 14885 245037
rect 14737 244260 14771 245036
rect 14771 244260 14851 245036
rect 14851 244260 14885 245036
rect 14947 245036 15095 245037
rect 14947 244260 14981 245036
rect 14981 244260 15061 245036
rect 15061 244260 15095 245036
rect 15157 245036 15305 245037
rect 15157 244260 15191 245036
rect 15191 244260 15271 245036
rect 15271 244260 15305 245036
rect 15367 245036 15515 245037
rect 15367 244260 15401 245036
rect 15401 244260 15481 245036
rect 15481 244260 15515 245036
rect 15577 245036 15725 245037
rect 15577 244260 15611 245036
rect 15611 244260 15691 245036
rect 15691 244260 15725 245036
rect 15787 245036 15935 245037
rect 15787 244260 15821 245036
rect 15821 244260 15901 245036
rect 15901 244260 15935 245036
rect 15997 245036 16145 245037
rect 15997 244260 16031 245036
rect 16031 244260 16111 245036
rect 16111 244260 16145 245036
rect 16207 245036 16355 245037
rect 16207 244260 16241 245036
rect 16241 244260 16321 245036
rect 16321 244260 16355 245036
rect 16417 245036 16565 245037
rect 16417 244260 16451 245036
rect 16451 244260 16531 245036
rect 16531 244260 16565 245036
rect 16627 245036 16775 245037
rect 16627 244260 16661 245036
rect 16661 244260 16741 245036
rect 16741 244260 16775 245036
rect 16837 245036 16985 245037
rect 16837 244260 16871 245036
rect 16871 244260 16951 245036
rect 16951 244260 16985 245036
rect 17047 245036 17195 245037
rect 17047 244260 17081 245036
rect 17081 244260 17161 245036
rect 17161 244260 17195 245036
rect 17257 245036 17405 245037
rect 17257 244260 17291 245036
rect 17291 244260 17371 245036
rect 17371 244260 17405 245036
rect 17467 245036 17615 245037
rect 17467 244260 17501 245036
rect 17501 244260 17581 245036
rect 17581 244260 17615 245036
rect 17677 245036 17825 245037
rect 17677 244260 17711 245036
rect 17711 244260 17791 245036
rect 17791 244260 17825 245036
rect 17887 245036 18035 245037
rect 17887 244260 17921 245036
rect 17921 244260 18001 245036
rect 18001 244260 18035 245036
rect 18097 245036 18245 245037
rect 18097 244260 18131 245036
rect 18131 244260 18211 245036
rect 18211 244260 18245 245036
rect 18307 245036 18455 245037
rect 18307 244260 18341 245036
rect 18341 244260 18421 245036
rect 18421 244260 18455 245036
rect 18517 245036 18665 245037
rect 18517 244260 18551 245036
rect 18551 244260 18631 245036
rect 18631 244260 18665 245036
rect 18727 245036 18875 245037
rect 18727 244260 18761 245036
rect 18761 244260 18841 245036
rect 18841 244260 18875 245036
rect 18937 245036 19085 245037
rect 18937 244260 18971 245036
rect 18971 244260 19051 245036
rect 19051 244260 19085 245036
rect 19147 245036 19295 245037
rect 19147 244260 19181 245036
rect 19181 244260 19261 245036
rect 19261 244260 19295 245036
rect 19357 245036 19505 245037
rect 19357 244260 19391 245036
rect 19391 244260 19471 245036
rect 19471 244260 19505 245036
rect 19567 245036 19715 245037
rect 19567 244260 19601 245036
rect 19601 244260 19681 245036
rect 19681 244260 19715 245036
rect 19777 245036 19925 245037
rect 19777 244260 19811 245036
rect 19811 244260 19891 245036
rect 19891 244260 19925 245036
rect 19987 245036 20135 245037
rect 19987 244260 20021 245036
rect 20021 244260 20101 245036
rect 20101 244260 20135 245036
rect 20197 245036 20345 245037
rect 20197 244260 20231 245036
rect 20231 244260 20311 245036
rect 20311 244260 20345 245036
rect 20407 245036 20555 245037
rect 20407 244260 20441 245036
rect 20441 244260 20521 245036
rect 20521 244260 20555 245036
rect 20617 245036 20765 245037
rect 20617 244260 20651 245036
rect 20651 244260 20731 245036
rect 20731 244260 20765 245036
rect 20827 245036 20975 245037
rect 20827 244260 20861 245036
rect 20861 244260 20941 245036
rect 20941 244260 20975 245036
rect 21037 245036 21185 245037
rect 21037 244260 21071 245036
rect 21071 244260 21151 245036
rect 21151 244260 21185 245036
rect 21247 245036 21395 245037
rect 21247 244260 21281 245036
rect 21281 244260 21361 245036
rect 21361 244260 21395 245036
rect 21457 245036 21605 245037
rect 21457 244260 21491 245036
rect 21491 244260 21571 245036
rect 21571 244260 21605 245036
rect 21667 245036 21815 245037
rect 21667 244260 21701 245036
rect 21701 244260 21781 245036
rect 21781 244260 21815 245036
rect 21877 245036 22025 245037
rect 21877 244260 21911 245036
rect 21911 244260 21991 245036
rect 21991 244260 22025 245036
rect 22087 245036 22235 245037
rect 22087 244260 22121 245036
rect 22121 244260 22201 245036
rect 22201 244260 22235 245036
rect 22297 245036 22445 245037
rect 22297 244260 22331 245036
rect 22331 244260 22411 245036
rect 22411 244260 22445 245036
rect 22507 245036 22655 245037
rect 22507 244260 22541 245036
rect 22541 244260 22621 245036
rect 22621 244260 22655 245036
rect 22717 245036 22865 245037
rect 22717 244260 22751 245036
rect 22751 244260 22831 245036
rect 22831 244260 22865 245036
rect 22927 245036 23075 245037
rect 22927 244260 22961 245036
rect 22961 244260 23041 245036
rect 23041 244260 23075 245036
rect 23137 245036 23285 245037
rect 23137 244260 23171 245036
rect 23171 244260 23251 245036
rect 23251 244260 23285 245036
rect 23347 245036 23495 245037
rect 23347 244260 23381 245036
rect 23381 244260 23461 245036
rect 23461 244260 23495 245036
rect 23557 245036 23705 245037
rect 23557 244260 23591 245036
rect 23591 244260 23671 245036
rect 23671 244260 23705 245036
rect 23767 245036 23915 245037
rect 23767 244260 23801 245036
rect 23801 244260 23881 245036
rect 23881 244260 23915 245036
rect 23977 245036 24125 245037
rect 23977 244260 24011 245036
rect 24011 244260 24091 245036
rect 24091 244260 24125 245036
rect 24187 245036 24335 245037
rect 24187 244260 24221 245036
rect 24221 244260 24301 245036
rect 24301 244260 24335 245036
rect 24397 245036 24545 245037
rect 24397 244260 24431 245036
rect 24431 244260 24511 245036
rect 24511 244260 24545 245036
rect 24607 245036 24755 245037
rect 24607 244260 24641 245036
rect 24641 244260 24721 245036
rect 24721 244260 24755 245036
rect 24817 245036 24965 245037
rect 24817 244260 24851 245036
rect 24851 244260 24931 245036
rect 24931 244260 24965 245036
rect 25027 245036 25175 245037
rect 25027 244260 25061 245036
rect 25061 244260 25141 245036
rect 25141 244260 25175 245036
rect 25237 245036 25385 245037
rect 25237 244260 25271 245036
rect 25271 244260 25351 245036
rect 25351 244260 25385 245036
rect 25447 245036 25595 245037
rect 25447 244260 25481 245036
rect 25481 244260 25561 245036
rect 25561 244260 25595 245036
rect 25657 245036 25805 245037
rect 25657 244260 25691 245036
rect 25691 244260 25771 245036
rect 25771 244260 25805 245036
rect 25867 245036 26015 245037
rect 25867 244260 25901 245036
rect 25901 244260 25981 245036
rect 25981 244260 26015 245036
rect 26077 245036 26225 245037
rect 26077 244260 26111 245036
rect 26111 244260 26191 245036
rect 26191 244260 26225 245036
rect 26287 245036 26435 245037
rect 26287 244260 26321 245036
rect 26321 244260 26401 245036
rect 26401 244260 26435 245036
rect 26497 245036 26645 245037
rect 26497 244260 26531 245036
rect 26531 244260 26611 245036
rect 26611 244260 26645 245036
rect 26707 245036 26855 245037
rect 26707 244260 26741 245036
rect 26741 244260 26821 245036
rect 26821 244260 26855 245036
rect 26917 245036 27065 245037
rect 26917 244260 26951 245036
rect 26951 244260 27031 245036
rect 27031 244260 27065 245036
rect 27127 245036 27275 245037
rect 27127 244260 27161 245036
rect 27161 244260 27241 245036
rect 27241 244260 27275 245036
rect -4163 243960 27485 244065
rect 27485 243960 27614 244041
rect 27414 243841 27614 243960
<< metal2 >>
rect -4179 264430 -3979 264440
rect -3770 264430 -3570 264440
rect -3979 264317 -3770 264327
rect -3350 264430 -3150 264440
rect -3570 264317 -3350 264327
rect -2930 264430 -2730 264440
rect -3150 264317 -2930 264327
rect -2510 264430 -2310 264440
rect -2730 264317 -2510 264327
rect -2090 264430 -1890 264440
rect -2310 264317 -2090 264327
rect -1670 264430 -1470 264440
rect -1890 264317 -1670 264327
rect -1250 264430 -1050 264440
rect -1470 264317 -1250 264327
rect -830 264430 -630 264440
rect -1050 264317 -830 264327
rect -410 264430 -210 264440
rect -630 264317 -410 264327
rect 10 264430 210 264440
rect -210 264317 10 264327
rect 430 264430 630 264440
rect 210 264317 430 264327
rect 850 264430 1050 264440
rect 630 264317 850 264327
rect 1270 264430 1470 264440
rect 1050 264317 1270 264327
rect 1690 264430 1890 264440
rect 1470 264317 1690 264327
rect 2110 264430 2310 264440
rect 1890 264317 2110 264327
rect 2530 264430 2730 264440
rect 2310 264317 2530 264327
rect 2950 264430 3150 264440
rect 2730 264317 2950 264327
rect 3370 264430 3570 264440
rect 3150 264317 3370 264327
rect 3790 264430 3990 264440
rect 3570 264317 3790 264327
rect 4210 264430 4410 264440
rect 3990 264317 4210 264327
rect 4630 264430 4830 264440
rect 4410 264317 4630 264327
rect 5050 264430 5250 264440
rect 4830 264317 5050 264327
rect 5470 264430 5670 264440
rect 5250 264317 5470 264327
rect 5890 264430 6090 264440
rect 5670 264317 5890 264327
rect 6310 264430 6510 264440
rect 6090 264317 6310 264327
rect 6730 264430 6930 264440
rect 6510 264317 6730 264327
rect 7150 264430 7350 264440
rect 6930 264317 7150 264327
rect 7570 264430 7770 264440
rect 7350 264317 7570 264327
rect 7990 264430 8190 264440
rect 7770 264317 7990 264327
rect 8410 264430 8610 264440
rect 8190 264317 8410 264327
rect 8830 264430 9030 264440
rect 8610 264317 8830 264327
rect 9250 264430 9450 264440
rect 9030 264317 9250 264327
rect 9670 264430 9870 264440
rect 9450 264317 9670 264327
rect 10090 264430 10290 264440
rect 9870 264317 10090 264327
rect 10510 264430 10710 264440
rect 10290 264317 10510 264327
rect 10930 264430 11130 264440
rect 10710 264317 10930 264327
rect 11350 264430 11550 264440
rect 11130 264317 11350 264327
rect 11770 264430 11970 264440
rect 11550 264317 11770 264327
rect 12190 264430 12390 264440
rect 11970 264317 12190 264327
rect 12610 264430 12810 264440
rect 12390 264317 12610 264327
rect 13030 264430 13230 264440
rect 12810 264317 13030 264327
rect 13450 264430 13650 264440
rect 13230 264317 13450 264327
rect 13870 264430 14070 264440
rect 13650 264317 13870 264327
rect 14290 264430 14490 264440
rect 14070 264317 14290 264327
rect 14710 264430 14910 264440
rect 14490 264317 14710 264327
rect 15130 264430 15330 264440
rect 14910 264317 15130 264327
rect 15550 264430 15750 264440
rect 15330 264317 15550 264327
rect 15970 264430 16170 264440
rect 15750 264317 15970 264327
rect 16390 264430 16590 264440
rect 16170 264317 16390 264327
rect 16810 264430 17010 264440
rect 16590 264317 16810 264327
rect 17230 264430 17430 264440
rect 17010 264317 17230 264327
rect 17650 264430 17850 264440
rect 17430 264317 17650 264327
rect 18070 264430 18270 264440
rect 17850 264317 18070 264327
rect 18490 264430 18690 264440
rect 18270 264317 18490 264327
rect 18910 264430 19110 264440
rect 18690 264317 18910 264327
rect 19330 264430 19530 264440
rect 19110 264317 19330 264327
rect 19750 264430 19950 264440
rect 19530 264317 19750 264327
rect 20170 264430 20370 264440
rect 19950 264317 20170 264327
rect 20590 264430 20790 264440
rect 20370 264317 20590 264327
rect 21010 264430 21210 264440
rect 20790 264317 21010 264327
rect 21430 264430 21630 264440
rect 21210 264317 21430 264327
rect 21850 264430 22050 264440
rect 21630 264317 21850 264327
rect 22270 264430 22470 264440
rect 22050 264317 22270 264327
rect 22690 264430 22890 264440
rect 22470 264317 22690 264327
rect 23110 264430 23310 264440
rect 22890 264317 23110 264327
rect 23530 264430 23730 264440
rect 23310 264317 23530 264327
rect 23950 264430 24150 264440
rect 23730 264317 23950 264327
rect 24370 264430 24570 264440
rect 24150 264317 24370 264327
rect 24790 264430 24990 264440
rect 24570 264317 24790 264327
rect 25210 264430 25410 264440
rect 24990 264317 25210 264327
rect 25630 264430 25830 264440
rect 25410 264317 25630 264327
rect 26050 264430 26250 264440
rect 25830 264317 26050 264327
rect 26470 264430 26670 264440
rect 26250 264317 26470 264327
rect 26890 264430 27090 264440
rect 26670 264317 26890 264327
rect 27310 264430 27510 264440
rect 27090 264317 27310 264327
rect -4179 264220 -4163 264230
rect 27486 264220 27510 264230
rect -4163 264202 27486 264212
rect -4070 264026 -4015 264202
rect -4070 263004 -4015 263250
rect -4070 262218 -4015 262228
rect -3963 264026 -3795 264038
rect -3963 263250 -3953 264026
rect -3805 263250 -3795 264026
rect -3963 263004 -3795 263250
rect -3963 262228 -3953 263004
rect -3805 262228 -3795 263004
rect -3963 261962 -3795 262228
rect -3753 264026 -3585 264202
rect -3753 263250 -3743 264026
rect -3595 263250 -3585 264026
rect -3753 263004 -3585 263250
rect -3753 262228 -3743 263004
rect -3595 262228 -3585 263004
rect -3753 262216 -3585 262228
rect -3543 264026 -3375 264038
rect -3543 263250 -3533 264026
rect -3385 263250 -3375 264026
rect -3543 263004 -3375 263250
rect -3543 262228 -3533 263004
rect -3385 262228 -3375 263004
rect -3543 261962 -3375 262228
rect -3333 264026 -3165 264202
rect -3333 263250 -3323 264026
rect -3175 263250 -3165 264026
rect -3333 263004 -3165 263250
rect -3333 262228 -3323 263004
rect -3175 262228 -3165 263004
rect -3333 262216 -3165 262228
rect -3123 264026 -2955 264038
rect -3123 263250 -3113 264026
rect -2965 263250 -2955 264026
rect -3123 263004 -2955 263250
rect -3123 262228 -3113 263004
rect -2965 262228 -2955 263004
rect -3123 261962 -2955 262228
rect -2913 264026 -2745 264202
rect -2913 263250 -2903 264026
rect -2755 263250 -2745 264026
rect -2913 263004 -2745 263250
rect -2913 262228 -2903 263004
rect -2755 262228 -2745 263004
rect -2913 262216 -2745 262228
rect -2703 264026 -2535 264038
rect -2703 263250 -2693 264026
rect -2545 263250 -2535 264026
rect -2703 263004 -2535 263250
rect -2703 262228 -2693 263004
rect -2545 262228 -2535 263004
rect -2703 261962 -2535 262228
rect -2493 264026 -2325 264202
rect -2493 263250 -2483 264026
rect -2335 263250 -2325 264026
rect -2493 263004 -2325 263250
rect -2493 262228 -2483 263004
rect -2335 262228 -2325 263004
rect -2493 262216 -2325 262228
rect -2283 264026 -2115 264038
rect -2283 263250 -2273 264026
rect -2125 263250 -2115 264026
rect -2283 263004 -2115 263250
rect -2283 262228 -2273 263004
rect -2125 262228 -2115 263004
rect -2283 261962 -2115 262228
rect -2073 264026 -1905 264202
rect -2073 263250 -2063 264026
rect -1915 263250 -1905 264026
rect -2073 263004 -1905 263250
rect -2073 262228 -2063 263004
rect -1915 262228 -1905 263004
rect -2073 262216 -1905 262228
rect -1863 264026 -1695 264038
rect -1863 263250 -1853 264026
rect -1705 263250 -1695 264026
rect -1863 263004 -1695 263250
rect -1863 262228 -1853 263004
rect -1705 262228 -1695 263004
rect -1863 261962 -1695 262228
rect -1653 264026 -1485 264202
rect -1653 263250 -1643 264026
rect -1495 263250 -1485 264026
rect -1653 263004 -1485 263250
rect -1653 262228 -1643 263004
rect -1495 262228 -1485 263004
rect -1653 262216 -1485 262228
rect -1443 264026 -1275 264038
rect -1443 263250 -1433 264026
rect -1285 263250 -1275 264026
rect -1443 263004 -1275 263250
rect -1443 262228 -1433 263004
rect -1285 262228 -1275 263004
rect -1443 261962 -1275 262228
rect -1233 264026 -1065 264202
rect -1233 263250 -1223 264026
rect -1075 263250 -1065 264026
rect -1233 263004 -1065 263250
rect -1233 262228 -1223 263004
rect -1075 262228 -1065 263004
rect -1233 262216 -1065 262228
rect -1023 264026 -855 264038
rect -1023 263250 -1013 264026
rect -865 263250 -855 264026
rect -1023 263004 -855 263250
rect -1023 262228 -1013 263004
rect -865 262228 -855 263004
rect -1023 261962 -855 262228
rect -813 264026 -645 264202
rect -813 263250 -803 264026
rect -655 263250 -645 264026
rect -813 263004 -645 263250
rect -813 262228 -803 263004
rect -655 262228 -645 263004
rect -813 262216 -645 262228
rect -603 264026 -435 264038
rect -603 263250 -593 264026
rect -445 263250 -435 264026
rect -603 263004 -435 263250
rect -603 262228 -593 263004
rect -445 262228 -435 263004
rect -603 261962 -435 262228
rect -393 264026 -225 264202
rect -393 263250 -383 264026
rect -235 263250 -225 264026
rect -393 263004 -225 263250
rect -393 262228 -383 263004
rect -235 262228 -225 263004
rect -393 262216 -225 262228
rect -183 264026 -15 264038
rect -183 263250 -173 264026
rect -25 263250 -15 264026
rect -183 263004 -15 263250
rect -183 262228 -173 263004
rect -25 262228 -15 263004
rect -183 261962 -15 262228
rect 27 264026 195 264202
rect 27 263250 37 264026
rect 185 263250 195 264026
rect 27 263004 195 263250
rect 27 262228 37 263004
rect 185 262228 195 263004
rect 27 262216 195 262228
rect 237 264026 405 264038
rect 237 263250 247 264026
rect 395 263250 405 264026
rect 237 263004 405 263250
rect 237 262228 247 263004
rect 395 262228 405 263004
rect 237 261962 405 262228
rect 447 264026 615 264202
rect 447 263250 457 264026
rect 605 263250 615 264026
rect 447 263004 615 263250
rect 447 262228 457 263004
rect 605 262228 615 263004
rect 447 262216 615 262228
rect 657 264026 825 264038
rect 657 263250 667 264026
rect 815 263250 825 264026
rect 657 263004 825 263250
rect 657 262228 667 263004
rect 815 262228 825 263004
rect 657 261962 825 262228
rect 867 264026 1035 264202
rect 867 263250 877 264026
rect 1025 263250 1035 264026
rect 867 263004 1035 263250
rect 867 262228 877 263004
rect 1025 262228 1035 263004
rect 867 262216 1035 262228
rect 1077 264026 1245 264038
rect 1077 263250 1087 264026
rect 1235 263250 1245 264026
rect 1077 263004 1245 263250
rect 1077 262228 1087 263004
rect 1235 262228 1245 263004
rect 1077 261962 1245 262228
rect 1287 264026 1455 264202
rect 1287 263250 1297 264026
rect 1445 263250 1455 264026
rect 1287 263004 1455 263250
rect 1287 262228 1297 263004
rect 1445 262228 1455 263004
rect 1287 262216 1455 262228
rect 1497 264026 1665 264038
rect 1497 263250 1507 264026
rect 1655 263250 1665 264026
rect 1497 263004 1665 263250
rect 1497 262228 1507 263004
rect 1655 262228 1665 263004
rect 1497 261962 1665 262228
rect 1707 264026 1875 264202
rect 1707 263250 1717 264026
rect 1865 263250 1875 264026
rect 1707 263004 1875 263250
rect 1707 262228 1717 263004
rect 1865 262228 1875 263004
rect 1707 262216 1875 262228
rect 1917 264026 2085 264038
rect 1917 263250 1927 264026
rect 2075 263250 2085 264026
rect 1917 263004 2085 263250
rect 1917 262228 1927 263004
rect 2075 262228 2085 263004
rect 1917 261962 2085 262228
rect 2127 264026 2295 264202
rect 2127 263250 2137 264026
rect 2285 263250 2295 264026
rect 2127 263004 2295 263250
rect 2127 262228 2137 263004
rect 2285 262228 2295 263004
rect 2127 262216 2295 262228
rect 2337 264026 2505 264038
rect 2337 263250 2347 264026
rect 2495 263250 2505 264026
rect 2337 263004 2505 263250
rect 2337 262228 2347 263004
rect 2495 262228 2505 263004
rect 2337 261962 2505 262228
rect 2547 264026 2715 264202
rect 2547 263250 2557 264026
rect 2705 263250 2715 264026
rect 2547 263004 2715 263250
rect 2547 262228 2557 263004
rect 2705 262228 2715 263004
rect 2547 262216 2715 262228
rect 2757 264026 2925 264038
rect 2757 263250 2767 264026
rect 2915 263250 2925 264026
rect 2757 263004 2925 263250
rect 2757 262228 2767 263004
rect 2915 262228 2925 263004
rect 2757 261962 2925 262228
rect 2967 264026 3135 264202
rect 2967 263250 2977 264026
rect 3125 263250 3135 264026
rect 2967 263004 3135 263250
rect 2967 262228 2977 263004
rect 3125 262228 3135 263004
rect 2967 262216 3135 262228
rect 3177 264026 3345 264038
rect 3177 263250 3187 264026
rect 3335 263250 3345 264026
rect 3177 263004 3345 263250
rect 3177 262228 3187 263004
rect 3335 262228 3345 263004
rect 3177 261962 3345 262228
rect 3387 264026 3555 264202
rect 3387 263250 3397 264026
rect 3545 263250 3555 264026
rect 3387 263004 3555 263250
rect 3387 262228 3397 263004
rect 3545 262228 3555 263004
rect 3387 262216 3555 262228
rect 3597 264026 3765 264038
rect 3597 263250 3607 264026
rect 3755 263250 3765 264026
rect 3597 263004 3765 263250
rect 3597 262228 3607 263004
rect 3755 262228 3765 263004
rect 3597 261962 3765 262228
rect 3807 264026 3975 264202
rect 3807 263250 3817 264026
rect 3965 263250 3975 264026
rect 3807 263004 3975 263250
rect 3807 262228 3817 263004
rect 3965 262228 3975 263004
rect 3807 262216 3975 262228
rect 4017 264026 4185 264038
rect 4017 263250 4027 264026
rect 4175 263250 4185 264026
rect 4017 263004 4185 263250
rect 4017 262228 4027 263004
rect 4175 262228 4185 263004
rect 4017 261962 4185 262228
rect 4227 264026 4395 264202
rect 4227 263250 4237 264026
rect 4385 263250 4395 264026
rect 4227 263004 4395 263250
rect 4227 262228 4237 263004
rect 4385 262228 4395 263004
rect 4227 262216 4395 262228
rect 4437 264026 4605 264038
rect 4437 263250 4447 264026
rect 4595 263250 4605 264026
rect 4437 263004 4605 263250
rect 4437 262228 4447 263004
rect 4595 262228 4605 263004
rect 4437 261962 4605 262228
rect 4647 264026 4815 264202
rect 4647 263250 4657 264026
rect 4805 263250 4815 264026
rect 4647 263004 4815 263250
rect 4647 262228 4657 263004
rect 4805 262228 4815 263004
rect 4647 262216 4815 262228
rect 4857 264026 5025 264038
rect 4857 263250 4867 264026
rect 5015 263250 5025 264026
rect 4857 263004 5025 263250
rect 4857 262228 4867 263004
rect 5015 262228 5025 263004
rect 4857 261962 5025 262228
rect 5067 264026 5235 264202
rect 5067 263250 5077 264026
rect 5225 263250 5235 264026
rect 5067 263004 5235 263250
rect 5067 262228 5077 263004
rect 5225 262228 5235 263004
rect 5067 262216 5235 262228
rect 5277 264026 5445 264038
rect 5277 263250 5287 264026
rect 5435 263250 5445 264026
rect 5277 263004 5445 263250
rect 5277 262228 5287 263004
rect 5435 262228 5445 263004
rect 5277 261962 5445 262228
rect 5487 264026 5655 264202
rect 5487 263250 5497 264026
rect 5645 263250 5655 264026
rect 5487 263004 5655 263250
rect 5487 262228 5497 263004
rect 5645 262228 5655 263004
rect 5487 262216 5655 262228
rect 5697 264026 5865 264038
rect 5697 263250 5707 264026
rect 5855 263250 5865 264026
rect 5697 263004 5865 263250
rect 5697 262228 5707 263004
rect 5855 262228 5865 263004
rect 5697 261962 5865 262228
rect 5907 264026 6075 264202
rect 5907 263250 5917 264026
rect 6065 263250 6075 264026
rect 5907 263004 6075 263250
rect 5907 262228 5917 263004
rect 6065 262228 6075 263004
rect 5907 262216 6075 262228
rect 6117 264026 6285 264038
rect 6117 263250 6127 264026
rect 6275 263250 6285 264026
rect 6117 263004 6285 263250
rect 6117 262228 6127 263004
rect 6275 262228 6285 263004
rect 6117 261962 6285 262228
rect 6327 264026 6495 264202
rect 6327 263250 6337 264026
rect 6485 263250 6495 264026
rect 6327 263004 6495 263250
rect 6327 262228 6337 263004
rect 6485 262228 6495 263004
rect 6327 262216 6495 262228
rect 6537 264026 6705 264038
rect 6537 263250 6547 264026
rect 6695 263250 6705 264026
rect 6537 263004 6705 263250
rect 6537 262228 6547 263004
rect 6695 262228 6705 263004
rect 6537 261962 6705 262228
rect 6747 264026 6915 264202
rect 6747 263250 6757 264026
rect 6905 263250 6915 264026
rect 6747 263004 6915 263250
rect 6747 262228 6757 263004
rect 6905 262228 6915 263004
rect 6747 262216 6915 262228
rect 6957 264026 7125 264038
rect 6957 263250 6967 264026
rect 7115 263250 7125 264026
rect 6957 263004 7125 263250
rect 6957 262228 6967 263004
rect 7115 262228 7125 263004
rect 6957 261962 7125 262228
rect 7167 264026 7335 264202
rect 7167 263250 7177 264026
rect 7325 263250 7335 264026
rect 7167 263004 7335 263250
rect 7167 262228 7177 263004
rect 7325 262228 7335 263004
rect 7167 262216 7335 262228
rect 7377 264026 7545 264038
rect 7377 263250 7387 264026
rect 7535 263250 7545 264026
rect 7377 263004 7545 263250
rect 7377 262228 7387 263004
rect 7535 262228 7545 263004
rect 7377 261962 7545 262228
rect 7587 264026 7755 264202
rect 7587 263250 7597 264026
rect 7745 263250 7755 264026
rect 7587 263004 7755 263250
rect 7587 262228 7597 263004
rect 7745 262228 7755 263004
rect 7587 262216 7755 262228
rect 7797 264026 7965 264038
rect 7797 263250 7807 264026
rect 7955 263250 7965 264026
rect 7797 263004 7965 263250
rect 7797 262228 7807 263004
rect 7955 262228 7965 263004
rect 7797 261962 7965 262228
rect 8007 264026 8175 264202
rect 8007 263250 8017 264026
rect 8165 263250 8175 264026
rect 8007 263004 8175 263250
rect 8007 262228 8017 263004
rect 8165 262228 8175 263004
rect 8007 262216 8175 262228
rect 8217 264026 8385 264038
rect 8217 263250 8227 264026
rect 8375 263250 8385 264026
rect 8217 263004 8385 263250
rect 8217 262228 8227 263004
rect 8375 262228 8385 263004
rect 8217 261962 8385 262228
rect 8427 264026 8595 264202
rect 8427 263250 8437 264026
rect 8585 263250 8595 264026
rect 8427 263004 8595 263250
rect 8427 262228 8437 263004
rect 8585 262228 8595 263004
rect 8427 262216 8595 262228
rect 8637 264026 8805 264038
rect 8637 263250 8647 264026
rect 8795 263250 8805 264026
rect 8637 263004 8805 263250
rect 8637 262228 8647 263004
rect 8795 262228 8805 263004
rect 8637 261962 8805 262228
rect 8847 264026 9015 264202
rect 8847 263250 8857 264026
rect 9005 263250 9015 264026
rect 8847 263004 9015 263250
rect 8847 262228 8857 263004
rect 9005 262228 9015 263004
rect 8847 262216 9015 262228
rect 9057 264026 9225 264038
rect 9057 263250 9067 264026
rect 9215 263250 9225 264026
rect 9057 263004 9225 263250
rect 9057 262228 9067 263004
rect 9215 262228 9225 263004
rect 9057 261962 9225 262228
rect 9267 264026 9435 264202
rect 9267 263250 9277 264026
rect 9425 263250 9435 264026
rect 9267 263004 9435 263250
rect 9267 262228 9277 263004
rect 9425 262228 9435 263004
rect 9267 262216 9435 262228
rect 9477 264026 9645 264038
rect 9477 263250 9487 264026
rect 9635 263250 9645 264026
rect 9477 263004 9645 263250
rect 9477 262228 9487 263004
rect 9635 262228 9645 263004
rect 9477 261962 9645 262228
rect 9687 264026 9855 264202
rect 9687 263250 9697 264026
rect 9845 263250 9855 264026
rect 9687 263004 9855 263250
rect 9687 262228 9697 263004
rect 9845 262228 9855 263004
rect 9687 262216 9855 262228
rect 9897 264026 10065 264038
rect 9897 263250 9907 264026
rect 10055 263250 10065 264026
rect 9897 263004 10065 263250
rect 9897 262228 9907 263004
rect 10055 262228 10065 263004
rect 9897 261962 10065 262228
rect 10107 264026 10275 264202
rect 10107 263250 10117 264026
rect 10265 263250 10275 264026
rect 10107 263004 10275 263250
rect 10107 262228 10117 263004
rect 10265 262228 10275 263004
rect 10107 262216 10275 262228
rect 10317 264026 10485 264038
rect 10317 263250 10327 264026
rect 10475 263250 10485 264026
rect 10317 263004 10485 263250
rect 10317 262228 10327 263004
rect 10475 262228 10485 263004
rect 10317 261962 10485 262228
rect 10527 264026 10695 264202
rect 10527 263250 10537 264026
rect 10685 263250 10695 264026
rect 10527 263004 10695 263250
rect 10527 262228 10537 263004
rect 10685 262228 10695 263004
rect 10527 262216 10695 262228
rect 10737 264026 10905 264038
rect 10737 263250 10747 264026
rect 10895 263250 10905 264026
rect 10737 263004 10905 263250
rect 10737 262228 10747 263004
rect 10895 262228 10905 263004
rect 10737 261962 10905 262228
rect 10947 264026 11115 264202
rect 10947 263250 10957 264026
rect 11105 263250 11115 264026
rect 10947 263004 11115 263250
rect 10947 262228 10957 263004
rect 11105 262228 11115 263004
rect 10947 262216 11115 262228
rect 11157 264026 11325 264038
rect 11157 263250 11167 264026
rect 11315 263250 11325 264026
rect 11157 263004 11325 263250
rect 11157 262228 11167 263004
rect 11315 262228 11325 263004
rect 11157 261962 11325 262228
rect 11367 264026 11535 264202
rect 11367 263250 11377 264026
rect 11525 263250 11535 264026
rect 11367 263004 11535 263250
rect 11367 262228 11377 263004
rect 11525 262228 11535 263004
rect 11367 262216 11535 262228
rect 11577 264026 11745 264038
rect 11577 263250 11587 264026
rect 11735 263250 11745 264026
rect 11577 263004 11745 263250
rect 11577 262228 11587 263004
rect 11735 262228 11745 263004
rect 11577 261962 11745 262228
rect 11787 264026 11955 264202
rect 11787 263250 11797 264026
rect 11945 263250 11955 264026
rect 11787 263004 11955 263250
rect 11787 262228 11797 263004
rect 11945 262228 11955 263004
rect 11787 262216 11955 262228
rect 11997 264026 12165 264038
rect 11997 263250 12007 264026
rect 12155 263250 12165 264026
rect 11997 263004 12165 263250
rect 11997 262228 12007 263004
rect 12155 262228 12165 263004
rect 11997 261962 12165 262228
rect 12207 264026 12375 264202
rect 12207 263250 12217 264026
rect 12365 263250 12375 264026
rect 12207 263004 12375 263250
rect 12207 262228 12217 263004
rect 12365 262228 12375 263004
rect 12207 262216 12375 262228
rect 12417 264026 12585 264038
rect 12417 263250 12427 264026
rect 12575 263250 12585 264026
rect 12417 263004 12585 263250
rect 12417 262228 12427 263004
rect 12575 262228 12585 263004
rect 12417 261962 12585 262228
rect 12627 264026 12795 264202
rect 12627 263250 12637 264026
rect 12785 263250 12795 264026
rect 12627 263004 12795 263250
rect 12627 262228 12637 263004
rect 12785 262228 12795 263004
rect 12627 262216 12795 262228
rect 12837 264026 13005 264038
rect 12837 263250 12847 264026
rect 12995 263250 13005 264026
rect 12837 263004 13005 263250
rect 12837 262228 12847 263004
rect 12995 262228 13005 263004
rect 12837 261962 13005 262228
rect 13047 264026 13215 264202
rect 13047 263250 13057 264026
rect 13205 263250 13215 264026
rect 13047 263004 13215 263250
rect 13047 262228 13057 263004
rect 13205 262228 13215 263004
rect 13047 262216 13215 262228
rect 13257 264026 13425 264038
rect 13257 263250 13267 264026
rect 13415 263250 13425 264026
rect 13257 263004 13425 263250
rect 13257 262228 13267 263004
rect 13415 262228 13425 263004
rect 13257 261962 13425 262228
rect 13467 264026 13635 264202
rect 13467 263250 13477 264026
rect 13625 263250 13635 264026
rect 13467 263004 13635 263250
rect 13467 262228 13477 263004
rect 13625 262228 13635 263004
rect 13467 262216 13635 262228
rect 13677 264026 13845 264038
rect 13677 263250 13687 264026
rect 13835 263250 13845 264026
rect 13677 263004 13845 263250
rect 13677 262228 13687 263004
rect 13835 262228 13845 263004
rect 13677 261962 13845 262228
rect 13887 264026 14055 264202
rect 13887 263250 13897 264026
rect 14045 263250 14055 264026
rect 13887 263004 14055 263250
rect 13887 262228 13897 263004
rect 14045 262228 14055 263004
rect 13887 262216 14055 262228
rect 14097 264026 14265 264038
rect 14097 263250 14107 264026
rect 14255 263250 14265 264026
rect 14097 263004 14265 263250
rect 14097 262228 14107 263004
rect 14255 262228 14265 263004
rect 14097 261962 14265 262228
rect 14307 264026 14475 264202
rect 14307 263250 14317 264026
rect 14465 263250 14475 264026
rect 14307 263004 14475 263250
rect 14307 262228 14317 263004
rect 14465 262228 14475 263004
rect 14307 262216 14475 262228
rect 14517 264026 14685 264038
rect 14517 263250 14527 264026
rect 14675 263250 14685 264026
rect 14517 263004 14685 263250
rect 14517 262228 14527 263004
rect 14675 262228 14685 263004
rect 14517 261962 14685 262228
rect 14727 264026 14895 264202
rect 14727 263250 14737 264026
rect 14885 263250 14895 264026
rect 14727 263004 14895 263250
rect 14727 262228 14737 263004
rect 14885 262228 14895 263004
rect 14727 262216 14895 262228
rect 14937 264026 15105 264038
rect 14937 263250 14947 264026
rect 15095 263250 15105 264026
rect 14937 263004 15105 263250
rect 14937 262228 14947 263004
rect 15095 262228 15105 263004
rect 14937 261962 15105 262228
rect 15147 264026 15315 264202
rect 15147 263250 15157 264026
rect 15305 263250 15315 264026
rect 15147 263004 15315 263250
rect 15147 262228 15157 263004
rect 15305 262228 15315 263004
rect 15147 262216 15315 262228
rect 15357 264026 15525 264038
rect 15357 263250 15367 264026
rect 15515 263250 15525 264026
rect 15357 263004 15525 263250
rect 15357 262228 15367 263004
rect 15515 262228 15525 263004
rect 15357 261962 15525 262228
rect 15567 264026 15735 264202
rect 15567 263250 15577 264026
rect 15725 263250 15735 264026
rect 15567 263004 15735 263250
rect 15567 262228 15577 263004
rect 15725 262228 15735 263004
rect 15567 262216 15735 262228
rect 15777 264026 15945 264038
rect 15777 263250 15787 264026
rect 15935 263250 15945 264026
rect 15777 263004 15945 263250
rect 15777 262228 15787 263004
rect 15935 262228 15945 263004
rect 15777 261962 15945 262228
rect 15987 264026 16155 264202
rect 15987 263250 15997 264026
rect 16145 263250 16155 264026
rect 15987 263004 16155 263250
rect 15987 262228 15997 263004
rect 16145 262228 16155 263004
rect 15987 262216 16155 262228
rect 16197 264026 16365 264038
rect 16197 263250 16207 264026
rect 16355 263250 16365 264026
rect 16197 263004 16365 263250
rect 16197 262228 16207 263004
rect 16355 262228 16365 263004
rect 16197 261962 16365 262228
rect 16407 264026 16575 264202
rect 16407 263250 16417 264026
rect 16565 263250 16575 264026
rect 16407 263004 16575 263250
rect 16407 262228 16417 263004
rect 16565 262228 16575 263004
rect 16407 262216 16575 262228
rect 16617 264026 16785 264038
rect 16617 263250 16627 264026
rect 16775 263250 16785 264026
rect 16617 263004 16785 263250
rect 16617 262228 16627 263004
rect 16775 262228 16785 263004
rect 16617 261962 16785 262228
rect 16827 264026 16995 264202
rect 16827 263250 16837 264026
rect 16985 263250 16995 264026
rect 16827 263004 16995 263250
rect 16827 262228 16837 263004
rect 16985 262228 16995 263004
rect 16827 262216 16995 262228
rect 17037 264026 17205 264038
rect 17037 263250 17047 264026
rect 17195 263250 17205 264026
rect 17037 263004 17205 263250
rect 17037 262228 17047 263004
rect 17195 262228 17205 263004
rect 17037 261962 17205 262228
rect 17247 264026 17415 264202
rect 17247 263250 17257 264026
rect 17405 263250 17415 264026
rect 17247 263004 17415 263250
rect 17247 262228 17257 263004
rect 17405 262228 17415 263004
rect 17247 262216 17415 262228
rect 17457 264026 17625 264038
rect 17457 263250 17467 264026
rect 17615 263250 17625 264026
rect 17457 263004 17625 263250
rect 17457 262228 17467 263004
rect 17615 262228 17625 263004
rect 17457 261962 17625 262228
rect 17667 264026 17835 264202
rect 17667 263250 17677 264026
rect 17825 263250 17835 264026
rect 17667 263004 17835 263250
rect 17667 262228 17677 263004
rect 17825 262228 17835 263004
rect 17667 262216 17835 262228
rect 17877 264026 18045 264038
rect 17877 263250 17887 264026
rect 18035 263250 18045 264026
rect 17877 263004 18045 263250
rect 17877 262228 17887 263004
rect 18035 262228 18045 263004
rect 17877 261962 18045 262228
rect 18087 264026 18255 264202
rect 18087 263250 18097 264026
rect 18245 263250 18255 264026
rect 18087 263004 18255 263250
rect 18087 262228 18097 263004
rect 18245 262228 18255 263004
rect 18087 262216 18255 262228
rect 18297 264026 18465 264038
rect 18297 263250 18307 264026
rect 18455 263250 18465 264026
rect 18297 263004 18465 263250
rect 18297 262228 18307 263004
rect 18455 262228 18465 263004
rect 18297 261962 18465 262228
rect 18507 264026 18675 264202
rect 18507 263250 18517 264026
rect 18665 263250 18675 264026
rect 18507 263004 18675 263250
rect 18507 262228 18517 263004
rect 18665 262228 18675 263004
rect 18507 262216 18675 262228
rect 18717 264026 18885 264038
rect 18717 263250 18727 264026
rect 18875 263250 18885 264026
rect 18717 263004 18885 263250
rect 18717 262228 18727 263004
rect 18875 262228 18885 263004
rect 18717 261962 18885 262228
rect 18927 264026 19095 264202
rect 18927 263250 18937 264026
rect 19085 263250 19095 264026
rect 18927 263004 19095 263250
rect 18927 262228 18937 263004
rect 19085 262228 19095 263004
rect 18927 262216 19095 262228
rect 19137 264026 19305 264038
rect 19137 263250 19147 264026
rect 19295 263250 19305 264026
rect 19137 263004 19305 263250
rect 19137 262228 19147 263004
rect 19295 262228 19305 263004
rect 19137 261962 19305 262228
rect 19347 264026 19515 264202
rect 19347 263250 19357 264026
rect 19505 263250 19515 264026
rect 19347 263004 19515 263250
rect 19347 262228 19357 263004
rect 19505 262228 19515 263004
rect 19347 262216 19515 262228
rect 19557 264026 19725 264038
rect 19557 263250 19567 264026
rect 19715 263250 19725 264026
rect 19557 263004 19725 263250
rect 19557 262228 19567 263004
rect 19715 262228 19725 263004
rect 19557 261962 19725 262228
rect 19767 264026 19935 264202
rect 19767 263250 19777 264026
rect 19925 263250 19935 264026
rect 19767 263004 19935 263250
rect 19767 262228 19777 263004
rect 19925 262228 19935 263004
rect 19767 262216 19935 262228
rect 19977 264026 20145 264038
rect 19977 263250 19987 264026
rect 20135 263250 20145 264026
rect 19977 263004 20145 263250
rect 19977 262228 19987 263004
rect 20135 262228 20145 263004
rect 19977 261962 20145 262228
rect 20187 264026 20355 264202
rect 20187 263250 20197 264026
rect 20345 263250 20355 264026
rect 20187 263004 20355 263250
rect 20187 262228 20197 263004
rect 20345 262228 20355 263004
rect 20187 262216 20355 262228
rect 20397 264026 20565 264038
rect 20397 263250 20407 264026
rect 20555 263250 20565 264026
rect 20397 263004 20565 263250
rect 20397 262228 20407 263004
rect 20555 262228 20565 263004
rect 20397 261962 20565 262228
rect 20607 264026 20775 264202
rect 20607 263250 20617 264026
rect 20765 263250 20775 264026
rect 20607 263004 20775 263250
rect 20607 262228 20617 263004
rect 20765 262228 20775 263004
rect 20607 262216 20775 262228
rect 20817 264026 20985 264038
rect 20817 263250 20827 264026
rect 20975 263250 20985 264026
rect 20817 263004 20985 263250
rect 20817 262228 20827 263004
rect 20975 262228 20985 263004
rect 20817 261962 20985 262228
rect 21027 264026 21195 264202
rect 21027 263250 21037 264026
rect 21185 263250 21195 264026
rect 21027 263004 21195 263250
rect 21027 262228 21037 263004
rect 21185 262228 21195 263004
rect 21027 262216 21195 262228
rect 21237 264026 21405 264038
rect 21237 263250 21247 264026
rect 21395 263250 21405 264026
rect 21237 263004 21405 263250
rect 21237 262228 21247 263004
rect 21395 262228 21405 263004
rect 21237 261962 21405 262228
rect 21447 264026 21615 264202
rect 21447 263250 21457 264026
rect 21605 263250 21615 264026
rect 21447 263004 21615 263250
rect 21447 262228 21457 263004
rect 21605 262228 21615 263004
rect 21447 262216 21615 262228
rect 21657 264026 21825 264038
rect 21657 263250 21667 264026
rect 21815 263250 21825 264026
rect 21657 263004 21825 263250
rect 21657 262228 21667 263004
rect 21815 262228 21825 263004
rect 21657 261962 21825 262228
rect 21867 264026 22035 264202
rect 21867 263250 21877 264026
rect 22025 263250 22035 264026
rect 21867 263004 22035 263250
rect 21867 262228 21877 263004
rect 22025 262228 22035 263004
rect 21867 262216 22035 262228
rect 22077 264026 22245 264038
rect 22077 263250 22087 264026
rect 22235 263250 22245 264026
rect 22077 263004 22245 263250
rect 22077 262228 22087 263004
rect 22235 262228 22245 263004
rect 22077 261962 22245 262228
rect 22287 264026 22455 264202
rect 22287 263250 22297 264026
rect 22445 263250 22455 264026
rect 22287 263004 22455 263250
rect 22287 262228 22297 263004
rect 22445 262228 22455 263004
rect 22287 262216 22455 262228
rect 22497 264026 22665 264038
rect 22497 263250 22507 264026
rect 22655 263250 22665 264026
rect 22497 263004 22665 263250
rect 22497 262228 22507 263004
rect 22655 262228 22665 263004
rect 22497 261962 22665 262228
rect 22707 264026 22875 264202
rect 22707 263250 22717 264026
rect 22865 263250 22875 264026
rect 22707 263004 22875 263250
rect 22707 262228 22717 263004
rect 22865 262228 22875 263004
rect 22707 262216 22875 262228
rect 22917 264026 23085 264038
rect 22917 263250 22927 264026
rect 23075 263250 23085 264026
rect 22917 263004 23085 263250
rect 22917 262228 22927 263004
rect 23075 262228 23085 263004
rect 22917 261962 23085 262228
rect 23127 264026 23295 264202
rect 23127 263250 23137 264026
rect 23285 263250 23295 264026
rect 23127 263004 23295 263250
rect 23127 262228 23137 263004
rect 23285 262228 23295 263004
rect 23127 262216 23295 262228
rect 23337 264026 23505 264038
rect 23337 263250 23347 264026
rect 23495 263250 23505 264026
rect 23337 263004 23505 263250
rect 23337 262228 23347 263004
rect 23495 262228 23505 263004
rect 23337 261962 23505 262228
rect 23547 264026 23715 264202
rect 23547 263250 23557 264026
rect 23705 263250 23715 264026
rect 23547 263004 23715 263250
rect 23547 262228 23557 263004
rect 23705 262228 23715 263004
rect 23547 262216 23715 262228
rect 23757 264026 23925 264038
rect 23757 263250 23767 264026
rect 23915 263250 23925 264026
rect 23757 263004 23925 263250
rect 23757 262228 23767 263004
rect 23915 262228 23925 263004
rect 23757 261962 23925 262228
rect 23967 264026 24135 264202
rect 23967 263250 23977 264026
rect 24125 263250 24135 264026
rect 23967 263004 24135 263250
rect 23967 262228 23977 263004
rect 24125 262228 24135 263004
rect 23967 262216 24135 262228
rect 24177 264026 24345 264038
rect 24177 263250 24187 264026
rect 24335 263250 24345 264026
rect 24177 263004 24345 263250
rect 24177 262228 24187 263004
rect 24335 262228 24345 263004
rect 24177 261962 24345 262228
rect 24387 264026 24555 264202
rect 24387 263250 24397 264026
rect 24545 263250 24555 264026
rect 24387 263004 24555 263250
rect 24387 262228 24397 263004
rect 24545 262228 24555 263004
rect 24387 262216 24555 262228
rect 24597 264026 24765 264038
rect 24597 263250 24607 264026
rect 24755 263250 24765 264026
rect 24597 263004 24765 263250
rect 24597 262228 24607 263004
rect 24755 262228 24765 263004
rect 24597 261962 24765 262228
rect 24807 264026 24975 264202
rect 24807 263250 24817 264026
rect 24965 263250 24975 264026
rect 24807 263004 24975 263250
rect 24807 262228 24817 263004
rect 24965 262228 24975 263004
rect 24807 262216 24975 262228
rect 25017 264026 25185 264038
rect 25017 263250 25027 264026
rect 25175 263250 25185 264026
rect 25017 263004 25185 263250
rect 25017 262228 25027 263004
rect 25175 262228 25185 263004
rect 25017 261962 25185 262228
rect 25227 264026 25395 264202
rect 25227 263250 25237 264026
rect 25385 263250 25395 264026
rect 25227 263004 25395 263250
rect 25227 262228 25237 263004
rect 25385 262228 25395 263004
rect 25227 262216 25395 262228
rect 25437 264026 25605 264038
rect 25437 263250 25447 264026
rect 25595 263250 25605 264026
rect 25437 263004 25605 263250
rect 25437 262228 25447 263004
rect 25595 262228 25605 263004
rect 25437 261962 25605 262228
rect 25647 264026 25815 264202
rect 25647 263250 25657 264026
rect 25805 263250 25815 264026
rect 25647 263004 25815 263250
rect 25647 262228 25657 263004
rect 25805 262228 25815 263004
rect 25647 262216 25815 262228
rect 25857 264026 26025 264038
rect 25857 263250 25867 264026
rect 26015 263250 26025 264026
rect 25857 263004 26025 263250
rect 25857 262228 25867 263004
rect 26015 262228 26025 263004
rect 25857 261962 26025 262228
rect 26067 264026 26235 264202
rect 26067 263250 26077 264026
rect 26225 263250 26235 264026
rect 26067 263004 26235 263250
rect 26067 262228 26077 263004
rect 26225 262228 26235 263004
rect 26067 262216 26235 262228
rect 26277 264026 26445 264038
rect 26277 263250 26287 264026
rect 26435 263250 26445 264026
rect 26277 263004 26445 263250
rect 26277 262228 26287 263004
rect 26435 262228 26445 263004
rect 26277 261962 26445 262228
rect 26487 264026 26655 264202
rect 26487 263250 26497 264026
rect 26645 263250 26655 264026
rect 26487 263004 26655 263250
rect 26487 262228 26497 263004
rect 26645 262228 26655 263004
rect 26487 262216 26655 262228
rect 26697 264026 26865 264038
rect 26697 263250 26707 264026
rect 26855 263250 26865 264026
rect 26697 263004 26865 263250
rect 26697 262228 26707 263004
rect 26855 262228 26865 263004
rect 26697 261962 26865 262228
rect 26907 264026 27075 264202
rect 26907 263250 26917 264026
rect 27065 263250 27075 264026
rect 26907 263004 27075 263250
rect 26907 262228 26917 263004
rect 27065 262228 27075 263004
rect 26907 262216 27075 262228
rect 27117 264026 27285 264038
rect 27117 263250 27127 264026
rect 27275 263250 27285 264026
rect 27117 263004 27285 263250
rect 27117 262228 27127 263004
rect 27275 262228 27285 263004
rect 27117 261962 27285 262228
rect -3980 261952 -3780 261962
rect -3980 261742 -3780 261752
rect -3560 261952 -3360 261962
rect -3560 261742 -3360 261752
rect -3140 261952 -2940 261962
rect -3140 261742 -2940 261752
rect -2720 261952 -2520 261962
rect -2720 261742 -2520 261752
rect -2300 261952 -2100 261962
rect -2300 261742 -2100 261752
rect -1880 261952 -1680 261962
rect -1880 261742 -1680 261752
rect -1460 261952 -1260 261962
rect -1460 261742 -1260 261752
rect -1040 261952 -840 261962
rect -1040 261742 -840 261752
rect -620 261952 -420 261962
rect -620 261742 -420 261752
rect -200 261952 0 261962
rect -200 261742 0 261752
rect 220 261952 420 261962
rect 220 261742 420 261752
rect 640 261952 840 261962
rect 640 261742 840 261752
rect 1060 261952 1260 261962
rect 1060 261742 1260 261752
rect 1480 261952 1680 261962
rect 1480 261742 1680 261752
rect 1900 261952 2100 261962
rect 1900 261742 2100 261752
rect 2320 261952 2520 261962
rect 2320 261742 2520 261752
rect 2740 261952 2940 261962
rect 2740 261742 2940 261752
rect 3160 261952 3360 261962
rect 3160 261742 3360 261752
rect 3580 261952 3780 261962
rect 3580 261742 3780 261752
rect 4000 261952 4200 261962
rect 4000 261742 4200 261752
rect 4420 261952 4620 261962
rect 4420 261742 4620 261752
rect 4840 261952 5040 261962
rect 4840 261742 5040 261752
rect 5260 261952 5460 261962
rect 5260 261742 5460 261752
rect 5680 261952 5880 261962
rect 5680 261742 5880 261752
rect 6100 261952 6300 261962
rect 6100 261742 6300 261752
rect 6520 261952 6720 261962
rect 6520 261742 6720 261752
rect 6940 261952 7140 261962
rect 6940 261742 7140 261752
rect 7360 261952 7560 261962
rect 7360 261742 7560 261752
rect 7780 261952 7980 261962
rect 7780 261742 7980 261752
rect 8200 261952 8400 261962
rect 8200 261742 8400 261752
rect 8620 261952 8820 261962
rect 8620 261742 8820 261752
rect 9040 261952 9240 261962
rect 9040 261742 9240 261752
rect 9460 261952 9660 261962
rect 9460 261742 9660 261752
rect 9880 261952 10080 261962
rect 9880 261742 10080 261752
rect 10300 261952 10500 261962
rect 10300 261742 10500 261752
rect 10720 261952 10920 261962
rect 10720 261742 10920 261752
rect 11140 261952 11340 261962
rect 11140 261742 11340 261752
rect 11560 261952 11760 261962
rect 11560 261742 11760 261752
rect 11980 261952 12180 261962
rect 11980 261742 12180 261752
rect 12400 261952 12600 261962
rect 12400 261742 12600 261752
rect 12820 261952 13020 261962
rect 12820 261742 13020 261752
rect 13240 261952 13440 261962
rect 13240 261742 13440 261752
rect 13660 261952 13860 261962
rect 13660 261742 13860 261752
rect 14080 261952 14280 261962
rect 14080 261742 14280 261752
rect 14500 261952 14700 261962
rect 14500 261742 14700 261752
rect 14920 261952 15120 261962
rect 14920 261742 15120 261752
rect 15340 261952 15540 261962
rect 15340 261742 15540 261752
rect 15760 261952 15960 261962
rect 15760 261742 15960 261752
rect 16180 261952 16380 261962
rect 16180 261742 16380 261752
rect 16600 261952 16800 261962
rect 16600 261742 16800 261752
rect 17020 261952 17220 261962
rect 17020 261742 17220 261752
rect 17440 261952 17640 261962
rect 17440 261742 17640 261752
rect 17860 261952 18060 261962
rect 17860 261742 18060 261752
rect 18280 261952 18480 261962
rect 18280 261742 18480 261752
rect 18700 261952 18900 261962
rect 18700 261742 18900 261752
rect 19120 261952 19320 261962
rect 19120 261742 19320 261752
rect 19540 261952 19740 261962
rect 19540 261742 19740 261752
rect 19960 261952 20160 261962
rect 19960 261742 20160 261752
rect 20380 261952 20580 261962
rect 20380 261742 20580 261752
rect 20800 261952 21000 261962
rect 20800 261742 21000 261752
rect 21220 261952 21420 261962
rect 21220 261742 21420 261752
rect 21640 261952 21840 261962
rect 21640 261742 21840 261752
rect 22060 261952 22260 261962
rect 22060 261742 22260 261752
rect 22480 261952 22680 261962
rect 22480 261742 22680 261752
rect 22900 261952 23100 261962
rect 22900 261742 23100 261752
rect 23320 261952 23520 261962
rect 23320 261742 23520 261752
rect 23740 261952 23940 261962
rect 23740 261742 23940 261752
rect 24160 261952 24360 261962
rect 24160 261742 24360 261752
rect 24580 261952 24780 261962
rect 24580 261742 24780 261752
rect 25000 261952 25200 261962
rect 25000 261742 25200 261752
rect 25420 261952 25620 261962
rect 25420 261742 25620 261752
rect 25840 261952 26040 261962
rect 25840 261742 26040 261752
rect 26260 261952 26460 261962
rect 26260 261742 26460 261752
rect 26680 261952 26880 261962
rect 26680 261742 26880 261752
rect 27100 261952 27300 261962
rect 27100 261742 27300 261752
rect -3979 254947 -3779 254957
rect -3979 254737 -3779 254747
rect -3559 254947 -3359 254957
rect -3559 254737 -3359 254747
rect -3139 254947 -2939 254957
rect -3139 254737 -2939 254747
rect -2719 254947 -2519 254957
rect -2719 254737 -2519 254747
rect -2299 254947 -2099 254957
rect -2299 254737 -2099 254747
rect -1879 254947 -1679 254957
rect -1879 254737 -1679 254747
rect -1459 254947 -1259 254957
rect -1459 254737 -1259 254747
rect -1039 254947 -839 254957
rect -1039 254737 -839 254747
rect -619 254947 -419 254957
rect -619 254737 -419 254747
rect -199 254947 1 254957
rect -199 254737 1 254747
rect 221 254947 421 254957
rect 221 254737 421 254747
rect 641 254947 841 254957
rect 641 254737 841 254747
rect 1061 254947 1261 254957
rect 1061 254737 1261 254747
rect 1481 254947 1681 254957
rect 1481 254737 1681 254747
rect 1901 254947 2101 254957
rect 1901 254737 2101 254747
rect 2321 254947 2521 254957
rect 2321 254737 2521 254747
rect 2741 254947 2941 254957
rect 2741 254737 2941 254747
rect 3161 254947 3361 254957
rect 3161 254737 3361 254747
rect 3581 254947 3781 254957
rect 3581 254737 3781 254747
rect 4001 254947 4201 254957
rect 4001 254737 4201 254747
rect 4421 254947 4621 254957
rect 4421 254737 4621 254747
rect 4841 254947 5041 254957
rect 4841 254737 5041 254747
rect 5261 254947 5461 254957
rect 5261 254737 5461 254747
rect 5681 254947 5881 254957
rect 5681 254737 5881 254747
rect 6101 254947 6301 254957
rect 6101 254737 6301 254747
rect 6521 254947 6721 254957
rect 6521 254737 6721 254747
rect 6941 254947 7141 254957
rect 6941 254737 7141 254747
rect 7361 254947 7561 254957
rect 7361 254737 7561 254747
rect 7781 254947 7981 254957
rect 7781 254737 7981 254747
rect 8201 254947 8401 254957
rect 8201 254737 8401 254747
rect 8621 254947 8821 254957
rect 8621 254737 8821 254747
rect 9041 254947 9241 254957
rect 9041 254737 9241 254747
rect 9461 254947 9661 254957
rect 9461 254737 9661 254747
rect 9881 254947 10081 254957
rect 9881 254737 10081 254747
rect 10301 254947 10501 254957
rect 10301 254737 10501 254747
rect 10721 254947 10921 254957
rect 10721 254737 10921 254747
rect 11141 254947 11341 254957
rect 11141 254737 11341 254747
rect 11561 254947 11761 254957
rect 11561 254737 11761 254747
rect 11981 254947 12181 254957
rect 11981 254737 12181 254747
rect 12401 254947 12601 254957
rect 12401 254737 12601 254747
rect 12821 254947 13021 254957
rect 12821 254737 13021 254747
rect 13241 254947 13441 254957
rect 13241 254737 13441 254747
rect 13661 254947 13861 254957
rect 13661 254737 13861 254747
rect 14081 254947 14281 254957
rect 14081 254737 14281 254747
rect 14501 254947 14701 254957
rect 14501 254737 14701 254747
rect 14921 254947 15121 254957
rect 14921 254737 15121 254747
rect 15341 254947 15541 254957
rect 15341 254737 15541 254747
rect 15761 254947 15961 254957
rect 15761 254737 15961 254747
rect 16181 254947 16381 254957
rect 16181 254737 16381 254747
rect 16601 254947 16801 254957
rect 16601 254737 16801 254747
rect 17021 254947 17221 254957
rect 17021 254737 17221 254747
rect 17441 254947 17641 254957
rect 17441 254737 17641 254747
rect 17861 254947 18061 254957
rect 17861 254737 18061 254747
rect 18281 254947 18481 254957
rect 18281 254737 18481 254747
rect 18701 254947 18901 254957
rect 18701 254737 18901 254747
rect 19121 254947 19321 254957
rect 19121 254737 19321 254747
rect 19541 254947 19741 254957
rect 19541 254737 19741 254747
rect 19961 254947 20161 254957
rect 19961 254737 20161 254747
rect 20381 254947 20581 254957
rect 20381 254737 20581 254747
rect 20801 254947 21001 254957
rect 20801 254737 21001 254747
rect 21221 254947 21421 254957
rect 21221 254737 21421 254747
rect 21641 254947 21841 254957
rect 21641 254737 21841 254747
rect 22061 254947 22261 254957
rect 22061 254737 22261 254747
rect 22481 254947 22681 254957
rect 22481 254737 22681 254747
rect 22901 254947 23101 254957
rect 22901 254737 23101 254747
rect 23321 254947 23521 254957
rect 23321 254737 23521 254747
rect 23741 254947 23941 254957
rect 23741 254737 23941 254747
rect 24161 254947 24361 254957
rect 24161 254737 24361 254747
rect 24581 254947 24781 254957
rect 24581 254737 24781 254747
rect 25001 254947 25201 254957
rect 25001 254737 25201 254747
rect 25421 254947 25621 254957
rect 25421 254737 25621 254747
rect 25841 254947 26041 254957
rect 25841 254737 26041 254747
rect 26261 254947 26461 254957
rect 26261 254737 26461 254747
rect 26681 254947 26881 254957
rect 26681 254737 26881 254747
rect 27101 254947 27301 254957
rect 27101 254737 27301 254747
rect -4075 254489 -4015 254499
rect -4075 253713 -4069 254489
rect -4075 253453 -4015 253713
rect -4075 252677 -4069 253453
rect -4075 252417 -4015 252677
rect -4075 251641 -4069 252417
rect -4075 251381 -4015 251641
rect -4075 250605 -4069 251381
rect -4075 250345 -4015 250605
rect -4075 249569 -4069 250345
rect -4075 249180 -4015 249569
rect -4075 248144 -4015 248404
rect -4075 247108 -4015 247368
rect -4075 246072 -4015 246332
rect -4075 245036 -4015 245296
rect -4075 244075 -4015 244260
rect -3963 254489 -3795 254737
rect -3963 253713 -3953 254489
rect -3805 253713 -3795 254489
rect -3963 253453 -3795 253713
rect -3963 252677 -3953 253453
rect -3805 252677 -3795 253453
rect -3963 252417 -3795 252677
rect -3963 251641 -3953 252417
rect -3805 251641 -3795 252417
rect -3963 251381 -3795 251641
rect -3963 250605 -3953 251381
rect -3805 250605 -3795 251381
rect -3963 250345 -3795 250605
rect -3963 249569 -3953 250345
rect -3805 249569 -3795 250345
rect -3963 249180 -3795 249569
rect -3963 248404 -3953 249180
rect -3805 248404 -3795 249180
rect -3963 248144 -3795 248404
rect -3963 247368 -3953 248144
rect -3805 247368 -3795 248144
rect -3963 247108 -3795 247368
rect -3963 246332 -3953 247108
rect -3805 246332 -3795 247108
rect -3963 246072 -3795 246332
rect -3963 245296 -3953 246072
rect -3805 245296 -3795 246072
rect -3963 245036 -3795 245296
rect -3963 244260 -3953 245036
rect -3805 244260 -3795 245036
rect -3963 244248 -3795 244260
rect -3753 254489 -3585 254501
rect -3753 253713 -3743 254489
rect -3595 253713 -3585 254489
rect -3753 253453 -3585 253713
rect -3753 252677 -3743 253453
rect -3595 252677 -3585 253453
rect -3753 252417 -3585 252677
rect -3753 251641 -3743 252417
rect -3595 251641 -3585 252417
rect -3753 251381 -3585 251641
rect -3753 250605 -3743 251381
rect -3595 250605 -3585 251381
rect -3753 250345 -3585 250605
rect -3753 249569 -3743 250345
rect -3595 249569 -3585 250345
rect -3753 249180 -3585 249569
rect -3753 248404 -3743 249180
rect -3595 248404 -3585 249180
rect -3753 248144 -3585 248404
rect -3753 247368 -3743 248144
rect -3595 247368 -3585 248144
rect -3753 247108 -3585 247368
rect -3753 246332 -3743 247108
rect -3595 246332 -3585 247108
rect -3753 246072 -3585 246332
rect -3753 245296 -3743 246072
rect -3595 245296 -3585 246072
rect -3753 245036 -3585 245296
rect -3753 244260 -3743 245036
rect -3595 244260 -3585 245036
rect -3753 244075 -3585 244260
rect -3543 254490 -3375 254737
rect -3543 253713 -3533 254490
rect -3385 253713 -3375 254490
rect -3543 253454 -3375 253713
rect -3543 252677 -3533 253454
rect -3385 252677 -3375 253454
rect -3543 252418 -3375 252677
rect -3543 251641 -3533 252418
rect -3385 251641 -3375 252418
rect -3543 251382 -3375 251641
rect -3543 250605 -3533 251382
rect -3385 250605 -3375 251382
rect -3543 250346 -3375 250605
rect -3543 249569 -3533 250346
rect -3385 249569 -3375 250346
rect -3543 249181 -3375 249569
rect -3543 248404 -3533 249181
rect -3385 248404 -3375 249181
rect -3543 248145 -3375 248404
rect -3543 247368 -3533 248145
rect -3385 247368 -3375 248145
rect -3543 247109 -3375 247368
rect -3543 246332 -3533 247109
rect -3385 246332 -3375 247109
rect -3543 246073 -3375 246332
rect -3543 245296 -3533 246073
rect -3385 245296 -3375 246073
rect -3543 245037 -3375 245296
rect -3543 244260 -3533 245037
rect -3385 244260 -3375 245037
rect -3543 244248 -3375 244260
rect -3333 254490 -3165 254501
rect -3333 253713 -3323 254490
rect -3175 253713 -3165 254490
rect -3333 253454 -3165 253713
rect -3333 252677 -3323 253454
rect -3175 252677 -3165 253454
rect -3333 252418 -3165 252677
rect -3333 251641 -3323 252418
rect -3175 251641 -3165 252418
rect -3333 251382 -3165 251641
rect -3333 250605 -3323 251382
rect -3175 250605 -3165 251382
rect -3333 250346 -3165 250605
rect -3333 249569 -3323 250346
rect -3175 249569 -3165 250346
rect -3333 249181 -3165 249569
rect -3333 248404 -3323 249181
rect -3175 248404 -3165 249181
rect -3333 248145 -3165 248404
rect -3333 247368 -3323 248145
rect -3175 247368 -3165 248145
rect -3333 247109 -3165 247368
rect -3333 246332 -3323 247109
rect -3175 246332 -3165 247109
rect -3333 246073 -3165 246332
rect -3333 245296 -3323 246073
rect -3175 245296 -3165 246073
rect -3333 245037 -3165 245296
rect -3333 244260 -3323 245037
rect -3175 244260 -3165 245037
rect -3333 244075 -3165 244260
rect -3123 254490 -2955 254737
rect -3123 253713 -3113 254490
rect -2965 253713 -2955 254490
rect -3123 253454 -2955 253713
rect -3123 252677 -3113 253454
rect -2965 252677 -2955 253454
rect -3123 252418 -2955 252677
rect -3123 251641 -3113 252418
rect -2965 251641 -2955 252418
rect -3123 251382 -2955 251641
rect -3123 250605 -3113 251382
rect -2965 250605 -2955 251382
rect -3123 250346 -2955 250605
rect -3123 249569 -3113 250346
rect -2965 249569 -2955 250346
rect -3123 249181 -2955 249569
rect -3123 248404 -3113 249181
rect -2965 248404 -2955 249181
rect -3123 248145 -2955 248404
rect -3123 247368 -3113 248145
rect -2965 247368 -2955 248145
rect -3123 247109 -2955 247368
rect -3123 246332 -3113 247109
rect -2965 246332 -2955 247109
rect -3123 246073 -2955 246332
rect -3123 245296 -3113 246073
rect -2965 245296 -2955 246073
rect -3123 245037 -2955 245296
rect -3123 244260 -3113 245037
rect -2965 244260 -2955 245037
rect -3123 244248 -2955 244260
rect -2913 254490 -2745 254501
rect -2913 253713 -2903 254490
rect -2755 253713 -2745 254490
rect -2913 253454 -2745 253713
rect -2913 252677 -2903 253454
rect -2755 252677 -2745 253454
rect -2913 252418 -2745 252677
rect -2913 251641 -2903 252418
rect -2755 251641 -2745 252418
rect -2913 251382 -2745 251641
rect -2913 250605 -2903 251382
rect -2755 250605 -2745 251382
rect -2913 250346 -2745 250605
rect -2913 249569 -2903 250346
rect -2755 249569 -2745 250346
rect -2913 249181 -2745 249569
rect -2913 248404 -2903 249181
rect -2755 248404 -2745 249181
rect -2913 248145 -2745 248404
rect -2913 247368 -2903 248145
rect -2755 247368 -2745 248145
rect -2913 247109 -2745 247368
rect -2913 246332 -2903 247109
rect -2755 246332 -2745 247109
rect -2913 246073 -2745 246332
rect -2913 245296 -2903 246073
rect -2755 245296 -2745 246073
rect -2913 245037 -2745 245296
rect -2913 244260 -2903 245037
rect -2755 244260 -2745 245037
rect -2913 244075 -2745 244260
rect -2703 254490 -2535 254737
rect -2703 253713 -2693 254490
rect -2545 253713 -2535 254490
rect -2703 253454 -2535 253713
rect -2703 252677 -2693 253454
rect -2545 252677 -2535 253454
rect -2703 252418 -2535 252677
rect -2703 251641 -2693 252418
rect -2545 251641 -2535 252418
rect -2703 251382 -2535 251641
rect -2703 250605 -2693 251382
rect -2545 250605 -2535 251382
rect -2703 250346 -2535 250605
rect -2703 249569 -2693 250346
rect -2545 249569 -2535 250346
rect -2703 249181 -2535 249569
rect -2703 248404 -2693 249181
rect -2545 248404 -2535 249181
rect -2703 248145 -2535 248404
rect -2703 247368 -2693 248145
rect -2545 247368 -2535 248145
rect -2703 247109 -2535 247368
rect -2703 246332 -2693 247109
rect -2545 246332 -2535 247109
rect -2703 246073 -2535 246332
rect -2703 245296 -2693 246073
rect -2545 245296 -2535 246073
rect -2703 245037 -2535 245296
rect -2703 244260 -2693 245037
rect -2545 244260 -2535 245037
rect -2703 244248 -2535 244260
rect -2493 254490 -2325 254501
rect -2493 253713 -2483 254490
rect -2335 253713 -2325 254490
rect -2493 253454 -2325 253713
rect -2493 252677 -2483 253454
rect -2335 252677 -2325 253454
rect -2493 252418 -2325 252677
rect -2493 251641 -2483 252418
rect -2335 251641 -2325 252418
rect -2493 251382 -2325 251641
rect -2493 250605 -2483 251382
rect -2335 250605 -2325 251382
rect -2493 250346 -2325 250605
rect -2493 249569 -2483 250346
rect -2335 249569 -2325 250346
rect -2493 249181 -2325 249569
rect -2493 248404 -2483 249181
rect -2335 248404 -2325 249181
rect -2493 248145 -2325 248404
rect -2493 247368 -2483 248145
rect -2335 247368 -2325 248145
rect -2493 247109 -2325 247368
rect -2493 246332 -2483 247109
rect -2335 246332 -2325 247109
rect -2493 246073 -2325 246332
rect -2493 245296 -2483 246073
rect -2335 245296 -2325 246073
rect -2493 245037 -2325 245296
rect -2493 244260 -2483 245037
rect -2335 244260 -2325 245037
rect -2493 244075 -2325 244260
rect -2283 254490 -2115 254737
rect -2283 253713 -2273 254490
rect -2125 253713 -2115 254490
rect -2283 253454 -2115 253713
rect -2283 252677 -2273 253454
rect -2125 252677 -2115 253454
rect -2283 252418 -2115 252677
rect -2283 251641 -2273 252418
rect -2125 251641 -2115 252418
rect -2283 251382 -2115 251641
rect -2283 250605 -2273 251382
rect -2125 250605 -2115 251382
rect -2283 250346 -2115 250605
rect -2283 249569 -2273 250346
rect -2125 249569 -2115 250346
rect -2283 249181 -2115 249569
rect -2283 248404 -2273 249181
rect -2125 248404 -2115 249181
rect -2283 248145 -2115 248404
rect -2283 247368 -2273 248145
rect -2125 247368 -2115 248145
rect -2283 247109 -2115 247368
rect -2283 246332 -2273 247109
rect -2125 246332 -2115 247109
rect -2283 246073 -2115 246332
rect -2283 245296 -2273 246073
rect -2125 245296 -2115 246073
rect -2283 245037 -2115 245296
rect -2283 244260 -2273 245037
rect -2125 244260 -2115 245037
rect -2283 244248 -2115 244260
rect -2073 254490 -1905 254501
rect -2073 253713 -2063 254490
rect -1915 253713 -1905 254490
rect -2073 253454 -1905 253713
rect -2073 252677 -2063 253454
rect -1915 252677 -1905 253454
rect -2073 252418 -1905 252677
rect -2073 251641 -2063 252418
rect -1915 251641 -1905 252418
rect -2073 251382 -1905 251641
rect -2073 250605 -2063 251382
rect -1915 250605 -1905 251382
rect -2073 250346 -1905 250605
rect -2073 249569 -2063 250346
rect -1915 249569 -1905 250346
rect -2073 249181 -1905 249569
rect -2073 248404 -2063 249181
rect -1915 248404 -1905 249181
rect -2073 248145 -1905 248404
rect -2073 247368 -2063 248145
rect -1915 247368 -1905 248145
rect -2073 247109 -1905 247368
rect -2073 246332 -2063 247109
rect -1915 246332 -1905 247109
rect -2073 246073 -1905 246332
rect -2073 245296 -2063 246073
rect -1915 245296 -1905 246073
rect -2073 245037 -1905 245296
rect -2073 244260 -2063 245037
rect -1915 244260 -1905 245037
rect -2073 244075 -1905 244260
rect -1863 254490 -1695 254737
rect -1863 253713 -1853 254490
rect -1705 253713 -1695 254490
rect -1863 253454 -1695 253713
rect -1863 252677 -1853 253454
rect -1705 252677 -1695 253454
rect -1863 252418 -1695 252677
rect -1863 251641 -1853 252418
rect -1705 251641 -1695 252418
rect -1863 251382 -1695 251641
rect -1863 250605 -1853 251382
rect -1705 250605 -1695 251382
rect -1863 250346 -1695 250605
rect -1863 249569 -1853 250346
rect -1705 249569 -1695 250346
rect -1863 249181 -1695 249569
rect -1863 248404 -1853 249181
rect -1705 248404 -1695 249181
rect -1863 248145 -1695 248404
rect -1863 247368 -1853 248145
rect -1705 247368 -1695 248145
rect -1863 247109 -1695 247368
rect -1863 246332 -1853 247109
rect -1705 246332 -1695 247109
rect -1863 246073 -1695 246332
rect -1863 245296 -1853 246073
rect -1705 245296 -1695 246073
rect -1863 245037 -1695 245296
rect -1863 244260 -1853 245037
rect -1705 244260 -1695 245037
rect -1863 244248 -1695 244260
rect -1653 254490 -1485 254501
rect -1653 253713 -1643 254490
rect -1495 253713 -1485 254490
rect -1653 253454 -1485 253713
rect -1653 252677 -1643 253454
rect -1495 252677 -1485 253454
rect -1653 252418 -1485 252677
rect -1653 251641 -1643 252418
rect -1495 251641 -1485 252418
rect -1653 251382 -1485 251641
rect -1653 250605 -1643 251382
rect -1495 250605 -1485 251382
rect -1653 250346 -1485 250605
rect -1653 249569 -1643 250346
rect -1495 249569 -1485 250346
rect -1653 249181 -1485 249569
rect -1653 248404 -1643 249181
rect -1495 248404 -1485 249181
rect -1653 248145 -1485 248404
rect -1653 247368 -1643 248145
rect -1495 247368 -1485 248145
rect -1653 247109 -1485 247368
rect -1653 246332 -1643 247109
rect -1495 246332 -1485 247109
rect -1653 246073 -1485 246332
rect -1653 245296 -1643 246073
rect -1495 245296 -1485 246073
rect -1653 245037 -1485 245296
rect -1653 244260 -1643 245037
rect -1495 244260 -1485 245037
rect -1653 244075 -1485 244260
rect -1443 254490 -1275 254737
rect -1443 253713 -1433 254490
rect -1285 253713 -1275 254490
rect -1443 253454 -1275 253713
rect -1443 252677 -1433 253454
rect -1285 252677 -1275 253454
rect -1443 252418 -1275 252677
rect -1443 251641 -1433 252418
rect -1285 251641 -1275 252418
rect -1443 251382 -1275 251641
rect -1443 250605 -1433 251382
rect -1285 250605 -1275 251382
rect -1443 250346 -1275 250605
rect -1443 249569 -1433 250346
rect -1285 249569 -1275 250346
rect -1443 249181 -1275 249569
rect -1443 248404 -1433 249181
rect -1285 248404 -1275 249181
rect -1443 248145 -1275 248404
rect -1443 247368 -1433 248145
rect -1285 247368 -1275 248145
rect -1443 247109 -1275 247368
rect -1443 246332 -1433 247109
rect -1285 246332 -1275 247109
rect -1443 246073 -1275 246332
rect -1443 245296 -1433 246073
rect -1285 245296 -1275 246073
rect -1443 245037 -1275 245296
rect -1443 244260 -1433 245037
rect -1285 244260 -1275 245037
rect -1443 244248 -1275 244260
rect -1233 254490 -1065 254501
rect -1233 253713 -1223 254490
rect -1075 253713 -1065 254490
rect -1233 253454 -1065 253713
rect -1233 252677 -1223 253454
rect -1075 252677 -1065 253454
rect -1233 252418 -1065 252677
rect -1233 251641 -1223 252418
rect -1075 251641 -1065 252418
rect -1233 251382 -1065 251641
rect -1233 250605 -1223 251382
rect -1075 250605 -1065 251382
rect -1233 250346 -1065 250605
rect -1233 249569 -1223 250346
rect -1075 249569 -1065 250346
rect -1233 249181 -1065 249569
rect -1233 248404 -1223 249181
rect -1075 248404 -1065 249181
rect -1233 248145 -1065 248404
rect -1233 247368 -1223 248145
rect -1075 247368 -1065 248145
rect -1233 247109 -1065 247368
rect -1233 246332 -1223 247109
rect -1075 246332 -1065 247109
rect -1233 246073 -1065 246332
rect -1233 245296 -1223 246073
rect -1075 245296 -1065 246073
rect -1233 245037 -1065 245296
rect -1233 244260 -1223 245037
rect -1075 244260 -1065 245037
rect -1233 244075 -1065 244260
rect -1023 254490 -855 254737
rect -1023 253713 -1013 254490
rect -865 253713 -855 254490
rect -1023 253454 -855 253713
rect -1023 252677 -1013 253454
rect -865 252677 -855 253454
rect -1023 252418 -855 252677
rect -1023 251641 -1013 252418
rect -865 251641 -855 252418
rect -1023 251382 -855 251641
rect -1023 250605 -1013 251382
rect -865 250605 -855 251382
rect -1023 250346 -855 250605
rect -1023 249569 -1013 250346
rect -865 249569 -855 250346
rect -1023 249181 -855 249569
rect -1023 248404 -1013 249181
rect -865 248404 -855 249181
rect -1023 248145 -855 248404
rect -1023 247368 -1013 248145
rect -865 247368 -855 248145
rect -1023 247109 -855 247368
rect -1023 246332 -1013 247109
rect -865 246332 -855 247109
rect -1023 246073 -855 246332
rect -1023 245296 -1013 246073
rect -865 245296 -855 246073
rect -1023 245037 -855 245296
rect -1023 244260 -1013 245037
rect -865 244260 -855 245037
rect -1023 244248 -855 244260
rect -813 254490 -645 254501
rect -813 253713 -803 254490
rect -655 253713 -645 254490
rect -813 253454 -645 253713
rect -813 252677 -803 253454
rect -655 252677 -645 253454
rect -813 252418 -645 252677
rect -813 251641 -803 252418
rect -655 251641 -645 252418
rect -813 251382 -645 251641
rect -813 250605 -803 251382
rect -655 250605 -645 251382
rect -813 250346 -645 250605
rect -813 249569 -803 250346
rect -655 249569 -645 250346
rect -813 249181 -645 249569
rect -813 248404 -803 249181
rect -655 248404 -645 249181
rect -813 248145 -645 248404
rect -813 247368 -803 248145
rect -655 247368 -645 248145
rect -813 247109 -645 247368
rect -813 246332 -803 247109
rect -655 246332 -645 247109
rect -813 246073 -645 246332
rect -813 245296 -803 246073
rect -655 245296 -645 246073
rect -813 245037 -645 245296
rect -813 244260 -803 245037
rect -655 244260 -645 245037
rect -813 244075 -645 244260
rect -603 254490 -435 254737
rect -603 253713 -593 254490
rect -445 253713 -435 254490
rect -603 253454 -435 253713
rect -603 252677 -593 253454
rect -445 252677 -435 253454
rect -603 252418 -435 252677
rect -603 251641 -593 252418
rect -445 251641 -435 252418
rect -603 251382 -435 251641
rect -603 250605 -593 251382
rect -445 250605 -435 251382
rect -603 250346 -435 250605
rect -603 249569 -593 250346
rect -445 249569 -435 250346
rect -603 249181 -435 249569
rect -603 248404 -593 249181
rect -445 248404 -435 249181
rect -603 248145 -435 248404
rect -603 247368 -593 248145
rect -445 247368 -435 248145
rect -603 247109 -435 247368
rect -603 246332 -593 247109
rect -445 246332 -435 247109
rect -603 246073 -435 246332
rect -603 245296 -593 246073
rect -445 245296 -435 246073
rect -603 245037 -435 245296
rect -603 244260 -593 245037
rect -445 244260 -435 245037
rect -603 244248 -435 244260
rect -393 254490 -225 254501
rect -393 253713 -383 254490
rect -235 253713 -225 254490
rect -393 253454 -225 253713
rect -393 252677 -383 253454
rect -235 252677 -225 253454
rect -393 252418 -225 252677
rect -393 251641 -383 252418
rect -235 251641 -225 252418
rect -393 251382 -225 251641
rect -393 250605 -383 251382
rect -235 250605 -225 251382
rect -393 250346 -225 250605
rect -393 249569 -383 250346
rect -235 249569 -225 250346
rect -393 249181 -225 249569
rect -393 248404 -383 249181
rect -235 248404 -225 249181
rect -393 248145 -225 248404
rect -393 247368 -383 248145
rect -235 247368 -225 248145
rect -393 247109 -225 247368
rect -393 246332 -383 247109
rect -235 246332 -225 247109
rect -393 246073 -225 246332
rect -393 245296 -383 246073
rect -235 245296 -225 246073
rect -393 245037 -225 245296
rect -393 244260 -383 245037
rect -235 244260 -225 245037
rect -393 244075 -225 244260
rect -183 254490 -15 254737
rect -183 253713 -173 254490
rect -25 253713 -15 254490
rect -183 253454 -15 253713
rect -183 252677 -173 253454
rect -25 252677 -15 253454
rect -183 252418 -15 252677
rect -183 251641 -173 252418
rect -25 251641 -15 252418
rect -183 251382 -15 251641
rect -183 250605 -173 251382
rect -25 250605 -15 251382
rect -183 250346 -15 250605
rect -183 249569 -173 250346
rect -25 249569 -15 250346
rect -183 249181 -15 249569
rect -183 248404 -173 249181
rect -25 248404 -15 249181
rect -183 248145 -15 248404
rect -183 247368 -173 248145
rect -25 247368 -15 248145
rect -183 247109 -15 247368
rect -183 246332 -173 247109
rect -25 246332 -15 247109
rect -183 246073 -15 246332
rect -183 245296 -173 246073
rect -25 245296 -15 246073
rect -183 245037 -15 245296
rect -183 244260 -173 245037
rect -25 244260 -15 245037
rect -183 244248 -15 244260
rect 27 254490 195 254501
rect 27 253713 37 254490
rect 185 253713 195 254490
rect 27 253454 195 253713
rect 27 252677 37 253454
rect 185 252677 195 253454
rect 27 252418 195 252677
rect 27 251641 37 252418
rect 185 251641 195 252418
rect 27 251382 195 251641
rect 27 250605 37 251382
rect 185 250605 195 251382
rect 27 250346 195 250605
rect 27 249569 37 250346
rect 185 249569 195 250346
rect 27 249181 195 249569
rect 27 248404 37 249181
rect 185 248404 195 249181
rect 27 248145 195 248404
rect 27 247368 37 248145
rect 185 247368 195 248145
rect 27 247109 195 247368
rect 27 246332 37 247109
rect 185 246332 195 247109
rect 27 246073 195 246332
rect 27 245296 37 246073
rect 185 245296 195 246073
rect 27 245037 195 245296
rect 27 244260 37 245037
rect 185 244260 195 245037
rect 27 244075 195 244260
rect 237 254490 405 254737
rect 237 253713 247 254490
rect 395 253713 405 254490
rect 237 253454 405 253713
rect 237 252677 247 253454
rect 395 252677 405 253454
rect 237 252418 405 252677
rect 237 251641 247 252418
rect 395 251641 405 252418
rect 237 251382 405 251641
rect 237 250605 247 251382
rect 395 250605 405 251382
rect 237 250346 405 250605
rect 237 249569 247 250346
rect 395 249569 405 250346
rect 237 249181 405 249569
rect 237 248404 247 249181
rect 395 248404 405 249181
rect 237 248145 405 248404
rect 237 247368 247 248145
rect 395 247368 405 248145
rect 237 247109 405 247368
rect 237 246332 247 247109
rect 395 246332 405 247109
rect 237 246073 405 246332
rect 237 245296 247 246073
rect 395 245296 405 246073
rect 237 245037 405 245296
rect 237 244260 247 245037
rect 395 244260 405 245037
rect 237 244248 405 244260
rect 447 254490 615 254501
rect 447 253713 457 254490
rect 605 253713 615 254490
rect 447 253454 615 253713
rect 447 252677 457 253454
rect 605 252677 615 253454
rect 447 252418 615 252677
rect 447 251641 457 252418
rect 605 251641 615 252418
rect 447 251382 615 251641
rect 447 250605 457 251382
rect 605 250605 615 251382
rect 447 250346 615 250605
rect 447 249569 457 250346
rect 605 249569 615 250346
rect 447 249181 615 249569
rect 447 248404 457 249181
rect 605 248404 615 249181
rect 447 248145 615 248404
rect 447 247368 457 248145
rect 605 247368 615 248145
rect 447 247109 615 247368
rect 447 246332 457 247109
rect 605 246332 615 247109
rect 447 246073 615 246332
rect 447 245296 457 246073
rect 605 245296 615 246073
rect 447 245037 615 245296
rect 447 244260 457 245037
rect 605 244260 615 245037
rect 447 244075 615 244260
rect 657 254490 825 254737
rect 657 253713 667 254490
rect 815 253713 825 254490
rect 657 253454 825 253713
rect 657 252677 667 253454
rect 815 252677 825 253454
rect 657 252418 825 252677
rect 657 251641 667 252418
rect 815 251641 825 252418
rect 657 251382 825 251641
rect 657 250605 667 251382
rect 815 250605 825 251382
rect 657 250346 825 250605
rect 657 249569 667 250346
rect 815 249569 825 250346
rect 657 249181 825 249569
rect 657 248404 667 249181
rect 815 248404 825 249181
rect 657 248145 825 248404
rect 657 247368 667 248145
rect 815 247368 825 248145
rect 657 247109 825 247368
rect 657 246332 667 247109
rect 815 246332 825 247109
rect 657 246073 825 246332
rect 657 245296 667 246073
rect 815 245296 825 246073
rect 657 245037 825 245296
rect 657 244260 667 245037
rect 815 244260 825 245037
rect 657 244248 825 244260
rect 867 254490 1035 254501
rect 867 253713 877 254490
rect 1025 253713 1035 254490
rect 867 253454 1035 253713
rect 867 252677 877 253454
rect 1025 252677 1035 253454
rect 867 252418 1035 252677
rect 867 251641 877 252418
rect 1025 251641 1035 252418
rect 867 251382 1035 251641
rect 867 250605 877 251382
rect 1025 250605 1035 251382
rect 867 250346 1035 250605
rect 867 249569 877 250346
rect 1025 249569 1035 250346
rect 867 249181 1035 249569
rect 867 248404 877 249181
rect 1025 248404 1035 249181
rect 867 248145 1035 248404
rect 867 247368 877 248145
rect 1025 247368 1035 248145
rect 867 247109 1035 247368
rect 867 246332 877 247109
rect 1025 246332 1035 247109
rect 867 246073 1035 246332
rect 867 245296 877 246073
rect 1025 245296 1035 246073
rect 867 245037 1035 245296
rect 867 244260 877 245037
rect 1025 244260 1035 245037
rect 867 244075 1035 244260
rect 1077 254490 1245 254737
rect 1077 253713 1087 254490
rect 1235 253713 1245 254490
rect 1077 253454 1245 253713
rect 1077 252677 1087 253454
rect 1235 252677 1245 253454
rect 1077 252418 1245 252677
rect 1077 251641 1087 252418
rect 1235 251641 1245 252418
rect 1077 251382 1245 251641
rect 1077 250605 1087 251382
rect 1235 250605 1245 251382
rect 1077 250346 1245 250605
rect 1077 249569 1087 250346
rect 1235 249569 1245 250346
rect 1077 249181 1245 249569
rect 1077 248404 1087 249181
rect 1235 248404 1245 249181
rect 1077 248145 1245 248404
rect 1077 247368 1087 248145
rect 1235 247368 1245 248145
rect 1077 247109 1245 247368
rect 1077 246332 1087 247109
rect 1235 246332 1245 247109
rect 1077 246073 1245 246332
rect 1077 245296 1087 246073
rect 1235 245296 1245 246073
rect 1077 245037 1245 245296
rect 1077 244260 1087 245037
rect 1235 244260 1245 245037
rect 1077 244248 1245 244260
rect 1287 254490 1455 254501
rect 1287 253713 1297 254490
rect 1445 253713 1455 254490
rect 1287 253454 1455 253713
rect 1287 252677 1297 253454
rect 1445 252677 1455 253454
rect 1287 252418 1455 252677
rect 1287 251641 1297 252418
rect 1445 251641 1455 252418
rect 1287 251382 1455 251641
rect 1287 250605 1297 251382
rect 1445 250605 1455 251382
rect 1287 250346 1455 250605
rect 1287 249569 1297 250346
rect 1445 249569 1455 250346
rect 1287 249181 1455 249569
rect 1287 248404 1297 249181
rect 1445 248404 1455 249181
rect 1287 248145 1455 248404
rect 1287 247368 1297 248145
rect 1445 247368 1455 248145
rect 1287 247109 1455 247368
rect 1287 246332 1297 247109
rect 1445 246332 1455 247109
rect 1287 246073 1455 246332
rect 1287 245296 1297 246073
rect 1445 245296 1455 246073
rect 1287 245037 1455 245296
rect 1287 244260 1297 245037
rect 1445 244260 1455 245037
rect 1287 244075 1455 244260
rect 1497 254490 1665 254737
rect 1497 253713 1507 254490
rect 1655 253713 1665 254490
rect 1497 253454 1665 253713
rect 1497 252677 1507 253454
rect 1655 252677 1665 253454
rect 1497 252418 1665 252677
rect 1497 251641 1507 252418
rect 1655 251641 1665 252418
rect 1497 251382 1665 251641
rect 1497 250605 1507 251382
rect 1655 250605 1665 251382
rect 1497 250346 1665 250605
rect 1497 249569 1507 250346
rect 1655 249569 1665 250346
rect 1497 249181 1665 249569
rect 1497 248404 1507 249181
rect 1655 248404 1665 249181
rect 1497 248145 1665 248404
rect 1497 247368 1507 248145
rect 1655 247368 1665 248145
rect 1497 247109 1665 247368
rect 1497 246332 1507 247109
rect 1655 246332 1665 247109
rect 1497 246073 1665 246332
rect 1497 245296 1507 246073
rect 1655 245296 1665 246073
rect 1497 245037 1665 245296
rect 1497 244260 1507 245037
rect 1655 244260 1665 245037
rect 1497 244248 1665 244260
rect 1707 254490 1875 254501
rect 1707 253713 1717 254490
rect 1865 253713 1875 254490
rect 1707 253454 1875 253713
rect 1707 252677 1717 253454
rect 1865 252677 1875 253454
rect 1707 252418 1875 252677
rect 1707 251641 1717 252418
rect 1865 251641 1875 252418
rect 1707 251382 1875 251641
rect 1707 250605 1717 251382
rect 1865 250605 1875 251382
rect 1707 250346 1875 250605
rect 1707 249569 1717 250346
rect 1865 249569 1875 250346
rect 1707 249181 1875 249569
rect 1707 248404 1717 249181
rect 1865 248404 1875 249181
rect 1707 248145 1875 248404
rect 1707 247368 1717 248145
rect 1865 247368 1875 248145
rect 1707 247109 1875 247368
rect 1707 246332 1717 247109
rect 1865 246332 1875 247109
rect 1707 246073 1875 246332
rect 1707 245296 1717 246073
rect 1865 245296 1875 246073
rect 1707 245037 1875 245296
rect 1707 244260 1717 245037
rect 1865 244260 1875 245037
rect 1707 244075 1875 244260
rect 1917 254490 2085 254737
rect 1917 253713 1927 254490
rect 2075 253713 2085 254490
rect 1917 253454 2085 253713
rect 1917 252677 1927 253454
rect 2075 252677 2085 253454
rect 1917 252418 2085 252677
rect 1917 251641 1927 252418
rect 2075 251641 2085 252418
rect 1917 251382 2085 251641
rect 1917 250605 1927 251382
rect 2075 250605 2085 251382
rect 1917 250346 2085 250605
rect 1917 249569 1927 250346
rect 2075 249569 2085 250346
rect 1917 249181 2085 249569
rect 1917 248404 1927 249181
rect 2075 248404 2085 249181
rect 1917 248145 2085 248404
rect 1917 247368 1927 248145
rect 2075 247368 2085 248145
rect 1917 247109 2085 247368
rect 1917 246332 1927 247109
rect 2075 246332 2085 247109
rect 1917 246073 2085 246332
rect 1917 245296 1927 246073
rect 2075 245296 2085 246073
rect 1917 245037 2085 245296
rect 1917 244260 1927 245037
rect 2075 244260 2085 245037
rect 1917 244248 2085 244260
rect 2127 254490 2295 254501
rect 2127 253713 2137 254490
rect 2285 253713 2295 254490
rect 2127 253454 2295 253713
rect 2127 252677 2137 253454
rect 2285 252677 2295 253454
rect 2127 252418 2295 252677
rect 2127 251641 2137 252418
rect 2285 251641 2295 252418
rect 2127 251382 2295 251641
rect 2127 250605 2137 251382
rect 2285 250605 2295 251382
rect 2127 250346 2295 250605
rect 2127 249569 2137 250346
rect 2285 249569 2295 250346
rect 2127 249181 2295 249569
rect 2127 248404 2137 249181
rect 2285 248404 2295 249181
rect 2127 248145 2295 248404
rect 2127 247368 2137 248145
rect 2285 247368 2295 248145
rect 2127 247109 2295 247368
rect 2127 246332 2137 247109
rect 2285 246332 2295 247109
rect 2127 246073 2295 246332
rect 2127 245296 2137 246073
rect 2285 245296 2295 246073
rect 2127 245037 2295 245296
rect 2127 244260 2137 245037
rect 2285 244260 2295 245037
rect 2127 244075 2295 244260
rect 2337 254490 2505 254737
rect 2337 253713 2347 254490
rect 2495 253713 2505 254490
rect 2337 253454 2505 253713
rect 2337 252677 2347 253454
rect 2495 252677 2505 253454
rect 2337 252418 2505 252677
rect 2337 251641 2347 252418
rect 2495 251641 2505 252418
rect 2337 251382 2505 251641
rect 2337 250605 2347 251382
rect 2495 250605 2505 251382
rect 2337 250346 2505 250605
rect 2337 249569 2347 250346
rect 2495 249569 2505 250346
rect 2337 249181 2505 249569
rect 2337 248404 2347 249181
rect 2495 248404 2505 249181
rect 2337 248145 2505 248404
rect 2337 247368 2347 248145
rect 2495 247368 2505 248145
rect 2337 247109 2505 247368
rect 2337 246332 2347 247109
rect 2495 246332 2505 247109
rect 2337 246073 2505 246332
rect 2337 245296 2347 246073
rect 2495 245296 2505 246073
rect 2337 245037 2505 245296
rect 2337 244260 2347 245037
rect 2495 244260 2505 245037
rect 2337 244248 2505 244260
rect 2547 254490 2715 254501
rect 2547 253713 2557 254490
rect 2705 253713 2715 254490
rect 2547 253454 2715 253713
rect 2547 252677 2557 253454
rect 2705 252677 2715 253454
rect 2547 252418 2715 252677
rect 2547 251641 2557 252418
rect 2705 251641 2715 252418
rect 2547 251382 2715 251641
rect 2547 250605 2557 251382
rect 2705 250605 2715 251382
rect 2547 250346 2715 250605
rect 2547 249569 2557 250346
rect 2705 249569 2715 250346
rect 2547 249181 2715 249569
rect 2547 248404 2557 249181
rect 2705 248404 2715 249181
rect 2547 248145 2715 248404
rect 2547 247368 2557 248145
rect 2705 247368 2715 248145
rect 2547 247109 2715 247368
rect 2547 246332 2557 247109
rect 2705 246332 2715 247109
rect 2547 246073 2715 246332
rect 2547 245296 2557 246073
rect 2705 245296 2715 246073
rect 2547 245037 2715 245296
rect 2547 244260 2557 245037
rect 2705 244260 2715 245037
rect 2547 244075 2715 244260
rect 2757 254490 2925 254737
rect 2757 253713 2767 254490
rect 2915 253713 2925 254490
rect 2757 253454 2925 253713
rect 2757 252677 2767 253454
rect 2915 252677 2925 253454
rect 2757 252418 2925 252677
rect 2757 251641 2767 252418
rect 2915 251641 2925 252418
rect 2757 251382 2925 251641
rect 2757 250605 2767 251382
rect 2915 250605 2925 251382
rect 2757 250346 2925 250605
rect 2757 249569 2767 250346
rect 2915 249569 2925 250346
rect 2757 249181 2925 249569
rect 2757 248404 2767 249181
rect 2915 248404 2925 249181
rect 2757 248145 2925 248404
rect 2757 247368 2767 248145
rect 2915 247368 2925 248145
rect 2757 247109 2925 247368
rect 2757 246332 2767 247109
rect 2915 246332 2925 247109
rect 2757 246073 2925 246332
rect 2757 245296 2767 246073
rect 2915 245296 2925 246073
rect 2757 245037 2925 245296
rect 2757 244260 2767 245037
rect 2915 244260 2925 245037
rect 2757 244248 2925 244260
rect 2967 254490 3135 254501
rect 2967 253713 2977 254490
rect 3125 253713 3135 254490
rect 2967 253454 3135 253713
rect 2967 252677 2977 253454
rect 3125 252677 3135 253454
rect 2967 252418 3135 252677
rect 2967 251641 2977 252418
rect 3125 251641 3135 252418
rect 2967 251382 3135 251641
rect 2967 250605 2977 251382
rect 3125 250605 3135 251382
rect 2967 250346 3135 250605
rect 2967 249569 2977 250346
rect 3125 249569 3135 250346
rect 2967 249181 3135 249569
rect 2967 248404 2977 249181
rect 3125 248404 3135 249181
rect 2967 248145 3135 248404
rect 2967 247368 2977 248145
rect 3125 247368 3135 248145
rect 2967 247109 3135 247368
rect 2967 246332 2977 247109
rect 3125 246332 3135 247109
rect 2967 246073 3135 246332
rect 2967 245296 2977 246073
rect 3125 245296 3135 246073
rect 2967 245037 3135 245296
rect 2967 244260 2977 245037
rect 3125 244260 3135 245037
rect 2967 244075 3135 244260
rect 3177 254490 3345 254737
rect 3177 253713 3187 254490
rect 3335 253713 3345 254490
rect 3177 253454 3345 253713
rect 3177 252677 3187 253454
rect 3335 252677 3345 253454
rect 3177 252418 3345 252677
rect 3177 251641 3187 252418
rect 3335 251641 3345 252418
rect 3177 251382 3345 251641
rect 3177 250605 3187 251382
rect 3335 250605 3345 251382
rect 3177 250346 3345 250605
rect 3177 249569 3187 250346
rect 3335 249569 3345 250346
rect 3177 249181 3345 249569
rect 3177 248404 3187 249181
rect 3335 248404 3345 249181
rect 3177 248145 3345 248404
rect 3177 247368 3187 248145
rect 3335 247368 3345 248145
rect 3177 247109 3345 247368
rect 3177 246332 3187 247109
rect 3335 246332 3345 247109
rect 3177 246073 3345 246332
rect 3177 245296 3187 246073
rect 3335 245296 3345 246073
rect 3177 245037 3345 245296
rect 3177 244260 3187 245037
rect 3335 244260 3345 245037
rect 3177 244248 3345 244260
rect 3387 254490 3555 254501
rect 3387 253713 3397 254490
rect 3545 253713 3555 254490
rect 3387 253454 3555 253713
rect 3387 252677 3397 253454
rect 3545 252677 3555 253454
rect 3387 252418 3555 252677
rect 3387 251641 3397 252418
rect 3545 251641 3555 252418
rect 3387 251382 3555 251641
rect 3387 250605 3397 251382
rect 3545 250605 3555 251382
rect 3387 250346 3555 250605
rect 3387 249569 3397 250346
rect 3545 249569 3555 250346
rect 3387 249181 3555 249569
rect 3387 248404 3397 249181
rect 3545 248404 3555 249181
rect 3387 248145 3555 248404
rect 3387 247368 3397 248145
rect 3545 247368 3555 248145
rect 3387 247109 3555 247368
rect 3387 246332 3397 247109
rect 3545 246332 3555 247109
rect 3387 246073 3555 246332
rect 3387 245296 3397 246073
rect 3545 245296 3555 246073
rect 3387 245037 3555 245296
rect 3387 244260 3397 245037
rect 3545 244260 3555 245037
rect 3387 244075 3555 244260
rect 3597 254490 3765 254737
rect 3597 253713 3607 254490
rect 3755 253713 3765 254490
rect 3597 253454 3765 253713
rect 3597 252677 3607 253454
rect 3755 252677 3765 253454
rect 3597 252418 3765 252677
rect 3597 251641 3607 252418
rect 3755 251641 3765 252418
rect 3597 251382 3765 251641
rect 3597 250605 3607 251382
rect 3755 250605 3765 251382
rect 3597 250346 3765 250605
rect 3597 249569 3607 250346
rect 3755 249569 3765 250346
rect 3597 249181 3765 249569
rect 3597 248404 3607 249181
rect 3755 248404 3765 249181
rect 3597 248145 3765 248404
rect 3597 247368 3607 248145
rect 3755 247368 3765 248145
rect 3597 247109 3765 247368
rect 3597 246332 3607 247109
rect 3755 246332 3765 247109
rect 3597 246073 3765 246332
rect 3597 245296 3607 246073
rect 3755 245296 3765 246073
rect 3597 245037 3765 245296
rect 3597 244260 3607 245037
rect 3755 244260 3765 245037
rect 3597 244248 3765 244260
rect 3807 254490 3975 254501
rect 3807 253713 3817 254490
rect 3965 253713 3975 254490
rect 3807 253454 3975 253713
rect 3807 252677 3817 253454
rect 3965 252677 3975 253454
rect 3807 252418 3975 252677
rect 3807 251641 3817 252418
rect 3965 251641 3975 252418
rect 3807 251382 3975 251641
rect 3807 250605 3817 251382
rect 3965 250605 3975 251382
rect 3807 250346 3975 250605
rect 3807 249569 3817 250346
rect 3965 249569 3975 250346
rect 3807 249181 3975 249569
rect 3807 248404 3817 249181
rect 3965 248404 3975 249181
rect 3807 248145 3975 248404
rect 3807 247368 3817 248145
rect 3965 247368 3975 248145
rect 3807 247109 3975 247368
rect 3807 246332 3817 247109
rect 3965 246332 3975 247109
rect 3807 246073 3975 246332
rect 3807 245296 3817 246073
rect 3965 245296 3975 246073
rect 3807 245037 3975 245296
rect 3807 244260 3817 245037
rect 3965 244260 3975 245037
rect 3807 244075 3975 244260
rect 4017 254490 4185 254737
rect 4017 253713 4027 254490
rect 4175 253713 4185 254490
rect 4017 253454 4185 253713
rect 4017 252677 4027 253454
rect 4175 252677 4185 253454
rect 4017 252418 4185 252677
rect 4017 251641 4027 252418
rect 4175 251641 4185 252418
rect 4017 251382 4185 251641
rect 4017 250605 4027 251382
rect 4175 250605 4185 251382
rect 4017 250346 4185 250605
rect 4017 249569 4027 250346
rect 4175 249569 4185 250346
rect 4017 249181 4185 249569
rect 4017 248404 4027 249181
rect 4175 248404 4185 249181
rect 4017 248145 4185 248404
rect 4017 247368 4027 248145
rect 4175 247368 4185 248145
rect 4017 247109 4185 247368
rect 4017 246332 4027 247109
rect 4175 246332 4185 247109
rect 4017 246073 4185 246332
rect 4017 245296 4027 246073
rect 4175 245296 4185 246073
rect 4017 245037 4185 245296
rect 4017 244260 4027 245037
rect 4175 244260 4185 245037
rect 4017 244248 4185 244260
rect 4227 254490 4395 254501
rect 4227 253713 4237 254490
rect 4385 253713 4395 254490
rect 4227 253454 4395 253713
rect 4227 252677 4237 253454
rect 4385 252677 4395 253454
rect 4227 252418 4395 252677
rect 4227 251641 4237 252418
rect 4385 251641 4395 252418
rect 4227 251382 4395 251641
rect 4227 250605 4237 251382
rect 4385 250605 4395 251382
rect 4227 250346 4395 250605
rect 4227 249569 4237 250346
rect 4385 249569 4395 250346
rect 4227 249181 4395 249569
rect 4227 248404 4237 249181
rect 4385 248404 4395 249181
rect 4227 248145 4395 248404
rect 4227 247368 4237 248145
rect 4385 247368 4395 248145
rect 4227 247109 4395 247368
rect 4227 246332 4237 247109
rect 4385 246332 4395 247109
rect 4227 246073 4395 246332
rect 4227 245296 4237 246073
rect 4385 245296 4395 246073
rect 4227 245037 4395 245296
rect 4227 244260 4237 245037
rect 4385 244260 4395 245037
rect 4227 244075 4395 244260
rect 4437 254490 4605 254737
rect 4437 253713 4447 254490
rect 4595 253713 4605 254490
rect 4437 253454 4605 253713
rect 4437 252677 4447 253454
rect 4595 252677 4605 253454
rect 4437 252418 4605 252677
rect 4437 251641 4447 252418
rect 4595 251641 4605 252418
rect 4437 251382 4605 251641
rect 4437 250605 4447 251382
rect 4595 250605 4605 251382
rect 4437 250346 4605 250605
rect 4437 249569 4447 250346
rect 4595 249569 4605 250346
rect 4437 249181 4605 249569
rect 4437 248404 4447 249181
rect 4595 248404 4605 249181
rect 4437 248145 4605 248404
rect 4437 247368 4447 248145
rect 4595 247368 4605 248145
rect 4437 247109 4605 247368
rect 4437 246332 4447 247109
rect 4595 246332 4605 247109
rect 4437 246073 4605 246332
rect 4437 245296 4447 246073
rect 4595 245296 4605 246073
rect 4437 245037 4605 245296
rect 4437 244260 4447 245037
rect 4595 244260 4605 245037
rect 4437 244248 4605 244260
rect 4647 254490 4815 254501
rect 4647 253713 4657 254490
rect 4805 253713 4815 254490
rect 4647 253454 4815 253713
rect 4647 252677 4657 253454
rect 4805 252677 4815 253454
rect 4647 252418 4815 252677
rect 4647 251641 4657 252418
rect 4805 251641 4815 252418
rect 4647 251382 4815 251641
rect 4647 250605 4657 251382
rect 4805 250605 4815 251382
rect 4647 250346 4815 250605
rect 4647 249569 4657 250346
rect 4805 249569 4815 250346
rect 4647 249181 4815 249569
rect 4647 248404 4657 249181
rect 4805 248404 4815 249181
rect 4647 248145 4815 248404
rect 4647 247368 4657 248145
rect 4805 247368 4815 248145
rect 4647 247109 4815 247368
rect 4647 246332 4657 247109
rect 4805 246332 4815 247109
rect 4647 246073 4815 246332
rect 4647 245296 4657 246073
rect 4805 245296 4815 246073
rect 4647 245037 4815 245296
rect 4647 244260 4657 245037
rect 4805 244260 4815 245037
rect 4647 244075 4815 244260
rect 4857 254490 5025 254737
rect 4857 253713 4867 254490
rect 5015 253713 5025 254490
rect 4857 253454 5025 253713
rect 4857 252677 4867 253454
rect 5015 252677 5025 253454
rect 4857 252418 5025 252677
rect 4857 251641 4867 252418
rect 5015 251641 5025 252418
rect 4857 251382 5025 251641
rect 4857 250605 4867 251382
rect 5015 250605 5025 251382
rect 4857 250346 5025 250605
rect 4857 249569 4867 250346
rect 5015 249569 5025 250346
rect 4857 249181 5025 249569
rect 4857 248404 4867 249181
rect 5015 248404 5025 249181
rect 4857 248145 5025 248404
rect 4857 247368 4867 248145
rect 5015 247368 5025 248145
rect 4857 247109 5025 247368
rect 4857 246332 4867 247109
rect 5015 246332 5025 247109
rect 4857 246073 5025 246332
rect 4857 245296 4867 246073
rect 5015 245296 5025 246073
rect 4857 245037 5025 245296
rect 4857 244260 4867 245037
rect 5015 244260 5025 245037
rect 4857 244248 5025 244260
rect 5067 254490 5235 254501
rect 5067 253713 5077 254490
rect 5225 253713 5235 254490
rect 5067 253454 5235 253713
rect 5067 252677 5077 253454
rect 5225 252677 5235 253454
rect 5067 252418 5235 252677
rect 5067 251641 5077 252418
rect 5225 251641 5235 252418
rect 5067 251382 5235 251641
rect 5067 250605 5077 251382
rect 5225 250605 5235 251382
rect 5067 250346 5235 250605
rect 5067 249569 5077 250346
rect 5225 249569 5235 250346
rect 5067 249181 5235 249569
rect 5067 248404 5077 249181
rect 5225 248404 5235 249181
rect 5067 248145 5235 248404
rect 5067 247368 5077 248145
rect 5225 247368 5235 248145
rect 5067 247109 5235 247368
rect 5067 246332 5077 247109
rect 5225 246332 5235 247109
rect 5067 246073 5235 246332
rect 5067 245296 5077 246073
rect 5225 245296 5235 246073
rect 5067 245037 5235 245296
rect 5067 244260 5077 245037
rect 5225 244260 5235 245037
rect 5067 244075 5235 244260
rect 5277 254490 5445 254737
rect 5277 253713 5287 254490
rect 5435 253713 5445 254490
rect 5277 253454 5445 253713
rect 5277 252677 5287 253454
rect 5435 252677 5445 253454
rect 5277 252418 5445 252677
rect 5277 251641 5287 252418
rect 5435 251641 5445 252418
rect 5277 251382 5445 251641
rect 5277 250605 5287 251382
rect 5435 250605 5445 251382
rect 5277 250346 5445 250605
rect 5277 249569 5287 250346
rect 5435 249569 5445 250346
rect 5277 249181 5445 249569
rect 5277 248404 5287 249181
rect 5435 248404 5445 249181
rect 5277 248145 5445 248404
rect 5277 247368 5287 248145
rect 5435 247368 5445 248145
rect 5277 247109 5445 247368
rect 5277 246332 5287 247109
rect 5435 246332 5445 247109
rect 5277 246073 5445 246332
rect 5277 245296 5287 246073
rect 5435 245296 5445 246073
rect 5277 245037 5445 245296
rect 5277 244260 5287 245037
rect 5435 244260 5445 245037
rect 5277 244248 5445 244260
rect 5487 254490 5655 254501
rect 5487 253713 5497 254490
rect 5645 253713 5655 254490
rect 5487 253454 5655 253713
rect 5487 252677 5497 253454
rect 5645 252677 5655 253454
rect 5487 252418 5655 252677
rect 5487 251641 5497 252418
rect 5645 251641 5655 252418
rect 5487 251382 5655 251641
rect 5487 250605 5497 251382
rect 5645 250605 5655 251382
rect 5487 250346 5655 250605
rect 5487 249569 5497 250346
rect 5645 249569 5655 250346
rect 5487 249181 5655 249569
rect 5487 248404 5497 249181
rect 5645 248404 5655 249181
rect 5487 248145 5655 248404
rect 5487 247368 5497 248145
rect 5645 247368 5655 248145
rect 5487 247109 5655 247368
rect 5487 246332 5497 247109
rect 5645 246332 5655 247109
rect 5487 246073 5655 246332
rect 5487 245296 5497 246073
rect 5645 245296 5655 246073
rect 5487 245037 5655 245296
rect 5487 244260 5497 245037
rect 5645 244260 5655 245037
rect 5487 244075 5655 244260
rect 5697 254490 5865 254737
rect 5697 253713 5707 254490
rect 5855 253713 5865 254490
rect 5697 253454 5865 253713
rect 5697 252677 5707 253454
rect 5855 252677 5865 253454
rect 5697 252418 5865 252677
rect 5697 251641 5707 252418
rect 5855 251641 5865 252418
rect 5697 251382 5865 251641
rect 5697 250605 5707 251382
rect 5855 250605 5865 251382
rect 5697 250346 5865 250605
rect 5697 249569 5707 250346
rect 5855 249569 5865 250346
rect 5697 249181 5865 249569
rect 5697 248404 5707 249181
rect 5855 248404 5865 249181
rect 5697 248145 5865 248404
rect 5697 247368 5707 248145
rect 5855 247368 5865 248145
rect 5697 247109 5865 247368
rect 5697 246332 5707 247109
rect 5855 246332 5865 247109
rect 5697 246073 5865 246332
rect 5697 245296 5707 246073
rect 5855 245296 5865 246073
rect 5697 245037 5865 245296
rect 5697 244260 5707 245037
rect 5855 244260 5865 245037
rect 5697 244248 5865 244260
rect 5907 254490 6075 254501
rect 5907 253713 5917 254490
rect 6065 253713 6075 254490
rect 5907 253454 6075 253713
rect 5907 252677 5917 253454
rect 6065 252677 6075 253454
rect 5907 252418 6075 252677
rect 5907 251641 5917 252418
rect 6065 251641 6075 252418
rect 5907 251382 6075 251641
rect 5907 250605 5917 251382
rect 6065 250605 6075 251382
rect 5907 250346 6075 250605
rect 5907 249569 5917 250346
rect 6065 249569 6075 250346
rect 5907 249181 6075 249569
rect 5907 248404 5917 249181
rect 6065 248404 6075 249181
rect 5907 248145 6075 248404
rect 5907 247368 5917 248145
rect 6065 247368 6075 248145
rect 5907 247109 6075 247368
rect 5907 246332 5917 247109
rect 6065 246332 6075 247109
rect 5907 246073 6075 246332
rect 5907 245296 5917 246073
rect 6065 245296 6075 246073
rect 5907 245037 6075 245296
rect 5907 244260 5917 245037
rect 6065 244260 6075 245037
rect 5907 244075 6075 244260
rect 6117 254490 6285 254737
rect 6117 253713 6127 254490
rect 6275 253713 6285 254490
rect 6117 253454 6285 253713
rect 6117 252677 6127 253454
rect 6275 252677 6285 253454
rect 6117 252418 6285 252677
rect 6117 251641 6127 252418
rect 6275 251641 6285 252418
rect 6117 251382 6285 251641
rect 6117 250605 6127 251382
rect 6275 250605 6285 251382
rect 6117 250346 6285 250605
rect 6117 249569 6127 250346
rect 6275 249569 6285 250346
rect 6117 249181 6285 249569
rect 6117 248404 6127 249181
rect 6275 248404 6285 249181
rect 6117 248145 6285 248404
rect 6117 247368 6127 248145
rect 6275 247368 6285 248145
rect 6117 247109 6285 247368
rect 6117 246332 6127 247109
rect 6275 246332 6285 247109
rect 6117 246073 6285 246332
rect 6117 245296 6127 246073
rect 6275 245296 6285 246073
rect 6117 245037 6285 245296
rect 6117 244260 6127 245037
rect 6275 244260 6285 245037
rect 6117 244248 6285 244260
rect 6327 254490 6495 254501
rect 6327 253713 6337 254490
rect 6485 253713 6495 254490
rect 6327 253454 6495 253713
rect 6327 252677 6337 253454
rect 6485 252677 6495 253454
rect 6327 252418 6495 252677
rect 6327 251641 6337 252418
rect 6485 251641 6495 252418
rect 6327 251382 6495 251641
rect 6327 250605 6337 251382
rect 6485 250605 6495 251382
rect 6327 250346 6495 250605
rect 6327 249569 6337 250346
rect 6485 249569 6495 250346
rect 6327 249181 6495 249569
rect 6327 248404 6337 249181
rect 6485 248404 6495 249181
rect 6327 248145 6495 248404
rect 6327 247368 6337 248145
rect 6485 247368 6495 248145
rect 6327 247109 6495 247368
rect 6327 246332 6337 247109
rect 6485 246332 6495 247109
rect 6327 246073 6495 246332
rect 6327 245296 6337 246073
rect 6485 245296 6495 246073
rect 6327 245037 6495 245296
rect 6327 244260 6337 245037
rect 6485 244260 6495 245037
rect 6327 244075 6495 244260
rect 6537 254490 6705 254737
rect 6537 253713 6547 254490
rect 6695 253713 6705 254490
rect 6537 253454 6705 253713
rect 6537 252677 6547 253454
rect 6695 252677 6705 253454
rect 6537 252418 6705 252677
rect 6537 251641 6547 252418
rect 6695 251641 6705 252418
rect 6537 251382 6705 251641
rect 6537 250605 6547 251382
rect 6695 250605 6705 251382
rect 6537 250346 6705 250605
rect 6537 249569 6547 250346
rect 6695 249569 6705 250346
rect 6537 249181 6705 249569
rect 6537 248404 6547 249181
rect 6695 248404 6705 249181
rect 6537 248145 6705 248404
rect 6537 247368 6547 248145
rect 6695 247368 6705 248145
rect 6537 247109 6705 247368
rect 6537 246332 6547 247109
rect 6695 246332 6705 247109
rect 6537 246073 6705 246332
rect 6537 245296 6547 246073
rect 6695 245296 6705 246073
rect 6537 245037 6705 245296
rect 6537 244260 6547 245037
rect 6695 244260 6705 245037
rect 6537 244248 6705 244260
rect 6747 254490 6915 254501
rect 6747 253713 6757 254490
rect 6905 253713 6915 254490
rect 6747 253454 6915 253713
rect 6747 252677 6757 253454
rect 6905 252677 6915 253454
rect 6747 252418 6915 252677
rect 6747 251641 6757 252418
rect 6905 251641 6915 252418
rect 6747 251382 6915 251641
rect 6747 250605 6757 251382
rect 6905 250605 6915 251382
rect 6747 250346 6915 250605
rect 6747 249569 6757 250346
rect 6905 249569 6915 250346
rect 6747 249181 6915 249569
rect 6747 248404 6757 249181
rect 6905 248404 6915 249181
rect 6747 248145 6915 248404
rect 6747 247368 6757 248145
rect 6905 247368 6915 248145
rect 6747 247109 6915 247368
rect 6747 246332 6757 247109
rect 6905 246332 6915 247109
rect 6747 246073 6915 246332
rect 6747 245296 6757 246073
rect 6905 245296 6915 246073
rect 6747 245037 6915 245296
rect 6747 244260 6757 245037
rect 6905 244260 6915 245037
rect 6747 244075 6915 244260
rect 6957 254490 7125 254737
rect 6957 253713 6967 254490
rect 7115 253713 7125 254490
rect 6957 253454 7125 253713
rect 6957 252677 6967 253454
rect 7115 252677 7125 253454
rect 6957 252418 7125 252677
rect 6957 251641 6967 252418
rect 7115 251641 7125 252418
rect 6957 251382 7125 251641
rect 6957 250605 6967 251382
rect 7115 250605 7125 251382
rect 6957 250346 7125 250605
rect 6957 249569 6967 250346
rect 7115 249569 7125 250346
rect 6957 249181 7125 249569
rect 6957 248404 6967 249181
rect 7115 248404 7125 249181
rect 6957 248145 7125 248404
rect 6957 247368 6967 248145
rect 7115 247368 7125 248145
rect 6957 247109 7125 247368
rect 6957 246332 6967 247109
rect 7115 246332 7125 247109
rect 6957 246073 7125 246332
rect 6957 245296 6967 246073
rect 7115 245296 7125 246073
rect 6957 245037 7125 245296
rect 6957 244260 6967 245037
rect 7115 244260 7125 245037
rect 6957 244248 7125 244260
rect 7167 254490 7335 254501
rect 7167 253713 7177 254490
rect 7325 253713 7335 254490
rect 7167 253454 7335 253713
rect 7167 252677 7177 253454
rect 7325 252677 7335 253454
rect 7167 252418 7335 252677
rect 7167 251641 7177 252418
rect 7325 251641 7335 252418
rect 7167 251382 7335 251641
rect 7167 250605 7177 251382
rect 7325 250605 7335 251382
rect 7167 250346 7335 250605
rect 7167 249569 7177 250346
rect 7325 249569 7335 250346
rect 7167 249181 7335 249569
rect 7167 248404 7177 249181
rect 7325 248404 7335 249181
rect 7167 248145 7335 248404
rect 7167 247368 7177 248145
rect 7325 247368 7335 248145
rect 7167 247109 7335 247368
rect 7167 246332 7177 247109
rect 7325 246332 7335 247109
rect 7167 246073 7335 246332
rect 7167 245296 7177 246073
rect 7325 245296 7335 246073
rect 7167 245037 7335 245296
rect 7167 244260 7177 245037
rect 7325 244260 7335 245037
rect 7167 244075 7335 244260
rect 7377 254490 7545 254737
rect 7377 253713 7387 254490
rect 7535 253713 7545 254490
rect 7377 253454 7545 253713
rect 7377 252677 7387 253454
rect 7535 252677 7545 253454
rect 7377 252418 7545 252677
rect 7377 251641 7387 252418
rect 7535 251641 7545 252418
rect 7377 251382 7545 251641
rect 7377 250605 7387 251382
rect 7535 250605 7545 251382
rect 7377 250346 7545 250605
rect 7377 249569 7387 250346
rect 7535 249569 7545 250346
rect 7377 249181 7545 249569
rect 7377 248404 7387 249181
rect 7535 248404 7545 249181
rect 7377 248145 7545 248404
rect 7377 247368 7387 248145
rect 7535 247368 7545 248145
rect 7377 247109 7545 247368
rect 7377 246332 7387 247109
rect 7535 246332 7545 247109
rect 7377 246073 7545 246332
rect 7377 245296 7387 246073
rect 7535 245296 7545 246073
rect 7377 245037 7545 245296
rect 7377 244260 7387 245037
rect 7535 244260 7545 245037
rect 7377 244248 7545 244260
rect 7587 254490 7755 254501
rect 7587 253713 7597 254490
rect 7745 253713 7755 254490
rect 7587 253454 7755 253713
rect 7587 252677 7597 253454
rect 7745 252677 7755 253454
rect 7587 252418 7755 252677
rect 7587 251641 7597 252418
rect 7745 251641 7755 252418
rect 7587 251382 7755 251641
rect 7587 250605 7597 251382
rect 7745 250605 7755 251382
rect 7587 250346 7755 250605
rect 7587 249569 7597 250346
rect 7745 249569 7755 250346
rect 7587 249181 7755 249569
rect 7587 248404 7597 249181
rect 7745 248404 7755 249181
rect 7587 248145 7755 248404
rect 7587 247368 7597 248145
rect 7745 247368 7755 248145
rect 7587 247109 7755 247368
rect 7587 246332 7597 247109
rect 7745 246332 7755 247109
rect 7587 246073 7755 246332
rect 7587 245296 7597 246073
rect 7745 245296 7755 246073
rect 7587 245037 7755 245296
rect 7587 244260 7597 245037
rect 7745 244260 7755 245037
rect 7587 244075 7755 244260
rect 7797 254490 7965 254737
rect 7797 253713 7807 254490
rect 7955 253713 7965 254490
rect 7797 253454 7965 253713
rect 7797 252677 7807 253454
rect 7955 252677 7965 253454
rect 7797 252418 7965 252677
rect 7797 251641 7807 252418
rect 7955 251641 7965 252418
rect 7797 251382 7965 251641
rect 7797 250605 7807 251382
rect 7955 250605 7965 251382
rect 7797 250346 7965 250605
rect 7797 249569 7807 250346
rect 7955 249569 7965 250346
rect 7797 249181 7965 249569
rect 7797 248404 7807 249181
rect 7955 248404 7965 249181
rect 7797 248145 7965 248404
rect 7797 247368 7807 248145
rect 7955 247368 7965 248145
rect 7797 247109 7965 247368
rect 7797 246332 7807 247109
rect 7955 246332 7965 247109
rect 7797 246073 7965 246332
rect 7797 245296 7807 246073
rect 7955 245296 7965 246073
rect 7797 245037 7965 245296
rect 7797 244260 7807 245037
rect 7955 244260 7965 245037
rect 7797 244248 7965 244260
rect 8007 254490 8175 254501
rect 8007 253713 8017 254490
rect 8165 253713 8175 254490
rect 8007 253454 8175 253713
rect 8007 252677 8017 253454
rect 8165 252677 8175 253454
rect 8007 252418 8175 252677
rect 8007 251641 8017 252418
rect 8165 251641 8175 252418
rect 8007 251382 8175 251641
rect 8007 250605 8017 251382
rect 8165 250605 8175 251382
rect 8007 250346 8175 250605
rect 8007 249569 8017 250346
rect 8165 249569 8175 250346
rect 8007 249181 8175 249569
rect 8007 248404 8017 249181
rect 8165 248404 8175 249181
rect 8007 248145 8175 248404
rect 8007 247368 8017 248145
rect 8165 247368 8175 248145
rect 8007 247109 8175 247368
rect 8007 246332 8017 247109
rect 8165 246332 8175 247109
rect 8007 246073 8175 246332
rect 8007 245296 8017 246073
rect 8165 245296 8175 246073
rect 8007 245037 8175 245296
rect 8007 244260 8017 245037
rect 8165 244260 8175 245037
rect 8007 244075 8175 244260
rect 8217 254490 8385 254737
rect 8217 253713 8227 254490
rect 8375 253713 8385 254490
rect 8217 253454 8385 253713
rect 8217 252677 8227 253454
rect 8375 252677 8385 253454
rect 8217 252418 8385 252677
rect 8217 251641 8227 252418
rect 8375 251641 8385 252418
rect 8217 251382 8385 251641
rect 8217 250605 8227 251382
rect 8375 250605 8385 251382
rect 8217 250346 8385 250605
rect 8217 249569 8227 250346
rect 8375 249569 8385 250346
rect 8217 249181 8385 249569
rect 8217 248404 8227 249181
rect 8375 248404 8385 249181
rect 8217 248145 8385 248404
rect 8217 247368 8227 248145
rect 8375 247368 8385 248145
rect 8217 247109 8385 247368
rect 8217 246332 8227 247109
rect 8375 246332 8385 247109
rect 8217 246073 8385 246332
rect 8217 245296 8227 246073
rect 8375 245296 8385 246073
rect 8217 245037 8385 245296
rect 8217 244260 8227 245037
rect 8375 244260 8385 245037
rect 8217 244248 8385 244260
rect 8427 254490 8595 254501
rect 8427 253713 8437 254490
rect 8585 253713 8595 254490
rect 8427 253454 8595 253713
rect 8427 252677 8437 253454
rect 8585 252677 8595 253454
rect 8427 252418 8595 252677
rect 8427 251641 8437 252418
rect 8585 251641 8595 252418
rect 8427 251382 8595 251641
rect 8427 250605 8437 251382
rect 8585 250605 8595 251382
rect 8427 250346 8595 250605
rect 8427 249569 8437 250346
rect 8585 249569 8595 250346
rect 8427 249181 8595 249569
rect 8427 248404 8437 249181
rect 8585 248404 8595 249181
rect 8427 248145 8595 248404
rect 8427 247368 8437 248145
rect 8585 247368 8595 248145
rect 8427 247109 8595 247368
rect 8427 246332 8437 247109
rect 8585 246332 8595 247109
rect 8427 246073 8595 246332
rect 8427 245296 8437 246073
rect 8585 245296 8595 246073
rect 8427 245037 8595 245296
rect 8427 244260 8437 245037
rect 8585 244260 8595 245037
rect 8427 244075 8595 244260
rect 8637 254490 8805 254737
rect 8637 253713 8647 254490
rect 8795 253713 8805 254490
rect 8637 253454 8805 253713
rect 8637 252677 8647 253454
rect 8795 252677 8805 253454
rect 8637 252418 8805 252677
rect 8637 251641 8647 252418
rect 8795 251641 8805 252418
rect 8637 251382 8805 251641
rect 8637 250605 8647 251382
rect 8795 250605 8805 251382
rect 8637 250346 8805 250605
rect 8637 249569 8647 250346
rect 8795 249569 8805 250346
rect 8637 249181 8805 249569
rect 8637 248404 8647 249181
rect 8795 248404 8805 249181
rect 8637 248145 8805 248404
rect 8637 247368 8647 248145
rect 8795 247368 8805 248145
rect 8637 247109 8805 247368
rect 8637 246332 8647 247109
rect 8795 246332 8805 247109
rect 8637 246073 8805 246332
rect 8637 245296 8647 246073
rect 8795 245296 8805 246073
rect 8637 245037 8805 245296
rect 8637 244260 8647 245037
rect 8795 244260 8805 245037
rect 8637 244248 8805 244260
rect 8847 254490 9015 254501
rect 8847 253713 8857 254490
rect 9005 253713 9015 254490
rect 8847 253454 9015 253713
rect 8847 252677 8857 253454
rect 9005 252677 9015 253454
rect 8847 252418 9015 252677
rect 8847 251641 8857 252418
rect 9005 251641 9015 252418
rect 8847 251382 9015 251641
rect 8847 250605 8857 251382
rect 9005 250605 9015 251382
rect 8847 250346 9015 250605
rect 8847 249569 8857 250346
rect 9005 249569 9015 250346
rect 8847 249181 9015 249569
rect 8847 248404 8857 249181
rect 9005 248404 9015 249181
rect 8847 248145 9015 248404
rect 8847 247368 8857 248145
rect 9005 247368 9015 248145
rect 8847 247109 9015 247368
rect 8847 246332 8857 247109
rect 9005 246332 9015 247109
rect 8847 246073 9015 246332
rect 8847 245296 8857 246073
rect 9005 245296 9015 246073
rect 8847 245037 9015 245296
rect 8847 244260 8857 245037
rect 9005 244260 9015 245037
rect 8847 244075 9015 244260
rect 9057 254490 9225 254737
rect 9057 253713 9067 254490
rect 9215 253713 9225 254490
rect 9057 253454 9225 253713
rect 9057 252677 9067 253454
rect 9215 252677 9225 253454
rect 9057 252418 9225 252677
rect 9057 251641 9067 252418
rect 9215 251641 9225 252418
rect 9057 251382 9225 251641
rect 9057 250605 9067 251382
rect 9215 250605 9225 251382
rect 9057 250346 9225 250605
rect 9057 249569 9067 250346
rect 9215 249569 9225 250346
rect 9057 249181 9225 249569
rect 9057 248404 9067 249181
rect 9215 248404 9225 249181
rect 9057 248145 9225 248404
rect 9057 247368 9067 248145
rect 9215 247368 9225 248145
rect 9057 247109 9225 247368
rect 9057 246332 9067 247109
rect 9215 246332 9225 247109
rect 9057 246073 9225 246332
rect 9057 245296 9067 246073
rect 9215 245296 9225 246073
rect 9057 245037 9225 245296
rect 9057 244260 9067 245037
rect 9215 244260 9225 245037
rect 9057 244248 9225 244260
rect 9267 254490 9435 254501
rect 9267 253713 9277 254490
rect 9425 253713 9435 254490
rect 9267 253454 9435 253713
rect 9267 252677 9277 253454
rect 9425 252677 9435 253454
rect 9267 252418 9435 252677
rect 9267 251641 9277 252418
rect 9425 251641 9435 252418
rect 9267 251382 9435 251641
rect 9267 250605 9277 251382
rect 9425 250605 9435 251382
rect 9267 250346 9435 250605
rect 9267 249569 9277 250346
rect 9425 249569 9435 250346
rect 9267 249181 9435 249569
rect 9267 248404 9277 249181
rect 9425 248404 9435 249181
rect 9267 248145 9435 248404
rect 9267 247368 9277 248145
rect 9425 247368 9435 248145
rect 9267 247109 9435 247368
rect 9267 246332 9277 247109
rect 9425 246332 9435 247109
rect 9267 246073 9435 246332
rect 9267 245296 9277 246073
rect 9425 245296 9435 246073
rect 9267 245037 9435 245296
rect 9267 244260 9277 245037
rect 9425 244260 9435 245037
rect 9267 244075 9435 244260
rect 9477 254490 9645 254737
rect 9477 253713 9487 254490
rect 9635 253713 9645 254490
rect 9477 253454 9645 253713
rect 9477 252677 9487 253454
rect 9635 252677 9645 253454
rect 9477 252418 9645 252677
rect 9477 251641 9487 252418
rect 9635 251641 9645 252418
rect 9477 251382 9645 251641
rect 9477 250605 9487 251382
rect 9635 250605 9645 251382
rect 9477 250346 9645 250605
rect 9477 249569 9487 250346
rect 9635 249569 9645 250346
rect 9477 249181 9645 249569
rect 9477 248404 9487 249181
rect 9635 248404 9645 249181
rect 9477 248145 9645 248404
rect 9477 247368 9487 248145
rect 9635 247368 9645 248145
rect 9477 247109 9645 247368
rect 9477 246332 9487 247109
rect 9635 246332 9645 247109
rect 9477 246073 9645 246332
rect 9477 245296 9487 246073
rect 9635 245296 9645 246073
rect 9477 245037 9645 245296
rect 9477 244260 9487 245037
rect 9635 244260 9645 245037
rect 9477 244248 9645 244260
rect 9687 254490 9855 254501
rect 9687 253713 9697 254490
rect 9845 253713 9855 254490
rect 9687 253454 9855 253713
rect 9687 252677 9697 253454
rect 9845 252677 9855 253454
rect 9687 252418 9855 252677
rect 9687 251641 9697 252418
rect 9845 251641 9855 252418
rect 9687 251382 9855 251641
rect 9687 250605 9697 251382
rect 9845 250605 9855 251382
rect 9687 250346 9855 250605
rect 9687 249569 9697 250346
rect 9845 249569 9855 250346
rect 9687 249181 9855 249569
rect 9687 248404 9697 249181
rect 9845 248404 9855 249181
rect 9687 248145 9855 248404
rect 9687 247368 9697 248145
rect 9845 247368 9855 248145
rect 9687 247109 9855 247368
rect 9687 246332 9697 247109
rect 9845 246332 9855 247109
rect 9687 246073 9855 246332
rect 9687 245296 9697 246073
rect 9845 245296 9855 246073
rect 9687 245037 9855 245296
rect 9687 244260 9697 245037
rect 9845 244260 9855 245037
rect 9687 244075 9855 244260
rect 9897 254490 10065 254737
rect 9897 253713 9907 254490
rect 10055 253713 10065 254490
rect 9897 253454 10065 253713
rect 9897 252677 9907 253454
rect 10055 252677 10065 253454
rect 9897 252418 10065 252677
rect 9897 251641 9907 252418
rect 10055 251641 10065 252418
rect 9897 251382 10065 251641
rect 9897 250605 9907 251382
rect 10055 250605 10065 251382
rect 9897 250346 10065 250605
rect 9897 249569 9907 250346
rect 10055 249569 10065 250346
rect 9897 249181 10065 249569
rect 9897 248404 9907 249181
rect 10055 248404 10065 249181
rect 9897 248145 10065 248404
rect 9897 247368 9907 248145
rect 10055 247368 10065 248145
rect 9897 247109 10065 247368
rect 9897 246332 9907 247109
rect 10055 246332 10065 247109
rect 9897 246073 10065 246332
rect 9897 245296 9907 246073
rect 10055 245296 10065 246073
rect 9897 245037 10065 245296
rect 9897 244260 9907 245037
rect 10055 244260 10065 245037
rect 9897 244248 10065 244260
rect 10107 254490 10275 254501
rect 10107 253713 10117 254490
rect 10265 253713 10275 254490
rect 10107 253454 10275 253713
rect 10107 252677 10117 253454
rect 10265 252677 10275 253454
rect 10107 252418 10275 252677
rect 10107 251641 10117 252418
rect 10265 251641 10275 252418
rect 10107 251382 10275 251641
rect 10107 250605 10117 251382
rect 10265 250605 10275 251382
rect 10107 250346 10275 250605
rect 10107 249569 10117 250346
rect 10265 249569 10275 250346
rect 10107 249181 10275 249569
rect 10107 248404 10117 249181
rect 10265 248404 10275 249181
rect 10107 248145 10275 248404
rect 10107 247368 10117 248145
rect 10265 247368 10275 248145
rect 10107 247109 10275 247368
rect 10107 246332 10117 247109
rect 10265 246332 10275 247109
rect 10107 246073 10275 246332
rect 10107 245296 10117 246073
rect 10265 245296 10275 246073
rect 10107 245037 10275 245296
rect 10107 244260 10117 245037
rect 10265 244260 10275 245037
rect 10107 244075 10275 244260
rect 10317 254490 10485 254737
rect 10317 253713 10327 254490
rect 10475 253713 10485 254490
rect 10317 253454 10485 253713
rect 10317 252677 10327 253454
rect 10475 252677 10485 253454
rect 10317 252418 10485 252677
rect 10317 251641 10327 252418
rect 10475 251641 10485 252418
rect 10317 251382 10485 251641
rect 10317 250605 10327 251382
rect 10475 250605 10485 251382
rect 10317 250346 10485 250605
rect 10317 249569 10327 250346
rect 10475 249569 10485 250346
rect 10317 249181 10485 249569
rect 10317 248404 10327 249181
rect 10475 248404 10485 249181
rect 10317 248145 10485 248404
rect 10317 247368 10327 248145
rect 10475 247368 10485 248145
rect 10317 247109 10485 247368
rect 10317 246332 10327 247109
rect 10475 246332 10485 247109
rect 10317 246073 10485 246332
rect 10317 245296 10327 246073
rect 10475 245296 10485 246073
rect 10317 245037 10485 245296
rect 10317 244260 10327 245037
rect 10475 244260 10485 245037
rect 10317 244248 10485 244260
rect 10527 254490 10695 254501
rect 10527 253713 10537 254490
rect 10685 253713 10695 254490
rect 10527 253454 10695 253713
rect 10527 252677 10537 253454
rect 10685 252677 10695 253454
rect 10527 252418 10695 252677
rect 10527 251641 10537 252418
rect 10685 251641 10695 252418
rect 10527 251382 10695 251641
rect 10527 250605 10537 251382
rect 10685 250605 10695 251382
rect 10527 250346 10695 250605
rect 10527 249569 10537 250346
rect 10685 249569 10695 250346
rect 10527 249181 10695 249569
rect 10527 248404 10537 249181
rect 10685 248404 10695 249181
rect 10527 248145 10695 248404
rect 10527 247368 10537 248145
rect 10685 247368 10695 248145
rect 10527 247109 10695 247368
rect 10527 246332 10537 247109
rect 10685 246332 10695 247109
rect 10527 246073 10695 246332
rect 10527 245296 10537 246073
rect 10685 245296 10695 246073
rect 10527 245037 10695 245296
rect 10527 244260 10537 245037
rect 10685 244260 10695 245037
rect 10527 244075 10695 244260
rect 10737 254490 10905 254737
rect 10737 253713 10747 254490
rect 10895 253713 10905 254490
rect 10737 253454 10905 253713
rect 10737 252677 10747 253454
rect 10895 252677 10905 253454
rect 10737 252418 10905 252677
rect 10737 251641 10747 252418
rect 10895 251641 10905 252418
rect 10737 251382 10905 251641
rect 10737 250605 10747 251382
rect 10895 250605 10905 251382
rect 10737 250346 10905 250605
rect 10737 249569 10747 250346
rect 10895 249569 10905 250346
rect 10737 249181 10905 249569
rect 10737 248404 10747 249181
rect 10895 248404 10905 249181
rect 10737 248145 10905 248404
rect 10737 247368 10747 248145
rect 10895 247368 10905 248145
rect 10737 247109 10905 247368
rect 10737 246332 10747 247109
rect 10895 246332 10905 247109
rect 10737 246073 10905 246332
rect 10737 245296 10747 246073
rect 10895 245296 10905 246073
rect 10737 245037 10905 245296
rect 10737 244260 10747 245037
rect 10895 244260 10905 245037
rect 10737 244248 10905 244260
rect 10947 254490 11115 254501
rect 10947 253713 10957 254490
rect 11105 253713 11115 254490
rect 10947 253454 11115 253713
rect 10947 252677 10957 253454
rect 11105 252677 11115 253454
rect 10947 252418 11115 252677
rect 10947 251641 10957 252418
rect 11105 251641 11115 252418
rect 10947 251382 11115 251641
rect 10947 250605 10957 251382
rect 11105 250605 11115 251382
rect 10947 250346 11115 250605
rect 10947 249569 10957 250346
rect 11105 249569 11115 250346
rect 10947 249181 11115 249569
rect 10947 248404 10957 249181
rect 11105 248404 11115 249181
rect 10947 248145 11115 248404
rect 10947 247368 10957 248145
rect 11105 247368 11115 248145
rect 10947 247109 11115 247368
rect 10947 246332 10957 247109
rect 11105 246332 11115 247109
rect 10947 246073 11115 246332
rect 10947 245296 10957 246073
rect 11105 245296 11115 246073
rect 10947 245037 11115 245296
rect 10947 244260 10957 245037
rect 11105 244260 11115 245037
rect 10947 244075 11115 244260
rect 11157 254490 11325 254737
rect 11157 253713 11167 254490
rect 11315 253713 11325 254490
rect 11157 253454 11325 253713
rect 11157 252677 11167 253454
rect 11315 252677 11325 253454
rect 11157 252418 11325 252677
rect 11157 251641 11167 252418
rect 11315 251641 11325 252418
rect 11157 251382 11325 251641
rect 11157 250605 11167 251382
rect 11315 250605 11325 251382
rect 11157 250346 11325 250605
rect 11157 249569 11167 250346
rect 11315 249569 11325 250346
rect 11157 249181 11325 249569
rect 11157 248404 11167 249181
rect 11315 248404 11325 249181
rect 11157 248145 11325 248404
rect 11157 247368 11167 248145
rect 11315 247368 11325 248145
rect 11157 247109 11325 247368
rect 11157 246332 11167 247109
rect 11315 246332 11325 247109
rect 11157 246073 11325 246332
rect 11157 245296 11167 246073
rect 11315 245296 11325 246073
rect 11157 245037 11325 245296
rect 11157 244260 11167 245037
rect 11315 244260 11325 245037
rect 11157 244248 11325 244260
rect 11367 254490 11535 254501
rect 11367 253713 11377 254490
rect 11525 253713 11535 254490
rect 11367 253454 11535 253713
rect 11367 252677 11377 253454
rect 11525 252677 11535 253454
rect 11367 252418 11535 252677
rect 11367 251641 11377 252418
rect 11525 251641 11535 252418
rect 11367 251382 11535 251641
rect 11367 250605 11377 251382
rect 11525 250605 11535 251382
rect 11367 250346 11535 250605
rect 11367 249569 11377 250346
rect 11525 249569 11535 250346
rect 11367 249181 11535 249569
rect 11367 248404 11377 249181
rect 11525 248404 11535 249181
rect 11367 248145 11535 248404
rect 11367 247368 11377 248145
rect 11525 247368 11535 248145
rect 11367 247109 11535 247368
rect 11367 246332 11377 247109
rect 11525 246332 11535 247109
rect 11367 246073 11535 246332
rect 11367 245296 11377 246073
rect 11525 245296 11535 246073
rect 11367 245037 11535 245296
rect 11367 244260 11377 245037
rect 11525 244260 11535 245037
rect 11367 244075 11535 244260
rect 11577 254490 11745 254737
rect 11577 253713 11587 254490
rect 11735 253713 11745 254490
rect 11577 253454 11745 253713
rect 11577 252677 11587 253454
rect 11735 252677 11745 253454
rect 11577 252418 11745 252677
rect 11577 251641 11587 252418
rect 11735 251641 11745 252418
rect 11577 251382 11745 251641
rect 11577 250605 11587 251382
rect 11735 250605 11745 251382
rect 11577 250346 11745 250605
rect 11577 249569 11587 250346
rect 11735 249569 11745 250346
rect 11577 249181 11745 249569
rect 11577 248404 11587 249181
rect 11735 248404 11745 249181
rect 11577 248145 11745 248404
rect 11577 247368 11587 248145
rect 11735 247368 11745 248145
rect 11577 247109 11745 247368
rect 11577 246332 11587 247109
rect 11735 246332 11745 247109
rect 11577 246073 11745 246332
rect 11577 245296 11587 246073
rect 11735 245296 11745 246073
rect 11577 245037 11745 245296
rect 11577 244260 11587 245037
rect 11735 244260 11745 245037
rect 11577 244248 11745 244260
rect 11787 254490 11955 254501
rect 11787 253713 11797 254490
rect 11945 253713 11955 254490
rect 11787 253454 11955 253713
rect 11787 252677 11797 253454
rect 11945 252677 11955 253454
rect 11787 252418 11955 252677
rect 11787 251641 11797 252418
rect 11945 251641 11955 252418
rect 11787 251382 11955 251641
rect 11787 250605 11797 251382
rect 11945 250605 11955 251382
rect 11787 250346 11955 250605
rect 11787 249569 11797 250346
rect 11945 249569 11955 250346
rect 11787 249181 11955 249569
rect 11787 248404 11797 249181
rect 11945 248404 11955 249181
rect 11787 248145 11955 248404
rect 11787 247368 11797 248145
rect 11945 247368 11955 248145
rect 11787 247109 11955 247368
rect 11787 246332 11797 247109
rect 11945 246332 11955 247109
rect 11787 246073 11955 246332
rect 11787 245296 11797 246073
rect 11945 245296 11955 246073
rect 11787 245037 11955 245296
rect 11787 244260 11797 245037
rect 11945 244260 11955 245037
rect 11787 244075 11955 244260
rect 11997 254490 12165 254737
rect 11997 253713 12007 254490
rect 12155 253713 12165 254490
rect 11997 253454 12165 253713
rect 11997 252677 12007 253454
rect 12155 252677 12165 253454
rect 11997 252418 12165 252677
rect 11997 251641 12007 252418
rect 12155 251641 12165 252418
rect 11997 251382 12165 251641
rect 11997 250605 12007 251382
rect 12155 250605 12165 251382
rect 11997 250346 12165 250605
rect 11997 249569 12007 250346
rect 12155 249569 12165 250346
rect 11997 249181 12165 249569
rect 11997 248404 12007 249181
rect 12155 248404 12165 249181
rect 11997 248145 12165 248404
rect 11997 247368 12007 248145
rect 12155 247368 12165 248145
rect 11997 247109 12165 247368
rect 11997 246332 12007 247109
rect 12155 246332 12165 247109
rect 11997 246073 12165 246332
rect 11997 245296 12007 246073
rect 12155 245296 12165 246073
rect 11997 245037 12165 245296
rect 11997 244260 12007 245037
rect 12155 244260 12165 245037
rect 11997 244248 12165 244260
rect 12207 254490 12375 254501
rect 12207 253713 12217 254490
rect 12365 253713 12375 254490
rect 12207 253454 12375 253713
rect 12207 252677 12217 253454
rect 12365 252677 12375 253454
rect 12207 252418 12375 252677
rect 12207 251641 12217 252418
rect 12365 251641 12375 252418
rect 12207 251382 12375 251641
rect 12207 250605 12217 251382
rect 12365 250605 12375 251382
rect 12207 250346 12375 250605
rect 12207 249569 12217 250346
rect 12365 249569 12375 250346
rect 12207 249181 12375 249569
rect 12207 248404 12217 249181
rect 12365 248404 12375 249181
rect 12207 248145 12375 248404
rect 12207 247368 12217 248145
rect 12365 247368 12375 248145
rect 12207 247109 12375 247368
rect 12207 246332 12217 247109
rect 12365 246332 12375 247109
rect 12207 246073 12375 246332
rect 12207 245296 12217 246073
rect 12365 245296 12375 246073
rect 12207 245037 12375 245296
rect 12207 244260 12217 245037
rect 12365 244260 12375 245037
rect 12207 244075 12375 244260
rect 12417 254490 12585 254737
rect 12417 253713 12427 254490
rect 12575 253713 12585 254490
rect 12417 253454 12585 253713
rect 12417 252677 12427 253454
rect 12575 252677 12585 253454
rect 12417 252418 12585 252677
rect 12417 251641 12427 252418
rect 12575 251641 12585 252418
rect 12417 251382 12585 251641
rect 12417 250605 12427 251382
rect 12575 250605 12585 251382
rect 12417 250346 12585 250605
rect 12417 249569 12427 250346
rect 12575 249569 12585 250346
rect 12417 249181 12585 249569
rect 12417 248404 12427 249181
rect 12575 248404 12585 249181
rect 12417 248145 12585 248404
rect 12417 247368 12427 248145
rect 12575 247368 12585 248145
rect 12417 247109 12585 247368
rect 12417 246332 12427 247109
rect 12575 246332 12585 247109
rect 12417 246073 12585 246332
rect 12417 245296 12427 246073
rect 12575 245296 12585 246073
rect 12417 245037 12585 245296
rect 12417 244260 12427 245037
rect 12575 244260 12585 245037
rect 12417 244248 12585 244260
rect 12627 254490 12795 254501
rect 12627 253713 12637 254490
rect 12785 253713 12795 254490
rect 12627 253454 12795 253713
rect 12627 252677 12637 253454
rect 12785 252677 12795 253454
rect 12627 252418 12795 252677
rect 12627 251641 12637 252418
rect 12785 251641 12795 252418
rect 12627 251382 12795 251641
rect 12627 250605 12637 251382
rect 12785 250605 12795 251382
rect 12627 250346 12795 250605
rect 12627 249569 12637 250346
rect 12785 249569 12795 250346
rect 12627 249181 12795 249569
rect 12627 248404 12637 249181
rect 12785 248404 12795 249181
rect 12627 248145 12795 248404
rect 12627 247368 12637 248145
rect 12785 247368 12795 248145
rect 12627 247109 12795 247368
rect 12627 246332 12637 247109
rect 12785 246332 12795 247109
rect 12627 246073 12795 246332
rect 12627 245296 12637 246073
rect 12785 245296 12795 246073
rect 12627 245037 12795 245296
rect 12627 244260 12637 245037
rect 12785 244260 12795 245037
rect 12627 244075 12795 244260
rect 12837 254490 13005 254737
rect 12837 253713 12847 254490
rect 12995 253713 13005 254490
rect 12837 253454 13005 253713
rect 12837 252677 12847 253454
rect 12995 252677 13005 253454
rect 12837 252418 13005 252677
rect 12837 251641 12847 252418
rect 12995 251641 13005 252418
rect 12837 251382 13005 251641
rect 12837 250605 12847 251382
rect 12995 250605 13005 251382
rect 12837 250346 13005 250605
rect 12837 249569 12847 250346
rect 12995 249569 13005 250346
rect 12837 249181 13005 249569
rect 12837 248404 12847 249181
rect 12995 248404 13005 249181
rect 12837 248145 13005 248404
rect 12837 247368 12847 248145
rect 12995 247368 13005 248145
rect 12837 247109 13005 247368
rect 12837 246332 12847 247109
rect 12995 246332 13005 247109
rect 12837 246073 13005 246332
rect 12837 245296 12847 246073
rect 12995 245296 13005 246073
rect 12837 245037 13005 245296
rect 12837 244260 12847 245037
rect 12995 244260 13005 245037
rect 12837 244248 13005 244260
rect 13047 254490 13215 254501
rect 13047 253713 13057 254490
rect 13205 253713 13215 254490
rect 13047 253454 13215 253713
rect 13047 252677 13057 253454
rect 13205 252677 13215 253454
rect 13047 252418 13215 252677
rect 13047 251641 13057 252418
rect 13205 251641 13215 252418
rect 13047 251382 13215 251641
rect 13047 250605 13057 251382
rect 13205 250605 13215 251382
rect 13047 250346 13215 250605
rect 13047 249569 13057 250346
rect 13205 249569 13215 250346
rect 13047 249181 13215 249569
rect 13047 248404 13057 249181
rect 13205 248404 13215 249181
rect 13047 248145 13215 248404
rect 13047 247368 13057 248145
rect 13205 247368 13215 248145
rect 13047 247109 13215 247368
rect 13047 246332 13057 247109
rect 13205 246332 13215 247109
rect 13047 246073 13215 246332
rect 13047 245296 13057 246073
rect 13205 245296 13215 246073
rect 13047 245037 13215 245296
rect 13047 244260 13057 245037
rect 13205 244260 13215 245037
rect 13047 244075 13215 244260
rect 13257 254490 13425 254737
rect 13257 253713 13267 254490
rect 13415 253713 13425 254490
rect 13257 253454 13425 253713
rect 13257 252677 13267 253454
rect 13415 252677 13425 253454
rect 13257 252418 13425 252677
rect 13257 251641 13267 252418
rect 13415 251641 13425 252418
rect 13257 251382 13425 251641
rect 13257 250605 13267 251382
rect 13415 250605 13425 251382
rect 13257 250346 13425 250605
rect 13257 249569 13267 250346
rect 13415 249569 13425 250346
rect 13257 249181 13425 249569
rect 13257 248404 13267 249181
rect 13415 248404 13425 249181
rect 13257 248145 13425 248404
rect 13257 247368 13267 248145
rect 13415 247368 13425 248145
rect 13257 247109 13425 247368
rect 13257 246332 13267 247109
rect 13415 246332 13425 247109
rect 13257 246073 13425 246332
rect 13257 245296 13267 246073
rect 13415 245296 13425 246073
rect 13257 245037 13425 245296
rect 13257 244260 13267 245037
rect 13415 244260 13425 245037
rect 13257 244248 13425 244260
rect 13467 254490 13635 254501
rect 13467 253713 13477 254490
rect 13625 253713 13635 254490
rect 13467 253454 13635 253713
rect 13467 252677 13477 253454
rect 13625 252677 13635 253454
rect 13467 252418 13635 252677
rect 13467 251641 13477 252418
rect 13625 251641 13635 252418
rect 13467 251382 13635 251641
rect 13467 250605 13477 251382
rect 13625 250605 13635 251382
rect 13467 250346 13635 250605
rect 13467 249569 13477 250346
rect 13625 249569 13635 250346
rect 13467 249181 13635 249569
rect 13467 248404 13477 249181
rect 13625 248404 13635 249181
rect 13467 248145 13635 248404
rect 13467 247368 13477 248145
rect 13625 247368 13635 248145
rect 13467 247109 13635 247368
rect 13467 246332 13477 247109
rect 13625 246332 13635 247109
rect 13467 246073 13635 246332
rect 13467 245296 13477 246073
rect 13625 245296 13635 246073
rect 13467 245037 13635 245296
rect 13467 244260 13477 245037
rect 13625 244260 13635 245037
rect 13467 244075 13635 244260
rect 13677 254490 13845 254737
rect 13677 253713 13687 254490
rect 13835 253713 13845 254490
rect 13677 253454 13845 253713
rect 13677 252677 13687 253454
rect 13835 252677 13845 253454
rect 13677 252418 13845 252677
rect 13677 251641 13687 252418
rect 13835 251641 13845 252418
rect 13677 251382 13845 251641
rect 13677 250605 13687 251382
rect 13835 250605 13845 251382
rect 13677 250346 13845 250605
rect 13677 249569 13687 250346
rect 13835 249569 13845 250346
rect 13677 249181 13845 249569
rect 13677 248404 13687 249181
rect 13835 248404 13845 249181
rect 13677 248145 13845 248404
rect 13677 247368 13687 248145
rect 13835 247368 13845 248145
rect 13677 247109 13845 247368
rect 13677 246332 13687 247109
rect 13835 246332 13845 247109
rect 13677 246073 13845 246332
rect 13677 245296 13687 246073
rect 13835 245296 13845 246073
rect 13677 245037 13845 245296
rect 13677 244260 13687 245037
rect 13835 244260 13845 245037
rect 13677 244248 13845 244260
rect 13887 254490 14055 254501
rect 13887 253713 13897 254490
rect 14045 253713 14055 254490
rect 13887 253454 14055 253713
rect 13887 252677 13897 253454
rect 14045 252677 14055 253454
rect 13887 252418 14055 252677
rect 13887 251641 13897 252418
rect 14045 251641 14055 252418
rect 13887 251382 14055 251641
rect 13887 250605 13897 251382
rect 14045 250605 14055 251382
rect 13887 250346 14055 250605
rect 13887 249569 13897 250346
rect 14045 249569 14055 250346
rect 13887 249181 14055 249569
rect 13887 248404 13897 249181
rect 14045 248404 14055 249181
rect 13887 248145 14055 248404
rect 13887 247368 13897 248145
rect 14045 247368 14055 248145
rect 13887 247109 14055 247368
rect 13887 246332 13897 247109
rect 14045 246332 14055 247109
rect 13887 246073 14055 246332
rect 13887 245296 13897 246073
rect 14045 245296 14055 246073
rect 13887 245037 14055 245296
rect 13887 244260 13897 245037
rect 14045 244260 14055 245037
rect 13887 244075 14055 244260
rect 14097 254490 14265 254737
rect 14097 253713 14107 254490
rect 14255 253713 14265 254490
rect 14097 253454 14265 253713
rect 14097 252677 14107 253454
rect 14255 252677 14265 253454
rect 14097 252418 14265 252677
rect 14097 251641 14107 252418
rect 14255 251641 14265 252418
rect 14097 251382 14265 251641
rect 14097 250605 14107 251382
rect 14255 250605 14265 251382
rect 14097 250346 14265 250605
rect 14097 249569 14107 250346
rect 14255 249569 14265 250346
rect 14097 249181 14265 249569
rect 14097 248404 14107 249181
rect 14255 248404 14265 249181
rect 14097 248145 14265 248404
rect 14097 247368 14107 248145
rect 14255 247368 14265 248145
rect 14097 247109 14265 247368
rect 14097 246332 14107 247109
rect 14255 246332 14265 247109
rect 14097 246073 14265 246332
rect 14097 245296 14107 246073
rect 14255 245296 14265 246073
rect 14097 245037 14265 245296
rect 14097 244260 14107 245037
rect 14255 244260 14265 245037
rect 14097 244248 14265 244260
rect 14307 254490 14475 254501
rect 14307 253713 14317 254490
rect 14465 253713 14475 254490
rect 14307 253454 14475 253713
rect 14307 252677 14317 253454
rect 14465 252677 14475 253454
rect 14307 252418 14475 252677
rect 14307 251641 14317 252418
rect 14465 251641 14475 252418
rect 14307 251382 14475 251641
rect 14307 250605 14317 251382
rect 14465 250605 14475 251382
rect 14307 250346 14475 250605
rect 14307 249569 14317 250346
rect 14465 249569 14475 250346
rect 14307 249181 14475 249569
rect 14307 248404 14317 249181
rect 14465 248404 14475 249181
rect 14307 248145 14475 248404
rect 14307 247368 14317 248145
rect 14465 247368 14475 248145
rect 14307 247109 14475 247368
rect 14307 246332 14317 247109
rect 14465 246332 14475 247109
rect 14307 246073 14475 246332
rect 14307 245296 14317 246073
rect 14465 245296 14475 246073
rect 14307 245037 14475 245296
rect 14307 244260 14317 245037
rect 14465 244260 14475 245037
rect 14307 244075 14475 244260
rect 14517 254490 14685 254737
rect 14517 253713 14527 254490
rect 14675 253713 14685 254490
rect 14517 253454 14685 253713
rect 14517 252677 14527 253454
rect 14675 252677 14685 253454
rect 14517 252418 14685 252677
rect 14517 251641 14527 252418
rect 14675 251641 14685 252418
rect 14517 251382 14685 251641
rect 14517 250605 14527 251382
rect 14675 250605 14685 251382
rect 14517 250346 14685 250605
rect 14517 249569 14527 250346
rect 14675 249569 14685 250346
rect 14517 249181 14685 249569
rect 14517 248404 14527 249181
rect 14675 248404 14685 249181
rect 14517 248145 14685 248404
rect 14517 247368 14527 248145
rect 14675 247368 14685 248145
rect 14517 247109 14685 247368
rect 14517 246332 14527 247109
rect 14675 246332 14685 247109
rect 14517 246073 14685 246332
rect 14517 245296 14527 246073
rect 14675 245296 14685 246073
rect 14517 245037 14685 245296
rect 14517 244260 14527 245037
rect 14675 244260 14685 245037
rect 14517 244248 14685 244260
rect 14727 254490 14895 254501
rect 14727 253713 14737 254490
rect 14885 253713 14895 254490
rect 14727 253454 14895 253713
rect 14727 252677 14737 253454
rect 14885 252677 14895 253454
rect 14727 252418 14895 252677
rect 14727 251641 14737 252418
rect 14885 251641 14895 252418
rect 14727 251382 14895 251641
rect 14727 250605 14737 251382
rect 14885 250605 14895 251382
rect 14727 250346 14895 250605
rect 14727 249569 14737 250346
rect 14885 249569 14895 250346
rect 14727 249181 14895 249569
rect 14727 248404 14737 249181
rect 14885 248404 14895 249181
rect 14727 248145 14895 248404
rect 14727 247368 14737 248145
rect 14885 247368 14895 248145
rect 14727 247109 14895 247368
rect 14727 246332 14737 247109
rect 14885 246332 14895 247109
rect 14727 246073 14895 246332
rect 14727 245296 14737 246073
rect 14885 245296 14895 246073
rect 14727 245037 14895 245296
rect 14727 244260 14737 245037
rect 14885 244260 14895 245037
rect 14727 244075 14895 244260
rect 14937 254490 15105 254737
rect 14937 253713 14947 254490
rect 15095 253713 15105 254490
rect 14937 253454 15105 253713
rect 14937 252677 14947 253454
rect 15095 252677 15105 253454
rect 14937 252418 15105 252677
rect 14937 251641 14947 252418
rect 15095 251641 15105 252418
rect 14937 251382 15105 251641
rect 14937 250605 14947 251382
rect 15095 250605 15105 251382
rect 14937 250346 15105 250605
rect 14937 249569 14947 250346
rect 15095 249569 15105 250346
rect 14937 249181 15105 249569
rect 14937 248404 14947 249181
rect 15095 248404 15105 249181
rect 14937 248145 15105 248404
rect 14937 247368 14947 248145
rect 15095 247368 15105 248145
rect 14937 247109 15105 247368
rect 14937 246332 14947 247109
rect 15095 246332 15105 247109
rect 14937 246073 15105 246332
rect 14937 245296 14947 246073
rect 15095 245296 15105 246073
rect 14937 245037 15105 245296
rect 14937 244260 14947 245037
rect 15095 244260 15105 245037
rect 14937 244248 15105 244260
rect 15147 254490 15315 254501
rect 15147 253713 15157 254490
rect 15305 253713 15315 254490
rect 15147 253454 15315 253713
rect 15147 252677 15157 253454
rect 15305 252677 15315 253454
rect 15147 252418 15315 252677
rect 15147 251641 15157 252418
rect 15305 251641 15315 252418
rect 15147 251382 15315 251641
rect 15147 250605 15157 251382
rect 15305 250605 15315 251382
rect 15147 250346 15315 250605
rect 15147 249569 15157 250346
rect 15305 249569 15315 250346
rect 15147 249181 15315 249569
rect 15147 248404 15157 249181
rect 15305 248404 15315 249181
rect 15147 248145 15315 248404
rect 15147 247368 15157 248145
rect 15305 247368 15315 248145
rect 15147 247109 15315 247368
rect 15147 246332 15157 247109
rect 15305 246332 15315 247109
rect 15147 246073 15315 246332
rect 15147 245296 15157 246073
rect 15305 245296 15315 246073
rect 15147 245037 15315 245296
rect 15147 244260 15157 245037
rect 15305 244260 15315 245037
rect 15147 244075 15315 244260
rect 15357 254490 15525 254737
rect 15357 253713 15367 254490
rect 15515 253713 15525 254490
rect 15357 253454 15525 253713
rect 15357 252677 15367 253454
rect 15515 252677 15525 253454
rect 15357 252418 15525 252677
rect 15357 251641 15367 252418
rect 15515 251641 15525 252418
rect 15357 251382 15525 251641
rect 15357 250605 15367 251382
rect 15515 250605 15525 251382
rect 15357 250346 15525 250605
rect 15357 249569 15367 250346
rect 15515 249569 15525 250346
rect 15357 249181 15525 249569
rect 15357 248404 15367 249181
rect 15515 248404 15525 249181
rect 15357 248145 15525 248404
rect 15357 247368 15367 248145
rect 15515 247368 15525 248145
rect 15357 247109 15525 247368
rect 15357 246332 15367 247109
rect 15515 246332 15525 247109
rect 15357 246073 15525 246332
rect 15357 245296 15367 246073
rect 15515 245296 15525 246073
rect 15357 245037 15525 245296
rect 15357 244260 15367 245037
rect 15515 244260 15525 245037
rect 15357 244248 15525 244260
rect 15567 254490 15735 254501
rect 15567 253713 15577 254490
rect 15725 253713 15735 254490
rect 15567 253454 15735 253713
rect 15567 252677 15577 253454
rect 15725 252677 15735 253454
rect 15567 252418 15735 252677
rect 15567 251641 15577 252418
rect 15725 251641 15735 252418
rect 15567 251382 15735 251641
rect 15567 250605 15577 251382
rect 15725 250605 15735 251382
rect 15567 250346 15735 250605
rect 15567 249569 15577 250346
rect 15725 249569 15735 250346
rect 15567 249181 15735 249569
rect 15567 248404 15577 249181
rect 15725 248404 15735 249181
rect 15567 248145 15735 248404
rect 15567 247368 15577 248145
rect 15725 247368 15735 248145
rect 15567 247109 15735 247368
rect 15567 246332 15577 247109
rect 15725 246332 15735 247109
rect 15567 246073 15735 246332
rect 15567 245296 15577 246073
rect 15725 245296 15735 246073
rect 15567 245037 15735 245296
rect 15567 244260 15577 245037
rect 15725 244260 15735 245037
rect 15567 244075 15735 244260
rect 15777 254490 15945 254737
rect 15777 253713 15787 254490
rect 15935 253713 15945 254490
rect 15777 253454 15945 253713
rect 15777 252677 15787 253454
rect 15935 252677 15945 253454
rect 15777 252418 15945 252677
rect 15777 251641 15787 252418
rect 15935 251641 15945 252418
rect 15777 251382 15945 251641
rect 15777 250605 15787 251382
rect 15935 250605 15945 251382
rect 15777 250346 15945 250605
rect 15777 249569 15787 250346
rect 15935 249569 15945 250346
rect 15777 249181 15945 249569
rect 15777 248404 15787 249181
rect 15935 248404 15945 249181
rect 15777 248145 15945 248404
rect 15777 247368 15787 248145
rect 15935 247368 15945 248145
rect 15777 247109 15945 247368
rect 15777 246332 15787 247109
rect 15935 246332 15945 247109
rect 15777 246073 15945 246332
rect 15777 245296 15787 246073
rect 15935 245296 15945 246073
rect 15777 245037 15945 245296
rect 15777 244260 15787 245037
rect 15935 244260 15945 245037
rect 15777 244248 15945 244260
rect 15987 254490 16155 254501
rect 15987 253713 15997 254490
rect 16145 253713 16155 254490
rect 15987 253454 16155 253713
rect 15987 252677 15997 253454
rect 16145 252677 16155 253454
rect 15987 252418 16155 252677
rect 15987 251641 15997 252418
rect 16145 251641 16155 252418
rect 15987 251382 16155 251641
rect 15987 250605 15997 251382
rect 16145 250605 16155 251382
rect 15987 250346 16155 250605
rect 15987 249569 15997 250346
rect 16145 249569 16155 250346
rect 15987 249181 16155 249569
rect 15987 248404 15997 249181
rect 16145 248404 16155 249181
rect 15987 248145 16155 248404
rect 15987 247368 15997 248145
rect 16145 247368 16155 248145
rect 15987 247109 16155 247368
rect 15987 246332 15997 247109
rect 16145 246332 16155 247109
rect 15987 246073 16155 246332
rect 15987 245296 15997 246073
rect 16145 245296 16155 246073
rect 15987 245037 16155 245296
rect 15987 244260 15997 245037
rect 16145 244260 16155 245037
rect 15987 244075 16155 244260
rect 16197 254490 16365 254737
rect 16197 253713 16207 254490
rect 16355 253713 16365 254490
rect 16197 253454 16365 253713
rect 16197 252677 16207 253454
rect 16355 252677 16365 253454
rect 16197 252418 16365 252677
rect 16197 251641 16207 252418
rect 16355 251641 16365 252418
rect 16197 251382 16365 251641
rect 16197 250605 16207 251382
rect 16355 250605 16365 251382
rect 16197 250346 16365 250605
rect 16197 249569 16207 250346
rect 16355 249569 16365 250346
rect 16197 249181 16365 249569
rect 16197 248404 16207 249181
rect 16355 248404 16365 249181
rect 16197 248145 16365 248404
rect 16197 247368 16207 248145
rect 16355 247368 16365 248145
rect 16197 247109 16365 247368
rect 16197 246332 16207 247109
rect 16355 246332 16365 247109
rect 16197 246073 16365 246332
rect 16197 245296 16207 246073
rect 16355 245296 16365 246073
rect 16197 245037 16365 245296
rect 16197 244260 16207 245037
rect 16355 244260 16365 245037
rect 16197 244248 16365 244260
rect 16407 254490 16575 254501
rect 16407 253713 16417 254490
rect 16565 253713 16575 254490
rect 16407 253454 16575 253713
rect 16407 252677 16417 253454
rect 16565 252677 16575 253454
rect 16407 252418 16575 252677
rect 16407 251641 16417 252418
rect 16565 251641 16575 252418
rect 16407 251382 16575 251641
rect 16407 250605 16417 251382
rect 16565 250605 16575 251382
rect 16407 250346 16575 250605
rect 16407 249569 16417 250346
rect 16565 249569 16575 250346
rect 16407 249181 16575 249569
rect 16407 248404 16417 249181
rect 16565 248404 16575 249181
rect 16407 248145 16575 248404
rect 16407 247368 16417 248145
rect 16565 247368 16575 248145
rect 16407 247109 16575 247368
rect 16407 246332 16417 247109
rect 16565 246332 16575 247109
rect 16407 246073 16575 246332
rect 16407 245296 16417 246073
rect 16565 245296 16575 246073
rect 16407 245037 16575 245296
rect 16407 244260 16417 245037
rect 16565 244260 16575 245037
rect 16407 244075 16575 244260
rect 16617 254490 16785 254737
rect 16617 253713 16627 254490
rect 16775 253713 16785 254490
rect 16617 253454 16785 253713
rect 16617 252677 16627 253454
rect 16775 252677 16785 253454
rect 16617 252418 16785 252677
rect 16617 251641 16627 252418
rect 16775 251641 16785 252418
rect 16617 251382 16785 251641
rect 16617 250605 16627 251382
rect 16775 250605 16785 251382
rect 16617 250346 16785 250605
rect 16617 249569 16627 250346
rect 16775 249569 16785 250346
rect 16617 249181 16785 249569
rect 16617 248404 16627 249181
rect 16775 248404 16785 249181
rect 16617 248145 16785 248404
rect 16617 247368 16627 248145
rect 16775 247368 16785 248145
rect 16617 247109 16785 247368
rect 16617 246332 16627 247109
rect 16775 246332 16785 247109
rect 16617 246073 16785 246332
rect 16617 245296 16627 246073
rect 16775 245296 16785 246073
rect 16617 245037 16785 245296
rect 16617 244260 16627 245037
rect 16775 244260 16785 245037
rect 16617 244248 16785 244260
rect 16827 254490 16995 254501
rect 16827 253713 16837 254490
rect 16985 253713 16995 254490
rect 16827 253454 16995 253713
rect 16827 252677 16837 253454
rect 16985 252677 16995 253454
rect 16827 252418 16995 252677
rect 16827 251641 16837 252418
rect 16985 251641 16995 252418
rect 16827 251382 16995 251641
rect 16827 250605 16837 251382
rect 16985 250605 16995 251382
rect 16827 250346 16995 250605
rect 16827 249569 16837 250346
rect 16985 249569 16995 250346
rect 16827 249181 16995 249569
rect 16827 248404 16837 249181
rect 16985 248404 16995 249181
rect 16827 248145 16995 248404
rect 16827 247368 16837 248145
rect 16985 247368 16995 248145
rect 16827 247109 16995 247368
rect 16827 246332 16837 247109
rect 16985 246332 16995 247109
rect 16827 246073 16995 246332
rect 16827 245296 16837 246073
rect 16985 245296 16995 246073
rect 16827 245037 16995 245296
rect 16827 244260 16837 245037
rect 16985 244260 16995 245037
rect 16827 244075 16995 244260
rect 17037 254490 17205 254737
rect 17037 253713 17047 254490
rect 17195 253713 17205 254490
rect 17037 253454 17205 253713
rect 17037 252677 17047 253454
rect 17195 252677 17205 253454
rect 17037 252418 17205 252677
rect 17037 251641 17047 252418
rect 17195 251641 17205 252418
rect 17037 251382 17205 251641
rect 17037 250605 17047 251382
rect 17195 250605 17205 251382
rect 17037 250346 17205 250605
rect 17037 249569 17047 250346
rect 17195 249569 17205 250346
rect 17037 249181 17205 249569
rect 17037 248404 17047 249181
rect 17195 248404 17205 249181
rect 17037 248145 17205 248404
rect 17037 247368 17047 248145
rect 17195 247368 17205 248145
rect 17037 247109 17205 247368
rect 17037 246332 17047 247109
rect 17195 246332 17205 247109
rect 17037 246073 17205 246332
rect 17037 245296 17047 246073
rect 17195 245296 17205 246073
rect 17037 245037 17205 245296
rect 17037 244260 17047 245037
rect 17195 244260 17205 245037
rect 17037 244248 17205 244260
rect 17247 254490 17415 254501
rect 17247 253713 17257 254490
rect 17405 253713 17415 254490
rect 17247 253454 17415 253713
rect 17247 252677 17257 253454
rect 17405 252677 17415 253454
rect 17247 252418 17415 252677
rect 17247 251641 17257 252418
rect 17405 251641 17415 252418
rect 17247 251382 17415 251641
rect 17247 250605 17257 251382
rect 17405 250605 17415 251382
rect 17247 250346 17415 250605
rect 17247 249569 17257 250346
rect 17405 249569 17415 250346
rect 17247 249181 17415 249569
rect 17247 248404 17257 249181
rect 17405 248404 17415 249181
rect 17247 248145 17415 248404
rect 17247 247368 17257 248145
rect 17405 247368 17415 248145
rect 17247 247109 17415 247368
rect 17247 246332 17257 247109
rect 17405 246332 17415 247109
rect 17247 246073 17415 246332
rect 17247 245296 17257 246073
rect 17405 245296 17415 246073
rect 17247 245037 17415 245296
rect 17247 244260 17257 245037
rect 17405 244260 17415 245037
rect 17247 244075 17415 244260
rect 17457 254490 17625 254737
rect 17457 253713 17467 254490
rect 17615 253713 17625 254490
rect 17457 253454 17625 253713
rect 17457 252677 17467 253454
rect 17615 252677 17625 253454
rect 17457 252418 17625 252677
rect 17457 251641 17467 252418
rect 17615 251641 17625 252418
rect 17457 251382 17625 251641
rect 17457 250605 17467 251382
rect 17615 250605 17625 251382
rect 17457 250346 17625 250605
rect 17457 249569 17467 250346
rect 17615 249569 17625 250346
rect 17457 249181 17625 249569
rect 17457 248404 17467 249181
rect 17615 248404 17625 249181
rect 17457 248145 17625 248404
rect 17457 247368 17467 248145
rect 17615 247368 17625 248145
rect 17457 247109 17625 247368
rect 17457 246332 17467 247109
rect 17615 246332 17625 247109
rect 17457 246073 17625 246332
rect 17457 245296 17467 246073
rect 17615 245296 17625 246073
rect 17457 245037 17625 245296
rect 17457 244260 17467 245037
rect 17615 244260 17625 245037
rect 17457 244248 17625 244260
rect 17667 254490 17835 254501
rect 17667 253713 17677 254490
rect 17825 253713 17835 254490
rect 17667 253454 17835 253713
rect 17667 252677 17677 253454
rect 17825 252677 17835 253454
rect 17667 252418 17835 252677
rect 17667 251641 17677 252418
rect 17825 251641 17835 252418
rect 17667 251382 17835 251641
rect 17667 250605 17677 251382
rect 17825 250605 17835 251382
rect 17667 250346 17835 250605
rect 17667 249569 17677 250346
rect 17825 249569 17835 250346
rect 17667 249181 17835 249569
rect 17667 248404 17677 249181
rect 17825 248404 17835 249181
rect 17667 248145 17835 248404
rect 17667 247368 17677 248145
rect 17825 247368 17835 248145
rect 17667 247109 17835 247368
rect 17667 246332 17677 247109
rect 17825 246332 17835 247109
rect 17667 246073 17835 246332
rect 17667 245296 17677 246073
rect 17825 245296 17835 246073
rect 17667 245037 17835 245296
rect 17667 244260 17677 245037
rect 17825 244260 17835 245037
rect 17667 244075 17835 244260
rect 17877 254490 18045 254737
rect 17877 253713 17887 254490
rect 18035 253713 18045 254490
rect 17877 253454 18045 253713
rect 17877 252677 17887 253454
rect 18035 252677 18045 253454
rect 17877 252418 18045 252677
rect 17877 251641 17887 252418
rect 18035 251641 18045 252418
rect 17877 251382 18045 251641
rect 17877 250605 17887 251382
rect 18035 250605 18045 251382
rect 17877 250346 18045 250605
rect 17877 249569 17887 250346
rect 18035 249569 18045 250346
rect 17877 249181 18045 249569
rect 17877 248404 17887 249181
rect 18035 248404 18045 249181
rect 17877 248145 18045 248404
rect 17877 247368 17887 248145
rect 18035 247368 18045 248145
rect 17877 247109 18045 247368
rect 17877 246332 17887 247109
rect 18035 246332 18045 247109
rect 17877 246073 18045 246332
rect 17877 245296 17887 246073
rect 18035 245296 18045 246073
rect 17877 245037 18045 245296
rect 17877 244260 17887 245037
rect 18035 244260 18045 245037
rect 17877 244248 18045 244260
rect 18087 254490 18255 254501
rect 18087 253713 18097 254490
rect 18245 253713 18255 254490
rect 18087 253454 18255 253713
rect 18087 252677 18097 253454
rect 18245 252677 18255 253454
rect 18087 252418 18255 252677
rect 18087 251641 18097 252418
rect 18245 251641 18255 252418
rect 18087 251382 18255 251641
rect 18087 250605 18097 251382
rect 18245 250605 18255 251382
rect 18087 250346 18255 250605
rect 18087 249569 18097 250346
rect 18245 249569 18255 250346
rect 18087 249181 18255 249569
rect 18087 248404 18097 249181
rect 18245 248404 18255 249181
rect 18087 248145 18255 248404
rect 18087 247368 18097 248145
rect 18245 247368 18255 248145
rect 18087 247109 18255 247368
rect 18087 246332 18097 247109
rect 18245 246332 18255 247109
rect 18087 246073 18255 246332
rect 18087 245296 18097 246073
rect 18245 245296 18255 246073
rect 18087 245037 18255 245296
rect 18087 244260 18097 245037
rect 18245 244260 18255 245037
rect 18087 244075 18255 244260
rect 18297 254490 18465 254737
rect 18297 253713 18307 254490
rect 18455 253713 18465 254490
rect 18297 253454 18465 253713
rect 18297 252677 18307 253454
rect 18455 252677 18465 253454
rect 18297 252418 18465 252677
rect 18297 251641 18307 252418
rect 18455 251641 18465 252418
rect 18297 251382 18465 251641
rect 18297 250605 18307 251382
rect 18455 250605 18465 251382
rect 18297 250346 18465 250605
rect 18297 249569 18307 250346
rect 18455 249569 18465 250346
rect 18297 249181 18465 249569
rect 18297 248404 18307 249181
rect 18455 248404 18465 249181
rect 18297 248145 18465 248404
rect 18297 247368 18307 248145
rect 18455 247368 18465 248145
rect 18297 247109 18465 247368
rect 18297 246332 18307 247109
rect 18455 246332 18465 247109
rect 18297 246073 18465 246332
rect 18297 245296 18307 246073
rect 18455 245296 18465 246073
rect 18297 245037 18465 245296
rect 18297 244260 18307 245037
rect 18455 244260 18465 245037
rect 18297 244248 18465 244260
rect 18507 254490 18675 254501
rect 18507 253713 18517 254490
rect 18665 253713 18675 254490
rect 18507 253454 18675 253713
rect 18507 252677 18517 253454
rect 18665 252677 18675 253454
rect 18507 252418 18675 252677
rect 18507 251641 18517 252418
rect 18665 251641 18675 252418
rect 18507 251382 18675 251641
rect 18507 250605 18517 251382
rect 18665 250605 18675 251382
rect 18507 250346 18675 250605
rect 18507 249569 18517 250346
rect 18665 249569 18675 250346
rect 18507 249181 18675 249569
rect 18507 248404 18517 249181
rect 18665 248404 18675 249181
rect 18507 248145 18675 248404
rect 18507 247368 18517 248145
rect 18665 247368 18675 248145
rect 18507 247109 18675 247368
rect 18507 246332 18517 247109
rect 18665 246332 18675 247109
rect 18507 246073 18675 246332
rect 18507 245296 18517 246073
rect 18665 245296 18675 246073
rect 18507 245037 18675 245296
rect 18507 244260 18517 245037
rect 18665 244260 18675 245037
rect 18507 244075 18675 244260
rect 18717 254490 18885 254737
rect 18717 253713 18727 254490
rect 18875 253713 18885 254490
rect 18717 253454 18885 253713
rect 18717 252677 18727 253454
rect 18875 252677 18885 253454
rect 18717 252418 18885 252677
rect 18717 251641 18727 252418
rect 18875 251641 18885 252418
rect 18717 251382 18885 251641
rect 18717 250605 18727 251382
rect 18875 250605 18885 251382
rect 18717 250346 18885 250605
rect 18717 249569 18727 250346
rect 18875 249569 18885 250346
rect 18717 249181 18885 249569
rect 18717 248404 18727 249181
rect 18875 248404 18885 249181
rect 18717 248145 18885 248404
rect 18717 247368 18727 248145
rect 18875 247368 18885 248145
rect 18717 247109 18885 247368
rect 18717 246332 18727 247109
rect 18875 246332 18885 247109
rect 18717 246073 18885 246332
rect 18717 245296 18727 246073
rect 18875 245296 18885 246073
rect 18717 245037 18885 245296
rect 18717 244260 18727 245037
rect 18875 244260 18885 245037
rect 18717 244248 18885 244260
rect 18927 254490 19095 254501
rect 18927 253713 18937 254490
rect 19085 253713 19095 254490
rect 18927 253454 19095 253713
rect 18927 252677 18937 253454
rect 19085 252677 19095 253454
rect 18927 252418 19095 252677
rect 18927 251641 18937 252418
rect 19085 251641 19095 252418
rect 18927 251382 19095 251641
rect 18927 250605 18937 251382
rect 19085 250605 19095 251382
rect 18927 250346 19095 250605
rect 18927 249569 18937 250346
rect 19085 249569 19095 250346
rect 18927 249181 19095 249569
rect 18927 248404 18937 249181
rect 19085 248404 19095 249181
rect 18927 248145 19095 248404
rect 18927 247368 18937 248145
rect 19085 247368 19095 248145
rect 18927 247109 19095 247368
rect 18927 246332 18937 247109
rect 19085 246332 19095 247109
rect 18927 246073 19095 246332
rect 18927 245296 18937 246073
rect 19085 245296 19095 246073
rect 18927 245037 19095 245296
rect 18927 244260 18937 245037
rect 19085 244260 19095 245037
rect 18927 244075 19095 244260
rect 19137 254490 19305 254737
rect 19137 253713 19147 254490
rect 19295 253713 19305 254490
rect 19137 253454 19305 253713
rect 19137 252677 19147 253454
rect 19295 252677 19305 253454
rect 19137 252418 19305 252677
rect 19137 251641 19147 252418
rect 19295 251641 19305 252418
rect 19137 251382 19305 251641
rect 19137 250605 19147 251382
rect 19295 250605 19305 251382
rect 19137 250346 19305 250605
rect 19137 249569 19147 250346
rect 19295 249569 19305 250346
rect 19137 249181 19305 249569
rect 19137 248404 19147 249181
rect 19295 248404 19305 249181
rect 19137 248145 19305 248404
rect 19137 247368 19147 248145
rect 19295 247368 19305 248145
rect 19137 247109 19305 247368
rect 19137 246332 19147 247109
rect 19295 246332 19305 247109
rect 19137 246073 19305 246332
rect 19137 245296 19147 246073
rect 19295 245296 19305 246073
rect 19137 245037 19305 245296
rect 19137 244260 19147 245037
rect 19295 244260 19305 245037
rect 19137 244248 19305 244260
rect 19347 254490 19515 254501
rect 19347 253713 19357 254490
rect 19505 253713 19515 254490
rect 19347 253454 19515 253713
rect 19347 252677 19357 253454
rect 19505 252677 19515 253454
rect 19347 252418 19515 252677
rect 19347 251641 19357 252418
rect 19505 251641 19515 252418
rect 19347 251382 19515 251641
rect 19347 250605 19357 251382
rect 19505 250605 19515 251382
rect 19347 250346 19515 250605
rect 19347 249569 19357 250346
rect 19505 249569 19515 250346
rect 19347 249181 19515 249569
rect 19347 248404 19357 249181
rect 19505 248404 19515 249181
rect 19347 248145 19515 248404
rect 19347 247368 19357 248145
rect 19505 247368 19515 248145
rect 19347 247109 19515 247368
rect 19347 246332 19357 247109
rect 19505 246332 19515 247109
rect 19347 246073 19515 246332
rect 19347 245296 19357 246073
rect 19505 245296 19515 246073
rect 19347 245037 19515 245296
rect 19347 244260 19357 245037
rect 19505 244260 19515 245037
rect 19347 244075 19515 244260
rect 19557 254490 19725 254737
rect 19557 253713 19567 254490
rect 19715 253713 19725 254490
rect 19557 253454 19725 253713
rect 19557 252677 19567 253454
rect 19715 252677 19725 253454
rect 19557 252418 19725 252677
rect 19557 251641 19567 252418
rect 19715 251641 19725 252418
rect 19557 251382 19725 251641
rect 19557 250605 19567 251382
rect 19715 250605 19725 251382
rect 19557 250346 19725 250605
rect 19557 249569 19567 250346
rect 19715 249569 19725 250346
rect 19557 249181 19725 249569
rect 19557 248404 19567 249181
rect 19715 248404 19725 249181
rect 19557 248145 19725 248404
rect 19557 247368 19567 248145
rect 19715 247368 19725 248145
rect 19557 247109 19725 247368
rect 19557 246332 19567 247109
rect 19715 246332 19725 247109
rect 19557 246073 19725 246332
rect 19557 245296 19567 246073
rect 19715 245296 19725 246073
rect 19557 245037 19725 245296
rect 19557 244260 19567 245037
rect 19715 244260 19725 245037
rect 19557 244248 19725 244260
rect 19767 254490 19935 254501
rect 19767 253713 19777 254490
rect 19925 253713 19935 254490
rect 19767 253454 19935 253713
rect 19767 252677 19777 253454
rect 19925 252677 19935 253454
rect 19767 252418 19935 252677
rect 19767 251641 19777 252418
rect 19925 251641 19935 252418
rect 19767 251382 19935 251641
rect 19767 250605 19777 251382
rect 19925 250605 19935 251382
rect 19767 250346 19935 250605
rect 19767 249569 19777 250346
rect 19925 249569 19935 250346
rect 19767 249181 19935 249569
rect 19767 248404 19777 249181
rect 19925 248404 19935 249181
rect 19767 248145 19935 248404
rect 19767 247368 19777 248145
rect 19925 247368 19935 248145
rect 19767 247109 19935 247368
rect 19767 246332 19777 247109
rect 19925 246332 19935 247109
rect 19767 246073 19935 246332
rect 19767 245296 19777 246073
rect 19925 245296 19935 246073
rect 19767 245037 19935 245296
rect 19767 244260 19777 245037
rect 19925 244260 19935 245037
rect 19767 244075 19935 244260
rect 19977 254490 20145 254737
rect 19977 253713 19987 254490
rect 20135 253713 20145 254490
rect 19977 253454 20145 253713
rect 19977 252677 19987 253454
rect 20135 252677 20145 253454
rect 19977 252418 20145 252677
rect 19977 251641 19987 252418
rect 20135 251641 20145 252418
rect 19977 251382 20145 251641
rect 19977 250605 19987 251382
rect 20135 250605 20145 251382
rect 19977 250346 20145 250605
rect 19977 249569 19987 250346
rect 20135 249569 20145 250346
rect 19977 249181 20145 249569
rect 19977 248404 19987 249181
rect 20135 248404 20145 249181
rect 19977 248145 20145 248404
rect 19977 247368 19987 248145
rect 20135 247368 20145 248145
rect 19977 247109 20145 247368
rect 19977 246332 19987 247109
rect 20135 246332 20145 247109
rect 19977 246073 20145 246332
rect 19977 245296 19987 246073
rect 20135 245296 20145 246073
rect 19977 245037 20145 245296
rect 19977 244260 19987 245037
rect 20135 244260 20145 245037
rect 19977 244248 20145 244260
rect 20187 254490 20355 254501
rect 20187 253713 20197 254490
rect 20345 253713 20355 254490
rect 20187 253454 20355 253713
rect 20187 252677 20197 253454
rect 20345 252677 20355 253454
rect 20187 252418 20355 252677
rect 20187 251641 20197 252418
rect 20345 251641 20355 252418
rect 20187 251382 20355 251641
rect 20187 250605 20197 251382
rect 20345 250605 20355 251382
rect 20187 250346 20355 250605
rect 20187 249569 20197 250346
rect 20345 249569 20355 250346
rect 20187 249181 20355 249569
rect 20187 248404 20197 249181
rect 20345 248404 20355 249181
rect 20187 248145 20355 248404
rect 20187 247368 20197 248145
rect 20345 247368 20355 248145
rect 20187 247109 20355 247368
rect 20187 246332 20197 247109
rect 20345 246332 20355 247109
rect 20187 246073 20355 246332
rect 20187 245296 20197 246073
rect 20345 245296 20355 246073
rect 20187 245037 20355 245296
rect 20187 244260 20197 245037
rect 20345 244260 20355 245037
rect 20187 244075 20355 244260
rect 20397 254490 20565 254737
rect 20397 253713 20407 254490
rect 20555 253713 20565 254490
rect 20397 253454 20565 253713
rect 20397 252677 20407 253454
rect 20555 252677 20565 253454
rect 20397 252418 20565 252677
rect 20397 251641 20407 252418
rect 20555 251641 20565 252418
rect 20397 251382 20565 251641
rect 20397 250605 20407 251382
rect 20555 250605 20565 251382
rect 20397 250346 20565 250605
rect 20397 249569 20407 250346
rect 20555 249569 20565 250346
rect 20397 249181 20565 249569
rect 20397 248404 20407 249181
rect 20555 248404 20565 249181
rect 20397 248145 20565 248404
rect 20397 247368 20407 248145
rect 20555 247368 20565 248145
rect 20397 247109 20565 247368
rect 20397 246332 20407 247109
rect 20555 246332 20565 247109
rect 20397 246073 20565 246332
rect 20397 245296 20407 246073
rect 20555 245296 20565 246073
rect 20397 245037 20565 245296
rect 20397 244260 20407 245037
rect 20555 244260 20565 245037
rect 20397 244248 20565 244260
rect 20607 254490 20775 254501
rect 20607 253713 20617 254490
rect 20765 253713 20775 254490
rect 20607 253454 20775 253713
rect 20607 252677 20617 253454
rect 20765 252677 20775 253454
rect 20607 252418 20775 252677
rect 20607 251641 20617 252418
rect 20765 251641 20775 252418
rect 20607 251382 20775 251641
rect 20607 250605 20617 251382
rect 20765 250605 20775 251382
rect 20607 250346 20775 250605
rect 20607 249569 20617 250346
rect 20765 249569 20775 250346
rect 20607 249181 20775 249569
rect 20607 248404 20617 249181
rect 20765 248404 20775 249181
rect 20607 248145 20775 248404
rect 20607 247368 20617 248145
rect 20765 247368 20775 248145
rect 20607 247109 20775 247368
rect 20607 246332 20617 247109
rect 20765 246332 20775 247109
rect 20607 246073 20775 246332
rect 20607 245296 20617 246073
rect 20765 245296 20775 246073
rect 20607 245037 20775 245296
rect 20607 244260 20617 245037
rect 20765 244260 20775 245037
rect 20607 244075 20775 244260
rect 20817 254490 20985 254737
rect 20817 253713 20827 254490
rect 20975 253713 20985 254490
rect 20817 253454 20985 253713
rect 20817 252677 20827 253454
rect 20975 252677 20985 253454
rect 20817 252418 20985 252677
rect 20817 251641 20827 252418
rect 20975 251641 20985 252418
rect 20817 251382 20985 251641
rect 20817 250605 20827 251382
rect 20975 250605 20985 251382
rect 20817 250346 20985 250605
rect 20817 249569 20827 250346
rect 20975 249569 20985 250346
rect 20817 249181 20985 249569
rect 20817 248404 20827 249181
rect 20975 248404 20985 249181
rect 20817 248145 20985 248404
rect 20817 247368 20827 248145
rect 20975 247368 20985 248145
rect 20817 247109 20985 247368
rect 20817 246332 20827 247109
rect 20975 246332 20985 247109
rect 20817 246073 20985 246332
rect 20817 245296 20827 246073
rect 20975 245296 20985 246073
rect 20817 245037 20985 245296
rect 20817 244260 20827 245037
rect 20975 244260 20985 245037
rect 20817 244248 20985 244260
rect 21027 254490 21195 254501
rect 21027 253713 21037 254490
rect 21185 253713 21195 254490
rect 21027 253454 21195 253713
rect 21027 252677 21037 253454
rect 21185 252677 21195 253454
rect 21027 252418 21195 252677
rect 21027 251641 21037 252418
rect 21185 251641 21195 252418
rect 21027 251382 21195 251641
rect 21027 250605 21037 251382
rect 21185 250605 21195 251382
rect 21027 250346 21195 250605
rect 21027 249569 21037 250346
rect 21185 249569 21195 250346
rect 21027 249181 21195 249569
rect 21027 248404 21037 249181
rect 21185 248404 21195 249181
rect 21027 248145 21195 248404
rect 21027 247368 21037 248145
rect 21185 247368 21195 248145
rect 21027 247109 21195 247368
rect 21027 246332 21037 247109
rect 21185 246332 21195 247109
rect 21027 246073 21195 246332
rect 21027 245296 21037 246073
rect 21185 245296 21195 246073
rect 21027 245037 21195 245296
rect 21027 244260 21037 245037
rect 21185 244260 21195 245037
rect 21027 244075 21195 244260
rect 21237 254490 21405 254737
rect 21237 253713 21247 254490
rect 21395 253713 21405 254490
rect 21237 253454 21405 253713
rect 21237 252677 21247 253454
rect 21395 252677 21405 253454
rect 21237 252418 21405 252677
rect 21237 251641 21247 252418
rect 21395 251641 21405 252418
rect 21237 251382 21405 251641
rect 21237 250605 21247 251382
rect 21395 250605 21405 251382
rect 21237 250346 21405 250605
rect 21237 249569 21247 250346
rect 21395 249569 21405 250346
rect 21237 249181 21405 249569
rect 21237 248404 21247 249181
rect 21395 248404 21405 249181
rect 21237 248145 21405 248404
rect 21237 247368 21247 248145
rect 21395 247368 21405 248145
rect 21237 247109 21405 247368
rect 21237 246332 21247 247109
rect 21395 246332 21405 247109
rect 21237 246073 21405 246332
rect 21237 245296 21247 246073
rect 21395 245296 21405 246073
rect 21237 245037 21405 245296
rect 21237 244260 21247 245037
rect 21395 244260 21405 245037
rect 21237 244248 21405 244260
rect 21447 254490 21615 254501
rect 21447 253713 21457 254490
rect 21605 253713 21615 254490
rect 21447 253454 21615 253713
rect 21447 252677 21457 253454
rect 21605 252677 21615 253454
rect 21447 252418 21615 252677
rect 21447 251641 21457 252418
rect 21605 251641 21615 252418
rect 21447 251382 21615 251641
rect 21447 250605 21457 251382
rect 21605 250605 21615 251382
rect 21447 250346 21615 250605
rect 21447 249569 21457 250346
rect 21605 249569 21615 250346
rect 21447 249181 21615 249569
rect 21447 248404 21457 249181
rect 21605 248404 21615 249181
rect 21447 248145 21615 248404
rect 21447 247368 21457 248145
rect 21605 247368 21615 248145
rect 21447 247109 21615 247368
rect 21447 246332 21457 247109
rect 21605 246332 21615 247109
rect 21447 246073 21615 246332
rect 21447 245296 21457 246073
rect 21605 245296 21615 246073
rect 21447 245037 21615 245296
rect 21447 244260 21457 245037
rect 21605 244260 21615 245037
rect 21447 244075 21615 244260
rect 21657 254490 21825 254737
rect 21657 253713 21667 254490
rect 21815 253713 21825 254490
rect 21657 253454 21825 253713
rect 21657 252677 21667 253454
rect 21815 252677 21825 253454
rect 21657 252418 21825 252677
rect 21657 251641 21667 252418
rect 21815 251641 21825 252418
rect 21657 251382 21825 251641
rect 21657 250605 21667 251382
rect 21815 250605 21825 251382
rect 21657 250346 21825 250605
rect 21657 249569 21667 250346
rect 21815 249569 21825 250346
rect 21657 249181 21825 249569
rect 21657 248404 21667 249181
rect 21815 248404 21825 249181
rect 21657 248145 21825 248404
rect 21657 247368 21667 248145
rect 21815 247368 21825 248145
rect 21657 247109 21825 247368
rect 21657 246332 21667 247109
rect 21815 246332 21825 247109
rect 21657 246073 21825 246332
rect 21657 245296 21667 246073
rect 21815 245296 21825 246073
rect 21657 245037 21825 245296
rect 21657 244260 21667 245037
rect 21815 244260 21825 245037
rect 21657 244248 21825 244260
rect 21867 254490 22035 254501
rect 21867 253713 21877 254490
rect 22025 253713 22035 254490
rect 21867 253454 22035 253713
rect 21867 252677 21877 253454
rect 22025 252677 22035 253454
rect 21867 252418 22035 252677
rect 21867 251641 21877 252418
rect 22025 251641 22035 252418
rect 21867 251382 22035 251641
rect 21867 250605 21877 251382
rect 22025 250605 22035 251382
rect 21867 250346 22035 250605
rect 21867 249569 21877 250346
rect 22025 249569 22035 250346
rect 21867 249181 22035 249569
rect 21867 248404 21877 249181
rect 22025 248404 22035 249181
rect 21867 248145 22035 248404
rect 21867 247368 21877 248145
rect 22025 247368 22035 248145
rect 21867 247109 22035 247368
rect 21867 246332 21877 247109
rect 22025 246332 22035 247109
rect 21867 246073 22035 246332
rect 21867 245296 21877 246073
rect 22025 245296 22035 246073
rect 21867 245037 22035 245296
rect 21867 244260 21877 245037
rect 22025 244260 22035 245037
rect 21867 244075 22035 244260
rect 22077 254490 22245 254737
rect 22077 253713 22087 254490
rect 22235 253713 22245 254490
rect 22077 253454 22245 253713
rect 22077 252677 22087 253454
rect 22235 252677 22245 253454
rect 22077 252418 22245 252677
rect 22077 251641 22087 252418
rect 22235 251641 22245 252418
rect 22077 251382 22245 251641
rect 22077 250605 22087 251382
rect 22235 250605 22245 251382
rect 22077 250346 22245 250605
rect 22077 249569 22087 250346
rect 22235 249569 22245 250346
rect 22077 249181 22245 249569
rect 22077 248404 22087 249181
rect 22235 248404 22245 249181
rect 22077 248145 22245 248404
rect 22077 247368 22087 248145
rect 22235 247368 22245 248145
rect 22077 247109 22245 247368
rect 22077 246332 22087 247109
rect 22235 246332 22245 247109
rect 22077 246073 22245 246332
rect 22077 245296 22087 246073
rect 22235 245296 22245 246073
rect 22077 245037 22245 245296
rect 22077 244260 22087 245037
rect 22235 244260 22245 245037
rect 22077 244248 22245 244260
rect 22287 254490 22455 254501
rect 22287 253713 22297 254490
rect 22445 253713 22455 254490
rect 22287 253454 22455 253713
rect 22287 252677 22297 253454
rect 22445 252677 22455 253454
rect 22287 252418 22455 252677
rect 22287 251641 22297 252418
rect 22445 251641 22455 252418
rect 22287 251382 22455 251641
rect 22287 250605 22297 251382
rect 22445 250605 22455 251382
rect 22287 250346 22455 250605
rect 22287 249569 22297 250346
rect 22445 249569 22455 250346
rect 22287 249181 22455 249569
rect 22287 248404 22297 249181
rect 22445 248404 22455 249181
rect 22287 248145 22455 248404
rect 22287 247368 22297 248145
rect 22445 247368 22455 248145
rect 22287 247109 22455 247368
rect 22287 246332 22297 247109
rect 22445 246332 22455 247109
rect 22287 246073 22455 246332
rect 22287 245296 22297 246073
rect 22445 245296 22455 246073
rect 22287 245037 22455 245296
rect 22287 244260 22297 245037
rect 22445 244260 22455 245037
rect 22287 244075 22455 244260
rect 22497 254490 22665 254737
rect 22497 253713 22507 254490
rect 22655 253713 22665 254490
rect 22497 253454 22665 253713
rect 22497 252677 22507 253454
rect 22655 252677 22665 253454
rect 22497 252418 22665 252677
rect 22497 251641 22507 252418
rect 22655 251641 22665 252418
rect 22497 251382 22665 251641
rect 22497 250605 22507 251382
rect 22655 250605 22665 251382
rect 22497 250346 22665 250605
rect 22497 249569 22507 250346
rect 22655 249569 22665 250346
rect 22497 249181 22665 249569
rect 22497 248404 22507 249181
rect 22655 248404 22665 249181
rect 22497 248145 22665 248404
rect 22497 247368 22507 248145
rect 22655 247368 22665 248145
rect 22497 247109 22665 247368
rect 22497 246332 22507 247109
rect 22655 246332 22665 247109
rect 22497 246073 22665 246332
rect 22497 245296 22507 246073
rect 22655 245296 22665 246073
rect 22497 245037 22665 245296
rect 22497 244260 22507 245037
rect 22655 244260 22665 245037
rect 22497 244248 22665 244260
rect 22707 254490 22875 254501
rect 22707 253713 22717 254490
rect 22865 253713 22875 254490
rect 22707 253454 22875 253713
rect 22707 252677 22717 253454
rect 22865 252677 22875 253454
rect 22707 252418 22875 252677
rect 22707 251641 22717 252418
rect 22865 251641 22875 252418
rect 22707 251382 22875 251641
rect 22707 250605 22717 251382
rect 22865 250605 22875 251382
rect 22707 250346 22875 250605
rect 22707 249569 22717 250346
rect 22865 249569 22875 250346
rect 22707 249181 22875 249569
rect 22707 248404 22717 249181
rect 22865 248404 22875 249181
rect 22707 248145 22875 248404
rect 22707 247368 22717 248145
rect 22865 247368 22875 248145
rect 22707 247109 22875 247368
rect 22707 246332 22717 247109
rect 22865 246332 22875 247109
rect 22707 246073 22875 246332
rect 22707 245296 22717 246073
rect 22865 245296 22875 246073
rect 22707 245037 22875 245296
rect 22707 244260 22717 245037
rect 22865 244260 22875 245037
rect 22707 244075 22875 244260
rect 22917 254490 23085 254737
rect 22917 253713 22927 254490
rect 23075 253713 23085 254490
rect 22917 253454 23085 253713
rect 22917 252677 22927 253454
rect 23075 252677 23085 253454
rect 22917 252418 23085 252677
rect 22917 251641 22927 252418
rect 23075 251641 23085 252418
rect 22917 251382 23085 251641
rect 22917 250605 22927 251382
rect 23075 250605 23085 251382
rect 22917 250346 23085 250605
rect 22917 249569 22927 250346
rect 23075 249569 23085 250346
rect 22917 249181 23085 249569
rect 22917 248404 22927 249181
rect 23075 248404 23085 249181
rect 22917 248145 23085 248404
rect 22917 247368 22927 248145
rect 23075 247368 23085 248145
rect 22917 247109 23085 247368
rect 22917 246332 22927 247109
rect 23075 246332 23085 247109
rect 22917 246073 23085 246332
rect 22917 245296 22927 246073
rect 23075 245296 23085 246073
rect 22917 245037 23085 245296
rect 22917 244260 22927 245037
rect 23075 244260 23085 245037
rect 22917 244248 23085 244260
rect 23127 254490 23295 254501
rect 23127 253713 23137 254490
rect 23285 253713 23295 254490
rect 23127 253454 23295 253713
rect 23127 252677 23137 253454
rect 23285 252677 23295 253454
rect 23127 252418 23295 252677
rect 23127 251641 23137 252418
rect 23285 251641 23295 252418
rect 23127 251382 23295 251641
rect 23127 250605 23137 251382
rect 23285 250605 23295 251382
rect 23127 250346 23295 250605
rect 23127 249569 23137 250346
rect 23285 249569 23295 250346
rect 23127 249181 23295 249569
rect 23127 248404 23137 249181
rect 23285 248404 23295 249181
rect 23127 248145 23295 248404
rect 23127 247368 23137 248145
rect 23285 247368 23295 248145
rect 23127 247109 23295 247368
rect 23127 246332 23137 247109
rect 23285 246332 23295 247109
rect 23127 246073 23295 246332
rect 23127 245296 23137 246073
rect 23285 245296 23295 246073
rect 23127 245037 23295 245296
rect 23127 244260 23137 245037
rect 23285 244260 23295 245037
rect 23127 244075 23295 244260
rect 23337 254490 23505 254737
rect 23337 253713 23347 254490
rect 23495 253713 23505 254490
rect 23337 253454 23505 253713
rect 23337 252677 23347 253454
rect 23495 252677 23505 253454
rect 23337 252418 23505 252677
rect 23337 251641 23347 252418
rect 23495 251641 23505 252418
rect 23337 251382 23505 251641
rect 23337 250605 23347 251382
rect 23495 250605 23505 251382
rect 23337 250346 23505 250605
rect 23337 249569 23347 250346
rect 23495 249569 23505 250346
rect 23337 249181 23505 249569
rect 23337 248404 23347 249181
rect 23495 248404 23505 249181
rect 23337 248145 23505 248404
rect 23337 247368 23347 248145
rect 23495 247368 23505 248145
rect 23337 247109 23505 247368
rect 23337 246332 23347 247109
rect 23495 246332 23505 247109
rect 23337 246073 23505 246332
rect 23337 245296 23347 246073
rect 23495 245296 23505 246073
rect 23337 245037 23505 245296
rect 23337 244260 23347 245037
rect 23495 244260 23505 245037
rect 23337 244248 23505 244260
rect 23547 254490 23715 254501
rect 23547 253713 23557 254490
rect 23705 253713 23715 254490
rect 23547 253454 23715 253713
rect 23547 252677 23557 253454
rect 23705 252677 23715 253454
rect 23547 252418 23715 252677
rect 23547 251641 23557 252418
rect 23705 251641 23715 252418
rect 23547 251382 23715 251641
rect 23547 250605 23557 251382
rect 23705 250605 23715 251382
rect 23547 250346 23715 250605
rect 23547 249569 23557 250346
rect 23705 249569 23715 250346
rect 23547 249181 23715 249569
rect 23547 248404 23557 249181
rect 23705 248404 23715 249181
rect 23547 248145 23715 248404
rect 23547 247368 23557 248145
rect 23705 247368 23715 248145
rect 23547 247109 23715 247368
rect 23547 246332 23557 247109
rect 23705 246332 23715 247109
rect 23547 246073 23715 246332
rect 23547 245296 23557 246073
rect 23705 245296 23715 246073
rect 23547 245037 23715 245296
rect 23547 244260 23557 245037
rect 23705 244260 23715 245037
rect 23547 244075 23715 244260
rect 23757 254490 23925 254737
rect 23757 253713 23767 254490
rect 23915 253713 23925 254490
rect 23757 253454 23925 253713
rect 23757 252677 23767 253454
rect 23915 252677 23925 253454
rect 23757 252418 23925 252677
rect 23757 251641 23767 252418
rect 23915 251641 23925 252418
rect 23757 251382 23925 251641
rect 23757 250605 23767 251382
rect 23915 250605 23925 251382
rect 23757 250346 23925 250605
rect 23757 249569 23767 250346
rect 23915 249569 23925 250346
rect 23757 249181 23925 249569
rect 23757 248404 23767 249181
rect 23915 248404 23925 249181
rect 23757 248145 23925 248404
rect 23757 247368 23767 248145
rect 23915 247368 23925 248145
rect 23757 247109 23925 247368
rect 23757 246332 23767 247109
rect 23915 246332 23925 247109
rect 23757 246073 23925 246332
rect 23757 245296 23767 246073
rect 23915 245296 23925 246073
rect 23757 245037 23925 245296
rect 23757 244260 23767 245037
rect 23915 244260 23925 245037
rect 23757 244248 23925 244260
rect 23967 254490 24135 254501
rect 23967 253713 23977 254490
rect 24125 253713 24135 254490
rect 23967 253454 24135 253713
rect 23967 252677 23977 253454
rect 24125 252677 24135 253454
rect 23967 252418 24135 252677
rect 23967 251641 23977 252418
rect 24125 251641 24135 252418
rect 23967 251382 24135 251641
rect 23967 250605 23977 251382
rect 24125 250605 24135 251382
rect 23967 250346 24135 250605
rect 23967 249569 23977 250346
rect 24125 249569 24135 250346
rect 23967 249181 24135 249569
rect 23967 248404 23977 249181
rect 24125 248404 24135 249181
rect 23967 248145 24135 248404
rect 23967 247368 23977 248145
rect 24125 247368 24135 248145
rect 23967 247109 24135 247368
rect 23967 246332 23977 247109
rect 24125 246332 24135 247109
rect 23967 246073 24135 246332
rect 23967 245296 23977 246073
rect 24125 245296 24135 246073
rect 23967 245037 24135 245296
rect 23967 244260 23977 245037
rect 24125 244260 24135 245037
rect 23967 244075 24135 244260
rect 24177 254490 24345 254737
rect 24177 253713 24187 254490
rect 24335 253713 24345 254490
rect 24177 253454 24345 253713
rect 24177 252677 24187 253454
rect 24335 252677 24345 253454
rect 24177 252418 24345 252677
rect 24177 251641 24187 252418
rect 24335 251641 24345 252418
rect 24177 251382 24345 251641
rect 24177 250605 24187 251382
rect 24335 250605 24345 251382
rect 24177 250346 24345 250605
rect 24177 249569 24187 250346
rect 24335 249569 24345 250346
rect 24177 249181 24345 249569
rect 24177 248404 24187 249181
rect 24335 248404 24345 249181
rect 24177 248145 24345 248404
rect 24177 247368 24187 248145
rect 24335 247368 24345 248145
rect 24177 247109 24345 247368
rect 24177 246332 24187 247109
rect 24335 246332 24345 247109
rect 24177 246073 24345 246332
rect 24177 245296 24187 246073
rect 24335 245296 24345 246073
rect 24177 245037 24345 245296
rect 24177 244260 24187 245037
rect 24335 244260 24345 245037
rect 24177 244248 24345 244260
rect 24387 254490 24555 254501
rect 24387 253713 24397 254490
rect 24545 253713 24555 254490
rect 24387 253454 24555 253713
rect 24387 252677 24397 253454
rect 24545 252677 24555 253454
rect 24387 252418 24555 252677
rect 24387 251641 24397 252418
rect 24545 251641 24555 252418
rect 24387 251382 24555 251641
rect 24387 250605 24397 251382
rect 24545 250605 24555 251382
rect 24387 250346 24555 250605
rect 24387 249569 24397 250346
rect 24545 249569 24555 250346
rect 24387 249181 24555 249569
rect 24387 248404 24397 249181
rect 24545 248404 24555 249181
rect 24387 248145 24555 248404
rect 24387 247368 24397 248145
rect 24545 247368 24555 248145
rect 24387 247109 24555 247368
rect 24387 246332 24397 247109
rect 24545 246332 24555 247109
rect 24387 246073 24555 246332
rect 24387 245296 24397 246073
rect 24545 245296 24555 246073
rect 24387 245037 24555 245296
rect 24387 244260 24397 245037
rect 24545 244260 24555 245037
rect 24387 244075 24555 244260
rect 24597 254490 24765 254737
rect 24597 253713 24607 254490
rect 24755 253713 24765 254490
rect 24597 253454 24765 253713
rect 24597 252677 24607 253454
rect 24755 252677 24765 253454
rect 24597 252418 24765 252677
rect 24597 251641 24607 252418
rect 24755 251641 24765 252418
rect 24597 251382 24765 251641
rect 24597 250605 24607 251382
rect 24755 250605 24765 251382
rect 24597 250346 24765 250605
rect 24597 249569 24607 250346
rect 24755 249569 24765 250346
rect 24597 249181 24765 249569
rect 24597 248404 24607 249181
rect 24755 248404 24765 249181
rect 24597 248145 24765 248404
rect 24597 247368 24607 248145
rect 24755 247368 24765 248145
rect 24597 247109 24765 247368
rect 24597 246332 24607 247109
rect 24755 246332 24765 247109
rect 24597 246073 24765 246332
rect 24597 245296 24607 246073
rect 24755 245296 24765 246073
rect 24597 245037 24765 245296
rect 24597 244260 24607 245037
rect 24755 244260 24765 245037
rect 24597 244248 24765 244260
rect 24807 254490 24975 254501
rect 24807 253713 24817 254490
rect 24965 253713 24975 254490
rect 24807 253454 24975 253713
rect 24807 252677 24817 253454
rect 24965 252677 24975 253454
rect 24807 252418 24975 252677
rect 24807 251641 24817 252418
rect 24965 251641 24975 252418
rect 24807 251382 24975 251641
rect 24807 250605 24817 251382
rect 24965 250605 24975 251382
rect 24807 250346 24975 250605
rect 24807 249569 24817 250346
rect 24965 249569 24975 250346
rect 24807 249181 24975 249569
rect 24807 248404 24817 249181
rect 24965 248404 24975 249181
rect 24807 248145 24975 248404
rect 24807 247368 24817 248145
rect 24965 247368 24975 248145
rect 24807 247109 24975 247368
rect 24807 246332 24817 247109
rect 24965 246332 24975 247109
rect 24807 246073 24975 246332
rect 24807 245296 24817 246073
rect 24965 245296 24975 246073
rect 24807 245037 24975 245296
rect 24807 244260 24817 245037
rect 24965 244260 24975 245037
rect 24807 244075 24975 244260
rect 25017 254490 25185 254737
rect 25017 253713 25027 254490
rect 25175 253713 25185 254490
rect 25017 253454 25185 253713
rect 25017 252677 25027 253454
rect 25175 252677 25185 253454
rect 25017 252418 25185 252677
rect 25017 251641 25027 252418
rect 25175 251641 25185 252418
rect 25017 251382 25185 251641
rect 25017 250605 25027 251382
rect 25175 250605 25185 251382
rect 25017 250346 25185 250605
rect 25017 249569 25027 250346
rect 25175 249569 25185 250346
rect 25017 249181 25185 249569
rect 25017 248404 25027 249181
rect 25175 248404 25185 249181
rect 25017 248145 25185 248404
rect 25017 247368 25027 248145
rect 25175 247368 25185 248145
rect 25017 247109 25185 247368
rect 25017 246332 25027 247109
rect 25175 246332 25185 247109
rect 25017 246073 25185 246332
rect 25017 245296 25027 246073
rect 25175 245296 25185 246073
rect 25017 245037 25185 245296
rect 25017 244260 25027 245037
rect 25175 244260 25185 245037
rect 25017 244248 25185 244260
rect 25227 254490 25395 254501
rect 25227 253713 25237 254490
rect 25385 253713 25395 254490
rect 25227 253454 25395 253713
rect 25227 252677 25237 253454
rect 25385 252677 25395 253454
rect 25227 252418 25395 252677
rect 25227 251641 25237 252418
rect 25385 251641 25395 252418
rect 25227 251382 25395 251641
rect 25227 250605 25237 251382
rect 25385 250605 25395 251382
rect 25227 250346 25395 250605
rect 25227 249569 25237 250346
rect 25385 249569 25395 250346
rect 25227 249181 25395 249569
rect 25227 248404 25237 249181
rect 25385 248404 25395 249181
rect 25227 248145 25395 248404
rect 25227 247368 25237 248145
rect 25385 247368 25395 248145
rect 25227 247109 25395 247368
rect 25227 246332 25237 247109
rect 25385 246332 25395 247109
rect 25227 246073 25395 246332
rect 25227 245296 25237 246073
rect 25385 245296 25395 246073
rect 25227 245037 25395 245296
rect 25227 244260 25237 245037
rect 25385 244260 25395 245037
rect 25227 244075 25395 244260
rect 25437 254490 25605 254737
rect 25437 253713 25447 254490
rect 25595 253713 25605 254490
rect 25437 253454 25605 253713
rect 25437 252677 25447 253454
rect 25595 252677 25605 253454
rect 25437 252418 25605 252677
rect 25437 251641 25447 252418
rect 25595 251641 25605 252418
rect 25437 251382 25605 251641
rect 25437 250605 25447 251382
rect 25595 250605 25605 251382
rect 25437 250346 25605 250605
rect 25437 249569 25447 250346
rect 25595 249569 25605 250346
rect 25437 249181 25605 249569
rect 25437 248404 25447 249181
rect 25595 248404 25605 249181
rect 25437 248145 25605 248404
rect 25437 247368 25447 248145
rect 25595 247368 25605 248145
rect 25437 247109 25605 247368
rect 25437 246332 25447 247109
rect 25595 246332 25605 247109
rect 25437 246073 25605 246332
rect 25437 245296 25447 246073
rect 25595 245296 25605 246073
rect 25437 245037 25605 245296
rect 25437 244260 25447 245037
rect 25595 244260 25605 245037
rect 25437 244248 25605 244260
rect 25647 254490 25815 254501
rect 25647 253713 25657 254490
rect 25805 253713 25815 254490
rect 25647 253454 25815 253713
rect 25647 252677 25657 253454
rect 25805 252677 25815 253454
rect 25647 252418 25815 252677
rect 25647 251641 25657 252418
rect 25805 251641 25815 252418
rect 25647 251382 25815 251641
rect 25647 250605 25657 251382
rect 25805 250605 25815 251382
rect 25647 250346 25815 250605
rect 25647 249569 25657 250346
rect 25805 249569 25815 250346
rect 25647 249181 25815 249569
rect 25647 248404 25657 249181
rect 25805 248404 25815 249181
rect 25647 248145 25815 248404
rect 25647 247368 25657 248145
rect 25805 247368 25815 248145
rect 25647 247109 25815 247368
rect 25647 246332 25657 247109
rect 25805 246332 25815 247109
rect 25647 246073 25815 246332
rect 25647 245296 25657 246073
rect 25805 245296 25815 246073
rect 25647 245037 25815 245296
rect 25647 244260 25657 245037
rect 25805 244260 25815 245037
rect 25647 244075 25815 244260
rect 25857 254490 26025 254737
rect 25857 253713 25867 254490
rect 26015 253713 26025 254490
rect 25857 253454 26025 253713
rect 25857 252677 25867 253454
rect 26015 252677 26025 253454
rect 25857 252418 26025 252677
rect 25857 251641 25867 252418
rect 26015 251641 26025 252418
rect 25857 251382 26025 251641
rect 25857 250605 25867 251382
rect 26015 250605 26025 251382
rect 25857 250346 26025 250605
rect 25857 249569 25867 250346
rect 26015 249569 26025 250346
rect 25857 249181 26025 249569
rect 25857 248404 25867 249181
rect 26015 248404 26025 249181
rect 25857 248145 26025 248404
rect 25857 247368 25867 248145
rect 26015 247368 26025 248145
rect 25857 247109 26025 247368
rect 25857 246332 25867 247109
rect 26015 246332 26025 247109
rect 25857 246073 26025 246332
rect 25857 245296 25867 246073
rect 26015 245296 26025 246073
rect 25857 245037 26025 245296
rect 25857 244260 25867 245037
rect 26015 244260 26025 245037
rect 25857 244248 26025 244260
rect 26067 254490 26235 254501
rect 26067 253713 26077 254490
rect 26225 253713 26235 254490
rect 26067 253454 26235 253713
rect 26067 252677 26077 253454
rect 26225 252677 26235 253454
rect 26067 252418 26235 252677
rect 26067 251641 26077 252418
rect 26225 251641 26235 252418
rect 26067 251382 26235 251641
rect 26067 250605 26077 251382
rect 26225 250605 26235 251382
rect 26067 250346 26235 250605
rect 26067 249569 26077 250346
rect 26225 249569 26235 250346
rect 26067 249181 26235 249569
rect 26067 248404 26077 249181
rect 26225 248404 26235 249181
rect 26067 248145 26235 248404
rect 26067 247368 26077 248145
rect 26225 247368 26235 248145
rect 26067 247109 26235 247368
rect 26067 246332 26077 247109
rect 26225 246332 26235 247109
rect 26067 246073 26235 246332
rect 26067 245296 26077 246073
rect 26225 245296 26235 246073
rect 26067 245037 26235 245296
rect 26067 244260 26077 245037
rect 26225 244260 26235 245037
rect 26067 244075 26235 244260
rect 26277 254490 26445 254737
rect 26277 253713 26287 254490
rect 26435 253713 26445 254490
rect 26277 253454 26445 253713
rect 26277 252677 26287 253454
rect 26435 252677 26445 253454
rect 26277 252418 26445 252677
rect 26277 251641 26287 252418
rect 26435 251641 26445 252418
rect 26277 251382 26445 251641
rect 26277 250605 26287 251382
rect 26435 250605 26445 251382
rect 26277 250346 26445 250605
rect 26277 249569 26287 250346
rect 26435 249569 26445 250346
rect 26277 249181 26445 249569
rect 26277 248404 26287 249181
rect 26435 248404 26445 249181
rect 26277 248145 26445 248404
rect 26277 247368 26287 248145
rect 26435 247368 26445 248145
rect 26277 247109 26445 247368
rect 26277 246332 26287 247109
rect 26435 246332 26445 247109
rect 26277 246073 26445 246332
rect 26277 245296 26287 246073
rect 26435 245296 26445 246073
rect 26277 245037 26445 245296
rect 26277 244260 26287 245037
rect 26435 244260 26445 245037
rect 26277 244248 26445 244260
rect 26487 254490 26655 254501
rect 26487 253713 26497 254490
rect 26645 253713 26655 254490
rect 26487 253454 26655 253713
rect 26487 252677 26497 253454
rect 26645 252677 26655 253454
rect 26487 252418 26655 252677
rect 26487 251641 26497 252418
rect 26645 251641 26655 252418
rect 26487 251382 26655 251641
rect 26487 250605 26497 251382
rect 26645 250605 26655 251382
rect 26487 250346 26655 250605
rect 26487 249569 26497 250346
rect 26645 249569 26655 250346
rect 26487 249181 26655 249569
rect 26487 248404 26497 249181
rect 26645 248404 26655 249181
rect 26487 248145 26655 248404
rect 26487 247368 26497 248145
rect 26645 247368 26655 248145
rect 26487 247109 26655 247368
rect 26487 246332 26497 247109
rect 26645 246332 26655 247109
rect 26487 246073 26655 246332
rect 26487 245296 26497 246073
rect 26645 245296 26655 246073
rect 26487 245037 26655 245296
rect 26487 244260 26497 245037
rect 26645 244260 26655 245037
rect 26487 244075 26655 244260
rect 26697 254490 26865 254737
rect 26697 253713 26707 254490
rect 26855 253713 26865 254490
rect 26697 253454 26865 253713
rect 26697 252677 26707 253454
rect 26855 252677 26865 253454
rect 26697 252418 26865 252677
rect 26697 251641 26707 252418
rect 26855 251641 26865 252418
rect 26697 251382 26865 251641
rect 26697 250605 26707 251382
rect 26855 250605 26865 251382
rect 26697 250346 26865 250605
rect 26697 249569 26707 250346
rect 26855 249569 26865 250346
rect 26697 249181 26865 249569
rect 26697 248404 26707 249181
rect 26855 248404 26865 249181
rect 26697 248145 26865 248404
rect 26697 247368 26707 248145
rect 26855 247368 26865 248145
rect 26697 247109 26865 247368
rect 26697 246332 26707 247109
rect 26855 246332 26865 247109
rect 26697 246073 26865 246332
rect 26697 245296 26707 246073
rect 26855 245296 26865 246073
rect 26697 245037 26865 245296
rect 26697 244260 26707 245037
rect 26855 244260 26865 245037
rect 26697 244248 26865 244260
rect 26907 254490 27075 254501
rect 26907 253713 26917 254490
rect 27065 253713 27075 254490
rect 26907 253454 27075 253713
rect 26907 252677 26917 253454
rect 27065 252677 27075 253454
rect 26907 252418 27075 252677
rect 26907 251641 26917 252418
rect 27065 251641 27075 252418
rect 26907 251382 27075 251641
rect 26907 250605 26917 251382
rect 27065 250605 27075 251382
rect 26907 250346 27075 250605
rect 26907 249569 26917 250346
rect 27065 249569 27075 250346
rect 26907 249181 27075 249569
rect 26907 248404 26917 249181
rect 27065 248404 27075 249181
rect 26907 248145 27075 248404
rect 26907 247368 26917 248145
rect 27065 247368 27075 248145
rect 26907 247109 27075 247368
rect 26907 246332 26917 247109
rect 27065 246332 27075 247109
rect 26907 246073 27075 246332
rect 26907 245296 26917 246073
rect 27065 245296 27075 246073
rect 26907 245037 27075 245296
rect 26907 244260 26917 245037
rect 27065 244260 27075 245037
rect 26907 244075 27075 244260
rect 27117 254490 27285 254737
rect 27117 253713 27127 254490
rect 27275 253713 27285 254490
rect 27117 253454 27285 253713
rect 27117 252677 27127 253454
rect 27275 252677 27285 253454
rect 27117 252418 27285 252677
rect 27117 251641 27127 252418
rect 27275 251641 27285 252418
rect 27117 251382 27285 251641
rect 27117 250605 27127 251382
rect 27275 250605 27285 251382
rect 27117 250346 27285 250605
rect 27117 249569 27127 250346
rect 27275 249569 27285 250346
rect 27117 249181 27285 249569
rect 27117 248404 27127 249181
rect 27275 248404 27285 249181
rect 27117 248145 27285 248404
rect 27117 247368 27127 248145
rect 27275 247368 27285 248145
rect 27117 247109 27285 247368
rect 27117 246332 27127 247109
rect 27275 246332 27285 247109
rect 27117 246073 27285 246332
rect 27117 245296 27127 246073
rect 27275 245296 27285 246073
rect 27117 245037 27285 245296
rect 27117 244260 27127 245037
rect 27275 244260 27285 245037
rect 27117 244248 27285 244260
rect -4163 244065 27485 244075
rect -4180 244041 -4163 244051
rect 27485 244041 27614 244051
rect -3980 243950 -3771 243960
rect -4180 243831 -3980 243841
rect -3571 243950 -3351 243960
rect -3771 243831 -3571 243841
rect -3151 243950 -2931 243960
rect -3351 243831 -3151 243841
rect -2731 243950 -2511 243960
rect -2931 243831 -2731 243841
rect -2311 243950 -2091 243960
rect -2511 243831 -2311 243841
rect -1891 243950 -1671 243960
rect -2091 243831 -1891 243841
rect -1471 243950 -1251 243960
rect -1671 243831 -1471 243841
rect -1051 243950 -831 243960
rect -1251 243831 -1051 243841
rect -631 243950 -411 243960
rect -831 243831 -631 243841
rect -211 243950 9 243960
rect -411 243831 -211 243841
rect 209 243950 429 243960
rect 9 243831 209 243841
rect 629 243950 849 243960
rect 429 243831 629 243841
rect 1049 243950 1269 243960
rect 849 243831 1049 243841
rect 1469 243950 1689 243960
rect 1269 243831 1469 243841
rect 1889 243950 2109 243960
rect 1689 243831 1889 243841
rect 2309 243950 2529 243960
rect 2109 243831 2309 243841
rect 2729 243950 2949 243960
rect 2529 243831 2729 243841
rect 3149 243950 3369 243960
rect 2949 243831 3149 243841
rect 3569 243950 3789 243960
rect 3369 243831 3569 243841
rect 3989 243950 4209 243960
rect 3789 243831 3989 243841
rect 4409 243950 4629 243960
rect 4209 243831 4409 243841
rect 4829 243950 5049 243960
rect 4629 243831 4829 243841
rect 5249 243950 5469 243960
rect 5049 243831 5249 243841
rect 5669 243950 5889 243960
rect 5469 243831 5669 243841
rect 6089 243950 6309 243960
rect 5889 243831 6089 243841
rect 6509 243950 6729 243960
rect 6309 243831 6509 243841
rect 6929 243950 7149 243960
rect 6729 243831 6929 243841
rect 7349 243950 7569 243960
rect 7149 243831 7349 243841
rect 7769 243950 7989 243960
rect 7569 243831 7769 243841
rect 8189 243950 8409 243960
rect 7989 243831 8189 243841
rect 8609 243950 8829 243960
rect 8409 243831 8609 243841
rect 9029 243950 9249 243960
rect 8829 243831 9029 243841
rect 9449 243950 9669 243960
rect 9249 243831 9449 243841
rect 9869 243950 10089 243960
rect 9669 243831 9869 243841
rect 10289 243950 10509 243960
rect 10089 243831 10289 243841
rect 10709 243950 10929 243960
rect 10509 243831 10709 243841
rect 11129 243950 11349 243960
rect 10929 243831 11129 243841
rect 11549 243950 11769 243960
rect 11349 243831 11549 243841
rect 11969 243950 12189 243960
rect 11769 243831 11969 243841
rect 12389 243950 12609 243960
rect 12189 243831 12389 243841
rect 12809 243950 13029 243960
rect 12609 243831 12809 243841
rect 13229 243950 13449 243960
rect 13029 243831 13229 243841
rect 13649 243950 13869 243960
rect 13449 243831 13649 243841
rect 14069 243950 14289 243960
rect 13869 243831 14069 243841
rect 14489 243950 14709 243960
rect 14289 243831 14489 243841
rect 14909 243950 15129 243960
rect 14709 243831 14909 243841
rect 15329 243950 15549 243960
rect 15129 243831 15329 243841
rect 15749 243950 15969 243960
rect 15549 243831 15749 243841
rect 16169 243950 16389 243960
rect 15969 243831 16169 243841
rect 16589 243950 16809 243960
rect 16389 243831 16589 243841
rect 17009 243950 17229 243960
rect 16809 243831 17009 243841
rect 17429 243950 17649 243960
rect 17229 243831 17429 243841
rect 17849 243950 18069 243960
rect 17649 243831 17849 243841
rect 18269 243950 18489 243960
rect 18069 243831 18269 243841
rect 18689 243950 18909 243960
rect 18489 243831 18689 243841
rect 19109 243950 19329 243960
rect 18909 243831 19109 243841
rect 19529 243950 19749 243960
rect 19329 243831 19529 243841
rect 19949 243950 20169 243960
rect 19749 243831 19949 243841
rect 20369 243950 20589 243960
rect 20169 243831 20369 243841
rect 20789 243950 21009 243960
rect 20589 243831 20789 243841
rect 21209 243950 21429 243960
rect 21009 243831 21209 243841
rect 21629 243950 21849 243960
rect 21429 243831 21629 243841
rect 22049 243950 22269 243960
rect 21849 243831 22049 243841
rect 22469 243950 22689 243960
rect 22269 243831 22469 243841
rect 22889 243950 23109 243960
rect 22689 243831 22889 243841
rect 23309 243950 23529 243960
rect 23109 243831 23309 243841
rect 23729 243950 23949 243960
rect 23529 243831 23729 243841
rect 24149 243950 24369 243960
rect 23949 243831 24149 243841
rect 24569 243950 24789 243960
rect 24369 243831 24569 243841
rect 24989 243950 25209 243960
rect 24789 243831 24989 243841
rect 25409 243950 25629 243960
rect 25209 243831 25409 243841
rect 25829 243950 26049 243960
rect 25629 243831 25829 243841
rect 26249 243950 26469 243960
rect 26049 243831 26249 243841
rect 26669 243950 26889 243960
rect 26469 243831 26669 243841
rect 27089 243950 27414 243960
rect 26889 243831 27089 243841
rect 27414 243831 27614 243841
<< via2 >>
rect -4179 264317 -3979 264430
rect -3770 264317 -3570 264430
rect -3350 264317 -3150 264430
rect -2930 264317 -2730 264430
rect -2510 264317 -2310 264430
rect -2090 264317 -1890 264430
rect -1670 264317 -1470 264430
rect -1250 264317 -1050 264430
rect -830 264317 -630 264430
rect -410 264317 -210 264430
rect 10 264317 210 264430
rect 430 264317 630 264430
rect 850 264317 1050 264430
rect 1270 264317 1470 264430
rect 1690 264317 1890 264430
rect 2110 264317 2310 264430
rect 2530 264317 2730 264430
rect 2950 264317 3150 264430
rect 3370 264317 3570 264430
rect 3790 264317 3990 264430
rect 4210 264317 4410 264430
rect 4630 264317 4830 264430
rect 5050 264317 5250 264430
rect 5470 264317 5670 264430
rect 5890 264317 6090 264430
rect 6310 264317 6510 264430
rect 6730 264317 6930 264430
rect 7150 264317 7350 264430
rect 7570 264317 7770 264430
rect 7990 264317 8190 264430
rect 8410 264317 8610 264430
rect 8830 264317 9030 264430
rect 9250 264317 9450 264430
rect 9670 264317 9870 264430
rect 10090 264317 10290 264430
rect 10510 264317 10710 264430
rect 10930 264317 11130 264430
rect 11350 264317 11550 264430
rect 11770 264317 11970 264430
rect 12190 264317 12390 264430
rect 12610 264317 12810 264430
rect 13030 264317 13230 264430
rect 13450 264317 13650 264430
rect 13870 264317 14070 264430
rect 14290 264317 14490 264430
rect 14710 264317 14910 264430
rect 15130 264317 15330 264430
rect 15550 264317 15750 264430
rect 15970 264317 16170 264430
rect 16390 264317 16590 264430
rect 16810 264317 17010 264430
rect 17230 264317 17430 264430
rect 17650 264317 17850 264430
rect 18070 264317 18270 264430
rect 18490 264317 18690 264430
rect 18910 264317 19110 264430
rect 19330 264317 19530 264430
rect 19750 264317 19950 264430
rect 20170 264317 20370 264430
rect 20590 264317 20790 264430
rect 21010 264317 21210 264430
rect 21430 264317 21630 264430
rect 21850 264317 22050 264430
rect 22270 264317 22470 264430
rect 22690 264317 22890 264430
rect 23110 264317 23310 264430
rect 23530 264317 23730 264430
rect 23950 264317 24150 264430
rect 24370 264317 24570 264430
rect 24790 264317 24990 264430
rect 25210 264317 25410 264430
rect 25630 264317 25830 264430
rect 26050 264317 26250 264430
rect 26470 264317 26670 264430
rect 26890 264317 27090 264430
rect -4179 264230 -4163 264317
rect -4163 264230 -3979 264317
rect -3770 264230 -3570 264317
rect -3350 264230 -3150 264317
rect -2930 264230 -2730 264317
rect -2510 264230 -2310 264317
rect -2090 264230 -1890 264317
rect -1670 264230 -1470 264317
rect -1250 264230 -1050 264317
rect -830 264230 -630 264317
rect -410 264230 -210 264317
rect 10 264230 210 264317
rect 430 264230 630 264317
rect 850 264230 1050 264317
rect 1270 264230 1470 264317
rect 1690 264230 1890 264317
rect 2110 264230 2310 264317
rect 2530 264230 2730 264317
rect 2950 264230 3150 264317
rect 3370 264230 3570 264317
rect 3790 264230 3990 264317
rect 4210 264230 4410 264317
rect 4630 264230 4830 264317
rect 5050 264230 5250 264317
rect 5470 264230 5670 264317
rect 5890 264230 6090 264317
rect 6310 264230 6510 264317
rect 6730 264230 6930 264317
rect 7150 264230 7350 264317
rect 7570 264230 7770 264317
rect 7990 264230 8190 264317
rect 8410 264230 8610 264317
rect 8830 264230 9030 264317
rect 9250 264230 9450 264317
rect 9670 264230 9870 264317
rect 10090 264230 10290 264317
rect 10510 264230 10710 264317
rect 10930 264230 11130 264317
rect 11350 264230 11550 264317
rect 11770 264230 11970 264317
rect 12190 264230 12390 264317
rect 12610 264230 12810 264317
rect 13030 264230 13230 264317
rect 13450 264230 13650 264317
rect 13870 264230 14070 264317
rect 14290 264230 14490 264317
rect 14710 264230 14910 264317
rect 15130 264230 15330 264317
rect 15550 264230 15750 264317
rect 15970 264230 16170 264317
rect 16390 264230 16590 264317
rect 16810 264230 17010 264317
rect 17230 264230 17430 264317
rect 17650 264230 17850 264317
rect 18070 264230 18270 264317
rect 18490 264230 18690 264317
rect 18910 264230 19110 264317
rect 19330 264230 19530 264317
rect 19750 264230 19950 264317
rect 20170 264230 20370 264317
rect 20590 264230 20790 264317
rect 21010 264230 21210 264317
rect 21430 264230 21630 264317
rect 21850 264230 22050 264317
rect 22270 264230 22470 264317
rect 22690 264230 22890 264317
rect 23110 264230 23310 264317
rect 23530 264230 23730 264317
rect 23950 264230 24150 264317
rect 24370 264230 24570 264317
rect 24790 264230 24990 264317
rect 25210 264230 25410 264317
rect 25630 264230 25830 264317
rect 26050 264230 26250 264317
rect 26470 264230 26670 264317
rect 26890 264230 27090 264317
rect 27310 264230 27510 264430
rect -3980 261752 -3780 261952
rect -3560 261752 -3360 261952
rect -3140 261752 -2940 261952
rect -2720 261752 -2520 261952
rect -2300 261752 -2100 261952
rect -1880 261752 -1680 261952
rect -1460 261752 -1260 261952
rect -1040 261752 -840 261952
rect -620 261752 -420 261952
rect -200 261752 0 261952
rect 220 261752 420 261952
rect 640 261752 840 261952
rect 1060 261752 1260 261952
rect 1480 261752 1680 261952
rect 1900 261752 2100 261952
rect 2320 261752 2520 261952
rect 2740 261752 2940 261952
rect 3160 261752 3360 261952
rect 3580 261752 3780 261952
rect 4000 261752 4200 261952
rect 4420 261752 4620 261952
rect 4840 261752 5040 261952
rect 5260 261752 5460 261952
rect 5680 261752 5880 261952
rect 6100 261752 6300 261952
rect 6520 261752 6720 261952
rect 6940 261752 7140 261952
rect 7360 261752 7560 261952
rect 7780 261752 7980 261952
rect 8200 261752 8400 261952
rect 8620 261752 8820 261952
rect 9040 261752 9240 261952
rect 9460 261752 9660 261952
rect 9880 261752 10080 261952
rect 10300 261752 10500 261952
rect 10720 261752 10920 261952
rect 11140 261752 11340 261952
rect 11560 261752 11760 261952
rect 11980 261752 12180 261952
rect 12400 261752 12600 261952
rect 12820 261752 13020 261952
rect 13240 261752 13440 261952
rect 13660 261752 13860 261952
rect 14080 261752 14280 261952
rect 14500 261752 14700 261952
rect 14920 261752 15120 261952
rect 15340 261752 15540 261952
rect 15760 261752 15960 261952
rect 16180 261752 16380 261952
rect 16600 261752 16800 261952
rect 17020 261752 17220 261952
rect 17440 261752 17640 261952
rect 17860 261752 18060 261952
rect 18280 261752 18480 261952
rect 18700 261752 18900 261952
rect 19120 261752 19320 261952
rect 19540 261752 19740 261952
rect 19960 261752 20160 261952
rect 20380 261752 20580 261952
rect 20800 261752 21000 261952
rect 21220 261752 21420 261952
rect 21640 261752 21840 261952
rect 22060 261752 22260 261952
rect 22480 261752 22680 261952
rect 22900 261752 23100 261952
rect 23320 261752 23520 261952
rect 23740 261752 23940 261952
rect 24160 261752 24360 261952
rect 24580 261752 24780 261952
rect 25000 261752 25200 261952
rect 25420 261752 25620 261952
rect 25840 261752 26040 261952
rect 26260 261752 26460 261952
rect 26680 261752 26880 261952
rect 27100 261752 27300 261952
rect -3979 254747 -3779 254947
rect -3559 254747 -3359 254947
rect -3139 254747 -2939 254947
rect -2719 254747 -2519 254947
rect -2299 254747 -2099 254947
rect -1879 254747 -1679 254947
rect -1459 254747 -1259 254947
rect -1039 254747 -839 254947
rect -619 254747 -419 254947
rect -199 254747 1 254947
rect 221 254747 421 254947
rect 641 254747 841 254947
rect 1061 254747 1261 254947
rect 1481 254747 1681 254947
rect 1901 254747 2101 254947
rect 2321 254747 2521 254947
rect 2741 254747 2941 254947
rect 3161 254747 3361 254947
rect 3581 254747 3781 254947
rect 4001 254747 4201 254947
rect 4421 254747 4621 254947
rect 4841 254747 5041 254947
rect 5261 254747 5461 254947
rect 5681 254747 5881 254947
rect 6101 254747 6301 254947
rect 6521 254747 6721 254947
rect 6941 254747 7141 254947
rect 7361 254747 7561 254947
rect 7781 254747 7981 254947
rect 8201 254747 8401 254947
rect 8621 254747 8821 254947
rect 9041 254747 9241 254947
rect 9461 254747 9661 254947
rect 9881 254747 10081 254947
rect 10301 254747 10501 254947
rect 10721 254747 10921 254947
rect 11141 254747 11341 254947
rect 11561 254747 11761 254947
rect 11981 254747 12181 254947
rect 12401 254747 12601 254947
rect 12821 254747 13021 254947
rect 13241 254747 13441 254947
rect 13661 254747 13861 254947
rect 14081 254747 14281 254947
rect 14501 254747 14701 254947
rect 14921 254747 15121 254947
rect 15341 254747 15541 254947
rect 15761 254747 15961 254947
rect 16181 254747 16381 254947
rect 16601 254747 16801 254947
rect 17021 254747 17221 254947
rect 17441 254747 17641 254947
rect 17861 254747 18061 254947
rect 18281 254747 18481 254947
rect 18701 254747 18901 254947
rect 19121 254747 19321 254947
rect 19541 254747 19741 254947
rect 19961 254747 20161 254947
rect 20381 254747 20581 254947
rect 20801 254747 21001 254947
rect 21221 254747 21421 254947
rect 21641 254747 21841 254947
rect 22061 254747 22261 254947
rect 22481 254747 22681 254947
rect 22901 254747 23101 254947
rect 23321 254747 23521 254947
rect 23741 254747 23941 254947
rect 24161 254747 24361 254947
rect 24581 254747 24781 254947
rect 25001 254747 25201 254947
rect 25421 254747 25621 254947
rect 25841 254747 26041 254947
rect 26261 254747 26461 254947
rect 26681 254747 26881 254947
rect 27101 254747 27301 254947
rect -4180 243960 -4163 244041
rect -4163 243960 -3980 244041
rect -3771 243960 -3571 244041
rect -3351 243960 -3151 244041
rect -2931 243960 -2731 244041
rect -2511 243960 -2311 244041
rect -2091 243960 -1891 244041
rect -1671 243960 -1471 244041
rect -1251 243960 -1051 244041
rect -831 243960 -631 244041
rect -411 243960 -211 244041
rect 9 243960 209 244041
rect 429 243960 629 244041
rect 849 243960 1049 244041
rect 1269 243960 1469 244041
rect 1689 243960 1889 244041
rect 2109 243960 2309 244041
rect 2529 243960 2729 244041
rect 2949 243960 3149 244041
rect 3369 243960 3569 244041
rect 3789 243960 3989 244041
rect 4209 243960 4409 244041
rect 4629 243960 4829 244041
rect 5049 243960 5249 244041
rect 5469 243960 5669 244041
rect 5889 243960 6089 244041
rect 6309 243960 6509 244041
rect 6729 243960 6929 244041
rect 7149 243960 7349 244041
rect 7569 243960 7769 244041
rect 7989 243960 8189 244041
rect 8409 243960 8609 244041
rect 8829 243960 9029 244041
rect 9249 243960 9449 244041
rect 9669 243960 9869 244041
rect 10089 243960 10289 244041
rect 10509 243960 10709 244041
rect 10929 243960 11129 244041
rect 11349 243960 11549 244041
rect 11769 243960 11969 244041
rect 12189 243960 12389 244041
rect 12609 243960 12809 244041
rect 13029 243960 13229 244041
rect 13449 243960 13649 244041
rect 13869 243960 14069 244041
rect 14289 243960 14489 244041
rect 14709 243960 14909 244041
rect 15129 243960 15329 244041
rect 15549 243960 15749 244041
rect 15969 243960 16169 244041
rect 16389 243960 16589 244041
rect 16809 243960 17009 244041
rect 17229 243960 17429 244041
rect 17649 243960 17849 244041
rect 18069 243960 18269 244041
rect 18489 243960 18689 244041
rect 18909 243960 19109 244041
rect 19329 243960 19529 244041
rect 19749 243960 19949 244041
rect 20169 243960 20369 244041
rect 20589 243960 20789 244041
rect 21009 243960 21209 244041
rect 21429 243960 21629 244041
rect 21849 243960 22049 244041
rect 22269 243960 22469 244041
rect 22689 243960 22889 244041
rect 23109 243960 23309 244041
rect 23529 243960 23729 244041
rect 23949 243960 24149 244041
rect 24369 243960 24569 244041
rect 24789 243960 24989 244041
rect 25209 243960 25409 244041
rect 25629 243960 25829 244041
rect 26049 243960 26249 244041
rect 26469 243960 26669 244041
rect 26889 243960 27089 244041
rect -4180 243841 -3980 243960
rect -3771 243841 -3571 243960
rect -3351 243841 -3151 243960
rect -2931 243841 -2731 243960
rect -2511 243841 -2311 243960
rect -2091 243841 -1891 243960
rect -1671 243841 -1471 243960
rect -1251 243841 -1051 243960
rect -831 243841 -631 243960
rect -411 243841 -211 243960
rect 9 243841 209 243960
rect 429 243841 629 243960
rect 849 243841 1049 243960
rect 1269 243841 1469 243960
rect 1689 243841 1889 243960
rect 2109 243841 2309 243960
rect 2529 243841 2729 243960
rect 2949 243841 3149 243960
rect 3369 243841 3569 243960
rect 3789 243841 3989 243960
rect 4209 243841 4409 243960
rect 4629 243841 4829 243960
rect 5049 243841 5249 243960
rect 5469 243841 5669 243960
rect 5889 243841 6089 243960
rect 6309 243841 6509 243960
rect 6729 243841 6929 243960
rect 7149 243841 7349 243960
rect 7569 243841 7769 243960
rect 7989 243841 8189 243960
rect 8409 243841 8609 243960
rect 8829 243841 9029 243960
rect 9249 243841 9449 243960
rect 9669 243841 9869 243960
rect 10089 243841 10289 243960
rect 10509 243841 10709 243960
rect 10929 243841 11129 243960
rect 11349 243841 11549 243960
rect 11769 243841 11969 243960
rect 12189 243841 12389 243960
rect 12609 243841 12809 243960
rect 13029 243841 13229 243960
rect 13449 243841 13649 243960
rect 13869 243841 14069 243960
rect 14289 243841 14489 243960
rect 14709 243841 14909 243960
rect 15129 243841 15329 243960
rect 15549 243841 15749 243960
rect 15969 243841 16169 243960
rect 16389 243841 16589 243960
rect 16809 243841 17009 243960
rect 17229 243841 17429 243960
rect 17649 243841 17849 243960
rect 18069 243841 18269 243960
rect 18489 243841 18689 243960
rect 18909 243841 19109 243960
rect 19329 243841 19529 243960
rect 19749 243841 19949 243960
rect 20169 243841 20369 243960
rect 20589 243841 20789 243960
rect 21009 243841 21209 243960
rect 21429 243841 21629 243960
rect 21849 243841 22049 243960
rect 22269 243841 22469 243960
rect 22689 243841 22889 243960
rect 23109 243841 23309 243960
rect 23529 243841 23729 243960
rect 23949 243841 24149 243960
rect 24369 243841 24569 243960
rect 24789 243841 24989 243960
rect 25209 243841 25409 243960
rect 25629 243841 25829 243960
rect 26049 243841 26249 243960
rect 26469 243841 26669 243960
rect 26889 243841 27089 243960
rect 27414 243841 27614 244041
<< metal3 >>
rect -4189 264430 -3969 264435
rect -4189 264230 -4179 264430
rect -3979 264230 -3969 264430
rect -4189 264225 -3969 264230
rect -3780 264430 -3560 264435
rect -3780 264230 -3770 264430
rect -3570 264230 -3560 264430
rect -3780 264225 -3560 264230
rect -3360 264430 -3140 264435
rect -3360 264230 -3350 264430
rect -3150 264230 -3140 264430
rect -3360 264225 -3140 264230
rect -2940 264430 -2720 264435
rect -2940 264230 -2930 264430
rect -2730 264230 -2720 264430
rect -2940 264225 -2720 264230
rect -2520 264430 -2300 264435
rect -2520 264230 -2510 264430
rect -2310 264230 -2300 264430
rect -2520 264225 -2300 264230
rect -2100 264430 -1880 264435
rect -2100 264230 -2090 264430
rect -1890 264230 -1880 264430
rect -2100 264225 -1880 264230
rect -1680 264430 -1460 264435
rect -1680 264230 -1670 264430
rect -1470 264230 -1460 264430
rect -1680 264225 -1460 264230
rect -1260 264430 -1040 264435
rect -1260 264230 -1250 264430
rect -1050 264230 -1040 264430
rect -1260 264225 -1040 264230
rect -840 264430 -620 264435
rect -840 264230 -830 264430
rect -630 264230 -620 264430
rect -840 264225 -620 264230
rect -420 264430 -200 264435
rect -420 264230 -410 264430
rect -210 264230 -200 264430
rect -420 264225 -200 264230
rect 0 264430 220 264435
rect 0 264230 10 264430
rect 210 264230 220 264430
rect 0 264225 220 264230
rect 420 264430 640 264435
rect 420 264230 430 264430
rect 630 264230 640 264430
rect 420 264225 640 264230
rect 840 264430 1060 264435
rect 840 264230 850 264430
rect 1050 264230 1060 264430
rect 840 264225 1060 264230
rect 1260 264430 1480 264435
rect 1260 264230 1270 264430
rect 1470 264230 1480 264430
rect 1260 264225 1480 264230
rect 1680 264430 1900 264435
rect 1680 264230 1690 264430
rect 1890 264230 1900 264430
rect 1680 264225 1900 264230
rect 2100 264430 2320 264435
rect 2100 264230 2110 264430
rect 2310 264230 2320 264430
rect 2100 264225 2320 264230
rect 2520 264430 2740 264435
rect 2520 264230 2530 264430
rect 2730 264230 2740 264430
rect 2520 264225 2740 264230
rect 2940 264430 3160 264435
rect 2940 264230 2950 264430
rect 3150 264230 3160 264430
rect 2940 264225 3160 264230
rect 3360 264430 3580 264435
rect 3360 264230 3370 264430
rect 3570 264230 3580 264430
rect 3360 264225 3580 264230
rect 3780 264430 4000 264435
rect 3780 264230 3790 264430
rect 3990 264230 4000 264430
rect 3780 264225 4000 264230
rect 4200 264430 4420 264435
rect 4200 264230 4210 264430
rect 4410 264230 4420 264430
rect 4200 264225 4420 264230
rect 4620 264430 4840 264435
rect 4620 264230 4630 264430
rect 4830 264230 4840 264430
rect 4620 264225 4840 264230
rect 5040 264430 5260 264435
rect 5040 264230 5050 264430
rect 5250 264230 5260 264430
rect 5040 264225 5260 264230
rect 5460 264430 5680 264435
rect 5460 264230 5470 264430
rect 5670 264230 5680 264430
rect 5460 264225 5680 264230
rect 5880 264430 6100 264435
rect 5880 264230 5890 264430
rect 6090 264230 6100 264430
rect 5880 264225 6100 264230
rect 6300 264430 6520 264435
rect 6300 264230 6310 264430
rect 6510 264230 6520 264430
rect 6300 264225 6520 264230
rect 6720 264430 6940 264435
rect 6720 264230 6730 264430
rect 6930 264230 6940 264430
rect 6720 264225 6940 264230
rect 7140 264430 7360 264435
rect 7140 264230 7150 264430
rect 7350 264230 7360 264430
rect 7140 264225 7360 264230
rect 7560 264430 7780 264435
rect 7560 264230 7570 264430
rect 7770 264230 7780 264430
rect 7560 264225 7780 264230
rect 7980 264430 8200 264435
rect 7980 264230 7990 264430
rect 8190 264230 8200 264430
rect 7980 264225 8200 264230
rect 8400 264430 8620 264435
rect 8400 264230 8410 264430
rect 8610 264230 8620 264430
rect 8400 264225 8620 264230
rect 8820 264430 9040 264435
rect 8820 264230 8830 264430
rect 9030 264230 9040 264430
rect 8820 264225 9040 264230
rect 9240 264430 9460 264435
rect 9240 264230 9250 264430
rect 9450 264230 9460 264430
rect 9240 264225 9460 264230
rect 9660 264430 9880 264435
rect 9660 264230 9670 264430
rect 9870 264230 9880 264430
rect 9660 264225 9880 264230
rect 10080 264430 10300 264435
rect 10080 264230 10090 264430
rect 10290 264230 10300 264430
rect 10080 264225 10300 264230
rect 10500 264430 10720 264435
rect 10500 264230 10510 264430
rect 10710 264230 10720 264430
rect 10500 264225 10720 264230
rect 10920 264430 11140 264435
rect 10920 264230 10930 264430
rect 11130 264230 11140 264430
rect 10920 264225 11140 264230
rect 11340 264430 11560 264435
rect 11340 264230 11350 264430
rect 11550 264230 11560 264430
rect 11340 264225 11560 264230
rect 11760 264430 11980 264435
rect 11760 264230 11770 264430
rect 11970 264230 11980 264430
rect 11760 264225 11980 264230
rect 12180 264430 12400 264435
rect 12180 264230 12190 264430
rect 12390 264230 12400 264430
rect 12180 264225 12400 264230
rect 12600 264430 12820 264435
rect 12600 264230 12610 264430
rect 12810 264230 12820 264430
rect 12600 264225 12820 264230
rect 13020 264430 13240 264435
rect 13020 264230 13030 264430
rect 13230 264230 13240 264430
rect 13020 264225 13240 264230
rect 13440 264430 13660 264435
rect 13440 264230 13450 264430
rect 13650 264230 13660 264430
rect 13440 264225 13660 264230
rect 13860 264430 14080 264435
rect 13860 264230 13870 264430
rect 14070 264230 14080 264430
rect 13860 264225 14080 264230
rect 14280 264430 14500 264435
rect 14280 264230 14290 264430
rect 14490 264230 14500 264430
rect 14280 264225 14500 264230
rect 14700 264430 14920 264435
rect 14700 264230 14710 264430
rect 14910 264230 14920 264430
rect 14700 264225 14920 264230
rect 15120 264430 15340 264435
rect 15120 264230 15130 264430
rect 15330 264230 15340 264430
rect 15120 264225 15340 264230
rect 15540 264430 15760 264435
rect 15540 264230 15550 264430
rect 15750 264230 15760 264430
rect 15540 264225 15760 264230
rect 15960 264430 16180 264435
rect 15960 264230 15970 264430
rect 16170 264230 16180 264430
rect 15960 264225 16180 264230
rect 16380 264430 16600 264435
rect 16380 264230 16390 264430
rect 16590 264230 16600 264430
rect 16380 264225 16600 264230
rect 16800 264430 17020 264435
rect 16800 264230 16810 264430
rect 17010 264230 17020 264430
rect 16800 264225 17020 264230
rect 17220 264430 17440 264435
rect 17220 264230 17230 264430
rect 17430 264230 17440 264430
rect 17220 264225 17440 264230
rect 17640 264430 17860 264435
rect 17640 264230 17650 264430
rect 17850 264230 17860 264430
rect 17640 264225 17860 264230
rect 18060 264430 18280 264435
rect 18060 264230 18070 264430
rect 18270 264230 18280 264430
rect 18060 264225 18280 264230
rect 18480 264430 18700 264435
rect 18480 264230 18490 264430
rect 18690 264230 18700 264430
rect 18480 264225 18700 264230
rect 18900 264430 19120 264435
rect 18900 264230 18910 264430
rect 19110 264230 19120 264430
rect 18900 264225 19120 264230
rect 19320 264430 19540 264435
rect 19320 264230 19330 264430
rect 19530 264230 19540 264430
rect 19320 264225 19540 264230
rect 19740 264430 19960 264435
rect 19740 264230 19750 264430
rect 19950 264230 19960 264430
rect 19740 264225 19960 264230
rect 20160 264430 20380 264435
rect 20160 264230 20170 264430
rect 20370 264230 20380 264430
rect 20160 264225 20380 264230
rect 20580 264430 20800 264435
rect 20580 264230 20590 264430
rect 20790 264230 20800 264430
rect 20580 264225 20800 264230
rect 21000 264430 21220 264435
rect 21000 264230 21010 264430
rect 21210 264230 21220 264430
rect 21000 264225 21220 264230
rect 21420 264430 21640 264435
rect 21420 264230 21430 264430
rect 21630 264230 21640 264430
rect 21420 264225 21640 264230
rect 21840 264430 22060 264435
rect 21840 264230 21850 264430
rect 22050 264230 22060 264430
rect 21840 264225 22060 264230
rect 22260 264430 22480 264435
rect 22260 264230 22270 264430
rect 22470 264230 22480 264430
rect 22260 264225 22480 264230
rect 22680 264430 22900 264435
rect 22680 264230 22690 264430
rect 22890 264230 22900 264430
rect 22680 264225 22900 264230
rect 23100 264430 23320 264435
rect 23100 264230 23110 264430
rect 23310 264230 23320 264430
rect 23100 264225 23320 264230
rect 23520 264430 23740 264435
rect 23520 264230 23530 264430
rect 23730 264230 23740 264430
rect 23520 264225 23740 264230
rect 23940 264430 24160 264435
rect 23940 264230 23950 264430
rect 24150 264230 24160 264430
rect 23940 264225 24160 264230
rect 24360 264430 24580 264435
rect 24360 264230 24370 264430
rect 24570 264230 24580 264430
rect 24360 264225 24580 264230
rect 24780 264430 25000 264435
rect 24780 264230 24790 264430
rect 24990 264230 25000 264430
rect 24780 264225 25000 264230
rect 25200 264430 25420 264435
rect 25200 264230 25210 264430
rect 25410 264230 25420 264430
rect 25200 264225 25420 264230
rect 25620 264430 25840 264435
rect 25620 264230 25630 264430
rect 25830 264230 25840 264430
rect 25620 264225 25840 264230
rect 26040 264430 26260 264435
rect 26040 264230 26050 264430
rect 26250 264230 26260 264430
rect 26040 264225 26260 264230
rect 26460 264430 26680 264435
rect 26460 264230 26470 264430
rect 26670 264230 26680 264430
rect 26460 264225 26680 264230
rect 26880 264430 27100 264435
rect 26880 264230 26890 264430
rect 27090 264230 27100 264430
rect 26880 264225 27100 264230
rect 27300 264430 27520 264435
rect 27300 264230 27310 264430
rect 27510 264230 27520 264430
rect 27300 264225 27520 264230
rect -3990 261952 27457 261957
rect -3990 261752 -3980 261952
rect -3780 261752 -3560 261952
rect -3360 261752 -3140 261952
rect -2940 261752 -2720 261952
rect -2520 261752 -2300 261952
rect -2100 261752 -1880 261952
rect -1680 261752 -1460 261952
rect -1260 261752 -1040 261952
rect -840 261752 -620 261952
rect -420 261752 -200 261952
rect 0 261752 220 261952
rect 420 261752 640 261952
rect 840 261752 1060 261952
rect 1260 261752 1480 261952
rect 1680 261752 1900 261952
rect 2100 261752 2320 261952
rect 2520 261752 2740 261952
rect 2940 261752 3160 261952
rect 3360 261752 3580 261952
rect 3780 261752 4000 261952
rect 4200 261752 4420 261952
rect 4620 261752 4840 261952
rect 5040 261752 5260 261952
rect 5460 261752 5680 261952
rect 5880 261752 6100 261952
rect 6300 261752 6520 261952
rect 6720 261752 6940 261952
rect 7140 261752 7360 261952
rect 7560 261752 7780 261952
rect 7980 261752 8200 261952
rect 8400 261752 8620 261952
rect 8820 261752 9040 261952
rect 9240 261752 9460 261952
rect 9660 261752 9880 261952
rect 10080 261752 10300 261952
rect 10500 261752 10720 261952
rect 10920 261752 11140 261952
rect 11340 261752 11560 261952
rect 11760 261752 11980 261952
rect 12180 261752 12400 261952
rect 12600 261752 12820 261952
rect 13020 261752 13240 261952
rect 13440 261752 13660 261952
rect 13860 261752 14080 261952
rect 14280 261752 14500 261952
rect 14700 261752 14920 261952
rect 15120 261752 15340 261952
rect 15540 261752 15760 261952
rect 15960 261752 16180 261952
rect 16380 261752 16600 261952
rect 16800 261752 17020 261952
rect 17220 261752 17440 261952
rect 17640 261752 17860 261952
rect 18060 261752 18280 261952
rect 18480 261752 18700 261952
rect 18900 261752 19120 261952
rect 19320 261752 19540 261952
rect 19740 261752 19960 261952
rect 20160 261752 20380 261952
rect 20580 261752 20800 261952
rect 21000 261752 21220 261952
rect 21420 261752 21640 261952
rect 21840 261752 22060 261952
rect 22260 261752 22480 261952
rect 22680 261752 22900 261952
rect 23100 261752 23320 261952
rect 23520 261752 23740 261952
rect 23940 261752 24160 261952
rect 24360 261752 24580 261952
rect 24780 261752 25000 261952
rect 25200 261752 25420 261952
rect 25620 261752 25840 261952
rect 26040 261752 26260 261952
rect 26460 261752 26680 261952
rect 26880 261752 27100 261952
rect 27300 261752 27457 261952
rect -3990 254947 27457 261752
rect -3990 254747 -3979 254947
rect -3779 254747 -3559 254947
rect -3359 254747 -3139 254947
rect -2939 254747 -2719 254947
rect -2519 254747 -2299 254947
rect -2099 254747 -1879 254947
rect -1679 254747 -1459 254947
rect -1259 254747 -1039 254947
rect -839 254747 -619 254947
rect -419 254747 -199 254947
rect 1 254747 221 254947
rect 421 254747 641 254947
rect 841 254747 1061 254947
rect 1261 254747 1481 254947
rect 1681 254747 1901 254947
rect 2101 254747 2321 254947
rect 2521 254747 2741 254947
rect 2941 254747 3161 254947
rect 3361 254747 3581 254947
rect 3781 254747 4001 254947
rect 4201 254747 4421 254947
rect 4621 254747 4841 254947
rect 5041 254747 5261 254947
rect 5461 254747 5681 254947
rect 5881 254747 6101 254947
rect 6301 254747 6521 254947
rect 6721 254747 6941 254947
rect 7141 254747 7361 254947
rect 7561 254747 7781 254947
rect 7981 254747 8201 254947
rect 8401 254747 8621 254947
rect 8821 254747 9041 254947
rect 9241 254747 9461 254947
rect 9661 254747 9881 254947
rect 10081 254747 10301 254947
rect 10501 254747 10721 254947
rect 10921 254747 11141 254947
rect 11341 254747 11561 254947
rect 11761 254747 11981 254947
rect 12181 254747 12401 254947
rect 12601 254747 12821 254947
rect 13021 254747 13241 254947
rect 13441 254747 13661 254947
rect 13861 254747 14081 254947
rect 14281 254747 14501 254947
rect 14701 254747 14921 254947
rect 15121 254747 15341 254947
rect 15541 254747 15761 254947
rect 15961 254747 16181 254947
rect 16381 254747 16601 254947
rect 16801 254747 17021 254947
rect 17221 254747 17441 254947
rect 17641 254747 17861 254947
rect 18061 254747 18281 254947
rect 18481 254747 18701 254947
rect 18901 254747 19121 254947
rect 19321 254747 19541 254947
rect 19741 254747 19961 254947
rect 20161 254747 20381 254947
rect 20581 254747 20801 254947
rect 21001 254747 21221 254947
rect 21421 254747 21641 254947
rect 21841 254747 22061 254947
rect 22261 254747 22481 254947
rect 22681 254747 22901 254947
rect 23101 254747 23321 254947
rect 23521 254747 23741 254947
rect 23941 254747 24161 254947
rect 24361 254747 24581 254947
rect 24781 254747 25001 254947
rect 25201 254747 25421 254947
rect 25621 254747 25841 254947
rect 26041 254747 26261 254947
rect 26461 254747 26681 254947
rect 26881 254747 27101 254947
rect 27301 254747 27457 254947
rect -3990 254742 27457 254747
rect -4190 244041 -3970 244046
rect -4190 243841 -4180 244041
rect -3980 243841 -3970 244041
rect -4190 243836 -3970 243841
rect -3781 244041 -3561 244046
rect -3781 243841 -3771 244041
rect -3571 243841 -3561 244041
rect -3781 243836 -3561 243841
rect -3361 244041 -3141 244046
rect -3361 243841 -3351 244041
rect -3151 243841 -3141 244041
rect -3361 243836 -3141 243841
rect -2941 244041 -2721 244046
rect -2941 243841 -2931 244041
rect -2731 243841 -2721 244041
rect -2941 243836 -2721 243841
rect -2521 244041 -2301 244046
rect -2521 243841 -2511 244041
rect -2311 243841 -2301 244041
rect -2521 243836 -2301 243841
rect -2101 244041 -1881 244046
rect -2101 243841 -2091 244041
rect -1891 243841 -1881 244041
rect -2101 243836 -1881 243841
rect -1681 244041 -1461 244046
rect -1681 243841 -1671 244041
rect -1471 243841 -1461 244041
rect -1681 243836 -1461 243841
rect -1261 244041 -1041 244046
rect -1261 243841 -1251 244041
rect -1051 243841 -1041 244041
rect -1261 243836 -1041 243841
rect -841 244041 -621 244046
rect -841 243841 -831 244041
rect -631 243841 -621 244041
rect -841 243836 -621 243841
rect -421 244041 -201 244046
rect -421 243841 -411 244041
rect -211 243841 -201 244041
rect -421 243836 -201 243841
rect -1 244041 219 244046
rect -1 243841 9 244041
rect 209 243841 219 244041
rect -1 243836 219 243841
rect 419 244041 639 244046
rect 419 243841 429 244041
rect 629 243841 639 244041
rect 419 243836 639 243841
rect 839 244041 1059 244046
rect 839 243841 849 244041
rect 1049 243841 1059 244041
rect 839 243836 1059 243841
rect 1259 244041 1479 244046
rect 1259 243841 1269 244041
rect 1469 243841 1479 244041
rect 1259 243836 1479 243841
rect 1679 244041 1899 244046
rect 1679 243841 1689 244041
rect 1889 243841 1899 244041
rect 1679 243836 1899 243841
rect 2099 244041 2319 244046
rect 2099 243841 2109 244041
rect 2309 243841 2319 244041
rect 2099 243836 2319 243841
rect 2519 244041 2739 244046
rect 2519 243841 2529 244041
rect 2729 243841 2739 244041
rect 2519 243836 2739 243841
rect 2939 244041 3159 244046
rect 2939 243841 2949 244041
rect 3149 243841 3159 244041
rect 2939 243836 3159 243841
rect 3359 244041 3579 244046
rect 3359 243841 3369 244041
rect 3569 243841 3579 244041
rect 3359 243836 3579 243841
rect 3779 244041 3999 244046
rect 3779 243841 3789 244041
rect 3989 243841 3999 244041
rect 3779 243836 3999 243841
rect 4199 244041 4419 244046
rect 4199 243841 4209 244041
rect 4409 243841 4419 244041
rect 4199 243836 4419 243841
rect 4619 244041 4839 244046
rect 4619 243841 4629 244041
rect 4829 243841 4839 244041
rect 4619 243836 4839 243841
rect 5039 244041 5259 244046
rect 5039 243841 5049 244041
rect 5249 243841 5259 244041
rect 5039 243836 5259 243841
rect 5459 244041 5679 244046
rect 5459 243841 5469 244041
rect 5669 243841 5679 244041
rect 5459 243836 5679 243841
rect 5879 244041 6099 244046
rect 5879 243841 5889 244041
rect 6089 243841 6099 244041
rect 5879 243836 6099 243841
rect 6299 244041 6519 244046
rect 6299 243841 6309 244041
rect 6509 243841 6519 244041
rect 6299 243836 6519 243841
rect 6719 244041 6939 244046
rect 6719 243841 6729 244041
rect 6929 243841 6939 244041
rect 6719 243836 6939 243841
rect 7139 244041 7359 244046
rect 7139 243841 7149 244041
rect 7349 243841 7359 244041
rect 7139 243836 7359 243841
rect 7559 244041 7779 244046
rect 7559 243841 7569 244041
rect 7769 243841 7779 244041
rect 7559 243836 7779 243841
rect 7979 244041 8199 244046
rect 7979 243841 7989 244041
rect 8189 243841 8199 244041
rect 7979 243836 8199 243841
rect 8399 244041 8619 244046
rect 8399 243841 8409 244041
rect 8609 243841 8619 244041
rect 8399 243836 8619 243841
rect 8819 244041 9039 244046
rect 8819 243841 8829 244041
rect 9029 243841 9039 244041
rect 8819 243836 9039 243841
rect 9239 244041 9459 244046
rect 9239 243841 9249 244041
rect 9449 243841 9459 244041
rect 9239 243836 9459 243841
rect 9659 244041 9879 244046
rect 9659 243841 9669 244041
rect 9869 243841 9879 244041
rect 9659 243836 9879 243841
rect 10079 244041 10299 244046
rect 10079 243841 10089 244041
rect 10289 243841 10299 244041
rect 10079 243836 10299 243841
rect 10499 244041 10719 244046
rect 10499 243841 10509 244041
rect 10709 243841 10719 244041
rect 10499 243836 10719 243841
rect 10919 244041 11139 244046
rect 10919 243841 10929 244041
rect 11129 243841 11139 244041
rect 10919 243836 11139 243841
rect 11339 244041 11559 244046
rect 11339 243841 11349 244041
rect 11549 243841 11559 244041
rect 11339 243836 11559 243841
rect 11759 244041 11979 244046
rect 11759 243841 11769 244041
rect 11969 243841 11979 244041
rect 11759 243836 11979 243841
rect 12179 244041 12399 244046
rect 12179 243841 12189 244041
rect 12389 243841 12399 244041
rect 12179 243836 12399 243841
rect 12599 244041 12819 244046
rect 12599 243841 12609 244041
rect 12809 243841 12819 244041
rect 12599 243836 12819 243841
rect 13019 244041 13239 244046
rect 13019 243841 13029 244041
rect 13229 243841 13239 244041
rect 13019 243836 13239 243841
rect 13439 244041 13659 244046
rect 13439 243841 13449 244041
rect 13649 243841 13659 244041
rect 13439 243836 13659 243841
rect 13859 244041 14079 244046
rect 13859 243841 13869 244041
rect 14069 243841 14079 244041
rect 13859 243836 14079 243841
rect 14279 244041 14499 244046
rect 14279 243841 14289 244041
rect 14489 243841 14499 244041
rect 14279 243836 14499 243841
rect 14699 244041 14919 244046
rect 14699 243841 14709 244041
rect 14909 243841 14919 244041
rect 14699 243836 14919 243841
rect 15119 244041 15339 244046
rect 15119 243841 15129 244041
rect 15329 243841 15339 244041
rect 15119 243836 15339 243841
rect 15539 244041 15759 244046
rect 15539 243841 15549 244041
rect 15749 243841 15759 244041
rect 15539 243836 15759 243841
rect 15959 244041 16179 244046
rect 15959 243841 15969 244041
rect 16169 243841 16179 244041
rect 15959 243836 16179 243841
rect 16379 244041 16599 244046
rect 16379 243841 16389 244041
rect 16589 243841 16599 244041
rect 16379 243836 16599 243841
rect 16799 244041 17019 244046
rect 16799 243841 16809 244041
rect 17009 243841 17019 244041
rect 16799 243836 17019 243841
rect 17219 244041 17439 244046
rect 17219 243841 17229 244041
rect 17429 243841 17439 244041
rect 17219 243836 17439 243841
rect 17639 244041 17859 244046
rect 17639 243841 17649 244041
rect 17849 243841 17859 244041
rect 17639 243836 17859 243841
rect 18059 244041 18279 244046
rect 18059 243841 18069 244041
rect 18269 243841 18279 244041
rect 18059 243836 18279 243841
rect 18479 244041 18699 244046
rect 18479 243841 18489 244041
rect 18689 243841 18699 244041
rect 18479 243836 18699 243841
rect 18899 244041 19119 244046
rect 18899 243841 18909 244041
rect 19109 243841 19119 244041
rect 18899 243836 19119 243841
rect 19319 244041 19539 244046
rect 19319 243841 19329 244041
rect 19529 243841 19539 244041
rect 19319 243836 19539 243841
rect 19739 244041 19959 244046
rect 19739 243841 19749 244041
rect 19949 243841 19959 244041
rect 19739 243836 19959 243841
rect 20159 244041 20379 244046
rect 20159 243841 20169 244041
rect 20369 243841 20379 244041
rect 20159 243836 20379 243841
rect 20579 244041 20799 244046
rect 20579 243841 20589 244041
rect 20789 243841 20799 244041
rect 20579 243836 20799 243841
rect 20999 244041 21219 244046
rect 20999 243841 21009 244041
rect 21209 243841 21219 244041
rect 20999 243836 21219 243841
rect 21419 244041 21639 244046
rect 21419 243841 21429 244041
rect 21629 243841 21639 244041
rect 21419 243836 21639 243841
rect 21839 244041 22059 244046
rect 21839 243841 21849 244041
rect 22049 243841 22059 244041
rect 21839 243836 22059 243841
rect 22259 244041 22479 244046
rect 22259 243841 22269 244041
rect 22469 243841 22479 244041
rect 22259 243836 22479 243841
rect 22679 244041 22899 244046
rect 22679 243841 22689 244041
rect 22889 243841 22899 244041
rect 22679 243836 22899 243841
rect 23099 244041 23319 244046
rect 23099 243841 23109 244041
rect 23309 243841 23319 244041
rect 23099 243836 23319 243841
rect 23519 244041 23739 244046
rect 23519 243841 23529 244041
rect 23729 243841 23739 244041
rect 23519 243836 23739 243841
rect 23939 244041 24159 244046
rect 23939 243841 23949 244041
rect 24149 243841 24159 244041
rect 23939 243836 24159 243841
rect 24359 244041 24579 244046
rect 24359 243841 24369 244041
rect 24569 243841 24579 244041
rect 24359 243836 24579 243841
rect 24779 244041 24999 244046
rect 24779 243841 24789 244041
rect 24989 243841 24999 244041
rect 24779 243836 24999 243841
rect 25199 244041 25419 244046
rect 25199 243841 25209 244041
rect 25409 243841 25419 244041
rect 25199 243836 25419 243841
rect 25619 244041 25839 244046
rect 25619 243841 25629 244041
rect 25829 243841 25839 244041
rect 25619 243836 25839 243841
rect 26039 244041 26259 244046
rect 26039 243841 26049 244041
rect 26249 243841 26259 244041
rect 26039 243836 26259 243841
rect 26459 244041 26679 244046
rect 26459 243841 26469 244041
rect 26669 243841 26679 244041
rect 26459 243836 26679 243841
rect 26879 244041 27099 244046
rect 26879 243841 26889 244041
rect 27089 243841 27099 244041
rect 26879 243836 27099 243841
rect 27404 244041 27624 244046
rect 27404 243841 27414 244041
rect 27614 243841 27624 244041
rect 27404 243836 27624 243841
<< via3 >>
rect -4179 264230 -3979 264430
rect -3770 264230 -3570 264430
rect -3350 264230 -3150 264430
rect -2930 264230 -2730 264430
rect -2510 264230 -2310 264430
rect -2090 264230 -1890 264430
rect -1670 264230 -1470 264430
rect -1250 264230 -1050 264430
rect -830 264230 -630 264430
rect -410 264230 -210 264430
rect 10 264230 210 264430
rect 430 264230 630 264430
rect 850 264230 1050 264430
rect 1270 264230 1470 264430
rect 1690 264230 1890 264430
rect 2110 264230 2310 264430
rect 2530 264230 2730 264430
rect 2950 264230 3150 264430
rect 3370 264230 3570 264430
rect 3790 264230 3990 264430
rect 4210 264230 4410 264430
rect 4630 264230 4830 264430
rect 5050 264230 5250 264430
rect 5470 264230 5670 264430
rect 5890 264230 6090 264430
rect 6310 264230 6510 264430
rect 6730 264230 6930 264430
rect 7150 264230 7350 264430
rect 7570 264230 7770 264430
rect 7990 264230 8190 264430
rect 8410 264230 8610 264430
rect 8830 264230 9030 264430
rect 9250 264230 9450 264430
rect 9670 264230 9870 264430
rect 10090 264230 10290 264430
rect 10510 264230 10710 264430
rect 10930 264230 11130 264430
rect 11350 264230 11550 264430
rect 11770 264230 11970 264430
rect 12190 264230 12390 264430
rect 12610 264230 12810 264430
rect 13030 264230 13230 264430
rect 13450 264230 13650 264430
rect 13870 264230 14070 264430
rect 14290 264230 14490 264430
rect 14710 264230 14910 264430
rect 15130 264230 15330 264430
rect 15550 264230 15750 264430
rect 15970 264230 16170 264430
rect 16390 264230 16590 264430
rect 16810 264230 17010 264430
rect 17230 264230 17430 264430
rect 17650 264230 17850 264430
rect 18070 264230 18270 264430
rect 18490 264230 18690 264430
rect 18910 264230 19110 264430
rect 19330 264230 19530 264430
rect 19750 264230 19950 264430
rect 20170 264230 20370 264430
rect 20590 264230 20790 264430
rect 21010 264230 21210 264430
rect 21430 264230 21630 264430
rect 21850 264230 22050 264430
rect 22270 264230 22470 264430
rect 22690 264230 22890 264430
rect 23110 264230 23310 264430
rect 23530 264230 23730 264430
rect 23950 264230 24150 264430
rect 24370 264230 24570 264430
rect 24790 264230 24990 264430
rect 25210 264230 25410 264430
rect 25630 264230 25830 264430
rect 26050 264230 26250 264430
rect 26470 264230 26670 264430
rect 26890 264230 27090 264430
rect 27310 264230 27510 264430
rect -4180 243841 -3980 244041
rect -3771 243841 -3571 244041
rect -3351 243841 -3151 244041
rect -2931 243841 -2731 244041
rect -2511 243841 -2311 244041
rect -2091 243841 -1891 244041
rect -1671 243841 -1471 244041
rect -1251 243841 -1051 244041
rect -831 243841 -631 244041
rect -411 243841 -211 244041
rect 9 243841 209 244041
rect 429 243841 629 244041
rect 849 243841 1049 244041
rect 1269 243841 1469 244041
rect 1689 243841 1889 244041
rect 2109 243841 2309 244041
rect 2529 243841 2729 244041
rect 2949 243841 3149 244041
rect 3369 243841 3569 244041
rect 3789 243841 3989 244041
rect 4209 243841 4409 244041
rect 4629 243841 4829 244041
rect 5049 243841 5249 244041
rect 5469 243841 5669 244041
rect 5889 243841 6089 244041
rect 6309 243841 6509 244041
rect 6729 243841 6929 244041
rect 7149 243841 7349 244041
rect 7569 243841 7769 244041
rect 7989 243841 8189 244041
rect 8409 243841 8609 244041
rect 8829 243841 9029 244041
rect 9249 243841 9449 244041
rect 9669 243841 9869 244041
rect 10089 243841 10289 244041
rect 10509 243841 10709 244041
rect 10929 243841 11129 244041
rect 11349 243841 11549 244041
rect 11769 243841 11969 244041
rect 12189 243841 12389 244041
rect 12609 243841 12809 244041
rect 13029 243841 13229 244041
rect 13449 243841 13649 244041
rect 13869 243841 14069 244041
rect 14289 243841 14489 244041
rect 14709 243841 14909 244041
rect 15129 243841 15329 244041
rect 15549 243841 15749 244041
rect 15969 243841 16169 244041
rect 16389 243841 16589 244041
rect 16809 243841 17009 244041
rect 17229 243841 17429 244041
rect 17649 243841 17849 244041
rect 18069 243841 18269 244041
rect 18489 243841 18689 244041
rect 18909 243841 19109 244041
rect 19329 243841 19529 244041
rect 19749 243841 19949 244041
rect 20169 243841 20369 244041
rect 20589 243841 20789 244041
rect 21009 243841 21209 244041
rect 21429 243841 21629 244041
rect 21849 243841 22049 244041
rect 22269 243841 22469 244041
rect 22689 243841 22889 244041
rect 23109 243841 23309 244041
rect 23529 243841 23729 244041
rect 23949 243841 24149 244041
rect 24369 243841 24569 244041
rect 24789 243841 24989 244041
rect 25209 243841 25409 244041
rect 25629 243841 25829 244041
rect 26049 243841 26249 244041
rect 26469 243841 26669 244041
rect 26889 243841 27089 244041
rect 27414 243841 27614 244041
<< metal4 >>
rect -4180 264430 27520 265028
rect -4180 264230 -4179 264430
rect -3979 264230 -3770 264430
rect -3570 264230 -3350 264430
rect -3150 264230 -2930 264430
rect -2730 264230 -2510 264430
rect -2310 264230 -2090 264430
rect -1890 264230 -1670 264430
rect -1470 264230 -1250 264430
rect -1050 264230 -830 264430
rect -630 264230 -410 264430
rect -210 264230 10 264430
rect 210 264230 430 264430
rect 630 264230 850 264430
rect 1050 264230 1270 264430
rect 1470 264230 1690 264430
rect 1890 264230 2110 264430
rect 2310 264230 2530 264430
rect 2730 264230 2950 264430
rect 3150 264230 3370 264430
rect 3570 264230 3790 264430
rect 3990 264230 4210 264430
rect 4410 264230 4630 264430
rect 4830 264230 5050 264430
rect 5250 264230 5470 264430
rect 5670 264230 5890 264430
rect 6090 264230 6310 264430
rect 6510 264230 6730 264430
rect 6930 264230 7150 264430
rect 7350 264230 7570 264430
rect 7770 264230 7990 264430
rect 8190 264230 8410 264430
rect 8610 264230 8830 264430
rect 9030 264230 9250 264430
rect 9450 264230 9670 264430
rect 9870 264230 10090 264430
rect 10290 264230 10510 264430
rect 10710 264230 10930 264430
rect 11130 264230 11350 264430
rect 11550 264230 11770 264430
rect 11970 264230 12190 264430
rect 12390 264230 12610 264430
rect 12810 264230 13030 264430
rect 13230 264230 13450 264430
rect 13650 264230 13870 264430
rect 14070 264230 14290 264430
rect 14490 264230 14710 264430
rect 14910 264230 15130 264430
rect 15330 264230 15550 264430
rect 15750 264230 15970 264430
rect 16170 264230 16390 264430
rect 16590 264230 16810 264430
rect 17010 264230 17230 264430
rect 17430 264230 17650 264430
rect 17850 264230 18070 264430
rect 18270 264230 18490 264430
rect 18690 264230 18910 264430
rect 19110 264230 19330 264430
rect 19530 264230 19750 264430
rect 19950 264230 20170 264430
rect 20370 264230 20590 264430
rect 20790 264230 21010 264430
rect 21210 264230 21430 264430
rect 21630 264230 21850 264430
rect 22050 264230 22270 264430
rect 22470 264230 22690 264430
rect 22890 264230 23110 264430
rect 23310 264230 23530 264430
rect 23730 264230 23950 264430
rect 24150 264230 24370 264430
rect 24570 264230 24790 264430
rect 24990 264230 25210 264430
rect 25410 264230 25630 264430
rect 25830 264230 26050 264430
rect 26250 264230 26470 264430
rect 26670 264230 26890 264430
rect 27090 264230 27310 264430
rect 27510 264230 27520 264430
rect -4180 264229 27520 264230
rect -4142 264225 27520 264229
rect -4181 244041 27615 244042
rect -4181 243841 -4180 244041
rect -3980 243841 -3771 244041
rect -3571 243841 -3351 244041
rect -3151 243841 -2931 244041
rect -2731 243841 -2511 244041
rect -2311 243841 -2091 244041
rect -1891 243841 -1671 244041
rect -1471 243841 -1251 244041
rect -1051 243841 -831 244041
rect -631 243841 -411 244041
rect -211 243841 9 244041
rect 209 243841 429 244041
rect 629 243841 849 244041
rect 1049 243841 1269 244041
rect 1469 243841 1689 244041
rect 1889 243841 2109 244041
rect 2309 243841 2529 244041
rect 2729 243841 2949 244041
rect 3149 243841 3369 244041
rect 3569 243841 3789 244041
rect 3989 243841 4209 244041
rect 4409 243841 4629 244041
rect 4829 243841 5049 244041
rect 5249 243841 5469 244041
rect 5669 243841 5889 244041
rect 6089 243841 6309 244041
rect 6509 243841 6729 244041
rect 6929 243841 7149 244041
rect 7349 243841 7569 244041
rect 7769 243841 7989 244041
rect 8189 243841 8409 244041
rect 8609 243841 8829 244041
rect 9029 243841 9249 244041
rect 9449 243841 9669 244041
rect 9869 243841 10089 244041
rect 10289 243841 10509 244041
rect 10709 243841 10929 244041
rect 11129 243841 11349 244041
rect 11549 243841 11769 244041
rect 11969 243841 12189 244041
rect 12389 243841 12609 244041
rect 12809 243841 13029 244041
rect 13229 243841 13449 244041
rect 13649 243841 13869 244041
rect 14069 243841 14289 244041
rect 14489 243841 14709 244041
rect 14909 243841 15129 244041
rect 15329 243841 15549 244041
rect 15749 243841 15969 244041
rect 16169 243841 16389 244041
rect 16589 243841 16809 244041
rect 17009 243841 17229 244041
rect 17429 243841 17649 244041
rect 17849 243841 18069 244041
rect 18269 243841 18489 244041
rect 18689 243841 18909 244041
rect 19109 243841 19329 244041
rect 19529 243841 19749 244041
rect 19949 243841 20169 244041
rect 20369 243841 20589 244041
rect 20789 243841 21009 244041
rect 21209 243841 21429 244041
rect 21629 243841 21849 244041
rect 22049 243841 22269 244041
rect 22469 243841 22689 244041
rect 22889 243841 23109 244041
rect 23309 243841 23529 244041
rect 23729 243841 23949 244041
rect 24149 243841 24369 244041
rect 24569 243841 24789 244041
rect 24989 243841 25209 244041
rect 25409 243841 25629 244041
rect 25829 243841 26049 244041
rect 26249 243841 26469 244041
rect 26669 243841 26889 244041
rect 27089 243841 27414 244041
rect 27614 243841 27615 244041
rect -4181 243446 27615 243841
<< labels >>
flabel metal3 21719 257630 21719 257630 0 FreeSans 8000 0 0 0 out_p
port 4 nsew
flabel metal1 -4399 263315 -4399 263315 0 FreeSans 8000 0 0 0 vp_n
port 2 nsew
flabel metal1 -4493 249296 -4493 249296 0 FreeSans 8000 0 0 0 vp_p
port 1 nsew
<< end >>
