magic
tech sky130A
magscale 1 2
timestamp 1629189150
<< nwell >>
rect -703 -859 11421 1251
rect 785 -5483 3981 -1137
<< pwell >>
rect 5949 -4589 6351 -3293
rect 785 -7705 9933 -5831
<< pmoslvt >>
rect -507 632 -307 1032
rect -135 632 65 1032
rect 237 632 437 1032
rect 609 632 809 1032
rect 981 632 1181 1032
rect 1353 632 1553 1032
rect 1725 632 1925 1032
rect 2097 632 2297 1032
rect 2469 632 2669 1032
rect 2841 632 3041 1032
rect 3213 632 3413 1032
rect 3585 632 3785 1032
rect 3957 632 4157 1032
rect 4329 632 4529 1032
rect 4701 632 4901 1032
rect 5073 632 5273 1032
rect 5445 632 5645 1032
rect 5817 632 6017 1032
rect 6189 632 6389 1032
rect 6561 632 6761 1032
rect 6933 632 7133 1032
rect 7305 632 7505 1032
rect 7677 632 7877 1032
rect 8049 632 8249 1032
rect 8421 632 8621 1032
rect 8793 632 8993 1032
rect 9165 632 9365 1032
rect 9537 632 9737 1032
rect 9909 632 10109 1032
rect 10281 632 10481 1032
rect 10653 632 10853 1032
rect 11025 632 11225 1032
rect -507 -4 -307 396
rect -135 -4 65 396
rect 237 -4 437 396
rect 609 -4 809 396
rect 981 -4 1181 396
rect 1353 -4 1553 396
rect 1725 -4 1925 396
rect 2097 -4 2297 396
rect 2469 -4 2669 396
rect 2841 -4 3041 396
rect 3213 -4 3413 396
rect 3585 -4 3785 396
rect 3957 -4 4157 396
rect 4329 -4 4529 396
rect 4701 -4 4901 396
rect 5073 -4 5273 396
rect 5445 -4 5645 396
rect 5817 -4 6017 396
rect 6189 -4 6389 396
rect 6561 -4 6761 396
rect 6933 -4 7133 396
rect 7305 -4 7505 396
rect 7677 -4 7877 396
rect 8049 -4 8249 396
rect 8421 -4 8621 396
rect 8793 -4 8993 396
rect 9165 -4 9365 396
rect 9537 -4 9737 396
rect 9909 -4 10109 396
rect 10281 -4 10481 396
rect 10653 -4 10853 396
rect 11025 -4 11225 396
rect -507 -640 -307 -240
rect -135 -640 65 -240
rect 237 -640 437 -240
rect 609 -640 809 -240
rect 981 -640 1181 -240
rect 1353 -640 1553 -240
rect 1725 -640 1925 -240
rect 2097 -640 2297 -240
rect 2469 -640 2669 -240
rect 2841 -640 3041 -240
rect 3213 -640 3413 -240
rect 3585 -640 3785 -240
rect 3957 -640 4157 -240
rect 4329 -640 4529 -240
rect 4701 -640 4901 -240
rect 5073 -640 5273 -240
rect 5445 -640 5645 -240
rect 5817 -640 6017 -240
rect 6189 -640 6389 -240
rect 6561 -640 6761 -240
rect 6933 -640 7133 -240
rect 7305 -640 7505 -240
rect 7677 -640 7877 -240
rect 8049 -640 8249 -240
rect 8421 -640 8621 -240
rect 8793 -640 8993 -240
rect 9165 -640 9365 -240
rect 9537 -640 9737 -240
rect 9909 -640 10109 -240
rect 10281 -640 10481 -240
rect 10653 -640 10853 -240
rect 11025 -640 11225 -240
rect 981 -2156 1181 -1356
rect 1353 -2156 1553 -1356
rect 1725 -2156 1925 -1356
rect 2097 -2156 2297 -1356
rect 2469 -2156 2669 -1356
rect 2841 -2156 3041 -1356
rect 3213 -2156 3413 -1356
rect 3585 -2156 3785 -1356
rect 981 -3192 1181 -2392
rect 1353 -3192 1553 -2392
rect 1725 -3192 1925 -2392
rect 2097 -3192 2297 -2392
rect 2469 -3192 2669 -2392
rect 2841 -3192 3041 -2392
rect 3213 -3192 3413 -2392
rect 3585 -3192 3785 -2392
rect 981 -4228 1181 -3428
rect 1353 -4228 1553 -3428
rect 1725 -4228 1925 -3428
rect 2097 -4228 2297 -3428
rect 2469 -4228 2669 -3428
rect 2841 -4228 3041 -3428
rect 3213 -4228 3413 -3428
rect 3585 -4228 3785 -3428
rect 981 -5264 1181 -4464
rect 1353 -5264 1553 -4464
rect 1725 -5264 1925 -4464
rect 2097 -5264 2297 -4464
rect 2469 -5264 2669 -4464
rect 2841 -5264 3041 -4464
rect 3213 -5264 3413 -4464
rect 3585 -5264 3785 -4464
<< nmoslvt >>
rect 981 -6241 1181 -6041
rect 1353 -6241 1553 -6041
rect 1725 -6241 1925 -6041
rect 2097 -6241 2297 -6041
rect 2469 -6241 2669 -6041
rect 2841 -6241 3041 -6041
rect 3213 -6241 3413 -6041
rect 3585 -6241 3785 -6041
rect 3957 -6241 4157 -6041
rect 4329 -6241 4529 -6041
rect 4701 -6241 4901 -6041
rect 5073 -6241 5273 -6041
rect 5445 -6241 5645 -6041
rect 5817 -6241 6017 -6041
rect 6189 -6241 6389 -6041
rect 6561 -6241 6761 -6041
rect 6933 -6241 7133 -6041
rect 7305 -6241 7505 -6041
rect 7677 -6241 7877 -6041
rect 8049 -6241 8249 -6041
rect 8421 -6241 8621 -6041
rect 8793 -6241 8993 -6041
rect 9165 -6241 9365 -6041
rect 9537 -6241 9737 -6041
rect 981 -6659 1181 -6459
rect 1353 -6659 1553 -6459
rect 1725 -6659 1925 -6459
rect 2097 -6659 2297 -6459
rect 2469 -6659 2669 -6459
rect 2841 -6659 3041 -6459
rect 3213 -6659 3413 -6459
rect 3585 -6659 3785 -6459
rect 3957 -6659 4157 -6459
rect 4329 -6659 4529 -6459
rect 4701 -6659 4901 -6459
rect 5073 -6659 5273 -6459
rect 5445 -6659 5645 -6459
rect 5817 -6659 6017 -6459
rect 6189 -6659 6389 -6459
rect 6561 -6659 6761 -6459
rect 6933 -6659 7133 -6459
rect 7305 -6659 7505 -6459
rect 7677 -6659 7877 -6459
rect 8049 -6659 8249 -6459
rect 8421 -6659 8621 -6459
rect 8793 -6659 8993 -6459
rect 9165 -6659 9365 -6459
rect 9537 -6659 9737 -6459
rect 981 -7077 1181 -6877
rect 1353 -7077 1553 -6877
rect 1725 -7077 1925 -6877
rect 2097 -7077 2297 -6877
rect 2469 -7077 2669 -6877
rect 2841 -7077 3041 -6877
rect 3213 -7077 3413 -6877
rect 3585 -7077 3785 -6877
rect 3957 -7077 4157 -6877
rect 4329 -7077 4529 -6877
rect 4701 -7077 4901 -6877
rect 5073 -7077 5273 -6877
rect 5445 -7077 5645 -6877
rect 5817 -7077 6017 -6877
rect 6189 -7077 6389 -6877
rect 6561 -7077 6761 -6877
rect 6933 -7077 7133 -6877
rect 7305 -7077 7505 -6877
rect 7677 -7077 7877 -6877
rect 8049 -7077 8249 -6877
rect 8421 -7077 8621 -6877
rect 8793 -7077 8993 -6877
rect 9165 -7077 9365 -6877
rect 9537 -7077 9737 -6877
rect 981 -7495 1181 -7295
rect 1353 -7495 1553 -7295
rect 1725 -7495 1925 -7295
rect 2097 -7495 2297 -7295
rect 2469 -7495 2669 -7295
rect 2841 -7495 3041 -7295
rect 3213 -7495 3413 -7295
rect 3585 -7495 3785 -7295
rect 3957 -7495 4157 -7295
rect 4329 -7495 4529 -7295
rect 4701 -7495 4901 -7295
rect 5073 -7495 5273 -7295
rect 5445 -7495 5645 -7295
rect 5817 -7495 6017 -7295
rect 6189 -7495 6389 -7295
rect 6561 -7495 6761 -7295
rect 6933 -7495 7133 -7295
rect 7305 -7495 7505 -7295
rect 7677 -7495 7877 -7295
rect 8049 -7495 8249 -7295
rect 8421 -7495 8621 -7295
rect 8793 -7495 8993 -7295
rect 9165 -7495 9365 -7295
rect 9537 -7495 9737 -7295
<< ndiff >>
rect 923 -6053 981 -6041
rect 923 -6229 935 -6053
rect 969 -6229 981 -6053
rect 923 -6241 981 -6229
rect 1181 -6053 1239 -6041
rect 1181 -6229 1193 -6053
rect 1227 -6229 1239 -6053
rect 1181 -6241 1239 -6229
rect 1295 -6053 1353 -6041
rect 1295 -6229 1307 -6053
rect 1341 -6229 1353 -6053
rect 1295 -6241 1353 -6229
rect 1553 -6053 1611 -6041
rect 1553 -6229 1565 -6053
rect 1599 -6229 1611 -6053
rect 1553 -6241 1611 -6229
rect 1667 -6053 1725 -6041
rect 1667 -6229 1679 -6053
rect 1713 -6229 1725 -6053
rect 1667 -6241 1725 -6229
rect 1925 -6053 1983 -6041
rect 1925 -6229 1937 -6053
rect 1971 -6229 1983 -6053
rect 1925 -6241 1983 -6229
rect 2039 -6053 2097 -6041
rect 2039 -6229 2051 -6053
rect 2085 -6229 2097 -6053
rect 2039 -6241 2097 -6229
rect 2297 -6053 2355 -6041
rect 2297 -6229 2309 -6053
rect 2343 -6229 2355 -6053
rect 2297 -6241 2355 -6229
rect 2411 -6053 2469 -6041
rect 2411 -6229 2423 -6053
rect 2457 -6229 2469 -6053
rect 2411 -6241 2469 -6229
rect 2669 -6053 2727 -6041
rect 2669 -6229 2681 -6053
rect 2715 -6229 2727 -6053
rect 2669 -6241 2727 -6229
rect 2783 -6053 2841 -6041
rect 2783 -6229 2795 -6053
rect 2829 -6229 2841 -6053
rect 2783 -6241 2841 -6229
rect 3041 -6053 3099 -6041
rect 3041 -6229 3053 -6053
rect 3087 -6229 3099 -6053
rect 3041 -6241 3099 -6229
rect 3155 -6053 3213 -6041
rect 3155 -6229 3167 -6053
rect 3201 -6229 3213 -6053
rect 3155 -6241 3213 -6229
rect 3413 -6053 3471 -6041
rect 3413 -6229 3425 -6053
rect 3459 -6229 3471 -6053
rect 3413 -6241 3471 -6229
rect 3527 -6053 3585 -6041
rect 3527 -6229 3539 -6053
rect 3573 -6229 3585 -6053
rect 3527 -6241 3585 -6229
rect 3785 -6053 3843 -6041
rect 3785 -6229 3797 -6053
rect 3831 -6229 3843 -6053
rect 3785 -6241 3843 -6229
rect 3899 -6053 3957 -6041
rect 3899 -6229 3911 -6053
rect 3945 -6229 3957 -6053
rect 3899 -6241 3957 -6229
rect 4157 -6053 4215 -6041
rect 4157 -6229 4169 -6053
rect 4203 -6229 4215 -6053
rect 4157 -6241 4215 -6229
rect 4271 -6053 4329 -6041
rect 4271 -6229 4283 -6053
rect 4317 -6229 4329 -6053
rect 4271 -6241 4329 -6229
rect 4529 -6053 4587 -6041
rect 4529 -6229 4541 -6053
rect 4575 -6229 4587 -6053
rect 4529 -6241 4587 -6229
rect 4643 -6053 4701 -6041
rect 4643 -6229 4655 -6053
rect 4689 -6229 4701 -6053
rect 4643 -6241 4701 -6229
rect 4901 -6053 4959 -6041
rect 4901 -6229 4913 -6053
rect 4947 -6229 4959 -6053
rect 4901 -6241 4959 -6229
rect 5015 -6053 5073 -6041
rect 5015 -6229 5027 -6053
rect 5061 -6229 5073 -6053
rect 5015 -6241 5073 -6229
rect 5273 -6053 5331 -6041
rect 5273 -6229 5285 -6053
rect 5319 -6229 5331 -6053
rect 5273 -6241 5331 -6229
rect 5387 -6053 5445 -6041
rect 5387 -6229 5399 -6053
rect 5433 -6229 5445 -6053
rect 5387 -6241 5445 -6229
rect 5645 -6053 5703 -6041
rect 5645 -6229 5657 -6053
rect 5691 -6229 5703 -6053
rect 5645 -6241 5703 -6229
rect 5759 -6053 5817 -6041
rect 5759 -6229 5771 -6053
rect 5805 -6229 5817 -6053
rect 5759 -6241 5817 -6229
rect 6017 -6053 6075 -6041
rect 6017 -6229 6029 -6053
rect 6063 -6229 6075 -6053
rect 6017 -6241 6075 -6229
rect 6131 -6053 6189 -6041
rect 6131 -6229 6143 -6053
rect 6177 -6229 6189 -6053
rect 6131 -6241 6189 -6229
rect 6389 -6053 6447 -6041
rect 6389 -6229 6401 -6053
rect 6435 -6229 6447 -6053
rect 6389 -6241 6447 -6229
rect 6503 -6053 6561 -6041
rect 6503 -6229 6515 -6053
rect 6549 -6229 6561 -6053
rect 6503 -6241 6561 -6229
rect 6761 -6053 6819 -6041
rect 6761 -6229 6773 -6053
rect 6807 -6229 6819 -6053
rect 6761 -6241 6819 -6229
rect 6875 -6053 6933 -6041
rect 6875 -6229 6887 -6053
rect 6921 -6229 6933 -6053
rect 6875 -6241 6933 -6229
rect 7133 -6053 7191 -6041
rect 7133 -6229 7145 -6053
rect 7179 -6229 7191 -6053
rect 7133 -6241 7191 -6229
rect 7247 -6053 7305 -6041
rect 7247 -6229 7259 -6053
rect 7293 -6229 7305 -6053
rect 7247 -6241 7305 -6229
rect 7505 -6053 7563 -6041
rect 7505 -6229 7517 -6053
rect 7551 -6229 7563 -6053
rect 7505 -6241 7563 -6229
rect 7619 -6053 7677 -6041
rect 7619 -6229 7631 -6053
rect 7665 -6229 7677 -6053
rect 7619 -6241 7677 -6229
rect 7877 -6053 7935 -6041
rect 7877 -6229 7889 -6053
rect 7923 -6229 7935 -6053
rect 7877 -6241 7935 -6229
rect 7991 -6053 8049 -6041
rect 7991 -6229 8003 -6053
rect 8037 -6229 8049 -6053
rect 7991 -6241 8049 -6229
rect 8249 -6053 8307 -6041
rect 8249 -6229 8261 -6053
rect 8295 -6229 8307 -6053
rect 8249 -6241 8307 -6229
rect 8363 -6053 8421 -6041
rect 8363 -6229 8375 -6053
rect 8409 -6229 8421 -6053
rect 8363 -6241 8421 -6229
rect 8621 -6053 8679 -6041
rect 8621 -6229 8633 -6053
rect 8667 -6229 8679 -6053
rect 8621 -6241 8679 -6229
rect 8735 -6053 8793 -6041
rect 8735 -6229 8747 -6053
rect 8781 -6229 8793 -6053
rect 8735 -6241 8793 -6229
rect 8993 -6053 9051 -6041
rect 8993 -6229 9005 -6053
rect 9039 -6229 9051 -6053
rect 8993 -6241 9051 -6229
rect 9107 -6053 9165 -6041
rect 9107 -6229 9119 -6053
rect 9153 -6229 9165 -6053
rect 9107 -6241 9165 -6229
rect 9365 -6053 9423 -6041
rect 9365 -6229 9377 -6053
rect 9411 -6229 9423 -6053
rect 9365 -6241 9423 -6229
rect 9479 -6053 9537 -6041
rect 9479 -6229 9491 -6053
rect 9525 -6229 9537 -6053
rect 9479 -6241 9537 -6229
rect 9737 -6053 9795 -6041
rect 9737 -6229 9749 -6053
rect 9783 -6229 9795 -6053
rect 9737 -6241 9795 -6229
rect 923 -6471 981 -6459
rect 923 -6647 935 -6471
rect 969 -6647 981 -6471
rect 923 -6659 981 -6647
rect 1181 -6471 1239 -6459
rect 1181 -6647 1193 -6471
rect 1227 -6647 1239 -6471
rect 1181 -6659 1239 -6647
rect 1295 -6471 1353 -6459
rect 1295 -6647 1307 -6471
rect 1341 -6647 1353 -6471
rect 1295 -6659 1353 -6647
rect 1553 -6471 1611 -6459
rect 1553 -6647 1565 -6471
rect 1599 -6647 1611 -6471
rect 1553 -6659 1611 -6647
rect 1667 -6471 1725 -6459
rect 1667 -6647 1679 -6471
rect 1713 -6647 1725 -6471
rect 1667 -6659 1725 -6647
rect 1925 -6471 1983 -6459
rect 1925 -6647 1937 -6471
rect 1971 -6647 1983 -6471
rect 1925 -6659 1983 -6647
rect 2039 -6471 2097 -6459
rect 2039 -6647 2051 -6471
rect 2085 -6647 2097 -6471
rect 2039 -6659 2097 -6647
rect 2297 -6471 2355 -6459
rect 2297 -6647 2309 -6471
rect 2343 -6647 2355 -6471
rect 2297 -6659 2355 -6647
rect 2411 -6471 2469 -6459
rect 2411 -6647 2423 -6471
rect 2457 -6647 2469 -6471
rect 2411 -6659 2469 -6647
rect 2669 -6471 2727 -6459
rect 2669 -6647 2681 -6471
rect 2715 -6647 2727 -6471
rect 2669 -6659 2727 -6647
rect 2783 -6471 2841 -6459
rect 2783 -6647 2795 -6471
rect 2829 -6647 2841 -6471
rect 2783 -6659 2841 -6647
rect 3041 -6471 3099 -6459
rect 3041 -6647 3053 -6471
rect 3087 -6647 3099 -6471
rect 3041 -6659 3099 -6647
rect 3155 -6471 3213 -6459
rect 3155 -6647 3167 -6471
rect 3201 -6647 3213 -6471
rect 3155 -6659 3213 -6647
rect 3413 -6471 3471 -6459
rect 3413 -6647 3425 -6471
rect 3459 -6647 3471 -6471
rect 3413 -6659 3471 -6647
rect 3527 -6471 3585 -6459
rect 3527 -6647 3539 -6471
rect 3573 -6647 3585 -6471
rect 3527 -6659 3585 -6647
rect 3785 -6471 3843 -6459
rect 3785 -6647 3797 -6471
rect 3831 -6647 3843 -6471
rect 3785 -6659 3843 -6647
rect 3899 -6471 3957 -6459
rect 3899 -6647 3911 -6471
rect 3945 -6647 3957 -6471
rect 3899 -6659 3957 -6647
rect 4157 -6471 4215 -6459
rect 4157 -6647 4169 -6471
rect 4203 -6647 4215 -6471
rect 4157 -6659 4215 -6647
rect 4271 -6471 4329 -6459
rect 4271 -6647 4283 -6471
rect 4317 -6647 4329 -6471
rect 4271 -6659 4329 -6647
rect 4529 -6471 4587 -6459
rect 4529 -6647 4541 -6471
rect 4575 -6647 4587 -6471
rect 4529 -6659 4587 -6647
rect 4643 -6471 4701 -6459
rect 4643 -6647 4655 -6471
rect 4689 -6647 4701 -6471
rect 4643 -6659 4701 -6647
rect 4901 -6471 4959 -6459
rect 4901 -6647 4913 -6471
rect 4947 -6647 4959 -6471
rect 4901 -6659 4959 -6647
rect 5015 -6471 5073 -6459
rect 5015 -6647 5027 -6471
rect 5061 -6647 5073 -6471
rect 5015 -6659 5073 -6647
rect 5273 -6471 5331 -6459
rect 5273 -6647 5285 -6471
rect 5319 -6647 5331 -6471
rect 5273 -6659 5331 -6647
rect 5387 -6471 5445 -6459
rect 5387 -6647 5399 -6471
rect 5433 -6647 5445 -6471
rect 5387 -6659 5445 -6647
rect 5645 -6471 5703 -6459
rect 5645 -6647 5657 -6471
rect 5691 -6647 5703 -6471
rect 5645 -6659 5703 -6647
rect 5759 -6471 5817 -6459
rect 5759 -6647 5771 -6471
rect 5805 -6647 5817 -6471
rect 5759 -6659 5817 -6647
rect 6017 -6471 6075 -6459
rect 6017 -6647 6029 -6471
rect 6063 -6647 6075 -6471
rect 6017 -6659 6075 -6647
rect 6131 -6471 6189 -6459
rect 6131 -6647 6143 -6471
rect 6177 -6647 6189 -6471
rect 6131 -6659 6189 -6647
rect 6389 -6471 6447 -6459
rect 6389 -6647 6401 -6471
rect 6435 -6647 6447 -6471
rect 6389 -6659 6447 -6647
rect 6503 -6471 6561 -6459
rect 6503 -6647 6515 -6471
rect 6549 -6647 6561 -6471
rect 6503 -6659 6561 -6647
rect 6761 -6471 6819 -6459
rect 6761 -6647 6773 -6471
rect 6807 -6647 6819 -6471
rect 6761 -6659 6819 -6647
rect 6875 -6471 6933 -6459
rect 6875 -6647 6887 -6471
rect 6921 -6647 6933 -6471
rect 6875 -6659 6933 -6647
rect 7133 -6471 7191 -6459
rect 7133 -6647 7145 -6471
rect 7179 -6647 7191 -6471
rect 7133 -6659 7191 -6647
rect 7247 -6471 7305 -6459
rect 7247 -6647 7259 -6471
rect 7293 -6647 7305 -6471
rect 7247 -6659 7305 -6647
rect 7505 -6471 7563 -6459
rect 7505 -6647 7517 -6471
rect 7551 -6647 7563 -6471
rect 7505 -6659 7563 -6647
rect 7619 -6471 7677 -6459
rect 7619 -6647 7631 -6471
rect 7665 -6647 7677 -6471
rect 7619 -6659 7677 -6647
rect 7877 -6471 7935 -6459
rect 7877 -6647 7889 -6471
rect 7923 -6647 7935 -6471
rect 7877 -6659 7935 -6647
rect 7991 -6471 8049 -6459
rect 7991 -6647 8003 -6471
rect 8037 -6647 8049 -6471
rect 7991 -6659 8049 -6647
rect 8249 -6471 8307 -6459
rect 8249 -6647 8261 -6471
rect 8295 -6647 8307 -6471
rect 8249 -6659 8307 -6647
rect 8363 -6471 8421 -6459
rect 8363 -6647 8375 -6471
rect 8409 -6647 8421 -6471
rect 8363 -6659 8421 -6647
rect 8621 -6471 8679 -6459
rect 8621 -6647 8633 -6471
rect 8667 -6647 8679 -6471
rect 8621 -6659 8679 -6647
rect 8735 -6471 8793 -6459
rect 8735 -6647 8747 -6471
rect 8781 -6647 8793 -6471
rect 8735 -6659 8793 -6647
rect 8993 -6471 9051 -6459
rect 8993 -6647 9005 -6471
rect 9039 -6647 9051 -6471
rect 8993 -6659 9051 -6647
rect 9107 -6471 9165 -6459
rect 9107 -6647 9119 -6471
rect 9153 -6647 9165 -6471
rect 9107 -6659 9165 -6647
rect 9365 -6471 9423 -6459
rect 9365 -6647 9377 -6471
rect 9411 -6647 9423 -6471
rect 9365 -6659 9423 -6647
rect 9479 -6471 9537 -6459
rect 9479 -6647 9491 -6471
rect 9525 -6647 9537 -6471
rect 9479 -6659 9537 -6647
rect 9737 -6471 9795 -6459
rect 9737 -6647 9749 -6471
rect 9783 -6647 9795 -6471
rect 9737 -6659 9795 -6647
rect 923 -6889 981 -6877
rect 923 -7065 935 -6889
rect 969 -7065 981 -6889
rect 923 -7077 981 -7065
rect 1181 -6889 1239 -6877
rect 1181 -7065 1193 -6889
rect 1227 -7065 1239 -6889
rect 1181 -7077 1239 -7065
rect 1295 -6889 1353 -6877
rect 1295 -7065 1307 -6889
rect 1341 -7065 1353 -6889
rect 1295 -7077 1353 -7065
rect 1553 -6889 1611 -6877
rect 1553 -7065 1565 -6889
rect 1599 -7065 1611 -6889
rect 1553 -7077 1611 -7065
rect 1667 -6889 1725 -6877
rect 1667 -7065 1679 -6889
rect 1713 -7065 1725 -6889
rect 1667 -7077 1725 -7065
rect 1925 -6889 1983 -6877
rect 1925 -7065 1937 -6889
rect 1971 -7065 1983 -6889
rect 1925 -7077 1983 -7065
rect 2039 -6889 2097 -6877
rect 2039 -7065 2051 -6889
rect 2085 -7065 2097 -6889
rect 2039 -7077 2097 -7065
rect 2297 -6889 2355 -6877
rect 2297 -7065 2309 -6889
rect 2343 -7065 2355 -6889
rect 2297 -7077 2355 -7065
rect 2411 -6889 2469 -6877
rect 2411 -7065 2423 -6889
rect 2457 -7065 2469 -6889
rect 2411 -7077 2469 -7065
rect 2669 -6889 2727 -6877
rect 2669 -7065 2681 -6889
rect 2715 -7065 2727 -6889
rect 2669 -7077 2727 -7065
rect 2783 -6889 2841 -6877
rect 2783 -7065 2795 -6889
rect 2829 -7065 2841 -6889
rect 2783 -7077 2841 -7065
rect 3041 -6889 3099 -6877
rect 3041 -7065 3053 -6889
rect 3087 -7065 3099 -6889
rect 3041 -7077 3099 -7065
rect 3155 -6889 3213 -6877
rect 3155 -7065 3167 -6889
rect 3201 -7065 3213 -6889
rect 3155 -7077 3213 -7065
rect 3413 -6889 3471 -6877
rect 3413 -7065 3425 -6889
rect 3459 -7065 3471 -6889
rect 3413 -7077 3471 -7065
rect 3527 -6889 3585 -6877
rect 3527 -7065 3539 -6889
rect 3573 -7065 3585 -6889
rect 3527 -7077 3585 -7065
rect 3785 -6889 3843 -6877
rect 3785 -7065 3797 -6889
rect 3831 -7065 3843 -6889
rect 3785 -7077 3843 -7065
rect 3899 -6889 3957 -6877
rect 3899 -7065 3911 -6889
rect 3945 -7065 3957 -6889
rect 3899 -7077 3957 -7065
rect 4157 -6889 4215 -6877
rect 4157 -7065 4169 -6889
rect 4203 -7065 4215 -6889
rect 4157 -7077 4215 -7065
rect 4271 -6889 4329 -6877
rect 4271 -7065 4283 -6889
rect 4317 -7065 4329 -6889
rect 4271 -7077 4329 -7065
rect 4529 -6889 4587 -6877
rect 4529 -7065 4541 -6889
rect 4575 -7065 4587 -6889
rect 4529 -7077 4587 -7065
rect 4643 -6889 4701 -6877
rect 4643 -7065 4655 -6889
rect 4689 -7065 4701 -6889
rect 4643 -7077 4701 -7065
rect 4901 -6889 4959 -6877
rect 4901 -7065 4913 -6889
rect 4947 -7065 4959 -6889
rect 4901 -7077 4959 -7065
rect 5015 -6889 5073 -6877
rect 5015 -7065 5027 -6889
rect 5061 -7065 5073 -6889
rect 5015 -7077 5073 -7065
rect 5273 -6889 5331 -6877
rect 5273 -7065 5285 -6889
rect 5319 -7065 5331 -6889
rect 5273 -7077 5331 -7065
rect 5387 -6889 5445 -6877
rect 5387 -7065 5399 -6889
rect 5433 -7065 5445 -6889
rect 5387 -7077 5445 -7065
rect 5645 -6889 5703 -6877
rect 5645 -7065 5657 -6889
rect 5691 -7065 5703 -6889
rect 5645 -7077 5703 -7065
rect 5759 -6889 5817 -6877
rect 5759 -7065 5771 -6889
rect 5805 -7065 5817 -6889
rect 5759 -7077 5817 -7065
rect 6017 -6889 6075 -6877
rect 6017 -7065 6029 -6889
rect 6063 -7065 6075 -6889
rect 6017 -7077 6075 -7065
rect 6131 -6889 6189 -6877
rect 6131 -7065 6143 -6889
rect 6177 -7065 6189 -6889
rect 6131 -7077 6189 -7065
rect 6389 -6889 6447 -6877
rect 6389 -7065 6401 -6889
rect 6435 -7065 6447 -6889
rect 6389 -7077 6447 -7065
rect 6503 -6889 6561 -6877
rect 6503 -7065 6515 -6889
rect 6549 -7065 6561 -6889
rect 6503 -7077 6561 -7065
rect 6761 -6889 6819 -6877
rect 6761 -7065 6773 -6889
rect 6807 -7065 6819 -6889
rect 6761 -7077 6819 -7065
rect 6875 -6889 6933 -6877
rect 6875 -7065 6887 -6889
rect 6921 -7065 6933 -6889
rect 6875 -7077 6933 -7065
rect 7133 -6889 7191 -6877
rect 7133 -7065 7145 -6889
rect 7179 -7065 7191 -6889
rect 7133 -7077 7191 -7065
rect 7247 -6889 7305 -6877
rect 7247 -7065 7259 -6889
rect 7293 -7065 7305 -6889
rect 7247 -7077 7305 -7065
rect 7505 -6889 7563 -6877
rect 7505 -7065 7517 -6889
rect 7551 -7065 7563 -6889
rect 7505 -7077 7563 -7065
rect 7619 -6889 7677 -6877
rect 7619 -7065 7631 -6889
rect 7665 -7065 7677 -6889
rect 7619 -7077 7677 -7065
rect 7877 -6889 7935 -6877
rect 7877 -7065 7889 -6889
rect 7923 -7065 7935 -6889
rect 7877 -7077 7935 -7065
rect 7991 -6889 8049 -6877
rect 7991 -7065 8003 -6889
rect 8037 -7065 8049 -6889
rect 7991 -7077 8049 -7065
rect 8249 -6889 8307 -6877
rect 8249 -7065 8261 -6889
rect 8295 -7065 8307 -6889
rect 8249 -7077 8307 -7065
rect 8363 -6889 8421 -6877
rect 8363 -7065 8375 -6889
rect 8409 -7065 8421 -6889
rect 8363 -7077 8421 -7065
rect 8621 -6889 8679 -6877
rect 8621 -7065 8633 -6889
rect 8667 -7065 8679 -6889
rect 8621 -7077 8679 -7065
rect 8735 -6889 8793 -6877
rect 8735 -7065 8747 -6889
rect 8781 -7065 8793 -6889
rect 8735 -7077 8793 -7065
rect 8993 -6889 9051 -6877
rect 8993 -7065 9005 -6889
rect 9039 -7065 9051 -6889
rect 8993 -7077 9051 -7065
rect 9107 -6889 9165 -6877
rect 9107 -7065 9119 -6889
rect 9153 -7065 9165 -6889
rect 9107 -7077 9165 -7065
rect 9365 -6889 9423 -6877
rect 9365 -7065 9377 -6889
rect 9411 -7065 9423 -6889
rect 9365 -7077 9423 -7065
rect 9479 -6889 9537 -6877
rect 9479 -7065 9491 -6889
rect 9525 -7065 9537 -6889
rect 9479 -7077 9537 -7065
rect 9737 -6889 9795 -6877
rect 9737 -7065 9749 -6889
rect 9783 -7065 9795 -6889
rect 9737 -7077 9795 -7065
rect 923 -7307 981 -7295
rect 923 -7483 935 -7307
rect 969 -7483 981 -7307
rect 923 -7495 981 -7483
rect 1181 -7307 1239 -7295
rect 1181 -7483 1193 -7307
rect 1227 -7483 1239 -7307
rect 1181 -7495 1239 -7483
rect 1295 -7307 1353 -7295
rect 1295 -7483 1307 -7307
rect 1341 -7483 1353 -7307
rect 1295 -7495 1353 -7483
rect 1553 -7307 1611 -7295
rect 1553 -7483 1565 -7307
rect 1599 -7483 1611 -7307
rect 1553 -7495 1611 -7483
rect 1667 -7307 1725 -7295
rect 1667 -7483 1679 -7307
rect 1713 -7483 1725 -7307
rect 1667 -7495 1725 -7483
rect 1925 -7307 1983 -7295
rect 1925 -7483 1937 -7307
rect 1971 -7483 1983 -7307
rect 1925 -7495 1983 -7483
rect 2039 -7307 2097 -7295
rect 2039 -7483 2051 -7307
rect 2085 -7483 2097 -7307
rect 2039 -7495 2097 -7483
rect 2297 -7307 2355 -7295
rect 2297 -7483 2309 -7307
rect 2343 -7483 2355 -7307
rect 2297 -7495 2355 -7483
rect 2411 -7307 2469 -7295
rect 2411 -7483 2423 -7307
rect 2457 -7483 2469 -7307
rect 2411 -7495 2469 -7483
rect 2669 -7307 2727 -7295
rect 2669 -7483 2681 -7307
rect 2715 -7483 2727 -7307
rect 2669 -7495 2727 -7483
rect 2783 -7307 2841 -7295
rect 2783 -7483 2795 -7307
rect 2829 -7483 2841 -7307
rect 2783 -7495 2841 -7483
rect 3041 -7307 3099 -7295
rect 3041 -7483 3053 -7307
rect 3087 -7483 3099 -7307
rect 3041 -7495 3099 -7483
rect 3155 -7307 3213 -7295
rect 3155 -7483 3167 -7307
rect 3201 -7483 3213 -7307
rect 3155 -7495 3213 -7483
rect 3413 -7307 3471 -7295
rect 3413 -7483 3425 -7307
rect 3459 -7483 3471 -7307
rect 3413 -7495 3471 -7483
rect 3527 -7307 3585 -7295
rect 3527 -7483 3539 -7307
rect 3573 -7483 3585 -7307
rect 3527 -7495 3585 -7483
rect 3785 -7307 3843 -7295
rect 3785 -7483 3797 -7307
rect 3831 -7483 3843 -7307
rect 3785 -7495 3843 -7483
rect 3899 -7307 3957 -7295
rect 3899 -7483 3911 -7307
rect 3945 -7483 3957 -7307
rect 3899 -7495 3957 -7483
rect 4157 -7307 4215 -7295
rect 4157 -7483 4169 -7307
rect 4203 -7483 4215 -7307
rect 4157 -7495 4215 -7483
rect 4271 -7307 4329 -7295
rect 4271 -7483 4283 -7307
rect 4317 -7483 4329 -7307
rect 4271 -7495 4329 -7483
rect 4529 -7307 4587 -7295
rect 4529 -7483 4541 -7307
rect 4575 -7483 4587 -7307
rect 4529 -7495 4587 -7483
rect 4643 -7307 4701 -7295
rect 4643 -7483 4655 -7307
rect 4689 -7483 4701 -7307
rect 4643 -7495 4701 -7483
rect 4901 -7307 4959 -7295
rect 4901 -7483 4913 -7307
rect 4947 -7483 4959 -7307
rect 4901 -7495 4959 -7483
rect 5015 -7307 5073 -7295
rect 5015 -7483 5027 -7307
rect 5061 -7483 5073 -7307
rect 5015 -7495 5073 -7483
rect 5273 -7307 5331 -7295
rect 5273 -7483 5285 -7307
rect 5319 -7483 5331 -7307
rect 5273 -7495 5331 -7483
rect 5387 -7307 5445 -7295
rect 5387 -7483 5399 -7307
rect 5433 -7483 5445 -7307
rect 5387 -7495 5445 -7483
rect 5645 -7307 5703 -7295
rect 5645 -7483 5657 -7307
rect 5691 -7483 5703 -7307
rect 5645 -7495 5703 -7483
rect 5759 -7307 5817 -7295
rect 5759 -7483 5771 -7307
rect 5805 -7483 5817 -7307
rect 5759 -7495 5817 -7483
rect 6017 -7307 6075 -7295
rect 6017 -7483 6029 -7307
rect 6063 -7483 6075 -7307
rect 6017 -7495 6075 -7483
rect 6131 -7307 6189 -7295
rect 6131 -7483 6143 -7307
rect 6177 -7483 6189 -7307
rect 6131 -7495 6189 -7483
rect 6389 -7307 6447 -7295
rect 6389 -7483 6401 -7307
rect 6435 -7483 6447 -7307
rect 6389 -7495 6447 -7483
rect 6503 -7307 6561 -7295
rect 6503 -7483 6515 -7307
rect 6549 -7483 6561 -7307
rect 6503 -7495 6561 -7483
rect 6761 -7307 6819 -7295
rect 6761 -7483 6773 -7307
rect 6807 -7483 6819 -7307
rect 6761 -7495 6819 -7483
rect 6875 -7307 6933 -7295
rect 6875 -7483 6887 -7307
rect 6921 -7483 6933 -7307
rect 6875 -7495 6933 -7483
rect 7133 -7307 7191 -7295
rect 7133 -7483 7145 -7307
rect 7179 -7483 7191 -7307
rect 7133 -7495 7191 -7483
rect 7247 -7307 7305 -7295
rect 7247 -7483 7259 -7307
rect 7293 -7483 7305 -7307
rect 7247 -7495 7305 -7483
rect 7505 -7307 7563 -7295
rect 7505 -7483 7517 -7307
rect 7551 -7483 7563 -7307
rect 7505 -7495 7563 -7483
rect 7619 -7307 7677 -7295
rect 7619 -7483 7631 -7307
rect 7665 -7483 7677 -7307
rect 7619 -7495 7677 -7483
rect 7877 -7307 7935 -7295
rect 7877 -7483 7889 -7307
rect 7923 -7483 7935 -7307
rect 7877 -7495 7935 -7483
rect 7991 -7307 8049 -7295
rect 7991 -7483 8003 -7307
rect 8037 -7483 8049 -7307
rect 7991 -7495 8049 -7483
rect 8249 -7307 8307 -7295
rect 8249 -7483 8261 -7307
rect 8295 -7483 8307 -7307
rect 8249 -7495 8307 -7483
rect 8363 -7307 8421 -7295
rect 8363 -7483 8375 -7307
rect 8409 -7483 8421 -7307
rect 8363 -7495 8421 -7483
rect 8621 -7307 8679 -7295
rect 8621 -7483 8633 -7307
rect 8667 -7483 8679 -7307
rect 8621 -7495 8679 -7483
rect 8735 -7307 8793 -7295
rect 8735 -7483 8747 -7307
rect 8781 -7483 8793 -7307
rect 8735 -7495 8793 -7483
rect 8993 -7307 9051 -7295
rect 8993 -7483 9005 -7307
rect 9039 -7483 9051 -7307
rect 8993 -7495 9051 -7483
rect 9107 -7307 9165 -7295
rect 9107 -7483 9119 -7307
rect 9153 -7483 9165 -7307
rect 9107 -7495 9165 -7483
rect 9365 -7307 9423 -7295
rect 9365 -7483 9377 -7307
rect 9411 -7483 9423 -7307
rect 9365 -7495 9423 -7483
rect 9479 -7307 9537 -7295
rect 9479 -7483 9491 -7307
rect 9525 -7483 9537 -7307
rect 9479 -7495 9537 -7483
rect 9737 -7307 9795 -7295
rect 9737 -7483 9749 -7307
rect 9783 -7483 9795 -7307
rect 9737 -7495 9795 -7483
<< pdiff >>
rect -565 1020 -507 1032
rect -565 644 -553 1020
rect -519 644 -507 1020
rect -565 632 -507 644
rect -307 1020 -249 1032
rect -307 644 -295 1020
rect -261 644 -249 1020
rect -307 632 -249 644
rect -193 1020 -135 1032
rect -193 644 -181 1020
rect -147 644 -135 1020
rect -193 632 -135 644
rect 65 1020 123 1032
rect 65 644 77 1020
rect 111 644 123 1020
rect 65 632 123 644
rect 179 1020 237 1032
rect 179 644 191 1020
rect 225 644 237 1020
rect 179 632 237 644
rect 437 1020 495 1032
rect 437 644 449 1020
rect 483 644 495 1020
rect 437 632 495 644
rect 551 1020 609 1032
rect 551 644 563 1020
rect 597 644 609 1020
rect 551 632 609 644
rect 809 1020 867 1032
rect 809 644 821 1020
rect 855 644 867 1020
rect 809 632 867 644
rect 923 1020 981 1032
rect 923 644 935 1020
rect 969 644 981 1020
rect 923 632 981 644
rect 1181 1020 1239 1032
rect 1181 644 1193 1020
rect 1227 644 1239 1020
rect 1181 632 1239 644
rect 1295 1020 1353 1032
rect 1295 644 1307 1020
rect 1341 644 1353 1020
rect 1295 632 1353 644
rect 1553 1020 1611 1032
rect 1553 644 1565 1020
rect 1599 644 1611 1020
rect 1553 632 1611 644
rect 1667 1020 1725 1032
rect 1667 644 1679 1020
rect 1713 644 1725 1020
rect 1667 632 1725 644
rect 1925 1020 1983 1032
rect 1925 644 1937 1020
rect 1971 644 1983 1020
rect 1925 632 1983 644
rect 2039 1020 2097 1032
rect 2039 644 2051 1020
rect 2085 644 2097 1020
rect 2039 632 2097 644
rect 2297 1020 2355 1032
rect 2297 644 2309 1020
rect 2343 644 2355 1020
rect 2297 632 2355 644
rect 2411 1020 2469 1032
rect 2411 644 2423 1020
rect 2457 644 2469 1020
rect 2411 632 2469 644
rect 2669 1020 2727 1032
rect 2669 644 2681 1020
rect 2715 644 2727 1020
rect 2669 632 2727 644
rect 2783 1020 2841 1032
rect 2783 644 2795 1020
rect 2829 644 2841 1020
rect 2783 632 2841 644
rect 3041 1020 3099 1032
rect 3041 644 3053 1020
rect 3087 644 3099 1020
rect 3041 632 3099 644
rect 3155 1020 3213 1032
rect 3155 644 3167 1020
rect 3201 644 3213 1020
rect 3155 632 3213 644
rect 3413 1020 3471 1032
rect 3413 644 3425 1020
rect 3459 644 3471 1020
rect 3413 632 3471 644
rect 3527 1020 3585 1032
rect 3527 644 3539 1020
rect 3573 644 3585 1020
rect 3527 632 3585 644
rect 3785 1020 3843 1032
rect 3785 644 3797 1020
rect 3831 644 3843 1020
rect 3785 632 3843 644
rect 3899 1020 3957 1032
rect 3899 644 3911 1020
rect 3945 644 3957 1020
rect 3899 632 3957 644
rect 4157 1020 4215 1032
rect 4157 644 4169 1020
rect 4203 644 4215 1020
rect 4157 632 4215 644
rect 4271 1020 4329 1032
rect 4271 644 4283 1020
rect 4317 644 4329 1020
rect 4271 632 4329 644
rect 4529 1020 4587 1032
rect 4529 644 4541 1020
rect 4575 644 4587 1020
rect 4529 632 4587 644
rect 4643 1020 4701 1032
rect 4643 644 4655 1020
rect 4689 644 4701 1020
rect 4643 632 4701 644
rect 4901 1020 4959 1032
rect 4901 644 4913 1020
rect 4947 644 4959 1020
rect 4901 632 4959 644
rect 5015 1020 5073 1032
rect 5015 644 5027 1020
rect 5061 644 5073 1020
rect 5015 632 5073 644
rect 5273 1020 5331 1032
rect 5273 644 5285 1020
rect 5319 644 5331 1020
rect 5273 632 5331 644
rect 5387 1020 5445 1032
rect 5387 644 5399 1020
rect 5433 644 5445 1020
rect 5387 632 5445 644
rect 5645 1020 5703 1032
rect 5645 644 5657 1020
rect 5691 644 5703 1020
rect 5645 632 5703 644
rect 5759 1020 5817 1032
rect 5759 644 5771 1020
rect 5805 644 5817 1020
rect 5759 632 5817 644
rect 6017 1020 6075 1032
rect 6017 644 6029 1020
rect 6063 644 6075 1020
rect 6017 632 6075 644
rect 6131 1020 6189 1032
rect 6131 644 6143 1020
rect 6177 644 6189 1020
rect 6131 632 6189 644
rect 6389 1020 6447 1032
rect 6389 644 6401 1020
rect 6435 644 6447 1020
rect 6389 632 6447 644
rect 6503 1020 6561 1032
rect 6503 644 6515 1020
rect 6549 644 6561 1020
rect 6503 632 6561 644
rect 6761 1020 6819 1032
rect 6761 644 6773 1020
rect 6807 644 6819 1020
rect 6761 632 6819 644
rect 6875 1020 6933 1032
rect 6875 644 6887 1020
rect 6921 644 6933 1020
rect 6875 632 6933 644
rect 7133 1020 7191 1032
rect 7133 644 7145 1020
rect 7179 644 7191 1020
rect 7133 632 7191 644
rect 7247 1020 7305 1032
rect 7247 644 7259 1020
rect 7293 644 7305 1020
rect 7247 632 7305 644
rect 7505 1020 7563 1032
rect 7505 644 7517 1020
rect 7551 644 7563 1020
rect 7505 632 7563 644
rect 7619 1020 7677 1032
rect 7619 644 7631 1020
rect 7665 644 7677 1020
rect 7619 632 7677 644
rect 7877 1020 7935 1032
rect 7877 644 7889 1020
rect 7923 644 7935 1020
rect 7877 632 7935 644
rect 7991 1020 8049 1032
rect 7991 644 8003 1020
rect 8037 644 8049 1020
rect 7991 632 8049 644
rect 8249 1020 8307 1032
rect 8249 644 8261 1020
rect 8295 644 8307 1020
rect 8249 632 8307 644
rect 8363 1020 8421 1032
rect 8363 644 8375 1020
rect 8409 644 8421 1020
rect 8363 632 8421 644
rect 8621 1020 8679 1032
rect 8621 644 8633 1020
rect 8667 644 8679 1020
rect 8621 632 8679 644
rect 8735 1020 8793 1032
rect 8735 644 8747 1020
rect 8781 644 8793 1020
rect 8735 632 8793 644
rect 8993 1020 9051 1032
rect 8993 644 9005 1020
rect 9039 644 9051 1020
rect 8993 632 9051 644
rect 9107 1020 9165 1032
rect 9107 644 9119 1020
rect 9153 644 9165 1020
rect 9107 632 9165 644
rect 9365 1020 9423 1032
rect 9365 644 9377 1020
rect 9411 644 9423 1020
rect 9365 632 9423 644
rect 9479 1020 9537 1032
rect 9479 644 9491 1020
rect 9525 644 9537 1020
rect 9479 632 9537 644
rect 9737 1020 9795 1032
rect 9737 644 9749 1020
rect 9783 644 9795 1020
rect 9737 632 9795 644
rect 9851 1020 9909 1032
rect 9851 644 9863 1020
rect 9897 644 9909 1020
rect 9851 632 9909 644
rect 10109 1020 10167 1032
rect 10109 644 10121 1020
rect 10155 644 10167 1020
rect 10109 632 10167 644
rect 10223 1020 10281 1032
rect 10223 644 10235 1020
rect 10269 644 10281 1020
rect 10223 632 10281 644
rect 10481 1020 10539 1032
rect 10481 644 10493 1020
rect 10527 644 10539 1020
rect 10481 632 10539 644
rect 10595 1020 10653 1032
rect 10595 644 10607 1020
rect 10641 644 10653 1020
rect 10595 632 10653 644
rect 10853 1020 10911 1032
rect 10853 644 10865 1020
rect 10899 644 10911 1020
rect 10853 632 10911 644
rect 10967 1020 11025 1032
rect 10967 644 10979 1020
rect 11013 644 11025 1020
rect 10967 632 11025 644
rect 11225 1020 11283 1032
rect 11225 644 11237 1020
rect 11271 644 11283 1020
rect 11225 632 11283 644
rect -565 384 -507 396
rect -565 8 -553 384
rect -519 8 -507 384
rect -565 -4 -507 8
rect -307 384 -249 396
rect -307 8 -295 384
rect -261 8 -249 384
rect -307 -4 -249 8
rect -193 384 -135 396
rect -193 8 -181 384
rect -147 8 -135 384
rect -193 -4 -135 8
rect 65 384 123 396
rect 65 8 77 384
rect 111 8 123 384
rect 65 -4 123 8
rect 179 384 237 396
rect 179 8 191 384
rect 225 8 237 384
rect 179 -4 237 8
rect 437 384 495 396
rect 437 8 449 384
rect 483 8 495 384
rect 437 -4 495 8
rect 551 384 609 396
rect 551 8 563 384
rect 597 8 609 384
rect 551 -4 609 8
rect 809 384 867 396
rect 809 8 821 384
rect 855 8 867 384
rect 809 -4 867 8
rect 923 384 981 396
rect 923 8 935 384
rect 969 8 981 384
rect 923 -4 981 8
rect 1181 384 1239 396
rect 1181 8 1193 384
rect 1227 8 1239 384
rect 1181 -4 1239 8
rect 1295 384 1353 396
rect 1295 8 1307 384
rect 1341 8 1353 384
rect 1295 -4 1353 8
rect 1553 384 1611 396
rect 1553 8 1565 384
rect 1599 8 1611 384
rect 1553 -4 1611 8
rect 1667 384 1725 396
rect 1667 8 1679 384
rect 1713 8 1725 384
rect 1667 -4 1725 8
rect 1925 384 1983 396
rect 1925 8 1937 384
rect 1971 8 1983 384
rect 1925 -4 1983 8
rect 2039 384 2097 396
rect 2039 8 2051 384
rect 2085 8 2097 384
rect 2039 -4 2097 8
rect 2297 384 2355 396
rect 2297 8 2309 384
rect 2343 8 2355 384
rect 2297 -4 2355 8
rect 2411 384 2469 396
rect 2411 8 2423 384
rect 2457 8 2469 384
rect 2411 -4 2469 8
rect 2669 384 2727 396
rect 2669 8 2681 384
rect 2715 8 2727 384
rect 2669 -4 2727 8
rect 2783 384 2841 396
rect 2783 8 2795 384
rect 2829 8 2841 384
rect 2783 -4 2841 8
rect 3041 384 3099 396
rect 3041 8 3053 384
rect 3087 8 3099 384
rect 3041 -4 3099 8
rect 3155 384 3213 396
rect 3155 8 3167 384
rect 3201 8 3213 384
rect 3155 -4 3213 8
rect 3413 384 3471 396
rect 3413 8 3425 384
rect 3459 8 3471 384
rect 3413 -4 3471 8
rect 3527 384 3585 396
rect 3527 8 3539 384
rect 3573 8 3585 384
rect 3527 -4 3585 8
rect 3785 384 3843 396
rect 3785 8 3797 384
rect 3831 8 3843 384
rect 3785 -4 3843 8
rect 3899 384 3957 396
rect 3899 8 3911 384
rect 3945 8 3957 384
rect 3899 -4 3957 8
rect 4157 384 4215 396
rect 4157 8 4169 384
rect 4203 8 4215 384
rect 4157 -4 4215 8
rect 4271 384 4329 396
rect 4271 8 4283 384
rect 4317 8 4329 384
rect 4271 -4 4329 8
rect 4529 384 4587 396
rect 4529 8 4541 384
rect 4575 8 4587 384
rect 4529 -4 4587 8
rect 4643 384 4701 396
rect 4643 8 4655 384
rect 4689 8 4701 384
rect 4643 -4 4701 8
rect 4901 384 4959 396
rect 4901 8 4913 384
rect 4947 8 4959 384
rect 4901 -4 4959 8
rect 5015 384 5073 396
rect 5015 8 5027 384
rect 5061 8 5073 384
rect 5015 -4 5073 8
rect 5273 384 5331 396
rect 5273 8 5285 384
rect 5319 8 5331 384
rect 5273 -4 5331 8
rect 5387 384 5445 396
rect 5387 8 5399 384
rect 5433 8 5445 384
rect 5387 -4 5445 8
rect 5645 384 5703 396
rect 5645 8 5657 384
rect 5691 8 5703 384
rect 5645 -4 5703 8
rect 5759 384 5817 396
rect 5759 8 5771 384
rect 5805 8 5817 384
rect 5759 -4 5817 8
rect 6017 384 6075 396
rect 6017 8 6029 384
rect 6063 8 6075 384
rect 6017 -4 6075 8
rect 6131 384 6189 396
rect 6131 8 6143 384
rect 6177 8 6189 384
rect 6131 -4 6189 8
rect 6389 384 6447 396
rect 6389 8 6401 384
rect 6435 8 6447 384
rect 6389 -4 6447 8
rect 6503 384 6561 396
rect 6503 8 6515 384
rect 6549 8 6561 384
rect 6503 -4 6561 8
rect 6761 384 6819 396
rect 6761 8 6773 384
rect 6807 8 6819 384
rect 6761 -4 6819 8
rect 6875 384 6933 396
rect 6875 8 6887 384
rect 6921 8 6933 384
rect 6875 -4 6933 8
rect 7133 384 7191 396
rect 7133 8 7145 384
rect 7179 8 7191 384
rect 7133 -4 7191 8
rect 7247 384 7305 396
rect 7247 8 7259 384
rect 7293 8 7305 384
rect 7247 -4 7305 8
rect 7505 384 7563 396
rect 7505 8 7517 384
rect 7551 8 7563 384
rect 7505 -4 7563 8
rect 7619 384 7677 396
rect 7619 8 7631 384
rect 7665 8 7677 384
rect 7619 -4 7677 8
rect 7877 384 7935 396
rect 7877 8 7889 384
rect 7923 8 7935 384
rect 7877 -4 7935 8
rect 7991 384 8049 396
rect 7991 8 8003 384
rect 8037 8 8049 384
rect 7991 -4 8049 8
rect 8249 384 8307 396
rect 8249 8 8261 384
rect 8295 8 8307 384
rect 8249 -4 8307 8
rect 8363 384 8421 396
rect 8363 8 8375 384
rect 8409 8 8421 384
rect 8363 -4 8421 8
rect 8621 384 8679 396
rect 8621 8 8633 384
rect 8667 8 8679 384
rect 8621 -4 8679 8
rect 8735 384 8793 396
rect 8735 8 8747 384
rect 8781 8 8793 384
rect 8735 -4 8793 8
rect 8993 384 9051 396
rect 8993 8 9005 384
rect 9039 8 9051 384
rect 8993 -4 9051 8
rect 9107 384 9165 396
rect 9107 8 9119 384
rect 9153 8 9165 384
rect 9107 -4 9165 8
rect 9365 384 9423 396
rect 9365 8 9377 384
rect 9411 8 9423 384
rect 9365 -4 9423 8
rect 9479 384 9537 396
rect 9479 8 9491 384
rect 9525 8 9537 384
rect 9479 -4 9537 8
rect 9737 384 9795 396
rect 9737 8 9749 384
rect 9783 8 9795 384
rect 9737 -4 9795 8
rect 9851 384 9909 396
rect 9851 8 9863 384
rect 9897 8 9909 384
rect 9851 -4 9909 8
rect 10109 384 10167 396
rect 10109 8 10121 384
rect 10155 8 10167 384
rect 10109 -4 10167 8
rect 10223 384 10281 396
rect 10223 8 10235 384
rect 10269 8 10281 384
rect 10223 -4 10281 8
rect 10481 384 10539 396
rect 10481 8 10493 384
rect 10527 8 10539 384
rect 10481 -4 10539 8
rect 10595 384 10653 396
rect 10595 8 10607 384
rect 10641 8 10653 384
rect 10595 -4 10653 8
rect 10853 384 10911 396
rect 10853 8 10865 384
rect 10899 8 10911 384
rect 10853 -4 10911 8
rect 10967 384 11025 396
rect 10967 8 10979 384
rect 11013 8 11025 384
rect 10967 -4 11025 8
rect 11225 384 11283 396
rect 11225 8 11237 384
rect 11271 8 11283 384
rect 11225 -4 11283 8
rect -565 -252 -507 -240
rect -565 -628 -553 -252
rect -519 -628 -507 -252
rect -565 -640 -507 -628
rect -307 -252 -249 -240
rect -307 -628 -295 -252
rect -261 -628 -249 -252
rect -307 -640 -249 -628
rect -193 -252 -135 -240
rect -193 -628 -181 -252
rect -147 -628 -135 -252
rect -193 -640 -135 -628
rect 65 -252 123 -240
rect 65 -628 77 -252
rect 111 -628 123 -252
rect 65 -640 123 -628
rect 179 -252 237 -240
rect 179 -628 191 -252
rect 225 -628 237 -252
rect 179 -640 237 -628
rect 437 -252 495 -240
rect 437 -628 449 -252
rect 483 -628 495 -252
rect 437 -640 495 -628
rect 551 -252 609 -240
rect 551 -628 563 -252
rect 597 -628 609 -252
rect 551 -640 609 -628
rect 809 -252 867 -240
rect 809 -628 821 -252
rect 855 -628 867 -252
rect 809 -640 867 -628
rect 923 -252 981 -240
rect 923 -628 935 -252
rect 969 -628 981 -252
rect 923 -640 981 -628
rect 1181 -252 1239 -240
rect 1181 -628 1193 -252
rect 1227 -628 1239 -252
rect 1181 -640 1239 -628
rect 1295 -252 1353 -240
rect 1295 -628 1307 -252
rect 1341 -628 1353 -252
rect 1295 -640 1353 -628
rect 1553 -252 1611 -240
rect 1553 -628 1565 -252
rect 1599 -628 1611 -252
rect 1553 -640 1611 -628
rect 1667 -252 1725 -240
rect 1667 -628 1679 -252
rect 1713 -628 1725 -252
rect 1667 -640 1725 -628
rect 1925 -252 1983 -240
rect 1925 -628 1937 -252
rect 1971 -628 1983 -252
rect 1925 -640 1983 -628
rect 2039 -252 2097 -240
rect 2039 -628 2051 -252
rect 2085 -628 2097 -252
rect 2039 -640 2097 -628
rect 2297 -252 2355 -240
rect 2297 -628 2309 -252
rect 2343 -628 2355 -252
rect 2297 -640 2355 -628
rect 2411 -252 2469 -240
rect 2411 -628 2423 -252
rect 2457 -628 2469 -252
rect 2411 -640 2469 -628
rect 2669 -252 2727 -240
rect 2669 -628 2681 -252
rect 2715 -628 2727 -252
rect 2669 -640 2727 -628
rect 2783 -252 2841 -240
rect 2783 -628 2795 -252
rect 2829 -628 2841 -252
rect 2783 -640 2841 -628
rect 3041 -252 3099 -240
rect 3041 -628 3053 -252
rect 3087 -628 3099 -252
rect 3041 -640 3099 -628
rect 3155 -252 3213 -240
rect 3155 -628 3167 -252
rect 3201 -628 3213 -252
rect 3155 -640 3213 -628
rect 3413 -252 3471 -240
rect 3413 -628 3425 -252
rect 3459 -628 3471 -252
rect 3413 -640 3471 -628
rect 3527 -252 3585 -240
rect 3527 -628 3539 -252
rect 3573 -628 3585 -252
rect 3527 -640 3585 -628
rect 3785 -252 3843 -240
rect 3785 -628 3797 -252
rect 3831 -628 3843 -252
rect 3785 -640 3843 -628
rect 3899 -252 3957 -240
rect 3899 -628 3911 -252
rect 3945 -628 3957 -252
rect 3899 -640 3957 -628
rect 4157 -252 4215 -240
rect 4157 -628 4169 -252
rect 4203 -628 4215 -252
rect 4157 -640 4215 -628
rect 4271 -252 4329 -240
rect 4271 -628 4283 -252
rect 4317 -628 4329 -252
rect 4271 -640 4329 -628
rect 4529 -252 4587 -240
rect 4529 -628 4541 -252
rect 4575 -628 4587 -252
rect 4529 -640 4587 -628
rect 4643 -252 4701 -240
rect 4643 -628 4655 -252
rect 4689 -628 4701 -252
rect 4643 -640 4701 -628
rect 4901 -252 4959 -240
rect 4901 -628 4913 -252
rect 4947 -628 4959 -252
rect 4901 -640 4959 -628
rect 5015 -252 5073 -240
rect 5015 -628 5027 -252
rect 5061 -628 5073 -252
rect 5015 -640 5073 -628
rect 5273 -252 5331 -240
rect 5273 -628 5285 -252
rect 5319 -628 5331 -252
rect 5273 -640 5331 -628
rect 5387 -252 5445 -240
rect 5387 -628 5399 -252
rect 5433 -628 5445 -252
rect 5387 -640 5445 -628
rect 5645 -252 5703 -240
rect 5645 -628 5657 -252
rect 5691 -628 5703 -252
rect 5645 -640 5703 -628
rect 5759 -252 5817 -240
rect 5759 -628 5771 -252
rect 5805 -628 5817 -252
rect 5759 -640 5817 -628
rect 6017 -252 6075 -240
rect 6017 -628 6029 -252
rect 6063 -628 6075 -252
rect 6017 -640 6075 -628
rect 6131 -252 6189 -240
rect 6131 -628 6143 -252
rect 6177 -628 6189 -252
rect 6131 -640 6189 -628
rect 6389 -252 6447 -240
rect 6389 -628 6401 -252
rect 6435 -628 6447 -252
rect 6389 -640 6447 -628
rect 6503 -252 6561 -240
rect 6503 -628 6515 -252
rect 6549 -628 6561 -252
rect 6503 -640 6561 -628
rect 6761 -252 6819 -240
rect 6761 -628 6773 -252
rect 6807 -628 6819 -252
rect 6761 -640 6819 -628
rect 6875 -252 6933 -240
rect 6875 -628 6887 -252
rect 6921 -628 6933 -252
rect 6875 -640 6933 -628
rect 7133 -252 7191 -240
rect 7133 -628 7145 -252
rect 7179 -628 7191 -252
rect 7133 -640 7191 -628
rect 7247 -252 7305 -240
rect 7247 -628 7259 -252
rect 7293 -628 7305 -252
rect 7247 -640 7305 -628
rect 7505 -252 7563 -240
rect 7505 -628 7517 -252
rect 7551 -628 7563 -252
rect 7505 -640 7563 -628
rect 7619 -252 7677 -240
rect 7619 -628 7631 -252
rect 7665 -628 7677 -252
rect 7619 -640 7677 -628
rect 7877 -252 7935 -240
rect 7877 -628 7889 -252
rect 7923 -628 7935 -252
rect 7877 -640 7935 -628
rect 7991 -252 8049 -240
rect 7991 -628 8003 -252
rect 8037 -628 8049 -252
rect 7991 -640 8049 -628
rect 8249 -252 8307 -240
rect 8249 -628 8261 -252
rect 8295 -628 8307 -252
rect 8249 -640 8307 -628
rect 8363 -252 8421 -240
rect 8363 -628 8375 -252
rect 8409 -628 8421 -252
rect 8363 -640 8421 -628
rect 8621 -252 8679 -240
rect 8621 -628 8633 -252
rect 8667 -628 8679 -252
rect 8621 -640 8679 -628
rect 8735 -252 8793 -240
rect 8735 -628 8747 -252
rect 8781 -628 8793 -252
rect 8735 -640 8793 -628
rect 8993 -252 9051 -240
rect 8993 -628 9005 -252
rect 9039 -628 9051 -252
rect 8993 -640 9051 -628
rect 9107 -252 9165 -240
rect 9107 -628 9119 -252
rect 9153 -628 9165 -252
rect 9107 -640 9165 -628
rect 9365 -252 9423 -240
rect 9365 -628 9377 -252
rect 9411 -628 9423 -252
rect 9365 -640 9423 -628
rect 9479 -252 9537 -240
rect 9479 -628 9491 -252
rect 9525 -628 9537 -252
rect 9479 -640 9537 -628
rect 9737 -252 9795 -240
rect 9737 -628 9749 -252
rect 9783 -628 9795 -252
rect 9737 -640 9795 -628
rect 9851 -252 9909 -240
rect 9851 -628 9863 -252
rect 9897 -628 9909 -252
rect 9851 -640 9909 -628
rect 10109 -252 10167 -240
rect 10109 -628 10121 -252
rect 10155 -628 10167 -252
rect 10109 -640 10167 -628
rect 10223 -252 10281 -240
rect 10223 -628 10235 -252
rect 10269 -628 10281 -252
rect 10223 -640 10281 -628
rect 10481 -252 10539 -240
rect 10481 -628 10493 -252
rect 10527 -628 10539 -252
rect 10481 -640 10539 -628
rect 10595 -252 10653 -240
rect 10595 -628 10607 -252
rect 10641 -628 10653 -252
rect 10595 -640 10653 -628
rect 10853 -252 10911 -240
rect 10853 -628 10865 -252
rect 10899 -628 10911 -252
rect 10853 -640 10911 -628
rect 10967 -252 11025 -240
rect 10967 -628 10979 -252
rect 11013 -628 11025 -252
rect 10967 -640 11025 -628
rect 11225 -252 11283 -240
rect 11225 -628 11237 -252
rect 11271 -628 11283 -252
rect 11225 -640 11283 -628
rect 923 -1368 981 -1356
rect 923 -2144 935 -1368
rect 969 -2144 981 -1368
rect 923 -2156 981 -2144
rect 1181 -1368 1239 -1356
rect 1181 -2144 1193 -1368
rect 1227 -2144 1239 -1368
rect 1181 -2156 1239 -2144
rect 1295 -1368 1353 -1356
rect 1295 -2144 1307 -1368
rect 1341 -2144 1353 -1368
rect 1295 -2156 1353 -2144
rect 1553 -1368 1611 -1356
rect 1553 -2144 1565 -1368
rect 1599 -2144 1611 -1368
rect 1553 -2156 1611 -2144
rect 1667 -1368 1725 -1356
rect 1667 -2144 1679 -1368
rect 1713 -2144 1725 -1368
rect 1667 -2156 1725 -2144
rect 1925 -1368 1983 -1356
rect 1925 -2144 1937 -1368
rect 1971 -2144 1983 -1368
rect 1925 -2156 1983 -2144
rect 2039 -1368 2097 -1356
rect 2039 -2144 2051 -1368
rect 2085 -2144 2097 -1368
rect 2039 -2156 2097 -2144
rect 2297 -1368 2355 -1356
rect 2297 -2144 2309 -1368
rect 2343 -2144 2355 -1368
rect 2297 -2156 2355 -2144
rect 2411 -1368 2469 -1356
rect 2411 -2144 2423 -1368
rect 2457 -2144 2469 -1368
rect 2411 -2156 2469 -2144
rect 2669 -1368 2727 -1356
rect 2669 -2144 2681 -1368
rect 2715 -2144 2727 -1368
rect 2669 -2156 2727 -2144
rect 2783 -1368 2841 -1356
rect 2783 -2144 2795 -1368
rect 2829 -2144 2841 -1368
rect 2783 -2156 2841 -2144
rect 3041 -1368 3099 -1356
rect 3041 -2144 3053 -1368
rect 3087 -2144 3099 -1368
rect 3041 -2156 3099 -2144
rect 3155 -1368 3213 -1356
rect 3155 -2144 3167 -1368
rect 3201 -2144 3213 -1368
rect 3155 -2156 3213 -2144
rect 3413 -1368 3471 -1356
rect 3413 -2144 3425 -1368
rect 3459 -2144 3471 -1368
rect 3413 -2156 3471 -2144
rect 3527 -1368 3585 -1356
rect 3527 -2144 3539 -1368
rect 3573 -2144 3585 -1368
rect 3527 -2156 3585 -2144
rect 3785 -1368 3843 -1356
rect 3785 -2144 3797 -1368
rect 3831 -2144 3843 -1368
rect 3785 -2156 3843 -2144
rect 923 -2404 981 -2392
rect 923 -3180 935 -2404
rect 969 -3180 981 -2404
rect 923 -3192 981 -3180
rect 1181 -2404 1239 -2392
rect 1181 -3180 1193 -2404
rect 1227 -3180 1239 -2404
rect 1181 -3192 1239 -3180
rect 1295 -2404 1353 -2392
rect 1295 -3180 1307 -2404
rect 1341 -3180 1353 -2404
rect 1295 -3192 1353 -3180
rect 1553 -2404 1611 -2392
rect 1553 -3180 1565 -2404
rect 1599 -3180 1611 -2404
rect 1553 -3192 1611 -3180
rect 1667 -2404 1725 -2392
rect 1667 -3180 1679 -2404
rect 1713 -3180 1725 -2404
rect 1667 -3192 1725 -3180
rect 1925 -2404 1983 -2392
rect 1925 -3180 1937 -2404
rect 1971 -3180 1983 -2404
rect 1925 -3192 1983 -3180
rect 2039 -2404 2097 -2392
rect 2039 -3180 2051 -2404
rect 2085 -3180 2097 -2404
rect 2039 -3192 2097 -3180
rect 2297 -2404 2355 -2392
rect 2297 -3180 2309 -2404
rect 2343 -3180 2355 -2404
rect 2297 -3192 2355 -3180
rect 2411 -2404 2469 -2392
rect 2411 -3180 2423 -2404
rect 2457 -3180 2469 -2404
rect 2411 -3192 2469 -3180
rect 2669 -2404 2727 -2392
rect 2669 -3180 2681 -2404
rect 2715 -3180 2727 -2404
rect 2669 -3192 2727 -3180
rect 2783 -2404 2841 -2392
rect 2783 -3180 2795 -2404
rect 2829 -3180 2841 -2404
rect 2783 -3192 2841 -3180
rect 3041 -2404 3099 -2392
rect 3041 -3180 3053 -2404
rect 3087 -3180 3099 -2404
rect 3041 -3192 3099 -3180
rect 3155 -2404 3213 -2392
rect 3155 -3180 3167 -2404
rect 3201 -3180 3213 -2404
rect 3155 -3192 3213 -3180
rect 3413 -2404 3471 -2392
rect 3413 -3180 3425 -2404
rect 3459 -3180 3471 -2404
rect 3413 -3192 3471 -3180
rect 3527 -2404 3585 -2392
rect 3527 -3180 3539 -2404
rect 3573 -3180 3585 -2404
rect 3527 -3192 3585 -3180
rect 3785 -2404 3843 -2392
rect 3785 -3180 3797 -2404
rect 3831 -3180 3843 -2404
rect 3785 -3192 3843 -3180
rect 923 -3440 981 -3428
rect 923 -4216 935 -3440
rect 969 -4216 981 -3440
rect 923 -4228 981 -4216
rect 1181 -3440 1239 -3428
rect 1181 -4216 1193 -3440
rect 1227 -4216 1239 -3440
rect 1181 -4228 1239 -4216
rect 1295 -3440 1353 -3428
rect 1295 -4216 1307 -3440
rect 1341 -4216 1353 -3440
rect 1295 -4228 1353 -4216
rect 1553 -3440 1611 -3428
rect 1553 -4216 1565 -3440
rect 1599 -4216 1611 -3440
rect 1553 -4228 1611 -4216
rect 1667 -3440 1725 -3428
rect 1667 -4216 1679 -3440
rect 1713 -4216 1725 -3440
rect 1667 -4228 1725 -4216
rect 1925 -3440 1983 -3428
rect 1925 -4216 1937 -3440
rect 1971 -4216 1983 -3440
rect 1925 -4228 1983 -4216
rect 2039 -3440 2097 -3428
rect 2039 -4216 2051 -3440
rect 2085 -4216 2097 -3440
rect 2039 -4228 2097 -4216
rect 2297 -3440 2355 -3428
rect 2297 -4216 2309 -3440
rect 2343 -4216 2355 -3440
rect 2297 -4228 2355 -4216
rect 2411 -3440 2469 -3428
rect 2411 -4216 2423 -3440
rect 2457 -4216 2469 -3440
rect 2411 -4228 2469 -4216
rect 2669 -3440 2727 -3428
rect 2669 -4216 2681 -3440
rect 2715 -4216 2727 -3440
rect 2669 -4228 2727 -4216
rect 2783 -3440 2841 -3428
rect 2783 -4216 2795 -3440
rect 2829 -4216 2841 -3440
rect 2783 -4228 2841 -4216
rect 3041 -3440 3099 -3428
rect 3041 -4216 3053 -3440
rect 3087 -4216 3099 -3440
rect 3041 -4228 3099 -4216
rect 3155 -3440 3213 -3428
rect 3155 -4216 3167 -3440
rect 3201 -4216 3213 -3440
rect 3155 -4228 3213 -4216
rect 3413 -3440 3471 -3428
rect 3413 -4216 3425 -3440
rect 3459 -4216 3471 -3440
rect 3413 -4228 3471 -4216
rect 3527 -3440 3585 -3428
rect 3527 -4216 3539 -3440
rect 3573 -4216 3585 -3440
rect 3527 -4228 3585 -4216
rect 3785 -3440 3843 -3428
rect 3785 -4216 3797 -3440
rect 3831 -4216 3843 -3440
rect 3785 -4228 3843 -4216
rect 923 -4476 981 -4464
rect 923 -5252 935 -4476
rect 969 -5252 981 -4476
rect 923 -5264 981 -5252
rect 1181 -4476 1239 -4464
rect 1181 -5252 1193 -4476
rect 1227 -5252 1239 -4476
rect 1181 -5264 1239 -5252
rect 1295 -4476 1353 -4464
rect 1295 -5252 1307 -4476
rect 1341 -5252 1353 -4476
rect 1295 -5264 1353 -5252
rect 1553 -4476 1611 -4464
rect 1553 -5252 1565 -4476
rect 1599 -5252 1611 -4476
rect 1553 -5264 1611 -5252
rect 1667 -4476 1725 -4464
rect 1667 -5252 1679 -4476
rect 1713 -5252 1725 -4476
rect 1667 -5264 1725 -5252
rect 1925 -4476 1983 -4464
rect 1925 -5252 1937 -4476
rect 1971 -5252 1983 -4476
rect 1925 -5264 1983 -5252
rect 2039 -4476 2097 -4464
rect 2039 -5252 2051 -4476
rect 2085 -5252 2097 -4476
rect 2039 -5264 2097 -5252
rect 2297 -4476 2355 -4464
rect 2297 -5252 2309 -4476
rect 2343 -5252 2355 -4476
rect 2297 -5264 2355 -5252
rect 2411 -4476 2469 -4464
rect 2411 -5252 2423 -4476
rect 2457 -5252 2469 -4476
rect 2411 -5264 2469 -5252
rect 2669 -4476 2727 -4464
rect 2669 -5252 2681 -4476
rect 2715 -5252 2727 -4476
rect 2669 -5264 2727 -5252
rect 2783 -4476 2841 -4464
rect 2783 -5252 2795 -4476
rect 2829 -5252 2841 -4476
rect 2783 -5264 2841 -5252
rect 3041 -4476 3099 -4464
rect 3041 -5252 3053 -4476
rect 3087 -5252 3099 -4476
rect 3041 -5264 3099 -5252
rect 3155 -4476 3213 -4464
rect 3155 -5252 3167 -4476
rect 3201 -5252 3213 -4476
rect 3155 -5264 3213 -5252
rect 3413 -4476 3471 -4464
rect 3413 -5252 3425 -4476
rect 3459 -5252 3471 -4476
rect 3413 -5264 3471 -5252
rect 3527 -4476 3585 -4464
rect 3527 -5252 3539 -4476
rect 3573 -5252 3585 -4476
rect 3527 -5264 3585 -5252
rect 3785 -4476 3843 -4464
rect 3785 -5252 3797 -4476
rect 3831 -5252 3843 -4476
rect 3785 -5264 3843 -5252
<< ndiffc >>
rect 935 -6229 969 -6053
rect 1193 -6229 1227 -6053
rect 1307 -6229 1341 -6053
rect 1565 -6229 1599 -6053
rect 1679 -6229 1713 -6053
rect 1937 -6229 1971 -6053
rect 2051 -6229 2085 -6053
rect 2309 -6229 2343 -6053
rect 2423 -6229 2457 -6053
rect 2681 -6229 2715 -6053
rect 2795 -6229 2829 -6053
rect 3053 -6229 3087 -6053
rect 3167 -6229 3201 -6053
rect 3425 -6229 3459 -6053
rect 3539 -6229 3573 -6053
rect 3797 -6229 3831 -6053
rect 3911 -6229 3945 -6053
rect 4169 -6229 4203 -6053
rect 4283 -6229 4317 -6053
rect 4541 -6229 4575 -6053
rect 4655 -6229 4689 -6053
rect 4913 -6229 4947 -6053
rect 5027 -6229 5061 -6053
rect 5285 -6229 5319 -6053
rect 5399 -6229 5433 -6053
rect 5657 -6229 5691 -6053
rect 5771 -6229 5805 -6053
rect 6029 -6229 6063 -6053
rect 6143 -6229 6177 -6053
rect 6401 -6229 6435 -6053
rect 6515 -6229 6549 -6053
rect 6773 -6229 6807 -6053
rect 6887 -6229 6921 -6053
rect 7145 -6229 7179 -6053
rect 7259 -6229 7293 -6053
rect 7517 -6229 7551 -6053
rect 7631 -6229 7665 -6053
rect 7889 -6229 7923 -6053
rect 8003 -6229 8037 -6053
rect 8261 -6229 8295 -6053
rect 8375 -6229 8409 -6053
rect 8633 -6229 8667 -6053
rect 8747 -6229 8781 -6053
rect 9005 -6229 9039 -6053
rect 9119 -6229 9153 -6053
rect 9377 -6229 9411 -6053
rect 9491 -6229 9525 -6053
rect 9749 -6229 9783 -6053
rect 935 -6647 969 -6471
rect 1193 -6647 1227 -6471
rect 1307 -6647 1341 -6471
rect 1565 -6647 1599 -6471
rect 1679 -6647 1713 -6471
rect 1937 -6647 1971 -6471
rect 2051 -6647 2085 -6471
rect 2309 -6647 2343 -6471
rect 2423 -6647 2457 -6471
rect 2681 -6647 2715 -6471
rect 2795 -6647 2829 -6471
rect 3053 -6647 3087 -6471
rect 3167 -6647 3201 -6471
rect 3425 -6647 3459 -6471
rect 3539 -6647 3573 -6471
rect 3797 -6647 3831 -6471
rect 3911 -6647 3945 -6471
rect 4169 -6647 4203 -6471
rect 4283 -6647 4317 -6471
rect 4541 -6647 4575 -6471
rect 4655 -6647 4689 -6471
rect 4913 -6647 4947 -6471
rect 5027 -6647 5061 -6471
rect 5285 -6647 5319 -6471
rect 5399 -6647 5433 -6471
rect 5657 -6647 5691 -6471
rect 5771 -6647 5805 -6471
rect 6029 -6647 6063 -6471
rect 6143 -6647 6177 -6471
rect 6401 -6647 6435 -6471
rect 6515 -6647 6549 -6471
rect 6773 -6647 6807 -6471
rect 6887 -6647 6921 -6471
rect 7145 -6647 7179 -6471
rect 7259 -6647 7293 -6471
rect 7517 -6647 7551 -6471
rect 7631 -6647 7665 -6471
rect 7889 -6647 7923 -6471
rect 8003 -6647 8037 -6471
rect 8261 -6647 8295 -6471
rect 8375 -6647 8409 -6471
rect 8633 -6647 8667 -6471
rect 8747 -6647 8781 -6471
rect 9005 -6647 9039 -6471
rect 9119 -6647 9153 -6471
rect 9377 -6647 9411 -6471
rect 9491 -6647 9525 -6471
rect 9749 -6647 9783 -6471
rect 935 -7065 969 -6889
rect 1193 -7065 1227 -6889
rect 1307 -7065 1341 -6889
rect 1565 -7065 1599 -6889
rect 1679 -7065 1713 -6889
rect 1937 -7065 1971 -6889
rect 2051 -7065 2085 -6889
rect 2309 -7065 2343 -6889
rect 2423 -7065 2457 -6889
rect 2681 -7065 2715 -6889
rect 2795 -7065 2829 -6889
rect 3053 -7065 3087 -6889
rect 3167 -7065 3201 -6889
rect 3425 -7065 3459 -6889
rect 3539 -7065 3573 -6889
rect 3797 -7065 3831 -6889
rect 3911 -7065 3945 -6889
rect 4169 -7065 4203 -6889
rect 4283 -7065 4317 -6889
rect 4541 -7065 4575 -6889
rect 4655 -7065 4689 -6889
rect 4913 -7065 4947 -6889
rect 5027 -7065 5061 -6889
rect 5285 -7065 5319 -6889
rect 5399 -7065 5433 -6889
rect 5657 -7065 5691 -6889
rect 5771 -7065 5805 -6889
rect 6029 -7065 6063 -6889
rect 6143 -7065 6177 -6889
rect 6401 -7065 6435 -6889
rect 6515 -7065 6549 -6889
rect 6773 -7065 6807 -6889
rect 6887 -7065 6921 -6889
rect 7145 -7065 7179 -6889
rect 7259 -7065 7293 -6889
rect 7517 -7065 7551 -6889
rect 7631 -7065 7665 -6889
rect 7889 -7065 7923 -6889
rect 8003 -7065 8037 -6889
rect 8261 -7065 8295 -6889
rect 8375 -7065 8409 -6889
rect 8633 -7065 8667 -6889
rect 8747 -7065 8781 -6889
rect 9005 -7065 9039 -6889
rect 9119 -7065 9153 -6889
rect 9377 -7065 9411 -6889
rect 9491 -7065 9525 -6889
rect 9749 -7065 9783 -6889
rect 935 -7483 969 -7307
rect 1193 -7483 1227 -7307
rect 1307 -7483 1341 -7307
rect 1565 -7483 1599 -7307
rect 1679 -7483 1713 -7307
rect 1937 -7483 1971 -7307
rect 2051 -7483 2085 -7307
rect 2309 -7483 2343 -7307
rect 2423 -7483 2457 -7307
rect 2681 -7483 2715 -7307
rect 2795 -7483 2829 -7307
rect 3053 -7483 3087 -7307
rect 3167 -7483 3201 -7307
rect 3425 -7483 3459 -7307
rect 3539 -7483 3573 -7307
rect 3797 -7483 3831 -7307
rect 3911 -7483 3945 -7307
rect 4169 -7483 4203 -7307
rect 4283 -7483 4317 -7307
rect 4541 -7483 4575 -7307
rect 4655 -7483 4689 -7307
rect 4913 -7483 4947 -7307
rect 5027 -7483 5061 -7307
rect 5285 -7483 5319 -7307
rect 5399 -7483 5433 -7307
rect 5657 -7483 5691 -7307
rect 5771 -7483 5805 -7307
rect 6029 -7483 6063 -7307
rect 6143 -7483 6177 -7307
rect 6401 -7483 6435 -7307
rect 6515 -7483 6549 -7307
rect 6773 -7483 6807 -7307
rect 6887 -7483 6921 -7307
rect 7145 -7483 7179 -7307
rect 7259 -7483 7293 -7307
rect 7517 -7483 7551 -7307
rect 7631 -7483 7665 -7307
rect 7889 -7483 7923 -7307
rect 8003 -7483 8037 -7307
rect 8261 -7483 8295 -7307
rect 8375 -7483 8409 -7307
rect 8633 -7483 8667 -7307
rect 8747 -7483 8781 -7307
rect 9005 -7483 9039 -7307
rect 9119 -7483 9153 -7307
rect 9377 -7483 9411 -7307
rect 9491 -7483 9525 -7307
rect 9749 -7483 9783 -7307
<< pdiffc >>
rect -553 644 -519 1020
rect -295 644 -261 1020
rect -181 644 -147 1020
rect 77 644 111 1020
rect 191 644 225 1020
rect 449 644 483 1020
rect 563 644 597 1020
rect 821 644 855 1020
rect 935 644 969 1020
rect 1193 644 1227 1020
rect 1307 644 1341 1020
rect 1565 644 1599 1020
rect 1679 644 1713 1020
rect 1937 644 1971 1020
rect 2051 644 2085 1020
rect 2309 644 2343 1020
rect 2423 644 2457 1020
rect 2681 644 2715 1020
rect 2795 644 2829 1020
rect 3053 644 3087 1020
rect 3167 644 3201 1020
rect 3425 644 3459 1020
rect 3539 644 3573 1020
rect 3797 644 3831 1020
rect 3911 644 3945 1020
rect 4169 644 4203 1020
rect 4283 644 4317 1020
rect 4541 644 4575 1020
rect 4655 644 4689 1020
rect 4913 644 4947 1020
rect 5027 644 5061 1020
rect 5285 644 5319 1020
rect 5399 644 5433 1020
rect 5657 644 5691 1020
rect 5771 644 5805 1020
rect 6029 644 6063 1020
rect 6143 644 6177 1020
rect 6401 644 6435 1020
rect 6515 644 6549 1020
rect 6773 644 6807 1020
rect 6887 644 6921 1020
rect 7145 644 7179 1020
rect 7259 644 7293 1020
rect 7517 644 7551 1020
rect 7631 644 7665 1020
rect 7889 644 7923 1020
rect 8003 644 8037 1020
rect 8261 644 8295 1020
rect 8375 644 8409 1020
rect 8633 644 8667 1020
rect 8747 644 8781 1020
rect 9005 644 9039 1020
rect 9119 644 9153 1020
rect 9377 644 9411 1020
rect 9491 644 9525 1020
rect 9749 644 9783 1020
rect 9863 644 9897 1020
rect 10121 644 10155 1020
rect 10235 644 10269 1020
rect 10493 644 10527 1020
rect 10607 644 10641 1020
rect 10865 644 10899 1020
rect 10979 644 11013 1020
rect 11237 644 11271 1020
rect -553 8 -519 384
rect -295 8 -261 384
rect -181 8 -147 384
rect 77 8 111 384
rect 191 8 225 384
rect 449 8 483 384
rect 563 8 597 384
rect 821 8 855 384
rect 935 8 969 384
rect 1193 8 1227 384
rect 1307 8 1341 384
rect 1565 8 1599 384
rect 1679 8 1713 384
rect 1937 8 1971 384
rect 2051 8 2085 384
rect 2309 8 2343 384
rect 2423 8 2457 384
rect 2681 8 2715 384
rect 2795 8 2829 384
rect 3053 8 3087 384
rect 3167 8 3201 384
rect 3425 8 3459 384
rect 3539 8 3573 384
rect 3797 8 3831 384
rect 3911 8 3945 384
rect 4169 8 4203 384
rect 4283 8 4317 384
rect 4541 8 4575 384
rect 4655 8 4689 384
rect 4913 8 4947 384
rect 5027 8 5061 384
rect 5285 8 5319 384
rect 5399 8 5433 384
rect 5657 8 5691 384
rect 5771 8 5805 384
rect 6029 8 6063 384
rect 6143 8 6177 384
rect 6401 8 6435 384
rect 6515 8 6549 384
rect 6773 8 6807 384
rect 6887 8 6921 384
rect 7145 8 7179 384
rect 7259 8 7293 384
rect 7517 8 7551 384
rect 7631 8 7665 384
rect 7889 8 7923 384
rect 8003 8 8037 384
rect 8261 8 8295 384
rect 8375 8 8409 384
rect 8633 8 8667 384
rect 8747 8 8781 384
rect 9005 8 9039 384
rect 9119 8 9153 384
rect 9377 8 9411 384
rect 9491 8 9525 384
rect 9749 8 9783 384
rect 9863 8 9897 384
rect 10121 8 10155 384
rect 10235 8 10269 384
rect 10493 8 10527 384
rect 10607 8 10641 384
rect 10865 8 10899 384
rect 10979 8 11013 384
rect 11237 8 11271 384
rect -553 -628 -519 -252
rect -295 -628 -261 -252
rect -181 -628 -147 -252
rect 77 -628 111 -252
rect 191 -628 225 -252
rect 449 -628 483 -252
rect 563 -628 597 -252
rect 821 -628 855 -252
rect 935 -628 969 -252
rect 1193 -628 1227 -252
rect 1307 -628 1341 -252
rect 1565 -628 1599 -252
rect 1679 -628 1713 -252
rect 1937 -628 1971 -252
rect 2051 -628 2085 -252
rect 2309 -628 2343 -252
rect 2423 -628 2457 -252
rect 2681 -628 2715 -252
rect 2795 -628 2829 -252
rect 3053 -628 3087 -252
rect 3167 -628 3201 -252
rect 3425 -628 3459 -252
rect 3539 -628 3573 -252
rect 3797 -628 3831 -252
rect 3911 -628 3945 -252
rect 4169 -628 4203 -252
rect 4283 -628 4317 -252
rect 4541 -628 4575 -252
rect 4655 -628 4689 -252
rect 4913 -628 4947 -252
rect 5027 -628 5061 -252
rect 5285 -628 5319 -252
rect 5399 -628 5433 -252
rect 5657 -628 5691 -252
rect 5771 -628 5805 -252
rect 6029 -628 6063 -252
rect 6143 -628 6177 -252
rect 6401 -628 6435 -252
rect 6515 -628 6549 -252
rect 6773 -628 6807 -252
rect 6887 -628 6921 -252
rect 7145 -628 7179 -252
rect 7259 -628 7293 -252
rect 7517 -628 7551 -252
rect 7631 -628 7665 -252
rect 7889 -628 7923 -252
rect 8003 -628 8037 -252
rect 8261 -628 8295 -252
rect 8375 -628 8409 -252
rect 8633 -628 8667 -252
rect 8747 -628 8781 -252
rect 9005 -628 9039 -252
rect 9119 -628 9153 -252
rect 9377 -628 9411 -252
rect 9491 -628 9525 -252
rect 9749 -628 9783 -252
rect 9863 -628 9897 -252
rect 10121 -628 10155 -252
rect 10235 -628 10269 -252
rect 10493 -628 10527 -252
rect 10607 -628 10641 -252
rect 10865 -628 10899 -252
rect 10979 -628 11013 -252
rect 11237 -628 11271 -252
rect 935 -2144 969 -1368
rect 1193 -2144 1227 -1368
rect 1307 -2144 1341 -1368
rect 1565 -2144 1599 -1368
rect 1679 -2144 1713 -1368
rect 1937 -2144 1971 -1368
rect 2051 -2144 2085 -1368
rect 2309 -2144 2343 -1368
rect 2423 -2144 2457 -1368
rect 2681 -2144 2715 -1368
rect 2795 -2144 2829 -1368
rect 3053 -2144 3087 -1368
rect 3167 -2144 3201 -1368
rect 3425 -2144 3459 -1368
rect 3539 -2144 3573 -1368
rect 3797 -2144 3831 -1368
rect 935 -3180 969 -2404
rect 1193 -3180 1227 -2404
rect 1307 -3180 1341 -2404
rect 1565 -3180 1599 -2404
rect 1679 -3180 1713 -2404
rect 1937 -3180 1971 -2404
rect 2051 -3180 2085 -2404
rect 2309 -3180 2343 -2404
rect 2423 -3180 2457 -2404
rect 2681 -3180 2715 -2404
rect 2795 -3180 2829 -2404
rect 3053 -3180 3087 -2404
rect 3167 -3180 3201 -2404
rect 3425 -3180 3459 -2404
rect 3539 -3180 3573 -2404
rect 3797 -3180 3831 -2404
rect 935 -4216 969 -3440
rect 1193 -4216 1227 -3440
rect 1307 -4216 1341 -3440
rect 1565 -4216 1599 -3440
rect 1679 -4216 1713 -3440
rect 1937 -4216 1971 -3440
rect 2051 -4216 2085 -3440
rect 2309 -4216 2343 -3440
rect 2423 -4216 2457 -3440
rect 2681 -4216 2715 -3440
rect 2795 -4216 2829 -3440
rect 3053 -4216 3087 -3440
rect 3167 -4216 3201 -3440
rect 3425 -4216 3459 -3440
rect 3539 -4216 3573 -3440
rect 3797 -4216 3831 -3440
rect 935 -5252 969 -4476
rect 1193 -5252 1227 -4476
rect 1307 -5252 1341 -4476
rect 1565 -5252 1599 -4476
rect 1679 -5252 1713 -4476
rect 1937 -5252 1971 -4476
rect 2051 -5252 2085 -4476
rect 2309 -5252 2343 -4476
rect 2423 -5252 2457 -4476
rect 2681 -5252 2715 -4476
rect 2795 -5252 2829 -4476
rect 3053 -5252 3087 -4476
rect 3167 -5252 3201 -4476
rect 3425 -5252 3459 -4476
rect 3539 -5252 3573 -4476
rect 3797 -5252 3831 -4476
<< psubdiff >>
rect 5985 -3363 6081 -3329
rect 6219 -3363 6315 -3329
rect 5985 -3425 6019 -3363
rect 6281 -3425 6315 -3363
rect 5985 -4519 6019 -4457
rect 6281 -4519 6315 -4457
rect 5985 -4553 6081 -4519
rect 6219 -4553 6315 -4519
rect 821 -5901 917 -5867
rect 9801 -5901 9897 -5867
rect 821 -5963 855 -5901
rect 9863 -5963 9897 -5901
rect 821 -7635 855 -7573
rect 9863 -7635 9897 -7573
rect 821 -7669 917 -7635
rect 9801 -7669 9897 -7635
<< nsubdiff >>
rect -667 1181 -571 1215
rect 11289 1181 11385 1215
rect -667 1119 -633 1181
rect 11351 1119 11385 1181
rect -667 -789 -633 -727
rect 11351 -789 11385 -727
rect -667 -823 -571 -789
rect 11289 -823 11385 -789
rect 821 -1207 917 -1173
rect 3849 -1207 3945 -1173
rect 821 -1269 855 -1207
rect 3911 -1269 3945 -1207
rect 821 -5413 855 -5351
rect 3911 -5413 3945 -5351
rect 821 -5447 917 -5413
rect 3849 -5447 3945 -5413
<< psubdiffcont >>
rect 6081 -3363 6219 -3329
rect 5985 -4457 6019 -3425
rect 6281 -4457 6315 -3425
rect 6081 -4553 6219 -4519
rect 917 -5901 9801 -5867
rect 821 -7573 855 -5963
rect 9863 -7573 9897 -5963
rect 917 -7669 9801 -7635
<< nsubdiffcont >>
rect -571 1181 11289 1215
rect -667 -727 -633 1119
rect 11351 -727 11385 1119
rect -571 -823 11289 -789
rect 917 -1207 3849 -1173
rect 821 -5351 855 -1269
rect 3911 -5351 3945 -1269
rect 917 -5447 3849 -5413
<< poly >>
rect -507 1113 -307 1129
rect -507 1079 -491 1113
rect -323 1079 -307 1113
rect -507 1032 -307 1079
rect -135 1113 65 1129
rect -135 1079 -119 1113
rect 49 1079 65 1113
rect -135 1032 65 1079
rect 237 1113 437 1129
rect 237 1079 253 1113
rect 421 1079 437 1113
rect 237 1032 437 1079
rect 609 1113 809 1129
rect 609 1079 625 1113
rect 793 1079 809 1113
rect 609 1032 809 1079
rect 981 1113 1181 1129
rect 981 1079 997 1113
rect 1165 1079 1181 1113
rect 981 1032 1181 1079
rect 1353 1113 1553 1129
rect 1353 1079 1369 1113
rect 1537 1079 1553 1113
rect 1353 1032 1553 1079
rect 1725 1113 1925 1129
rect 1725 1079 1741 1113
rect 1909 1079 1925 1113
rect 1725 1032 1925 1079
rect 2097 1113 2297 1129
rect 2097 1079 2113 1113
rect 2281 1079 2297 1113
rect 2097 1032 2297 1079
rect 2469 1113 2669 1129
rect 2469 1079 2485 1113
rect 2653 1079 2669 1113
rect 2469 1032 2669 1079
rect 2841 1113 3041 1129
rect 2841 1079 2857 1113
rect 3025 1079 3041 1113
rect 2841 1032 3041 1079
rect 3213 1113 3413 1129
rect 3213 1079 3229 1113
rect 3397 1079 3413 1113
rect 3213 1032 3413 1079
rect 3585 1113 3785 1129
rect 3585 1079 3601 1113
rect 3769 1079 3785 1113
rect 3585 1032 3785 1079
rect 3957 1113 4157 1129
rect 3957 1079 3973 1113
rect 4141 1079 4157 1113
rect 3957 1032 4157 1079
rect 4329 1113 4529 1129
rect 4329 1079 4345 1113
rect 4513 1079 4529 1113
rect 4329 1032 4529 1079
rect 4701 1113 4901 1129
rect 4701 1079 4717 1113
rect 4885 1079 4901 1113
rect 4701 1032 4901 1079
rect 5073 1113 5273 1129
rect 5073 1079 5089 1113
rect 5257 1079 5273 1113
rect 5073 1032 5273 1079
rect 5445 1113 5645 1129
rect 5445 1079 5461 1113
rect 5629 1079 5645 1113
rect 5445 1032 5645 1079
rect 5817 1113 6017 1129
rect 5817 1079 5833 1113
rect 6001 1079 6017 1113
rect 5817 1032 6017 1079
rect 6189 1113 6389 1129
rect 6189 1079 6205 1113
rect 6373 1079 6389 1113
rect 6189 1032 6389 1079
rect 6561 1113 6761 1129
rect 6561 1079 6577 1113
rect 6745 1079 6761 1113
rect 6561 1032 6761 1079
rect 6933 1113 7133 1129
rect 6933 1079 6949 1113
rect 7117 1079 7133 1113
rect 6933 1032 7133 1079
rect 7305 1113 7505 1129
rect 7305 1079 7321 1113
rect 7489 1079 7505 1113
rect 7305 1032 7505 1079
rect 7677 1113 7877 1129
rect 7677 1079 7693 1113
rect 7861 1079 7877 1113
rect 7677 1032 7877 1079
rect 8049 1113 8249 1129
rect 8049 1079 8065 1113
rect 8233 1079 8249 1113
rect 8049 1032 8249 1079
rect 8421 1113 8621 1129
rect 8421 1079 8437 1113
rect 8605 1079 8621 1113
rect 8421 1032 8621 1079
rect 8793 1113 8993 1129
rect 8793 1079 8809 1113
rect 8977 1079 8993 1113
rect 8793 1032 8993 1079
rect 9165 1113 9365 1129
rect 9165 1079 9181 1113
rect 9349 1079 9365 1113
rect 9165 1032 9365 1079
rect 9537 1113 9737 1129
rect 9537 1079 9553 1113
rect 9721 1079 9737 1113
rect 9537 1032 9737 1079
rect 9909 1113 10109 1129
rect 9909 1079 9925 1113
rect 10093 1079 10109 1113
rect 9909 1032 10109 1079
rect 10281 1113 10481 1129
rect 10281 1079 10297 1113
rect 10465 1079 10481 1113
rect 10281 1032 10481 1079
rect 10653 1113 10853 1129
rect 10653 1079 10669 1113
rect 10837 1079 10853 1113
rect 10653 1032 10853 1079
rect 11025 1113 11225 1129
rect 11025 1079 11041 1113
rect 11209 1079 11225 1113
rect 11025 1032 11225 1079
rect -507 585 -307 632
rect -507 551 -491 585
rect -323 551 -307 585
rect -507 535 -307 551
rect -135 585 65 632
rect -135 551 -119 585
rect 49 551 65 585
rect -135 535 65 551
rect 237 585 437 632
rect 237 551 253 585
rect 421 551 437 585
rect 237 535 437 551
rect 609 585 809 632
rect 609 551 625 585
rect 793 551 809 585
rect 609 535 809 551
rect 981 585 1181 632
rect 981 551 997 585
rect 1165 551 1181 585
rect 981 535 1181 551
rect 1353 585 1553 632
rect 1353 551 1369 585
rect 1537 551 1553 585
rect 1353 535 1553 551
rect 1725 585 1925 632
rect 1725 551 1741 585
rect 1909 551 1925 585
rect 1725 535 1925 551
rect 2097 585 2297 632
rect 2097 551 2113 585
rect 2281 551 2297 585
rect 2097 535 2297 551
rect 2469 585 2669 632
rect 2469 551 2485 585
rect 2653 551 2669 585
rect 2469 535 2669 551
rect 2841 585 3041 632
rect 2841 551 2857 585
rect 3025 551 3041 585
rect 2841 535 3041 551
rect 3213 585 3413 632
rect 3213 551 3229 585
rect 3397 551 3413 585
rect 3213 535 3413 551
rect 3585 585 3785 632
rect 3585 551 3601 585
rect 3769 551 3785 585
rect 3585 535 3785 551
rect 3957 585 4157 632
rect 3957 551 3973 585
rect 4141 551 4157 585
rect 3957 535 4157 551
rect 4329 585 4529 632
rect 4329 551 4345 585
rect 4513 551 4529 585
rect 4329 535 4529 551
rect 4701 585 4901 632
rect 4701 551 4717 585
rect 4885 551 4901 585
rect 4701 535 4901 551
rect 5073 585 5273 632
rect 5073 551 5089 585
rect 5257 551 5273 585
rect 5073 535 5273 551
rect 5445 585 5645 632
rect 5445 551 5461 585
rect 5629 551 5645 585
rect 5445 535 5645 551
rect 5817 585 6017 632
rect 5817 551 5833 585
rect 6001 551 6017 585
rect 5817 535 6017 551
rect 6189 585 6389 632
rect 6189 551 6205 585
rect 6373 551 6389 585
rect 6189 535 6389 551
rect 6561 585 6761 632
rect 6561 551 6577 585
rect 6745 551 6761 585
rect 6561 535 6761 551
rect 6933 585 7133 632
rect 6933 551 6949 585
rect 7117 551 7133 585
rect 6933 535 7133 551
rect 7305 585 7505 632
rect 7305 551 7321 585
rect 7489 551 7505 585
rect 7305 535 7505 551
rect 7677 585 7877 632
rect 7677 551 7693 585
rect 7861 551 7877 585
rect 7677 535 7877 551
rect 8049 585 8249 632
rect 8049 551 8065 585
rect 8233 551 8249 585
rect 8049 535 8249 551
rect 8421 585 8621 632
rect 8421 551 8437 585
rect 8605 551 8621 585
rect 8421 535 8621 551
rect 8793 585 8993 632
rect 8793 551 8809 585
rect 8977 551 8993 585
rect 8793 535 8993 551
rect 9165 585 9365 632
rect 9165 551 9181 585
rect 9349 551 9365 585
rect 9165 535 9365 551
rect 9537 585 9737 632
rect 9537 551 9553 585
rect 9721 551 9737 585
rect 9537 535 9737 551
rect 9909 585 10109 632
rect 9909 551 9925 585
rect 10093 551 10109 585
rect 9909 535 10109 551
rect 10281 585 10481 632
rect 10281 551 10297 585
rect 10465 551 10481 585
rect 10281 535 10481 551
rect 10653 585 10853 632
rect 10653 551 10669 585
rect 10837 551 10853 585
rect 10653 535 10853 551
rect 11025 585 11225 632
rect 11025 551 11041 585
rect 11209 551 11225 585
rect 11025 535 11225 551
rect -507 477 -307 493
rect -507 443 -491 477
rect -323 443 -307 477
rect -507 396 -307 443
rect -135 477 65 493
rect -135 443 -119 477
rect 49 443 65 477
rect -135 396 65 443
rect 237 477 437 493
rect 237 443 253 477
rect 421 443 437 477
rect 237 396 437 443
rect 609 477 809 493
rect 609 443 625 477
rect 793 443 809 477
rect 609 396 809 443
rect 981 477 1181 493
rect 981 443 997 477
rect 1165 443 1181 477
rect 981 396 1181 443
rect 1353 477 1553 493
rect 1353 443 1369 477
rect 1537 443 1553 477
rect 1353 396 1553 443
rect 1725 477 1925 493
rect 1725 443 1741 477
rect 1909 443 1925 477
rect 1725 396 1925 443
rect 2097 477 2297 493
rect 2097 443 2113 477
rect 2281 443 2297 477
rect 2097 396 2297 443
rect 2469 477 2669 493
rect 2469 443 2485 477
rect 2653 443 2669 477
rect 2469 396 2669 443
rect 2841 477 3041 493
rect 2841 443 2857 477
rect 3025 443 3041 477
rect 2841 396 3041 443
rect 3213 477 3413 493
rect 3213 443 3229 477
rect 3397 443 3413 477
rect 3213 396 3413 443
rect 3585 477 3785 493
rect 3585 443 3601 477
rect 3769 443 3785 477
rect 3585 396 3785 443
rect 3957 477 4157 493
rect 3957 443 3973 477
rect 4141 443 4157 477
rect 3957 396 4157 443
rect 4329 477 4529 493
rect 4329 443 4345 477
rect 4513 443 4529 477
rect 4329 396 4529 443
rect 4701 477 4901 493
rect 4701 443 4717 477
rect 4885 443 4901 477
rect 4701 396 4901 443
rect 5073 477 5273 493
rect 5073 443 5089 477
rect 5257 443 5273 477
rect 5073 396 5273 443
rect 5445 477 5645 493
rect 5445 443 5461 477
rect 5629 443 5645 477
rect 5445 396 5645 443
rect 5817 477 6017 493
rect 5817 443 5833 477
rect 6001 443 6017 477
rect 5817 396 6017 443
rect 6189 477 6389 493
rect 6189 443 6205 477
rect 6373 443 6389 477
rect 6189 396 6389 443
rect 6561 477 6761 493
rect 6561 443 6577 477
rect 6745 443 6761 477
rect 6561 396 6761 443
rect 6933 477 7133 493
rect 6933 443 6949 477
rect 7117 443 7133 477
rect 6933 396 7133 443
rect 7305 477 7505 493
rect 7305 443 7321 477
rect 7489 443 7505 477
rect 7305 396 7505 443
rect 7677 477 7877 493
rect 7677 443 7693 477
rect 7861 443 7877 477
rect 7677 396 7877 443
rect 8049 477 8249 493
rect 8049 443 8065 477
rect 8233 443 8249 477
rect 8049 396 8249 443
rect 8421 477 8621 493
rect 8421 443 8437 477
rect 8605 443 8621 477
rect 8421 396 8621 443
rect 8793 477 8993 493
rect 8793 443 8809 477
rect 8977 443 8993 477
rect 8793 396 8993 443
rect 9165 477 9365 493
rect 9165 443 9181 477
rect 9349 443 9365 477
rect 9165 396 9365 443
rect 9537 477 9737 493
rect 9537 443 9553 477
rect 9721 443 9737 477
rect 9537 396 9737 443
rect 9909 477 10109 493
rect 9909 443 9925 477
rect 10093 443 10109 477
rect 9909 396 10109 443
rect 10281 477 10481 493
rect 10281 443 10297 477
rect 10465 443 10481 477
rect 10281 396 10481 443
rect 10653 477 10853 493
rect 10653 443 10669 477
rect 10837 443 10853 477
rect 10653 396 10853 443
rect 11025 477 11225 493
rect 11025 443 11041 477
rect 11209 443 11225 477
rect 11025 396 11225 443
rect -507 -51 -307 -4
rect -507 -85 -491 -51
rect -323 -85 -307 -51
rect -507 -101 -307 -85
rect -135 -51 65 -4
rect -135 -85 -119 -51
rect 49 -85 65 -51
rect -135 -101 65 -85
rect 237 -51 437 -4
rect 237 -85 253 -51
rect 421 -85 437 -51
rect 237 -101 437 -85
rect 609 -51 809 -4
rect 609 -85 625 -51
rect 793 -85 809 -51
rect 609 -101 809 -85
rect 981 -51 1181 -4
rect 981 -85 997 -51
rect 1165 -85 1181 -51
rect 981 -101 1181 -85
rect 1353 -51 1553 -4
rect 1353 -85 1369 -51
rect 1537 -85 1553 -51
rect 1353 -101 1553 -85
rect 1725 -51 1925 -4
rect 1725 -85 1741 -51
rect 1909 -85 1925 -51
rect 1725 -101 1925 -85
rect 2097 -51 2297 -4
rect 2097 -85 2113 -51
rect 2281 -85 2297 -51
rect 2097 -101 2297 -85
rect 2469 -51 2669 -4
rect 2469 -85 2485 -51
rect 2653 -85 2669 -51
rect 2469 -101 2669 -85
rect 2841 -51 3041 -4
rect 2841 -85 2857 -51
rect 3025 -85 3041 -51
rect 2841 -101 3041 -85
rect 3213 -51 3413 -4
rect 3213 -85 3229 -51
rect 3397 -85 3413 -51
rect 3213 -101 3413 -85
rect 3585 -51 3785 -4
rect 3585 -85 3601 -51
rect 3769 -85 3785 -51
rect 3585 -101 3785 -85
rect 3957 -51 4157 -4
rect 3957 -85 3973 -51
rect 4141 -85 4157 -51
rect 3957 -101 4157 -85
rect 4329 -51 4529 -4
rect 4329 -85 4345 -51
rect 4513 -85 4529 -51
rect 4329 -101 4529 -85
rect 4701 -51 4901 -4
rect 4701 -85 4717 -51
rect 4885 -85 4901 -51
rect 4701 -101 4901 -85
rect 5073 -51 5273 -4
rect 5073 -85 5089 -51
rect 5257 -85 5273 -51
rect 5073 -101 5273 -85
rect 5445 -51 5645 -4
rect 5445 -85 5461 -51
rect 5629 -85 5645 -51
rect 5445 -101 5645 -85
rect 5817 -51 6017 -4
rect 5817 -85 5833 -51
rect 6001 -85 6017 -51
rect 5817 -101 6017 -85
rect 6189 -51 6389 -4
rect 6189 -85 6205 -51
rect 6373 -85 6389 -51
rect 6189 -101 6389 -85
rect 6561 -51 6761 -4
rect 6561 -85 6577 -51
rect 6745 -85 6761 -51
rect 6561 -101 6761 -85
rect 6933 -51 7133 -4
rect 6933 -85 6949 -51
rect 7117 -85 7133 -51
rect 6933 -101 7133 -85
rect 7305 -51 7505 -4
rect 7305 -85 7321 -51
rect 7489 -85 7505 -51
rect 7305 -101 7505 -85
rect 7677 -51 7877 -4
rect 7677 -85 7693 -51
rect 7861 -85 7877 -51
rect 7677 -101 7877 -85
rect 8049 -51 8249 -4
rect 8049 -85 8065 -51
rect 8233 -85 8249 -51
rect 8049 -101 8249 -85
rect 8421 -51 8621 -4
rect 8421 -85 8437 -51
rect 8605 -85 8621 -51
rect 8421 -101 8621 -85
rect 8793 -51 8993 -4
rect 8793 -85 8809 -51
rect 8977 -85 8993 -51
rect 8793 -101 8993 -85
rect 9165 -51 9365 -4
rect 9165 -85 9181 -51
rect 9349 -85 9365 -51
rect 9165 -101 9365 -85
rect 9537 -51 9737 -4
rect 9537 -85 9553 -51
rect 9721 -85 9737 -51
rect 9537 -101 9737 -85
rect 9909 -51 10109 -4
rect 9909 -85 9925 -51
rect 10093 -85 10109 -51
rect 9909 -101 10109 -85
rect 10281 -51 10481 -4
rect 10281 -85 10297 -51
rect 10465 -85 10481 -51
rect 10281 -101 10481 -85
rect 10653 -51 10853 -4
rect 10653 -85 10669 -51
rect 10837 -85 10853 -51
rect 10653 -101 10853 -85
rect 11025 -51 11225 -4
rect 11025 -85 11041 -51
rect 11209 -85 11225 -51
rect 11025 -101 11225 -85
rect -507 -159 -307 -143
rect -507 -193 -491 -159
rect -323 -193 -307 -159
rect -507 -240 -307 -193
rect -135 -159 65 -143
rect -135 -193 -119 -159
rect 49 -193 65 -159
rect -135 -240 65 -193
rect 237 -159 437 -143
rect 237 -193 253 -159
rect 421 -193 437 -159
rect 237 -240 437 -193
rect 609 -159 809 -143
rect 609 -193 625 -159
rect 793 -193 809 -159
rect 609 -240 809 -193
rect 981 -159 1181 -143
rect 981 -193 997 -159
rect 1165 -193 1181 -159
rect 981 -240 1181 -193
rect 1353 -159 1553 -143
rect 1353 -193 1369 -159
rect 1537 -193 1553 -159
rect 1353 -240 1553 -193
rect 1725 -159 1925 -143
rect 1725 -193 1741 -159
rect 1909 -193 1925 -159
rect 1725 -240 1925 -193
rect 2097 -159 2297 -143
rect 2097 -193 2113 -159
rect 2281 -193 2297 -159
rect 2097 -240 2297 -193
rect 2469 -159 2669 -143
rect 2469 -193 2485 -159
rect 2653 -193 2669 -159
rect 2469 -240 2669 -193
rect 2841 -159 3041 -143
rect 2841 -193 2857 -159
rect 3025 -193 3041 -159
rect 2841 -240 3041 -193
rect 3213 -159 3413 -143
rect 3213 -193 3229 -159
rect 3397 -193 3413 -159
rect 3213 -240 3413 -193
rect 3585 -159 3785 -143
rect 3585 -193 3601 -159
rect 3769 -193 3785 -159
rect 3585 -240 3785 -193
rect 3957 -159 4157 -143
rect 3957 -193 3973 -159
rect 4141 -193 4157 -159
rect 3957 -240 4157 -193
rect 4329 -159 4529 -143
rect 4329 -193 4345 -159
rect 4513 -193 4529 -159
rect 4329 -240 4529 -193
rect 4701 -159 4901 -143
rect 4701 -193 4717 -159
rect 4885 -193 4901 -159
rect 4701 -240 4901 -193
rect 5073 -159 5273 -143
rect 5073 -193 5089 -159
rect 5257 -193 5273 -159
rect 5073 -240 5273 -193
rect 5445 -159 5645 -143
rect 5445 -193 5461 -159
rect 5629 -193 5645 -159
rect 5445 -240 5645 -193
rect 5817 -159 6017 -143
rect 5817 -193 5833 -159
rect 6001 -193 6017 -159
rect 5817 -240 6017 -193
rect 6189 -159 6389 -143
rect 6189 -193 6205 -159
rect 6373 -193 6389 -159
rect 6189 -240 6389 -193
rect 6561 -159 6761 -143
rect 6561 -193 6577 -159
rect 6745 -193 6761 -159
rect 6561 -240 6761 -193
rect 6933 -159 7133 -143
rect 6933 -193 6949 -159
rect 7117 -193 7133 -159
rect 6933 -240 7133 -193
rect 7305 -159 7505 -143
rect 7305 -193 7321 -159
rect 7489 -193 7505 -159
rect 7305 -240 7505 -193
rect 7677 -159 7877 -143
rect 7677 -193 7693 -159
rect 7861 -193 7877 -159
rect 7677 -240 7877 -193
rect 8049 -159 8249 -143
rect 8049 -193 8065 -159
rect 8233 -193 8249 -159
rect 8049 -240 8249 -193
rect 8421 -159 8621 -143
rect 8421 -193 8437 -159
rect 8605 -193 8621 -159
rect 8421 -240 8621 -193
rect 8793 -159 8993 -143
rect 8793 -193 8809 -159
rect 8977 -193 8993 -159
rect 8793 -240 8993 -193
rect 9165 -159 9365 -143
rect 9165 -193 9181 -159
rect 9349 -193 9365 -159
rect 9165 -240 9365 -193
rect 9537 -159 9737 -143
rect 9537 -193 9553 -159
rect 9721 -193 9737 -159
rect 9537 -240 9737 -193
rect 9909 -159 10109 -143
rect 9909 -193 9925 -159
rect 10093 -193 10109 -159
rect 9909 -240 10109 -193
rect 10281 -159 10481 -143
rect 10281 -193 10297 -159
rect 10465 -193 10481 -159
rect 10281 -240 10481 -193
rect 10653 -159 10853 -143
rect 10653 -193 10669 -159
rect 10837 -193 10853 -159
rect 10653 -240 10853 -193
rect 11025 -159 11225 -143
rect 11025 -193 11041 -159
rect 11209 -193 11225 -159
rect 11025 -240 11225 -193
rect -507 -687 -307 -640
rect -507 -721 -491 -687
rect -323 -721 -307 -687
rect -507 -737 -307 -721
rect -135 -687 65 -640
rect -135 -721 -119 -687
rect 49 -721 65 -687
rect -135 -737 65 -721
rect 237 -687 437 -640
rect 237 -721 253 -687
rect 421 -721 437 -687
rect 237 -737 437 -721
rect 609 -687 809 -640
rect 609 -721 625 -687
rect 793 -721 809 -687
rect 609 -737 809 -721
rect 981 -687 1181 -640
rect 981 -721 997 -687
rect 1165 -721 1181 -687
rect 981 -737 1181 -721
rect 1353 -687 1553 -640
rect 1353 -721 1369 -687
rect 1537 -721 1553 -687
rect 1353 -737 1553 -721
rect 1725 -687 1925 -640
rect 1725 -721 1741 -687
rect 1909 -721 1925 -687
rect 1725 -737 1925 -721
rect 2097 -687 2297 -640
rect 2097 -721 2113 -687
rect 2281 -721 2297 -687
rect 2097 -737 2297 -721
rect 2469 -687 2669 -640
rect 2469 -721 2485 -687
rect 2653 -721 2669 -687
rect 2469 -737 2669 -721
rect 2841 -687 3041 -640
rect 2841 -721 2857 -687
rect 3025 -721 3041 -687
rect 2841 -737 3041 -721
rect 3213 -687 3413 -640
rect 3213 -721 3229 -687
rect 3397 -721 3413 -687
rect 3213 -737 3413 -721
rect 3585 -687 3785 -640
rect 3585 -721 3601 -687
rect 3769 -721 3785 -687
rect 3585 -737 3785 -721
rect 3957 -687 4157 -640
rect 3957 -721 3973 -687
rect 4141 -721 4157 -687
rect 3957 -737 4157 -721
rect 4329 -687 4529 -640
rect 4329 -721 4345 -687
rect 4513 -721 4529 -687
rect 4329 -737 4529 -721
rect 4701 -687 4901 -640
rect 4701 -721 4717 -687
rect 4885 -721 4901 -687
rect 4701 -737 4901 -721
rect 5073 -687 5273 -640
rect 5073 -721 5089 -687
rect 5257 -721 5273 -687
rect 5073 -737 5273 -721
rect 5445 -687 5645 -640
rect 5445 -721 5461 -687
rect 5629 -721 5645 -687
rect 5445 -737 5645 -721
rect 5817 -687 6017 -640
rect 5817 -721 5833 -687
rect 6001 -721 6017 -687
rect 5817 -737 6017 -721
rect 6189 -687 6389 -640
rect 6189 -721 6205 -687
rect 6373 -721 6389 -687
rect 6189 -737 6389 -721
rect 6561 -687 6761 -640
rect 6561 -721 6577 -687
rect 6745 -721 6761 -687
rect 6561 -737 6761 -721
rect 6933 -687 7133 -640
rect 6933 -721 6949 -687
rect 7117 -721 7133 -687
rect 6933 -737 7133 -721
rect 7305 -687 7505 -640
rect 7305 -721 7321 -687
rect 7489 -721 7505 -687
rect 7305 -737 7505 -721
rect 7677 -687 7877 -640
rect 7677 -721 7693 -687
rect 7861 -721 7877 -687
rect 7677 -737 7877 -721
rect 8049 -687 8249 -640
rect 8049 -721 8065 -687
rect 8233 -721 8249 -687
rect 8049 -737 8249 -721
rect 8421 -687 8621 -640
rect 8421 -721 8437 -687
rect 8605 -721 8621 -687
rect 8421 -737 8621 -721
rect 8793 -687 8993 -640
rect 8793 -721 8809 -687
rect 8977 -721 8993 -687
rect 8793 -737 8993 -721
rect 9165 -687 9365 -640
rect 9165 -721 9181 -687
rect 9349 -721 9365 -687
rect 9165 -737 9365 -721
rect 9537 -687 9737 -640
rect 9537 -721 9553 -687
rect 9721 -721 9737 -687
rect 9537 -737 9737 -721
rect 9909 -687 10109 -640
rect 9909 -721 9925 -687
rect 10093 -721 10109 -687
rect 9909 -737 10109 -721
rect 10281 -687 10481 -640
rect 10281 -721 10297 -687
rect 10465 -721 10481 -687
rect 10281 -737 10481 -721
rect 10653 -687 10853 -640
rect 10653 -721 10669 -687
rect 10837 -721 10853 -687
rect 10653 -737 10853 -721
rect 11025 -687 11225 -640
rect 11025 -721 11041 -687
rect 11209 -721 11225 -687
rect 11025 -737 11225 -721
rect 981 -1275 1181 -1259
rect 981 -1309 997 -1275
rect 1165 -1309 1181 -1275
rect 981 -1356 1181 -1309
rect 1353 -1275 1553 -1259
rect 1353 -1309 1369 -1275
rect 1537 -1309 1553 -1275
rect 1353 -1356 1553 -1309
rect 1725 -1275 1925 -1259
rect 1725 -1309 1741 -1275
rect 1909 -1309 1925 -1275
rect 1725 -1356 1925 -1309
rect 2097 -1275 2297 -1259
rect 2097 -1309 2113 -1275
rect 2281 -1309 2297 -1275
rect 2097 -1356 2297 -1309
rect 2469 -1275 2669 -1259
rect 2469 -1309 2485 -1275
rect 2653 -1309 2669 -1275
rect 2469 -1356 2669 -1309
rect 2841 -1275 3041 -1259
rect 2841 -1309 2857 -1275
rect 3025 -1309 3041 -1275
rect 2841 -1356 3041 -1309
rect 3213 -1275 3413 -1259
rect 3213 -1309 3229 -1275
rect 3397 -1309 3413 -1275
rect 3213 -1356 3413 -1309
rect 3585 -1275 3785 -1259
rect 3585 -1309 3601 -1275
rect 3769 -1309 3785 -1275
rect 3585 -1356 3785 -1309
rect 981 -2203 1181 -2156
rect 981 -2237 997 -2203
rect 1165 -2237 1181 -2203
rect 981 -2253 1181 -2237
rect 1353 -2203 1553 -2156
rect 1353 -2237 1369 -2203
rect 1537 -2237 1553 -2203
rect 1353 -2253 1553 -2237
rect 1725 -2203 1925 -2156
rect 1725 -2237 1741 -2203
rect 1909 -2237 1925 -2203
rect 1725 -2253 1925 -2237
rect 2097 -2203 2297 -2156
rect 2097 -2237 2113 -2203
rect 2281 -2237 2297 -2203
rect 2097 -2253 2297 -2237
rect 2469 -2203 2669 -2156
rect 2469 -2237 2485 -2203
rect 2653 -2237 2669 -2203
rect 2469 -2253 2669 -2237
rect 2841 -2203 3041 -2156
rect 2841 -2237 2857 -2203
rect 3025 -2237 3041 -2203
rect 2841 -2253 3041 -2237
rect 3213 -2203 3413 -2156
rect 3213 -2237 3229 -2203
rect 3397 -2237 3413 -2203
rect 3213 -2253 3413 -2237
rect 3585 -2203 3785 -2156
rect 3585 -2237 3601 -2203
rect 3769 -2237 3785 -2203
rect 3585 -2253 3785 -2237
rect 981 -2311 1181 -2295
rect 981 -2345 997 -2311
rect 1165 -2345 1181 -2311
rect 981 -2392 1181 -2345
rect 1353 -2311 1553 -2295
rect 1353 -2345 1369 -2311
rect 1537 -2345 1553 -2311
rect 1353 -2392 1553 -2345
rect 1725 -2311 1925 -2295
rect 1725 -2345 1741 -2311
rect 1909 -2345 1925 -2311
rect 1725 -2392 1925 -2345
rect 2097 -2311 2297 -2295
rect 2097 -2345 2113 -2311
rect 2281 -2345 2297 -2311
rect 2097 -2392 2297 -2345
rect 2469 -2311 2669 -2295
rect 2469 -2345 2485 -2311
rect 2653 -2345 2669 -2311
rect 2469 -2392 2669 -2345
rect 2841 -2311 3041 -2295
rect 2841 -2345 2857 -2311
rect 3025 -2345 3041 -2311
rect 2841 -2392 3041 -2345
rect 3213 -2311 3413 -2295
rect 3213 -2345 3229 -2311
rect 3397 -2345 3413 -2311
rect 3213 -2392 3413 -2345
rect 3585 -2311 3785 -2295
rect 3585 -2345 3601 -2311
rect 3769 -2345 3785 -2311
rect 3585 -2392 3785 -2345
rect 981 -3239 1181 -3192
rect 981 -3273 997 -3239
rect 1165 -3273 1181 -3239
rect 981 -3289 1181 -3273
rect 1353 -3239 1553 -3192
rect 1353 -3273 1369 -3239
rect 1537 -3273 1553 -3239
rect 1353 -3289 1553 -3273
rect 1725 -3239 1925 -3192
rect 1725 -3273 1741 -3239
rect 1909 -3273 1925 -3239
rect 1725 -3289 1925 -3273
rect 2097 -3239 2297 -3192
rect 2097 -3273 2113 -3239
rect 2281 -3273 2297 -3239
rect 2097 -3289 2297 -3273
rect 2469 -3239 2669 -3192
rect 2469 -3273 2485 -3239
rect 2653 -3273 2669 -3239
rect 2469 -3289 2669 -3273
rect 2841 -3239 3041 -3192
rect 2841 -3273 2857 -3239
rect 3025 -3273 3041 -3239
rect 2841 -3289 3041 -3273
rect 3213 -3239 3413 -3192
rect 3213 -3273 3229 -3239
rect 3397 -3273 3413 -3239
rect 3213 -3289 3413 -3273
rect 3585 -3239 3785 -3192
rect 3585 -3273 3601 -3239
rect 3769 -3273 3785 -3239
rect 3585 -3289 3785 -3273
rect 981 -3347 1181 -3331
rect 981 -3381 997 -3347
rect 1165 -3381 1181 -3347
rect 981 -3428 1181 -3381
rect 1353 -3347 1553 -3331
rect 1353 -3381 1369 -3347
rect 1537 -3381 1553 -3347
rect 1353 -3428 1553 -3381
rect 1725 -3347 1925 -3331
rect 1725 -3381 1741 -3347
rect 1909 -3381 1925 -3347
rect 1725 -3428 1925 -3381
rect 2097 -3347 2297 -3331
rect 2097 -3381 2113 -3347
rect 2281 -3381 2297 -3347
rect 2097 -3428 2297 -3381
rect 2469 -3347 2669 -3331
rect 2469 -3381 2485 -3347
rect 2653 -3381 2669 -3347
rect 2469 -3428 2669 -3381
rect 2841 -3347 3041 -3331
rect 2841 -3381 2857 -3347
rect 3025 -3381 3041 -3347
rect 2841 -3428 3041 -3381
rect 3213 -3347 3413 -3331
rect 3213 -3381 3229 -3347
rect 3397 -3381 3413 -3347
rect 3213 -3428 3413 -3381
rect 3585 -3347 3785 -3331
rect 3585 -3381 3601 -3347
rect 3769 -3381 3785 -3347
rect 3585 -3428 3785 -3381
rect 981 -4275 1181 -4228
rect 981 -4309 997 -4275
rect 1165 -4309 1181 -4275
rect 981 -4325 1181 -4309
rect 1353 -4275 1553 -4228
rect 1353 -4309 1369 -4275
rect 1537 -4309 1553 -4275
rect 1353 -4325 1553 -4309
rect 1725 -4275 1925 -4228
rect 1725 -4309 1741 -4275
rect 1909 -4309 1925 -4275
rect 1725 -4325 1925 -4309
rect 2097 -4275 2297 -4228
rect 2097 -4309 2113 -4275
rect 2281 -4309 2297 -4275
rect 2097 -4325 2297 -4309
rect 2469 -4275 2669 -4228
rect 2469 -4309 2485 -4275
rect 2653 -4309 2669 -4275
rect 2469 -4325 2669 -4309
rect 2841 -4275 3041 -4228
rect 2841 -4309 2857 -4275
rect 3025 -4309 3041 -4275
rect 2841 -4325 3041 -4309
rect 3213 -4275 3413 -4228
rect 3213 -4309 3229 -4275
rect 3397 -4309 3413 -4275
rect 3213 -4325 3413 -4309
rect 3585 -4275 3785 -4228
rect 3585 -4309 3601 -4275
rect 3769 -4309 3785 -4275
rect 3585 -4325 3785 -4309
rect 981 -4383 1181 -4367
rect 981 -4417 997 -4383
rect 1165 -4417 1181 -4383
rect 981 -4464 1181 -4417
rect 1353 -4383 1553 -4367
rect 1353 -4417 1369 -4383
rect 1537 -4417 1553 -4383
rect 1353 -4464 1553 -4417
rect 1725 -4383 1925 -4367
rect 1725 -4417 1741 -4383
rect 1909 -4417 1925 -4383
rect 1725 -4464 1925 -4417
rect 2097 -4383 2297 -4367
rect 2097 -4417 2113 -4383
rect 2281 -4417 2297 -4383
rect 2097 -4464 2297 -4417
rect 2469 -4383 2669 -4367
rect 2469 -4417 2485 -4383
rect 2653 -4417 2669 -4383
rect 2469 -4464 2669 -4417
rect 2841 -4383 3041 -4367
rect 2841 -4417 2857 -4383
rect 3025 -4417 3041 -4383
rect 2841 -4464 3041 -4417
rect 3213 -4383 3413 -4367
rect 3213 -4417 3229 -4383
rect 3397 -4417 3413 -4383
rect 3213 -4464 3413 -4417
rect 3585 -4383 3785 -4367
rect 3585 -4417 3601 -4383
rect 3769 -4417 3785 -4383
rect 3585 -4464 3785 -4417
rect 981 -5311 1181 -5264
rect 981 -5345 997 -5311
rect 1165 -5345 1181 -5311
rect 981 -5361 1181 -5345
rect 1353 -5311 1553 -5264
rect 1353 -5345 1369 -5311
rect 1537 -5345 1553 -5311
rect 1353 -5361 1553 -5345
rect 1725 -5311 1925 -5264
rect 1725 -5345 1741 -5311
rect 1909 -5345 1925 -5311
rect 1725 -5361 1925 -5345
rect 2097 -5311 2297 -5264
rect 2097 -5345 2113 -5311
rect 2281 -5345 2297 -5311
rect 2097 -5361 2297 -5345
rect 2469 -5311 2669 -5264
rect 2469 -5345 2485 -5311
rect 2653 -5345 2669 -5311
rect 2469 -5361 2669 -5345
rect 2841 -5311 3041 -5264
rect 2841 -5345 2857 -5311
rect 3025 -5345 3041 -5311
rect 2841 -5361 3041 -5345
rect 3213 -5311 3413 -5264
rect 3213 -5345 3229 -5311
rect 3397 -5345 3413 -5311
rect 3213 -5361 3413 -5345
rect 3585 -5311 3785 -5264
rect 3585 -5345 3601 -5311
rect 3769 -5345 3785 -5311
rect 3585 -5361 3785 -5345
rect 981 -5969 1181 -5953
rect 981 -6003 997 -5969
rect 1165 -6003 1181 -5969
rect 981 -6041 1181 -6003
rect 1353 -5969 1553 -5953
rect 1353 -6003 1369 -5969
rect 1537 -6003 1553 -5969
rect 1353 -6041 1553 -6003
rect 1725 -5969 1925 -5953
rect 1725 -6003 1741 -5969
rect 1909 -6003 1925 -5969
rect 1725 -6041 1925 -6003
rect 2097 -5969 2297 -5953
rect 2097 -6003 2113 -5969
rect 2281 -6003 2297 -5969
rect 2097 -6041 2297 -6003
rect 2469 -5969 2669 -5953
rect 2469 -6003 2485 -5969
rect 2653 -6003 2669 -5969
rect 2469 -6041 2669 -6003
rect 2841 -5969 3041 -5953
rect 2841 -6003 2857 -5969
rect 3025 -6003 3041 -5969
rect 2841 -6041 3041 -6003
rect 3213 -5969 3413 -5953
rect 3213 -6003 3229 -5969
rect 3397 -6003 3413 -5969
rect 3213 -6041 3413 -6003
rect 3585 -5969 3785 -5953
rect 3585 -6003 3601 -5969
rect 3769 -6003 3785 -5969
rect 3585 -6041 3785 -6003
rect 3957 -5969 4157 -5953
rect 3957 -6003 3973 -5969
rect 4141 -6003 4157 -5969
rect 3957 -6041 4157 -6003
rect 4329 -5969 4529 -5953
rect 4329 -6003 4345 -5969
rect 4513 -6003 4529 -5969
rect 4329 -6041 4529 -6003
rect 4701 -5969 4901 -5953
rect 4701 -6003 4717 -5969
rect 4885 -6003 4901 -5969
rect 4701 -6041 4901 -6003
rect 5073 -5969 5273 -5953
rect 5073 -6003 5089 -5969
rect 5257 -6003 5273 -5969
rect 5073 -6041 5273 -6003
rect 5445 -5969 5645 -5953
rect 5445 -6003 5461 -5969
rect 5629 -6003 5645 -5969
rect 5445 -6041 5645 -6003
rect 5817 -5969 6017 -5953
rect 5817 -6003 5833 -5969
rect 6001 -6003 6017 -5969
rect 5817 -6041 6017 -6003
rect 6189 -5969 6389 -5953
rect 6189 -6003 6205 -5969
rect 6373 -6003 6389 -5969
rect 6189 -6041 6389 -6003
rect 6561 -5969 6761 -5953
rect 6561 -6003 6577 -5969
rect 6745 -6003 6761 -5969
rect 6561 -6041 6761 -6003
rect 6933 -5969 7133 -5953
rect 6933 -6003 6949 -5969
rect 7117 -6003 7133 -5969
rect 6933 -6041 7133 -6003
rect 7305 -5969 7505 -5953
rect 7305 -6003 7321 -5969
rect 7489 -6003 7505 -5969
rect 7305 -6041 7505 -6003
rect 7677 -5969 7877 -5953
rect 7677 -6003 7693 -5969
rect 7861 -6003 7877 -5969
rect 7677 -6041 7877 -6003
rect 8049 -5969 8249 -5953
rect 8049 -6003 8065 -5969
rect 8233 -6003 8249 -5969
rect 8049 -6041 8249 -6003
rect 8421 -5969 8621 -5953
rect 8421 -6003 8437 -5969
rect 8605 -6003 8621 -5969
rect 8421 -6041 8621 -6003
rect 8793 -5969 8993 -5953
rect 8793 -6003 8809 -5969
rect 8977 -6003 8993 -5969
rect 8793 -6041 8993 -6003
rect 9165 -5969 9365 -5953
rect 9165 -6003 9181 -5969
rect 9349 -6003 9365 -5969
rect 9165 -6041 9365 -6003
rect 9537 -5969 9737 -5953
rect 9537 -6003 9553 -5969
rect 9721 -6003 9737 -5969
rect 9537 -6041 9737 -6003
rect 981 -6279 1181 -6241
rect 981 -6313 997 -6279
rect 1165 -6313 1181 -6279
rect 981 -6329 1181 -6313
rect 1353 -6279 1553 -6241
rect 1353 -6313 1369 -6279
rect 1537 -6313 1553 -6279
rect 1353 -6329 1553 -6313
rect 1725 -6279 1925 -6241
rect 1725 -6313 1741 -6279
rect 1909 -6313 1925 -6279
rect 1725 -6329 1925 -6313
rect 2097 -6279 2297 -6241
rect 2097 -6313 2113 -6279
rect 2281 -6313 2297 -6279
rect 2097 -6329 2297 -6313
rect 2469 -6279 2669 -6241
rect 2469 -6313 2485 -6279
rect 2653 -6313 2669 -6279
rect 2469 -6329 2669 -6313
rect 2841 -6279 3041 -6241
rect 2841 -6313 2857 -6279
rect 3025 -6313 3041 -6279
rect 2841 -6329 3041 -6313
rect 3213 -6279 3413 -6241
rect 3213 -6313 3229 -6279
rect 3397 -6313 3413 -6279
rect 3213 -6329 3413 -6313
rect 3585 -6279 3785 -6241
rect 3585 -6313 3601 -6279
rect 3769 -6313 3785 -6279
rect 3585 -6329 3785 -6313
rect 3957 -6279 4157 -6241
rect 3957 -6313 3973 -6279
rect 4141 -6313 4157 -6279
rect 3957 -6329 4157 -6313
rect 4329 -6279 4529 -6241
rect 4329 -6313 4345 -6279
rect 4513 -6313 4529 -6279
rect 4329 -6329 4529 -6313
rect 4701 -6279 4901 -6241
rect 4701 -6313 4717 -6279
rect 4885 -6313 4901 -6279
rect 4701 -6329 4901 -6313
rect 5073 -6279 5273 -6241
rect 5073 -6313 5089 -6279
rect 5257 -6313 5273 -6279
rect 5073 -6329 5273 -6313
rect 5445 -6279 5645 -6241
rect 5445 -6313 5461 -6279
rect 5629 -6313 5645 -6279
rect 5445 -6329 5645 -6313
rect 5817 -6279 6017 -6241
rect 5817 -6313 5833 -6279
rect 6001 -6313 6017 -6279
rect 5817 -6329 6017 -6313
rect 6189 -6279 6389 -6241
rect 6189 -6313 6205 -6279
rect 6373 -6313 6389 -6279
rect 6189 -6329 6389 -6313
rect 6561 -6279 6761 -6241
rect 6561 -6313 6577 -6279
rect 6745 -6313 6761 -6279
rect 6561 -6329 6761 -6313
rect 6933 -6279 7133 -6241
rect 6933 -6313 6949 -6279
rect 7117 -6313 7133 -6279
rect 6933 -6329 7133 -6313
rect 7305 -6279 7505 -6241
rect 7305 -6313 7321 -6279
rect 7489 -6313 7505 -6279
rect 7305 -6329 7505 -6313
rect 7677 -6279 7877 -6241
rect 7677 -6313 7693 -6279
rect 7861 -6313 7877 -6279
rect 7677 -6329 7877 -6313
rect 8049 -6279 8249 -6241
rect 8049 -6313 8065 -6279
rect 8233 -6313 8249 -6279
rect 8049 -6329 8249 -6313
rect 8421 -6279 8621 -6241
rect 8421 -6313 8437 -6279
rect 8605 -6313 8621 -6279
rect 8421 -6329 8621 -6313
rect 8793 -6279 8993 -6241
rect 8793 -6313 8809 -6279
rect 8977 -6313 8993 -6279
rect 8793 -6329 8993 -6313
rect 9165 -6279 9365 -6241
rect 9165 -6313 9181 -6279
rect 9349 -6313 9365 -6279
rect 9165 -6329 9365 -6313
rect 9537 -6279 9737 -6241
rect 9537 -6313 9553 -6279
rect 9721 -6313 9737 -6279
rect 9537 -6329 9737 -6313
rect 981 -6387 1181 -6371
rect 981 -6421 997 -6387
rect 1165 -6421 1181 -6387
rect 981 -6459 1181 -6421
rect 1353 -6387 1553 -6371
rect 1353 -6421 1369 -6387
rect 1537 -6421 1553 -6387
rect 1353 -6459 1553 -6421
rect 1725 -6387 1925 -6371
rect 1725 -6421 1741 -6387
rect 1909 -6421 1925 -6387
rect 1725 -6459 1925 -6421
rect 2097 -6387 2297 -6371
rect 2097 -6421 2113 -6387
rect 2281 -6421 2297 -6387
rect 2097 -6459 2297 -6421
rect 2469 -6387 2669 -6371
rect 2469 -6421 2485 -6387
rect 2653 -6421 2669 -6387
rect 2469 -6459 2669 -6421
rect 2841 -6387 3041 -6371
rect 2841 -6421 2857 -6387
rect 3025 -6421 3041 -6387
rect 2841 -6459 3041 -6421
rect 3213 -6387 3413 -6371
rect 3213 -6421 3229 -6387
rect 3397 -6421 3413 -6387
rect 3213 -6459 3413 -6421
rect 3585 -6387 3785 -6371
rect 3585 -6421 3601 -6387
rect 3769 -6421 3785 -6387
rect 3585 -6459 3785 -6421
rect 3957 -6387 4157 -6371
rect 3957 -6421 3973 -6387
rect 4141 -6421 4157 -6387
rect 3957 -6459 4157 -6421
rect 4329 -6387 4529 -6371
rect 4329 -6421 4345 -6387
rect 4513 -6421 4529 -6387
rect 4329 -6459 4529 -6421
rect 4701 -6387 4901 -6371
rect 4701 -6421 4717 -6387
rect 4885 -6421 4901 -6387
rect 4701 -6459 4901 -6421
rect 5073 -6387 5273 -6371
rect 5073 -6421 5089 -6387
rect 5257 -6421 5273 -6387
rect 5073 -6459 5273 -6421
rect 5445 -6387 5645 -6371
rect 5445 -6421 5461 -6387
rect 5629 -6421 5645 -6387
rect 5445 -6459 5645 -6421
rect 5817 -6387 6017 -6371
rect 5817 -6421 5833 -6387
rect 6001 -6421 6017 -6387
rect 5817 -6459 6017 -6421
rect 6189 -6387 6389 -6371
rect 6189 -6421 6205 -6387
rect 6373 -6421 6389 -6387
rect 6189 -6459 6389 -6421
rect 6561 -6387 6761 -6371
rect 6561 -6421 6577 -6387
rect 6745 -6421 6761 -6387
rect 6561 -6459 6761 -6421
rect 6933 -6387 7133 -6371
rect 6933 -6421 6949 -6387
rect 7117 -6421 7133 -6387
rect 6933 -6459 7133 -6421
rect 7305 -6387 7505 -6371
rect 7305 -6421 7321 -6387
rect 7489 -6421 7505 -6387
rect 7305 -6459 7505 -6421
rect 7677 -6387 7877 -6371
rect 7677 -6421 7693 -6387
rect 7861 -6421 7877 -6387
rect 7677 -6459 7877 -6421
rect 8049 -6387 8249 -6371
rect 8049 -6421 8065 -6387
rect 8233 -6421 8249 -6387
rect 8049 -6459 8249 -6421
rect 8421 -6387 8621 -6371
rect 8421 -6421 8437 -6387
rect 8605 -6421 8621 -6387
rect 8421 -6459 8621 -6421
rect 8793 -6387 8993 -6371
rect 8793 -6421 8809 -6387
rect 8977 -6421 8993 -6387
rect 8793 -6459 8993 -6421
rect 9165 -6387 9365 -6371
rect 9165 -6421 9181 -6387
rect 9349 -6421 9365 -6387
rect 9165 -6459 9365 -6421
rect 9537 -6387 9737 -6371
rect 9537 -6421 9553 -6387
rect 9721 -6421 9737 -6387
rect 9537 -6459 9737 -6421
rect 981 -6697 1181 -6659
rect 981 -6731 997 -6697
rect 1165 -6731 1181 -6697
rect 981 -6747 1181 -6731
rect 1353 -6697 1553 -6659
rect 1353 -6731 1369 -6697
rect 1537 -6731 1553 -6697
rect 1353 -6747 1553 -6731
rect 1725 -6697 1925 -6659
rect 1725 -6731 1741 -6697
rect 1909 -6731 1925 -6697
rect 1725 -6747 1925 -6731
rect 2097 -6697 2297 -6659
rect 2097 -6731 2113 -6697
rect 2281 -6731 2297 -6697
rect 2097 -6747 2297 -6731
rect 2469 -6697 2669 -6659
rect 2469 -6731 2485 -6697
rect 2653 -6731 2669 -6697
rect 2469 -6747 2669 -6731
rect 2841 -6697 3041 -6659
rect 2841 -6731 2857 -6697
rect 3025 -6731 3041 -6697
rect 2841 -6747 3041 -6731
rect 3213 -6697 3413 -6659
rect 3213 -6731 3229 -6697
rect 3397 -6731 3413 -6697
rect 3213 -6747 3413 -6731
rect 3585 -6697 3785 -6659
rect 3585 -6731 3601 -6697
rect 3769 -6731 3785 -6697
rect 3585 -6747 3785 -6731
rect 3957 -6697 4157 -6659
rect 3957 -6731 3973 -6697
rect 4141 -6731 4157 -6697
rect 3957 -6747 4157 -6731
rect 4329 -6697 4529 -6659
rect 4329 -6731 4345 -6697
rect 4513 -6731 4529 -6697
rect 4329 -6747 4529 -6731
rect 4701 -6697 4901 -6659
rect 4701 -6731 4717 -6697
rect 4885 -6731 4901 -6697
rect 4701 -6747 4901 -6731
rect 5073 -6697 5273 -6659
rect 5073 -6731 5089 -6697
rect 5257 -6731 5273 -6697
rect 5073 -6747 5273 -6731
rect 5445 -6697 5645 -6659
rect 5445 -6731 5461 -6697
rect 5629 -6731 5645 -6697
rect 5445 -6747 5645 -6731
rect 5817 -6697 6017 -6659
rect 5817 -6731 5833 -6697
rect 6001 -6731 6017 -6697
rect 5817 -6747 6017 -6731
rect 6189 -6697 6389 -6659
rect 6189 -6731 6205 -6697
rect 6373 -6731 6389 -6697
rect 6189 -6747 6389 -6731
rect 6561 -6697 6761 -6659
rect 6561 -6731 6577 -6697
rect 6745 -6731 6761 -6697
rect 6561 -6747 6761 -6731
rect 6933 -6697 7133 -6659
rect 6933 -6731 6949 -6697
rect 7117 -6731 7133 -6697
rect 6933 -6747 7133 -6731
rect 7305 -6697 7505 -6659
rect 7305 -6731 7321 -6697
rect 7489 -6731 7505 -6697
rect 7305 -6747 7505 -6731
rect 7677 -6697 7877 -6659
rect 7677 -6731 7693 -6697
rect 7861 -6731 7877 -6697
rect 7677 -6747 7877 -6731
rect 8049 -6697 8249 -6659
rect 8049 -6731 8065 -6697
rect 8233 -6731 8249 -6697
rect 8049 -6747 8249 -6731
rect 8421 -6697 8621 -6659
rect 8421 -6731 8437 -6697
rect 8605 -6731 8621 -6697
rect 8421 -6747 8621 -6731
rect 8793 -6697 8993 -6659
rect 8793 -6731 8809 -6697
rect 8977 -6731 8993 -6697
rect 8793 -6747 8993 -6731
rect 9165 -6697 9365 -6659
rect 9165 -6731 9181 -6697
rect 9349 -6731 9365 -6697
rect 9165 -6747 9365 -6731
rect 9537 -6697 9737 -6659
rect 9537 -6731 9553 -6697
rect 9721 -6731 9737 -6697
rect 9537 -6747 9737 -6731
rect 981 -6805 1181 -6789
rect 981 -6839 997 -6805
rect 1165 -6839 1181 -6805
rect 981 -6877 1181 -6839
rect 1353 -6805 1553 -6789
rect 1353 -6839 1369 -6805
rect 1537 -6839 1553 -6805
rect 1353 -6877 1553 -6839
rect 1725 -6805 1925 -6789
rect 1725 -6839 1741 -6805
rect 1909 -6839 1925 -6805
rect 1725 -6877 1925 -6839
rect 2097 -6805 2297 -6789
rect 2097 -6839 2113 -6805
rect 2281 -6839 2297 -6805
rect 2097 -6877 2297 -6839
rect 2469 -6805 2669 -6789
rect 2469 -6839 2485 -6805
rect 2653 -6839 2669 -6805
rect 2469 -6877 2669 -6839
rect 2841 -6805 3041 -6789
rect 2841 -6839 2857 -6805
rect 3025 -6839 3041 -6805
rect 2841 -6877 3041 -6839
rect 3213 -6805 3413 -6789
rect 3213 -6839 3229 -6805
rect 3397 -6839 3413 -6805
rect 3213 -6877 3413 -6839
rect 3585 -6805 3785 -6789
rect 3585 -6839 3601 -6805
rect 3769 -6839 3785 -6805
rect 3585 -6877 3785 -6839
rect 3957 -6805 4157 -6789
rect 3957 -6839 3973 -6805
rect 4141 -6839 4157 -6805
rect 3957 -6877 4157 -6839
rect 4329 -6805 4529 -6789
rect 4329 -6839 4345 -6805
rect 4513 -6839 4529 -6805
rect 4329 -6877 4529 -6839
rect 4701 -6805 4901 -6789
rect 4701 -6839 4717 -6805
rect 4885 -6839 4901 -6805
rect 4701 -6877 4901 -6839
rect 5073 -6805 5273 -6789
rect 5073 -6839 5089 -6805
rect 5257 -6839 5273 -6805
rect 5073 -6877 5273 -6839
rect 5445 -6805 5645 -6789
rect 5445 -6839 5461 -6805
rect 5629 -6839 5645 -6805
rect 5445 -6877 5645 -6839
rect 5817 -6805 6017 -6789
rect 5817 -6839 5833 -6805
rect 6001 -6839 6017 -6805
rect 5817 -6877 6017 -6839
rect 6189 -6805 6389 -6789
rect 6189 -6839 6205 -6805
rect 6373 -6839 6389 -6805
rect 6189 -6877 6389 -6839
rect 6561 -6805 6761 -6789
rect 6561 -6839 6577 -6805
rect 6745 -6839 6761 -6805
rect 6561 -6877 6761 -6839
rect 6933 -6805 7133 -6789
rect 6933 -6839 6949 -6805
rect 7117 -6839 7133 -6805
rect 6933 -6877 7133 -6839
rect 7305 -6805 7505 -6789
rect 7305 -6839 7321 -6805
rect 7489 -6839 7505 -6805
rect 7305 -6877 7505 -6839
rect 7677 -6805 7877 -6789
rect 7677 -6839 7693 -6805
rect 7861 -6839 7877 -6805
rect 7677 -6877 7877 -6839
rect 8049 -6805 8249 -6789
rect 8049 -6839 8065 -6805
rect 8233 -6839 8249 -6805
rect 8049 -6877 8249 -6839
rect 8421 -6805 8621 -6789
rect 8421 -6839 8437 -6805
rect 8605 -6839 8621 -6805
rect 8421 -6877 8621 -6839
rect 8793 -6805 8993 -6789
rect 8793 -6839 8809 -6805
rect 8977 -6839 8993 -6805
rect 8793 -6877 8993 -6839
rect 9165 -6805 9365 -6789
rect 9165 -6839 9181 -6805
rect 9349 -6839 9365 -6805
rect 9165 -6877 9365 -6839
rect 9537 -6805 9737 -6789
rect 9537 -6839 9553 -6805
rect 9721 -6839 9737 -6805
rect 9537 -6877 9737 -6839
rect 981 -7115 1181 -7077
rect 981 -7149 997 -7115
rect 1165 -7149 1181 -7115
rect 981 -7165 1181 -7149
rect 1353 -7115 1553 -7077
rect 1353 -7149 1369 -7115
rect 1537 -7149 1553 -7115
rect 1353 -7165 1553 -7149
rect 1725 -7115 1925 -7077
rect 1725 -7149 1741 -7115
rect 1909 -7149 1925 -7115
rect 1725 -7165 1925 -7149
rect 2097 -7115 2297 -7077
rect 2097 -7149 2113 -7115
rect 2281 -7149 2297 -7115
rect 2097 -7165 2297 -7149
rect 2469 -7115 2669 -7077
rect 2469 -7149 2485 -7115
rect 2653 -7149 2669 -7115
rect 2469 -7165 2669 -7149
rect 2841 -7115 3041 -7077
rect 2841 -7149 2857 -7115
rect 3025 -7149 3041 -7115
rect 2841 -7165 3041 -7149
rect 3213 -7115 3413 -7077
rect 3213 -7149 3229 -7115
rect 3397 -7149 3413 -7115
rect 3213 -7165 3413 -7149
rect 3585 -7115 3785 -7077
rect 3585 -7149 3601 -7115
rect 3769 -7149 3785 -7115
rect 3585 -7165 3785 -7149
rect 3957 -7115 4157 -7077
rect 3957 -7149 3973 -7115
rect 4141 -7149 4157 -7115
rect 3957 -7165 4157 -7149
rect 4329 -7115 4529 -7077
rect 4329 -7149 4345 -7115
rect 4513 -7149 4529 -7115
rect 4329 -7165 4529 -7149
rect 4701 -7115 4901 -7077
rect 4701 -7149 4717 -7115
rect 4885 -7149 4901 -7115
rect 4701 -7165 4901 -7149
rect 5073 -7115 5273 -7077
rect 5073 -7149 5089 -7115
rect 5257 -7149 5273 -7115
rect 5073 -7165 5273 -7149
rect 5445 -7115 5645 -7077
rect 5445 -7149 5461 -7115
rect 5629 -7149 5645 -7115
rect 5445 -7165 5645 -7149
rect 5817 -7115 6017 -7077
rect 5817 -7149 5833 -7115
rect 6001 -7149 6017 -7115
rect 5817 -7165 6017 -7149
rect 6189 -7115 6389 -7077
rect 6189 -7149 6205 -7115
rect 6373 -7149 6389 -7115
rect 6189 -7165 6389 -7149
rect 6561 -7115 6761 -7077
rect 6561 -7149 6577 -7115
rect 6745 -7149 6761 -7115
rect 6561 -7165 6761 -7149
rect 6933 -7115 7133 -7077
rect 6933 -7149 6949 -7115
rect 7117 -7149 7133 -7115
rect 6933 -7165 7133 -7149
rect 7305 -7115 7505 -7077
rect 7305 -7149 7321 -7115
rect 7489 -7149 7505 -7115
rect 7305 -7165 7505 -7149
rect 7677 -7115 7877 -7077
rect 7677 -7149 7693 -7115
rect 7861 -7149 7877 -7115
rect 7677 -7165 7877 -7149
rect 8049 -7115 8249 -7077
rect 8049 -7149 8065 -7115
rect 8233 -7149 8249 -7115
rect 8049 -7165 8249 -7149
rect 8421 -7115 8621 -7077
rect 8421 -7149 8437 -7115
rect 8605 -7149 8621 -7115
rect 8421 -7165 8621 -7149
rect 8793 -7115 8993 -7077
rect 8793 -7149 8809 -7115
rect 8977 -7149 8993 -7115
rect 8793 -7165 8993 -7149
rect 9165 -7115 9365 -7077
rect 9165 -7149 9181 -7115
rect 9349 -7149 9365 -7115
rect 9165 -7165 9365 -7149
rect 9537 -7115 9737 -7077
rect 9537 -7149 9553 -7115
rect 9721 -7149 9737 -7115
rect 9537 -7165 9737 -7149
rect 981 -7223 1181 -7207
rect 981 -7257 997 -7223
rect 1165 -7257 1181 -7223
rect 981 -7295 1181 -7257
rect 1353 -7223 1553 -7207
rect 1353 -7257 1369 -7223
rect 1537 -7257 1553 -7223
rect 1353 -7295 1553 -7257
rect 1725 -7223 1925 -7207
rect 1725 -7257 1741 -7223
rect 1909 -7257 1925 -7223
rect 1725 -7295 1925 -7257
rect 2097 -7223 2297 -7207
rect 2097 -7257 2113 -7223
rect 2281 -7257 2297 -7223
rect 2097 -7295 2297 -7257
rect 2469 -7223 2669 -7207
rect 2469 -7257 2485 -7223
rect 2653 -7257 2669 -7223
rect 2469 -7295 2669 -7257
rect 2841 -7223 3041 -7207
rect 2841 -7257 2857 -7223
rect 3025 -7257 3041 -7223
rect 2841 -7295 3041 -7257
rect 3213 -7223 3413 -7207
rect 3213 -7257 3229 -7223
rect 3397 -7257 3413 -7223
rect 3213 -7295 3413 -7257
rect 3585 -7223 3785 -7207
rect 3585 -7257 3601 -7223
rect 3769 -7257 3785 -7223
rect 3585 -7295 3785 -7257
rect 3957 -7223 4157 -7207
rect 3957 -7257 3973 -7223
rect 4141 -7257 4157 -7223
rect 3957 -7295 4157 -7257
rect 4329 -7223 4529 -7207
rect 4329 -7257 4345 -7223
rect 4513 -7257 4529 -7223
rect 4329 -7295 4529 -7257
rect 4701 -7223 4901 -7207
rect 4701 -7257 4717 -7223
rect 4885 -7257 4901 -7223
rect 4701 -7295 4901 -7257
rect 5073 -7223 5273 -7207
rect 5073 -7257 5089 -7223
rect 5257 -7257 5273 -7223
rect 5073 -7295 5273 -7257
rect 5445 -7223 5645 -7207
rect 5445 -7257 5461 -7223
rect 5629 -7257 5645 -7223
rect 5445 -7295 5645 -7257
rect 5817 -7223 6017 -7207
rect 5817 -7257 5833 -7223
rect 6001 -7257 6017 -7223
rect 5817 -7295 6017 -7257
rect 6189 -7223 6389 -7207
rect 6189 -7257 6205 -7223
rect 6373 -7257 6389 -7223
rect 6189 -7295 6389 -7257
rect 6561 -7223 6761 -7207
rect 6561 -7257 6577 -7223
rect 6745 -7257 6761 -7223
rect 6561 -7295 6761 -7257
rect 6933 -7223 7133 -7207
rect 6933 -7257 6949 -7223
rect 7117 -7257 7133 -7223
rect 6933 -7295 7133 -7257
rect 7305 -7223 7505 -7207
rect 7305 -7257 7321 -7223
rect 7489 -7257 7505 -7223
rect 7305 -7295 7505 -7257
rect 7677 -7223 7877 -7207
rect 7677 -7257 7693 -7223
rect 7861 -7257 7877 -7223
rect 7677 -7295 7877 -7257
rect 8049 -7223 8249 -7207
rect 8049 -7257 8065 -7223
rect 8233 -7257 8249 -7223
rect 8049 -7295 8249 -7257
rect 8421 -7223 8621 -7207
rect 8421 -7257 8437 -7223
rect 8605 -7257 8621 -7223
rect 8421 -7295 8621 -7257
rect 8793 -7223 8993 -7207
rect 8793 -7257 8809 -7223
rect 8977 -7257 8993 -7223
rect 8793 -7295 8993 -7257
rect 9165 -7223 9365 -7207
rect 9165 -7257 9181 -7223
rect 9349 -7257 9365 -7223
rect 9165 -7295 9365 -7257
rect 9537 -7223 9737 -7207
rect 9537 -7257 9553 -7223
rect 9721 -7257 9737 -7223
rect 9537 -7295 9737 -7257
rect 981 -7533 1181 -7495
rect 981 -7567 997 -7533
rect 1165 -7567 1181 -7533
rect 981 -7583 1181 -7567
rect 1353 -7533 1553 -7495
rect 1353 -7567 1369 -7533
rect 1537 -7567 1553 -7533
rect 1353 -7583 1553 -7567
rect 1725 -7533 1925 -7495
rect 1725 -7567 1741 -7533
rect 1909 -7567 1925 -7533
rect 1725 -7583 1925 -7567
rect 2097 -7533 2297 -7495
rect 2097 -7567 2113 -7533
rect 2281 -7567 2297 -7533
rect 2097 -7583 2297 -7567
rect 2469 -7533 2669 -7495
rect 2469 -7567 2485 -7533
rect 2653 -7567 2669 -7533
rect 2469 -7583 2669 -7567
rect 2841 -7533 3041 -7495
rect 2841 -7567 2857 -7533
rect 3025 -7567 3041 -7533
rect 2841 -7583 3041 -7567
rect 3213 -7533 3413 -7495
rect 3213 -7567 3229 -7533
rect 3397 -7567 3413 -7533
rect 3213 -7583 3413 -7567
rect 3585 -7533 3785 -7495
rect 3585 -7567 3601 -7533
rect 3769 -7567 3785 -7533
rect 3585 -7583 3785 -7567
rect 3957 -7533 4157 -7495
rect 3957 -7567 3973 -7533
rect 4141 -7567 4157 -7533
rect 3957 -7583 4157 -7567
rect 4329 -7533 4529 -7495
rect 4329 -7567 4345 -7533
rect 4513 -7567 4529 -7533
rect 4329 -7583 4529 -7567
rect 4701 -7533 4901 -7495
rect 4701 -7567 4717 -7533
rect 4885 -7567 4901 -7533
rect 4701 -7583 4901 -7567
rect 5073 -7533 5273 -7495
rect 5073 -7567 5089 -7533
rect 5257 -7567 5273 -7533
rect 5073 -7583 5273 -7567
rect 5445 -7533 5645 -7495
rect 5445 -7567 5461 -7533
rect 5629 -7567 5645 -7533
rect 5445 -7583 5645 -7567
rect 5817 -7533 6017 -7495
rect 5817 -7567 5833 -7533
rect 6001 -7567 6017 -7533
rect 5817 -7583 6017 -7567
rect 6189 -7533 6389 -7495
rect 6189 -7567 6205 -7533
rect 6373 -7567 6389 -7533
rect 6189 -7583 6389 -7567
rect 6561 -7533 6761 -7495
rect 6561 -7567 6577 -7533
rect 6745 -7567 6761 -7533
rect 6561 -7583 6761 -7567
rect 6933 -7533 7133 -7495
rect 6933 -7567 6949 -7533
rect 7117 -7567 7133 -7533
rect 6933 -7583 7133 -7567
rect 7305 -7533 7505 -7495
rect 7305 -7567 7321 -7533
rect 7489 -7567 7505 -7533
rect 7305 -7583 7505 -7567
rect 7677 -7533 7877 -7495
rect 7677 -7567 7693 -7533
rect 7861 -7567 7877 -7533
rect 7677 -7583 7877 -7567
rect 8049 -7533 8249 -7495
rect 8049 -7567 8065 -7533
rect 8233 -7567 8249 -7533
rect 8049 -7583 8249 -7567
rect 8421 -7533 8621 -7495
rect 8421 -7567 8437 -7533
rect 8605 -7567 8621 -7533
rect 8421 -7583 8621 -7567
rect 8793 -7533 8993 -7495
rect 8793 -7567 8809 -7533
rect 8977 -7567 8993 -7533
rect 8793 -7583 8993 -7567
rect 9165 -7533 9365 -7495
rect 9165 -7567 9181 -7533
rect 9349 -7567 9365 -7533
rect 9165 -7583 9365 -7567
rect 9537 -7533 9737 -7495
rect 9537 -7567 9553 -7533
rect 9721 -7567 9737 -7533
rect 9537 -7583 9737 -7567
<< polycont >>
rect -491 1079 -323 1113
rect -119 1079 49 1113
rect 253 1079 421 1113
rect 625 1079 793 1113
rect 997 1079 1165 1113
rect 1369 1079 1537 1113
rect 1741 1079 1909 1113
rect 2113 1079 2281 1113
rect 2485 1079 2653 1113
rect 2857 1079 3025 1113
rect 3229 1079 3397 1113
rect 3601 1079 3769 1113
rect 3973 1079 4141 1113
rect 4345 1079 4513 1113
rect 4717 1079 4885 1113
rect 5089 1079 5257 1113
rect 5461 1079 5629 1113
rect 5833 1079 6001 1113
rect 6205 1079 6373 1113
rect 6577 1079 6745 1113
rect 6949 1079 7117 1113
rect 7321 1079 7489 1113
rect 7693 1079 7861 1113
rect 8065 1079 8233 1113
rect 8437 1079 8605 1113
rect 8809 1079 8977 1113
rect 9181 1079 9349 1113
rect 9553 1079 9721 1113
rect 9925 1079 10093 1113
rect 10297 1079 10465 1113
rect 10669 1079 10837 1113
rect 11041 1079 11209 1113
rect -491 551 -323 585
rect -119 551 49 585
rect 253 551 421 585
rect 625 551 793 585
rect 997 551 1165 585
rect 1369 551 1537 585
rect 1741 551 1909 585
rect 2113 551 2281 585
rect 2485 551 2653 585
rect 2857 551 3025 585
rect 3229 551 3397 585
rect 3601 551 3769 585
rect 3973 551 4141 585
rect 4345 551 4513 585
rect 4717 551 4885 585
rect 5089 551 5257 585
rect 5461 551 5629 585
rect 5833 551 6001 585
rect 6205 551 6373 585
rect 6577 551 6745 585
rect 6949 551 7117 585
rect 7321 551 7489 585
rect 7693 551 7861 585
rect 8065 551 8233 585
rect 8437 551 8605 585
rect 8809 551 8977 585
rect 9181 551 9349 585
rect 9553 551 9721 585
rect 9925 551 10093 585
rect 10297 551 10465 585
rect 10669 551 10837 585
rect 11041 551 11209 585
rect -491 443 -323 477
rect -119 443 49 477
rect 253 443 421 477
rect 625 443 793 477
rect 997 443 1165 477
rect 1369 443 1537 477
rect 1741 443 1909 477
rect 2113 443 2281 477
rect 2485 443 2653 477
rect 2857 443 3025 477
rect 3229 443 3397 477
rect 3601 443 3769 477
rect 3973 443 4141 477
rect 4345 443 4513 477
rect 4717 443 4885 477
rect 5089 443 5257 477
rect 5461 443 5629 477
rect 5833 443 6001 477
rect 6205 443 6373 477
rect 6577 443 6745 477
rect 6949 443 7117 477
rect 7321 443 7489 477
rect 7693 443 7861 477
rect 8065 443 8233 477
rect 8437 443 8605 477
rect 8809 443 8977 477
rect 9181 443 9349 477
rect 9553 443 9721 477
rect 9925 443 10093 477
rect 10297 443 10465 477
rect 10669 443 10837 477
rect 11041 443 11209 477
rect -491 -85 -323 -51
rect -119 -85 49 -51
rect 253 -85 421 -51
rect 625 -85 793 -51
rect 997 -85 1165 -51
rect 1369 -85 1537 -51
rect 1741 -85 1909 -51
rect 2113 -85 2281 -51
rect 2485 -85 2653 -51
rect 2857 -85 3025 -51
rect 3229 -85 3397 -51
rect 3601 -85 3769 -51
rect 3973 -85 4141 -51
rect 4345 -85 4513 -51
rect 4717 -85 4885 -51
rect 5089 -85 5257 -51
rect 5461 -85 5629 -51
rect 5833 -85 6001 -51
rect 6205 -85 6373 -51
rect 6577 -85 6745 -51
rect 6949 -85 7117 -51
rect 7321 -85 7489 -51
rect 7693 -85 7861 -51
rect 8065 -85 8233 -51
rect 8437 -85 8605 -51
rect 8809 -85 8977 -51
rect 9181 -85 9349 -51
rect 9553 -85 9721 -51
rect 9925 -85 10093 -51
rect 10297 -85 10465 -51
rect 10669 -85 10837 -51
rect 11041 -85 11209 -51
rect -491 -193 -323 -159
rect -119 -193 49 -159
rect 253 -193 421 -159
rect 625 -193 793 -159
rect 997 -193 1165 -159
rect 1369 -193 1537 -159
rect 1741 -193 1909 -159
rect 2113 -193 2281 -159
rect 2485 -193 2653 -159
rect 2857 -193 3025 -159
rect 3229 -193 3397 -159
rect 3601 -193 3769 -159
rect 3973 -193 4141 -159
rect 4345 -193 4513 -159
rect 4717 -193 4885 -159
rect 5089 -193 5257 -159
rect 5461 -193 5629 -159
rect 5833 -193 6001 -159
rect 6205 -193 6373 -159
rect 6577 -193 6745 -159
rect 6949 -193 7117 -159
rect 7321 -193 7489 -159
rect 7693 -193 7861 -159
rect 8065 -193 8233 -159
rect 8437 -193 8605 -159
rect 8809 -193 8977 -159
rect 9181 -193 9349 -159
rect 9553 -193 9721 -159
rect 9925 -193 10093 -159
rect 10297 -193 10465 -159
rect 10669 -193 10837 -159
rect 11041 -193 11209 -159
rect -491 -721 -323 -687
rect -119 -721 49 -687
rect 253 -721 421 -687
rect 625 -721 793 -687
rect 997 -721 1165 -687
rect 1369 -721 1537 -687
rect 1741 -721 1909 -687
rect 2113 -721 2281 -687
rect 2485 -721 2653 -687
rect 2857 -721 3025 -687
rect 3229 -721 3397 -687
rect 3601 -721 3769 -687
rect 3973 -721 4141 -687
rect 4345 -721 4513 -687
rect 4717 -721 4885 -687
rect 5089 -721 5257 -687
rect 5461 -721 5629 -687
rect 5833 -721 6001 -687
rect 6205 -721 6373 -687
rect 6577 -721 6745 -687
rect 6949 -721 7117 -687
rect 7321 -721 7489 -687
rect 7693 -721 7861 -687
rect 8065 -721 8233 -687
rect 8437 -721 8605 -687
rect 8809 -721 8977 -687
rect 9181 -721 9349 -687
rect 9553 -721 9721 -687
rect 9925 -721 10093 -687
rect 10297 -721 10465 -687
rect 10669 -721 10837 -687
rect 11041 -721 11209 -687
rect 997 -1309 1165 -1275
rect 1369 -1309 1537 -1275
rect 1741 -1309 1909 -1275
rect 2113 -1309 2281 -1275
rect 2485 -1309 2653 -1275
rect 2857 -1309 3025 -1275
rect 3229 -1309 3397 -1275
rect 3601 -1309 3769 -1275
rect 997 -2237 1165 -2203
rect 1369 -2237 1537 -2203
rect 1741 -2237 1909 -2203
rect 2113 -2237 2281 -2203
rect 2485 -2237 2653 -2203
rect 2857 -2237 3025 -2203
rect 3229 -2237 3397 -2203
rect 3601 -2237 3769 -2203
rect 997 -2345 1165 -2311
rect 1369 -2345 1537 -2311
rect 1741 -2345 1909 -2311
rect 2113 -2345 2281 -2311
rect 2485 -2345 2653 -2311
rect 2857 -2345 3025 -2311
rect 3229 -2345 3397 -2311
rect 3601 -2345 3769 -2311
rect 997 -3273 1165 -3239
rect 1369 -3273 1537 -3239
rect 1741 -3273 1909 -3239
rect 2113 -3273 2281 -3239
rect 2485 -3273 2653 -3239
rect 2857 -3273 3025 -3239
rect 3229 -3273 3397 -3239
rect 3601 -3273 3769 -3239
rect 997 -3381 1165 -3347
rect 1369 -3381 1537 -3347
rect 1741 -3381 1909 -3347
rect 2113 -3381 2281 -3347
rect 2485 -3381 2653 -3347
rect 2857 -3381 3025 -3347
rect 3229 -3381 3397 -3347
rect 3601 -3381 3769 -3347
rect 997 -4309 1165 -4275
rect 1369 -4309 1537 -4275
rect 1741 -4309 1909 -4275
rect 2113 -4309 2281 -4275
rect 2485 -4309 2653 -4275
rect 2857 -4309 3025 -4275
rect 3229 -4309 3397 -4275
rect 3601 -4309 3769 -4275
rect 997 -4417 1165 -4383
rect 1369 -4417 1537 -4383
rect 1741 -4417 1909 -4383
rect 2113 -4417 2281 -4383
rect 2485 -4417 2653 -4383
rect 2857 -4417 3025 -4383
rect 3229 -4417 3397 -4383
rect 3601 -4417 3769 -4383
rect 997 -5345 1165 -5311
rect 1369 -5345 1537 -5311
rect 1741 -5345 1909 -5311
rect 2113 -5345 2281 -5311
rect 2485 -5345 2653 -5311
rect 2857 -5345 3025 -5311
rect 3229 -5345 3397 -5311
rect 3601 -5345 3769 -5311
rect 997 -6003 1165 -5969
rect 1369 -6003 1537 -5969
rect 1741 -6003 1909 -5969
rect 2113 -6003 2281 -5969
rect 2485 -6003 2653 -5969
rect 2857 -6003 3025 -5969
rect 3229 -6003 3397 -5969
rect 3601 -6003 3769 -5969
rect 3973 -6003 4141 -5969
rect 4345 -6003 4513 -5969
rect 4717 -6003 4885 -5969
rect 5089 -6003 5257 -5969
rect 5461 -6003 5629 -5969
rect 5833 -6003 6001 -5969
rect 6205 -6003 6373 -5969
rect 6577 -6003 6745 -5969
rect 6949 -6003 7117 -5969
rect 7321 -6003 7489 -5969
rect 7693 -6003 7861 -5969
rect 8065 -6003 8233 -5969
rect 8437 -6003 8605 -5969
rect 8809 -6003 8977 -5969
rect 9181 -6003 9349 -5969
rect 9553 -6003 9721 -5969
rect 997 -6313 1165 -6279
rect 1369 -6313 1537 -6279
rect 1741 -6313 1909 -6279
rect 2113 -6313 2281 -6279
rect 2485 -6313 2653 -6279
rect 2857 -6313 3025 -6279
rect 3229 -6313 3397 -6279
rect 3601 -6313 3769 -6279
rect 3973 -6313 4141 -6279
rect 4345 -6313 4513 -6279
rect 4717 -6313 4885 -6279
rect 5089 -6313 5257 -6279
rect 5461 -6313 5629 -6279
rect 5833 -6313 6001 -6279
rect 6205 -6313 6373 -6279
rect 6577 -6313 6745 -6279
rect 6949 -6313 7117 -6279
rect 7321 -6313 7489 -6279
rect 7693 -6313 7861 -6279
rect 8065 -6313 8233 -6279
rect 8437 -6313 8605 -6279
rect 8809 -6313 8977 -6279
rect 9181 -6313 9349 -6279
rect 9553 -6313 9721 -6279
rect 997 -6421 1165 -6387
rect 1369 -6421 1537 -6387
rect 1741 -6421 1909 -6387
rect 2113 -6421 2281 -6387
rect 2485 -6421 2653 -6387
rect 2857 -6421 3025 -6387
rect 3229 -6421 3397 -6387
rect 3601 -6421 3769 -6387
rect 3973 -6421 4141 -6387
rect 4345 -6421 4513 -6387
rect 4717 -6421 4885 -6387
rect 5089 -6421 5257 -6387
rect 5461 -6421 5629 -6387
rect 5833 -6421 6001 -6387
rect 6205 -6421 6373 -6387
rect 6577 -6421 6745 -6387
rect 6949 -6421 7117 -6387
rect 7321 -6421 7489 -6387
rect 7693 -6421 7861 -6387
rect 8065 -6421 8233 -6387
rect 8437 -6421 8605 -6387
rect 8809 -6421 8977 -6387
rect 9181 -6421 9349 -6387
rect 9553 -6421 9721 -6387
rect 997 -6731 1165 -6697
rect 1369 -6731 1537 -6697
rect 1741 -6731 1909 -6697
rect 2113 -6731 2281 -6697
rect 2485 -6731 2653 -6697
rect 2857 -6731 3025 -6697
rect 3229 -6731 3397 -6697
rect 3601 -6731 3769 -6697
rect 3973 -6731 4141 -6697
rect 4345 -6731 4513 -6697
rect 4717 -6731 4885 -6697
rect 5089 -6731 5257 -6697
rect 5461 -6731 5629 -6697
rect 5833 -6731 6001 -6697
rect 6205 -6731 6373 -6697
rect 6577 -6731 6745 -6697
rect 6949 -6731 7117 -6697
rect 7321 -6731 7489 -6697
rect 7693 -6731 7861 -6697
rect 8065 -6731 8233 -6697
rect 8437 -6731 8605 -6697
rect 8809 -6731 8977 -6697
rect 9181 -6731 9349 -6697
rect 9553 -6731 9721 -6697
rect 997 -6839 1165 -6805
rect 1369 -6839 1537 -6805
rect 1741 -6839 1909 -6805
rect 2113 -6839 2281 -6805
rect 2485 -6839 2653 -6805
rect 2857 -6839 3025 -6805
rect 3229 -6839 3397 -6805
rect 3601 -6839 3769 -6805
rect 3973 -6839 4141 -6805
rect 4345 -6839 4513 -6805
rect 4717 -6839 4885 -6805
rect 5089 -6839 5257 -6805
rect 5461 -6839 5629 -6805
rect 5833 -6839 6001 -6805
rect 6205 -6839 6373 -6805
rect 6577 -6839 6745 -6805
rect 6949 -6839 7117 -6805
rect 7321 -6839 7489 -6805
rect 7693 -6839 7861 -6805
rect 8065 -6839 8233 -6805
rect 8437 -6839 8605 -6805
rect 8809 -6839 8977 -6805
rect 9181 -6839 9349 -6805
rect 9553 -6839 9721 -6805
rect 997 -7149 1165 -7115
rect 1369 -7149 1537 -7115
rect 1741 -7149 1909 -7115
rect 2113 -7149 2281 -7115
rect 2485 -7149 2653 -7115
rect 2857 -7149 3025 -7115
rect 3229 -7149 3397 -7115
rect 3601 -7149 3769 -7115
rect 3973 -7149 4141 -7115
rect 4345 -7149 4513 -7115
rect 4717 -7149 4885 -7115
rect 5089 -7149 5257 -7115
rect 5461 -7149 5629 -7115
rect 5833 -7149 6001 -7115
rect 6205 -7149 6373 -7115
rect 6577 -7149 6745 -7115
rect 6949 -7149 7117 -7115
rect 7321 -7149 7489 -7115
rect 7693 -7149 7861 -7115
rect 8065 -7149 8233 -7115
rect 8437 -7149 8605 -7115
rect 8809 -7149 8977 -7115
rect 9181 -7149 9349 -7115
rect 9553 -7149 9721 -7115
rect 997 -7257 1165 -7223
rect 1369 -7257 1537 -7223
rect 1741 -7257 1909 -7223
rect 2113 -7257 2281 -7223
rect 2485 -7257 2653 -7223
rect 2857 -7257 3025 -7223
rect 3229 -7257 3397 -7223
rect 3601 -7257 3769 -7223
rect 3973 -7257 4141 -7223
rect 4345 -7257 4513 -7223
rect 4717 -7257 4885 -7223
rect 5089 -7257 5257 -7223
rect 5461 -7257 5629 -7223
rect 5833 -7257 6001 -7223
rect 6205 -7257 6373 -7223
rect 6577 -7257 6745 -7223
rect 6949 -7257 7117 -7223
rect 7321 -7257 7489 -7223
rect 7693 -7257 7861 -7223
rect 8065 -7257 8233 -7223
rect 8437 -7257 8605 -7223
rect 8809 -7257 8977 -7223
rect 9181 -7257 9349 -7223
rect 9553 -7257 9721 -7223
rect 997 -7567 1165 -7533
rect 1369 -7567 1537 -7533
rect 1741 -7567 1909 -7533
rect 2113 -7567 2281 -7533
rect 2485 -7567 2653 -7533
rect 2857 -7567 3025 -7533
rect 3229 -7567 3397 -7533
rect 3601 -7567 3769 -7533
rect 3973 -7567 4141 -7533
rect 4345 -7567 4513 -7533
rect 4717 -7567 4885 -7533
rect 5089 -7567 5257 -7533
rect 5461 -7567 5629 -7533
rect 5833 -7567 6001 -7533
rect 6205 -7567 6373 -7533
rect 6577 -7567 6745 -7533
rect 6949 -7567 7117 -7533
rect 7321 -7567 7489 -7533
rect 7693 -7567 7861 -7533
rect 8065 -7567 8233 -7533
rect 8437 -7567 8605 -7533
rect 8809 -7567 8977 -7533
rect 9181 -7567 9349 -7533
rect 9553 -7567 9721 -7533
<< xpolycontact >>
rect 6115 -3891 6185 -3459
rect 6115 -4423 6185 -3991
<< xpolyres >>
rect 6115 -3991 6185 -3891
<< locali >>
rect -667 1181 -571 1215
rect 11292 1181 11385 1215
rect -667 1119 -633 1181
rect 11351 1119 11385 1181
rect -507 1079 -491 1113
rect -323 1079 -307 1113
rect -135 1079 -119 1113
rect 49 1079 65 1113
rect 237 1079 253 1113
rect 421 1079 437 1113
rect 609 1079 625 1113
rect 793 1079 809 1113
rect 981 1079 997 1113
rect 1165 1079 1181 1113
rect 1353 1079 1369 1113
rect 1537 1079 1553 1113
rect 1725 1079 1741 1113
rect 1909 1079 1925 1113
rect 2097 1079 2113 1113
rect 2281 1079 2297 1113
rect 2469 1079 2485 1113
rect 2653 1079 2669 1113
rect 2841 1079 2857 1113
rect 3025 1079 3041 1113
rect 3213 1079 3229 1113
rect 3397 1079 3413 1113
rect 3585 1079 3601 1113
rect 3769 1079 3785 1113
rect 3957 1079 3973 1113
rect 4141 1079 4157 1113
rect 4329 1079 4345 1113
rect 4513 1079 4529 1113
rect 4701 1079 4717 1113
rect 4885 1079 4901 1113
rect 5073 1079 5089 1113
rect 5257 1079 5273 1113
rect 5445 1079 5461 1113
rect 5629 1079 5645 1113
rect 5817 1079 5833 1113
rect 6001 1079 6017 1113
rect 6189 1079 6205 1113
rect 6373 1079 6389 1113
rect 6561 1079 6577 1113
rect 6745 1079 6761 1113
rect 6933 1079 6949 1113
rect 7117 1079 7133 1113
rect 7305 1079 7321 1113
rect 7489 1079 7505 1113
rect 7677 1079 7693 1113
rect 7861 1079 7877 1113
rect 8049 1079 8065 1113
rect 8233 1079 8249 1113
rect 8421 1079 8437 1113
rect 8605 1079 8621 1113
rect 8793 1079 8809 1113
rect 8977 1079 8993 1113
rect 9165 1079 9181 1113
rect 9349 1079 9365 1113
rect 9537 1079 9553 1113
rect 9721 1079 9737 1113
rect 9909 1079 9925 1113
rect 10093 1079 10109 1113
rect 10281 1079 10297 1113
rect 10465 1079 10481 1113
rect 10653 1079 10669 1113
rect 10837 1079 10853 1113
rect 11025 1079 11041 1113
rect 11209 1079 11225 1113
rect -553 1020 -519 1036
rect -553 628 -519 644
rect -295 1020 -261 1036
rect -295 628 -261 644
rect -181 1020 -147 1036
rect -181 628 -147 644
rect 77 1020 111 1036
rect 77 628 111 644
rect 191 1020 225 1036
rect 191 628 225 644
rect 449 1020 483 1036
rect 449 628 483 644
rect 563 1020 597 1036
rect 563 628 597 644
rect 821 1020 855 1036
rect 821 628 855 644
rect 935 1020 969 1036
rect 935 628 969 644
rect 1193 1020 1227 1036
rect 1193 628 1227 644
rect 1307 1020 1341 1036
rect 1307 628 1341 644
rect 1565 1020 1599 1036
rect 1565 628 1599 644
rect 1679 1020 1713 1036
rect 1679 628 1713 644
rect 1937 1020 1971 1036
rect 1937 628 1971 644
rect 2051 1020 2085 1036
rect 2051 628 2085 644
rect 2309 1020 2343 1036
rect 2309 628 2343 644
rect 2423 1020 2457 1036
rect 2423 628 2457 644
rect 2681 1020 2715 1036
rect 2681 628 2715 644
rect 2795 1020 2829 1036
rect 2795 628 2829 644
rect 3053 1020 3087 1036
rect 3053 628 3087 644
rect 3167 1020 3201 1036
rect 3167 628 3201 644
rect 3425 1020 3459 1036
rect 3425 628 3459 644
rect 3539 1020 3573 1036
rect 3539 628 3573 644
rect 3797 1020 3831 1036
rect 3797 628 3831 644
rect 3911 1020 3945 1036
rect 3911 628 3945 644
rect 4169 1020 4203 1036
rect 4169 628 4203 644
rect 4283 1020 4317 1036
rect 4283 628 4317 644
rect 4541 1020 4575 1036
rect 4541 628 4575 644
rect 4655 1020 4689 1036
rect 4655 628 4689 644
rect 4913 1020 4947 1036
rect 4913 628 4947 644
rect 5027 1020 5061 1036
rect 5027 628 5061 644
rect 5285 1020 5319 1036
rect 5285 628 5319 644
rect 5399 1020 5433 1036
rect 5399 628 5433 644
rect 5657 1020 5691 1036
rect 5657 628 5691 644
rect 5771 1020 5805 1036
rect 5771 628 5805 644
rect 6029 1020 6063 1036
rect 6029 628 6063 644
rect 6143 1020 6177 1036
rect 6143 628 6177 644
rect 6401 1020 6435 1036
rect 6401 628 6435 644
rect 6515 1020 6549 1036
rect 6515 628 6549 644
rect 6773 1020 6807 1036
rect 6773 628 6807 644
rect 6887 1020 6921 1036
rect 6887 628 6921 644
rect 7145 1020 7179 1036
rect 7145 628 7179 644
rect 7259 1020 7293 1036
rect 7259 628 7293 644
rect 7517 1020 7551 1036
rect 7517 628 7551 644
rect 7631 1020 7665 1036
rect 7631 628 7665 644
rect 7889 1020 7923 1036
rect 7889 628 7923 644
rect 8003 1020 8037 1036
rect 8003 628 8037 644
rect 8261 1020 8295 1036
rect 8261 628 8295 644
rect 8375 1020 8409 1036
rect 8375 628 8409 644
rect 8633 1020 8667 1036
rect 8633 628 8667 644
rect 8747 1020 8781 1036
rect 8747 628 8781 644
rect 9005 1020 9039 1036
rect 9005 628 9039 644
rect 9119 1020 9153 1036
rect 9119 628 9153 644
rect 9377 1020 9411 1036
rect 9377 628 9411 644
rect 9491 1020 9525 1036
rect 9491 628 9525 644
rect 9749 1020 9783 1036
rect 9749 628 9783 644
rect 9863 1020 9897 1036
rect 9863 628 9897 644
rect 10121 1020 10155 1036
rect 10121 628 10155 644
rect 10235 1020 10269 1036
rect 10235 628 10269 644
rect 10493 1020 10527 1036
rect 10493 628 10527 644
rect 10607 1020 10641 1036
rect 10607 628 10641 644
rect 10865 1020 10899 1036
rect 10865 628 10899 644
rect 10979 1020 11013 1036
rect 10979 628 11013 644
rect 11237 1020 11271 1036
rect 11237 628 11271 644
rect -507 551 -491 585
rect -323 551 -307 585
rect -135 551 -119 585
rect 49 551 65 585
rect 237 551 253 585
rect 421 551 437 585
rect 609 551 625 585
rect 793 551 809 585
rect 981 551 997 585
rect 1165 551 1181 585
rect 1353 551 1369 585
rect 1537 551 1553 585
rect 1725 551 1741 585
rect 1909 551 1925 585
rect 2097 551 2113 585
rect 2281 551 2297 585
rect 2469 551 2485 585
rect 2653 551 2669 585
rect 2841 551 2857 585
rect 3025 551 3041 585
rect 3213 551 3229 585
rect 3397 551 3413 585
rect 3585 551 3601 585
rect 3769 551 3785 585
rect 3957 551 3973 585
rect 4141 551 4157 585
rect 4329 551 4345 585
rect 4513 551 4529 585
rect 4701 551 4717 585
rect 4885 551 4901 585
rect 5073 551 5089 585
rect 5257 551 5273 585
rect 5445 551 5461 585
rect 5629 551 5645 585
rect 5817 551 5833 585
rect 6001 551 6017 585
rect 6189 551 6205 585
rect 6373 551 6389 585
rect 6561 551 6577 585
rect 6745 551 6761 585
rect 6933 551 6949 585
rect 7117 551 7133 585
rect 7305 551 7321 585
rect 7489 551 7505 585
rect 7677 551 7693 585
rect 7861 551 7877 585
rect 8049 551 8065 585
rect 8233 551 8249 585
rect 8421 551 8437 585
rect 8605 551 8621 585
rect 8793 551 8809 585
rect 8977 551 8993 585
rect 9165 551 9181 585
rect 9349 551 9365 585
rect 9537 551 9553 585
rect 9721 551 9737 585
rect 9909 551 9925 585
rect 10093 551 10109 585
rect 10281 551 10297 585
rect 10465 551 10481 585
rect 10653 551 10669 585
rect 10837 551 10853 585
rect 11025 551 11041 585
rect 11209 551 11225 585
rect -507 443 -491 477
rect -323 443 -307 477
rect -135 443 -119 477
rect 49 443 65 477
rect 237 443 253 477
rect 421 443 437 477
rect 609 443 625 477
rect 793 443 809 477
rect 981 443 997 477
rect 1165 443 1181 477
rect 1353 443 1369 477
rect 1537 443 1553 477
rect 1725 443 1741 477
rect 1909 443 1925 477
rect 2097 443 2113 477
rect 2281 443 2297 477
rect 2469 443 2485 477
rect 2653 443 2669 477
rect 2841 443 2857 477
rect 3025 443 3041 477
rect 3213 443 3229 477
rect 3397 443 3413 477
rect 3585 443 3601 477
rect 3769 443 3785 477
rect 3957 443 3973 477
rect 4141 443 4157 477
rect 4329 443 4345 477
rect 4513 443 4529 477
rect 4701 443 4717 477
rect 4885 443 4901 477
rect 5073 443 5089 477
rect 5257 443 5273 477
rect 5445 443 5461 477
rect 5629 443 5645 477
rect 5817 443 5833 477
rect 6001 443 6017 477
rect 6189 443 6205 477
rect 6373 443 6389 477
rect 6561 443 6577 477
rect 6745 443 6761 477
rect 6933 443 6949 477
rect 7117 443 7133 477
rect 7305 443 7321 477
rect 7489 443 7505 477
rect 7677 443 7693 477
rect 7861 443 7877 477
rect 8049 443 8065 477
rect 8233 443 8249 477
rect 8421 443 8437 477
rect 8605 443 8621 477
rect 8793 443 8809 477
rect 8977 443 8993 477
rect 9165 443 9181 477
rect 9349 443 9365 477
rect 9537 443 9553 477
rect 9721 443 9737 477
rect 9909 443 9925 477
rect 10093 443 10109 477
rect 10281 443 10297 477
rect 10465 443 10481 477
rect 10653 443 10669 477
rect 10837 443 10853 477
rect 11025 443 11041 477
rect 11209 443 11225 477
rect -553 384 -519 400
rect -553 -8 -519 8
rect -295 384 -261 400
rect -295 -8 -261 8
rect -181 384 -147 400
rect -181 -8 -147 8
rect 77 384 111 400
rect 77 -8 111 8
rect 191 384 225 400
rect 191 -8 225 8
rect 449 384 483 400
rect 449 -8 483 8
rect 563 384 597 400
rect 563 -8 597 8
rect 821 384 855 400
rect 821 -8 855 8
rect 935 384 969 400
rect 935 -8 969 8
rect 1193 384 1227 400
rect 1193 -8 1227 8
rect 1307 384 1341 400
rect 1307 -8 1341 8
rect 1565 384 1599 400
rect 1565 -8 1599 8
rect 1679 384 1713 400
rect 1679 -8 1713 8
rect 1937 384 1971 400
rect 1937 -8 1971 8
rect 2051 384 2085 400
rect 2051 -8 2085 8
rect 2309 384 2343 400
rect 2309 -8 2343 8
rect 2423 384 2457 400
rect 2423 -8 2457 8
rect 2681 384 2715 400
rect 2681 -8 2715 8
rect 2795 384 2829 400
rect 2795 -8 2829 8
rect 3053 384 3087 400
rect 3053 -8 3087 8
rect 3167 384 3201 400
rect 3167 -8 3201 8
rect 3425 384 3459 400
rect 3425 -8 3459 8
rect 3539 384 3573 400
rect 3539 -8 3573 8
rect 3797 384 3831 400
rect 3797 -8 3831 8
rect 3911 384 3945 400
rect 3911 -8 3945 8
rect 4169 384 4203 400
rect 4169 -8 4203 8
rect 4283 384 4317 400
rect 4283 -8 4317 8
rect 4541 384 4575 400
rect 4541 -8 4575 8
rect 4655 384 4689 400
rect 4655 -8 4689 8
rect 4913 384 4947 400
rect 4913 -8 4947 8
rect 5027 384 5061 400
rect 5027 -8 5061 8
rect 5285 384 5319 400
rect 5285 -8 5319 8
rect 5399 384 5433 400
rect 5399 -8 5433 8
rect 5657 384 5691 400
rect 5657 -8 5691 8
rect 5771 384 5805 400
rect 5771 -8 5805 8
rect 6029 384 6063 400
rect 6029 -8 6063 8
rect 6143 384 6177 400
rect 6143 -8 6177 8
rect 6401 384 6435 400
rect 6401 -8 6435 8
rect 6515 384 6549 400
rect 6515 -8 6549 8
rect 6773 384 6807 400
rect 6773 -8 6807 8
rect 6887 384 6921 400
rect 6887 -8 6921 8
rect 7145 384 7179 400
rect 7145 -8 7179 8
rect 7259 384 7293 400
rect 7259 -8 7293 8
rect 7517 384 7551 400
rect 7517 -8 7551 8
rect 7631 384 7665 400
rect 7631 -8 7665 8
rect 7889 384 7923 400
rect 7889 -8 7923 8
rect 8003 384 8037 400
rect 8003 -8 8037 8
rect 8261 384 8295 400
rect 8261 -8 8295 8
rect 8375 384 8409 400
rect 8375 -8 8409 8
rect 8633 384 8667 400
rect 8633 -8 8667 8
rect 8747 384 8781 400
rect 8747 -8 8781 8
rect 9005 384 9039 400
rect 9005 -8 9039 8
rect 9119 384 9153 400
rect 9119 -8 9153 8
rect 9377 384 9411 400
rect 9377 -8 9411 8
rect 9491 384 9525 400
rect 9491 -8 9525 8
rect 9749 384 9783 400
rect 9749 -8 9783 8
rect 9863 384 9897 400
rect 9863 -8 9897 8
rect 10121 384 10155 400
rect 10121 -8 10155 8
rect 10235 384 10269 400
rect 10235 -8 10269 8
rect 10493 384 10527 400
rect 10493 -8 10527 8
rect 10607 384 10641 400
rect 10607 -8 10641 8
rect 10865 384 10899 400
rect 10865 -8 10899 8
rect 10979 384 11013 400
rect 10979 -8 11013 8
rect 11237 384 11271 400
rect 11237 -8 11271 8
rect -507 -85 -491 -51
rect -323 -85 -307 -51
rect -135 -85 -119 -51
rect 49 -85 65 -51
rect 237 -85 253 -51
rect 421 -85 437 -51
rect 609 -85 625 -51
rect 793 -85 809 -51
rect 981 -85 997 -51
rect 1165 -85 1181 -51
rect 1353 -85 1369 -51
rect 1537 -85 1553 -51
rect 1725 -85 1741 -51
rect 1909 -85 1925 -51
rect 2097 -85 2113 -51
rect 2281 -85 2297 -51
rect 2469 -85 2485 -51
rect 2653 -85 2669 -51
rect 2841 -85 2857 -51
rect 3025 -85 3041 -51
rect 3213 -85 3229 -51
rect 3397 -85 3413 -51
rect 3585 -85 3601 -51
rect 3769 -85 3785 -51
rect 3957 -85 3973 -51
rect 4141 -85 4157 -51
rect 4329 -85 4345 -51
rect 4513 -85 4529 -51
rect 4701 -85 4717 -51
rect 4885 -85 4901 -51
rect 5073 -85 5089 -51
rect 5257 -85 5273 -51
rect 5445 -85 5461 -51
rect 5629 -85 5645 -51
rect 5817 -85 5833 -51
rect 6001 -85 6017 -51
rect 6189 -85 6205 -51
rect 6373 -85 6389 -51
rect 6561 -85 6577 -51
rect 6745 -85 6761 -51
rect 6933 -85 6949 -51
rect 7117 -85 7133 -51
rect 7305 -85 7321 -51
rect 7489 -85 7505 -51
rect 7677 -85 7693 -51
rect 7861 -85 7877 -51
rect 8049 -85 8065 -51
rect 8233 -85 8249 -51
rect 8421 -85 8437 -51
rect 8605 -85 8621 -51
rect 8793 -85 8809 -51
rect 8977 -85 8993 -51
rect 9165 -85 9181 -51
rect 9349 -85 9365 -51
rect 9537 -85 9553 -51
rect 9721 -85 9737 -51
rect 9909 -85 9925 -51
rect 10093 -85 10109 -51
rect 10281 -85 10297 -51
rect 10465 -85 10481 -51
rect 10653 -85 10669 -51
rect 10837 -85 10853 -51
rect 11025 -85 11041 -51
rect 11209 -85 11225 -51
rect -507 -193 -491 -159
rect -323 -193 -307 -159
rect -135 -193 -119 -159
rect 49 -193 65 -159
rect 237 -193 253 -159
rect 421 -193 437 -159
rect 609 -193 625 -159
rect 793 -193 809 -159
rect 981 -193 997 -159
rect 1165 -193 1181 -159
rect 1353 -193 1369 -159
rect 1537 -193 1553 -159
rect 1725 -193 1741 -159
rect 1909 -193 1925 -159
rect 2097 -193 2113 -159
rect 2281 -193 2297 -159
rect 2469 -193 2485 -159
rect 2653 -193 2669 -159
rect 2841 -193 2857 -159
rect 3025 -193 3041 -159
rect 3213 -193 3229 -159
rect 3397 -193 3413 -159
rect 3585 -193 3601 -159
rect 3769 -193 3785 -159
rect 3957 -193 3973 -159
rect 4141 -193 4157 -159
rect 4329 -193 4345 -159
rect 4513 -193 4529 -159
rect 4701 -193 4717 -159
rect 4885 -193 4901 -159
rect 5073 -193 5089 -159
rect 5257 -193 5273 -159
rect 5445 -193 5461 -159
rect 5629 -193 5645 -159
rect 5817 -193 5833 -159
rect 6001 -193 6017 -159
rect 6189 -193 6205 -159
rect 6373 -193 6389 -159
rect 6561 -193 6577 -159
rect 6745 -193 6761 -159
rect 6933 -193 6949 -159
rect 7117 -193 7133 -159
rect 7305 -193 7321 -159
rect 7489 -193 7505 -159
rect 7677 -193 7693 -159
rect 7861 -193 7877 -159
rect 8049 -193 8065 -159
rect 8233 -193 8249 -159
rect 8421 -193 8437 -159
rect 8605 -193 8621 -159
rect 8793 -193 8809 -159
rect 8977 -193 8993 -159
rect 9165 -193 9181 -159
rect 9349 -193 9365 -159
rect 9537 -193 9553 -159
rect 9721 -193 9737 -159
rect 9909 -193 9925 -159
rect 10093 -193 10109 -159
rect 10281 -193 10297 -159
rect 10465 -193 10481 -159
rect 10653 -193 10669 -159
rect 10837 -193 10853 -159
rect 11025 -193 11041 -159
rect 11209 -193 11225 -159
rect -553 -252 -519 -236
rect -553 -644 -519 -628
rect -295 -252 -261 -236
rect -295 -644 -261 -628
rect -181 -252 -147 -236
rect -181 -644 -147 -628
rect 77 -252 111 -236
rect 77 -644 111 -628
rect 191 -252 225 -236
rect 191 -644 225 -628
rect 449 -252 483 -236
rect 449 -644 483 -628
rect 563 -252 597 -236
rect 563 -644 597 -628
rect 821 -252 855 -236
rect 821 -644 855 -628
rect 935 -252 969 -236
rect 935 -644 969 -628
rect 1193 -252 1227 -236
rect 1193 -644 1227 -628
rect 1307 -252 1341 -236
rect 1307 -644 1341 -628
rect 1565 -252 1599 -236
rect 1565 -644 1599 -628
rect 1679 -252 1713 -236
rect 1679 -644 1713 -628
rect 1937 -252 1971 -236
rect 1937 -644 1971 -628
rect 2051 -252 2085 -236
rect 2051 -644 2085 -628
rect 2309 -252 2343 -236
rect 2309 -644 2343 -628
rect 2423 -252 2457 -236
rect 2423 -644 2457 -628
rect 2681 -252 2715 -236
rect 2681 -644 2715 -628
rect 2795 -252 2829 -236
rect 2795 -644 2829 -628
rect 3053 -252 3087 -236
rect 3053 -644 3087 -628
rect 3167 -252 3201 -236
rect 3167 -644 3201 -628
rect 3425 -252 3459 -236
rect 3425 -644 3459 -628
rect 3539 -252 3573 -236
rect 3539 -644 3573 -628
rect 3797 -252 3831 -236
rect 3797 -644 3831 -628
rect 3911 -252 3945 -236
rect 3911 -644 3945 -628
rect 4169 -252 4203 -236
rect 4169 -644 4203 -628
rect 4283 -252 4317 -236
rect 4283 -644 4317 -628
rect 4541 -252 4575 -236
rect 4541 -644 4575 -628
rect 4655 -252 4689 -236
rect 4655 -644 4689 -628
rect 4913 -252 4947 -236
rect 4913 -644 4947 -628
rect 5027 -252 5061 -236
rect 5027 -644 5061 -628
rect 5285 -252 5319 -236
rect 5285 -644 5319 -628
rect 5399 -252 5433 -236
rect 5399 -644 5433 -628
rect 5657 -252 5691 -236
rect 5657 -644 5691 -628
rect 5771 -252 5805 -236
rect 5771 -644 5805 -628
rect 6029 -252 6063 -236
rect 6029 -644 6063 -628
rect 6143 -252 6177 -236
rect 6143 -644 6177 -628
rect 6401 -252 6435 -236
rect 6401 -644 6435 -628
rect 6515 -252 6549 -236
rect 6515 -644 6549 -628
rect 6773 -252 6807 -236
rect 6773 -644 6807 -628
rect 6887 -252 6921 -236
rect 6887 -644 6921 -628
rect 7145 -252 7179 -236
rect 7145 -644 7179 -628
rect 7259 -252 7293 -236
rect 7259 -644 7293 -628
rect 7517 -252 7551 -236
rect 7517 -644 7551 -628
rect 7631 -252 7665 -236
rect 7631 -644 7665 -628
rect 7889 -252 7923 -236
rect 7889 -644 7923 -628
rect 8003 -252 8037 -236
rect 8003 -644 8037 -628
rect 8261 -252 8295 -236
rect 8261 -644 8295 -628
rect 8375 -252 8409 -236
rect 8375 -644 8409 -628
rect 8633 -252 8667 -236
rect 8633 -644 8667 -628
rect 8747 -252 8781 -236
rect 8747 -644 8781 -628
rect 9005 -252 9039 -236
rect 9005 -644 9039 -628
rect 9119 -252 9153 -236
rect 9119 -644 9153 -628
rect 9377 -252 9411 -236
rect 9377 -644 9411 -628
rect 9491 -252 9525 -236
rect 9491 -644 9525 -628
rect 9749 -252 9783 -236
rect 9749 -644 9783 -628
rect 9863 -252 9897 -236
rect 9863 -644 9897 -628
rect 10121 -252 10155 -236
rect 10121 -644 10155 -628
rect 10235 -252 10269 -236
rect 10235 -644 10269 -628
rect 10493 -252 10527 -236
rect 10493 -644 10527 -628
rect 10607 -252 10641 -236
rect 10607 -644 10641 -628
rect 10865 -252 10899 -236
rect 10865 -644 10899 -628
rect 10979 -252 11013 -236
rect 10979 -644 11013 -628
rect 11237 -252 11271 -236
rect 11237 -644 11271 -628
rect -507 -721 -491 -687
rect -323 -721 -307 -687
rect -135 -721 -119 -687
rect 49 -721 65 -687
rect 237 -721 253 -687
rect 421 -721 437 -687
rect 609 -721 625 -687
rect 793 -721 809 -687
rect 981 -721 997 -687
rect 1165 -721 1181 -687
rect 1353 -721 1369 -687
rect 1537 -721 1553 -687
rect 1725 -721 1741 -687
rect 1909 -721 1925 -687
rect 2097 -721 2113 -687
rect 2281 -721 2297 -687
rect 2469 -721 2485 -687
rect 2653 -721 2669 -687
rect 2841 -721 2857 -687
rect 3025 -721 3041 -687
rect 3213 -721 3229 -687
rect 3397 -721 3413 -687
rect 3585 -721 3601 -687
rect 3769 -721 3785 -687
rect 3957 -721 3973 -687
rect 4141 -721 4157 -687
rect 4329 -721 4345 -687
rect 4513 -721 4529 -687
rect 4701 -721 4717 -687
rect 4885 -721 4901 -687
rect 5073 -721 5089 -687
rect 5257 -721 5273 -687
rect 5445 -721 5461 -687
rect 5629 -721 5645 -687
rect 5817 -721 5833 -687
rect 6001 -721 6017 -687
rect 6189 -721 6205 -687
rect 6373 -721 6389 -687
rect 6561 -721 6577 -687
rect 6745 -721 6761 -687
rect 6933 -721 6949 -687
rect 7117 -721 7133 -687
rect 7305 -721 7321 -687
rect 7489 -721 7505 -687
rect 7677 -721 7693 -687
rect 7861 -721 7877 -687
rect 8049 -721 8065 -687
rect 8233 -721 8249 -687
rect 8421 -721 8437 -687
rect 8605 -721 8621 -687
rect 8793 -721 8809 -687
rect 8977 -721 8993 -687
rect 9165 -721 9181 -687
rect 9349 -721 9365 -687
rect 9537 -721 9553 -687
rect 9721 -721 9737 -687
rect 9909 -721 9925 -687
rect 10093 -721 10109 -687
rect 10281 -721 10297 -687
rect 10465 -721 10481 -687
rect 10653 -721 10669 -687
rect 10837 -721 10853 -687
rect 11025 -721 11041 -687
rect 11209 -721 11225 -687
rect -667 -789 -633 -727
rect 11351 -789 11385 -727
rect -667 -823 -571 -789
rect 11289 -823 11385 -789
rect 821 -1207 906 -1173
rect 3849 -1207 3945 -1173
rect 821 -1269 855 -1207
rect 3911 -1269 3945 -1207
rect 981 -1309 997 -1275
rect 1165 -1309 1181 -1275
rect 1353 -1309 1369 -1275
rect 1537 -1309 1553 -1275
rect 1725 -1309 1741 -1275
rect 1909 -1309 1925 -1275
rect 2097 -1309 2113 -1275
rect 2281 -1309 2297 -1275
rect 2469 -1309 2485 -1275
rect 2653 -1309 2669 -1275
rect 2841 -1309 2857 -1275
rect 3025 -1309 3041 -1275
rect 3213 -1309 3229 -1275
rect 3397 -1309 3413 -1275
rect 3585 -1309 3601 -1275
rect 3769 -1309 3785 -1275
rect 935 -1368 969 -1352
rect 935 -2160 969 -2144
rect 1193 -1368 1227 -1352
rect 1193 -2160 1227 -2144
rect 1307 -1368 1341 -1352
rect 1307 -2160 1341 -2144
rect 1565 -1368 1599 -1352
rect 1565 -2160 1599 -2144
rect 1679 -1368 1713 -1352
rect 1679 -2160 1713 -2144
rect 1937 -1368 1971 -1352
rect 1937 -2160 1971 -2144
rect 2051 -1368 2085 -1352
rect 2051 -2160 2085 -2144
rect 2309 -1368 2343 -1352
rect 2309 -2160 2343 -2144
rect 2423 -1368 2457 -1352
rect 2423 -2160 2457 -2144
rect 2681 -1368 2715 -1352
rect 2681 -2160 2715 -2144
rect 2795 -1368 2829 -1352
rect 2795 -2160 2829 -2144
rect 3053 -1368 3087 -1352
rect 3053 -2160 3087 -2144
rect 3167 -1368 3201 -1352
rect 3167 -2160 3201 -2144
rect 3425 -1368 3459 -1352
rect 3425 -2160 3459 -2144
rect 3539 -1368 3573 -1352
rect 3539 -2160 3573 -2144
rect 3797 -1368 3831 -1352
rect 3797 -2160 3831 -2144
rect 981 -2237 997 -2203
rect 1165 -2237 1181 -2203
rect 1353 -2237 1369 -2203
rect 1537 -2237 1553 -2203
rect 1725 -2237 1741 -2203
rect 1909 -2237 1925 -2203
rect 2097 -2237 2113 -2203
rect 2281 -2237 2297 -2203
rect 2469 -2237 2485 -2203
rect 2653 -2237 2669 -2203
rect 2841 -2237 2857 -2203
rect 3025 -2237 3041 -2203
rect 3213 -2237 3229 -2203
rect 3397 -2237 3413 -2203
rect 3585 -2237 3601 -2203
rect 3769 -2237 3785 -2203
rect 981 -2345 997 -2311
rect 1165 -2345 1181 -2311
rect 1353 -2345 1369 -2311
rect 1537 -2345 1553 -2311
rect 1725 -2345 1741 -2311
rect 1909 -2345 1925 -2311
rect 2097 -2345 2113 -2311
rect 2281 -2345 2297 -2311
rect 2469 -2345 2485 -2311
rect 2653 -2345 2669 -2311
rect 2841 -2345 2857 -2311
rect 3025 -2345 3041 -2311
rect 3213 -2345 3229 -2311
rect 3397 -2345 3413 -2311
rect 3585 -2345 3601 -2311
rect 3769 -2345 3785 -2311
rect 935 -2404 969 -2388
rect 935 -3196 969 -3180
rect 1193 -2404 1227 -2388
rect 1193 -3196 1227 -3180
rect 1307 -2404 1341 -2388
rect 1307 -3196 1341 -3180
rect 1565 -2404 1599 -2388
rect 1565 -3196 1599 -3180
rect 1679 -2404 1713 -2388
rect 1679 -3196 1713 -3180
rect 1937 -2404 1971 -2388
rect 1937 -3196 1971 -3180
rect 2051 -2404 2085 -2388
rect 2051 -3196 2085 -3180
rect 2309 -2404 2343 -2388
rect 2309 -3196 2343 -3180
rect 2423 -2404 2457 -2388
rect 2423 -3196 2457 -3180
rect 2681 -2404 2715 -2388
rect 2681 -3196 2715 -3180
rect 2795 -2404 2829 -2388
rect 2795 -3196 2829 -3180
rect 3053 -2404 3087 -2388
rect 3053 -3196 3087 -3180
rect 3167 -2404 3201 -2388
rect 3167 -3196 3201 -3180
rect 3425 -2404 3459 -2388
rect 3425 -3196 3459 -3180
rect 3539 -2404 3573 -2388
rect 3539 -3196 3573 -3180
rect 3797 -2404 3831 -2388
rect 3797 -3196 3831 -3180
rect 981 -3273 997 -3239
rect 1165 -3273 1181 -3239
rect 1353 -3273 1369 -3239
rect 1537 -3273 1553 -3239
rect 1725 -3273 1741 -3239
rect 1909 -3273 1925 -3239
rect 2097 -3273 2113 -3239
rect 2281 -3273 2297 -3239
rect 2469 -3273 2485 -3239
rect 2653 -3273 2669 -3239
rect 2841 -3273 2857 -3239
rect 3025 -3273 3041 -3239
rect 3213 -3273 3229 -3239
rect 3397 -3273 3413 -3239
rect 3585 -3273 3601 -3239
rect 3769 -3273 3785 -3239
rect 981 -3381 997 -3347
rect 1165 -3381 1181 -3347
rect 1353 -3381 1369 -3347
rect 1537 -3381 1553 -3347
rect 1725 -3381 1741 -3347
rect 1909 -3381 1925 -3347
rect 2097 -3381 2113 -3347
rect 2281 -3381 2297 -3347
rect 2469 -3381 2485 -3347
rect 2653 -3381 2669 -3347
rect 2841 -3381 2857 -3347
rect 3025 -3381 3041 -3347
rect 3213 -3381 3229 -3347
rect 3397 -3381 3413 -3347
rect 3585 -3381 3601 -3347
rect 3769 -3381 3785 -3347
rect 935 -3440 969 -3424
rect 935 -4232 969 -4216
rect 1193 -3440 1227 -3424
rect 1193 -4232 1227 -4216
rect 1307 -3440 1341 -3424
rect 1307 -4232 1341 -4216
rect 1565 -3440 1599 -3424
rect 1565 -4232 1599 -4216
rect 1679 -3440 1713 -3424
rect 1679 -4232 1713 -4216
rect 1937 -3440 1971 -3424
rect 1937 -4232 1971 -4216
rect 2051 -3440 2085 -3424
rect 2051 -4232 2085 -4216
rect 2309 -3440 2343 -3424
rect 2309 -4232 2343 -4216
rect 2423 -3440 2457 -3424
rect 2423 -4232 2457 -4216
rect 2681 -3440 2715 -3424
rect 2681 -4232 2715 -4216
rect 2795 -3440 2829 -3424
rect 2795 -4232 2829 -4216
rect 3053 -3440 3087 -3424
rect 3053 -4232 3087 -4216
rect 3167 -3440 3201 -3424
rect 3167 -4232 3201 -4216
rect 3425 -3440 3459 -3424
rect 3425 -4232 3459 -4216
rect 3539 -3440 3573 -3424
rect 3539 -4232 3573 -4216
rect 3797 -3440 3831 -3424
rect 3797 -4232 3831 -4216
rect 981 -4309 997 -4275
rect 1165 -4309 1181 -4275
rect 1353 -4309 1369 -4275
rect 1537 -4309 1553 -4275
rect 1725 -4309 1741 -4275
rect 1909 -4309 1925 -4275
rect 2097 -4309 2113 -4275
rect 2281 -4309 2297 -4275
rect 2469 -4309 2485 -4275
rect 2653 -4309 2669 -4275
rect 2841 -4309 2857 -4275
rect 3025 -4309 3041 -4275
rect 3213 -4309 3229 -4275
rect 3397 -4309 3413 -4275
rect 3585 -4309 3601 -4275
rect 3769 -4309 3785 -4275
rect 981 -4417 997 -4383
rect 1165 -4417 1181 -4383
rect 1353 -4417 1369 -4383
rect 1537 -4417 1553 -4383
rect 1725 -4417 1741 -4383
rect 1909 -4417 1925 -4383
rect 2097 -4417 2113 -4383
rect 2281 -4417 2297 -4383
rect 2469 -4417 2485 -4383
rect 2653 -4417 2669 -4383
rect 2841 -4417 2857 -4383
rect 3025 -4417 3041 -4383
rect 3213 -4417 3229 -4383
rect 3397 -4417 3413 -4383
rect 3585 -4417 3601 -4383
rect 3769 -4417 3785 -4383
rect 935 -4476 969 -4460
rect 935 -5268 969 -5252
rect 1193 -4476 1227 -4460
rect 1193 -5268 1227 -5252
rect 1307 -4476 1341 -4460
rect 1307 -5268 1341 -5252
rect 1565 -4476 1599 -4460
rect 1565 -5268 1599 -5252
rect 1679 -4476 1713 -4460
rect 1679 -5268 1713 -5252
rect 1937 -4476 1971 -4460
rect 1937 -5268 1971 -5252
rect 2051 -4476 2085 -4460
rect 2051 -5268 2085 -5252
rect 2309 -4476 2343 -4460
rect 2309 -5268 2343 -5252
rect 2423 -4476 2457 -4460
rect 2423 -5268 2457 -5252
rect 2681 -4476 2715 -4460
rect 2681 -5268 2715 -5252
rect 2795 -4476 2829 -4460
rect 2795 -5268 2829 -5252
rect 3053 -4476 3087 -4460
rect 3053 -5268 3087 -5252
rect 3167 -4476 3201 -4460
rect 3167 -5268 3201 -5252
rect 3425 -4476 3459 -4460
rect 3425 -5268 3459 -5252
rect 3539 -4476 3573 -4460
rect 3539 -5268 3573 -5252
rect 3797 -4476 3831 -4460
rect 3797 -5268 3831 -5252
rect 981 -5345 997 -5311
rect 1165 -5345 1181 -5311
rect 1353 -5345 1369 -5311
rect 1537 -5345 1553 -5311
rect 1725 -5345 1741 -5311
rect 1909 -5345 1925 -5311
rect 2097 -5345 2113 -5311
rect 2281 -5345 2297 -5311
rect 2469 -5345 2485 -5311
rect 2653 -5345 2669 -5311
rect 2841 -5345 2857 -5311
rect 3025 -5345 3041 -5311
rect 3213 -5345 3229 -5311
rect 3397 -5345 3413 -5311
rect 3585 -5345 3601 -5311
rect 3769 -5345 3785 -5311
rect 821 -5413 855 -5351
rect 5985 -3363 6081 -3329
rect 6219 -3363 6315 -3329
rect 5985 -3425 6019 -3363
rect 6281 -3425 6315 -3363
rect 5985 -4519 6019 -4457
rect 6281 -4519 6315 -4457
rect 5985 -4553 6081 -4519
rect 6219 -4553 6315 -4519
rect 3911 -5413 3945 -5351
rect 821 -5447 917 -5413
rect 3849 -5447 3945 -5413
rect 821 -5901 917 -5867
rect 9801 -5901 9897 -5867
rect 821 -5963 855 -5901
rect 9863 -5963 9897 -5901
rect 981 -6003 997 -5969
rect 1165 -6003 1181 -5969
rect 1353 -6003 1369 -5969
rect 1537 -6003 1553 -5969
rect 1725 -6003 1741 -5969
rect 1909 -6003 1925 -5969
rect 2097 -6003 2113 -5969
rect 2281 -6003 2297 -5969
rect 2469 -6003 2485 -5969
rect 2653 -6003 2669 -5969
rect 2841 -6003 2857 -5969
rect 3025 -6003 3041 -5969
rect 3213 -6003 3229 -5969
rect 3397 -6003 3413 -5969
rect 3585 -6003 3601 -5969
rect 3769 -6003 3785 -5969
rect 3957 -6003 3973 -5969
rect 4141 -6003 4157 -5969
rect 4329 -6003 4345 -5969
rect 4513 -6003 4529 -5969
rect 4701 -6003 4717 -5969
rect 4885 -6003 4901 -5969
rect 5073 -6003 5089 -5969
rect 5257 -6003 5273 -5969
rect 5445 -6003 5461 -5969
rect 5629 -6003 5645 -5969
rect 5817 -6003 5833 -5969
rect 6001 -6003 6017 -5969
rect 6189 -6003 6205 -5969
rect 6373 -6003 6389 -5969
rect 6561 -6003 6577 -5969
rect 6745 -6003 6761 -5969
rect 6933 -6003 6949 -5969
rect 7117 -6003 7133 -5969
rect 7305 -6003 7321 -5969
rect 7489 -6003 7505 -5969
rect 7677 -6003 7693 -5969
rect 7861 -6003 7877 -5969
rect 8049 -6003 8065 -5969
rect 8233 -6003 8249 -5969
rect 8421 -6003 8437 -5969
rect 8605 -6003 8621 -5969
rect 8793 -6003 8809 -5969
rect 8977 -6003 8993 -5969
rect 9165 -6003 9181 -5969
rect 9349 -6003 9365 -5969
rect 9537 -6003 9553 -5969
rect 9721 -6003 9737 -5969
rect 935 -6053 969 -6037
rect 935 -6245 969 -6229
rect 1193 -6053 1227 -6037
rect 1193 -6245 1227 -6229
rect 1307 -6053 1341 -6037
rect 1307 -6245 1341 -6229
rect 1565 -6053 1599 -6037
rect 1565 -6245 1599 -6229
rect 1679 -6053 1713 -6037
rect 1679 -6245 1713 -6229
rect 1937 -6053 1971 -6037
rect 1937 -6245 1971 -6229
rect 2051 -6053 2085 -6037
rect 2051 -6245 2085 -6229
rect 2309 -6053 2343 -6037
rect 2309 -6245 2343 -6229
rect 2423 -6053 2457 -6037
rect 2423 -6245 2457 -6229
rect 2681 -6053 2715 -6037
rect 2681 -6245 2715 -6229
rect 2795 -6053 2829 -6037
rect 2795 -6245 2829 -6229
rect 3053 -6053 3087 -6037
rect 3053 -6245 3087 -6229
rect 3167 -6053 3201 -6037
rect 3167 -6245 3201 -6229
rect 3425 -6053 3459 -6037
rect 3425 -6245 3459 -6229
rect 3539 -6053 3573 -6037
rect 3539 -6245 3573 -6229
rect 3797 -6053 3831 -6037
rect 3797 -6245 3831 -6229
rect 3911 -6053 3945 -6037
rect 3911 -6245 3945 -6229
rect 4169 -6053 4203 -6037
rect 4169 -6245 4203 -6229
rect 4283 -6053 4317 -6037
rect 4283 -6245 4317 -6229
rect 4541 -6053 4575 -6037
rect 4541 -6245 4575 -6229
rect 4655 -6053 4689 -6037
rect 4655 -6245 4689 -6229
rect 4913 -6053 4947 -6037
rect 4913 -6245 4947 -6229
rect 5027 -6053 5061 -6037
rect 5027 -6245 5061 -6229
rect 5285 -6053 5319 -6037
rect 5285 -6245 5319 -6229
rect 5399 -6053 5433 -6037
rect 5399 -6245 5433 -6229
rect 5657 -6053 5691 -6037
rect 5657 -6245 5691 -6229
rect 5771 -6053 5805 -6037
rect 5771 -6245 5805 -6229
rect 6029 -6053 6063 -6037
rect 6029 -6245 6063 -6229
rect 6143 -6053 6177 -6037
rect 6143 -6245 6177 -6229
rect 6401 -6053 6435 -6037
rect 6401 -6245 6435 -6229
rect 6515 -6053 6549 -6037
rect 6515 -6245 6549 -6229
rect 6773 -6053 6807 -6037
rect 6773 -6245 6807 -6229
rect 6887 -6053 6921 -6037
rect 6887 -6245 6921 -6229
rect 7145 -6053 7179 -6037
rect 7145 -6245 7179 -6229
rect 7259 -6053 7293 -6037
rect 7259 -6245 7293 -6229
rect 7517 -6053 7551 -6037
rect 7517 -6245 7551 -6229
rect 7631 -6053 7665 -6037
rect 7631 -6245 7665 -6229
rect 7889 -6053 7923 -6037
rect 7889 -6245 7923 -6229
rect 8003 -6053 8037 -6037
rect 8003 -6245 8037 -6229
rect 8261 -6053 8295 -6037
rect 8261 -6245 8295 -6229
rect 8375 -6053 8409 -6037
rect 8375 -6245 8409 -6229
rect 8633 -6053 8667 -6037
rect 8633 -6245 8667 -6229
rect 8747 -6053 8781 -6037
rect 8747 -6245 8781 -6229
rect 9005 -6053 9039 -6037
rect 9005 -6245 9039 -6229
rect 9119 -6053 9153 -6037
rect 9119 -6245 9153 -6229
rect 9377 -6053 9411 -6037
rect 9377 -6245 9411 -6229
rect 9491 -6053 9525 -6037
rect 9491 -6245 9525 -6229
rect 9749 -6053 9783 -6037
rect 9749 -6245 9783 -6229
rect 981 -6313 997 -6279
rect 1165 -6313 1181 -6279
rect 1353 -6313 1369 -6279
rect 1537 -6313 1553 -6279
rect 1725 -6313 1741 -6279
rect 1909 -6313 1925 -6279
rect 2097 -6313 2113 -6279
rect 2281 -6313 2297 -6279
rect 2469 -6313 2485 -6279
rect 2653 -6313 2669 -6279
rect 2841 -6313 2857 -6279
rect 3025 -6313 3041 -6279
rect 3213 -6313 3229 -6279
rect 3397 -6313 3413 -6279
rect 3585 -6313 3601 -6279
rect 3769 -6313 3785 -6279
rect 3957 -6313 3973 -6279
rect 4141 -6313 4157 -6279
rect 4329 -6313 4345 -6279
rect 4513 -6313 4529 -6279
rect 4701 -6313 4717 -6279
rect 4885 -6313 4901 -6279
rect 5073 -6313 5089 -6279
rect 5257 -6313 5273 -6279
rect 5445 -6313 5461 -6279
rect 5629 -6313 5645 -6279
rect 5817 -6313 5833 -6279
rect 6001 -6313 6017 -6279
rect 6189 -6313 6205 -6279
rect 6373 -6313 6389 -6279
rect 6561 -6313 6577 -6279
rect 6745 -6313 6761 -6279
rect 6933 -6313 6949 -6279
rect 7117 -6313 7133 -6279
rect 7305 -6313 7321 -6279
rect 7489 -6313 7505 -6279
rect 7677 -6313 7693 -6279
rect 7861 -6313 7877 -6279
rect 8049 -6313 8065 -6279
rect 8233 -6313 8249 -6279
rect 8421 -6313 8437 -6279
rect 8605 -6313 8621 -6279
rect 8793 -6313 8809 -6279
rect 8977 -6313 8993 -6279
rect 9165 -6313 9181 -6279
rect 9349 -6313 9365 -6279
rect 9537 -6313 9553 -6279
rect 9721 -6313 9737 -6279
rect 981 -6421 997 -6387
rect 1165 -6421 1181 -6387
rect 1353 -6421 1369 -6387
rect 1537 -6421 1553 -6387
rect 1725 -6421 1741 -6387
rect 1909 -6421 1925 -6387
rect 2097 -6421 2113 -6387
rect 2281 -6421 2297 -6387
rect 2469 -6421 2485 -6387
rect 2653 -6421 2669 -6387
rect 2841 -6421 2857 -6387
rect 3025 -6421 3041 -6387
rect 3213 -6421 3229 -6387
rect 3397 -6421 3413 -6387
rect 3585 -6421 3601 -6387
rect 3769 -6421 3785 -6387
rect 3957 -6421 3973 -6387
rect 4141 -6421 4157 -6387
rect 4329 -6421 4345 -6387
rect 4513 -6421 4529 -6387
rect 4701 -6421 4717 -6387
rect 4885 -6421 4901 -6387
rect 5073 -6421 5089 -6387
rect 5257 -6421 5273 -6387
rect 5445 -6421 5461 -6387
rect 5629 -6421 5645 -6387
rect 5817 -6421 5833 -6387
rect 6001 -6421 6017 -6387
rect 6189 -6421 6205 -6387
rect 6373 -6421 6389 -6387
rect 6561 -6421 6577 -6387
rect 6745 -6421 6761 -6387
rect 6933 -6421 6949 -6387
rect 7117 -6421 7133 -6387
rect 7305 -6421 7321 -6387
rect 7489 -6421 7505 -6387
rect 7677 -6421 7693 -6387
rect 7861 -6421 7877 -6387
rect 8049 -6421 8065 -6387
rect 8233 -6421 8249 -6387
rect 8421 -6421 8437 -6387
rect 8605 -6421 8621 -6387
rect 8793 -6421 8809 -6387
rect 8977 -6421 8993 -6387
rect 9165 -6421 9181 -6387
rect 9349 -6421 9365 -6387
rect 9537 -6421 9553 -6387
rect 9721 -6421 9737 -6387
rect 935 -6471 969 -6455
rect 935 -6663 969 -6647
rect 1193 -6471 1227 -6455
rect 1193 -6663 1227 -6647
rect 1307 -6471 1341 -6455
rect 1307 -6663 1341 -6647
rect 1565 -6471 1599 -6455
rect 1565 -6663 1599 -6647
rect 1679 -6471 1713 -6455
rect 1679 -6663 1713 -6647
rect 1937 -6471 1971 -6455
rect 1937 -6663 1971 -6647
rect 2051 -6471 2085 -6455
rect 2051 -6663 2085 -6647
rect 2309 -6471 2343 -6455
rect 2309 -6663 2343 -6647
rect 2423 -6471 2457 -6455
rect 2423 -6663 2457 -6647
rect 2681 -6471 2715 -6455
rect 2681 -6663 2715 -6647
rect 2795 -6471 2829 -6455
rect 2795 -6663 2829 -6647
rect 3053 -6471 3087 -6455
rect 3053 -6663 3087 -6647
rect 3167 -6471 3201 -6455
rect 3167 -6663 3201 -6647
rect 3425 -6471 3459 -6455
rect 3425 -6663 3459 -6647
rect 3539 -6471 3573 -6455
rect 3539 -6663 3573 -6647
rect 3797 -6471 3831 -6455
rect 3797 -6663 3831 -6647
rect 3911 -6471 3945 -6455
rect 3911 -6663 3945 -6647
rect 4169 -6471 4203 -6455
rect 4169 -6663 4203 -6647
rect 4283 -6471 4317 -6455
rect 4283 -6663 4317 -6647
rect 4541 -6471 4575 -6455
rect 4541 -6663 4575 -6647
rect 4655 -6471 4689 -6455
rect 4655 -6663 4689 -6647
rect 4913 -6471 4947 -6455
rect 4913 -6663 4947 -6647
rect 5027 -6471 5061 -6455
rect 5027 -6663 5061 -6647
rect 5285 -6471 5319 -6455
rect 5285 -6663 5319 -6647
rect 5399 -6471 5433 -6455
rect 5399 -6663 5433 -6647
rect 5657 -6471 5691 -6455
rect 5657 -6663 5691 -6647
rect 5771 -6471 5805 -6455
rect 5771 -6663 5805 -6647
rect 6029 -6471 6063 -6455
rect 6029 -6663 6063 -6647
rect 6143 -6471 6177 -6455
rect 6143 -6663 6177 -6647
rect 6401 -6471 6435 -6455
rect 6401 -6663 6435 -6647
rect 6515 -6471 6549 -6455
rect 6515 -6663 6549 -6647
rect 6773 -6471 6807 -6455
rect 6773 -6663 6807 -6647
rect 6887 -6471 6921 -6455
rect 6887 -6663 6921 -6647
rect 7145 -6471 7179 -6455
rect 7145 -6663 7179 -6647
rect 7259 -6471 7293 -6455
rect 7259 -6663 7293 -6647
rect 7517 -6471 7551 -6455
rect 7517 -6663 7551 -6647
rect 7631 -6471 7665 -6455
rect 7631 -6663 7665 -6647
rect 7889 -6471 7923 -6455
rect 7889 -6663 7923 -6647
rect 8003 -6471 8037 -6455
rect 8003 -6663 8037 -6647
rect 8261 -6471 8295 -6455
rect 8261 -6663 8295 -6647
rect 8375 -6471 8409 -6455
rect 8375 -6663 8409 -6647
rect 8633 -6471 8667 -6455
rect 8633 -6663 8667 -6647
rect 8747 -6471 8781 -6455
rect 8747 -6663 8781 -6647
rect 9005 -6471 9039 -6455
rect 9005 -6663 9039 -6647
rect 9119 -6471 9153 -6455
rect 9119 -6663 9153 -6647
rect 9377 -6471 9411 -6455
rect 9377 -6663 9411 -6647
rect 9491 -6471 9525 -6455
rect 9491 -6663 9525 -6647
rect 9749 -6471 9783 -6455
rect 9749 -6663 9783 -6647
rect 981 -6731 997 -6697
rect 1165 -6731 1181 -6697
rect 1353 -6731 1369 -6697
rect 1537 -6731 1553 -6697
rect 1725 -6731 1741 -6697
rect 1909 -6731 1925 -6697
rect 2097 -6731 2113 -6697
rect 2281 -6731 2297 -6697
rect 2469 -6731 2485 -6697
rect 2653 -6731 2669 -6697
rect 2841 -6731 2857 -6697
rect 3025 -6731 3041 -6697
rect 3213 -6731 3229 -6697
rect 3397 -6731 3413 -6697
rect 3585 -6731 3601 -6697
rect 3769 -6731 3785 -6697
rect 3957 -6731 3973 -6697
rect 4141 -6731 4157 -6697
rect 4329 -6731 4345 -6697
rect 4513 -6731 4529 -6697
rect 4701 -6731 4717 -6697
rect 4885 -6731 4901 -6697
rect 5073 -6731 5089 -6697
rect 5257 -6731 5273 -6697
rect 5445 -6731 5461 -6697
rect 5629 -6731 5645 -6697
rect 5817 -6731 5833 -6697
rect 6001 -6731 6017 -6697
rect 6189 -6731 6205 -6697
rect 6373 -6731 6389 -6697
rect 6561 -6731 6577 -6697
rect 6745 -6731 6761 -6697
rect 6933 -6731 6949 -6697
rect 7117 -6731 7133 -6697
rect 7305 -6731 7321 -6697
rect 7489 -6731 7505 -6697
rect 7677 -6731 7693 -6697
rect 7861 -6731 7877 -6697
rect 8049 -6731 8065 -6697
rect 8233 -6731 8249 -6697
rect 8421 -6731 8437 -6697
rect 8605 -6731 8621 -6697
rect 8793 -6731 8809 -6697
rect 8977 -6731 8993 -6697
rect 9165 -6731 9181 -6697
rect 9349 -6731 9365 -6697
rect 9537 -6731 9553 -6697
rect 9721 -6731 9737 -6697
rect 981 -6839 997 -6805
rect 1165 -6839 1181 -6805
rect 1353 -6839 1369 -6805
rect 1537 -6839 1553 -6805
rect 1725 -6839 1741 -6805
rect 1909 -6839 1925 -6805
rect 2097 -6839 2113 -6805
rect 2281 -6839 2297 -6805
rect 2469 -6839 2485 -6805
rect 2653 -6839 2669 -6805
rect 2841 -6839 2857 -6805
rect 3025 -6839 3041 -6805
rect 3213 -6839 3229 -6805
rect 3397 -6839 3413 -6805
rect 3585 -6839 3601 -6805
rect 3769 -6839 3785 -6805
rect 3957 -6839 3973 -6805
rect 4141 -6839 4157 -6805
rect 4329 -6839 4345 -6805
rect 4513 -6839 4529 -6805
rect 4701 -6839 4717 -6805
rect 4885 -6839 4901 -6805
rect 5073 -6839 5089 -6805
rect 5257 -6839 5273 -6805
rect 5445 -6839 5461 -6805
rect 5629 -6839 5645 -6805
rect 5817 -6839 5833 -6805
rect 6001 -6839 6017 -6805
rect 6189 -6839 6205 -6805
rect 6373 -6839 6389 -6805
rect 6561 -6839 6577 -6805
rect 6745 -6839 6761 -6805
rect 6933 -6839 6949 -6805
rect 7117 -6839 7133 -6805
rect 7305 -6839 7321 -6805
rect 7489 -6839 7505 -6805
rect 7677 -6839 7693 -6805
rect 7861 -6839 7877 -6805
rect 8049 -6839 8065 -6805
rect 8233 -6839 8249 -6805
rect 8421 -6839 8437 -6805
rect 8605 -6839 8621 -6805
rect 8793 -6839 8809 -6805
rect 8977 -6839 8993 -6805
rect 9165 -6839 9181 -6805
rect 9349 -6839 9365 -6805
rect 9537 -6839 9553 -6805
rect 9721 -6839 9737 -6805
rect 935 -6889 969 -6873
rect 935 -7081 969 -7065
rect 1193 -6889 1227 -6873
rect 1193 -7081 1227 -7065
rect 1307 -6889 1341 -6873
rect 1307 -7081 1341 -7065
rect 1565 -6889 1599 -6873
rect 1565 -7081 1599 -7065
rect 1679 -6889 1713 -6873
rect 1679 -7081 1713 -7065
rect 1937 -6889 1971 -6873
rect 1937 -7081 1971 -7065
rect 2051 -6889 2085 -6873
rect 2051 -7081 2085 -7065
rect 2309 -6889 2343 -6873
rect 2309 -7081 2343 -7065
rect 2423 -6889 2457 -6873
rect 2423 -7081 2457 -7065
rect 2681 -6889 2715 -6873
rect 2681 -7081 2715 -7065
rect 2795 -6889 2829 -6873
rect 2795 -7081 2829 -7065
rect 3053 -6889 3087 -6873
rect 3053 -7081 3087 -7065
rect 3167 -6889 3201 -6873
rect 3167 -7081 3201 -7065
rect 3425 -6889 3459 -6873
rect 3425 -7081 3459 -7065
rect 3539 -6889 3573 -6873
rect 3539 -7081 3573 -7065
rect 3797 -6889 3831 -6873
rect 3797 -7081 3831 -7065
rect 3911 -6889 3945 -6873
rect 3911 -7081 3945 -7065
rect 4169 -6889 4203 -6873
rect 4169 -7081 4203 -7065
rect 4283 -6889 4317 -6873
rect 4283 -7081 4317 -7065
rect 4541 -6889 4575 -6873
rect 4541 -7081 4575 -7065
rect 4655 -6889 4689 -6873
rect 4655 -7081 4689 -7065
rect 4913 -6889 4947 -6873
rect 4913 -7081 4947 -7065
rect 5027 -6889 5061 -6873
rect 5027 -7081 5061 -7065
rect 5285 -6889 5319 -6873
rect 5285 -7081 5319 -7065
rect 5399 -6889 5433 -6873
rect 5399 -7081 5433 -7065
rect 5657 -6889 5691 -6873
rect 5657 -7081 5691 -7065
rect 5771 -6889 5805 -6873
rect 5771 -7081 5805 -7065
rect 6029 -6889 6063 -6873
rect 6029 -7081 6063 -7065
rect 6143 -6889 6177 -6873
rect 6143 -7081 6177 -7065
rect 6401 -6889 6435 -6873
rect 6401 -7081 6435 -7065
rect 6515 -6889 6549 -6873
rect 6515 -7081 6549 -7065
rect 6773 -6889 6807 -6873
rect 6773 -7081 6807 -7065
rect 6887 -6889 6921 -6873
rect 6887 -7081 6921 -7065
rect 7145 -6889 7179 -6873
rect 7145 -7081 7179 -7065
rect 7259 -6889 7293 -6873
rect 7259 -7081 7293 -7065
rect 7517 -6889 7551 -6873
rect 7517 -7081 7551 -7065
rect 7631 -6889 7665 -6873
rect 7631 -7081 7665 -7065
rect 7889 -6889 7923 -6873
rect 7889 -7081 7923 -7065
rect 8003 -6889 8037 -6873
rect 8003 -7081 8037 -7065
rect 8261 -6889 8295 -6873
rect 8261 -7081 8295 -7065
rect 8375 -6889 8409 -6873
rect 8375 -7081 8409 -7065
rect 8633 -6889 8667 -6873
rect 8633 -7081 8667 -7065
rect 8747 -6889 8781 -6873
rect 8747 -7081 8781 -7065
rect 9005 -6889 9039 -6873
rect 9005 -7081 9039 -7065
rect 9119 -6889 9153 -6873
rect 9119 -7081 9153 -7065
rect 9377 -6889 9411 -6873
rect 9377 -7081 9411 -7065
rect 9491 -6889 9525 -6873
rect 9491 -7081 9525 -7065
rect 9749 -6889 9783 -6873
rect 9749 -7081 9783 -7065
rect 981 -7149 997 -7115
rect 1165 -7149 1181 -7115
rect 1353 -7149 1369 -7115
rect 1537 -7149 1553 -7115
rect 1725 -7149 1741 -7115
rect 1909 -7149 1925 -7115
rect 2097 -7149 2113 -7115
rect 2281 -7149 2297 -7115
rect 2469 -7149 2485 -7115
rect 2653 -7149 2669 -7115
rect 2841 -7149 2857 -7115
rect 3025 -7149 3041 -7115
rect 3213 -7149 3229 -7115
rect 3397 -7149 3413 -7115
rect 3585 -7149 3601 -7115
rect 3769 -7149 3785 -7115
rect 3957 -7149 3973 -7115
rect 4141 -7149 4157 -7115
rect 4329 -7149 4345 -7115
rect 4513 -7149 4529 -7115
rect 4701 -7149 4717 -7115
rect 4885 -7149 4901 -7115
rect 5073 -7149 5089 -7115
rect 5257 -7149 5273 -7115
rect 5445 -7149 5461 -7115
rect 5629 -7149 5645 -7115
rect 5817 -7149 5833 -7115
rect 6001 -7149 6017 -7115
rect 6189 -7149 6205 -7115
rect 6373 -7149 6389 -7115
rect 6561 -7149 6577 -7115
rect 6745 -7149 6761 -7115
rect 6933 -7149 6949 -7115
rect 7117 -7149 7133 -7115
rect 7305 -7149 7321 -7115
rect 7489 -7149 7505 -7115
rect 7677 -7149 7693 -7115
rect 7861 -7149 7877 -7115
rect 8049 -7149 8065 -7115
rect 8233 -7149 8249 -7115
rect 8421 -7149 8437 -7115
rect 8605 -7149 8621 -7115
rect 8793 -7149 8809 -7115
rect 8977 -7149 8993 -7115
rect 9165 -7149 9181 -7115
rect 9349 -7149 9365 -7115
rect 9537 -7149 9553 -7115
rect 9721 -7149 9737 -7115
rect 981 -7257 997 -7223
rect 1165 -7257 1181 -7223
rect 1353 -7257 1369 -7223
rect 1537 -7257 1553 -7223
rect 1725 -7257 1741 -7223
rect 1909 -7257 1925 -7223
rect 2097 -7257 2113 -7223
rect 2281 -7257 2297 -7223
rect 2469 -7257 2485 -7223
rect 2653 -7257 2669 -7223
rect 2841 -7257 2857 -7223
rect 3025 -7257 3041 -7223
rect 3213 -7257 3229 -7223
rect 3397 -7257 3413 -7223
rect 3585 -7257 3601 -7223
rect 3769 -7257 3785 -7223
rect 3957 -7257 3973 -7223
rect 4141 -7257 4157 -7223
rect 4329 -7257 4345 -7223
rect 4513 -7257 4529 -7223
rect 4701 -7257 4717 -7223
rect 4885 -7257 4901 -7223
rect 5073 -7257 5089 -7223
rect 5257 -7257 5273 -7223
rect 5445 -7257 5461 -7223
rect 5629 -7257 5645 -7223
rect 5817 -7257 5833 -7223
rect 6001 -7257 6017 -7223
rect 6189 -7257 6205 -7223
rect 6373 -7257 6389 -7223
rect 6561 -7257 6577 -7223
rect 6745 -7257 6761 -7223
rect 6933 -7257 6949 -7223
rect 7117 -7257 7133 -7223
rect 7305 -7257 7321 -7223
rect 7489 -7257 7505 -7223
rect 7677 -7257 7693 -7223
rect 7861 -7257 7877 -7223
rect 8049 -7257 8065 -7223
rect 8233 -7257 8249 -7223
rect 8421 -7257 8437 -7223
rect 8605 -7257 8621 -7223
rect 8793 -7257 8809 -7223
rect 8977 -7257 8993 -7223
rect 9165 -7257 9181 -7223
rect 9349 -7257 9365 -7223
rect 9537 -7257 9553 -7223
rect 9721 -7257 9737 -7223
rect 935 -7307 969 -7291
rect 935 -7499 969 -7483
rect 1193 -7307 1227 -7291
rect 1193 -7499 1227 -7483
rect 1307 -7307 1341 -7291
rect 1307 -7499 1341 -7483
rect 1565 -7307 1599 -7291
rect 1565 -7499 1599 -7483
rect 1679 -7307 1713 -7291
rect 1679 -7499 1713 -7483
rect 1937 -7307 1971 -7291
rect 1937 -7499 1971 -7483
rect 2051 -7307 2085 -7291
rect 2051 -7499 2085 -7483
rect 2309 -7307 2343 -7291
rect 2309 -7499 2343 -7483
rect 2423 -7307 2457 -7291
rect 2423 -7499 2457 -7483
rect 2681 -7307 2715 -7291
rect 2681 -7499 2715 -7483
rect 2795 -7307 2829 -7291
rect 2795 -7499 2829 -7483
rect 3053 -7307 3087 -7291
rect 3053 -7499 3087 -7483
rect 3167 -7307 3201 -7291
rect 3167 -7499 3201 -7483
rect 3425 -7307 3459 -7291
rect 3425 -7499 3459 -7483
rect 3539 -7307 3573 -7291
rect 3539 -7499 3573 -7483
rect 3797 -7307 3831 -7291
rect 3797 -7499 3831 -7483
rect 3911 -7307 3945 -7291
rect 3911 -7499 3945 -7483
rect 4169 -7307 4203 -7291
rect 4169 -7499 4203 -7483
rect 4283 -7307 4317 -7291
rect 4283 -7499 4317 -7483
rect 4541 -7307 4575 -7291
rect 4541 -7499 4575 -7483
rect 4655 -7307 4689 -7291
rect 4655 -7499 4689 -7483
rect 4913 -7307 4947 -7291
rect 4913 -7499 4947 -7483
rect 5027 -7307 5061 -7291
rect 5027 -7499 5061 -7483
rect 5285 -7307 5319 -7291
rect 5285 -7499 5319 -7483
rect 5399 -7307 5433 -7291
rect 5399 -7499 5433 -7483
rect 5657 -7307 5691 -7291
rect 5657 -7499 5691 -7483
rect 5771 -7307 5805 -7291
rect 5771 -7499 5805 -7483
rect 6029 -7307 6063 -7291
rect 6029 -7499 6063 -7483
rect 6143 -7307 6177 -7291
rect 6143 -7499 6177 -7483
rect 6401 -7307 6435 -7291
rect 6401 -7499 6435 -7483
rect 6515 -7307 6549 -7291
rect 6515 -7499 6549 -7483
rect 6773 -7307 6807 -7291
rect 6773 -7499 6807 -7483
rect 6887 -7307 6921 -7291
rect 6887 -7499 6921 -7483
rect 7145 -7307 7179 -7291
rect 7145 -7499 7179 -7483
rect 7259 -7307 7293 -7291
rect 7259 -7499 7293 -7483
rect 7517 -7307 7551 -7291
rect 7517 -7499 7551 -7483
rect 7631 -7307 7665 -7291
rect 7631 -7499 7665 -7483
rect 7889 -7307 7923 -7291
rect 7889 -7499 7923 -7483
rect 8003 -7307 8037 -7291
rect 8003 -7499 8037 -7483
rect 8261 -7307 8295 -7291
rect 8261 -7499 8295 -7483
rect 8375 -7307 8409 -7291
rect 8375 -7499 8409 -7483
rect 8633 -7307 8667 -7291
rect 8633 -7499 8667 -7483
rect 8747 -7307 8781 -7291
rect 8747 -7499 8781 -7483
rect 9005 -7307 9039 -7291
rect 9005 -7499 9039 -7483
rect 9119 -7307 9153 -7291
rect 9119 -7499 9153 -7483
rect 9377 -7307 9411 -7291
rect 9377 -7499 9411 -7483
rect 9491 -7307 9525 -7291
rect 9491 -7499 9525 -7483
rect 9749 -7307 9783 -7291
rect 9749 -7499 9783 -7483
rect 981 -7567 997 -7533
rect 1165 -7567 1181 -7533
rect 1353 -7567 1369 -7533
rect 1537 -7567 1553 -7533
rect 1725 -7567 1741 -7533
rect 1909 -7567 1925 -7533
rect 2097 -7567 2113 -7533
rect 2281 -7567 2297 -7533
rect 2469 -7567 2485 -7533
rect 2653 -7567 2669 -7533
rect 2841 -7567 2857 -7533
rect 3025 -7567 3041 -7533
rect 3213 -7567 3229 -7533
rect 3397 -7567 3413 -7533
rect 3585 -7567 3601 -7533
rect 3769 -7567 3785 -7533
rect 3957 -7567 3973 -7533
rect 4141 -7567 4157 -7533
rect 4329 -7567 4345 -7533
rect 4513 -7567 4529 -7533
rect 4701 -7567 4717 -7533
rect 4885 -7567 4901 -7533
rect 5073 -7567 5089 -7533
rect 5257 -7567 5273 -7533
rect 5445 -7567 5461 -7533
rect 5629 -7567 5645 -7533
rect 5817 -7567 5833 -7533
rect 6001 -7567 6017 -7533
rect 6189 -7567 6205 -7533
rect 6373 -7567 6389 -7533
rect 6561 -7567 6577 -7533
rect 6745 -7567 6761 -7533
rect 6933 -7567 6949 -7533
rect 7117 -7567 7133 -7533
rect 7305 -7567 7321 -7533
rect 7489 -7567 7505 -7533
rect 7677 -7567 7693 -7533
rect 7861 -7567 7877 -7533
rect 8049 -7567 8065 -7533
rect 8233 -7567 8249 -7533
rect 8421 -7567 8437 -7533
rect 8605 -7567 8621 -7533
rect 8793 -7567 8809 -7533
rect 8977 -7567 8993 -7533
rect 9165 -7567 9181 -7533
rect 9349 -7567 9365 -7533
rect 9537 -7567 9553 -7533
rect 9721 -7567 9737 -7533
rect 821 -7635 855 -7573
rect 9863 -7635 9897 -7573
rect 821 -7669 917 -7635
rect 9801 -7669 9897 -7635
<< viali >>
rect -256 1215 -186 1232
rect 488 1215 558 1232
rect 1232 1215 1302 1232
rect 1976 1215 2046 1232
rect 2720 1215 2790 1232
rect 3464 1215 3534 1232
rect 4208 1215 4278 1232
rect 4952 1215 5022 1232
rect 5324 1215 5394 1232
rect 6068 1215 6138 1232
rect 6812 1215 6882 1232
rect 7556 1215 7626 1232
rect 8300 1215 8370 1232
rect 9044 1215 9114 1232
rect 9788 1215 9858 1232
rect 10532 1215 10602 1232
rect 11222 1215 11292 1232
rect -256 1181 -186 1215
rect 488 1181 558 1215
rect 1232 1181 1302 1215
rect 1976 1181 2046 1215
rect 2720 1181 2790 1215
rect 3464 1181 3534 1215
rect 4208 1181 4278 1215
rect 4952 1181 5022 1215
rect 5324 1181 5394 1215
rect 6068 1181 6138 1215
rect 6812 1181 6882 1215
rect 7556 1181 7626 1215
rect 8300 1181 8370 1215
rect 9044 1181 9114 1215
rect 9788 1181 9858 1215
rect 10532 1181 10602 1215
rect 11222 1181 11289 1215
rect 11289 1181 11292 1215
rect -256 1162 -186 1181
rect 488 1162 558 1181
rect 1232 1162 1302 1181
rect 1976 1162 2046 1181
rect 2720 1162 2790 1181
rect 3464 1162 3534 1181
rect 4208 1162 4278 1181
rect 4952 1162 5022 1181
rect 5324 1162 5394 1181
rect 6068 1162 6138 1181
rect 6812 1162 6882 1181
rect 7556 1162 7626 1181
rect 8300 1162 8370 1181
rect 9044 1162 9114 1181
rect 9788 1162 9858 1181
rect 10532 1162 10602 1181
rect 11222 1162 11292 1181
rect -491 1079 -323 1113
rect -119 1079 49 1113
rect 253 1079 421 1113
rect 625 1079 793 1113
rect 997 1079 1165 1113
rect 1369 1079 1537 1113
rect 1741 1079 1909 1113
rect 2113 1079 2281 1113
rect 2485 1079 2653 1113
rect 2857 1079 3025 1113
rect 3229 1079 3397 1113
rect 3601 1079 3769 1113
rect 3973 1079 4141 1113
rect 4345 1079 4513 1113
rect 4717 1079 4885 1113
rect 5089 1079 5257 1113
rect 5461 1079 5629 1113
rect 5833 1079 6001 1113
rect 6205 1079 6373 1113
rect 6577 1079 6745 1113
rect 6949 1079 7117 1113
rect 7321 1079 7489 1113
rect 7693 1079 7861 1113
rect 8065 1079 8233 1113
rect 8437 1079 8605 1113
rect 8809 1079 8977 1113
rect 9181 1079 9349 1113
rect 9553 1079 9721 1113
rect 9925 1079 10093 1113
rect 10297 1079 10465 1113
rect 10669 1079 10837 1113
rect 11041 1079 11209 1113
rect -553 644 -519 1020
rect -295 644 -261 1020
rect -181 644 -147 1020
rect 77 644 111 1020
rect 191 644 225 1020
rect 449 644 483 1020
rect 563 644 597 1020
rect 821 644 855 1020
rect 935 644 969 1020
rect 1193 644 1227 1020
rect 1307 644 1341 1020
rect 1565 644 1599 1020
rect 1679 644 1713 1020
rect 1937 644 1971 1020
rect 2051 644 2085 1020
rect 2309 644 2343 1020
rect 2423 644 2457 1020
rect 2681 644 2715 1020
rect 2795 644 2829 1020
rect 3053 644 3087 1020
rect 3167 644 3201 1020
rect 3425 644 3459 1020
rect 3539 644 3573 1020
rect 3797 644 3831 1020
rect 3911 644 3945 1020
rect 4169 644 4203 1020
rect 4283 644 4317 1020
rect 4541 644 4575 1020
rect 4655 644 4689 1020
rect 4913 644 4947 1020
rect 5027 644 5061 1020
rect 5285 644 5319 1020
rect 5399 644 5433 1020
rect 5657 644 5691 1020
rect 5771 644 5805 1020
rect 6029 644 6063 1020
rect 6143 644 6177 1020
rect 6401 644 6435 1020
rect 6515 644 6549 1020
rect 6773 644 6807 1020
rect 6887 644 6921 1020
rect 7145 644 7179 1020
rect 7259 644 7293 1020
rect 7517 644 7551 1020
rect 7631 644 7665 1020
rect 7889 644 7923 1020
rect 8003 644 8037 1020
rect 8261 644 8295 1020
rect 8375 644 8409 1020
rect 8633 644 8667 1020
rect 8747 644 8781 1020
rect 9005 644 9039 1020
rect 9119 644 9153 1020
rect 9377 644 9411 1020
rect 9491 644 9525 1020
rect 9749 644 9783 1020
rect 9863 644 9897 1020
rect 10121 644 10155 1020
rect 10235 644 10269 1020
rect 10493 644 10527 1020
rect 10607 644 10641 1020
rect 10865 644 10899 1020
rect 10979 644 11013 1020
rect 11237 644 11271 1020
rect -491 551 -323 585
rect -119 551 49 585
rect 253 551 421 585
rect 625 551 793 585
rect 997 551 1165 585
rect 1369 551 1537 585
rect 1741 551 1909 585
rect 2113 551 2281 585
rect 2485 551 2653 585
rect 2857 551 3025 585
rect 3229 551 3397 585
rect 3601 551 3769 585
rect 3973 551 4141 585
rect 4345 551 4513 585
rect 4717 551 4885 585
rect 5089 551 5257 585
rect 5461 551 5629 585
rect 5833 551 6001 585
rect 6205 551 6373 585
rect 6577 551 6745 585
rect 6949 551 7117 585
rect 7321 551 7489 585
rect 7693 551 7861 585
rect 8065 551 8233 585
rect 8437 551 8605 585
rect 8809 551 8977 585
rect 9181 551 9349 585
rect 9553 551 9721 585
rect 9925 551 10093 585
rect 10297 551 10465 585
rect 10669 551 10837 585
rect 11041 551 11209 585
rect -491 443 -323 477
rect -119 443 49 477
rect 253 443 421 477
rect 625 443 793 477
rect 997 443 1165 477
rect 1369 443 1537 477
rect 1741 443 1909 477
rect 2113 443 2281 477
rect 2485 443 2653 477
rect 2857 443 3025 477
rect 3229 443 3397 477
rect 3601 443 3769 477
rect 3973 443 4141 477
rect 4345 443 4513 477
rect 4717 443 4885 477
rect 5089 443 5257 477
rect 5461 443 5629 477
rect 5833 443 6001 477
rect 6205 443 6373 477
rect 6577 443 6745 477
rect 6949 443 7117 477
rect 7321 443 7489 477
rect 7693 443 7861 477
rect 8065 443 8233 477
rect 8437 443 8605 477
rect 8809 443 8977 477
rect 9181 443 9349 477
rect 9553 443 9721 477
rect 9925 443 10093 477
rect 10297 443 10465 477
rect 10669 443 10837 477
rect 11041 443 11209 477
rect -553 8 -519 384
rect -295 8 -261 384
rect -181 8 -147 384
rect 77 8 111 384
rect 191 8 225 384
rect 449 8 483 384
rect 563 8 597 384
rect 821 8 855 384
rect 935 8 969 384
rect 1193 8 1227 384
rect 1307 8 1341 384
rect 1565 8 1599 384
rect 1679 8 1713 384
rect 1937 8 1971 384
rect 2051 8 2085 384
rect 2309 8 2343 384
rect 2423 8 2457 384
rect 2681 8 2715 384
rect 2795 8 2829 384
rect 3053 8 3087 384
rect 3167 8 3201 384
rect 3425 8 3459 384
rect 3539 8 3573 384
rect 3797 8 3831 384
rect 3911 8 3945 384
rect 4169 8 4203 384
rect 4283 8 4317 384
rect 4541 8 4575 384
rect 4655 8 4689 384
rect 4913 8 4947 384
rect 5027 8 5061 384
rect 5285 8 5319 384
rect 5399 8 5433 384
rect 5657 8 5691 384
rect 5771 8 5805 384
rect 6029 8 6063 384
rect 6143 8 6177 384
rect 6401 8 6435 384
rect 6515 8 6549 384
rect 6773 8 6807 384
rect 6887 8 6921 384
rect 7145 8 7179 384
rect 7259 8 7293 384
rect 7517 8 7551 384
rect 7631 8 7665 384
rect 7889 8 7923 384
rect 8003 8 8037 384
rect 8261 8 8295 384
rect 8375 8 8409 384
rect 8633 8 8667 384
rect 8747 8 8781 384
rect 9005 8 9039 384
rect 9119 8 9153 384
rect 9377 8 9411 384
rect 9491 8 9525 384
rect 9749 8 9783 384
rect 9863 8 9897 384
rect 10121 8 10155 384
rect 10235 8 10269 384
rect 10493 8 10527 384
rect 10607 8 10641 384
rect 10865 8 10899 384
rect 10979 8 11013 384
rect 11237 8 11271 384
rect -491 -85 -323 -51
rect -119 -85 49 -51
rect 253 -85 421 -51
rect 625 -85 793 -51
rect 997 -85 1165 -51
rect 1369 -85 1537 -51
rect 1741 -85 1909 -51
rect 2113 -85 2281 -51
rect 2485 -85 2653 -51
rect 2857 -85 3025 -51
rect 3229 -85 3397 -51
rect 3601 -85 3769 -51
rect 3973 -85 4141 -51
rect 4345 -85 4513 -51
rect 4717 -85 4885 -51
rect 5089 -85 5257 -51
rect 5461 -85 5629 -51
rect 5833 -85 6001 -51
rect 6205 -85 6373 -51
rect 6577 -85 6745 -51
rect 6949 -85 7117 -51
rect 7321 -85 7489 -51
rect 7693 -85 7861 -51
rect 8065 -85 8233 -51
rect 8437 -85 8605 -51
rect 8809 -85 8977 -51
rect 9181 -85 9349 -51
rect 9553 -85 9721 -51
rect 9925 -85 10093 -51
rect 10297 -85 10465 -51
rect 10669 -85 10837 -51
rect 11041 -85 11209 -51
rect -491 -193 -323 -159
rect -119 -193 49 -159
rect 253 -193 421 -159
rect 625 -193 793 -159
rect 997 -193 1165 -159
rect 1369 -193 1537 -159
rect 1741 -193 1909 -159
rect 2113 -193 2281 -159
rect 2485 -193 2653 -159
rect 2857 -193 3025 -159
rect 3229 -193 3397 -159
rect 3601 -193 3769 -159
rect 3973 -193 4141 -159
rect 4345 -193 4513 -159
rect 4717 -193 4885 -159
rect 5089 -193 5257 -159
rect 5461 -193 5629 -159
rect 5833 -193 6001 -159
rect 6205 -193 6373 -159
rect 6577 -193 6745 -159
rect 6949 -193 7117 -159
rect 7321 -193 7489 -159
rect 7693 -193 7861 -159
rect 8065 -193 8233 -159
rect 8437 -193 8605 -159
rect 8809 -193 8977 -159
rect 9181 -193 9349 -159
rect 9553 -193 9721 -159
rect 9925 -193 10093 -159
rect 10297 -193 10465 -159
rect 10669 -193 10837 -159
rect 11041 -193 11209 -159
rect -553 -628 -519 -252
rect -295 -628 -261 -252
rect -181 -628 -147 -252
rect 77 -628 111 -252
rect 191 -628 225 -252
rect 449 -628 483 -252
rect 563 -628 597 -252
rect 821 -628 855 -252
rect 935 -628 969 -252
rect 1193 -628 1227 -252
rect 1307 -628 1341 -252
rect 1565 -628 1599 -252
rect 1679 -628 1713 -252
rect 1937 -628 1971 -252
rect 2051 -628 2085 -252
rect 2309 -628 2343 -252
rect 2423 -628 2457 -252
rect 2681 -628 2715 -252
rect 2795 -628 2829 -252
rect 3053 -628 3087 -252
rect 3167 -628 3201 -252
rect 3425 -628 3459 -252
rect 3539 -628 3573 -252
rect 3797 -628 3831 -252
rect 3911 -628 3945 -252
rect 4169 -628 4203 -252
rect 4283 -628 4317 -252
rect 4541 -628 4575 -252
rect 4655 -628 4689 -252
rect 4913 -628 4947 -252
rect 5027 -628 5061 -252
rect 5285 -628 5319 -252
rect 5399 -628 5433 -252
rect 5657 -628 5691 -252
rect 5771 -628 5805 -252
rect 6029 -628 6063 -252
rect 6143 -628 6177 -252
rect 6401 -628 6435 -252
rect 6515 -628 6549 -252
rect 6773 -628 6807 -252
rect 6887 -628 6921 -252
rect 7145 -628 7179 -252
rect 7259 -628 7293 -252
rect 7517 -628 7551 -252
rect 7631 -628 7665 -252
rect 7889 -628 7923 -252
rect 8003 -628 8037 -252
rect 8261 -628 8295 -252
rect 8375 -628 8409 -252
rect 8633 -628 8667 -252
rect 8747 -628 8781 -252
rect 9005 -628 9039 -252
rect 9119 -628 9153 -252
rect 9377 -628 9411 -252
rect 9491 -628 9525 -252
rect 9749 -628 9783 -252
rect 9863 -628 9897 -252
rect 10121 -628 10155 -252
rect 10235 -628 10269 -252
rect 10493 -628 10527 -252
rect 10607 -628 10641 -252
rect 10865 -628 10899 -252
rect 10979 -628 11013 -252
rect 11237 -628 11271 -252
rect -491 -721 -323 -687
rect -119 -721 49 -687
rect 253 -721 421 -687
rect 625 -721 793 -687
rect 997 -721 1165 -687
rect 1369 -721 1537 -687
rect 1741 -721 1909 -687
rect 2113 -721 2281 -687
rect 2485 -721 2653 -687
rect 2857 -721 3025 -687
rect 3229 -721 3397 -687
rect 3601 -721 3769 -687
rect 3973 -721 4141 -687
rect 4345 -721 4513 -687
rect 4717 -721 4885 -687
rect 5089 -721 5257 -687
rect 5461 -721 5629 -687
rect 5833 -721 6001 -687
rect 6205 -721 6373 -687
rect 6577 -721 6745 -687
rect 6949 -721 7117 -687
rect 7321 -721 7489 -687
rect 7693 -721 7861 -687
rect 8065 -721 8233 -687
rect 8437 -721 8605 -687
rect 8809 -721 8977 -687
rect 9181 -721 9349 -687
rect 9553 -721 9721 -687
rect 9925 -721 10093 -687
rect 10297 -721 10465 -687
rect 10669 -721 10837 -687
rect 11041 -721 11209 -687
rect 906 -1173 976 -1156
rect 1278 -1173 1348 -1156
rect 1650 -1173 1720 -1156
rect 2022 -1173 2092 -1156
rect 2394 -1173 2464 -1156
rect 2766 -1173 2836 -1156
rect 3138 -1173 3208 -1156
rect 3510 -1173 3580 -1156
rect 3772 -1173 3842 -1156
rect 906 -1207 917 -1173
rect 917 -1207 976 -1173
rect 1278 -1207 1348 -1173
rect 1650 -1207 1720 -1173
rect 2022 -1207 2092 -1173
rect 2394 -1207 2464 -1173
rect 2766 -1207 2836 -1173
rect 3138 -1207 3208 -1173
rect 3510 -1207 3580 -1173
rect 3772 -1207 3842 -1173
rect 906 -1226 976 -1207
rect 1278 -1226 1348 -1207
rect 1650 -1226 1720 -1207
rect 2022 -1226 2092 -1207
rect 2394 -1226 2464 -1207
rect 2766 -1226 2836 -1207
rect 3138 -1226 3208 -1207
rect 3510 -1226 3580 -1207
rect 3772 -1226 3842 -1207
rect 997 -1309 1165 -1275
rect 1369 -1309 1537 -1275
rect 1741 -1309 1909 -1275
rect 2113 -1309 2281 -1275
rect 2485 -1309 2653 -1275
rect 2857 -1309 3025 -1275
rect 3229 -1309 3397 -1275
rect 3601 -1309 3769 -1275
rect 935 -2144 969 -1368
rect 1193 -2144 1227 -1368
rect 1307 -2144 1341 -1368
rect 1565 -2144 1599 -1368
rect 1679 -2144 1713 -1368
rect 1937 -2144 1971 -1368
rect 2051 -2144 2085 -1368
rect 2309 -2144 2343 -1368
rect 2423 -2144 2457 -1368
rect 2681 -2144 2715 -1368
rect 2795 -2144 2829 -1368
rect 3053 -2144 3087 -1368
rect 3167 -2144 3201 -1368
rect 3425 -2144 3459 -1368
rect 3539 -2144 3573 -1368
rect 3797 -2144 3831 -1368
rect 997 -2237 1165 -2203
rect 1369 -2237 1537 -2203
rect 1741 -2237 1909 -2203
rect 2113 -2237 2281 -2203
rect 2485 -2237 2653 -2203
rect 2857 -2237 3025 -2203
rect 3229 -2237 3397 -2203
rect 3601 -2237 3769 -2203
rect 997 -2345 1165 -2311
rect 1369 -2345 1537 -2311
rect 1741 -2345 1909 -2311
rect 2113 -2345 2281 -2311
rect 2485 -2345 2653 -2311
rect 2857 -2345 3025 -2311
rect 3229 -2345 3397 -2311
rect 3601 -2345 3769 -2311
rect 935 -3180 969 -2404
rect 1193 -3180 1227 -2404
rect 1307 -3180 1341 -2404
rect 1565 -3180 1599 -2404
rect 1679 -3180 1713 -2404
rect 1937 -3180 1971 -2404
rect 2051 -3180 2085 -2404
rect 2309 -3180 2343 -2404
rect 2423 -3180 2457 -2404
rect 2681 -3180 2715 -2404
rect 2795 -3180 2829 -2404
rect 3053 -3180 3087 -2404
rect 3167 -3180 3201 -2404
rect 3425 -3180 3459 -2404
rect 3539 -3180 3573 -2404
rect 3797 -3180 3831 -2404
rect 997 -3273 1165 -3239
rect 1369 -3273 1537 -3239
rect 1741 -3273 1909 -3239
rect 2113 -3273 2281 -3239
rect 2485 -3273 2653 -3239
rect 2857 -3273 3025 -3239
rect 3229 -3273 3397 -3239
rect 3601 -3273 3769 -3239
rect 997 -3381 1165 -3347
rect 1369 -3381 1537 -3347
rect 1741 -3381 1909 -3347
rect 2113 -3381 2281 -3347
rect 2485 -3381 2653 -3347
rect 2857 -3381 3025 -3347
rect 3229 -3381 3397 -3347
rect 3601 -3381 3769 -3347
rect 935 -4216 969 -3440
rect 1193 -4216 1227 -3440
rect 1307 -4216 1341 -3440
rect 1565 -4216 1599 -3440
rect 1679 -4216 1713 -3440
rect 1937 -4216 1971 -3440
rect 2051 -4216 2085 -3440
rect 2309 -4216 2343 -3440
rect 2423 -4216 2457 -3440
rect 2681 -4216 2715 -3440
rect 2795 -4216 2829 -3440
rect 3053 -4216 3087 -3440
rect 3167 -4216 3201 -3440
rect 3425 -4216 3459 -3440
rect 3539 -4216 3573 -3440
rect 3797 -4216 3831 -3440
rect 997 -4309 1165 -4275
rect 1369 -4309 1537 -4275
rect 1741 -4309 1909 -4275
rect 2113 -4309 2281 -4275
rect 2485 -4309 2653 -4275
rect 2857 -4309 3025 -4275
rect 3229 -4309 3397 -4275
rect 3601 -4309 3769 -4275
rect 997 -4417 1165 -4383
rect 1369 -4417 1537 -4383
rect 1741 -4417 1909 -4383
rect 2113 -4417 2281 -4383
rect 2485 -4417 2653 -4383
rect 2857 -4417 3025 -4383
rect 3229 -4417 3397 -4383
rect 3601 -4417 3769 -4383
rect 935 -5252 969 -4476
rect 1193 -5252 1227 -4476
rect 1307 -5252 1341 -4476
rect 1565 -5252 1599 -4476
rect 1679 -5252 1713 -4476
rect 1937 -5252 1971 -4476
rect 2051 -5252 2085 -4476
rect 2309 -5252 2343 -4476
rect 2423 -5252 2457 -4476
rect 2681 -5252 2715 -4476
rect 2795 -5252 2829 -4476
rect 3053 -5252 3087 -4476
rect 3167 -5252 3201 -4476
rect 3425 -5252 3459 -4476
rect 3539 -5252 3573 -4476
rect 3797 -5252 3831 -4476
rect 997 -5345 1165 -5311
rect 1369 -5345 1537 -5311
rect 1741 -5345 1909 -5311
rect 2113 -5345 2281 -5311
rect 2485 -5345 2653 -5311
rect 2857 -5345 3025 -5311
rect 3229 -5345 3397 -5311
rect 3601 -5345 3769 -5311
rect 5974 -3634 5985 -3584
rect 5985 -3634 6019 -3584
rect 6019 -3634 6030 -3584
rect 6131 -3874 6169 -3477
rect 5974 -4034 5985 -3984
rect 5985 -4034 6019 -3984
rect 6019 -4034 6030 -3984
rect 5974 -4434 5985 -4384
rect 5985 -4434 6019 -4384
rect 6019 -4434 6030 -4384
rect 6131 -4405 6169 -4008
rect 997 -6003 1165 -5969
rect 1369 -6003 1537 -5969
rect 1741 -6003 1909 -5969
rect 2113 -6003 2281 -5969
rect 2485 -6003 2653 -5969
rect 2857 -6003 3025 -5969
rect 3229 -6003 3397 -5969
rect 3601 -6003 3769 -5969
rect 3973 -6003 4141 -5969
rect 4345 -6003 4513 -5969
rect 4717 -6003 4885 -5969
rect 5089 -6003 5257 -5969
rect 5461 -6003 5629 -5969
rect 5833 -6003 6001 -5969
rect 6205 -6003 6373 -5969
rect 6577 -6003 6745 -5969
rect 6949 -6003 7117 -5969
rect 7321 -6003 7489 -5969
rect 7693 -6003 7861 -5969
rect 8065 -6003 8233 -5969
rect 8437 -6003 8605 -5969
rect 8809 -6003 8977 -5969
rect 9181 -6003 9349 -5969
rect 9553 -6003 9721 -5969
rect 935 -6229 969 -6053
rect 1193 -6229 1227 -6053
rect 1307 -6229 1341 -6053
rect 1565 -6229 1599 -6053
rect 1679 -6229 1713 -6053
rect 1937 -6229 1971 -6053
rect 2051 -6229 2085 -6053
rect 2309 -6229 2343 -6053
rect 2423 -6229 2457 -6053
rect 2681 -6229 2715 -6053
rect 2795 -6229 2829 -6053
rect 3053 -6229 3087 -6053
rect 3167 -6229 3201 -6053
rect 3425 -6229 3459 -6053
rect 3539 -6229 3573 -6053
rect 3797 -6229 3831 -6053
rect 3911 -6229 3945 -6053
rect 4169 -6229 4203 -6053
rect 4283 -6229 4317 -6053
rect 4541 -6229 4575 -6053
rect 4655 -6229 4689 -6053
rect 4913 -6229 4947 -6053
rect 5027 -6229 5061 -6053
rect 5285 -6229 5319 -6053
rect 5399 -6229 5433 -6053
rect 5657 -6229 5691 -6053
rect 5771 -6229 5805 -6053
rect 6029 -6229 6063 -6053
rect 6143 -6229 6177 -6053
rect 6401 -6229 6435 -6053
rect 6515 -6229 6549 -6053
rect 6773 -6229 6807 -6053
rect 6887 -6229 6921 -6053
rect 7145 -6229 7179 -6053
rect 7259 -6229 7293 -6053
rect 7517 -6229 7551 -6053
rect 7631 -6229 7665 -6053
rect 7889 -6229 7923 -6053
rect 8003 -6229 8037 -6053
rect 8261 -6229 8295 -6053
rect 8375 -6229 8409 -6053
rect 8633 -6229 8667 -6053
rect 8747 -6229 8781 -6053
rect 9005 -6229 9039 -6053
rect 9119 -6229 9153 -6053
rect 9377 -6229 9411 -6053
rect 9491 -6229 9525 -6053
rect 9749 -6229 9783 -6053
rect 997 -6313 1165 -6279
rect 1369 -6313 1537 -6279
rect 1741 -6313 1909 -6279
rect 2113 -6313 2281 -6279
rect 2485 -6313 2653 -6279
rect 2857 -6313 3025 -6279
rect 3229 -6313 3397 -6279
rect 3601 -6313 3769 -6279
rect 3973 -6313 4141 -6279
rect 4345 -6313 4513 -6279
rect 4717 -6313 4885 -6279
rect 5089 -6313 5257 -6279
rect 5461 -6313 5629 -6279
rect 5833 -6313 6001 -6279
rect 6205 -6313 6373 -6279
rect 6577 -6313 6745 -6279
rect 6949 -6313 7117 -6279
rect 7321 -6313 7489 -6279
rect 7693 -6313 7861 -6279
rect 8065 -6313 8233 -6279
rect 8437 -6313 8605 -6279
rect 8809 -6313 8977 -6279
rect 9181 -6313 9349 -6279
rect 9553 -6313 9721 -6279
rect 997 -6421 1165 -6387
rect 1369 -6421 1537 -6387
rect 1741 -6421 1909 -6387
rect 2113 -6421 2281 -6387
rect 2485 -6421 2653 -6387
rect 2857 -6421 3025 -6387
rect 3229 -6421 3397 -6387
rect 3601 -6421 3769 -6387
rect 3973 -6421 4141 -6387
rect 4345 -6421 4513 -6387
rect 4717 -6421 4885 -6387
rect 5089 -6421 5257 -6387
rect 5461 -6421 5629 -6387
rect 5833 -6421 6001 -6387
rect 6205 -6421 6373 -6387
rect 6577 -6421 6745 -6387
rect 6949 -6421 7117 -6387
rect 7321 -6421 7489 -6387
rect 7693 -6421 7861 -6387
rect 8065 -6421 8233 -6387
rect 8437 -6421 8605 -6387
rect 8809 -6421 8977 -6387
rect 9181 -6421 9349 -6387
rect 9553 -6421 9721 -6387
rect 935 -6647 969 -6471
rect 1193 -6647 1227 -6471
rect 1307 -6647 1341 -6471
rect 1565 -6647 1599 -6471
rect 1679 -6647 1713 -6471
rect 1937 -6647 1971 -6471
rect 2051 -6647 2085 -6471
rect 2309 -6647 2343 -6471
rect 2423 -6647 2457 -6471
rect 2681 -6647 2715 -6471
rect 2795 -6647 2829 -6471
rect 3053 -6647 3087 -6471
rect 3167 -6647 3201 -6471
rect 3425 -6647 3459 -6471
rect 3539 -6647 3573 -6471
rect 3797 -6647 3831 -6471
rect 3911 -6647 3945 -6471
rect 4169 -6647 4203 -6471
rect 4283 -6647 4317 -6471
rect 4541 -6647 4575 -6471
rect 4655 -6647 4689 -6471
rect 4913 -6647 4947 -6471
rect 5027 -6647 5061 -6471
rect 5285 -6647 5319 -6471
rect 5399 -6647 5433 -6471
rect 5657 -6647 5691 -6471
rect 5771 -6647 5805 -6471
rect 6029 -6647 6063 -6471
rect 6143 -6647 6177 -6471
rect 6401 -6647 6435 -6471
rect 6515 -6647 6549 -6471
rect 6773 -6647 6807 -6471
rect 6887 -6647 6921 -6471
rect 7145 -6647 7179 -6471
rect 7259 -6647 7293 -6471
rect 7517 -6647 7551 -6471
rect 7631 -6647 7665 -6471
rect 7889 -6647 7923 -6471
rect 8003 -6647 8037 -6471
rect 8261 -6647 8295 -6471
rect 8375 -6647 8409 -6471
rect 8633 -6647 8667 -6471
rect 8747 -6647 8781 -6471
rect 9005 -6647 9039 -6471
rect 9119 -6647 9153 -6471
rect 9377 -6647 9411 -6471
rect 9491 -6647 9525 -6471
rect 9749 -6647 9783 -6471
rect 997 -6731 1165 -6697
rect 1369 -6731 1537 -6697
rect 1741 -6731 1909 -6697
rect 2113 -6731 2281 -6697
rect 2485 -6731 2653 -6697
rect 2857 -6731 3025 -6697
rect 3229 -6731 3397 -6697
rect 3601 -6731 3769 -6697
rect 3973 -6731 4141 -6697
rect 4345 -6731 4513 -6697
rect 4717 -6731 4885 -6697
rect 5089 -6731 5257 -6697
rect 5461 -6731 5629 -6697
rect 5833 -6731 6001 -6697
rect 6205 -6731 6373 -6697
rect 6577 -6731 6745 -6697
rect 6949 -6731 7117 -6697
rect 7321 -6731 7489 -6697
rect 7693 -6731 7861 -6697
rect 8065 -6731 8233 -6697
rect 8437 -6731 8605 -6697
rect 8809 -6731 8977 -6697
rect 9181 -6731 9349 -6697
rect 9553 -6731 9721 -6697
rect 997 -6839 1165 -6805
rect 1369 -6839 1537 -6805
rect 1741 -6839 1909 -6805
rect 2113 -6839 2281 -6805
rect 2485 -6839 2653 -6805
rect 2857 -6839 3025 -6805
rect 3229 -6839 3397 -6805
rect 3601 -6839 3769 -6805
rect 3973 -6839 4141 -6805
rect 4345 -6839 4513 -6805
rect 4717 -6839 4885 -6805
rect 5089 -6839 5257 -6805
rect 5461 -6839 5629 -6805
rect 5833 -6839 6001 -6805
rect 6205 -6839 6373 -6805
rect 6577 -6839 6745 -6805
rect 6949 -6839 7117 -6805
rect 7321 -6839 7489 -6805
rect 7693 -6839 7861 -6805
rect 8065 -6839 8233 -6805
rect 8437 -6839 8605 -6805
rect 8809 -6839 8977 -6805
rect 9181 -6839 9349 -6805
rect 9553 -6839 9721 -6805
rect 935 -7065 969 -6889
rect 1193 -7065 1227 -6889
rect 1307 -7065 1341 -6889
rect 1565 -7065 1599 -6889
rect 1679 -7065 1713 -6889
rect 1937 -7065 1971 -6889
rect 2051 -7065 2085 -6889
rect 2309 -7065 2343 -6889
rect 2423 -7065 2457 -6889
rect 2681 -7065 2715 -6889
rect 2795 -7065 2829 -6889
rect 3053 -7065 3087 -6889
rect 3167 -7065 3201 -6889
rect 3425 -7065 3459 -6889
rect 3539 -7065 3573 -6889
rect 3797 -7065 3831 -6889
rect 3911 -7065 3945 -6889
rect 4169 -7065 4203 -6889
rect 4283 -7065 4317 -6889
rect 4541 -7065 4575 -6889
rect 4655 -7065 4689 -6889
rect 4913 -7065 4947 -6889
rect 5027 -7065 5061 -6889
rect 5285 -7065 5319 -6889
rect 5399 -7065 5433 -6889
rect 5657 -7065 5691 -6889
rect 5771 -7065 5805 -6889
rect 6029 -7065 6063 -6889
rect 6143 -7065 6177 -6889
rect 6401 -7065 6435 -6889
rect 6515 -7065 6549 -6889
rect 6773 -7065 6807 -6889
rect 6887 -7065 6921 -6889
rect 7145 -7065 7179 -6889
rect 7259 -7065 7293 -6889
rect 7517 -7065 7551 -6889
rect 7631 -7065 7665 -6889
rect 7889 -7065 7923 -6889
rect 8003 -7065 8037 -6889
rect 8261 -7065 8295 -6889
rect 8375 -7065 8409 -6889
rect 8633 -7065 8667 -6889
rect 8747 -7065 8781 -6889
rect 9005 -7065 9039 -6889
rect 9119 -7065 9153 -6889
rect 9377 -7065 9411 -6889
rect 9491 -7065 9525 -6889
rect 9749 -7065 9783 -6889
rect 997 -7149 1165 -7115
rect 1369 -7149 1537 -7115
rect 1741 -7149 1909 -7115
rect 2113 -7149 2281 -7115
rect 2485 -7149 2653 -7115
rect 2857 -7149 3025 -7115
rect 3229 -7149 3397 -7115
rect 3601 -7149 3769 -7115
rect 3973 -7149 4141 -7115
rect 4345 -7149 4513 -7115
rect 4717 -7149 4885 -7115
rect 5089 -7149 5257 -7115
rect 5461 -7149 5629 -7115
rect 5833 -7149 6001 -7115
rect 6205 -7149 6373 -7115
rect 6577 -7149 6745 -7115
rect 6949 -7149 7117 -7115
rect 7321 -7149 7489 -7115
rect 7693 -7149 7861 -7115
rect 8065 -7149 8233 -7115
rect 8437 -7149 8605 -7115
rect 8809 -7149 8977 -7115
rect 9181 -7149 9349 -7115
rect 9553 -7149 9721 -7115
rect 997 -7257 1165 -7223
rect 1369 -7257 1537 -7223
rect 1741 -7257 1909 -7223
rect 2113 -7257 2281 -7223
rect 2485 -7257 2653 -7223
rect 2857 -7257 3025 -7223
rect 3229 -7257 3397 -7223
rect 3601 -7257 3769 -7223
rect 3973 -7257 4141 -7223
rect 4345 -7257 4513 -7223
rect 4717 -7257 4885 -7223
rect 5089 -7257 5257 -7223
rect 5461 -7257 5629 -7223
rect 5833 -7257 6001 -7223
rect 6205 -7257 6373 -7223
rect 6577 -7257 6745 -7223
rect 6949 -7257 7117 -7223
rect 7321 -7257 7489 -7223
rect 7693 -7257 7861 -7223
rect 8065 -7257 8233 -7223
rect 8437 -7257 8605 -7223
rect 8809 -7257 8977 -7223
rect 9181 -7257 9349 -7223
rect 9553 -7257 9721 -7223
rect 935 -7483 969 -7307
rect 1193 -7483 1227 -7307
rect 1307 -7483 1341 -7307
rect 1565 -7483 1599 -7307
rect 1679 -7483 1713 -7307
rect 1937 -7483 1971 -7307
rect 2051 -7483 2085 -7307
rect 2309 -7483 2343 -7307
rect 2423 -7483 2457 -7307
rect 2681 -7483 2715 -7307
rect 2795 -7483 2829 -7307
rect 3053 -7483 3087 -7307
rect 3167 -7483 3201 -7307
rect 3425 -7483 3459 -7307
rect 3539 -7483 3573 -7307
rect 3797 -7483 3831 -7307
rect 3911 -7483 3945 -7307
rect 4169 -7483 4203 -7307
rect 4283 -7483 4317 -7307
rect 4541 -7483 4575 -7307
rect 4655 -7483 4689 -7307
rect 4913 -7483 4947 -7307
rect 5027 -7483 5061 -7307
rect 5285 -7483 5319 -7307
rect 5399 -7483 5433 -7307
rect 5657 -7483 5691 -7307
rect 5771 -7483 5805 -7307
rect 6029 -7483 6063 -7307
rect 6143 -7483 6177 -7307
rect 6401 -7483 6435 -7307
rect 6515 -7483 6549 -7307
rect 6773 -7483 6807 -7307
rect 6887 -7483 6921 -7307
rect 7145 -7483 7179 -7307
rect 7259 -7483 7293 -7307
rect 7517 -7483 7551 -7307
rect 7631 -7483 7665 -7307
rect 7889 -7483 7923 -7307
rect 8003 -7483 8037 -7307
rect 8261 -7483 8295 -7307
rect 8375 -7483 8409 -7307
rect 8633 -7483 8667 -7307
rect 8747 -7483 8781 -7307
rect 9005 -7483 9039 -7307
rect 9119 -7483 9153 -7307
rect 9377 -7483 9411 -7307
rect 9491 -7483 9525 -7307
rect 9749 -7483 9783 -7307
rect 997 -7567 1165 -7533
rect 1369 -7567 1537 -7533
rect 1741 -7567 1909 -7533
rect 2113 -7567 2281 -7533
rect 2485 -7567 2653 -7533
rect 2857 -7567 3025 -7533
rect 3229 -7567 3397 -7533
rect 3601 -7567 3769 -7533
rect 3973 -7567 4141 -7533
rect 4345 -7567 4513 -7533
rect 4717 -7567 4885 -7533
rect 5089 -7567 5257 -7533
rect 5461 -7567 5629 -7533
rect 5833 -7567 6001 -7533
rect 6205 -7567 6373 -7533
rect 6577 -7567 6745 -7533
rect 6949 -7567 7117 -7533
rect 7321 -7567 7489 -7533
rect 7693 -7567 7861 -7533
rect 8065 -7567 8233 -7533
rect 8437 -7567 8605 -7533
rect 8809 -7567 8977 -7533
rect 9181 -7567 9349 -7533
rect 9553 -7567 9721 -7533
rect 936 -7635 1006 -7624
rect 1604 -7635 1674 -7616
rect 2348 -7635 2418 -7616
rect 3092 -7635 3162 -7616
rect 3836 -7635 3906 -7616
rect 4580 -7635 4650 -7616
rect 5324 -7635 5394 -7616
rect 6068 -7635 6138 -7616
rect 6812 -7635 6882 -7616
rect 7556 -7635 7626 -7616
rect 8300 -7635 8370 -7616
rect 9044 -7635 9114 -7616
rect 9706 -7635 9776 -7620
rect 936 -7669 1006 -7635
rect 1604 -7669 1674 -7635
rect 2348 -7669 2418 -7635
rect 3092 -7669 3162 -7635
rect 3836 -7669 3906 -7635
rect 4580 -7669 4650 -7635
rect 5324 -7669 5394 -7635
rect 6068 -7669 6138 -7635
rect 6812 -7669 6882 -7635
rect 7556 -7669 7626 -7635
rect 8300 -7669 8370 -7635
rect 9044 -7669 9114 -7635
rect 9706 -7669 9776 -7635
rect 936 -7694 1006 -7669
rect 1604 -7686 1674 -7669
rect 2348 -7686 2418 -7669
rect 3092 -7686 3162 -7669
rect 3836 -7686 3906 -7669
rect 4580 -7686 4650 -7669
rect 5324 -7686 5394 -7669
rect 6068 -7686 6138 -7669
rect 6812 -7686 6882 -7669
rect 7556 -7686 7626 -7669
rect 8300 -7686 8370 -7669
rect 9044 -7686 9114 -7669
rect 9706 -7690 9776 -7669
<< metal1 >>
rect -332 1314 -322 1514
rect -122 1314 -112 1514
rect 412 1314 422 1514
rect 622 1314 632 1514
rect 1156 1314 1166 1514
rect 1366 1314 1376 1514
rect 1900 1314 1910 1514
rect 2110 1314 2120 1514
rect 2644 1314 2654 1514
rect 2854 1314 2864 1514
rect 3388 1314 3398 1514
rect 3598 1314 3608 1514
rect 4132 1314 4142 1514
rect 4342 1314 4352 1514
rect 4876 1314 4886 1514
rect 5086 1314 5096 1514
rect 5248 1314 5258 1514
rect 5458 1314 5468 1514
rect 5992 1314 6002 1514
rect 6202 1314 6212 1514
rect 6736 1314 6746 1514
rect 6946 1314 6956 1514
rect 7480 1314 7490 1514
rect 7690 1314 7700 1514
rect 8224 1314 8234 1514
rect 8434 1314 8444 1514
rect 8968 1314 8978 1514
rect 9178 1314 9188 1514
rect 9712 1314 9722 1514
rect 9922 1314 9932 1514
rect 10456 1314 10466 1514
rect 10666 1314 10676 1514
rect 11200 1314 11210 1514
rect 11410 1314 11420 1514
rect -250 1238 -192 1314
rect 494 1238 552 1314
rect 1238 1238 1296 1314
rect 1982 1238 2040 1314
rect 2726 1238 2784 1314
rect 3470 1238 3528 1314
rect 4214 1238 4272 1314
rect 4938 1304 5016 1314
rect 4958 1238 5016 1304
rect 5368 1238 5420 1314
rect 6074 1238 6132 1314
rect 6818 1238 6876 1314
rect 7562 1238 7620 1314
rect 8306 1238 8364 1314
rect 9050 1238 9108 1314
rect 9794 1238 9852 1314
rect 10538 1238 10596 1314
rect 11264 1298 11340 1314
rect 11264 1238 11322 1298
rect -268 1232 -174 1238
rect -268 1162 -256 1232
rect -186 1162 -174 1232
rect -268 1156 -174 1162
rect 476 1232 570 1238
rect 476 1162 488 1232
rect 558 1162 570 1232
rect 476 1156 570 1162
rect 1220 1232 1314 1238
rect 1220 1162 1232 1232
rect 1302 1162 1314 1232
rect 1220 1156 1314 1162
rect 1964 1232 2058 1238
rect 1964 1162 1976 1232
rect 2046 1162 2058 1232
rect 1964 1156 2058 1162
rect 2708 1232 2802 1238
rect 2708 1162 2720 1232
rect 2790 1162 2802 1232
rect 2708 1156 2802 1162
rect 3452 1232 3546 1238
rect 3452 1162 3464 1232
rect 3534 1162 3546 1232
rect 3452 1156 3546 1162
rect 4196 1232 4290 1238
rect 4196 1162 4208 1232
rect 4278 1162 4290 1232
rect 4196 1156 4290 1162
rect 4940 1232 5034 1238
rect 4940 1162 4952 1232
rect 5022 1162 5034 1232
rect 4940 1156 5034 1162
rect 5312 1232 5420 1238
rect 5312 1162 5324 1232
rect 5394 1162 5420 1232
rect 5312 1156 5420 1162
rect 6056 1232 6150 1238
rect 6056 1162 6068 1232
rect 6138 1162 6150 1232
rect 6056 1156 6150 1162
rect 6800 1232 6894 1238
rect 6800 1162 6812 1232
rect 6882 1162 6894 1232
rect 6800 1156 6894 1162
rect 7544 1232 7638 1238
rect 7544 1162 7556 1232
rect 7626 1162 7638 1232
rect 7544 1156 7638 1162
rect 8288 1232 8382 1238
rect 8288 1162 8300 1232
rect 8370 1162 8382 1232
rect 8288 1156 8382 1162
rect 9032 1232 9126 1238
rect 9032 1162 9044 1232
rect 9114 1162 9126 1232
rect 9032 1156 9126 1162
rect 9776 1232 9870 1238
rect 9776 1162 9788 1232
rect 9858 1162 9870 1232
rect 9776 1156 9870 1162
rect 10520 1232 10614 1238
rect 10520 1162 10532 1232
rect 10602 1162 10614 1232
rect 10520 1156 10614 1162
rect 11210 1232 11322 1238
rect 11210 1162 11222 1232
rect 11292 1162 11322 1232
rect 11210 1156 11322 1162
rect -560 1066 -492 1126
rect -322 1119 -312 1126
rect -322 1073 -311 1119
rect -322 1066 -312 1073
rect -560 1020 -512 1066
rect -250 1032 -192 1156
rect -130 1119 -120 1126
rect -131 1073 -120 1119
rect 50 1119 60 1126
rect 242 1119 252 1126
rect -130 1066 -120 1073
rect 50 1073 61 1119
rect 241 1073 252 1119
rect 422 1119 432 1126
rect 50 1066 60 1073
rect 242 1066 252 1073
rect 422 1073 433 1119
rect 422 1066 432 1073
rect 494 1032 552 1156
rect 614 1119 624 1126
rect 613 1073 624 1119
rect 614 1066 624 1073
rect 794 1066 996 1126
rect 1166 1119 1176 1126
rect 1166 1073 1177 1119
rect 1166 1066 1176 1073
rect 866 1032 924 1066
rect 1238 1032 1296 1156
rect 1358 1119 1368 1126
rect 1357 1073 1368 1119
rect 1538 1119 1548 1126
rect 1730 1119 1740 1126
rect 1358 1066 1368 1073
rect 1538 1073 1549 1119
rect 1729 1073 1740 1119
rect 1910 1119 1920 1126
rect 1538 1066 1548 1073
rect 1730 1066 1740 1073
rect 1910 1073 1921 1119
rect 1910 1066 1920 1073
rect 1982 1032 2040 1156
rect 2102 1119 2112 1126
rect 2101 1073 2112 1119
rect 2102 1066 2112 1073
rect 2282 1066 2484 1126
rect 2654 1119 2664 1126
rect 2654 1073 2665 1119
rect 2654 1066 2664 1073
rect 2354 1032 2412 1066
rect 2726 1032 2784 1156
rect 2846 1119 2856 1126
rect 2845 1073 2856 1119
rect 3026 1119 3036 1126
rect 3218 1119 3228 1126
rect 2846 1066 2856 1073
rect 3026 1073 3037 1119
rect 3217 1073 3228 1119
rect 3398 1119 3408 1126
rect 3026 1066 3036 1073
rect 3218 1066 3228 1073
rect 3398 1073 3409 1119
rect 3398 1066 3408 1073
rect 3470 1032 3528 1156
rect 3590 1119 3600 1126
rect 3589 1073 3600 1119
rect 3590 1066 3600 1073
rect 3770 1066 3972 1126
rect 4142 1119 4152 1126
rect 4142 1073 4153 1119
rect 4142 1066 4152 1073
rect 3842 1032 3900 1066
rect 4214 1032 4272 1156
rect 4334 1119 4344 1126
rect 4333 1073 4344 1119
rect 4514 1119 4524 1126
rect 4706 1119 4716 1126
rect 4334 1066 4344 1073
rect 4514 1073 4525 1119
rect 4705 1073 4716 1119
rect 4886 1119 4896 1126
rect 4514 1066 4524 1073
rect 4706 1066 4716 1073
rect 4886 1073 4897 1119
rect 4886 1066 4896 1073
rect 4958 1032 5016 1156
rect 5078 1119 5088 1126
rect 5077 1073 5088 1119
rect 5078 1066 5088 1073
rect 5258 1066 5330 1126
rect -560 644 -553 1020
rect -519 644 -512 1020
rect -560 592 -512 644
rect -301 1020 -141 1032
rect -301 644 -295 1020
rect -261 644 -181 1020
rect -147 644 -141 1020
rect -301 632 -141 644
rect 71 1020 231 1032
rect 71 644 77 1020
rect 111 644 191 1020
rect 225 644 231 1020
rect 71 632 231 644
rect 443 1020 603 1032
rect 443 644 449 1020
rect 483 644 563 1020
rect 597 644 603 1020
rect 443 632 603 644
rect 815 1020 975 1032
rect 815 644 821 1020
rect 855 644 935 1020
rect 969 644 975 1020
rect 815 632 975 644
rect 1187 1020 1347 1032
rect 1187 644 1193 1020
rect 1227 644 1307 1020
rect 1341 644 1347 1020
rect 1187 632 1347 644
rect 1559 1020 1719 1032
rect 1559 644 1565 1020
rect 1599 644 1679 1020
rect 1713 644 1719 1020
rect 1559 632 1719 644
rect 1931 1020 2091 1032
rect 1931 644 1937 1020
rect 1971 644 2051 1020
rect 2085 644 2091 1020
rect 1931 632 2091 644
rect 2303 1020 2463 1032
rect 2303 644 2309 1020
rect 2343 644 2423 1020
rect 2457 644 2463 1020
rect 2303 632 2463 644
rect 2675 1020 2835 1032
rect 2675 644 2681 1020
rect 2715 644 2795 1020
rect 2829 644 2835 1020
rect 2675 632 2835 644
rect 3047 1020 3207 1032
rect 3047 644 3053 1020
rect 3087 644 3167 1020
rect 3201 644 3207 1020
rect 3047 632 3207 644
rect 3419 1020 3579 1032
rect 3419 644 3425 1020
rect 3459 644 3539 1020
rect 3573 644 3579 1020
rect 3419 632 3579 644
rect 3791 1020 3951 1032
rect 3791 644 3797 1020
rect 3831 644 3911 1020
rect 3945 644 3951 1020
rect 3791 632 3951 644
rect 4163 1020 4323 1032
rect 4163 644 4169 1020
rect 4203 644 4283 1020
rect 4317 644 4323 1020
rect 4163 632 4323 644
rect 4535 1020 4695 1032
rect 4535 644 4541 1020
rect 4575 644 4655 1020
rect 4689 644 4695 1020
rect 4535 632 4695 644
rect 4907 1020 5067 1032
rect 4907 644 4913 1020
rect 4947 644 5027 1020
rect 5061 644 5067 1020
rect 4907 632 5067 644
rect 5278 1020 5330 1066
rect 5278 644 5285 1020
rect 5319 644 5330 1020
rect -560 591 -472 592
rect -560 586 -311 591
rect -560 442 -492 586
rect -322 545 -311 586
rect -322 483 -312 545
rect -322 442 -311 483
rect -560 437 -311 442
rect -560 436 -474 437
rect -560 384 -512 436
rect -256 396 -186 632
rect -131 586 61 591
rect -131 545 -120 586
rect -130 483 -120 545
rect -131 442 -120 483
rect 50 545 61 586
rect 50 483 60 545
rect 50 442 61 483
rect -131 437 61 442
rect 116 396 186 632
rect 241 586 433 591
rect 241 545 252 586
rect 242 483 252 545
rect 241 442 252 483
rect 422 545 433 586
rect 422 483 432 545
rect 422 442 433 483
rect 241 437 433 442
rect 488 396 558 632
rect 613 590 805 591
rect 860 590 930 632
rect 985 590 1177 591
rect 613 586 1177 590
rect 613 545 624 586
rect 614 483 624 545
rect 613 442 624 483
rect 794 442 996 586
rect 1166 545 1177 586
rect 1166 483 1176 545
rect 1166 442 1177 483
rect 613 438 1177 442
rect 613 437 805 438
rect 860 396 930 438
rect 985 437 1177 438
rect 1232 396 1302 632
rect 1357 586 1549 591
rect 1357 545 1368 586
rect 1358 483 1368 545
rect 1357 442 1368 483
rect 1538 545 1549 586
rect 1538 483 1548 545
rect 1538 442 1549 483
rect 1357 437 1549 442
rect 1604 396 1674 632
rect 1729 586 1921 591
rect 1729 545 1740 586
rect 1730 483 1740 545
rect 1729 442 1740 483
rect 1910 545 1921 586
rect 1910 483 1920 545
rect 1910 442 1921 483
rect 1729 437 1921 442
rect 1976 396 2046 632
rect 2348 592 2418 632
rect 2156 591 2574 592
rect 2101 586 2665 591
rect 2101 545 2112 586
rect 2102 483 2112 545
rect 2101 442 2112 483
rect 2282 442 2484 586
rect 2654 545 2665 586
rect 2654 483 2664 545
rect 2654 442 2665 483
rect 2101 437 2665 442
rect 2156 436 2574 437
rect 2348 396 2418 436
rect 2720 396 2790 632
rect 2845 586 3037 591
rect 2845 545 2856 586
rect 2846 483 2856 545
rect 2845 442 2856 483
rect 3026 545 3037 586
rect 3026 483 3036 545
rect 3026 442 3037 483
rect 2845 437 3037 442
rect 3092 396 3162 632
rect 3217 586 3409 591
rect 3217 545 3228 586
rect 3218 483 3228 545
rect 3217 442 3228 483
rect 3398 545 3409 586
rect 3398 483 3408 545
rect 3398 442 3409 483
rect 3217 437 3409 442
rect 3464 396 3534 632
rect 3836 592 3906 632
rect 3684 591 4060 592
rect 3589 586 4153 591
rect 3589 545 3600 586
rect 3590 483 3600 545
rect 3589 442 3600 483
rect 3770 442 3972 586
rect 4142 545 4153 586
rect 4142 483 4152 545
rect 4142 442 4153 483
rect 3589 437 4153 442
rect 3684 436 4060 437
rect 3836 396 3906 436
rect 4208 396 4278 632
rect 4333 586 4525 591
rect 4333 545 4344 586
rect 4334 483 4344 545
rect 4333 442 4344 483
rect 4514 545 4525 586
rect 4514 483 4524 545
rect 4514 442 4525 483
rect 4333 437 4525 442
rect 4580 396 4650 632
rect 4705 586 4897 591
rect 4705 545 4716 586
rect 4706 483 4716 545
rect 4705 442 4716 483
rect 4886 545 4897 586
rect 4886 483 4896 545
rect 4886 442 4897 483
rect 4705 437 4897 442
rect 4952 396 5022 632
rect 5278 592 5330 644
rect 5172 591 5330 592
rect 5077 586 5330 591
rect 5077 545 5088 586
rect 5078 483 5088 545
rect 5077 442 5088 483
rect 5258 442 5330 586
rect 5077 437 5330 442
rect 5172 436 5330 437
rect -560 8 -553 384
rect -519 8 -512 384
rect -560 -44 -512 8
rect -301 384 -141 396
rect -301 8 -295 384
rect -261 8 -181 384
rect -147 8 -141 384
rect -301 -4 -141 8
rect 71 384 231 396
rect 71 8 77 384
rect 111 8 191 384
rect 225 8 231 384
rect 71 -4 231 8
rect 443 384 603 396
rect 443 8 449 384
rect 483 8 563 384
rect 597 8 603 384
rect 443 -4 603 8
rect 815 384 975 396
rect 815 8 821 384
rect 855 8 935 384
rect 969 8 975 384
rect 815 -4 975 8
rect 1187 384 1347 396
rect 1187 8 1193 384
rect 1227 8 1307 384
rect 1341 8 1347 384
rect 1187 -4 1347 8
rect 1559 384 1719 396
rect 1559 8 1565 384
rect 1599 8 1679 384
rect 1713 8 1719 384
rect 1559 -4 1719 8
rect 1931 384 2091 396
rect 1931 8 1937 384
rect 1971 8 2051 384
rect 2085 8 2091 384
rect 1931 -4 2091 8
rect 2303 384 2463 396
rect 2303 8 2309 384
rect 2343 8 2423 384
rect 2457 8 2463 384
rect 2303 -4 2463 8
rect 2675 384 2835 396
rect 2675 8 2681 384
rect 2715 8 2795 384
rect 2829 8 2835 384
rect 2675 -4 2835 8
rect 3047 384 3207 396
rect 3047 8 3053 384
rect 3087 8 3167 384
rect 3201 8 3207 384
rect 3047 -4 3207 8
rect 3419 384 3579 396
rect 3419 8 3425 384
rect 3459 8 3539 384
rect 3573 8 3579 384
rect 3419 -4 3579 8
rect 3791 384 3951 396
rect 3791 8 3797 384
rect 3831 8 3911 384
rect 3945 8 3951 384
rect 3791 -4 3951 8
rect 4163 384 4323 396
rect 4163 8 4169 384
rect 4203 8 4283 384
rect 4317 8 4323 384
rect 4163 -4 4323 8
rect 4535 384 4695 396
rect 4535 8 4541 384
rect 4575 8 4655 384
rect 4689 8 4695 384
rect 4535 -4 4695 8
rect 4907 384 5067 396
rect 4907 8 4913 384
rect 4947 8 5027 384
rect 5061 8 5067 384
rect 4907 -4 5067 8
rect 5278 384 5330 436
rect 5278 8 5285 384
rect 5319 8 5330 384
rect -560 -45 -470 -44
rect -560 -50 -311 -45
rect -560 -194 -492 -50
rect -322 -91 -311 -50
rect -322 -153 -312 -91
rect -322 -194 -311 -153
rect -560 -199 -311 -194
rect -560 -204 -470 -199
rect -560 -252 -512 -204
rect -256 -240 -186 -4
rect -131 -50 61 -45
rect -131 -91 -120 -50
rect -130 -153 -120 -91
rect -131 -194 -120 -153
rect 50 -91 61 -50
rect 50 -153 60 -91
rect 50 -194 61 -153
rect -131 -199 61 -194
rect 116 -240 186 -4
rect 241 -50 433 -45
rect 241 -91 252 -50
rect 242 -153 252 -91
rect 241 -194 252 -153
rect 422 -91 433 -50
rect 422 -153 432 -91
rect 422 -194 433 -153
rect 241 -199 433 -194
rect 488 -240 558 -4
rect 613 -48 805 -45
rect 860 -48 930 -4
rect 985 -48 1177 -45
rect 613 -50 1177 -48
rect 613 -91 624 -50
rect 614 -153 624 -91
rect 613 -194 624 -153
rect 794 -194 996 -50
rect 1166 -91 1177 -50
rect 1166 -153 1176 -91
rect 1166 -194 1177 -153
rect 613 -199 1177 -194
rect 654 -200 1130 -199
rect 860 -240 930 -200
rect 1232 -240 1302 -4
rect 1357 -50 1549 -45
rect 1357 -91 1368 -50
rect 1358 -153 1368 -91
rect 1357 -194 1368 -153
rect 1538 -91 1549 -50
rect 1538 -153 1548 -91
rect 1538 -194 1549 -153
rect 1357 -199 1549 -194
rect 1604 -240 1674 -4
rect 1729 -50 1921 -45
rect 1729 -91 1740 -50
rect 1730 -153 1740 -91
rect 1729 -194 1740 -153
rect 1910 -91 1921 -50
rect 1910 -153 1920 -91
rect 1910 -194 1921 -153
rect 1729 -199 1921 -194
rect 1976 -240 2046 -4
rect 2348 -44 2418 -4
rect 2176 -45 2594 -44
rect 2101 -50 2665 -45
rect 2101 -91 2112 -50
rect 2102 -153 2112 -91
rect 2101 -194 2112 -153
rect 2282 -194 2484 -50
rect 2654 -91 2665 -50
rect 2654 -153 2664 -91
rect 2654 -194 2665 -153
rect 2101 -199 2665 -194
rect 2176 -200 2594 -199
rect 2348 -240 2418 -200
rect 2720 -240 2790 -4
rect 2845 -50 3037 -45
rect 2845 -91 2856 -50
rect 2846 -153 2856 -91
rect 2845 -194 2856 -153
rect 3026 -91 3037 -50
rect 3026 -153 3036 -91
rect 3026 -194 3037 -153
rect 2845 -199 3037 -194
rect 3092 -240 3162 -4
rect 3217 -50 3409 -45
rect 3217 -91 3228 -50
rect 3218 -153 3228 -91
rect 3217 -194 3228 -153
rect 3398 -91 3409 -50
rect 3398 -153 3408 -91
rect 3398 -194 3409 -153
rect 3217 -199 3409 -194
rect 3464 -240 3534 -4
rect 3836 -44 3906 -4
rect 3672 -45 4048 -44
rect 3589 -50 4153 -45
rect 3589 -91 3600 -50
rect 3590 -153 3600 -91
rect 3589 -194 3600 -153
rect 3770 -194 3972 -50
rect 4142 -91 4153 -50
rect 4142 -153 4152 -91
rect 4142 -194 4153 -153
rect 3589 -199 4153 -194
rect 3672 -200 4048 -199
rect 3836 -240 3906 -200
rect 4208 -240 4278 -4
rect 4333 -50 4525 -45
rect 4333 -91 4344 -50
rect 4334 -153 4344 -91
rect 4333 -194 4344 -153
rect 4514 -91 4525 -50
rect 4514 -153 4524 -91
rect 4514 -194 4525 -153
rect 4333 -199 4525 -194
rect 4580 -240 4650 -4
rect 4705 -50 4897 -45
rect 4705 -91 4716 -50
rect 4706 -153 4716 -91
rect 4705 -194 4716 -153
rect 4886 -91 4897 -50
rect 4886 -153 4896 -91
rect 4886 -194 4897 -153
rect 4705 -199 4897 -194
rect 4952 -240 5022 -4
rect 5278 -44 5330 8
rect 5188 -45 5330 -44
rect 5077 -50 5330 -45
rect 5077 -91 5088 -50
rect 5078 -153 5088 -91
rect 5077 -194 5088 -153
rect 5258 -194 5330 -50
rect 5077 -199 5330 -194
rect 5188 -200 5330 -199
rect -560 -628 -553 -252
rect -519 -628 -512 -252
rect -560 -674 -512 -628
rect -301 -252 -141 -240
rect -301 -628 -295 -252
rect -261 -628 -181 -252
rect -147 -628 -141 -252
rect -301 -640 -141 -628
rect 71 -252 231 -240
rect 71 -628 77 -252
rect 111 -628 191 -252
rect 225 -628 231 -252
rect 71 -640 231 -628
rect 443 -252 603 -240
rect 443 -628 449 -252
rect 483 -628 563 -252
rect 597 -628 603 -252
rect 443 -640 603 -628
rect 815 -252 975 -240
rect 815 -628 821 -252
rect 855 -628 935 -252
rect 969 -628 975 -252
rect 815 -640 975 -628
rect 1187 -252 1347 -240
rect 1187 -628 1193 -252
rect 1227 -628 1307 -252
rect 1341 -628 1347 -252
rect 1187 -640 1347 -628
rect 1559 -252 1719 -240
rect 1559 -628 1565 -252
rect 1599 -628 1679 -252
rect 1713 -628 1719 -252
rect 1559 -640 1719 -628
rect 1931 -252 2091 -240
rect 1931 -628 1937 -252
rect 1971 -628 2051 -252
rect 2085 -628 2091 -252
rect 1931 -640 2091 -628
rect 2303 -252 2463 -240
rect 2303 -628 2309 -252
rect 2343 -628 2423 -252
rect 2457 -628 2463 -252
rect 2303 -640 2463 -628
rect 2675 -252 2835 -240
rect 2675 -628 2681 -252
rect 2715 -628 2795 -252
rect 2829 -628 2835 -252
rect 2675 -640 2835 -628
rect 3047 -252 3207 -240
rect 3047 -628 3053 -252
rect 3087 -628 3167 -252
rect 3201 -628 3207 -252
rect 3047 -640 3207 -628
rect 3419 -252 3579 -240
rect 3419 -628 3425 -252
rect 3459 -628 3539 -252
rect 3573 -628 3579 -252
rect 3419 -640 3579 -628
rect 3791 -252 3951 -240
rect 3791 -628 3797 -252
rect 3831 -628 3911 -252
rect 3945 -628 3951 -252
rect 3791 -640 3951 -628
rect 4163 -252 4323 -240
rect 4163 -628 4169 -252
rect 4203 -628 4283 -252
rect 4317 -628 4323 -252
rect 4163 -640 4323 -628
rect 4535 -252 4695 -240
rect 4535 -628 4541 -252
rect 4575 -628 4655 -252
rect 4689 -628 4695 -252
rect 4535 -640 4695 -628
rect 4907 -252 5067 -240
rect 4907 -628 4913 -252
rect 4947 -628 5027 -252
rect 5061 -628 5067 -252
rect 4907 -640 5067 -628
rect 5278 -252 5330 -200
rect 5278 -628 5285 -252
rect 5319 -628 5330 -252
rect -560 -734 -492 -674
rect -322 -681 -312 -674
rect -130 -681 -120 -674
rect -322 -727 -311 -681
rect -131 -727 -120 -681
rect 50 -681 60 -674
rect -322 -734 -312 -727
rect -130 -734 -120 -727
rect 50 -727 61 -681
rect 50 -734 60 -727
rect 122 -982 180 -640
rect 866 -674 924 -640
rect 242 -681 252 -674
rect 241 -727 252 -681
rect 422 -681 432 -674
rect 614 -681 624 -674
rect 242 -734 252 -727
rect 422 -727 433 -681
rect 613 -727 624 -681
rect 422 -734 432 -727
rect 614 -734 624 -727
rect 794 -734 996 -674
rect 1166 -681 1176 -674
rect 1358 -681 1368 -674
rect 1166 -727 1177 -681
rect 1357 -727 1368 -681
rect 1538 -681 1548 -674
rect 1166 -734 1176 -727
rect 1358 -734 1368 -727
rect 1538 -727 1549 -681
rect 1538 -734 1548 -727
rect 740 -736 1070 -734
rect 1610 -982 1668 -640
rect 2354 -674 2412 -640
rect 1730 -681 1740 -674
rect 1729 -727 1740 -681
rect 1910 -681 1920 -674
rect 2102 -681 2112 -674
rect 1730 -734 1740 -727
rect 1910 -727 1921 -681
rect 2101 -727 2112 -681
rect 1910 -734 1920 -727
rect 2102 -734 2112 -727
rect 2282 -734 2484 -674
rect 2654 -681 2664 -674
rect 2846 -681 2856 -674
rect 2654 -727 2665 -681
rect 2845 -727 2856 -681
rect 3026 -681 3036 -674
rect 2654 -734 2664 -727
rect 2846 -734 2856 -727
rect 3026 -727 3037 -681
rect 3026 -734 3036 -727
rect 3098 -982 3156 -640
rect 3842 -674 3900 -640
rect 3218 -681 3228 -674
rect 3217 -727 3228 -681
rect 3398 -681 3408 -674
rect 3590 -681 3600 -674
rect 3218 -734 3228 -727
rect 3398 -727 3409 -681
rect 3589 -727 3600 -681
rect 3398 -734 3408 -727
rect 3590 -734 3600 -727
rect 3770 -734 3972 -674
rect 4142 -681 4152 -674
rect 4334 -681 4344 -674
rect 4142 -727 4153 -681
rect 4333 -727 4344 -681
rect 4514 -681 4524 -674
rect 4142 -734 4152 -727
rect 4334 -734 4344 -727
rect 4514 -727 4525 -681
rect 4514 -734 4524 -727
rect 4586 -982 4644 -640
rect 5278 -674 5330 -628
rect 5368 1032 5420 1156
rect 5454 1066 5460 1126
rect 5630 1119 5640 1126
rect 5822 1119 5832 1126
rect 5630 1073 5641 1119
rect 5821 1073 5832 1119
rect 6002 1119 6012 1126
rect 5630 1066 5640 1073
rect 5822 1066 5832 1073
rect 6002 1073 6013 1119
rect 6002 1066 6012 1073
rect 6074 1032 6132 1156
rect 6194 1119 6204 1126
rect 6193 1073 6204 1119
rect 6374 1119 6384 1126
rect 6566 1119 6576 1126
rect 6194 1066 6204 1073
rect 6374 1073 6385 1119
rect 6565 1073 6576 1119
rect 6746 1119 6756 1126
rect 6374 1066 6384 1073
rect 6566 1066 6576 1073
rect 6746 1073 6757 1119
rect 6746 1066 6756 1073
rect 6818 1032 6876 1156
rect 6938 1119 6948 1126
rect 6937 1073 6948 1119
rect 7118 1119 7128 1126
rect 7310 1119 7320 1126
rect 6938 1066 6948 1073
rect 7118 1073 7129 1119
rect 7309 1073 7320 1119
rect 7490 1119 7500 1126
rect 7118 1066 7128 1073
rect 7310 1066 7320 1073
rect 7490 1073 7501 1119
rect 7490 1066 7500 1073
rect 7562 1032 7620 1156
rect 7682 1119 7692 1126
rect 7681 1073 7692 1119
rect 7862 1119 7872 1126
rect 8054 1119 8064 1126
rect 7682 1066 7692 1073
rect 7862 1073 7873 1119
rect 8053 1073 8064 1119
rect 8234 1119 8244 1126
rect 7862 1066 7872 1073
rect 8054 1066 8064 1073
rect 8234 1073 8245 1119
rect 8234 1066 8244 1073
rect 8306 1032 8364 1156
rect 8426 1119 8436 1126
rect 8425 1073 8436 1119
rect 8606 1119 8616 1126
rect 8798 1119 8808 1126
rect 8426 1066 8436 1073
rect 8606 1073 8617 1119
rect 8797 1073 8808 1119
rect 8978 1119 8988 1126
rect 8606 1066 8616 1073
rect 8798 1066 8808 1073
rect 8978 1073 8989 1119
rect 8978 1066 8988 1073
rect 9050 1032 9108 1156
rect 9170 1119 9180 1126
rect 9169 1073 9180 1119
rect 9350 1119 9360 1126
rect 9542 1119 9552 1126
rect 9170 1066 9180 1073
rect 9350 1073 9361 1119
rect 9541 1073 9552 1119
rect 9722 1119 9732 1126
rect 9350 1066 9360 1073
rect 9542 1066 9552 1073
rect 9722 1073 9733 1119
rect 9722 1066 9732 1073
rect 9794 1032 9852 1156
rect 9914 1119 9924 1126
rect 9913 1073 9924 1119
rect 10094 1119 10104 1126
rect 10286 1119 10296 1126
rect 9914 1066 9924 1073
rect 10094 1073 10105 1119
rect 10285 1073 10296 1119
rect 10466 1119 10476 1126
rect 10094 1066 10104 1073
rect 10286 1066 10296 1073
rect 10466 1073 10477 1119
rect 10466 1066 10476 1073
rect 10538 1032 10596 1156
rect 10658 1119 10668 1126
rect 10657 1073 10668 1119
rect 10838 1119 10848 1126
rect 11030 1119 11040 1126
rect 10658 1066 10668 1073
rect 10838 1073 10849 1119
rect 11029 1073 11040 1119
rect 11210 1119 11220 1126
rect 10838 1066 10848 1073
rect 11030 1066 11040 1073
rect 11210 1073 11221 1119
rect 11210 1066 11220 1073
rect 11264 1032 11322 1156
rect 5368 1020 5439 1032
rect 5368 644 5399 1020
rect 5433 644 5439 1020
rect 5368 632 5439 644
rect 5651 1020 5811 1032
rect 5651 644 5657 1020
rect 5691 644 5771 1020
rect 5805 644 5811 1020
rect 5651 632 5811 644
rect 6023 1020 6183 1032
rect 6023 644 6029 1020
rect 6063 644 6143 1020
rect 6177 644 6183 1020
rect 6023 632 6183 644
rect 6395 1020 6555 1032
rect 6395 644 6401 1020
rect 6435 644 6515 1020
rect 6549 644 6555 1020
rect 6395 632 6555 644
rect 6767 1020 6927 1032
rect 6767 644 6773 1020
rect 6807 644 6887 1020
rect 6921 644 6927 1020
rect 6767 632 6927 644
rect 7139 1020 7299 1032
rect 7139 644 7145 1020
rect 7179 644 7259 1020
rect 7293 644 7299 1020
rect 7139 632 7299 644
rect 7511 1020 7671 1032
rect 7511 644 7517 1020
rect 7551 644 7631 1020
rect 7665 644 7671 1020
rect 7511 632 7671 644
rect 7883 1020 8043 1032
rect 7883 644 7889 1020
rect 7923 644 8003 1020
rect 8037 644 8043 1020
rect 7883 632 8043 644
rect 8255 1020 8415 1032
rect 8255 644 8261 1020
rect 8295 644 8375 1020
rect 8409 644 8415 1020
rect 8255 632 8415 644
rect 8627 1020 8787 1032
rect 8627 644 8633 1020
rect 8667 644 8747 1020
rect 8781 644 8787 1020
rect 8627 632 8787 644
rect 8999 1020 9159 1032
rect 8999 644 9005 1020
rect 9039 644 9119 1020
rect 9153 644 9159 1020
rect 8999 632 9159 644
rect 9371 1020 9531 1032
rect 9371 644 9377 1020
rect 9411 644 9491 1020
rect 9525 644 9531 1020
rect 9371 632 9531 644
rect 9743 1020 9903 1032
rect 9743 644 9749 1020
rect 9783 644 9863 1020
rect 9897 644 9903 1020
rect 9743 632 9903 644
rect 10115 1020 10275 1032
rect 10115 644 10121 1020
rect 10155 644 10235 1020
rect 10269 644 10275 1020
rect 10115 632 10275 644
rect 10487 1020 10647 1032
rect 10487 644 10493 1020
rect 10527 644 10607 1020
rect 10641 644 10647 1020
rect 10487 632 10647 644
rect 10859 1020 11019 1032
rect 10859 644 10865 1020
rect 10899 644 10979 1020
rect 11013 644 11019 1020
rect 10859 632 11019 644
rect 11231 1020 11322 1032
rect 11231 644 11237 1020
rect 11271 644 11322 1020
rect 11231 632 11322 644
rect 5368 396 5420 632
rect 5448 591 5574 592
rect 5448 586 5641 591
rect 5448 442 5460 586
rect 5630 545 5641 586
rect 5630 483 5640 545
rect 5630 442 5641 483
rect 5448 437 5641 442
rect 5448 436 5574 437
rect 5696 396 5766 632
rect 5821 586 6013 591
rect 5821 545 5832 586
rect 5822 483 5832 545
rect 5821 442 5832 483
rect 6002 545 6013 586
rect 6002 483 6012 545
rect 6002 442 6013 483
rect 5821 437 6013 442
rect 6068 396 6138 632
rect 6193 586 6385 591
rect 6193 545 6204 586
rect 6194 483 6204 545
rect 6193 442 6204 483
rect 6374 545 6385 586
rect 6374 483 6384 545
rect 6374 442 6385 483
rect 6193 437 6385 442
rect 6440 396 6510 632
rect 6565 586 6757 591
rect 6565 545 6576 586
rect 6566 483 6576 545
rect 6565 442 6576 483
rect 6746 545 6757 586
rect 6746 483 6756 545
rect 6746 442 6757 483
rect 6565 437 6757 442
rect 6812 396 6882 632
rect 6937 586 7129 591
rect 6937 545 6948 586
rect 6938 483 6948 545
rect 6937 442 6948 483
rect 7118 545 7129 586
rect 7118 483 7128 545
rect 7118 442 7129 483
rect 6937 437 7129 442
rect 7184 396 7254 632
rect 7309 586 7501 591
rect 7309 545 7320 586
rect 7310 483 7320 545
rect 7309 442 7320 483
rect 7490 545 7501 586
rect 7490 483 7500 545
rect 7490 442 7501 483
rect 7309 437 7501 442
rect 7556 396 7626 632
rect 7681 586 7873 591
rect 7681 545 7692 586
rect 7682 483 7692 545
rect 7681 442 7692 483
rect 7862 545 7873 586
rect 7862 483 7872 545
rect 7862 442 7873 483
rect 7681 437 7873 442
rect 7928 396 7998 632
rect 8053 586 8245 591
rect 8053 545 8064 586
rect 8054 483 8064 545
rect 8053 442 8064 483
rect 8234 545 8245 586
rect 8234 483 8244 545
rect 8234 442 8245 483
rect 8053 437 8245 442
rect 8300 396 8370 632
rect 8425 586 8617 591
rect 8425 545 8436 586
rect 8426 483 8436 545
rect 8425 442 8436 483
rect 8606 545 8617 586
rect 8606 483 8616 545
rect 8606 442 8617 483
rect 8425 437 8617 442
rect 8672 396 8742 632
rect 8797 586 8989 591
rect 8797 545 8808 586
rect 8798 483 8808 545
rect 8797 442 8808 483
rect 8978 545 8989 586
rect 8978 483 8988 545
rect 8978 442 8989 483
rect 8797 437 8989 442
rect 9044 396 9114 632
rect 9169 586 9361 591
rect 9169 545 9180 586
rect 9170 483 9180 545
rect 9169 442 9180 483
rect 9350 545 9361 586
rect 9350 483 9360 545
rect 9350 442 9361 483
rect 9169 437 9361 442
rect 9416 396 9486 632
rect 9541 586 9733 591
rect 9541 545 9552 586
rect 9542 483 9552 545
rect 9541 442 9552 483
rect 9722 545 9733 586
rect 9722 483 9732 545
rect 9722 442 9733 483
rect 9541 437 9733 442
rect 9788 396 9858 632
rect 9913 586 10105 591
rect 9913 545 9924 586
rect 9914 483 9924 545
rect 9913 442 9924 483
rect 10094 545 10105 586
rect 10094 483 10104 545
rect 10094 442 10105 483
rect 9913 437 10105 442
rect 10160 396 10230 632
rect 10285 586 10477 591
rect 10285 545 10296 586
rect 10286 483 10296 545
rect 10285 442 10296 483
rect 10466 545 10477 586
rect 10466 483 10476 545
rect 10466 442 10477 483
rect 10285 437 10477 442
rect 10532 396 10602 632
rect 10657 586 10849 591
rect 10657 545 10668 586
rect 10658 483 10668 545
rect 10657 442 10668 483
rect 10838 545 10849 586
rect 10838 483 10848 545
rect 10838 442 10849 483
rect 10657 437 10849 442
rect 10904 396 10974 632
rect 11029 586 11221 591
rect 11029 545 11040 586
rect 11030 483 11040 545
rect 11029 442 11040 483
rect 11210 545 11221 586
rect 11210 483 11220 545
rect 11210 442 11221 483
rect 11029 437 11221 442
rect 11264 396 11322 632
rect 5368 384 5439 396
rect 5368 8 5399 384
rect 5433 8 5439 384
rect 5368 -4 5439 8
rect 5651 384 5811 396
rect 5651 8 5657 384
rect 5691 8 5771 384
rect 5805 8 5811 384
rect 5651 -4 5811 8
rect 6023 384 6183 396
rect 6023 8 6029 384
rect 6063 8 6143 384
rect 6177 8 6183 384
rect 6023 -4 6183 8
rect 6395 384 6555 396
rect 6395 8 6401 384
rect 6435 8 6515 384
rect 6549 8 6555 384
rect 6395 -4 6555 8
rect 6767 384 6927 396
rect 6767 8 6773 384
rect 6807 8 6887 384
rect 6921 8 6927 384
rect 6767 -4 6927 8
rect 7139 384 7299 396
rect 7139 8 7145 384
rect 7179 8 7259 384
rect 7293 8 7299 384
rect 7139 -4 7299 8
rect 7511 384 7671 396
rect 7511 8 7517 384
rect 7551 8 7631 384
rect 7665 8 7671 384
rect 7511 -4 7671 8
rect 7883 384 8043 396
rect 7883 8 7889 384
rect 7923 8 8003 384
rect 8037 8 8043 384
rect 7883 -4 8043 8
rect 8255 384 8415 396
rect 8255 8 8261 384
rect 8295 8 8375 384
rect 8409 8 8415 384
rect 8255 -4 8415 8
rect 8627 384 8787 396
rect 8627 8 8633 384
rect 8667 8 8747 384
rect 8781 8 8787 384
rect 8627 -4 8787 8
rect 8999 384 9159 396
rect 8999 8 9005 384
rect 9039 8 9119 384
rect 9153 8 9159 384
rect 8999 -4 9159 8
rect 9371 384 9531 396
rect 9371 8 9377 384
rect 9411 8 9491 384
rect 9525 8 9531 384
rect 9371 -4 9531 8
rect 9743 384 9903 396
rect 9743 8 9749 384
rect 9783 8 9863 384
rect 9897 8 9903 384
rect 9743 -4 9903 8
rect 10115 384 10275 396
rect 10115 8 10121 384
rect 10155 8 10235 384
rect 10269 8 10275 384
rect 10115 -4 10275 8
rect 10487 384 10647 396
rect 10487 8 10493 384
rect 10527 8 10607 384
rect 10641 8 10647 384
rect 10487 -4 10647 8
rect 10859 384 11019 396
rect 10859 8 10865 384
rect 10899 8 10979 384
rect 11013 8 11019 384
rect 10859 -4 11019 8
rect 11231 384 11322 396
rect 11231 8 11237 384
rect 11271 8 11322 384
rect 11231 -4 11322 8
rect 5368 -240 5420 -4
rect 5448 -45 5590 -44
rect 5448 -50 5641 -45
rect 5448 -194 5460 -50
rect 5630 -91 5641 -50
rect 5630 -153 5640 -91
rect 5630 -194 5641 -153
rect 5448 -199 5641 -194
rect 5448 -200 5590 -199
rect 5696 -240 5766 -4
rect 5821 -50 6013 -45
rect 5821 -91 5832 -50
rect 5822 -153 5832 -91
rect 5821 -194 5832 -153
rect 6002 -91 6013 -50
rect 6002 -153 6012 -91
rect 6002 -194 6013 -153
rect 5821 -199 6013 -194
rect 6068 -240 6138 -4
rect 6193 -50 6385 -45
rect 6193 -91 6204 -50
rect 6194 -153 6204 -91
rect 6193 -194 6204 -153
rect 6374 -91 6385 -50
rect 6374 -153 6384 -91
rect 6374 -194 6385 -153
rect 6193 -199 6385 -194
rect 6440 -240 6510 -4
rect 6565 -50 6757 -45
rect 6565 -91 6576 -50
rect 6566 -153 6576 -91
rect 6565 -194 6576 -153
rect 6746 -91 6757 -50
rect 6746 -153 6756 -91
rect 6746 -194 6757 -153
rect 6565 -199 6757 -194
rect 6812 -240 6882 -4
rect 6937 -50 7129 -45
rect 6937 -91 6948 -50
rect 6938 -153 6948 -91
rect 6937 -194 6948 -153
rect 7118 -91 7129 -50
rect 7118 -153 7128 -91
rect 7118 -194 7129 -153
rect 6937 -199 7129 -194
rect 7184 -240 7254 -4
rect 7309 -50 7501 -45
rect 7309 -91 7320 -50
rect 7310 -153 7320 -91
rect 7309 -194 7320 -153
rect 7490 -91 7501 -50
rect 7490 -153 7500 -91
rect 7490 -194 7501 -153
rect 7309 -199 7501 -194
rect 7556 -240 7626 -4
rect 7681 -50 7873 -45
rect 7681 -91 7692 -50
rect 7682 -153 7692 -91
rect 7681 -194 7692 -153
rect 7862 -91 7873 -50
rect 7862 -153 7872 -91
rect 7862 -194 7873 -153
rect 7681 -199 7873 -194
rect 7928 -240 7998 -4
rect 8053 -50 8245 -45
rect 8053 -91 8064 -50
rect 8054 -153 8064 -91
rect 8053 -194 8064 -153
rect 8234 -91 8245 -50
rect 8234 -153 8244 -91
rect 8234 -194 8245 -153
rect 8053 -199 8245 -194
rect 8300 -240 8370 -4
rect 8425 -50 8617 -45
rect 8425 -91 8436 -50
rect 8426 -153 8436 -91
rect 8425 -194 8436 -153
rect 8606 -91 8617 -50
rect 8606 -153 8616 -91
rect 8606 -194 8617 -153
rect 8425 -199 8617 -194
rect 8672 -240 8742 -4
rect 8797 -50 8989 -45
rect 8797 -91 8808 -50
rect 8798 -153 8808 -91
rect 8797 -194 8808 -153
rect 8978 -91 8989 -50
rect 8978 -153 8988 -91
rect 8978 -194 8989 -153
rect 8797 -199 8989 -194
rect 9044 -240 9114 -4
rect 9169 -50 9361 -45
rect 9169 -91 9180 -50
rect 9170 -153 9180 -91
rect 9169 -194 9180 -153
rect 9350 -91 9361 -50
rect 9350 -153 9360 -91
rect 9350 -194 9361 -153
rect 9169 -199 9361 -194
rect 9416 -240 9486 -4
rect 9541 -50 9733 -45
rect 9541 -91 9552 -50
rect 9542 -153 9552 -91
rect 9541 -194 9552 -153
rect 9722 -91 9733 -50
rect 9722 -153 9732 -91
rect 9722 -194 9733 -153
rect 9541 -199 9733 -194
rect 9788 -240 9858 -4
rect 9913 -50 10105 -45
rect 9913 -91 9924 -50
rect 9914 -153 9924 -91
rect 9913 -194 9924 -153
rect 10094 -91 10105 -50
rect 10094 -153 10104 -91
rect 10094 -194 10105 -153
rect 9913 -199 10105 -194
rect 10160 -240 10230 -4
rect 10285 -50 10477 -45
rect 10285 -91 10296 -50
rect 10286 -153 10296 -91
rect 10285 -194 10296 -153
rect 10466 -91 10477 -50
rect 10466 -153 10476 -91
rect 10466 -194 10477 -153
rect 10285 -199 10477 -194
rect 10532 -240 10602 -4
rect 10657 -50 10849 -45
rect 10657 -91 10668 -50
rect 10658 -153 10668 -91
rect 10657 -194 10668 -153
rect 10838 -91 10849 -50
rect 10838 -153 10848 -91
rect 10838 -194 10849 -153
rect 10657 -199 10849 -194
rect 10904 -240 10974 -4
rect 11029 -50 11221 -45
rect 11029 -91 11040 -50
rect 11030 -153 11040 -91
rect 11029 -194 11040 -153
rect 11210 -91 11221 -50
rect 11210 -153 11220 -91
rect 11210 -194 11221 -153
rect 11029 -199 11221 -194
rect 11264 -240 11322 -4
rect 5368 -252 5439 -240
rect 5368 -628 5399 -252
rect 5433 -628 5439 -252
rect 5368 -640 5439 -628
rect 5651 -252 5811 -240
rect 5651 -628 5657 -252
rect 5691 -628 5771 -252
rect 5805 -628 5811 -252
rect 5651 -640 5811 -628
rect 6023 -252 6183 -240
rect 6023 -628 6029 -252
rect 6063 -628 6143 -252
rect 6177 -628 6183 -252
rect 6023 -640 6183 -628
rect 6395 -252 6555 -240
rect 6395 -628 6401 -252
rect 6435 -628 6515 -252
rect 6549 -628 6555 -252
rect 6395 -640 6555 -628
rect 6767 -252 6927 -240
rect 6767 -628 6773 -252
rect 6807 -628 6887 -252
rect 6921 -628 6927 -252
rect 6767 -640 6927 -628
rect 7139 -252 7299 -240
rect 7139 -628 7145 -252
rect 7179 -628 7259 -252
rect 7293 -628 7299 -252
rect 7139 -640 7299 -628
rect 7511 -252 7671 -240
rect 7511 -628 7517 -252
rect 7551 -628 7631 -252
rect 7665 -628 7671 -252
rect 7511 -640 7671 -628
rect 7883 -252 8043 -240
rect 7883 -628 7889 -252
rect 7923 -628 8003 -252
rect 8037 -628 8043 -252
rect 7883 -640 8043 -628
rect 8255 -252 8415 -240
rect 8255 -628 8261 -252
rect 8295 -628 8375 -252
rect 8409 -628 8415 -252
rect 8255 -640 8415 -628
rect 8627 -252 8787 -240
rect 8627 -628 8633 -252
rect 8667 -628 8747 -252
rect 8781 -628 8787 -252
rect 8627 -640 8787 -628
rect 8999 -252 9159 -240
rect 8999 -628 9005 -252
rect 9039 -628 9119 -252
rect 9153 -628 9159 -252
rect 8999 -640 9159 -628
rect 9371 -252 9531 -240
rect 9371 -628 9377 -252
rect 9411 -628 9491 -252
rect 9525 -628 9531 -252
rect 9371 -640 9531 -628
rect 9743 -252 9903 -240
rect 9743 -628 9749 -252
rect 9783 -628 9863 -252
rect 9897 -628 9903 -252
rect 9743 -640 9903 -628
rect 10115 -252 10275 -240
rect 10115 -628 10121 -252
rect 10155 -628 10235 -252
rect 10269 -628 10275 -252
rect 10115 -640 10275 -628
rect 10487 -252 10647 -240
rect 10487 -628 10493 -252
rect 10527 -628 10607 -252
rect 10641 -628 10647 -252
rect 10487 -640 10647 -628
rect 10859 -252 11019 -240
rect 10859 -628 10865 -252
rect 10899 -628 10979 -252
rect 11013 -628 11019 -252
rect 10859 -640 11019 -628
rect 11231 -252 11322 -240
rect 11231 -628 11237 -252
rect 11271 -628 11322 -252
rect 11231 -640 11322 -628
rect 4706 -681 4716 -674
rect 4705 -727 4716 -681
rect 4886 -681 4896 -674
rect 5078 -681 5088 -674
rect 4706 -734 4716 -727
rect 4886 -727 4897 -681
rect 5077 -727 5088 -681
rect 4886 -734 4896 -727
rect 5078 -734 5088 -727
rect 5258 -734 5330 -674
rect 5446 -734 5460 -674
rect 5630 -681 5640 -674
rect 5630 -727 5641 -681
rect 5630 -734 5640 -727
rect 122 -1046 4644 -982
rect 5696 -1042 5766 -640
rect 5822 -681 5832 -674
rect 5821 -727 5832 -681
rect 6002 -681 6012 -674
rect 6194 -681 6204 -674
rect 5822 -734 5832 -727
rect 6002 -727 6013 -681
rect 6193 -727 6204 -681
rect 6374 -681 6384 -674
rect 6002 -734 6012 -727
rect 6194 -734 6204 -727
rect 6374 -727 6385 -681
rect 6374 -734 6384 -727
rect 6440 -1042 6510 -640
rect 6566 -681 6576 -674
rect 6565 -727 6576 -681
rect 6746 -681 6756 -674
rect 6938 -681 6948 -674
rect 6566 -734 6576 -727
rect 6746 -727 6757 -681
rect 6937 -727 6948 -681
rect 7118 -681 7128 -674
rect 6746 -734 6756 -727
rect 6938 -734 6948 -727
rect 7118 -727 7129 -681
rect 7118 -734 7128 -727
rect 7184 -1042 7254 -640
rect 7310 -681 7320 -674
rect 7309 -727 7320 -681
rect 7490 -681 7500 -674
rect 7682 -681 7692 -674
rect 7310 -734 7320 -727
rect 7490 -727 7501 -681
rect 7681 -727 7692 -681
rect 7862 -681 7872 -674
rect 7490 -734 7500 -727
rect 7682 -734 7692 -727
rect 7862 -727 7873 -681
rect 7862 -734 7872 -727
rect 7928 -1042 7998 -640
rect 8054 -681 8064 -674
rect 8053 -727 8064 -681
rect 8234 -681 8244 -674
rect 8426 -681 8436 -674
rect 8054 -734 8064 -727
rect 8234 -727 8245 -681
rect 8425 -727 8436 -681
rect 8606 -681 8616 -674
rect 8234 -734 8244 -727
rect 8426 -734 8436 -727
rect 8606 -727 8617 -681
rect 8606 -734 8616 -727
rect 8672 -1042 8742 -640
rect 8798 -681 8808 -674
rect 8797 -727 8808 -681
rect 8978 -681 8988 -674
rect 9170 -681 9180 -674
rect 8798 -734 8808 -727
rect 8978 -727 8989 -681
rect 9169 -727 9180 -681
rect 9350 -681 9360 -674
rect 8978 -734 8988 -727
rect 9170 -734 9180 -727
rect 9350 -727 9361 -681
rect 9350 -734 9360 -727
rect 9416 -1042 9486 -640
rect 9542 -681 9552 -674
rect 9541 -727 9552 -681
rect 9722 -681 9732 -674
rect 9914 -681 9924 -674
rect 9542 -734 9552 -727
rect 9722 -727 9733 -681
rect 9913 -727 9924 -681
rect 10094 -681 10104 -674
rect 9722 -734 9732 -727
rect 9914 -734 9924 -727
rect 10094 -727 10105 -681
rect 10094 -734 10104 -727
rect 10160 -1042 10230 -640
rect 10286 -681 10296 -674
rect 10285 -727 10296 -681
rect 10466 -681 10476 -674
rect 10658 -681 10668 -674
rect 10286 -734 10296 -727
rect 10466 -727 10477 -681
rect 10657 -727 10668 -681
rect 10838 -681 10848 -674
rect 10466 -734 10476 -727
rect 10658 -734 10668 -727
rect 10838 -727 10849 -681
rect 10838 -734 10848 -727
rect 10904 -1042 10974 -640
rect 11030 -681 11040 -674
rect 11029 -727 11040 -681
rect 11210 -681 11220 -674
rect 11030 -734 11040 -727
rect 11210 -727 11221 -681
rect 11210 -734 11220 -727
rect 882 -1150 936 -1046
rect 1278 -1150 1348 -1046
rect 1610 -1150 1668 -1046
rect 2022 -1150 2092 -1046
rect 2354 -1150 2412 -1046
rect 2766 -1150 2836 -1046
rect 3098 -1150 3156 -1046
rect 3510 -1150 3580 -1046
rect 3830 -1150 3884 -1046
rect 882 -1156 988 -1150
rect 882 -1226 906 -1156
rect 976 -1226 988 -1156
rect 882 -1232 988 -1226
rect 1266 -1156 1360 -1150
rect 1266 -1226 1278 -1156
rect 1348 -1226 1360 -1156
rect 1266 -1232 1360 -1226
rect 1610 -1156 1732 -1150
rect 1610 -1226 1650 -1156
rect 1720 -1226 1732 -1156
rect 1610 -1232 1732 -1226
rect 2010 -1156 2104 -1150
rect 2010 -1226 2022 -1156
rect 2092 -1226 2104 -1156
rect 2010 -1232 2104 -1226
rect 2354 -1156 2476 -1150
rect 2354 -1226 2394 -1156
rect 2464 -1226 2476 -1156
rect 2354 -1232 2476 -1226
rect 2754 -1156 2848 -1150
rect 2754 -1226 2766 -1156
rect 2836 -1226 2848 -1156
rect 2754 -1232 2848 -1226
rect 3098 -1156 3220 -1150
rect 3098 -1226 3138 -1156
rect 3208 -1226 3220 -1156
rect 3098 -1232 3220 -1226
rect 3498 -1156 3592 -1150
rect 3498 -1226 3510 -1156
rect 3580 -1226 3592 -1156
rect 3498 -1232 3592 -1226
rect 3760 -1156 3884 -1150
rect 3760 -1226 3772 -1156
rect 3842 -1226 3884 -1156
rect 3760 -1232 3884 -1226
rect 882 -1356 936 -1232
rect 986 -1269 996 -1260
rect 985 -1315 996 -1269
rect 1166 -1269 1176 -1260
rect 1358 -1269 1368 -1260
rect 986 -1324 996 -1315
rect 1166 -1315 1177 -1269
rect 1357 -1315 1368 -1269
rect 1538 -1269 1548 -1260
rect 1166 -1324 1176 -1315
rect 1358 -1324 1368 -1315
rect 1538 -1315 1549 -1269
rect 1538 -1324 1548 -1315
rect 1610 -1356 1668 -1232
rect 1730 -1269 1740 -1260
rect 1729 -1315 1740 -1269
rect 1910 -1269 1920 -1260
rect 2102 -1269 2112 -1260
rect 1730 -1324 1740 -1315
rect 1910 -1315 1921 -1269
rect 2101 -1315 2112 -1269
rect 2282 -1269 2292 -1260
rect 1910 -1324 1920 -1315
rect 2102 -1324 2112 -1315
rect 2282 -1315 2293 -1269
rect 2282 -1324 2292 -1315
rect 2354 -1356 2412 -1232
rect 2474 -1269 2484 -1260
rect 2473 -1315 2484 -1269
rect 2654 -1269 2664 -1260
rect 2846 -1269 2856 -1260
rect 2474 -1324 2484 -1315
rect 2654 -1315 2665 -1269
rect 2845 -1315 2856 -1269
rect 3026 -1269 3036 -1260
rect 2654 -1324 2664 -1315
rect 2846 -1324 2856 -1315
rect 3026 -1315 3037 -1269
rect 3026 -1324 3036 -1315
rect 3098 -1356 3156 -1232
rect 3218 -1269 3228 -1260
rect 3217 -1315 3228 -1269
rect 3398 -1269 3408 -1260
rect 3590 -1269 3600 -1260
rect 3218 -1324 3228 -1315
rect 3398 -1315 3409 -1269
rect 3589 -1315 3600 -1269
rect 3770 -1269 3780 -1260
rect 3398 -1324 3408 -1315
rect 3590 -1324 3600 -1315
rect 3770 -1315 3781 -1269
rect 3770 -1324 3780 -1315
rect 3830 -1356 3884 -1232
rect 5582 -1314 5592 -1042
rect 5874 -1314 5884 -1042
rect 6326 -1314 6336 -1042
rect 6618 -1314 6628 -1042
rect 7070 -1314 7080 -1042
rect 7362 -1314 7372 -1042
rect 7814 -1314 7824 -1042
rect 8106 -1314 8116 -1042
rect 8558 -1314 8568 -1042
rect 8850 -1314 8860 -1042
rect 9302 -1314 9312 -1042
rect 9594 -1314 9604 -1042
rect 10046 -1314 10056 -1042
rect 10338 -1314 10348 -1042
rect 10790 -1314 10800 -1042
rect 11082 -1314 11092 -1042
rect 882 -1368 975 -1356
rect 882 -2144 935 -1368
rect 969 -2144 975 -1368
rect 882 -2156 975 -2144
rect 1187 -1368 1347 -1356
rect 1187 -2144 1193 -1368
rect 1227 -2144 1307 -1368
rect 1341 -2144 1347 -1368
rect 1187 -2156 1347 -2144
rect 1559 -1368 1719 -1356
rect 1559 -2144 1565 -1368
rect 1599 -2144 1679 -1368
rect 1713 -2144 1719 -1368
rect 1559 -2156 1719 -2144
rect 1931 -1368 2091 -1356
rect 1931 -2144 1937 -1368
rect 1971 -2144 2051 -1368
rect 2085 -2144 2091 -1368
rect 1931 -2156 2091 -2144
rect 2303 -1368 2463 -1356
rect 2303 -2144 2309 -1368
rect 2343 -2144 2423 -1368
rect 2457 -2144 2463 -1368
rect 2303 -2156 2463 -2144
rect 2675 -1368 2835 -1356
rect 2675 -2144 2681 -1368
rect 2715 -2144 2795 -1368
rect 2829 -2144 2835 -1368
rect 2675 -2156 2835 -2144
rect 3047 -1368 3207 -1356
rect 3047 -2144 3053 -1368
rect 3087 -2144 3167 -1368
rect 3201 -2144 3207 -1368
rect 3047 -2156 3207 -2144
rect 3419 -1368 3579 -1356
rect 3419 -2144 3425 -1368
rect 3459 -2144 3539 -1368
rect 3573 -2144 3579 -1368
rect 3419 -2156 3579 -2144
rect 3791 -1368 3884 -1356
rect 3791 -2144 3797 -1368
rect 3831 -2144 3884 -1368
rect 3791 -2156 3884 -2144
rect 882 -2392 930 -2156
rect 985 -2202 1177 -2197
rect 985 -2243 996 -2202
rect 986 -2305 996 -2243
rect 985 -2346 996 -2305
rect 1166 -2243 1177 -2202
rect 1166 -2305 1176 -2243
rect 1166 -2346 1177 -2305
rect 985 -2351 1177 -2346
rect 1232 -2392 1302 -2156
rect 1357 -2202 1549 -2197
rect 1357 -2243 1368 -2202
rect 1358 -2305 1368 -2243
rect 1357 -2346 1368 -2305
rect 1538 -2243 1549 -2202
rect 1538 -2305 1548 -2243
rect 1538 -2346 1549 -2305
rect 1357 -2351 1549 -2346
rect 1604 -2392 1674 -2156
rect 1729 -2202 1921 -2197
rect 1729 -2243 1740 -2202
rect 1730 -2305 1740 -2243
rect 1729 -2346 1740 -2305
rect 1910 -2243 1921 -2202
rect 1910 -2305 1920 -2243
rect 1910 -2346 1921 -2305
rect 1729 -2351 1921 -2346
rect 1976 -2392 2046 -2156
rect 2101 -2202 2293 -2197
rect 2101 -2243 2112 -2202
rect 2102 -2305 2112 -2243
rect 2101 -2346 2112 -2305
rect 2282 -2243 2293 -2202
rect 2282 -2305 2292 -2243
rect 2282 -2346 2293 -2305
rect 2101 -2351 2293 -2346
rect 2348 -2392 2418 -2156
rect 2473 -2202 2665 -2197
rect 2473 -2243 2484 -2202
rect 2474 -2305 2484 -2243
rect 2473 -2346 2484 -2305
rect 2654 -2243 2665 -2202
rect 2654 -2305 2664 -2243
rect 2654 -2346 2665 -2305
rect 2473 -2351 2665 -2346
rect 2720 -2392 2790 -2156
rect 2845 -2202 3037 -2197
rect 2845 -2243 2856 -2202
rect 2846 -2305 2856 -2243
rect 2845 -2346 2856 -2305
rect 3026 -2243 3037 -2202
rect 3026 -2305 3036 -2243
rect 3026 -2346 3037 -2305
rect 2845 -2351 3037 -2346
rect 3092 -2392 3162 -2156
rect 3217 -2202 3409 -2197
rect 3217 -2243 3228 -2202
rect 3218 -2305 3228 -2243
rect 3217 -2346 3228 -2305
rect 3398 -2243 3409 -2202
rect 3398 -2305 3408 -2243
rect 3398 -2346 3409 -2305
rect 3217 -2351 3409 -2346
rect 3464 -2392 3534 -2156
rect 3589 -2202 3781 -2197
rect 3589 -2243 3600 -2202
rect 3590 -2305 3600 -2243
rect 3589 -2346 3600 -2305
rect 3770 -2243 3781 -2202
rect 3770 -2305 3780 -2243
rect 3770 -2346 3781 -2305
rect 3589 -2351 3781 -2346
rect 3830 -2392 3884 -2156
rect 882 -2404 975 -2392
rect 882 -3180 935 -2404
rect 969 -3180 975 -2404
rect 882 -3192 975 -3180
rect 1187 -2404 1347 -2392
rect 1187 -3180 1193 -2404
rect 1227 -3180 1307 -2404
rect 1341 -3180 1347 -2404
rect 1187 -3192 1347 -3180
rect 1559 -2404 1719 -2392
rect 1559 -3180 1565 -2404
rect 1599 -3180 1679 -2404
rect 1713 -3180 1719 -2404
rect 1559 -3192 1719 -3180
rect 1931 -2404 2091 -2392
rect 1931 -3180 1937 -2404
rect 1971 -3180 2051 -2404
rect 2085 -3180 2091 -2404
rect 1931 -3192 2091 -3180
rect 2303 -2404 2463 -2392
rect 2303 -3180 2309 -2404
rect 2343 -3180 2423 -2404
rect 2457 -3180 2463 -2404
rect 2303 -3192 2463 -3180
rect 2675 -2404 2835 -2392
rect 2675 -3180 2681 -2404
rect 2715 -3180 2795 -2404
rect 2829 -3180 2835 -2404
rect 2675 -3192 2835 -3180
rect 3047 -2404 3207 -2392
rect 3047 -3180 3053 -2404
rect 3087 -3180 3167 -2404
rect 3201 -3180 3207 -2404
rect 3047 -3192 3207 -3180
rect 3419 -2404 3579 -2392
rect 3419 -3180 3425 -2404
rect 3459 -3180 3539 -2404
rect 3573 -3180 3579 -2404
rect 3419 -3192 3579 -3180
rect 3791 -2404 3884 -2392
rect 3791 -3180 3797 -2404
rect 3831 -3180 3884 -2404
rect 6002 -3088 6012 -2816
rect 6294 -3088 6304 -2816
rect 3791 -3192 3884 -3180
rect 882 -3428 930 -3192
rect 985 -3238 1177 -3233
rect 985 -3279 996 -3238
rect 986 -3341 996 -3279
rect 985 -3382 996 -3341
rect 1166 -3279 1177 -3238
rect 1166 -3341 1176 -3279
rect 1166 -3382 1177 -3341
rect 985 -3387 1177 -3382
rect 1232 -3428 1302 -3192
rect 1357 -3238 1549 -3233
rect 1357 -3279 1368 -3238
rect 1358 -3341 1368 -3279
rect 1357 -3382 1368 -3341
rect 1538 -3279 1549 -3238
rect 1538 -3341 1548 -3279
rect 1538 -3382 1549 -3341
rect 1357 -3387 1549 -3382
rect 1604 -3428 1674 -3192
rect 1729 -3238 1921 -3233
rect 1729 -3279 1740 -3238
rect 1730 -3341 1740 -3279
rect 1729 -3382 1740 -3341
rect 1910 -3279 1921 -3238
rect 1910 -3341 1920 -3279
rect 1910 -3382 1921 -3341
rect 1729 -3387 1921 -3382
rect 1976 -3428 2046 -3192
rect 2101 -3238 2293 -3233
rect 2101 -3279 2112 -3238
rect 2102 -3341 2112 -3279
rect 2101 -3382 2112 -3341
rect 2282 -3279 2293 -3238
rect 2282 -3341 2292 -3279
rect 2282 -3382 2293 -3341
rect 2101 -3387 2293 -3382
rect 2348 -3428 2418 -3192
rect 2473 -3238 2665 -3233
rect 2473 -3279 2484 -3238
rect 2474 -3341 2484 -3279
rect 2473 -3382 2484 -3341
rect 2654 -3279 2665 -3238
rect 2654 -3341 2664 -3279
rect 2654 -3382 2665 -3341
rect 2473 -3387 2665 -3382
rect 2720 -3428 2790 -3192
rect 2845 -3238 3037 -3233
rect 2845 -3279 2856 -3238
rect 2846 -3341 2856 -3279
rect 2845 -3382 2856 -3341
rect 3026 -3279 3037 -3238
rect 3026 -3341 3036 -3279
rect 3026 -3382 3037 -3341
rect 2845 -3387 3037 -3382
rect 3092 -3428 3162 -3192
rect 3217 -3238 3409 -3233
rect 3217 -3279 3228 -3238
rect 3218 -3341 3228 -3279
rect 3217 -3382 3228 -3341
rect 3398 -3279 3409 -3238
rect 3398 -3341 3408 -3279
rect 3398 -3382 3409 -3341
rect 3217 -3387 3409 -3382
rect 3464 -3428 3534 -3192
rect 3589 -3238 3781 -3233
rect 3589 -3279 3600 -3238
rect 3590 -3341 3600 -3279
rect 3589 -3382 3600 -3341
rect 3770 -3279 3781 -3238
rect 3770 -3341 3780 -3279
rect 3770 -3382 3781 -3341
rect 3589 -3387 3781 -3382
rect 3830 -3428 3884 -3192
rect 882 -3440 975 -3428
rect 882 -4216 935 -3440
rect 969 -4216 975 -3440
rect 882 -4228 975 -4216
rect 1187 -3440 1347 -3428
rect 1187 -4216 1193 -3440
rect 1227 -4216 1307 -3440
rect 1341 -4216 1347 -3440
rect 1187 -4228 1347 -4216
rect 1559 -3440 1719 -3428
rect 1559 -4216 1565 -3440
rect 1599 -4216 1679 -3440
rect 1713 -4216 1719 -3440
rect 1559 -4228 1719 -4216
rect 1931 -3440 2091 -3428
rect 1931 -4216 1937 -3440
rect 1971 -4216 2051 -3440
rect 2085 -4216 2091 -3440
rect 1931 -4228 2091 -4216
rect 2303 -3440 2463 -3428
rect 2303 -4216 2309 -3440
rect 2343 -4216 2423 -3440
rect 2457 -4216 2463 -3440
rect 2303 -4228 2463 -4216
rect 2675 -3440 2835 -3428
rect 2675 -4216 2681 -3440
rect 2715 -4216 2795 -3440
rect 2829 -4216 2835 -3440
rect 2675 -4228 2835 -4216
rect 3047 -3440 3207 -3428
rect 3047 -4216 3053 -3440
rect 3087 -4216 3167 -3440
rect 3201 -4216 3207 -3440
rect 3047 -4228 3207 -4216
rect 3419 -3440 3579 -3428
rect 3419 -4216 3425 -3440
rect 3459 -4216 3539 -3440
rect 3573 -4216 3579 -3440
rect 3419 -4228 3579 -4216
rect 3791 -3440 3884 -3428
rect 3791 -4216 3797 -3440
rect 3831 -4216 3884 -3440
rect 6114 -3477 6186 -3088
rect 5676 -3690 5686 -3528
rect 5846 -3578 5856 -3528
rect 5846 -3584 6042 -3578
rect 5846 -3634 5974 -3584
rect 6030 -3634 6042 -3584
rect 5846 -3640 6042 -3634
rect 5846 -3690 5856 -3640
rect 6114 -3874 6131 -3477
rect 6169 -3874 6186 -3477
rect 6114 -3892 6186 -3874
rect 5676 -4090 5686 -3928
rect 5846 -3978 5856 -3928
rect 5846 -3984 6042 -3978
rect 5846 -4034 5974 -3984
rect 6030 -4034 6042 -3984
rect 5846 -4040 6042 -4034
rect 6114 -4008 6186 -3990
rect 5846 -4090 5856 -4040
rect 3791 -4228 3884 -4216
rect 882 -4464 930 -4228
rect 985 -4274 1177 -4269
rect 985 -4315 996 -4274
rect 986 -4377 996 -4315
rect 985 -4418 996 -4377
rect 1166 -4315 1177 -4274
rect 1166 -4377 1176 -4315
rect 1166 -4418 1177 -4377
rect 985 -4423 1177 -4418
rect 1232 -4464 1302 -4228
rect 1357 -4274 1549 -4269
rect 1357 -4315 1368 -4274
rect 1358 -4377 1368 -4315
rect 1357 -4418 1368 -4377
rect 1538 -4315 1549 -4274
rect 1538 -4377 1548 -4315
rect 1538 -4418 1549 -4377
rect 1357 -4423 1549 -4418
rect 1604 -4464 1674 -4228
rect 1729 -4274 1921 -4269
rect 1729 -4315 1740 -4274
rect 1730 -4377 1740 -4315
rect 1729 -4418 1740 -4377
rect 1910 -4315 1921 -4274
rect 1910 -4377 1920 -4315
rect 1910 -4418 1921 -4377
rect 1729 -4423 1921 -4418
rect 1976 -4464 2046 -4228
rect 2101 -4274 2293 -4269
rect 2101 -4315 2112 -4274
rect 2102 -4377 2112 -4315
rect 2101 -4418 2112 -4377
rect 2282 -4315 2293 -4274
rect 2282 -4377 2292 -4315
rect 2282 -4418 2293 -4377
rect 2101 -4423 2293 -4418
rect 2348 -4464 2418 -4228
rect 2473 -4274 2665 -4269
rect 2473 -4315 2484 -4274
rect 2474 -4377 2484 -4315
rect 2473 -4418 2484 -4377
rect 2654 -4315 2665 -4274
rect 2654 -4377 2664 -4315
rect 2654 -4418 2665 -4377
rect 2473 -4423 2665 -4418
rect 2720 -4464 2790 -4228
rect 2845 -4274 3037 -4269
rect 2845 -4315 2856 -4274
rect 2846 -4377 2856 -4315
rect 2845 -4418 2856 -4377
rect 3026 -4315 3037 -4274
rect 3026 -4377 3036 -4315
rect 3026 -4418 3037 -4377
rect 2845 -4423 3037 -4418
rect 3092 -4464 3162 -4228
rect 3217 -4274 3409 -4269
rect 3217 -4315 3228 -4274
rect 3218 -4377 3228 -4315
rect 3217 -4418 3228 -4377
rect 3398 -4315 3409 -4274
rect 3398 -4377 3408 -4315
rect 3398 -4418 3409 -4377
rect 3217 -4423 3409 -4418
rect 3464 -4464 3534 -4228
rect 3589 -4274 3781 -4269
rect 3589 -4315 3600 -4274
rect 3590 -4377 3600 -4315
rect 3589 -4418 3600 -4377
rect 3770 -4315 3781 -4274
rect 3770 -4377 3780 -4315
rect 3770 -4418 3781 -4377
rect 3589 -4423 3781 -4418
rect 3830 -4464 3884 -4228
rect 882 -4476 975 -4464
rect 882 -5252 935 -4476
rect 969 -5252 975 -4476
rect 882 -5264 975 -5252
rect 1187 -4476 1347 -4464
rect 1187 -5252 1193 -4476
rect 1227 -5252 1307 -4476
rect 1341 -5252 1347 -4476
rect 1187 -5264 1347 -5252
rect 1559 -4476 1719 -4464
rect 1559 -5252 1565 -4476
rect 1599 -5252 1679 -4476
rect 1713 -5252 1719 -4476
rect 1559 -5264 1719 -5252
rect 1931 -4476 2091 -4464
rect 1931 -5252 1937 -4476
rect 1971 -5252 2051 -4476
rect 2085 -5252 2091 -4476
rect 1931 -5264 2091 -5252
rect 2303 -4476 2463 -4464
rect 2303 -5252 2309 -4476
rect 2343 -5252 2423 -4476
rect 2457 -5252 2463 -4476
rect 2303 -5264 2463 -5252
rect 2675 -4476 2835 -4464
rect 2675 -5252 2681 -4476
rect 2715 -5252 2795 -4476
rect 2829 -5252 2835 -4476
rect 2675 -5264 2835 -5252
rect 3047 -4476 3207 -4464
rect 3047 -5252 3053 -4476
rect 3087 -5252 3167 -4476
rect 3201 -5252 3207 -4476
rect 3047 -5264 3207 -5252
rect 3419 -4476 3579 -4464
rect 3419 -5252 3425 -4476
rect 3459 -5252 3539 -4476
rect 3573 -5252 3579 -4476
rect 3419 -5264 3579 -5252
rect 3791 -4476 3884 -4464
rect 3791 -5252 3797 -4476
rect 3831 -5252 3884 -4476
rect 5676 -4490 5686 -4328
rect 5846 -4378 5856 -4328
rect 5846 -4384 6042 -4378
rect 5846 -4434 5974 -4384
rect 6030 -4434 6042 -4384
rect 5846 -4440 6042 -4434
rect 6114 -4405 6131 -4008
rect 6169 -4405 6186 -4008
rect 5846 -4490 5856 -4440
rect 3791 -5264 3884 -5252
rect 986 -5305 996 -5300
rect 985 -5351 996 -5305
rect 1166 -5305 1176 -5300
rect 986 -5354 996 -5351
rect 1166 -5351 1177 -5305
rect 1166 -5354 1176 -5351
rect 1232 -5948 1302 -5264
rect 1358 -5305 1368 -5300
rect 1357 -5351 1368 -5305
rect 1538 -5305 1548 -5300
rect 1730 -5305 1740 -5300
rect 1358 -5354 1368 -5351
rect 1538 -5351 1549 -5305
rect 1729 -5351 1740 -5305
rect 1910 -5305 1920 -5300
rect 1538 -5354 1548 -5351
rect 1730 -5354 1740 -5351
rect 1910 -5351 1921 -5305
rect 1910 -5354 1920 -5351
rect 1976 -5640 2046 -5264
rect 2102 -5305 2112 -5300
rect 2101 -5351 2112 -5305
rect 2282 -5305 2292 -5300
rect 2474 -5305 2484 -5300
rect 2102 -5354 2112 -5351
rect 2282 -5351 2293 -5305
rect 2473 -5351 2484 -5305
rect 2654 -5305 2664 -5300
rect 2282 -5354 2292 -5351
rect 2474 -5354 2484 -5351
rect 2654 -5351 2665 -5305
rect 2654 -5354 2664 -5351
rect 2720 -5640 2790 -5264
rect 2846 -5305 2856 -5300
rect 2845 -5351 2856 -5305
rect 3026 -5305 3036 -5300
rect 3218 -5305 3228 -5300
rect 2846 -5354 2856 -5351
rect 3026 -5351 3037 -5305
rect 3217 -5351 3228 -5305
rect 3398 -5305 3408 -5300
rect 3026 -5354 3036 -5351
rect 3218 -5354 3228 -5351
rect 3398 -5351 3409 -5305
rect 3398 -5354 3408 -5351
rect 1966 -5820 1976 -5640
rect 2790 -5820 2800 -5640
rect 984 -5958 1550 -5948
rect 984 -6004 996 -5958
rect 985 -6009 996 -6004
rect 986 -6014 996 -6009
rect 1166 -6004 1368 -5958
rect 1166 -6009 1177 -6004
rect 1166 -6014 1176 -6009
rect 880 -6041 954 -6040
rect 1232 -6041 1302 -6004
rect 1357 -6009 1368 -6004
rect 1358 -6014 1368 -6009
rect 1538 -6004 1550 -5958
rect 1730 -5963 1740 -5958
rect 1538 -6009 1549 -6004
rect 1729 -6009 1740 -5963
rect 1910 -5963 1920 -5958
rect 1538 -6014 1548 -6009
rect 1730 -6014 1740 -6009
rect 1910 -6009 1921 -5963
rect 1910 -6014 1920 -6009
rect 1604 -6041 1674 -6040
rect 1976 -6041 2046 -5820
rect 2102 -5963 2112 -5958
rect 2101 -6009 2112 -5963
rect 2282 -5963 2292 -5958
rect 2474 -5963 2484 -5958
rect 2102 -6014 2112 -6009
rect 2282 -6009 2293 -5963
rect 2473 -6009 2484 -5963
rect 2654 -5963 2664 -5958
rect 2282 -6014 2292 -6009
rect 2474 -6014 2484 -6009
rect 2654 -6009 2665 -5963
rect 2654 -6014 2664 -6009
rect 2348 -6041 2418 -6040
rect 2720 -6041 2790 -5820
rect 3464 -5948 3534 -5264
rect 3590 -5305 3600 -5300
rect 3589 -5351 3600 -5305
rect 3770 -5305 3780 -5300
rect 3590 -5354 3600 -5351
rect 3770 -5351 3781 -5305
rect 3770 -5354 3780 -5351
rect 4092 -5496 4102 -5224
rect 4384 -5496 4394 -5224
rect 4836 -5496 4846 -5224
rect 5128 -5496 5138 -5224
rect 5580 -5496 5590 -5224
rect 5872 -5496 5882 -5224
rect 6114 -5452 6186 -4405
rect 3216 -5958 3782 -5948
rect 2846 -5963 2856 -5958
rect 2845 -6009 2856 -5963
rect 3026 -5963 3036 -5958
rect 2846 -6014 2856 -6009
rect 3026 -6009 3037 -5963
rect 3216 -6004 3228 -5958
rect 3217 -6009 3228 -6004
rect 3026 -6014 3036 -6009
rect 3218 -6014 3228 -6009
rect 3398 -6004 3600 -5958
rect 3398 -6009 3409 -6004
rect 3398 -6014 3408 -6009
rect 3092 -6041 3162 -6040
rect 3464 -6041 3534 -6004
rect 3589 -6009 3600 -6004
rect 3590 -6014 3600 -6009
rect 3770 -6004 3782 -5958
rect 3962 -5963 3972 -5958
rect 3770 -6009 3781 -6004
rect 3961 -6009 3972 -5963
rect 4142 -5963 4152 -5958
rect 3770 -6014 3780 -6009
rect 3962 -6014 3972 -6009
rect 4142 -6009 4153 -5963
rect 4142 -6014 4152 -6009
rect 3836 -6041 3906 -6040
rect 4208 -6041 4278 -5496
rect 4334 -5963 4344 -5958
rect 4333 -6009 4344 -5963
rect 4514 -5963 4524 -5958
rect 4706 -5963 4716 -5958
rect 4334 -6014 4344 -6009
rect 4514 -6009 4525 -5963
rect 4705 -6009 4716 -5963
rect 4886 -5963 4896 -5958
rect 4514 -6014 4524 -6009
rect 4706 -6014 4716 -6009
rect 4886 -6009 4897 -5963
rect 4886 -6014 4896 -6009
rect 4580 -6041 4650 -6040
rect 4952 -6041 5022 -5496
rect 5078 -5963 5088 -5958
rect 5077 -6009 5088 -5963
rect 5258 -5963 5268 -5958
rect 5450 -5963 5460 -5958
rect 5078 -6014 5088 -6009
rect 5258 -6009 5269 -5963
rect 5449 -6009 5460 -5963
rect 5630 -5963 5640 -5958
rect 5258 -6014 5268 -6009
rect 5450 -6014 5460 -6009
rect 5630 -6009 5641 -5963
rect 5630 -6014 5640 -6009
rect 5324 -6041 5394 -6040
rect 5696 -6041 5766 -5496
rect 6112 -5500 6186 -5452
rect 6324 -5496 6334 -5224
rect 6616 -5496 6626 -5224
rect 7068 -5496 7078 -5224
rect 7360 -5496 7370 -5224
rect 7812 -5496 7822 -5224
rect 8104 -5496 8114 -5224
rect 8556 -5496 8566 -5224
rect 8848 -5496 8858 -5224
rect 9300 -5496 9310 -5224
rect 9592 -5496 9602 -5224
rect 6072 -5512 6186 -5500
rect 5976 -5786 5986 -5512
rect 6264 -5786 6274 -5512
rect 5822 -5963 5832 -5958
rect 5821 -6009 5832 -5963
rect 6002 -5963 6012 -5958
rect 6194 -5963 6204 -5958
rect 5822 -6014 5832 -6009
rect 6002 -6009 6013 -5963
rect 6193 -6009 6204 -5963
rect 6374 -5963 6384 -5958
rect 6002 -6014 6012 -6009
rect 6194 -6014 6204 -6009
rect 6374 -6009 6385 -5963
rect 6374 -6014 6384 -6009
rect 6068 -6041 6138 -6040
rect 6440 -6041 6510 -5496
rect 6566 -5963 6576 -5958
rect 6565 -6009 6576 -5963
rect 6746 -5963 6756 -5958
rect 6938 -5963 6948 -5958
rect 6566 -6014 6576 -6009
rect 6746 -6009 6757 -5963
rect 6937 -6009 6948 -5963
rect 7118 -5963 7128 -5958
rect 6746 -6014 6756 -6009
rect 6938 -6014 6948 -6009
rect 7118 -6009 7129 -5963
rect 7118 -6014 7128 -6009
rect 6812 -6041 6882 -6040
rect 7184 -6041 7254 -5496
rect 7310 -5963 7320 -5958
rect 7309 -6009 7320 -5963
rect 7490 -5963 7500 -5958
rect 7682 -5963 7692 -5958
rect 7310 -6014 7320 -6009
rect 7490 -6009 7501 -5963
rect 7681 -6009 7692 -5963
rect 7862 -5963 7872 -5958
rect 7490 -6014 7500 -6009
rect 7682 -6014 7692 -6009
rect 7862 -6009 7873 -5963
rect 7862 -6014 7872 -6009
rect 7556 -6041 7626 -6040
rect 7928 -6041 7998 -5496
rect 8054 -5963 8064 -5958
rect 8053 -6009 8064 -5963
rect 8234 -5963 8244 -5958
rect 8426 -5963 8436 -5958
rect 8054 -6014 8064 -6009
rect 8234 -6009 8245 -5963
rect 8425 -6009 8436 -5963
rect 8606 -5963 8616 -5958
rect 8234 -6014 8244 -6009
rect 8426 -6014 8436 -6009
rect 8606 -6009 8617 -5963
rect 8606 -6014 8616 -6009
rect 8300 -6041 8370 -6040
rect 8672 -6041 8742 -5496
rect 8798 -5963 8808 -5958
rect 8797 -6009 8808 -5963
rect 8978 -5963 8988 -5958
rect 9170 -5963 9180 -5958
rect 8798 -6014 8808 -6009
rect 8978 -6009 8989 -5963
rect 9169 -6009 9180 -5963
rect 9350 -5963 9360 -5958
rect 8978 -6014 8988 -6009
rect 9170 -6014 9180 -6009
rect 9350 -6009 9361 -5963
rect 9350 -6014 9360 -6009
rect 9044 -6041 9114 -6040
rect 9416 -6041 9486 -5496
rect 9542 -5963 9552 -5958
rect 9541 -6009 9552 -5963
rect 9722 -5963 9732 -5958
rect 9542 -6014 9552 -6009
rect 9722 -6009 9733 -5963
rect 9722 -6014 9732 -6009
rect 9764 -6041 9838 -6028
rect 880 -6053 975 -6041
rect 880 -6229 935 -6053
rect 969 -6229 975 -6053
rect 880 -6241 975 -6229
rect 1187 -6053 1347 -6041
rect 1187 -6229 1193 -6053
rect 1227 -6229 1307 -6053
rect 1341 -6229 1347 -6053
rect 1187 -6241 1347 -6229
rect 1559 -6053 1719 -6041
rect 1559 -6229 1565 -6053
rect 1599 -6229 1679 -6053
rect 1713 -6229 1719 -6053
rect 1559 -6241 1719 -6229
rect 1931 -6053 2091 -6041
rect 1931 -6229 1937 -6053
rect 1971 -6229 2051 -6053
rect 2085 -6229 2091 -6053
rect 1931 -6241 2091 -6229
rect 2303 -6053 2463 -6041
rect 2303 -6229 2309 -6053
rect 2343 -6229 2423 -6053
rect 2457 -6229 2463 -6053
rect 2303 -6241 2463 -6229
rect 2675 -6053 2835 -6041
rect 2675 -6229 2681 -6053
rect 2715 -6229 2795 -6053
rect 2829 -6229 2835 -6053
rect 2675 -6241 2835 -6229
rect 3047 -6053 3207 -6041
rect 3047 -6229 3053 -6053
rect 3087 -6229 3167 -6053
rect 3201 -6229 3207 -6053
rect 3047 -6241 3207 -6229
rect 3419 -6053 3579 -6041
rect 3419 -6229 3425 -6053
rect 3459 -6229 3539 -6053
rect 3573 -6229 3579 -6053
rect 3419 -6241 3579 -6229
rect 3791 -6053 3951 -6041
rect 3791 -6229 3797 -6053
rect 3831 -6229 3911 -6053
rect 3945 -6229 3951 -6053
rect 3791 -6241 3951 -6229
rect 4163 -6053 4323 -6041
rect 4163 -6229 4169 -6053
rect 4203 -6229 4283 -6053
rect 4317 -6229 4323 -6053
rect 4163 -6241 4323 -6229
rect 4535 -6053 4695 -6041
rect 4535 -6229 4541 -6053
rect 4575 -6229 4655 -6053
rect 4689 -6229 4695 -6053
rect 4535 -6241 4695 -6229
rect 4907 -6053 5067 -6041
rect 4907 -6229 4913 -6053
rect 4947 -6229 5027 -6053
rect 5061 -6229 5067 -6053
rect 4907 -6241 5067 -6229
rect 5279 -6053 5439 -6041
rect 5279 -6229 5285 -6053
rect 5319 -6229 5399 -6053
rect 5433 -6229 5439 -6053
rect 5279 -6241 5439 -6229
rect 5651 -6053 5811 -6041
rect 5651 -6229 5657 -6053
rect 5691 -6229 5771 -6053
rect 5805 -6229 5811 -6053
rect 5651 -6241 5811 -6229
rect 6023 -6053 6183 -6041
rect 6023 -6229 6029 -6053
rect 6063 -6229 6143 -6053
rect 6177 -6229 6183 -6053
rect 6023 -6241 6183 -6229
rect 6395 -6053 6555 -6041
rect 6395 -6229 6401 -6053
rect 6435 -6229 6515 -6053
rect 6549 -6229 6555 -6053
rect 6395 -6241 6555 -6229
rect 6767 -6053 6927 -6041
rect 6767 -6229 6773 -6053
rect 6807 -6229 6887 -6053
rect 6921 -6229 6927 -6053
rect 6767 -6241 6927 -6229
rect 7139 -6053 7299 -6041
rect 7139 -6229 7145 -6053
rect 7179 -6229 7259 -6053
rect 7293 -6229 7299 -6053
rect 7139 -6241 7299 -6229
rect 7511 -6053 7671 -6041
rect 7511 -6229 7517 -6053
rect 7551 -6229 7631 -6053
rect 7665 -6229 7671 -6053
rect 7511 -6241 7671 -6229
rect 7883 -6053 8043 -6041
rect 7883 -6229 7889 -6053
rect 7923 -6229 8003 -6053
rect 8037 -6229 8043 -6053
rect 7883 -6241 8043 -6229
rect 8255 -6053 8415 -6041
rect 8255 -6229 8261 -6053
rect 8295 -6229 8375 -6053
rect 8409 -6229 8415 -6053
rect 8255 -6241 8415 -6229
rect 8627 -6053 8787 -6041
rect 8627 -6229 8633 -6053
rect 8667 -6229 8747 -6053
rect 8781 -6229 8787 -6053
rect 8627 -6241 8787 -6229
rect 8999 -6053 9159 -6041
rect 8999 -6229 9005 -6053
rect 9039 -6229 9119 -6053
rect 9153 -6229 9159 -6053
rect 8999 -6241 9159 -6229
rect 9371 -6053 9531 -6041
rect 9371 -6229 9377 -6053
rect 9411 -6229 9491 -6053
rect 9525 -6229 9531 -6053
rect 9371 -6241 9531 -6229
rect 9743 -6053 9838 -6041
rect 9743 -6229 9749 -6053
rect 9783 -6229 9838 -6053
rect 9743 -6241 9838 -6229
rect 880 -6459 954 -6241
rect 1232 -6272 1302 -6241
rect 984 -6278 1550 -6272
rect 984 -6422 996 -6278
rect 1166 -6422 1368 -6278
rect 1538 -6422 1550 -6278
rect 984 -6428 1550 -6422
rect 1232 -6459 1302 -6428
rect 1604 -6459 1674 -6241
rect 1729 -6278 1921 -6273
rect 1729 -6319 1740 -6278
rect 1730 -6381 1740 -6319
rect 1729 -6422 1740 -6381
rect 1910 -6319 1921 -6278
rect 1910 -6381 1920 -6319
rect 1910 -6422 1921 -6381
rect 1729 -6427 1921 -6422
rect 1976 -6459 2046 -6241
rect 2101 -6278 2293 -6273
rect 2101 -6319 2112 -6278
rect 2102 -6381 2112 -6319
rect 2101 -6422 2112 -6381
rect 2282 -6319 2293 -6278
rect 2282 -6381 2292 -6319
rect 2282 -6422 2293 -6381
rect 2101 -6427 2293 -6422
rect 2348 -6459 2418 -6241
rect 2473 -6278 2665 -6273
rect 2473 -6319 2484 -6278
rect 2474 -6381 2484 -6319
rect 2473 -6422 2484 -6381
rect 2654 -6319 2665 -6278
rect 2654 -6381 2664 -6319
rect 2654 -6422 2665 -6381
rect 2473 -6427 2665 -6422
rect 2720 -6459 2790 -6241
rect 2845 -6278 3037 -6273
rect 2845 -6319 2856 -6278
rect 2846 -6381 2856 -6319
rect 2845 -6422 2856 -6381
rect 3026 -6319 3037 -6278
rect 3026 -6381 3036 -6319
rect 3026 -6422 3037 -6381
rect 2845 -6427 3037 -6422
rect 3092 -6459 3162 -6241
rect 3464 -6272 3534 -6241
rect 3216 -6278 3782 -6272
rect 3216 -6422 3228 -6278
rect 3398 -6422 3600 -6278
rect 3770 -6422 3782 -6278
rect 3216 -6428 3782 -6422
rect 3464 -6459 3534 -6428
rect 3836 -6459 3906 -6241
rect 3961 -6278 4153 -6273
rect 3961 -6319 3972 -6278
rect 3962 -6381 3972 -6319
rect 3961 -6422 3972 -6381
rect 4142 -6319 4153 -6278
rect 4142 -6381 4152 -6319
rect 4142 -6422 4153 -6381
rect 3961 -6427 4153 -6422
rect 4208 -6459 4278 -6241
rect 4333 -6278 4525 -6273
rect 4333 -6319 4344 -6278
rect 4334 -6381 4344 -6319
rect 4333 -6422 4344 -6381
rect 4514 -6319 4525 -6278
rect 4514 -6381 4524 -6319
rect 4514 -6422 4525 -6381
rect 4333 -6427 4525 -6422
rect 4580 -6459 4650 -6241
rect 4705 -6278 4897 -6273
rect 4705 -6319 4716 -6278
rect 4706 -6381 4716 -6319
rect 4705 -6422 4716 -6381
rect 4886 -6319 4897 -6278
rect 4886 -6381 4896 -6319
rect 4886 -6422 4897 -6381
rect 4705 -6427 4897 -6422
rect 4952 -6459 5022 -6241
rect 5077 -6278 5269 -6273
rect 5077 -6319 5088 -6278
rect 5078 -6381 5088 -6319
rect 5077 -6422 5088 -6381
rect 5258 -6319 5269 -6278
rect 5258 -6381 5268 -6319
rect 5258 -6422 5269 -6381
rect 5077 -6427 5269 -6422
rect 5324 -6459 5394 -6241
rect 5449 -6278 5641 -6273
rect 5449 -6319 5460 -6278
rect 5450 -6381 5460 -6319
rect 5449 -6422 5460 -6381
rect 5630 -6319 5641 -6278
rect 5630 -6381 5640 -6319
rect 5630 -6422 5641 -6381
rect 5449 -6427 5641 -6422
rect 5696 -6459 5766 -6241
rect 5821 -6278 6013 -6273
rect 5821 -6319 5832 -6278
rect 5822 -6381 5832 -6319
rect 5821 -6422 5832 -6381
rect 6002 -6319 6013 -6278
rect 6002 -6381 6012 -6319
rect 6002 -6422 6013 -6381
rect 5821 -6427 6013 -6422
rect 6068 -6459 6138 -6241
rect 6193 -6278 6385 -6273
rect 6193 -6319 6204 -6278
rect 6194 -6381 6204 -6319
rect 6193 -6422 6204 -6381
rect 6374 -6319 6385 -6278
rect 6374 -6381 6384 -6319
rect 6374 -6422 6385 -6381
rect 6193 -6427 6385 -6422
rect 6440 -6459 6510 -6241
rect 6565 -6278 6757 -6273
rect 6565 -6319 6576 -6278
rect 6566 -6381 6576 -6319
rect 6565 -6422 6576 -6381
rect 6746 -6319 6757 -6278
rect 6746 -6381 6756 -6319
rect 6746 -6422 6757 -6381
rect 6565 -6427 6757 -6422
rect 6812 -6459 6882 -6241
rect 6937 -6278 7129 -6273
rect 6937 -6319 6948 -6278
rect 6938 -6381 6948 -6319
rect 6937 -6422 6948 -6381
rect 7118 -6319 7129 -6278
rect 7118 -6381 7128 -6319
rect 7118 -6422 7129 -6381
rect 6937 -6427 7129 -6422
rect 7184 -6459 7254 -6241
rect 7309 -6278 7501 -6273
rect 7309 -6319 7320 -6278
rect 7310 -6381 7320 -6319
rect 7309 -6422 7320 -6381
rect 7490 -6319 7501 -6278
rect 7490 -6381 7500 -6319
rect 7490 -6422 7501 -6381
rect 7309 -6427 7501 -6422
rect 7556 -6459 7626 -6241
rect 7681 -6278 7873 -6273
rect 7681 -6319 7692 -6278
rect 7682 -6381 7692 -6319
rect 7681 -6422 7692 -6381
rect 7862 -6319 7873 -6278
rect 7862 -6381 7872 -6319
rect 7862 -6422 7873 -6381
rect 7681 -6427 7873 -6422
rect 7928 -6459 7998 -6241
rect 8053 -6278 8245 -6273
rect 8053 -6319 8064 -6278
rect 8054 -6381 8064 -6319
rect 8053 -6422 8064 -6381
rect 8234 -6319 8245 -6278
rect 8234 -6381 8244 -6319
rect 8234 -6422 8245 -6381
rect 8053 -6427 8245 -6422
rect 8300 -6459 8370 -6241
rect 8425 -6278 8617 -6273
rect 8425 -6319 8436 -6278
rect 8426 -6381 8436 -6319
rect 8425 -6422 8436 -6381
rect 8606 -6319 8617 -6278
rect 8606 -6381 8616 -6319
rect 8606 -6422 8617 -6381
rect 8425 -6427 8617 -6422
rect 8672 -6459 8742 -6241
rect 8797 -6278 8989 -6273
rect 8797 -6319 8808 -6278
rect 8798 -6381 8808 -6319
rect 8797 -6422 8808 -6381
rect 8978 -6319 8989 -6278
rect 8978 -6381 8988 -6319
rect 8978 -6422 8989 -6381
rect 8797 -6427 8989 -6422
rect 9044 -6459 9114 -6241
rect 9169 -6278 9361 -6273
rect 9169 -6319 9180 -6278
rect 9170 -6381 9180 -6319
rect 9169 -6422 9180 -6381
rect 9350 -6319 9361 -6278
rect 9350 -6381 9360 -6319
rect 9350 -6422 9361 -6381
rect 9169 -6427 9361 -6422
rect 9416 -6459 9486 -6241
rect 9541 -6278 9733 -6273
rect 9541 -6319 9552 -6278
rect 9542 -6381 9552 -6319
rect 9541 -6422 9552 -6381
rect 9722 -6319 9733 -6278
rect 9722 -6381 9732 -6319
rect 9722 -6422 9733 -6381
rect 9541 -6427 9733 -6422
rect 9764 -6459 9838 -6241
rect 880 -6471 975 -6459
rect 880 -6647 935 -6471
rect 969 -6647 975 -6471
rect 880 -6659 975 -6647
rect 1187 -6471 1347 -6459
rect 1187 -6647 1193 -6471
rect 1227 -6647 1307 -6471
rect 1341 -6647 1347 -6471
rect 1187 -6659 1347 -6647
rect 1559 -6471 1719 -6459
rect 1559 -6647 1565 -6471
rect 1599 -6647 1679 -6471
rect 1713 -6647 1719 -6471
rect 1559 -6659 1719 -6647
rect 1931 -6471 2091 -6459
rect 1931 -6647 1937 -6471
rect 1971 -6647 2051 -6471
rect 2085 -6647 2091 -6471
rect 1931 -6659 2091 -6647
rect 2303 -6471 2463 -6459
rect 2303 -6647 2309 -6471
rect 2343 -6647 2423 -6471
rect 2457 -6647 2463 -6471
rect 2303 -6659 2463 -6647
rect 2675 -6471 2835 -6459
rect 2675 -6647 2681 -6471
rect 2715 -6647 2795 -6471
rect 2829 -6647 2835 -6471
rect 2675 -6659 2835 -6647
rect 3047 -6471 3207 -6459
rect 3047 -6647 3053 -6471
rect 3087 -6647 3167 -6471
rect 3201 -6647 3207 -6471
rect 3047 -6659 3207 -6647
rect 3419 -6471 3579 -6459
rect 3419 -6647 3425 -6471
rect 3459 -6647 3539 -6471
rect 3573 -6647 3579 -6471
rect 3419 -6659 3579 -6647
rect 3791 -6471 3951 -6459
rect 3791 -6647 3797 -6471
rect 3831 -6647 3911 -6471
rect 3945 -6647 3951 -6471
rect 3791 -6659 3951 -6647
rect 4163 -6471 4323 -6459
rect 4163 -6647 4169 -6471
rect 4203 -6647 4283 -6471
rect 4317 -6647 4323 -6471
rect 4163 -6659 4323 -6647
rect 4535 -6471 4695 -6459
rect 4535 -6647 4541 -6471
rect 4575 -6647 4655 -6471
rect 4689 -6647 4695 -6471
rect 4535 -6659 4695 -6647
rect 4907 -6471 5067 -6459
rect 4907 -6647 4913 -6471
rect 4947 -6647 5027 -6471
rect 5061 -6647 5067 -6471
rect 4907 -6659 5067 -6647
rect 5279 -6471 5439 -6459
rect 5279 -6647 5285 -6471
rect 5319 -6647 5399 -6471
rect 5433 -6647 5439 -6471
rect 5279 -6659 5439 -6647
rect 5651 -6471 5811 -6459
rect 5651 -6647 5657 -6471
rect 5691 -6647 5771 -6471
rect 5805 -6647 5811 -6471
rect 5651 -6659 5811 -6647
rect 6023 -6471 6183 -6459
rect 6023 -6647 6029 -6471
rect 6063 -6647 6143 -6471
rect 6177 -6647 6183 -6471
rect 6023 -6659 6183 -6647
rect 6395 -6471 6555 -6459
rect 6395 -6647 6401 -6471
rect 6435 -6647 6515 -6471
rect 6549 -6647 6555 -6471
rect 6395 -6659 6555 -6647
rect 6767 -6471 6927 -6459
rect 6767 -6647 6773 -6471
rect 6807 -6647 6887 -6471
rect 6921 -6647 6927 -6471
rect 6767 -6659 6927 -6647
rect 7139 -6471 7299 -6459
rect 7139 -6647 7145 -6471
rect 7179 -6647 7259 -6471
rect 7293 -6647 7299 -6471
rect 7139 -6659 7299 -6647
rect 7511 -6471 7671 -6459
rect 7511 -6647 7517 -6471
rect 7551 -6647 7631 -6471
rect 7665 -6647 7671 -6471
rect 7511 -6659 7671 -6647
rect 7883 -6471 8043 -6459
rect 7883 -6647 7889 -6471
rect 7923 -6647 8003 -6471
rect 8037 -6647 8043 -6471
rect 7883 -6659 8043 -6647
rect 8255 -6471 8415 -6459
rect 8255 -6647 8261 -6471
rect 8295 -6647 8375 -6471
rect 8409 -6647 8415 -6471
rect 8255 -6659 8415 -6647
rect 8627 -6471 8787 -6459
rect 8627 -6647 8633 -6471
rect 8667 -6647 8747 -6471
rect 8781 -6647 8787 -6471
rect 8627 -6659 8787 -6647
rect 8999 -6471 9159 -6459
rect 8999 -6647 9005 -6471
rect 9039 -6647 9119 -6471
rect 9153 -6647 9159 -6471
rect 8999 -6659 9159 -6647
rect 9371 -6471 9531 -6459
rect 9371 -6647 9377 -6471
rect 9411 -6647 9491 -6471
rect 9525 -6647 9531 -6471
rect 9371 -6659 9531 -6647
rect 9743 -6471 9838 -6459
rect 9743 -6647 9749 -6471
rect 9783 -6647 9838 -6471
rect 9743 -6659 9838 -6647
rect 880 -6877 954 -6659
rect 1232 -6690 1302 -6659
rect 984 -6696 1550 -6690
rect 984 -6840 996 -6696
rect 1166 -6840 1368 -6696
rect 1538 -6840 1550 -6696
rect 984 -6846 1550 -6840
rect 1232 -6877 1302 -6846
rect 1604 -6877 1674 -6659
rect 1729 -6696 1921 -6691
rect 1729 -6737 1740 -6696
rect 1730 -6799 1740 -6737
rect 1729 -6840 1740 -6799
rect 1910 -6737 1921 -6696
rect 1910 -6799 1920 -6737
rect 1910 -6840 1921 -6799
rect 1729 -6845 1921 -6840
rect 1976 -6877 2046 -6659
rect 2101 -6696 2293 -6691
rect 2101 -6737 2112 -6696
rect 2102 -6799 2112 -6737
rect 2101 -6840 2112 -6799
rect 2282 -6737 2293 -6696
rect 2282 -6799 2292 -6737
rect 2282 -6840 2293 -6799
rect 2101 -6845 2293 -6840
rect 2348 -6877 2418 -6659
rect 2473 -6696 2665 -6691
rect 2473 -6737 2484 -6696
rect 2474 -6799 2484 -6737
rect 2473 -6840 2484 -6799
rect 2654 -6737 2665 -6696
rect 2654 -6799 2664 -6737
rect 2654 -6840 2665 -6799
rect 2473 -6845 2665 -6840
rect 2720 -6877 2790 -6659
rect 2845 -6696 3037 -6691
rect 2845 -6737 2856 -6696
rect 2846 -6799 2856 -6737
rect 2845 -6840 2856 -6799
rect 3026 -6737 3037 -6696
rect 3026 -6799 3036 -6737
rect 3026 -6840 3037 -6799
rect 2845 -6845 3037 -6840
rect 3092 -6877 3162 -6659
rect 3464 -6690 3534 -6659
rect 3216 -6696 3782 -6690
rect 3216 -6840 3228 -6696
rect 3398 -6840 3600 -6696
rect 3770 -6840 3782 -6696
rect 3216 -6846 3782 -6840
rect 3464 -6877 3534 -6846
rect 3836 -6877 3906 -6659
rect 3961 -6696 4153 -6691
rect 3961 -6737 3972 -6696
rect 3962 -6799 3972 -6737
rect 3961 -6840 3972 -6799
rect 4142 -6737 4153 -6696
rect 4142 -6799 4152 -6737
rect 4142 -6840 4153 -6799
rect 3961 -6845 4153 -6840
rect 4208 -6877 4278 -6659
rect 4333 -6696 4525 -6691
rect 4333 -6737 4344 -6696
rect 4334 -6799 4344 -6737
rect 4333 -6840 4344 -6799
rect 4514 -6737 4525 -6696
rect 4514 -6799 4524 -6737
rect 4514 -6840 4525 -6799
rect 4333 -6845 4525 -6840
rect 4580 -6877 4650 -6659
rect 4705 -6696 4897 -6691
rect 4705 -6737 4716 -6696
rect 4706 -6799 4716 -6737
rect 4705 -6840 4716 -6799
rect 4886 -6737 4897 -6696
rect 4886 -6799 4896 -6737
rect 4886 -6840 4897 -6799
rect 4705 -6845 4897 -6840
rect 4952 -6877 5022 -6659
rect 5077 -6696 5269 -6691
rect 5077 -6737 5088 -6696
rect 5078 -6799 5088 -6737
rect 5077 -6840 5088 -6799
rect 5258 -6737 5269 -6696
rect 5258 -6799 5268 -6737
rect 5258 -6840 5269 -6799
rect 5077 -6845 5269 -6840
rect 5324 -6877 5394 -6659
rect 5449 -6696 5641 -6691
rect 5449 -6737 5460 -6696
rect 5450 -6799 5460 -6737
rect 5449 -6840 5460 -6799
rect 5630 -6737 5641 -6696
rect 5630 -6799 5640 -6737
rect 5630 -6840 5641 -6799
rect 5449 -6845 5641 -6840
rect 5696 -6877 5766 -6659
rect 5821 -6696 6013 -6691
rect 5821 -6737 5832 -6696
rect 5822 -6799 5832 -6737
rect 5821 -6840 5832 -6799
rect 6002 -6737 6013 -6696
rect 6002 -6799 6012 -6737
rect 6002 -6840 6013 -6799
rect 5821 -6845 6013 -6840
rect 6068 -6877 6138 -6659
rect 6193 -6696 6385 -6691
rect 6193 -6737 6204 -6696
rect 6194 -6799 6204 -6737
rect 6193 -6840 6204 -6799
rect 6374 -6737 6385 -6696
rect 6374 -6799 6384 -6737
rect 6374 -6840 6385 -6799
rect 6193 -6845 6385 -6840
rect 6440 -6877 6510 -6659
rect 6565 -6696 6757 -6691
rect 6565 -6737 6576 -6696
rect 6566 -6799 6576 -6737
rect 6565 -6840 6576 -6799
rect 6746 -6737 6757 -6696
rect 6746 -6799 6756 -6737
rect 6746 -6840 6757 -6799
rect 6565 -6845 6757 -6840
rect 6812 -6877 6882 -6659
rect 6937 -6696 7129 -6691
rect 6937 -6737 6948 -6696
rect 6938 -6799 6948 -6737
rect 6937 -6840 6948 -6799
rect 7118 -6737 7129 -6696
rect 7118 -6799 7128 -6737
rect 7118 -6840 7129 -6799
rect 6937 -6845 7129 -6840
rect 7184 -6877 7254 -6659
rect 7309 -6696 7501 -6691
rect 7309 -6737 7320 -6696
rect 7310 -6799 7320 -6737
rect 7309 -6840 7320 -6799
rect 7490 -6737 7501 -6696
rect 7490 -6799 7500 -6737
rect 7490 -6840 7501 -6799
rect 7309 -6845 7501 -6840
rect 7556 -6877 7626 -6659
rect 7681 -6696 7873 -6691
rect 7681 -6737 7692 -6696
rect 7682 -6799 7692 -6737
rect 7681 -6840 7692 -6799
rect 7862 -6737 7873 -6696
rect 7862 -6799 7872 -6737
rect 7862 -6840 7873 -6799
rect 7681 -6845 7873 -6840
rect 7928 -6877 7998 -6659
rect 8053 -6696 8245 -6691
rect 8053 -6737 8064 -6696
rect 8054 -6799 8064 -6737
rect 8053 -6840 8064 -6799
rect 8234 -6737 8245 -6696
rect 8234 -6799 8244 -6737
rect 8234 -6840 8245 -6799
rect 8053 -6845 8245 -6840
rect 8300 -6877 8370 -6659
rect 8425 -6696 8617 -6691
rect 8425 -6737 8436 -6696
rect 8426 -6799 8436 -6737
rect 8425 -6840 8436 -6799
rect 8606 -6737 8617 -6696
rect 8606 -6799 8616 -6737
rect 8606 -6840 8617 -6799
rect 8425 -6845 8617 -6840
rect 8672 -6877 8742 -6659
rect 8797 -6696 8989 -6691
rect 8797 -6737 8808 -6696
rect 8798 -6799 8808 -6737
rect 8797 -6840 8808 -6799
rect 8978 -6737 8989 -6696
rect 8978 -6799 8988 -6737
rect 8978 -6840 8989 -6799
rect 8797 -6845 8989 -6840
rect 9044 -6877 9114 -6659
rect 9169 -6696 9361 -6691
rect 9169 -6737 9180 -6696
rect 9170 -6799 9180 -6737
rect 9169 -6840 9180 -6799
rect 9350 -6737 9361 -6696
rect 9350 -6799 9360 -6737
rect 9350 -6840 9361 -6799
rect 9169 -6845 9361 -6840
rect 9416 -6877 9486 -6659
rect 9541 -6696 9733 -6691
rect 9541 -6737 9552 -6696
rect 9542 -6799 9552 -6737
rect 9541 -6840 9552 -6799
rect 9722 -6737 9733 -6696
rect 9722 -6799 9732 -6737
rect 9722 -6840 9733 -6799
rect 9541 -6845 9733 -6840
rect 9764 -6877 9838 -6659
rect 880 -6889 975 -6877
rect 880 -7065 935 -6889
rect 969 -7065 975 -6889
rect 880 -7077 975 -7065
rect 1187 -6889 1347 -6877
rect 1187 -7065 1193 -6889
rect 1227 -7065 1307 -6889
rect 1341 -7065 1347 -6889
rect 1187 -7077 1347 -7065
rect 1559 -6889 1719 -6877
rect 1559 -7065 1565 -6889
rect 1599 -7065 1679 -6889
rect 1713 -7065 1719 -6889
rect 1559 -7077 1719 -7065
rect 1931 -6889 2091 -6877
rect 1931 -7065 1937 -6889
rect 1971 -7065 2051 -6889
rect 2085 -7065 2091 -6889
rect 1931 -7077 2091 -7065
rect 2303 -6889 2463 -6877
rect 2303 -7065 2309 -6889
rect 2343 -7065 2423 -6889
rect 2457 -7065 2463 -6889
rect 2303 -7077 2463 -7065
rect 2675 -6889 2835 -6877
rect 2675 -7065 2681 -6889
rect 2715 -7065 2795 -6889
rect 2829 -7065 2835 -6889
rect 2675 -7077 2835 -7065
rect 3047 -6889 3207 -6877
rect 3047 -7065 3053 -6889
rect 3087 -7065 3167 -6889
rect 3201 -7065 3207 -6889
rect 3047 -7077 3207 -7065
rect 3419 -6889 3579 -6877
rect 3419 -7065 3425 -6889
rect 3459 -7065 3539 -6889
rect 3573 -7065 3579 -6889
rect 3419 -7077 3579 -7065
rect 3791 -6889 3951 -6877
rect 3791 -7065 3797 -6889
rect 3831 -7065 3911 -6889
rect 3945 -7065 3951 -6889
rect 3791 -7077 3951 -7065
rect 4163 -6889 4323 -6877
rect 4163 -7065 4169 -6889
rect 4203 -7065 4283 -6889
rect 4317 -7065 4323 -6889
rect 4163 -7077 4323 -7065
rect 4535 -6889 4695 -6877
rect 4535 -7065 4541 -6889
rect 4575 -7065 4655 -6889
rect 4689 -7065 4695 -6889
rect 4535 -7077 4695 -7065
rect 4907 -6889 5067 -6877
rect 4907 -7065 4913 -6889
rect 4947 -7065 5027 -6889
rect 5061 -7065 5067 -6889
rect 4907 -7077 5067 -7065
rect 5279 -6889 5439 -6877
rect 5279 -7065 5285 -6889
rect 5319 -7065 5399 -6889
rect 5433 -7065 5439 -6889
rect 5279 -7077 5439 -7065
rect 5651 -6889 5811 -6877
rect 5651 -7065 5657 -6889
rect 5691 -7065 5771 -6889
rect 5805 -7065 5811 -6889
rect 5651 -7077 5811 -7065
rect 6023 -6889 6183 -6877
rect 6023 -7065 6029 -6889
rect 6063 -7065 6143 -6889
rect 6177 -7065 6183 -6889
rect 6023 -7077 6183 -7065
rect 6395 -6889 6555 -6877
rect 6395 -7065 6401 -6889
rect 6435 -7065 6515 -6889
rect 6549 -7065 6555 -6889
rect 6395 -7077 6555 -7065
rect 6767 -6889 6927 -6877
rect 6767 -7065 6773 -6889
rect 6807 -7065 6887 -6889
rect 6921 -7065 6927 -6889
rect 6767 -7077 6927 -7065
rect 7139 -6889 7299 -6877
rect 7139 -7065 7145 -6889
rect 7179 -7065 7259 -6889
rect 7293 -7065 7299 -6889
rect 7139 -7077 7299 -7065
rect 7511 -6889 7671 -6877
rect 7511 -7065 7517 -6889
rect 7551 -7065 7631 -6889
rect 7665 -7065 7671 -6889
rect 7511 -7077 7671 -7065
rect 7883 -6889 8043 -6877
rect 7883 -7065 7889 -6889
rect 7923 -7065 8003 -6889
rect 8037 -7065 8043 -6889
rect 7883 -7077 8043 -7065
rect 8255 -6889 8415 -6877
rect 8255 -7065 8261 -6889
rect 8295 -7065 8375 -6889
rect 8409 -7065 8415 -6889
rect 8255 -7077 8415 -7065
rect 8627 -6889 8787 -6877
rect 8627 -7065 8633 -6889
rect 8667 -7065 8747 -6889
rect 8781 -7065 8787 -6889
rect 8627 -7077 8787 -7065
rect 8999 -6889 9159 -6877
rect 8999 -7065 9005 -6889
rect 9039 -7065 9119 -6889
rect 9153 -7065 9159 -6889
rect 8999 -7077 9159 -7065
rect 9371 -6889 9531 -6877
rect 9371 -7065 9377 -6889
rect 9411 -7065 9491 -6889
rect 9525 -7065 9531 -6889
rect 9371 -7077 9531 -7065
rect 9743 -6889 9838 -6877
rect 9743 -7065 9749 -6889
rect 9783 -7065 9838 -6889
rect 9743 -7077 9838 -7065
rect 880 -7295 954 -7077
rect 1232 -7108 1302 -7077
rect 984 -7114 1550 -7108
rect 984 -7258 996 -7114
rect 1166 -7258 1368 -7114
rect 1538 -7258 1550 -7114
rect 984 -7264 1550 -7258
rect 1232 -7295 1302 -7264
rect 1604 -7295 1674 -7077
rect 1729 -7114 1921 -7109
rect 1729 -7155 1740 -7114
rect 1730 -7217 1740 -7155
rect 1729 -7258 1740 -7217
rect 1910 -7155 1921 -7114
rect 1910 -7217 1920 -7155
rect 1910 -7258 1921 -7217
rect 1729 -7263 1921 -7258
rect 1976 -7295 2046 -7077
rect 2101 -7114 2293 -7109
rect 2101 -7155 2112 -7114
rect 2102 -7217 2112 -7155
rect 2101 -7258 2112 -7217
rect 2282 -7155 2293 -7114
rect 2282 -7217 2292 -7155
rect 2282 -7258 2293 -7217
rect 2101 -7263 2293 -7258
rect 2348 -7295 2418 -7077
rect 2473 -7114 2665 -7109
rect 2473 -7155 2484 -7114
rect 2474 -7217 2484 -7155
rect 2473 -7258 2484 -7217
rect 2654 -7155 2665 -7114
rect 2654 -7217 2664 -7155
rect 2654 -7258 2665 -7217
rect 2473 -7263 2665 -7258
rect 2720 -7295 2790 -7077
rect 2845 -7114 3037 -7109
rect 2845 -7155 2856 -7114
rect 2846 -7217 2856 -7155
rect 2845 -7258 2856 -7217
rect 3026 -7155 3037 -7114
rect 3026 -7217 3036 -7155
rect 3026 -7258 3037 -7217
rect 2845 -7263 3037 -7258
rect 3092 -7295 3162 -7077
rect 3464 -7108 3534 -7077
rect 3216 -7114 3782 -7108
rect 3216 -7258 3228 -7114
rect 3398 -7258 3600 -7114
rect 3770 -7258 3782 -7114
rect 3216 -7264 3782 -7258
rect 3464 -7295 3534 -7264
rect 3836 -7295 3906 -7077
rect 3961 -7114 4153 -7109
rect 3961 -7155 3972 -7114
rect 3962 -7217 3972 -7155
rect 3961 -7258 3972 -7217
rect 4142 -7155 4153 -7114
rect 4142 -7217 4152 -7155
rect 4142 -7258 4153 -7217
rect 3961 -7263 4153 -7258
rect 4208 -7295 4278 -7077
rect 4333 -7114 4525 -7109
rect 4333 -7155 4344 -7114
rect 4334 -7217 4344 -7155
rect 4333 -7258 4344 -7217
rect 4514 -7155 4525 -7114
rect 4514 -7217 4524 -7155
rect 4514 -7258 4525 -7217
rect 4333 -7263 4525 -7258
rect 4580 -7295 4650 -7077
rect 4705 -7114 4897 -7109
rect 4705 -7155 4716 -7114
rect 4706 -7217 4716 -7155
rect 4705 -7258 4716 -7217
rect 4886 -7155 4897 -7114
rect 4886 -7217 4896 -7155
rect 4886 -7258 4897 -7217
rect 4705 -7263 4897 -7258
rect 4952 -7295 5022 -7077
rect 5077 -7114 5269 -7109
rect 5077 -7155 5088 -7114
rect 5078 -7217 5088 -7155
rect 5077 -7258 5088 -7217
rect 5258 -7155 5269 -7114
rect 5258 -7217 5268 -7155
rect 5258 -7258 5269 -7217
rect 5077 -7263 5269 -7258
rect 5324 -7295 5394 -7077
rect 5449 -7114 5641 -7109
rect 5449 -7155 5460 -7114
rect 5450 -7217 5460 -7155
rect 5449 -7258 5460 -7217
rect 5630 -7155 5641 -7114
rect 5630 -7217 5640 -7155
rect 5630 -7258 5641 -7217
rect 5449 -7263 5641 -7258
rect 5696 -7295 5766 -7077
rect 5821 -7114 6013 -7109
rect 5821 -7155 5832 -7114
rect 5822 -7217 5832 -7155
rect 5821 -7258 5832 -7217
rect 6002 -7155 6013 -7114
rect 6002 -7217 6012 -7155
rect 6002 -7258 6013 -7217
rect 5821 -7263 6013 -7258
rect 6068 -7295 6138 -7077
rect 6193 -7114 6385 -7109
rect 6193 -7155 6204 -7114
rect 6194 -7217 6204 -7155
rect 6193 -7258 6204 -7217
rect 6374 -7155 6385 -7114
rect 6374 -7217 6384 -7155
rect 6374 -7258 6385 -7217
rect 6193 -7263 6385 -7258
rect 6440 -7295 6510 -7077
rect 6565 -7114 6757 -7109
rect 6565 -7155 6576 -7114
rect 6566 -7217 6576 -7155
rect 6565 -7258 6576 -7217
rect 6746 -7155 6757 -7114
rect 6746 -7217 6756 -7155
rect 6746 -7258 6757 -7217
rect 6565 -7263 6757 -7258
rect 6812 -7295 6882 -7077
rect 6937 -7114 7129 -7109
rect 6937 -7155 6948 -7114
rect 6938 -7217 6948 -7155
rect 6937 -7258 6948 -7217
rect 7118 -7155 7129 -7114
rect 7118 -7217 7128 -7155
rect 7118 -7258 7129 -7217
rect 6937 -7263 7129 -7258
rect 7184 -7295 7254 -7077
rect 7309 -7114 7501 -7109
rect 7309 -7155 7320 -7114
rect 7310 -7217 7320 -7155
rect 7309 -7258 7320 -7217
rect 7490 -7155 7501 -7114
rect 7490 -7217 7500 -7155
rect 7490 -7258 7501 -7217
rect 7309 -7263 7501 -7258
rect 7556 -7295 7626 -7077
rect 7681 -7114 7873 -7109
rect 7681 -7155 7692 -7114
rect 7682 -7217 7692 -7155
rect 7681 -7258 7692 -7217
rect 7862 -7155 7873 -7114
rect 7862 -7217 7872 -7155
rect 7862 -7258 7873 -7217
rect 7681 -7263 7873 -7258
rect 7928 -7295 7998 -7077
rect 8053 -7114 8245 -7109
rect 8053 -7155 8064 -7114
rect 8054 -7217 8064 -7155
rect 8053 -7258 8064 -7217
rect 8234 -7155 8245 -7114
rect 8234 -7217 8244 -7155
rect 8234 -7258 8245 -7217
rect 8053 -7263 8245 -7258
rect 8300 -7295 8370 -7077
rect 8425 -7114 8617 -7109
rect 8425 -7155 8436 -7114
rect 8426 -7217 8436 -7155
rect 8425 -7258 8436 -7217
rect 8606 -7155 8617 -7114
rect 8606 -7217 8616 -7155
rect 8606 -7258 8617 -7217
rect 8425 -7263 8617 -7258
rect 8672 -7295 8742 -7077
rect 8797 -7114 8989 -7109
rect 8797 -7155 8808 -7114
rect 8798 -7217 8808 -7155
rect 8797 -7258 8808 -7217
rect 8978 -7155 8989 -7114
rect 8978 -7217 8988 -7155
rect 8978 -7258 8989 -7217
rect 8797 -7263 8989 -7258
rect 9044 -7295 9114 -7077
rect 9169 -7114 9361 -7109
rect 9169 -7155 9180 -7114
rect 9170 -7217 9180 -7155
rect 9169 -7258 9180 -7217
rect 9350 -7155 9361 -7114
rect 9350 -7217 9360 -7155
rect 9350 -7258 9361 -7217
rect 9169 -7263 9361 -7258
rect 9416 -7295 9486 -7077
rect 9541 -7114 9733 -7109
rect 9541 -7155 9552 -7114
rect 9542 -7217 9552 -7155
rect 9541 -7258 9552 -7217
rect 9722 -7155 9733 -7114
rect 9722 -7217 9732 -7155
rect 9722 -7258 9733 -7217
rect 9541 -7263 9733 -7258
rect 9764 -7295 9838 -7077
rect 880 -7307 975 -7295
rect 880 -7483 935 -7307
rect 969 -7483 975 -7307
rect 880 -7495 975 -7483
rect 1187 -7307 1347 -7295
rect 1187 -7483 1193 -7307
rect 1227 -7483 1307 -7307
rect 1341 -7483 1347 -7307
rect 1187 -7495 1347 -7483
rect 1559 -7307 1719 -7295
rect 1559 -7483 1565 -7307
rect 1599 -7483 1679 -7307
rect 1713 -7483 1719 -7307
rect 1559 -7495 1719 -7483
rect 1931 -7307 2091 -7295
rect 1931 -7483 1937 -7307
rect 1971 -7483 2051 -7307
rect 2085 -7483 2091 -7307
rect 1931 -7495 2091 -7483
rect 2303 -7307 2463 -7295
rect 2303 -7483 2309 -7307
rect 2343 -7483 2423 -7307
rect 2457 -7483 2463 -7307
rect 2303 -7495 2463 -7483
rect 2675 -7307 2835 -7295
rect 2675 -7483 2681 -7307
rect 2715 -7483 2795 -7307
rect 2829 -7483 2835 -7307
rect 2675 -7495 2835 -7483
rect 3047 -7307 3207 -7295
rect 3047 -7483 3053 -7307
rect 3087 -7483 3167 -7307
rect 3201 -7483 3207 -7307
rect 3047 -7495 3207 -7483
rect 3419 -7307 3579 -7295
rect 3419 -7483 3425 -7307
rect 3459 -7483 3539 -7307
rect 3573 -7483 3579 -7307
rect 3419 -7495 3579 -7483
rect 3791 -7307 3951 -7295
rect 3791 -7483 3797 -7307
rect 3831 -7483 3911 -7307
rect 3945 -7483 3951 -7307
rect 3791 -7495 3951 -7483
rect 4163 -7307 4323 -7295
rect 4163 -7483 4169 -7307
rect 4203 -7483 4283 -7307
rect 4317 -7483 4323 -7307
rect 4163 -7495 4323 -7483
rect 4535 -7307 4695 -7295
rect 4535 -7483 4541 -7307
rect 4575 -7483 4655 -7307
rect 4689 -7483 4695 -7307
rect 4535 -7495 4695 -7483
rect 4907 -7307 5067 -7295
rect 4907 -7483 4913 -7307
rect 4947 -7483 5027 -7307
rect 5061 -7483 5067 -7307
rect 4907 -7495 5067 -7483
rect 5279 -7307 5439 -7295
rect 5279 -7483 5285 -7307
rect 5319 -7483 5399 -7307
rect 5433 -7483 5439 -7307
rect 5279 -7495 5439 -7483
rect 5651 -7307 5811 -7295
rect 5651 -7483 5657 -7307
rect 5691 -7483 5771 -7307
rect 5805 -7483 5811 -7307
rect 5651 -7495 5811 -7483
rect 6023 -7307 6183 -7295
rect 6023 -7483 6029 -7307
rect 6063 -7483 6143 -7307
rect 6177 -7483 6183 -7307
rect 6023 -7495 6183 -7483
rect 6395 -7307 6555 -7295
rect 6395 -7483 6401 -7307
rect 6435 -7483 6515 -7307
rect 6549 -7483 6555 -7307
rect 6395 -7495 6555 -7483
rect 6767 -7307 6927 -7295
rect 6767 -7483 6773 -7307
rect 6807 -7483 6887 -7307
rect 6921 -7483 6927 -7307
rect 6767 -7495 6927 -7483
rect 7139 -7307 7299 -7295
rect 7139 -7483 7145 -7307
rect 7179 -7483 7259 -7307
rect 7293 -7483 7299 -7307
rect 7139 -7495 7299 -7483
rect 7511 -7307 7671 -7295
rect 7511 -7483 7517 -7307
rect 7551 -7483 7631 -7307
rect 7665 -7483 7671 -7307
rect 7511 -7495 7671 -7483
rect 7883 -7307 8043 -7295
rect 7883 -7483 7889 -7307
rect 7923 -7483 8003 -7307
rect 8037 -7483 8043 -7307
rect 7883 -7495 8043 -7483
rect 8255 -7307 8415 -7295
rect 8255 -7483 8261 -7307
rect 8295 -7483 8375 -7307
rect 8409 -7483 8415 -7307
rect 8255 -7495 8415 -7483
rect 8627 -7307 8787 -7295
rect 8627 -7483 8633 -7307
rect 8667 -7483 8747 -7307
rect 8781 -7483 8787 -7307
rect 8627 -7495 8787 -7483
rect 8999 -7307 9159 -7295
rect 8999 -7483 9005 -7307
rect 9039 -7483 9119 -7307
rect 9153 -7483 9159 -7307
rect 8999 -7495 9159 -7483
rect 9371 -7307 9531 -7295
rect 9371 -7483 9377 -7307
rect 9411 -7483 9491 -7307
rect 9525 -7483 9531 -7307
rect 9371 -7495 9531 -7483
rect 9743 -7307 9838 -7295
rect 9743 -7483 9749 -7307
rect 9783 -7483 9838 -7307
rect 9743 -7495 9838 -7483
rect 880 -7618 954 -7495
rect 986 -7527 996 -7522
rect 985 -7532 996 -7527
rect 984 -7578 996 -7532
rect 1166 -7527 1176 -7522
rect 1166 -7532 1177 -7527
rect 1232 -7532 1302 -7495
rect 1604 -7496 1674 -7495
rect 1976 -7496 2046 -7495
rect 2348 -7496 2418 -7495
rect 2720 -7496 2790 -7495
rect 3092 -7496 3162 -7495
rect 1358 -7527 1368 -7522
rect 1357 -7532 1368 -7527
rect 1166 -7578 1368 -7532
rect 1538 -7527 1548 -7522
rect 1538 -7532 1549 -7527
rect 1538 -7578 1550 -7532
rect 984 -7590 1550 -7578
rect 1610 -7610 1668 -7496
rect 1730 -7527 1740 -7522
rect 1729 -7573 1740 -7527
rect 1910 -7527 1920 -7522
rect 2102 -7527 2112 -7522
rect 1730 -7578 1740 -7573
rect 1910 -7573 1921 -7527
rect 2101 -7573 2112 -7527
rect 2282 -7527 2292 -7522
rect 1910 -7578 1920 -7573
rect 2102 -7578 2112 -7573
rect 2282 -7573 2293 -7527
rect 2282 -7578 2292 -7573
rect 2354 -7610 2412 -7496
rect 2474 -7527 2484 -7522
rect 2473 -7573 2484 -7527
rect 2654 -7527 2664 -7522
rect 2846 -7527 2856 -7522
rect 2474 -7578 2484 -7573
rect 2654 -7573 2665 -7527
rect 2845 -7573 2856 -7527
rect 3026 -7527 3036 -7522
rect 2654 -7578 2664 -7573
rect 2846 -7578 2856 -7573
rect 3026 -7573 3037 -7527
rect 3026 -7578 3036 -7573
rect 3098 -7610 3156 -7496
rect 3218 -7527 3228 -7522
rect 3217 -7532 3228 -7527
rect 3216 -7578 3228 -7532
rect 3398 -7527 3408 -7522
rect 3398 -7532 3409 -7527
rect 3464 -7532 3534 -7495
rect 3836 -7496 3906 -7495
rect 4208 -7496 4278 -7495
rect 4580 -7496 4650 -7495
rect 4952 -7496 5022 -7495
rect 5324 -7496 5394 -7495
rect 5696 -7496 5766 -7495
rect 6068 -7496 6138 -7495
rect 6440 -7496 6510 -7495
rect 6812 -7496 6882 -7495
rect 7184 -7496 7254 -7495
rect 7556 -7496 7626 -7495
rect 7928 -7496 7998 -7495
rect 8300 -7496 8370 -7495
rect 8672 -7496 8742 -7495
rect 9044 -7496 9114 -7495
rect 9416 -7496 9486 -7495
rect 3590 -7527 3600 -7522
rect 3589 -7532 3600 -7527
rect 3398 -7578 3600 -7532
rect 3770 -7527 3780 -7522
rect 3770 -7532 3781 -7527
rect 3770 -7578 3782 -7532
rect 3216 -7590 3782 -7578
rect 3842 -7610 3900 -7496
rect 3962 -7527 3972 -7522
rect 3961 -7573 3972 -7527
rect 4142 -7527 4152 -7522
rect 4334 -7527 4344 -7522
rect 3962 -7578 3972 -7573
rect 4142 -7573 4153 -7527
rect 4333 -7573 4344 -7527
rect 4514 -7527 4524 -7522
rect 4142 -7578 4152 -7573
rect 4334 -7578 4344 -7573
rect 4514 -7573 4525 -7527
rect 4514 -7578 4524 -7573
rect 4586 -7610 4644 -7496
rect 4706 -7527 4716 -7522
rect 4705 -7573 4716 -7527
rect 4886 -7527 4896 -7522
rect 5078 -7527 5088 -7522
rect 4706 -7578 4716 -7573
rect 4886 -7573 4897 -7527
rect 5077 -7573 5088 -7527
rect 5258 -7527 5268 -7522
rect 4886 -7578 4896 -7573
rect 5078 -7578 5088 -7573
rect 5258 -7573 5269 -7527
rect 5258 -7578 5268 -7573
rect 5330 -7610 5388 -7496
rect 5450 -7527 5460 -7522
rect 5449 -7573 5460 -7527
rect 5630 -7527 5640 -7522
rect 5822 -7527 5832 -7522
rect 5450 -7578 5460 -7573
rect 5630 -7573 5641 -7527
rect 5821 -7573 5832 -7527
rect 6002 -7527 6012 -7522
rect 5630 -7578 5640 -7573
rect 5822 -7578 5832 -7573
rect 6002 -7573 6013 -7527
rect 6002 -7578 6012 -7573
rect 6074 -7610 6132 -7496
rect 6194 -7527 6204 -7522
rect 6193 -7573 6204 -7527
rect 6374 -7527 6384 -7522
rect 6566 -7527 6576 -7522
rect 6194 -7578 6204 -7573
rect 6374 -7573 6385 -7527
rect 6565 -7573 6576 -7527
rect 6746 -7527 6756 -7522
rect 6374 -7578 6384 -7573
rect 6566 -7578 6576 -7573
rect 6746 -7573 6757 -7527
rect 6746 -7578 6756 -7573
rect 6818 -7610 6876 -7496
rect 6938 -7527 6948 -7522
rect 6937 -7573 6948 -7527
rect 7118 -7527 7128 -7522
rect 7310 -7527 7320 -7522
rect 6938 -7578 6948 -7573
rect 7118 -7573 7129 -7527
rect 7309 -7573 7320 -7527
rect 7490 -7527 7500 -7522
rect 7118 -7578 7128 -7573
rect 7310 -7578 7320 -7573
rect 7490 -7573 7501 -7527
rect 7490 -7578 7500 -7573
rect 7562 -7610 7620 -7496
rect 7682 -7527 7692 -7522
rect 7681 -7573 7692 -7527
rect 7862 -7527 7872 -7522
rect 8054 -7527 8064 -7522
rect 7682 -7578 7692 -7573
rect 7862 -7573 7873 -7527
rect 8053 -7573 8064 -7527
rect 8234 -7527 8244 -7522
rect 7862 -7578 7872 -7573
rect 8054 -7578 8064 -7573
rect 8234 -7573 8245 -7527
rect 8234 -7578 8244 -7573
rect 8306 -7610 8364 -7496
rect 8426 -7527 8436 -7522
rect 8425 -7573 8436 -7527
rect 8606 -7527 8616 -7522
rect 8798 -7527 8808 -7522
rect 8426 -7578 8436 -7573
rect 8606 -7573 8617 -7527
rect 8797 -7573 8808 -7527
rect 8978 -7527 8988 -7522
rect 8606 -7578 8616 -7573
rect 8798 -7578 8808 -7573
rect 8978 -7573 8989 -7527
rect 8978 -7578 8988 -7573
rect 9050 -7610 9108 -7496
rect 9170 -7527 9180 -7522
rect 9169 -7573 9180 -7527
rect 9350 -7527 9360 -7522
rect 9542 -7527 9552 -7522
rect 9170 -7578 9180 -7573
rect 9350 -7573 9361 -7527
rect 9541 -7573 9552 -7527
rect 9722 -7527 9732 -7522
rect 9350 -7578 9360 -7573
rect 9542 -7578 9552 -7573
rect 9722 -7573 9733 -7527
rect 9722 -7578 9732 -7573
rect 1592 -7616 1686 -7610
rect 880 -7624 1018 -7618
rect 880 -7694 936 -7624
rect 1006 -7694 1018 -7624
rect 1592 -7686 1604 -7616
rect 1674 -7686 1686 -7616
rect 1592 -7692 1686 -7686
rect 2336 -7616 2430 -7610
rect 2336 -7686 2348 -7616
rect 2418 -7686 2430 -7616
rect 2336 -7692 2430 -7686
rect 3080 -7616 3174 -7610
rect 3080 -7686 3092 -7616
rect 3162 -7686 3174 -7616
rect 3080 -7692 3174 -7686
rect 3824 -7616 3918 -7610
rect 3824 -7686 3836 -7616
rect 3906 -7686 3918 -7616
rect 3824 -7692 3918 -7686
rect 4568 -7616 4662 -7610
rect 4568 -7686 4580 -7616
rect 4650 -7686 4662 -7616
rect 4568 -7692 4662 -7686
rect 5312 -7616 5406 -7610
rect 5312 -7686 5324 -7616
rect 5394 -7686 5406 -7616
rect 5312 -7692 5406 -7686
rect 6056 -7616 6150 -7610
rect 6056 -7686 6068 -7616
rect 6138 -7686 6150 -7616
rect 6056 -7692 6150 -7686
rect 6800 -7616 6894 -7610
rect 6800 -7686 6812 -7616
rect 6882 -7686 6894 -7616
rect 6800 -7692 6894 -7686
rect 7544 -7616 7638 -7610
rect 7544 -7686 7556 -7616
rect 7626 -7686 7638 -7616
rect 7544 -7692 7638 -7686
rect 8288 -7616 8382 -7610
rect 8288 -7686 8300 -7616
rect 8370 -7686 8382 -7616
rect 8288 -7692 8382 -7686
rect 9032 -7616 9126 -7610
rect 9764 -7614 9838 -7495
rect 9032 -7686 9044 -7616
rect 9114 -7686 9126 -7616
rect 9032 -7692 9126 -7686
rect 9694 -7620 9838 -7614
rect 9694 -7690 9706 -7620
rect 9776 -7690 9838 -7620
rect 880 -7700 1018 -7694
rect 880 -7732 954 -7700
rect 1610 -7732 1668 -7692
rect 2354 -7732 2412 -7692
rect 3098 -7732 3156 -7692
rect 3842 -7732 3900 -7692
rect 4586 -7732 4644 -7692
rect 5330 -7732 5388 -7692
rect 6074 -7732 6132 -7692
rect 6818 -7732 6876 -7692
rect 7562 -7732 7620 -7692
rect 8306 -7732 8364 -7692
rect 9050 -7732 9108 -7692
rect 9694 -7696 9838 -7690
rect 9764 -7720 9838 -7696
rect 9764 -7732 9852 -7720
rect 806 -7932 816 -7732
rect 1016 -7932 1026 -7732
rect 1530 -7932 1540 -7732
rect 1740 -7932 1750 -7732
rect 2274 -7932 2284 -7732
rect 2484 -7932 2494 -7732
rect 3018 -7932 3028 -7732
rect 3228 -7932 3238 -7732
rect 3762 -7932 3772 -7732
rect 3972 -7932 3982 -7732
rect 4506 -7932 4516 -7732
rect 4716 -7932 4726 -7732
rect 5250 -7932 5260 -7732
rect 5460 -7932 5470 -7732
rect 5994 -7932 6004 -7732
rect 6204 -7932 6214 -7732
rect 6738 -7932 6748 -7732
rect 6948 -7932 6958 -7732
rect 7482 -7932 7492 -7732
rect 7692 -7932 7702 -7732
rect 8226 -7932 8236 -7732
rect 8436 -7932 8446 -7732
rect 8970 -7932 8980 -7732
rect 9180 -7932 9190 -7732
rect 9714 -7932 9724 -7732
rect 9924 -7932 9934 -7732
<< via1 >>
rect -322 1314 -122 1514
rect 422 1314 622 1514
rect 1166 1314 1366 1514
rect 1910 1314 2110 1514
rect 2654 1314 2854 1514
rect 3398 1314 3598 1514
rect 4142 1314 4342 1514
rect 4886 1314 5086 1514
rect 5258 1314 5458 1514
rect 6002 1314 6202 1514
rect 6746 1314 6946 1514
rect 7490 1314 7690 1514
rect 8234 1314 8434 1514
rect 8978 1314 9178 1514
rect 9722 1314 9922 1514
rect 10466 1314 10666 1514
rect 11210 1314 11410 1514
rect -492 1113 -322 1126
rect -492 1079 -491 1113
rect -491 1079 -323 1113
rect -323 1079 -322 1113
rect -492 1066 -322 1079
rect -120 1113 50 1126
rect -120 1079 -119 1113
rect -119 1079 49 1113
rect 49 1079 50 1113
rect -120 1066 50 1079
rect 252 1113 422 1126
rect 252 1079 253 1113
rect 253 1079 421 1113
rect 421 1079 422 1113
rect 252 1066 422 1079
rect 624 1113 794 1126
rect 624 1079 625 1113
rect 625 1079 793 1113
rect 793 1079 794 1113
rect 624 1066 794 1079
rect 996 1113 1166 1126
rect 996 1079 997 1113
rect 997 1079 1165 1113
rect 1165 1079 1166 1113
rect 996 1066 1166 1079
rect 1368 1113 1538 1126
rect 1368 1079 1369 1113
rect 1369 1079 1537 1113
rect 1537 1079 1538 1113
rect 1368 1066 1538 1079
rect 1740 1113 1910 1126
rect 1740 1079 1741 1113
rect 1741 1079 1909 1113
rect 1909 1079 1910 1113
rect 1740 1066 1910 1079
rect 2112 1113 2282 1126
rect 2112 1079 2113 1113
rect 2113 1079 2281 1113
rect 2281 1079 2282 1113
rect 2112 1066 2282 1079
rect 2484 1113 2654 1126
rect 2484 1079 2485 1113
rect 2485 1079 2653 1113
rect 2653 1079 2654 1113
rect 2484 1066 2654 1079
rect 2856 1113 3026 1126
rect 2856 1079 2857 1113
rect 2857 1079 3025 1113
rect 3025 1079 3026 1113
rect 2856 1066 3026 1079
rect 3228 1113 3398 1126
rect 3228 1079 3229 1113
rect 3229 1079 3397 1113
rect 3397 1079 3398 1113
rect 3228 1066 3398 1079
rect 3600 1113 3770 1126
rect 3600 1079 3601 1113
rect 3601 1079 3769 1113
rect 3769 1079 3770 1113
rect 3600 1066 3770 1079
rect 3972 1113 4142 1126
rect 3972 1079 3973 1113
rect 3973 1079 4141 1113
rect 4141 1079 4142 1113
rect 3972 1066 4142 1079
rect 4344 1113 4514 1126
rect 4344 1079 4345 1113
rect 4345 1079 4513 1113
rect 4513 1079 4514 1113
rect 4344 1066 4514 1079
rect 4716 1113 4886 1126
rect 4716 1079 4717 1113
rect 4717 1079 4885 1113
rect 4885 1079 4886 1113
rect 4716 1066 4886 1079
rect 5088 1113 5258 1126
rect 5088 1079 5089 1113
rect 5089 1079 5257 1113
rect 5257 1079 5258 1113
rect 5088 1066 5258 1079
rect -492 585 -322 586
rect -492 551 -491 585
rect -491 551 -323 585
rect -323 551 -322 585
rect -492 477 -322 551
rect -492 443 -491 477
rect -491 443 -323 477
rect -323 443 -322 477
rect -492 442 -322 443
rect -120 585 50 586
rect -120 551 -119 585
rect -119 551 49 585
rect 49 551 50 585
rect -120 477 50 551
rect -120 443 -119 477
rect -119 443 49 477
rect 49 443 50 477
rect -120 442 50 443
rect 252 585 422 586
rect 252 551 253 585
rect 253 551 421 585
rect 421 551 422 585
rect 252 477 422 551
rect 252 443 253 477
rect 253 443 421 477
rect 421 443 422 477
rect 252 442 422 443
rect 624 585 794 586
rect 624 551 625 585
rect 625 551 793 585
rect 793 551 794 585
rect 624 477 794 551
rect 624 443 625 477
rect 625 443 793 477
rect 793 443 794 477
rect 624 442 794 443
rect 996 585 1166 586
rect 996 551 997 585
rect 997 551 1165 585
rect 1165 551 1166 585
rect 996 477 1166 551
rect 996 443 997 477
rect 997 443 1165 477
rect 1165 443 1166 477
rect 996 442 1166 443
rect 1368 585 1538 586
rect 1368 551 1369 585
rect 1369 551 1537 585
rect 1537 551 1538 585
rect 1368 477 1538 551
rect 1368 443 1369 477
rect 1369 443 1537 477
rect 1537 443 1538 477
rect 1368 442 1538 443
rect 1740 585 1910 586
rect 1740 551 1741 585
rect 1741 551 1909 585
rect 1909 551 1910 585
rect 1740 477 1910 551
rect 1740 443 1741 477
rect 1741 443 1909 477
rect 1909 443 1910 477
rect 1740 442 1910 443
rect 2112 585 2282 586
rect 2112 551 2113 585
rect 2113 551 2281 585
rect 2281 551 2282 585
rect 2112 477 2282 551
rect 2112 443 2113 477
rect 2113 443 2281 477
rect 2281 443 2282 477
rect 2112 442 2282 443
rect 2484 585 2654 586
rect 2484 551 2485 585
rect 2485 551 2653 585
rect 2653 551 2654 585
rect 2484 477 2654 551
rect 2484 443 2485 477
rect 2485 443 2653 477
rect 2653 443 2654 477
rect 2484 442 2654 443
rect 2856 585 3026 586
rect 2856 551 2857 585
rect 2857 551 3025 585
rect 3025 551 3026 585
rect 2856 477 3026 551
rect 2856 443 2857 477
rect 2857 443 3025 477
rect 3025 443 3026 477
rect 2856 442 3026 443
rect 3228 585 3398 586
rect 3228 551 3229 585
rect 3229 551 3397 585
rect 3397 551 3398 585
rect 3228 477 3398 551
rect 3228 443 3229 477
rect 3229 443 3397 477
rect 3397 443 3398 477
rect 3228 442 3398 443
rect 3600 585 3770 586
rect 3600 551 3601 585
rect 3601 551 3769 585
rect 3769 551 3770 585
rect 3600 477 3770 551
rect 3600 443 3601 477
rect 3601 443 3769 477
rect 3769 443 3770 477
rect 3600 442 3770 443
rect 3972 585 4142 586
rect 3972 551 3973 585
rect 3973 551 4141 585
rect 4141 551 4142 585
rect 3972 477 4142 551
rect 3972 443 3973 477
rect 3973 443 4141 477
rect 4141 443 4142 477
rect 3972 442 4142 443
rect 4344 585 4514 586
rect 4344 551 4345 585
rect 4345 551 4513 585
rect 4513 551 4514 585
rect 4344 477 4514 551
rect 4344 443 4345 477
rect 4345 443 4513 477
rect 4513 443 4514 477
rect 4344 442 4514 443
rect 4716 585 4886 586
rect 4716 551 4717 585
rect 4717 551 4885 585
rect 4885 551 4886 585
rect 4716 477 4886 551
rect 4716 443 4717 477
rect 4717 443 4885 477
rect 4885 443 4886 477
rect 4716 442 4886 443
rect 5088 585 5258 586
rect 5088 551 5089 585
rect 5089 551 5257 585
rect 5257 551 5258 585
rect 5088 477 5258 551
rect 5088 443 5089 477
rect 5089 443 5257 477
rect 5257 443 5258 477
rect 5088 442 5258 443
rect -492 -51 -322 -50
rect -492 -85 -491 -51
rect -491 -85 -323 -51
rect -323 -85 -322 -51
rect -492 -159 -322 -85
rect -492 -193 -491 -159
rect -491 -193 -323 -159
rect -323 -193 -322 -159
rect -492 -194 -322 -193
rect -120 -51 50 -50
rect -120 -85 -119 -51
rect -119 -85 49 -51
rect 49 -85 50 -51
rect -120 -159 50 -85
rect -120 -193 -119 -159
rect -119 -193 49 -159
rect 49 -193 50 -159
rect -120 -194 50 -193
rect 252 -51 422 -50
rect 252 -85 253 -51
rect 253 -85 421 -51
rect 421 -85 422 -51
rect 252 -159 422 -85
rect 252 -193 253 -159
rect 253 -193 421 -159
rect 421 -193 422 -159
rect 252 -194 422 -193
rect 624 -51 794 -50
rect 624 -85 625 -51
rect 625 -85 793 -51
rect 793 -85 794 -51
rect 624 -159 794 -85
rect 624 -193 625 -159
rect 625 -193 793 -159
rect 793 -193 794 -159
rect 624 -194 794 -193
rect 996 -51 1166 -50
rect 996 -85 997 -51
rect 997 -85 1165 -51
rect 1165 -85 1166 -51
rect 996 -159 1166 -85
rect 996 -193 997 -159
rect 997 -193 1165 -159
rect 1165 -193 1166 -159
rect 996 -194 1166 -193
rect 1368 -51 1538 -50
rect 1368 -85 1369 -51
rect 1369 -85 1537 -51
rect 1537 -85 1538 -51
rect 1368 -159 1538 -85
rect 1368 -193 1369 -159
rect 1369 -193 1537 -159
rect 1537 -193 1538 -159
rect 1368 -194 1538 -193
rect 1740 -51 1910 -50
rect 1740 -85 1741 -51
rect 1741 -85 1909 -51
rect 1909 -85 1910 -51
rect 1740 -159 1910 -85
rect 1740 -193 1741 -159
rect 1741 -193 1909 -159
rect 1909 -193 1910 -159
rect 1740 -194 1910 -193
rect 2112 -51 2282 -50
rect 2112 -85 2113 -51
rect 2113 -85 2281 -51
rect 2281 -85 2282 -51
rect 2112 -159 2282 -85
rect 2112 -193 2113 -159
rect 2113 -193 2281 -159
rect 2281 -193 2282 -159
rect 2112 -194 2282 -193
rect 2484 -51 2654 -50
rect 2484 -85 2485 -51
rect 2485 -85 2653 -51
rect 2653 -85 2654 -51
rect 2484 -159 2654 -85
rect 2484 -193 2485 -159
rect 2485 -193 2653 -159
rect 2653 -193 2654 -159
rect 2484 -194 2654 -193
rect 2856 -51 3026 -50
rect 2856 -85 2857 -51
rect 2857 -85 3025 -51
rect 3025 -85 3026 -51
rect 2856 -159 3026 -85
rect 2856 -193 2857 -159
rect 2857 -193 3025 -159
rect 3025 -193 3026 -159
rect 2856 -194 3026 -193
rect 3228 -51 3398 -50
rect 3228 -85 3229 -51
rect 3229 -85 3397 -51
rect 3397 -85 3398 -51
rect 3228 -159 3398 -85
rect 3228 -193 3229 -159
rect 3229 -193 3397 -159
rect 3397 -193 3398 -159
rect 3228 -194 3398 -193
rect 3600 -51 3770 -50
rect 3600 -85 3601 -51
rect 3601 -85 3769 -51
rect 3769 -85 3770 -51
rect 3600 -159 3770 -85
rect 3600 -193 3601 -159
rect 3601 -193 3769 -159
rect 3769 -193 3770 -159
rect 3600 -194 3770 -193
rect 3972 -51 4142 -50
rect 3972 -85 3973 -51
rect 3973 -85 4141 -51
rect 4141 -85 4142 -51
rect 3972 -159 4142 -85
rect 3972 -193 3973 -159
rect 3973 -193 4141 -159
rect 4141 -193 4142 -159
rect 3972 -194 4142 -193
rect 4344 -51 4514 -50
rect 4344 -85 4345 -51
rect 4345 -85 4513 -51
rect 4513 -85 4514 -51
rect 4344 -159 4514 -85
rect 4344 -193 4345 -159
rect 4345 -193 4513 -159
rect 4513 -193 4514 -159
rect 4344 -194 4514 -193
rect 4716 -51 4886 -50
rect 4716 -85 4717 -51
rect 4717 -85 4885 -51
rect 4885 -85 4886 -51
rect 4716 -159 4886 -85
rect 4716 -193 4717 -159
rect 4717 -193 4885 -159
rect 4885 -193 4886 -159
rect 4716 -194 4886 -193
rect 5088 -51 5258 -50
rect 5088 -85 5089 -51
rect 5089 -85 5257 -51
rect 5257 -85 5258 -51
rect 5088 -159 5258 -85
rect 5088 -193 5089 -159
rect 5089 -193 5257 -159
rect 5257 -193 5258 -159
rect 5088 -194 5258 -193
rect -492 -687 -322 -674
rect -492 -721 -491 -687
rect -491 -721 -323 -687
rect -323 -721 -322 -687
rect -492 -734 -322 -721
rect -120 -687 50 -674
rect -120 -721 -119 -687
rect -119 -721 49 -687
rect 49 -721 50 -687
rect -120 -734 50 -721
rect 252 -687 422 -674
rect 252 -721 253 -687
rect 253 -721 421 -687
rect 421 -721 422 -687
rect 252 -734 422 -721
rect 624 -687 794 -674
rect 624 -721 625 -687
rect 625 -721 793 -687
rect 793 -721 794 -687
rect 624 -734 794 -721
rect 996 -687 1166 -674
rect 996 -721 997 -687
rect 997 -721 1165 -687
rect 1165 -721 1166 -687
rect 996 -734 1166 -721
rect 1368 -687 1538 -674
rect 1368 -721 1369 -687
rect 1369 -721 1537 -687
rect 1537 -721 1538 -687
rect 1368 -734 1538 -721
rect 1740 -687 1910 -674
rect 1740 -721 1741 -687
rect 1741 -721 1909 -687
rect 1909 -721 1910 -687
rect 1740 -734 1910 -721
rect 2112 -687 2282 -674
rect 2112 -721 2113 -687
rect 2113 -721 2281 -687
rect 2281 -721 2282 -687
rect 2112 -734 2282 -721
rect 2484 -687 2654 -674
rect 2484 -721 2485 -687
rect 2485 -721 2653 -687
rect 2653 -721 2654 -687
rect 2484 -734 2654 -721
rect 2856 -687 3026 -674
rect 2856 -721 2857 -687
rect 2857 -721 3025 -687
rect 3025 -721 3026 -687
rect 2856 -734 3026 -721
rect 3228 -687 3398 -674
rect 3228 -721 3229 -687
rect 3229 -721 3397 -687
rect 3397 -721 3398 -687
rect 3228 -734 3398 -721
rect 3600 -687 3770 -674
rect 3600 -721 3601 -687
rect 3601 -721 3769 -687
rect 3769 -721 3770 -687
rect 3600 -734 3770 -721
rect 3972 -687 4142 -674
rect 3972 -721 3973 -687
rect 3973 -721 4141 -687
rect 4141 -721 4142 -687
rect 3972 -734 4142 -721
rect 4344 -687 4514 -674
rect 4344 -721 4345 -687
rect 4345 -721 4513 -687
rect 4513 -721 4514 -687
rect 4344 -734 4514 -721
rect 5460 1113 5630 1126
rect 5460 1079 5461 1113
rect 5461 1079 5629 1113
rect 5629 1079 5630 1113
rect 5460 1066 5630 1079
rect 5832 1113 6002 1126
rect 5832 1079 5833 1113
rect 5833 1079 6001 1113
rect 6001 1079 6002 1113
rect 5832 1066 6002 1079
rect 6204 1113 6374 1126
rect 6204 1079 6205 1113
rect 6205 1079 6373 1113
rect 6373 1079 6374 1113
rect 6204 1066 6374 1079
rect 6576 1113 6746 1126
rect 6576 1079 6577 1113
rect 6577 1079 6745 1113
rect 6745 1079 6746 1113
rect 6576 1066 6746 1079
rect 6948 1113 7118 1126
rect 6948 1079 6949 1113
rect 6949 1079 7117 1113
rect 7117 1079 7118 1113
rect 6948 1066 7118 1079
rect 7320 1113 7490 1126
rect 7320 1079 7321 1113
rect 7321 1079 7489 1113
rect 7489 1079 7490 1113
rect 7320 1066 7490 1079
rect 7692 1113 7862 1126
rect 7692 1079 7693 1113
rect 7693 1079 7861 1113
rect 7861 1079 7862 1113
rect 7692 1066 7862 1079
rect 8064 1113 8234 1126
rect 8064 1079 8065 1113
rect 8065 1079 8233 1113
rect 8233 1079 8234 1113
rect 8064 1066 8234 1079
rect 8436 1113 8606 1126
rect 8436 1079 8437 1113
rect 8437 1079 8605 1113
rect 8605 1079 8606 1113
rect 8436 1066 8606 1079
rect 8808 1113 8978 1126
rect 8808 1079 8809 1113
rect 8809 1079 8977 1113
rect 8977 1079 8978 1113
rect 8808 1066 8978 1079
rect 9180 1113 9350 1126
rect 9180 1079 9181 1113
rect 9181 1079 9349 1113
rect 9349 1079 9350 1113
rect 9180 1066 9350 1079
rect 9552 1113 9722 1126
rect 9552 1079 9553 1113
rect 9553 1079 9721 1113
rect 9721 1079 9722 1113
rect 9552 1066 9722 1079
rect 9924 1113 10094 1126
rect 9924 1079 9925 1113
rect 9925 1079 10093 1113
rect 10093 1079 10094 1113
rect 9924 1066 10094 1079
rect 10296 1113 10466 1126
rect 10296 1079 10297 1113
rect 10297 1079 10465 1113
rect 10465 1079 10466 1113
rect 10296 1066 10466 1079
rect 10668 1113 10838 1126
rect 10668 1079 10669 1113
rect 10669 1079 10837 1113
rect 10837 1079 10838 1113
rect 10668 1066 10838 1079
rect 11040 1113 11210 1126
rect 11040 1079 11041 1113
rect 11041 1079 11209 1113
rect 11209 1079 11210 1113
rect 11040 1066 11210 1079
rect 5460 585 5630 586
rect 5460 551 5461 585
rect 5461 551 5629 585
rect 5629 551 5630 585
rect 5460 477 5630 551
rect 5460 443 5461 477
rect 5461 443 5629 477
rect 5629 443 5630 477
rect 5460 442 5630 443
rect 5832 585 6002 586
rect 5832 551 5833 585
rect 5833 551 6001 585
rect 6001 551 6002 585
rect 5832 477 6002 551
rect 5832 443 5833 477
rect 5833 443 6001 477
rect 6001 443 6002 477
rect 5832 442 6002 443
rect 6204 585 6374 586
rect 6204 551 6205 585
rect 6205 551 6373 585
rect 6373 551 6374 585
rect 6204 477 6374 551
rect 6204 443 6205 477
rect 6205 443 6373 477
rect 6373 443 6374 477
rect 6204 442 6374 443
rect 6576 585 6746 586
rect 6576 551 6577 585
rect 6577 551 6745 585
rect 6745 551 6746 585
rect 6576 477 6746 551
rect 6576 443 6577 477
rect 6577 443 6745 477
rect 6745 443 6746 477
rect 6576 442 6746 443
rect 6948 585 7118 586
rect 6948 551 6949 585
rect 6949 551 7117 585
rect 7117 551 7118 585
rect 6948 477 7118 551
rect 6948 443 6949 477
rect 6949 443 7117 477
rect 7117 443 7118 477
rect 6948 442 7118 443
rect 7320 585 7490 586
rect 7320 551 7321 585
rect 7321 551 7489 585
rect 7489 551 7490 585
rect 7320 477 7490 551
rect 7320 443 7321 477
rect 7321 443 7489 477
rect 7489 443 7490 477
rect 7320 442 7490 443
rect 7692 585 7862 586
rect 7692 551 7693 585
rect 7693 551 7861 585
rect 7861 551 7862 585
rect 7692 477 7862 551
rect 7692 443 7693 477
rect 7693 443 7861 477
rect 7861 443 7862 477
rect 7692 442 7862 443
rect 8064 585 8234 586
rect 8064 551 8065 585
rect 8065 551 8233 585
rect 8233 551 8234 585
rect 8064 477 8234 551
rect 8064 443 8065 477
rect 8065 443 8233 477
rect 8233 443 8234 477
rect 8064 442 8234 443
rect 8436 585 8606 586
rect 8436 551 8437 585
rect 8437 551 8605 585
rect 8605 551 8606 585
rect 8436 477 8606 551
rect 8436 443 8437 477
rect 8437 443 8605 477
rect 8605 443 8606 477
rect 8436 442 8606 443
rect 8808 585 8978 586
rect 8808 551 8809 585
rect 8809 551 8977 585
rect 8977 551 8978 585
rect 8808 477 8978 551
rect 8808 443 8809 477
rect 8809 443 8977 477
rect 8977 443 8978 477
rect 8808 442 8978 443
rect 9180 585 9350 586
rect 9180 551 9181 585
rect 9181 551 9349 585
rect 9349 551 9350 585
rect 9180 477 9350 551
rect 9180 443 9181 477
rect 9181 443 9349 477
rect 9349 443 9350 477
rect 9180 442 9350 443
rect 9552 585 9722 586
rect 9552 551 9553 585
rect 9553 551 9721 585
rect 9721 551 9722 585
rect 9552 477 9722 551
rect 9552 443 9553 477
rect 9553 443 9721 477
rect 9721 443 9722 477
rect 9552 442 9722 443
rect 9924 585 10094 586
rect 9924 551 9925 585
rect 9925 551 10093 585
rect 10093 551 10094 585
rect 9924 477 10094 551
rect 9924 443 9925 477
rect 9925 443 10093 477
rect 10093 443 10094 477
rect 9924 442 10094 443
rect 10296 585 10466 586
rect 10296 551 10297 585
rect 10297 551 10465 585
rect 10465 551 10466 585
rect 10296 477 10466 551
rect 10296 443 10297 477
rect 10297 443 10465 477
rect 10465 443 10466 477
rect 10296 442 10466 443
rect 10668 585 10838 586
rect 10668 551 10669 585
rect 10669 551 10837 585
rect 10837 551 10838 585
rect 10668 477 10838 551
rect 10668 443 10669 477
rect 10669 443 10837 477
rect 10837 443 10838 477
rect 10668 442 10838 443
rect 11040 585 11210 586
rect 11040 551 11041 585
rect 11041 551 11209 585
rect 11209 551 11210 585
rect 11040 477 11210 551
rect 11040 443 11041 477
rect 11041 443 11209 477
rect 11209 443 11210 477
rect 11040 442 11210 443
rect 5460 -51 5630 -50
rect 5460 -85 5461 -51
rect 5461 -85 5629 -51
rect 5629 -85 5630 -51
rect 5460 -159 5630 -85
rect 5460 -193 5461 -159
rect 5461 -193 5629 -159
rect 5629 -193 5630 -159
rect 5460 -194 5630 -193
rect 5832 -51 6002 -50
rect 5832 -85 5833 -51
rect 5833 -85 6001 -51
rect 6001 -85 6002 -51
rect 5832 -159 6002 -85
rect 5832 -193 5833 -159
rect 5833 -193 6001 -159
rect 6001 -193 6002 -159
rect 5832 -194 6002 -193
rect 6204 -51 6374 -50
rect 6204 -85 6205 -51
rect 6205 -85 6373 -51
rect 6373 -85 6374 -51
rect 6204 -159 6374 -85
rect 6204 -193 6205 -159
rect 6205 -193 6373 -159
rect 6373 -193 6374 -159
rect 6204 -194 6374 -193
rect 6576 -51 6746 -50
rect 6576 -85 6577 -51
rect 6577 -85 6745 -51
rect 6745 -85 6746 -51
rect 6576 -159 6746 -85
rect 6576 -193 6577 -159
rect 6577 -193 6745 -159
rect 6745 -193 6746 -159
rect 6576 -194 6746 -193
rect 6948 -51 7118 -50
rect 6948 -85 6949 -51
rect 6949 -85 7117 -51
rect 7117 -85 7118 -51
rect 6948 -159 7118 -85
rect 6948 -193 6949 -159
rect 6949 -193 7117 -159
rect 7117 -193 7118 -159
rect 6948 -194 7118 -193
rect 7320 -51 7490 -50
rect 7320 -85 7321 -51
rect 7321 -85 7489 -51
rect 7489 -85 7490 -51
rect 7320 -159 7490 -85
rect 7320 -193 7321 -159
rect 7321 -193 7489 -159
rect 7489 -193 7490 -159
rect 7320 -194 7490 -193
rect 7692 -51 7862 -50
rect 7692 -85 7693 -51
rect 7693 -85 7861 -51
rect 7861 -85 7862 -51
rect 7692 -159 7862 -85
rect 7692 -193 7693 -159
rect 7693 -193 7861 -159
rect 7861 -193 7862 -159
rect 7692 -194 7862 -193
rect 8064 -51 8234 -50
rect 8064 -85 8065 -51
rect 8065 -85 8233 -51
rect 8233 -85 8234 -51
rect 8064 -159 8234 -85
rect 8064 -193 8065 -159
rect 8065 -193 8233 -159
rect 8233 -193 8234 -159
rect 8064 -194 8234 -193
rect 8436 -51 8606 -50
rect 8436 -85 8437 -51
rect 8437 -85 8605 -51
rect 8605 -85 8606 -51
rect 8436 -159 8606 -85
rect 8436 -193 8437 -159
rect 8437 -193 8605 -159
rect 8605 -193 8606 -159
rect 8436 -194 8606 -193
rect 8808 -51 8978 -50
rect 8808 -85 8809 -51
rect 8809 -85 8977 -51
rect 8977 -85 8978 -51
rect 8808 -159 8978 -85
rect 8808 -193 8809 -159
rect 8809 -193 8977 -159
rect 8977 -193 8978 -159
rect 8808 -194 8978 -193
rect 9180 -51 9350 -50
rect 9180 -85 9181 -51
rect 9181 -85 9349 -51
rect 9349 -85 9350 -51
rect 9180 -159 9350 -85
rect 9180 -193 9181 -159
rect 9181 -193 9349 -159
rect 9349 -193 9350 -159
rect 9180 -194 9350 -193
rect 9552 -51 9722 -50
rect 9552 -85 9553 -51
rect 9553 -85 9721 -51
rect 9721 -85 9722 -51
rect 9552 -159 9722 -85
rect 9552 -193 9553 -159
rect 9553 -193 9721 -159
rect 9721 -193 9722 -159
rect 9552 -194 9722 -193
rect 9924 -51 10094 -50
rect 9924 -85 9925 -51
rect 9925 -85 10093 -51
rect 10093 -85 10094 -51
rect 9924 -159 10094 -85
rect 9924 -193 9925 -159
rect 9925 -193 10093 -159
rect 10093 -193 10094 -159
rect 9924 -194 10094 -193
rect 10296 -51 10466 -50
rect 10296 -85 10297 -51
rect 10297 -85 10465 -51
rect 10465 -85 10466 -51
rect 10296 -159 10466 -85
rect 10296 -193 10297 -159
rect 10297 -193 10465 -159
rect 10465 -193 10466 -159
rect 10296 -194 10466 -193
rect 10668 -51 10838 -50
rect 10668 -85 10669 -51
rect 10669 -85 10837 -51
rect 10837 -85 10838 -51
rect 10668 -159 10838 -85
rect 10668 -193 10669 -159
rect 10669 -193 10837 -159
rect 10837 -193 10838 -159
rect 10668 -194 10838 -193
rect 11040 -51 11210 -50
rect 11040 -85 11041 -51
rect 11041 -85 11209 -51
rect 11209 -85 11210 -51
rect 11040 -159 11210 -85
rect 11040 -193 11041 -159
rect 11041 -193 11209 -159
rect 11209 -193 11210 -159
rect 11040 -194 11210 -193
rect 4716 -687 4886 -674
rect 4716 -721 4717 -687
rect 4717 -721 4885 -687
rect 4885 -721 4886 -687
rect 4716 -734 4886 -721
rect 5088 -687 5258 -674
rect 5088 -721 5089 -687
rect 5089 -721 5257 -687
rect 5257 -721 5258 -687
rect 5088 -734 5258 -721
rect 5460 -687 5630 -674
rect 5460 -721 5461 -687
rect 5461 -721 5629 -687
rect 5629 -721 5630 -687
rect 5460 -734 5630 -721
rect 5832 -687 6002 -674
rect 5832 -721 5833 -687
rect 5833 -721 6001 -687
rect 6001 -721 6002 -687
rect 5832 -734 6002 -721
rect 6204 -687 6374 -674
rect 6204 -721 6205 -687
rect 6205 -721 6373 -687
rect 6373 -721 6374 -687
rect 6204 -734 6374 -721
rect 6576 -687 6746 -674
rect 6576 -721 6577 -687
rect 6577 -721 6745 -687
rect 6745 -721 6746 -687
rect 6576 -734 6746 -721
rect 6948 -687 7118 -674
rect 6948 -721 6949 -687
rect 6949 -721 7117 -687
rect 7117 -721 7118 -687
rect 6948 -734 7118 -721
rect 7320 -687 7490 -674
rect 7320 -721 7321 -687
rect 7321 -721 7489 -687
rect 7489 -721 7490 -687
rect 7320 -734 7490 -721
rect 7692 -687 7862 -674
rect 7692 -721 7693 -687
rect 7693 -721 7861 -687
rect 7861 -721 7862 -687
rect 7692 -734 7862 -721
rect 8064 -687 8234 -674
rect 8064 -721 8065 -687
rect 8065 -721 8233 -687
rect 8233 -721 8234 -687
rect 8064 -734 8234 -721
rect 8436 -687 8606 -674
rect 8436 -721 8437 -687
rect 8437 -721 8605 -687
rect 8605 -721 8606 -687
rect 8436 -734 8606 -721
rect 8808 -687 8978 -674
rect 8808 -721 8809 -687
rect 8809 -721 8977 -687
rect 8977 -721 8978 -687
rect 8808 -734 8978 -721
rect 9180 -687 9350 -674
rect 9180 -721 9181 -687
rect 9181 -721 9349 -687
rect 9349 -721 9350 -687
rect 9180 -734 9350 -721
rect 9552 -687 9722 -674
rect 9552 -721 9553 -687
rect 9553 -721 9721 -687
rect 9721 -721 9722 -687
rect 9552 -734 9722 -721
rect 9924 -687 10094 -674
rect 9924 -721 9925 -687
rect 9925 -721 10093 -687
rect 10093 -721 10094 -687
rect 9924 -734 10094 -721
rect 10296 -687 10466 -674
rect 10296 -721 10297 -687
rect 10297 -721 10465 -687
rect 10465 -721 10466 -687
rect 10296 -734 10466 -721
rect 10668 -687 10838 -674
rect 10668 -721 10669 -687
rect 10669 -721 10837 -687
rect 10837 -721 10838 -687
rect 10668 -734 10838 -721
rect 11040 -687 11210 -674
rect 11040 -721 11041 -687
rect 11041 -721 11209 -687
rect 11209 -721 11210 -687
rect 11040 -734 11210 -721
rect 996 -1275 1166 -1260
rect 996 -1309 997 -1275
rect 997 -1309 1165 -1275
rect 1165 -1309 1166 -1275
rect 996 -1324 1166 -1309
rect 1368 -1275 1538 -1260
rect 1368 -1309 1369 -1275
rect 1369 -1309 1537 -1275
rect 1537 -1309 1538 -1275
rect 1368 -1324 1538 -1309
rect 1740 -1275 1910 -1260
rect 1740 -1309 1741 -1275
rect 1741 -1309 1909 -1275
rect 1909 -1309 1910 -1275
rect 1740 -1324 1910 -1309
rect 2112 -1275 2282 -1260
rect 2112 -1309 2113 -1275
rect 2113 -1309 2281 -1275
rect 2281 -1309 2282 -1275
rect 2112 -1324 2282 -1309
rect 2484 -1275 2654 -1260
rect 2484 -1309 2485 -1275
rect 2485 -1309 2653 -1275
rect 2653 -1309 2654 -1275
rect 2484 -1324 2654 -1309
rect 2856 -1275 3026 -1260
rect 2856 -1309 2857 -1275
rect 2857 -1309 3025 -1275
rect 3025 -1309 3026 -1275
rect 2856 -1324 3026 -1309
rect 3228 -1275 3398 -1260
rect 3228 -1309 3229 -1275
rect 3229 -1309 3397 -1275
rect 3397 -1309 3398 -1275
rect 3228 -1324 3398 -1309
rect 3600 -1275 3770 -1260
rect 3600 -1309 3601 -1275
rect 3601 -1309 3769 -1275
rect 3769 -1309 3770 -1275
rect 3600 -1324 3770 -1309
rect 5592 -1314 5874 -1042
rect 6336 -1314 6618 -1042
rect 7080 -1314 7362 -1042
rect 7824 -1314 8106 -1042
rect 8568 -1314 8850 -1042
rect 9312 -1314 9594 -1042
rect 10056 -1314 10338 -1042
rect 10800 -1314 11082 -1042
rect 996 -2203 1166 -2202
rect 996 -2237 997 -2203
rect 997 -2237 1165 -2203
rect 1165 -2237 1166 -2203
rect 996 -2311 1166 -2237
rect 996 -2345 997 -2311
rect 997 -2345 1165 -2311
rect 1165 -2345 1166 -2311
rect 996 -2346 1166 -2345
rect 1368 -2203 1538 -2202
rect 1368 -2237 1369 -2203
rect 1369 -2237 1537 -2203
rect 1537 -2237 1538 -2203
rect 1368 -2311 1538 -2237
rect 1368 -2345 1369 -2311
rect 1369 -2345 1537 -2311
rect 1537 -2345 1538 -2311
rect 1368 -2346 1538 -2345
rect 1740 -2203 1910 -2202
rect 1740 -2237 1741 -2203
rect 1741 -2237 1909 -2203
rect 1909 -2237 1910 -2203
rect 1740 -2311 1910 -2237
rect 1740 -2345 1741 -2311
rect 1741 -2345 1909 -2311
rect 1909 -2345 1910 -2311
rect 1740 -2346 1910 -2345
rect 2112 -2203 2282 -2202
rect 2112 -2237 2113 -2203
rect 2113 -2237 2281 -2203
rect 2281 -2237 2282 -2203
rect 2112 -2311 2282 -2237
rect 2112 -2345 2113 -2311
rect 2113 -2345 2281 -2311
rect 2281 -2345 2282 -2311
rect 2112 -2346 2282 -2345
rect 2484 -2203 2654 -2202
rect 2484 -2237 2485 -2203
rect 2485 -2237 2653 -2203
rect 2653 -2237 2654 -2203
rect 2484 -2311 2654 -2237
rect 2484 -2345 2485 -2311
rect 2485 -2345 2653 -2311
rect 2653 -2345 2654 -2311
rect 2484 -2346 2654 -2345
rect 2856 -2203 3026 -2202
rect 2856 -2237 2857 -2203
rect 2857 -2237 3025 -2203
rect 3025 -2237 3026 -2203
rect 2856 -2311 3026 -2237
rect 2856 -2345 2857 -2311
rect 2857 -2345 3025 -2311
rect 3025 -2345 3026 -2311
rect 2856 -2346 3026 -2345
rect 3228 -2203 3398 -2202
rect 3228 -2237 3229 -2203
rect 3229 -2237 3397 -2203
rect 3397 -2237 3398 -2203
rect 3228 -2311 3398 -2237
rect 3228 -2345 3229 -2311
rect 3229 -2345 3397 -2311
rect 3397 -2345 3398 -2311
rect 3228 -2346 3398 -2345
rect 3600 -2203 3770 -2202
rect 3600 -2237 3601 -2203
rect 3601 -2237 3769 -2203
rect 3769 -2237 3770 -2203
rect 3600 -2311 3770 -2237
rect 3600 -2345 3601 -2311
rect 3601 -2345 3769 -2311
rect 3769 -2345 3770 -2311
rect 3600 -2346 3770 -2345
rect 6012 -3088 6294 -2816
rect 996 -3239 1166 -3238
rect 996 -3273 997 -3239
rect 997 -3273 1165 -3239
rect 1165 -3273 1166 -3239
rect 996 -3347 1166 -3273
rect 996 -3381 997 -3347
rect 997 -3381 1165 -3347
rect 1165 -3381 1166 -3347
rect 996 -3382 1166 -3381
rect 1368 -3239 1538 -3238
rect 1368 -3273 1369 -3239
rect 1369 -3273 1537 -3239
rect 1537 -3273 1538 -3239
rect 1368 -3347 1538 -3273
rect 1368 -3381 1369 -3347
rect 1369 -3381 1537 -3347
rect 1537 -3381 1538 -3347
rect 1368 -3382 1538 -3381
rect 1740 -3239 1910 -3238
rect 1740 -3273 1741 -3239
rect 1741 -3273 1909 -3239
rect 1909 -3273 1910 -3239
rect 1740 -3347 1910 -3273
rect 1740 -3381 1741 -3347
rect 1741 -3381 1909 -3347
rect 1909 -3381 1910 -3347
rect 1740 -3382 1910 -3381
rect 2112 -3239 2282 -3238
rect 2112 -3273 2113 -3239
rect 2113 -3273 2281 -3239
rect 2281 -3273 2282 -3239
rect 2112 -3347 2282 -3273
rect 2112 -3381 2113 -3347
rect 2113 -3381 2281 -3347
rect 2281 -3381 2282 -3347
rect 2112 -3382 2282 -3381
rect 2484 -3239 2654 -3238
rect 2484 -3273 2485 -3239
rect 2485 -3273 2653 -3239
rect 2653 -3273 2654 -3239
rect 2484 -3347 2654 -3273
rect 2484 -3381 2485 -3347
rect 2485 -3381 2653 -3347
rect 2653 -3381 2654 -3347
rect 2484 -3382 2654 -3381
rect 2856 -3239 3026 -3238
rect 2856 -3273 2857 -3239
rect 2857 -3273 3025 -3239
rect 3025 -3273 3026 -3239
rect 2856 -3347 3026 -3273
rect 2856 -3381 2857 -3347
rect 2857 -3381 3025 -3347
rect 3025 -3381 3026 -3347
rect 2856 -3382 3026 -3381
rect 3228 -3239 3398 -3238
rect 3228 -3273 3229 -3239
rect 3229 -3273 3397 -3239
rect 3397 -3273 3398 -3239
rect 3228 -3347 3398 -3273
rect 3228 -3381 3229 -3347
rect 3229 -3381 3397 -3347
rect 3397 -3381 3398 -3347
rect 3228 -3382 3398 -3381
rect 3600 -3239 3770 -3238
rect 3600 -3273 3601 -3239
rect 3601 -3273 3769 -3239
rect 3769 -3273 3770 -3239
rect 3600 -3347 3770 -3273
rect 3600 -3381 3601 -3347
rect 3601 -3381 3769 -3347
rect 3769 -3381 3770 -3347
rect 3600 -3382 3770 -3381
rect 5686 -3690 5846 -3528
rect 5686 -4090 5846 -3928
rect 996 -4275 1166 -4274
rect 996 -4309 997 -4275
rect 997 -4309 1165 -4275
rect 1165 -4309 1166 -4275
rect 996 -4383 1166 -4309
rect 996 -4417 997 -4383
rect 997 -4417 1165 -4383
rect 1165 -4417 1166 -4383
rect 996 -4418 1166 -4417
rect 1368 -4275 1538 -4274
rect 1368 -4309 1369 -4275
rect 1369 -4309 1537 -4275
rect 1537 -4309 1538 -4275
rect 1368 -4383 1538 -4309
rect 1368 -4417 1369 -4383
rect 1369 -4417 1537 -4383
rect 1537 -4417 1538 -4383
rect 1368 -4418 1538 -4417
rect 1740 -4275 1910 -4274
rect 1740 -4309 1741 -4275
rect 1741 -4309 1909 -4275
rect 1909 -4309 1910 -4275
rect 1740 -4383 1910 -4309
rect 1740 -4417 1741 -4383
rect 1741 -4417 1909 -4383
rect 1909 -4417 1910 -4383
rect 1740 -4418 1910 -4417
rect 2112 -4275 2282 -4274
rect 2112 -4309 2113 -4275
rect 2113 -4309 2281 -4275
rect 2281 -4309 2282 -4275
rect 2112 -4383 2282 -4309
rect 2112 -4417 2113 -4383
rect 2113 -4417 2281 -4383
rect 2281 -4417 2282 -4383
rect 2112 -4418 2282 -4417
rect 2484 -4275 2654 -4274
rect 2484 -4309 2485 -4275
rect 2485 -4309 2653 -4275
rect 2653 -4309 2654 -4275
rect 2484 -4383 2654 -4309
rect 2484 -4417 2485 -4383
rect 2485 -4417 2653 -4383
rect 2653 -4417 2654 -4383
rect 2484 -4418 2654 -4417
rect 2856 -4275 3026 -4274
rect 2856 -4309 2857 -4275
rect 2857 -4309 3025 -4275
rect 3025 -4309 3026 -4275
rect 2856 -4383 3026 -4309
rect 2856 -4417 2857 -4383
rect 2857 -4417 3025 -4383
rect 3025 -4417 3026 -4383
rect 2856 -4418 3026 -4417
rect 3228 -4275 3398 -4274
rect 3228 -4309 3229 -4275
rect 3229 -4309 3397 -4275
rect 3397 -4309 3398 -4275
rect 3228 -4383 3398 -4309
rect 3228 -4417 3229 -4383
rect 3229 -4417 3397 -4383
rect 3397 -4417 3398 -4383
rect 3228 -4418 3398 -4417
rect 3600 -4275 3770 -4274
rect 3600 -4309 3601 -4275
rect 3601 -4309 3769 -4275
rect 3769 -4309 3770 -4275
rect 3600 -4383 3770 -4309
rect 3600 -4417 3601 -4383
rect 3601 -4417 3769 -4383
rect 3769 -4417 3770 -4383
rect 3600 -4418 3770 -4417
rect 5686 -4490 5846 -4328
rect 996 -5311 1166 -5300
rect 996 -5345 997 -5311
rect 997 -5345 1165 -5311
rect 1165 -5345 1166 -5311
rect 996 -5354 1166 -5345
rect 1368 -5311 1538 -5300
rect 1368 -5345 1369 -5311
rect 1369 -5345 1537 -5311
rect 1537 -5345 1538 -5311
rect 1368 -5354 1538 -5345
rect 1740 -5311 1910 -5300
rect 1740 -5345 1741 -5311
rect 1741 -5345 1909 -5311
rect 1909 -5345 1910 -5311
rect 1740 -5354 1910 -5345
rect 2112 -5311 2282 -5300
rect 2112 -5345 2113 -5311
rect 2113 -5345 2281 -5311
rect 2281 -5345 2282 -5311
rect 2112 -5354 2282 -5345
rect 2484 -5311 2654 -5300
rect 2484 -5345 2485 -5311
rect 2485 -5345 2653 -5311
rect 2653 -5345 2654 -5311
rect 2484 -5354 2654 -5345
rect 2856 -5311 3026 -5300
rect 2856 -5345 2857 -5311
rect 2857 -5345 3025 -5311
rect 3025 -5345 3026 -5311
rect 2856 -5354 3026 -5345
rect 3228 -5311 3398 -5300
rect 3228 -5345 3229 -5311
rect 3229 -5345 3397 -5311
rect 3397 -5345 3398 -5311
rect 3228 -5354 3398 -5345
rect 1976 -5820 2790 -5640
rect 996 -5969 1166 -5958
rect 996 -6003 997 -5969
rect 997 -6003 1165 -5969
rect 1165 -6003 1166 -5969
rect 996 -6014 1166 -6003
rect 1368 -5969 1538 -5958
rect 1368 -6003 1369 -5969
rect 1369 -6003 1537 -5969
rect 1537 -6003 1538 -5969
rect 1368 -6014 1538 -6003
rect 1740 -5969 1910 -5958
rect 1740 -6003 1741 -5969
rect 1741 -6003 1909 -5969
rect 1909 -6003 1910 -5969
rect 1740 -6014 1910 -6003
rect 2112 -5969 2282 -5958
rect 2112 -6003 2113 -5969
rect 2113 -6003 2281 -5969
rect 2281 -6003 2282 -5969
rect 2112 -6014 2282 -6003
rect 2484 -5969 2654 -5958
rect 2484 -6003 2485 -5969
rect 2485 -6003 2653 -5969
rect 2653 -6003 2654 -5969
rect 2484 -6014 2654 -6003
rect 3600 -5311 3770 -5300
rect 3600 -5345 3601 -5311
rect 3601 -5345 3769 -5311
rect 3769 -5345 3770 -5311
rect 3600 -5354 3770 -5345
rect 4102 -5496 4384 -5224
rect 4846 -5496 5128 -5224
rect 5590 -5496 5872 -5224
rect 2856 -5969 3026 -5958
rect 2856 -6003 2857 -5969
rect 2857 -6003 3025 -5969
rect 3025 -6003 3026 -5969
rect 2856 -6014 3026 -6003
rect 3228 -5969 3398 -5958
rect 3228 -6003 3229 -5969
rect 3229 -6003 3397 -5969
rect 3397 -6003 3398 -5969
rect 3228 -6014 3398 -6003
rect 3600 -5969 3770 -5958
rect 3600 -6003 3601 -5969
rect 3601 -6003 3769 -5969
rect 3769 -6003 3770 -5969
rect 3600 -6014 3770 -6003
rect 3972 -5969 4142 -5958
rect 3972 -6003 3973 -5969
rect 3973 -6003 4141 -5969
rect 4141 -6003 4142 -5969
rect 3972 -6014 4142 -6003
rect 4344 -5969 4514 -5958
rect 4344 -6003 4345 -5969
rect 4345 -6003 4513 -5969
rect 4513 -6003 4514 -5969
rect 4344 -6014 4514 -6003
rect 4716 -5969 4886 -5958
rect 4716 -6003 4717 -5969
rect 4717 -6003 4885 -5969
rect 4885 -6003 4886 -5969
rect 4716 -6014 4886 -6003
rect 5088 -5969 5258 -5958
rect 5088 -6003 5089 -5969
rect 5089 -6003 5257 -5969
rect 5257 -6003 5258 -5969
rect 5088 -6014 5258 -6003
rect 5460 -5969 5630 -5958
rect 5460 -6003 5461 -5969
rect 5461 -6003 5629 -5969
rect 5629 -6003 5630 -5969
rect 5460 -6014 5630 -6003
rect 6334 -5496 6616 -5224
rect 7078 -5496 7360 -5224
rect 7822 -5496 8104 -5224
rect 8566 -5496 8848 -5224
rect 9310 -5496 9592 -5224
rect 5986 -5786 6264 -5512
rect 5832 -5969 6002 -5958
rect 5832 -6003 5833 -5969
rect 5833 -6003 6001 -5969
rect 6001 -6003 6002 -5969
rect 5832 -6014 6002 -6003
rect 6204 -5969 6374 -5958
rect 6204 -6003 6205 -5969
rect 6205 -6003 6373 -5969
rect 6373 -6003 6374 -5969
rect 6204 -6014 6374 -6003
rect 6576 -5969 6746 -5958
rect 6576 -6003 6577 -5969
rect 6577 -6003 6745 -5969
rect 6745 -6003 6746 -5969
rect 6576 -6014 6746 -6003
rect 6948 -5969 7118 -5958
rect 6948 -6003 6949 -5969
rect 6949 -6003 7117 -5969
rect 7117 -6003 7118 -5969
rect 6948 -6014 7118 -6003
rect 7320 -5969 7490 -5958
rect 7320 -6003 7321 -5969
rect 7321 -6003 7489 -5969
rect 7489 -6003 7490 -5969
rect 7320 -6014 7490 -6003
rect 7692 -5969 7862 -5958
rect 7692 -6003 7693 -5969
rect 7693 -6003 7861 -5969
rect 7861 -6003 7862 -5969
rect 7692 -6014 7862 -6003
rect 8064 -5969 8234 -5958
rect 8064 -6003 8065 -5969
rect 8065 -6003 8233 -5969
rect 8233 -6003 8234 -5969
rect 8064 -6014 8234 -6003
rect 8436 -5969 8606 -5958
rect 8436 -6003 8437 -5969
rect 8437 -6003 8605 -5969
rect 8605 -6003 8606 -5969
rect 8436 -6014 8606 -6003
rect 8808 -5969 8978 -5958
rect 8808 -6003 8809 -5969
rect 8809 -6003 8977 -5969
rect 8977 -6003 8978 -5969
rect 8808 -6014 8978 -6003
rect 9180 -5969 9350 -5958
rect 9180 -6003 9181 -5969
rect 9181 -6003 9349 -5969
rect 9349 -6003 9350 -5969
rect 9180 -6014 9350 -6003
rect 9552 -5969 9722 -5958
rect 9552 -6003 9553 -5969
rect 9553 -6003 9721 -5969
rect 9721 -6003 9722 -5969
rect 9552 -6014 9722 -6003
rect 996 -6279 1166 -6278
rect 996 -6313 997 -6279
rect 997 -6313 1165 -6279
rect 1165 -6313 1166 -6279
rect 996 -6387 1166 -6313
rect 996 -6421 997 -6387
rect 997 -6421 1165 -6387
rect 1165 -6421 1166 -6387
rect 996 -6422 1166 -6421
rect 1368 -6279 1538 -6278
rect 1368 -6313 1369 -6279
rect 1369 -6313 1537 -6279
rect 1537 -6313 1538 -6279
rect 1368 -6387 1538 -6313
rect 1368 -6421 1369 -6387
rect 1369 -6421 1537 -6387
rect 1537 -6421 1538 -6387
rect 1368 -6422 1538 -6421
rect 1740 -6279 1910 -6278
rect 1740 -6313 1741 -6279
rect 1741 -6313 1909 -6279
rect 1909 -6313 1910 -6279
rect 1740 -6387 1910 -6313
rect 1740 -6421 1741 -6387
rect 1741 -6421 1909 -6387
rect 1909 -6421 1910 -6387
rect 1740 -6422 1910 -6421
rect 2112 -6279 2282 -6278
rect 2112 -6313 2113 -6279
rect 2113 -6313 2281 -6279
rect 2281 -6313 2282 -6279
rect 2112 -6387 2282 -6313
rect 2112 -6421 2113 -6387
rect 2113 -6421 2281 -6387
rect 2281 -6421 2282 -6387
rect 2112 -6422 2282 -6421
rect 2484 -6279 2654 -6278
rect 2484 -6313 2485 -6279
rect 2485 -6313 2653 -6279
rect 2653 -6313 2654 -6279
rect 2484 -6387 2654 -6313
rect 2484 -6421 2485 -6387
rect 2485 -6421 2653 -6387
rect 2653 -6421 2654 -6387
rect 2484 -6422 2654 -6421
rect 2856 -6279 3026 -6278
rect 2856 -6313 2857 -6279
rect 2857 -6313 3025 -6279
rect 3025 -6313 3026 -6279
rect 2856 -6387 3026 -6313
rect 2856 -6421 2857 -6387
rect 2857 -6421 3025 -6387
rect 3025 -6421 3026 -6387
rect 2856 -6422 3026 -6421
rect 3228 -6279 3398 -6278
rect 3228 -6313 3229 -6279
rect 3229 -6313 3397 -6279
rect 3397 -6313 3398 -6279
rect 3228 -6387 3398 -6313
rect 3228 -6421 3229 -6387
rect 3229 -6421 3397 -6387
rect 3397 -6421 3398 -6387
rect 3228 -6422 3398 -6421
rect 3600 -6279 3770 -6278
rect 3600 -6313 3601 -6279
rect 3601 -6313 3769 -6279
rect 3769 -6313 3770 -6279
rect 3600 -6387 3770 -6313
rect 3600 -6421 3601 -6387
rect 3601 -6421 3769 -6387
rect 3769 -6421 3770 -6387
rect 3600 -6422 3770 -6421
rect 3972 -6279 4142 -6278
rect 3972 -6313 3973 -6279
rect 3973 -6313 4141 -6279
rect 4141 -6313 4142 -6279
rect 3972 -6387 4142 -6313
rect 3972 -6421 3973 -6387
rect 3973 -6421 4141 -6387
rect 4141 -6421 4142 -6387
rect 3972 -6422 4142 -6421
rect 4344 -6279 4514 -6278
rect 4344 -6313 4345 -6279
rect 4345 -6313 4513 -6279
rect 4513 -6313 4514 -6279
rect 4344 -6387 4514 -6313
rect 4344 -6421 4345 -6387
rect 4345 -6421 4513 -6387
rect 4513 -6421 4514 -6387
rect 4344 -6422 4514 -6421
rect 4716 -6279 4886 -6278
rect 4716 -6313 4717 -6279
rect 4717 -6313 4885 -6279
rect 4885 -6313 4886 -6279
rect 4716 -6387 4886 -6313
rect 4716 -6421 4717 -6387
rect 4717 -6421 4885 -6387
rect 4885 -6421 4886 -6387
rect 4716 -6422 4886 -6421
rect 5088 -6279 5258 -6278
rect 5088 -6313 5089 -6279
rect 5089 -6313 5257 -6279
rect 5257 -6313 5258 -6279
rect 5088 -6387 5258 -6313
rect 5088 -6421 5089 -6387
rect 5089 -6421 5257 -6387
rect 5257 -6421 5258 -6387
rect 5088 -6422 5258 -6421
rect 5460 -6279 5630 -6278
rect 5460 -6313 5461 -6279
rect 5461 -6313 5629 -6279
rect 5629 -6313 5630 -6279
rect 5460 -6387 5630 -6313
rect 5460 -6421 5461 -6387
rect 5461 -6421 5629 -6387
rect 5629 -6421 5630 -6387
rect 5460 -6422 5630 -6421
rect 5832 -6279 6002 -6278
rect 5832 -6313 5833 -6279
rect 5833 -6313 6001 -6279
rect 6001 -6313 6002 -6279
rect 5832 -6387 6002 -6313
rect 5832 -6421 5833 -6387
rect 5833 -6421 6001 -6387
rect 6001 -6421 6002 -6387
rect 5832 -6422 6002 -6421
rect 6204 -6279 6374 -6278
rect 6204 -6313 6205 -6279
rect 6205 -6313 6373 -6279
rect 6373 -6313 6374 -6279
rect 6204 -6387 6374 -6313
rect 6204 -6421 6205 -6387
rect 6205 -6421 6373 -6387
rect 6373 -6421 6374 -6387
rect 6204 -6422 6374 -6421
rect 6576 -6279 6746 -6278
rect 6576 -6313 6577 -6279
rect 6577 -6313 6745 -6279
rect 6745 -6313 6746 -6279
rect 6576 -6387 6746 -6313
rect 6576 -6421 6577 -6387
rect 6577 -6421 6745 -6387
rect 6745 -6421 6746 -6387
rect 6576 -6422 6746 -6421
rect 6948 -6279 7118 -6278
rect 6948 -6313 6949 -6279
rect 6949 -6313 7117 -6279
rect 7117 -6313 7118 -6279
rect 6948 -6387 7118 -6313
rect 6948 -6421 6949 -6387
rect 6949 -6421 7117 -6387
rect 7117 -6421 7118 -6387
rect 6948 -6422 7118 -6421
rect 7320 -6279 7490 -6278
rect 7320 -6313 7321 -6279
rect 7321 -6313 7489 -6279
rect 7489 -6313 7490 -6279
rect 7320 -6387 7490 -6313
rect 7320 -6421 7321 -6387
rect 7321 -6421 7489 -6387
rect 7489 -6421 7490 -6387
rect 7320 -6422 7490 -6421
rect 7692 -6279 7862 -6278
rect 7692 -6313 7693 -6279
rect 7693 -6313 7861 -6279
rect 7861 -6313 7862 -6279
rect 7692 -6387 7862 -6313
rect 7692 -6421 7693 -6387
rect 7693 -6421 7861 -6387
rect 7861 -6421 7862 -6387
rect 7692 -6422 7862 -6421
rect 8064 -6279 8234 -6278
rect 8064 -6313 8065 -6279
rect 8065 -6313 8233 -6279
rect 8233 -6313 8234 -6279
rect 8064 -6387 8234 -6313
rect 8064 -6421 8065 -6387
rect 8065 -6421 8233 -6387
rect 8233 -6421 8234 -6387
rect 8064 -6422 8234 -6421
rect 8436 -6279 8606 -6278
rect 8436 -6313 8437 -6279
rect 8437 -6313 8605 -6279
rect 8605 -6313 8606 -6279
rect 8436 -6387 8606 -6313
rect 8436 -6421 8437 -6387
rect 8437 -6421 8605 -6387
rect 8605 -6421 8606 -6387
rect 8436 -6422 8606 -6421
rect 8808 -6279 8978 -6278
rect 8808 -6313 8809 -6279
rect 8809 -6313 8977 -6279
rect 8977 -6313 8978 -6279
rect 8808 -6387 8978 -6313
rect 8808 -6421 8809 -6387
rect 8809 -6421 8977 -6387
rect 8977 -6421 8978 -6387
rect 8808 -6422 8978 -6421
rect 9180 -6279 9350 -6278
rect 9180 -6313 9181 -6279
rect 9181 -6313 9349 -6279
rect 9349 -6313 9350 -6279
rect 9180 -6387 9350 -6313
rect 9180 -6421 9181 -6387
rect 9181 -6421 9349 -6387
rect 9349 -6421 9350 -6387
rect 9180 -6422 9350 -6421
rect 9552 -6279 9722 -6278
rect 9552 -6313 9553 -6279
rect 9553 -6313 9721 -6279
rect 9721 -6313 9722 -6279
rect 9552 -6387 9722 -6313
rect 9552 -6421 9553 -6387
rect 9553 -6421 9721 -6387
rect 9721 -6421 9722 -6387
rect 9552 -6422 9722 -6421
rect 996 -6697 1166 -6696
rect 996 -6731 997 -6697
rect 997 -6731 1165 -6697
rect 1165 -6731 1166 -6697
rect 996 -6805 1166 -6731
rect 996 -6839 997 -6805
rect 997 -6839 1165 -6805
rect 1165 -6839 1166 -6805
rect 996 -6840 1166 -6839
rect 1368 -6697 1538 -6696
rect 1368 -6731 1369 -6697
rect 1369 -6731 1537 -6697
rect 1537 -6731 1538 -6697
rect 1368 -6805 1538 -6731
rect 1368 -6839 1369 -6805
rect 1369 -6839 1537 -6805
rect 1537 -6839 1538 -6805
rect 1368 -6840 1538 -6839
rect 1740 -6697 1910 -6696
rect 1740 -6731 1741 -6697
rect 1741 -6731 1909 -6697
rect 1909 -6731 1910 -6697
rect 1740 -6805 1910 -6731
rect 1740 -6839 1741 -6805
rect 1741 -6839 1909 -6805
rect 1909 -6839 1910 -6805
rect 1740 -6840 1910 -6839
rect 2112 -6697 2282 -6696
rect 2112 -6731 2113 -6697
rect 2113 -6731 2281 -6697
rect 2281 -6731 2282 -6697
rect 2112 -6805 2282 -6731
rect 2112 -6839 2113 -6805
rect 2113 -6839 2281 -6805
rect 2281 -6839 2282 -6805
rect 2112 -6840 2282 -6839
rect 2484 -6697 2654 -6696
rect 2484 -6731 2485 -6697
rect 2485 -6731 2653 -6697
rect 2653 -6731 2654 -6697
rect 2484 -6805 2654 -6731
rect 2484 -6839 2485 -6805
rect 2485 -6839 2653 -6805
rect 2653 -6839 2654 -6805
rect 2484 -6840 2654 -6839
rect 2856 -6697 3026 -6696
rect 2856 -6731 2857 -6697
rect 2857 -6731 3025 -6697
rect 3025 -6731 3026 -6697
rect 2856 -6805 3026 -6731
rect 2856 -6839 2857 -6805
rect 2857 -6839 3025 -6805
rect 3025 -6839 3026 -6805
rect 2856 -6840 3026 -6839
rect 3228 -6697 3398 -6696
rect 3228 -6731 3229 -6697
rect 3229 -6731 3397 -6697
rect 3397 -6731 3398 -6697
rect 3228 -6805 3398 -6731
rect 3228 -6839 3229 -6805
rect 3229 -6839 3397 -6805
rect 3397 -6839 3398 -6805
rect 3228 -6840 3398 -6839
rect 3600 -6697 3770 -6696
rect 3600 -6731 3601 -6697
rect 3601 -6731 3769 -6697
rect 3769 -6731 3770 -6697
rect 3600 -6805 3770 -6731
rect 3600 -6839 3601 -6805
rect 3601 -6839 3769 -6805
rect 3769 -6839 3770 -6805
rect 3600 -6840 3770 -6839
rect 3972 -6697 4142 -6696
rect 3972 -6731 3973 -6697
rect 3973 -6731 4141 -6697
rect 4141 -6731 4142 -6697
rect 3972 -6805 4142 -6731
rect 3972 -6839 3973 -6805
rect 3973 -6839 4141 -6805
rect 4141 -6839 4142 -6805
rect 3972 -6840 4142 -6839
rect 4344 -6697 4514 -6696
rect 4344 -6731 4345 -6697
rect 4345 -6731 4513 -6697
rect 4513 -6731 4514 -6697
rect 4344 -6805 4514 -6731
rect 4344 -6839 4345 -6805
rect 4345 -6839 4513 -6805
rect 4513 -6839 4514 -6805
rect 4344 -6840 4514 -6839
rect 4716 -6697 4886 -6696
rect 4716 -6731 4717 -6697
rect 4717 -6731 4885 -6697
rect 4885 -6731 4886 -6697
rect 4716 -6805 4886 -6731
rect 4716 -6839 4717 -6805
rect 4717 -6839 4885 -6805
rect 4885 -6839 4886 -6805
rect 4716 -6840 4886 -6839
rect 5088 -6697 5258 -6696
rect 5088 -6731 5089 -6697
rect 5089 -6731 5257 -6697
rect 5257 -6731 5258 -6697
rect 5088 -6805 5258 -6731
rect 5088 -6839 5089 -6805
rect 5089 -6839 5257 -6805
rect 5257 -6839 5258 -6805
rect 5088 -6840 5258 -6839
rect 5460 -6697 5630 -6696
rect 5460 -6731 5461 -6697
rect 5461 -6731 5629 -6697
rect 5629 -6731 5630 -6697
rect 5460 -6805 5630 -6731
rect 5460 -6839 5461 -6805
rect 5461 -6839 5629 -6805
rect 5629 -6839 5630 -6805
rect 5460 -6840 5630 -6839
rect 5832 -6697 6002 -6696
rect 5832 -6731 5833 -6697
rect 5833 -6731 6001 -6697
rect 6001 -6731 6002 -6697
rect 5832 -6805 6002 -6731
rect 5832 -6839 5833 -6805
rect 5833 -6839 6001 -6805
rect 6001 -6839 6002 -6805
rect 5832 -6840 6002 -6839
rect 6204 -6697 6374 -6696
rect 6204 -6731 6205 -6697
rect 6205 -6731 6373 -6697
rect 6373 -6731 6374 -6697
rect 6204 -6805 6374 -6731
rect 6204 -6839 6205 -6805
rect 6205 -6839 6373 -6805
rect 6373 -6839 6374 -6805
rect 6204 -6840 6374 -6839
rect 6576 -6697 6746 -6696
rect 6576 -6731 6577 -6697
rect 6577 -6731 6745 -6697
rect 6745 -6731 6746 -6697
rect 6576 -6805 6746 -6731
rect 6576 -6839 6577 -6805
rect 6577 -6839 6745 -6805
rect 6745 -6839 6746 -6805
rect 6576 -6840 6746 -6839
rect 6948 -6697 7118 -6696
rect 6948 -6731 6949 -6697
rect 6949 -6731 7117 -6697
rect 7117 -6731 7118 -6697
rect 6948 -6805 7118 -6731
rect 6948 -6839 6949 -6805
rect 6949 -6839 7117 -6805
rect 7117 -6839 7118 -6805
rect 6948 -6840 7118 -6839
rect 7320 -6697 7490 -6696
rect 7320 -6731 7321 -6697
rect 7321 -6731 7489 -6697
rect 7489 -6731 7490 -6697
rect 7320 -6805 7490 -6731
rect 7320 -6839 7321 -6805
rect 7321 -6839 7489 -6805
rect 7489 -6839 7490 -6805
rect 7320 -6840 7490 -6839
rect 7692 -6697 7862 -6696
rect 7692 -6731 7693 -6697
rect 7693 -6731 7861 -6697
rect 7861 -6731 7862 -6697
rect 7692 -6805 7862 -6731
rect 7692 -6839 7693 -6805
rect 7693 -6839 7861 -6805
rect 7861 -6839 7862 -6805
rect 7692 -6840 7862 -6839
rect 8064 -6697 8234 -6696
rect 8064 -6731 8065 -6697
rect 8065 -6731 8233 -6697
rect 8233 -6731 8234 -6697
rect 8064 -6805 8234 -6731
rect 8064 -6839 8065 -6805
rect 8065 -6839 8233 -6805
rect 8233 -6839 8234 -6805
rect 8064 -6840 8234 -6839
rect 8436 -6697 8606 -6696
rect 8436 -6731 8437 -6697
rect 8437 -6731 8605 -6697
rect 8605 -6731 8606 -6697
rect 8436 -6805 8606 -6731
rect 8436 -6839 8437 -6805
rect 8437 -6839 8605 -6805
rect 8605 -6839 8606 -6805
rect 8436 -6840 8606 -6839
rect 8808 -6697 8978 -6696
rect 8808 -6731 8809 -6697
rect 8809 -6731 8977 -6697
rect 8977 -6731 8978 -6697
rect 8808 -6805 8978 -6731
rect 8808 -6839 8809 -6805
rect 8809 -6839 8977 -6805
rect 8977 -6839 8978 -6805
rect 8808 -6840 8978 -6839
rect 9180 -6697 9350 -6696
rect 9180 -6731 9181 -6697
rect 9181 -6731 9349 -6697
rect 9349 -6731 9350 -6697
rect 9180 -6805 9350 -6731
rect 9180 -6839 9181 -6805
rect 9181 -6839 9349 -6805
rect 9349 -6839 9350 -6805
rect 9180 -6840 9350 -6839
rect 9552 -6697 9722 -6696
rect 9552 -6731 9553 -6697
rect 9553 -6731 9721 -6697
rect 9721 -6731 9722 -6697
rect 9552 -6805 9722 -6731
rect 9552 -6839 9553 -6805
rect 9553 -6839 9721 -6805
rect 9721 -6839 9722 -6805
rect 9552 -6840 9722 -6839
rect 996 -7115 1166 -7114
rect 996 -7149 997 -7115
rect 997 -7149 1165 -7115
rect 1165 -7149 1166 -7115
rect 996 -7223 1166 -7149
rect 996 -7257 997 -7223
rect 997 -7257 1165 -7223
rect 1165 -7257 1166 -7223
rect 996 -7258 1166 -7257
rect 1368 -7115 1538 -7114
rect 1368 -7149 1369 -7115
rect 1369 -7149 1537 -7115
rect 1537 -7149 1538 -7115
rect 1368 -7223 1538 -7149
rect 1368 -7257 1369 -7223
rect 1369 -7257 1537 -7223
rect 1537 -7257 1538 -7223
rect 1368 -7258 1538 -7257
rect 1740 -7115 1910 -7114
rect 1740 -7149 1741 -7115
rect 1741 -7149 1909 -7115
rect 1909 -7149 1910 -7115
rect 1740 -7223 1910 -7149
rect 1740 -7257 1741 -7223
rect 1741 -7257 1909 -7223
rect 1909 -7257 1910 -7223
rect 1740 -7258 1910 -7257
rect 2112 -7115 2282 -7114
rect 2112 -7149 2113 -7115
rect 2113 -7149 2281 -7115
rect 2281 -7149 2282 -7115
rect 2112 -7223 2282 -7149
rect 2112 -7257 2113 -7223
rect 2113 -7257 2281 -7223
rect 2281 -7257 2282 -7223
rect 2112 -7258 2282 -7257
rect 2484 -7115 2654 -7114
rect 2484 -7149 2485 -7115
rect 2485 -7149 2653 -7115
rect 2653 -7149 2654 -7115
rect 2484 -7223 2654 -7149
rect 2484 -7257 2485 -7223
rect 2485 -7257 2653 -7223
rect 2653 -7257 2654 -7223
rect 2484 -7258 2654 -7257
rect 2856 -7115 3026 -7114
rect 2856 -7149 2857 -7115
rect 2857 -7149 3025 -7115
rect 3025 -7149 3026 -7115
rect 2856 -7223 3026 -7149
rect 2856 -7257 2857 -7223
rect 2857 -7257 3025 -7223
rect 3025 -7257 3026 -7223
rect 2856 -7258 3026 -7257
rect 3228 -7115 3398 -7114
rect 3228 -7149 3229 -7115
rect 3229 -7149 3397 -7115
rect 3397 -7149 3398 -7115
rect 3228 -7223 3398 -7149
rect 3228 -7257 3229 -7223
rect 3229 -7257 3397 -7223
rect 3397 -7257 3398 -7223
rect 3228 -7258 3398 -7257
rect 3600 -7115 3770 -7114
rect 3600 -7149 3601 -7115
rect 3601 -7149 3769 -7115
rect 3769 -7149 3770 -7115
rect 3600 -7223 3770 -7149
rect 3600 -7257 3601 -7223
rect 3601 -7257 3769 -7223
rect 3769 -7257 3770 -7223
rect 3600 -7258 3770 -7257
rect 3972 -7115 4142 -7114
rect 3972 -7149 3973 -7115
rect 3973 -7149 4141 -7115
rect 4141 -7149 4142 -7115
rect 3972 -7223 4142 -7149
rect 3972 -7257 3973 -7223
rect 3973 -7257 4141 -7223
rect 4141 -7257 4142 -7223
rect 3972 -7258 4142 -7257
rect 4344 -7115 4514 -7114
rect 4344 -7149 4345 -7115
rect 4345 -7149 4513 -7115
rect 4513 -7149 4514 -7115
rect 4344 -7223 4514 -7149
rect 4344 -7257 4345 -7223
rect 4345 -7257 4513 -7223
rect 4513 -7257 4514 -7223
rect 4344 -7258 4514 -7257
rect 4716 -7115 4886 -7114
rect 4716 -7149 4717 -7115
rect 4717 -7149 4885 -7115
rect 4885 -7149 4886 -7115
rect 4716 -7223 4886 -7149
rect 4716 -7257 4717 -7223
rect 4717 -7257 4885 -7223
rect 4885 -7257 4886 -7223
rect 4716 -7258 4886 -7257
rect 5088 -7115 5258 -7114
rect 5088 -7149 5089 -7115
rect 5089 -7149 5257 -7115
rect 5257 -7149 5258 -7115
rect 5088 -7223 5258 -7149
rect 5088 -7257 5089 -7223
rect 5089 -7257 5257 -7223
rect 5257 -7257 5258 -7223
rect 5088 -7258 5258 -7257
rect 5460 -7115 5630 -7114
rect 5460 -7149 5461 -7115
rect 5461 -7149 5629 -7115
rect 5629 -7149 5630 -7115
rect 5460 -7223 5630 -7149
rect 5460 -7257 5461 -7223
rect 5461 -7257 5629 -7223
rect 5629 -7257 5630 -7223
rect 5460 -7258 5630 -7257
rect 5832 -7115 6002 -7114
rect 5832 -7149 5833 -7115
rect 5833 -7149 6001 -7115
rect 6001 -7149 6002 -7115
rect 5832 -7223 6002 -7149
rect 5832 -7257 5833 -7223
rect 5833 -7257 6001 -7223
rect 6001 -7257 6002 -7223
rect 5832 -7258 6002 -7257
rect 6204 -7115 6374 -7114
rect 6204 -7149 6205 -7115
rect 6205 -7149 6373 -7115
rect 6373 -7149 6374 -7115
rect 6204 -7223 6374 -7149
rect 6204 -7257 6205 -7223
rect 6205 -7257 6373 -7223
rect 6373 -7257 6374 -7223
rect 6204 -7258 6374 -7257
rect 6576 -7115 6746 -7114
rect 6576 -7149 6577 -7115
rect 6577 -7149 6745 -7115
rect 6745 -7149 6746 -7115
rect 6576 -7223 6746 -7149
rect 6576 -7257 6577 -7223
rect 6577 -7257 6745 -7223
rect 6745 -7257 6746 -7223
rect 6576 -7258 6746 -7257
rect 6948 -7115 7118 -7114
rect 6948 -7149 6949 -7115
rect 6949 -7149 7117 -7115
rect 7117 -7149 7118 -7115
rect 6948 -7223 7118 -7149
rect 6948 -7257 6949 -7223
rect 6949 -7257 7117 -7223
rect 7117 -7257 7118 -7223
rect 6948 -7258 7118 -7257
rect 7320 -7115 7490 -7114
rect 7320 -7149 7321 -7115
rect 7321 -7149 7489 -7115
rect 7489 -7149 7490 -7115
rect 7320 -7223 7490 -7149
rect 7320 -7257 7321 -7223
rect 7321 -7257 7489 -7223
rect 7489 -7257 7490 -7223
rect 7320 -7258 7490 -7257
rect 7692 -7115 7862 -7114
rect 7692 -7149 7693 -7115
rect 7693 -7149 7861 -7115
rect 7861 -7149 7862 -7115
rect 7692 -7223 7862 -7149
rect 7692 -7257 7693 -7223
rect 7693 -7257 7861 -7223
rect 7861 -7257 7862 -7223
rect 7692 -7258 7862 -7257
rect 8064 -7115 8234 -7114
rect 8064 -7149 8065 -7115
rect 8065 -7149 8233 -7115
rect 8233 -7149 8234 -7115
rect 8064 -7223 8234 -7149
rect 8064 -7257 8065 -7223
rect 8065 -7257 8233 -7223
rect 8233 -7257 8234 -7223
rect 8064 -7258 8234 -7257
rect 8436 -7115 8606 -7114
rect 8436 -7149 8437 -7115
rect 8437 -7149 8605 -7115
rect 8605 -7149 8606 -7115
rect 8436 -7223 8606 -7149
rect 8436 -7257 8437 -7223
rect 8437 -7257 8605 -7223
rect 8605 -7257 8606 -7223
rect 8436 -7258 8606 -7257
rect 8808 -7115 8978 -7114
rect 8808 -7149 8809 -7115
rect 8809 -7149 8977 -7115
rect 8977 -7149 8978 -7115
rect 8808 -7223 8978 -7149
rect 8808 -7257 8809 -7223
rect 8809 -7257 8977 -7223
rect 8977 -7257 8978 -7223
rect 8808 -7258 8978 -7257
rect 9180 -7115 9350 -7114
rect 9180 -7149 9181 -7115
rect 9181 -7149 9349 -7115
rect 9349 -7149 9350 -7115
rect 9180 -7223 9350 -7149
rect 9180 -7257 9181 -7223
rect 9181 -7257 9349 -7223
rect 9349 -7257 9350 -7223
rect 9180 -7258 9350 -7257
rect 9552 -7115 9722 -7114
rect 9552 -7149 9553 -7115
rect 9553 -7149 9721 -7115
rect 9721 -7149 9722 -7115
rect 9552 -7223 9722 -7149
rect 9552 -7257 9553 -7223
rect 9553 -7257 9721 -7223
rect 9721 -7257 9722 -7223
rect 9552 -7258 9722 -7257
rect 996 -7533 1166 -7522
rect 996 -7567 997 -7533
rect 997 -7567 1165 -7533
rect 1165 -7567 1166 -7533
rect 996 -7578 1166 -7567
rect 1368 -7533 1538 -7522
rect 1368 -7567 1369 -7533
rect 1369 -7567 1537 -7533
rect 1537 -7567 1538 -7533
rect 1368 -7578 1538 -7567
rect 1740 -7533 1910 -7522
rect 1740 -7567 1741 -7533
rect 1741 -7567 1909 -7533
rect 1909 -7567 1910 -7533
rect 1740 -7578 1910 -7567
rect 2112 -7533 2282 -7522
rect 2112 -7567 2113 -7533
rect 2113 -7567 2281 -7533
rect 2281 -7567 2282 -7533
rect 2112 -7578 2282 -7567
rect 2484 -7533 2654 -7522
rect 2484 -7567 2485 -7533
rect 2485 -7567 2653 -7533
rect 2653 -7567 2654 -7533
rect 2484 -7578 2654 -7567
rect 2856 -7533 3026 -7522
rect 2856 -7567 2857 -7533
rect 2857 -7567 3025 -7533
rect 3025 -7567 3026 -7533
rect 2856 -7578 3026 -7567
rect 3228 -7533 3398 -7522
rect 3228 -7567 3229 -7533
rect 3229 -7567 3397 -7533
rect 3397 -7567 3398 -7533
rect 3228 -7578 3398 -7567
rect 3600 -7533 3770 -7522
rect 3600 -7567 3601 -7533
rect 3601 -7567 3769 -7533
rect 3769 -7567 3770 -7533
rect 3600 -7578 3770 -7567
rect 3972 -7533 4142 -7522
rect 3972 -7567 3973 -7533
rect 3973 -7567 4141 -7533
rect 4141 -7567 4142 -7533
rect 3972 -7578 4142 -7567
rect 4344 -7533 4514 -7522
rect 4344 -7567 4345 -7533
rect 4345 -7567 4513 -7533
rect 4513 -7567 4514 -7533
rect 4344 -7578 4514 -7567
rect 4716 -7533 4886 -7522
rect 4716 -7567 4717 -7533
rect 4717 -7567 4885 -7533
rect 4885 -7567 4886 -7533
rect 4716 -7578 4886 -7567
rect 5088 -7533 5258 -7522
rect 5088 -7567 5089 -7533
rect 5089 -7567 5257 -7533
rect 5257 -7567 5258 -7533
rect 5088 -7578 5258 -7567
rect 5460 -7533 5630 -7522
rect 5460 -7567 5461 -7533
rect 5461 -7567 5629 -7533
rect 5629 -7567 5630 -7533
rect 5460 -7578 5630 -7567
rect 5832 -7533 6002 -7522
rect 5832 -7567 5833 -7533
rect 5833 -7567 6001 -7533
rect 6001 -7567 6002 -7533
rect 5832 -7578 6002 -7567
rect 6204 -7533 6374 -7522
rect 6204 -7567 6205 -7533
rect 6205 -7567 6373 -7533
rect 6373 -7567 6374 -7533
rect 6204 -7578 6374 -7567
rect 6576 -7533 6746 -7522
rect 6576 -7567 6577 -7533
rect 6577 -7567 6745 -7533
rect 6745 -7567 6746 -7533
rect 6576 -7578 6746 -7567
rect 6948 -7533 7118 -7522
rect 6948 -7567 6949 -7533
rect 6949 -7567 7117 -7533
rect 7117 -7567 7118 -7533
rect 6948 -7578 7118 -7567
rect 7320 -7533 7490 -7522
rect 7320 -7567 7321 -7533
rect 7321 -7567 7489 -7533
rect 7489 -7567 7490 -7533
rect 7320 -7578 7490 -7567
rect 7692 -7533 7862 -7522
rect 7692 -7567 7693 -7533
rect 7693 -7567 7861 -7533
rect 7861 -7567 7862 -7533
rect 7692 -7578 7862 -7567
rect 8064 -7533 8234 -7522
rect 8064 -7567 8065 -7533
rect 8065 -7567 8233 -7533
rect 8233 -7567 8234 -7533
rect 8064 -7578 8234 -7567
rect 8436 -7533 8606 -7522
rect 8436 -7567 8437 -7533
rect 8437 -7567 8605 -7533
rect 8605 -7567 8606 -7533
rect 8436 -7578 8606 -7567
rect 8808 -7533 8978 -7522
rect 8808 -7567 8809 -7533
rect 8809 -7567 8977 -7533
rect 8977 -7567 8978 -7533
rect 8808 -7578 8978 -7567
rect 9180 -7533 9350 -7522
rect 9180 -7567 9181 -7533
rect 9181 -7567 9349 -7533
rect 9349 -7567 9350 -7533
rect 9180 -7578 9350 -7567
rect 9552 -7533 9722 -7522
rect 9552 -7567 9553 -7533
rect 9553 -7567 9721 -7533
rect 9721 -7567 9722 -7533
rect 9552 -7578 9722 -7567
rect 816 -7932 1016 -7732
rect 1540 -7932 1740 -7732
rect 2284 -7932 2484 -7732
rect 3028 -7932 3228 -7732
rect 3772 -7932 3972 -7732
rect 4516 -7932 4716 -7732
rect 5260 -7932 5460 -7732
rect 6004 -7932 6204 -7732
rect 6748 -7932 6948 -7732
rect 7492 -7932 7692 -7732
rect 8236 -7932 8436 -7732
rect 8980 -7932 9180 -7732
rect 9724 -7932 9924 -7732
<< metal2 >>
rect -322 1514 -122 1524
rect -322 1304 -122 1314
rect 422 1514 622 1524
rect 422 1304 622 1314
rect 1166 1514 1366 1524
rect 1166 1304 1366 1314
rect 1910 1514 2110 1524
rect 1910 1304 2110 1314
rect 2654 1514 2854 1524
rect 2654 1304 2854 1314
rect 3398 1514 3598 1524
rect 3398 1304 3598 1314
rect 4142 1514 4342 1524
rect 4142 1304 4342 1314
rect 4886 1514 5086 1524
rect 4886 1304 5086 1314
rect 5258 1514 5458 1524
rect 5258 1304 5458 1314
rect 6002 1514 6202 1524
rect 6002 1304 6202 1314
rect 6746 1514 6946 1524
rect 6746 1304 6946 1314
rect 7490 1514 7690 1524
rect 7490 1304 7690 1314
rect 8234 1514 8434 1524
rect 8234 1304 8434 1314
rect 8978 1514 9178 1524
rect 8978 1304 9178 1314
rect 9722 1514 9922 1524
rect 9722 1304 9922 1314
rect 10466 1514 10666 1524
rect 10466 1304 10666 1314
rect 11210 1514 11410 1524
rect 11210 1304 11410 1314
rect -492 1126 11220 1136
rect -322 1066 -120 1126
rect 50 1066 252 1126
rect 422 1066 624 1126
rect 794 1066 996 1126
rect 1166 1066 1368 1126
rect 1538 1066 1740 1126
rect 1910 1066 2112 1126
rect 2282 1066 2484 1126
rect 2654 1066 2856 1126
rect 3026 1066 3228 1126
rect 3398 1066 3600 1126
rect 3770 1066 3972 1126
rect 4142 1066 4344 1126
rect 4514 1066 4716 1126
rect 4886 1066 5088 1126
rect 5258 1066 5460 1126
rect 5630 1066 5832 1126
rect 6002 1066 6204 1126
rect 6374 1066 6576 1126
rect 6746 1066 6948 1126
rect 7118 1066 7320 1126
rect 7490 1066 7692 1126
rect 7862 1066 8064 1126
rect 8234 1066 8436 1126
rect 8606 1066 8808 1126
rect 8978 1066 9180 1126
rect 9350 1066 9552 1126
rect 9722 1066 9924 1126
rect 10094 1066 10296 1126
rect 10466 1066 10668 1126
rect 10838 1066 11040 1126
rect 11210 1066 11220 1126
rect -492 1056 11220 1066
rect -492 586 11210 596
rect -322 442 -120 586
rect 50 442 252 586
rect 422 442 624 586
rect 794 442 996 586
rect 1166 442 1368 586
rect 1538 442 1740 586
rect 1910 442 2112 586
rect 2282 442 2484 586
rect 2654 442 2856 586
rect 3026 442 3228 586
rect 3398 442 3600 586
rect 3770 442 3972 586
rect 4142 442 4344 586
rect 4514 442 4716 586
rect 4886 442 5088 586
rect 5258 442 5460 586
rect 5630 442 5832 586
rect 6002 442 6204 586
rect 6374 442 6576 586
rect 6746 442 6948 586
rect 7118 442 7320 586
rect 7490 442 7692 586
rect 7862 442 8064 586
rect 8234 442 8436 586
rect 8606 442 8808 586
rect 8978 442 9180 586
rect 9350 442 9552 586
rect 9722 442 9924 586
rect 10094 442 10296 586
rect 10466 442 10668 586
rect 10838 442 11040 586
rect -492 432 11210 442
rect -492 -50 11210 -40
rect -322 -194 -120 -50
rect 50 -194 252 -50
rect 422 -194 624 -50
rect 794 -194 996 -50
rect 1166 -194 1368 -50
rect 1538 -194 1740 -50
rect 1910 -194 2112 -50
rect 2282 -194 2484 -50
rect 2654 -194 2856 -50
rect 3026 -194 3228 -50
rect 3398 -194 3600 -50
rect 3770 -194 3972 -50
rect 4142 -194 4344 -50
rect 4514 -194 4716 -50
rect 4886 -194 5088 -50
rect 5258 -194 5460 -50
rect 5630 -194 5832 -50
rect 6002 -194 6204 -50
rect 6374 -194 6576 -50
rect 6746 -194 6948 -50
rect 7118 -194 7320 -50
rect 7490 -194 7692 -50
rect 7862 -194 8064 -50
rect 8234 -194 8436 -50
rect 8606 -194 8808 -50
rect 8978 -194 9180 -50
rect 9350 -194 9552 -50
rect 9722 -194 9924 -50
rect 10094 -194 10296 -50
rect 10466 -194 10668 -50
rect 10838 -194 11040 -50
rect -492 -204 11210 -194
rect -492 -674 11210 -664
rect -322 -734 -120 -674
rect 50 -734 252 -674
rect 422 -734 624 -674
rect 794 -734 996 -674
rect 1166 -734 1368 -674
rect 1538 -734 1740 -674
rect 1910 -734 2112 -674
rect 2282 -734 2484 -674
rect 2654 -734 2856 -674
rect 3026 -734 3228 -674
rect 3398 -734 3600 -674
rect 3770 -734 3972 -674
rect 4142 -734 4344 -674
rect 4514 -734 4716 -674
rect 4886 -734 5088 -674
rect 5258 -734 5460 -674
rect 5630 -734 5832 -674
rect 6002 -734 6204 -674
rect 6374 -734 6576 -674
rect 6746 -734 6948 -674
rect 7118 -734 7320 -674
rect 7490 -734 7692 -674
rect 7862 -734 8064 -674
rect 8234 -734 8436 -674
rect 8606 -734 8808 -674
rect 8978 -734 9180 -674
rect 9350 -734 9552 -674
rect 9722 -734 9924 -674
rect 10094 -734 10296 -674
rect 10466 -734 10668 -674
rect 10838 -734 11040 -674
rect -492 -744 11210 -734
rect 5592 -1042 11082 -1032
rect 516 -1160 3584 -1062
rect 1182 -1250 1352 -1160
rect 3414 -1250 3584 -1160
rect 996 -1260 1538 -1250
rect 1166 -1324 1368 -1260
rect 996 -1334 1538 -1324
rect 1740 -1260 3026 -1250
rect 1910 -1324 2112 -1260
rect 2282 -1324 2484 -1260
rect 2654 -1324 2856 -1260
rect 1740 -1334 3026 -1324
rect 3228 -1260 3770 -1250
rect 3398 -1324 3600 -1260
rect 5874 -1314 6336 -1042
rect 6618 -1314 7080 -1042
rect 7362 -1314 7824 -1042
rect 8106 -1314 8568 -1042
rect 8850 -1314 9312 -1042
rect 9594 -1314 10056 -1042
rect 10338 -1314 10800 -1042
rect 5592 -1324 11082 -1314
rect 3228 -1334 3770 -1324
rect 1240 -2192 1294 -1334
rect 1984 -2192 2038 -1334
rect 2728 -2192 2782 -1334
rect 3472 -2192 3526 -1334
rect 996 -2202 1538 -2192
rect 1166 -2346 1368 -2202
rect 996 -2356 1538 -2346
rect 1740 -2202 3026 -2192
rect 1910 -2346 2112 -2202
rect 2282 -2346 2484 -2202
rect 2654 -2346 2856 -2202
rect 1740 -2356 3026 -2346
rect 3228 -2202 3770 -2192
rect 3398 -2346 3600 -2202
rect 3228 -2356 3770 -2346
rect 1240 -3228 1294 -2356
rect 1984 -3228 2038 -2356
rect 2728 -3228 2782 -2356
rect 3472 -3228 3526 -2356
rect 6012 -2816 6294 -2806
rect 6012 -3098 6294 -3088
rect 996 -3238 1538 -3228
rect 1166 -3382 1368 -3238
rect 996 -3392 1538 -3382
rect 1740 -3238 3026 -3228
rect 1910 -3382 2112 -3238
rect 2282 -3382 2484 -3238
rect 2654 -3382 2856 -3238
rect 1740 -3392 3026 -3382
rect 3228 -3238 3770 -3228
rect 3398 -3382 3600 -3238
rect 3228 -3392 3770 -3382
rect 1240 -4264 1294 -3392
rect 1984 -4264 2038 -3392
rect 2728 -4264 2782 -3392
rect 3472 -4264 3526 -3392
rect 5686 -3528 5846 -3518
rect 5686 -3700 5846 -3690
rect 5686 -3928 5846 -3918
rect 5686 -4100 5846 -4090
rect 996 -4274 1538 -4264
rect 1166 -4418 1368 -4274
rect 996 -4428 1538 -4418
rect 1740 -4274 3026 -4264
rect 1910 -4418 2112 -4274
rect 2282 -4418 2484 -4274
rect 2654 -4418 2856 -4274
rect 1740 -4428 3026 -4418
rect 3228 -4274 3770 -4264
rect 3398 -4418 3600 -4274
rect 3228 -4428 3770 -4418
rect 5686 -4328 5846 -4318
rect 1240 -5290 1294 -4428
rect 1984 -5290 2038 -4428
rect 2728 -5290 2782 -4428
rect 3472 -5290 3526 -4428
rect 5686 -4500 5846 -4490
rect 4102 -5224 9602 -5214
rect 996 -5300 1538 -5290
rect 1166 -5354 1368 -5300
rect 996 -5364 1538 -5354
rect 1740 -5300 3026 -5290
rect 1910 -5354 2112 -5300
rect 2282 -5354 2484 -5300
rect 2654 -5354 2856 -5300
rect 1740 -5364 3026 -5354
rect 3228 -5300 3770 -5290
rect 3398 -5354 3600 -5300
rect 3228 -5364 3770 -5354
rect 1926 -5464 2096 -5364
rect 2670 -5464 2840 -5364
rect 516 -5562 2840 -5464
rect 4384 -5388 4846 -5224
rect 4102 -5506 4384 -5496
rect 5128 -5388 5590 -5224
rect 4846 -5506 5128 -5496
rect 5872 -5388 6334 -5224
rect 5590 -5506 5872 -5496
rect 6616 -5388 7078 -5224
rect 5986 -5512 6264 -5502
rect 6334 -5506 6616 -5496
rect 7360 -5388 7822 -5224
rect 7078 -5506 7360 -5496
rect 8104 -5388 8566 -5224
rect 7822 -5506 8104 -5496
rect 8848 -5388 9310 -5224
rect 8566 -5506 8848 -5496
rect 9592 -5388 9602 -5224
rect 9310 -5506 9592 -5496
rect 1976 -5640 5986 -5630
rect 2790 -5774 5986 -5640
rect 2790 -5820 3956 -5774
rect 6264 -5774 6278 -5630
rect 5986 -5796 6264 -5786
rect 1976 -5830 3956 -5820
rect 3830 -5948 3956 -5830
rect 996 -5958 3782 -5948
rect 1166 -6014 1368 -5958
rect 1538 -6014 1740 -5958
rect 1910 -6014 2112 -5958
rect 2282 -6014 2484 -5958
rect 2654 -6014 2856 -5958
rect 3026 -6014 3228 -5958
rect 3398 -6014 3600 -5958
rect 3770 -6014 3782 -5958
rect 996 -6024 3782 -6014
rect 3830 -5958 9722 -5948
rect 3830 -6014 3972 -5958
rect 4142 -6014 4344 -5958
rect 4514 -6014 4716 -5958
rect 4886 -6014 5088 -5958
rect 5258 -6014 5460 -5958
rect 5630 -6014 5832 -5958
rect 6002 -6014 6204 -5958
rect 6374 -6014 6576 -5958
rect 6746 -6014 6948 -5958
rect 7118 -6014 7320 -5958
rect 7490 -6014 7692 -5958
rect 7862 -6014 8064 -5958
rect 8234 -6014 8436 -5958
rect 8606 -6014 8808 -5958
rect 8978 -6014 9180 -5958
rect 9350 -6014 9552 -5958
rect 3830 -6024 9722 -6014
rect 3830 -6268 3956 -6024
rect 996 -6278 3782 -6268
rect 1166 -6422 1368 -6278
rect 1538 -6422 1740 -6278
rect 1910 -6422 2112 -6278
rect 2282 -6422 2484 -6278
rect 2654 -6422 2856 -6278
rect 3026 -6422 3228 -6278
rect 3398 -6422 3600 -6278
rect 3770 -6422 3782 -6278
rect 996 -6432 3782 -6422
rect 3830 -6278 9722 -6268
rect 3830 -6422 3972 -6278
rect 4142 -6422 4344 -6278
rect 4514 -6422 4716 -6278
rect 4886 -6422 5088 -6278
rect 5258 -6422 5460 -6278
rect 5630 -6422 5832 -6278
rect 6002 -6422 6204 -6278
rect 6374 -6422 6576 -6278
rect 6746 -6422 6948 -6278
rect 7118 -6422 7320 -6278
rect 7490 -6422 7692 -6278
rect 7862 -6422 8064 -6278
rect 8234 -6422 8436 -6278
rect 8606 -6422 8808 -6278
rect 8978 -6422 9180 -6278
rect 9350 -6422 9552 -6278
rect 3830 -6432 9722 -6422
rect 3830 -6686 3956 -6432
rect 996 -6696 3782 -6686
rect 1166 -6840 1368 -6696
rect 1538 -6840 1740 -6696
rect 1910 -6840 2112 -6696
rect 2282 -6840 2484 -6696
rect 2654 -6840 2856 -6696
rect 3026 -6840 3228 -6696
rect 3398 -6840 3600 -6696
rect 3770 -6840 3782 -6696
rect 996 -6850 3782 -6840
rect 3830 -6696 9722 -6686
rect 3830 -6840 3972 -6696
rect 4142 -6840 4344 -6696
rect 4514 -6840 4716 -6696
rect 4886 -6840 5088 -6696
rect 5258 -6840 5460 -6696
rect 5630 -6840 5832 -6696
rect 6002 -6840 6204 -6696
rect 6374 -6840 6576 -6696
rect 6746 -6840 6948 -6696
rect 7118 -6840 7320 -6696
rect 7490 -6840 7692 -6696
rect 7862 -6840 8064 -6696
rect 8234 -6840 8436 -6696
rect 8606 -6840 8808 -6696
rect 8978 -6840 9180 -6696
rect 9350 -6840 9552 -6696
rect 3830 -6850 9722 -6840
rect 3830 -7104 3956 -6850
rect 996 -7114 3782 -7104
rect 1166 -7258 1368 -7114
rect 1538 -7258 1740 -7114
rect 1910 -7258 2112 -7114
rect 2282 -7258 2484 -7114
rect 2654 -7258 2856 -7114
rect 3026 -7258 3228 -7114
rect 3398 -7258 3600 -7114
rect 3770 -7258 3782 -7114
rect 996 -7268 3782 -7258
rect 3830 -7114 9722 -7104
rect 3830 -7258 3972 -7114
rect 4142 -7258 4344 -7114
rect 4514 -7258 4716 -7114
rect 4886 -7258 5088 -7114
rect 5258 -7258 5460 -7114
rect 5630 -7258 5832 -7114
rect 6002 -7258 6204 -7114
rect 6374 -7258 6576 -7114
rect 6746 -7258 6948 -7114
rect 7118 -7258 7320 -7114
rect 7490 -7258 7692 -7114
rect 7862 -7258 8064 -7114
rect 8234 -7258 8436 -7114
rect 8606 -7258 8808 -7114
rect 8978 -7258 9180 -7114
rect 9350 -7258 9552 -7114
rect 3830 -7268 9722 -7258
rect 3830 -7512 3956 -7268
rect 996 -7522 3782 -7512
rect 1166 -7578 1368 -7522
rect 1538 -7578 1740 -7522
rect 1910 -7578 2112 -7522
rect 2282 -7578 2484 -7522
rect 2654 -7578 2856 -7522
rect 3026 -7578 3228 -7522
rect 3398 -7578 3600 -7522
rect 3770 -7578 3782 -7522
rect 996 -7588 3782 -7578
rect 3830 -7522 9722 -7512
rect 3830 -7578 3972 -7522
rect 4142 -7578 4344 -7522
rect 4514 -7578 4716 -7522
rect 4886 -7578 5088 -7522
rect 5258 -7578 5460 -7522
rect 5630 -7578 5832 -7522
rect 6002 -7578 6204 -7522
rect 6374 -7578 6576 -7522
rect 6746 -7578 6948 -7522
rect 7118 -7578 7320 -7522
rect 7490 -7578 7692 -7522
rect 7862 -7578 8064 -7522
rect 8234 -7578 8436 -7522
rect 8606 -7578 8808 -7522
rect 8978 -7578 9180 -7522
rect 9350 -7578 9552 -7522
rect 3830 -7588 9722 -7578
rect 816 -7732 1016 -7722
rect 816 -7942 1016 -7932
rect 1540 -7732 1740 -7722
rect 1540 -7942 1740 -7932
rect 2284 -7732 2484 -7722
rect 2284 -7942 2484 -7932
rect 3028 -7732 3228 -7722
rect 3028 -7942 3228 -7932
rect 3772 -7732 3972 -7722
rect 3772 -7942 3972 -7932
rect 4516 -7732 4716 -7722
rect 4516 -7942 4716 -7932
rect 5260 -7732 5460 -7722
rect 5260 -7942 5460 -7932
rect 6004 -7732 6204 -7722
rect 6004 -7942 6204 -7932
rect 6748 -7732 6948 -7722
rect 6748 -7942 6948 -7932
rect 7492 -7732 7692 -7722
rect 7492 -7942 7692 -7932
rect 8236 -7732 8436 -7722
rect 8236 -7942 8436 -7932
rect 8980 -7732 9180 -7722
rect 8980 -7942 9180 -7932
rect 9724 -7732 9924 -7722
rect 9724 -7942 9924 -7932
<< via2 >>
rect -322 1314 -122 1514
rect 422 1314 622 1514
rect 1166 1314 1366 1514
rect 1910 1314 2110 1514
rect 2654 1314 2854 1514
rect 3398 1314 3598 1514
rect 4142 1314 4342 1514
rect 4886 1314 5086 1514
rect 5258 1314 5458 1514
rect 6002 1314 6202 1514
rect 6746 1314 6946 1514
rect 7490 1314 7690 1514
rect 8234 1314 8434 1514
rect 8978 1314 9178 1514
rect 9722 1314 9922 1514
rect 10466 1314 10666 1514
rect 11210 1314 11410 1514
rect 7080 -1314 7362 -1042
rect 7824 -1314 8106 -1042
rect 8568 -1314 8850 -1042
rect 9312 -1314 9594 -1042
rect 6012 -3088 6294 -2816
rect 5686 -3690 5846 -3528
rect 5686 -4090 5846 -3928
rect 5686 -4490 5846 -4328
rect 7078 -5496 7360 -5224
rect 7822 -5496 8104 -5224
rect 8566 -5496 8848 -5224
rect 9310 -5496 9592 -5224
rect 816 -7932 1016 -7732
rect 1540 -7932 1740 -7732
rect 2284 -7932 2484 -7732
rect 3028 -7932 3228 -7732
rect 3772 -7932 3972 -7732
rect 4516 -7932 4716 -7732
rect 5260 -7932 5460 -7732
rect 6004 -7932 6204 -7732
rect 6748 -7932 6948 -7732
rect 7492 -7932 7692 -7732
rect 8236 -7932 8436 -7732
rect 8980 -7932 9180 -7732
rect 9724 -7932 9924 -7732
<< metal3 >>
rect -332 1514 -112 1519
rect -332 1314 -322 1514
rect -122 1314 -112 1514
rect -332 1309 -112 1314
rect 412 1514 632 1519
rect 412 1314 422 1514
rect 622 1314 632 1514
rect 412 1309 632 1314
rect 1156 1514 1376 1519
rect 1156 1314 1166 1514
rect 1366 1314 1376 1514
rect 1156 1309 1376 1314
rect 1900 1514 2120 1519
rect 1900 1314 1910 1514
rect 2110 1314 2120 1514
rect 1900 1309 2120 1314
rect 2644 1514 2864 1519
rect 2644 1314 2654 1514
rect 2854 1314 2864 1514
rect 2644 1309 2864 1314
rect 3388 1514 3608 1519
rect 3388 1314 3398 1514
rect 3598 1314 3608 1514
rect 3388 1309 3608 1314
rect 4132 1514 4352 1519
rect 4132 1314 4142 1514
rect 4342 1314 4352 1514
rect 4132 1309 4352 1314
rect 4876 1514 5096 1519
rect 4876 1314 4886 1514
rect 5086 1314 5096 1514
rect 4876 1309 5096 1314
rect 5248 1514 5468 1519
rect 5248 1314 5258 1514
rect 5458 1314 5468 1514
rect 5248 1309 5468 1314
rect 5992 1514 6212 1519
rect 5992 1314 6002 1514
rect 6202 1314 6212 1514
rect 5992 1309 6212 1314
rect 6736 1514 6956 1519
rect 6736 1314 6746 1514
rect 6946 1314 6956 1514
rect 6736 1309 6956 1314
rect 7480 1514 7700 1519
rect 7480 1314 7490 1514
rect 7690 1314 7700 1514
rect 7480 1309 7700 1314
rect 8224 1514 8444 1519
rect 8224 1314 8234 1514
rect 8434 1314 8444 1514
rect 8224 1309 8444 1314
rect 8968 1514 9188 1519
rect 8968 1314 8978 1514
rect 9178 1314 9188 1514
rect 8968 1309 9188 1314
rect 9712 1514 9932 1519
rect 9712 1314 9722 1514
rect 9922 1314 9932 1514
rect 9712 1309 9932 1314
rect 10456 1514 10676 1519
rect 10456 1314 10466 1514
rect 10666 1314 10676 1514
rect 10456 1309 10676 1314
rect 11200 1514 11420 1519
rect 11200 1314 11210 1514
rect 11410 1314 11420 1514
rect 11200 1309 11420 1314
rect 7070 -1042 7372 -1037
rect 7070 -1314 7080 -1042
rect 7362 -1314 7372 -1042
rect 7070 -1556 7372 -1314
rect 7814 -1042 8116 -1037
rect 7814 -1314 7824 -1042
rect 8106 -1314 8116 -1042
rect 7814 -1556 8116 -1314
rect 8558 -1042 8860 -1037
rect 8558 -1314 8568 -1042
rect 8850 -1314 8860 -1042
rect 8558 -1556 8860 -1314
rect 9302 -1042 9604 -1037
rect 9302 -1314 9312 -1042
rect 9594 -1314 9604 -1042
rect 9302 -1556 9604 -1314
rect 6808 -2714 9792 -1556
rect 6002 -2816 6304 -2811
rect 6002 -3088 6012 -2816
rect 6294 -3088 6304 -2816
rect 6002 -3093 6304 -3088
rect 6808 -3454 10304 -2714
rect 5676 -3528 5856 -3523
rect 5676 -3690 5686 -3528
rect 5846 -3690 5856 -3528
rect 5676 -3695 5856 -3690
rect 5676 -3928 5856 -3923
rect 5676 -4090 5686 -3928
rect 5846 -4090 5856 -3928
rect 5676 -4095 5856 -4090
rect 5676 -4328 5856 -4323
rect 5676 -4490 5686 -4328
rect 5846 -4490 5856 -4328
rect 5676 -4495 5856 -4490
rect 6808 -4556 9792 -3454
rect 7068 -5224 7370 -4556
rect 7068 -5496 7078 -5224
rect 7360 -5496 7370 -5224
rect 7068 -5501 7370 -5496
rect 7812 -5224 8114 -4556
rect 7812 -5496 7822 -5224
rect 8104 -5496 8114 -5224
rect 7812 -5501 8114 -5496
rect 8556 -5224 8858 -4556
rect 8556 -5496 8566 -5224
rect 8848 -5496 8858 -5224
rect 8556 -5501 8858 -5496
rect 9300 -5224 9602 -4556
rect 9300 -5496 9310 -5224
rect 9592 -5496 9602 -5224
rect 9300 -5501 9602 -5496
rect 806 -7732 1026 -7727
rect 806 -7932 816 -7732
rect 1016 -7932 1026 -7732
rect 806 -7937 1026 -7932
rect 1530 -7732 1750 -7727
rect 1530 -7932 1540 -7732
rect 1740 -7932 1750 -7732
rect 1530 -7937 1750 -7932
rect 2274 -7732 2494 -7727
rect 2274 -7932 2284 -7732
rect 2484 -7932 2494 -7732
rect 2274 -7937 2494 -7932
rect 3018 -7732 3238 -7727
rect 3018 -7932 3028 -7732
rect 3228 -7932 3238 -7732
rect 3018 -7937 3238 -7932
rect 3762 -7732 3982 -7727
rect 3762 -7932 3772 -7732
rect 3972 -7932 3982 -7732
rect 3762 -7937 3982 -7932
rect 4506 -7732 4726 -7727
rect 4506 -7932 4516 -7732
rect 4716 -7932 4726 -7732
rect 4506 -7937 4726 -7932
rect 5250 -7732 5470 -7727
rect 5250 -7932 5260 -7732
rect 5460 -7932 5470 -7732
rect 5250 -7937 5470 -7932
rect 5994 -7732 6214 -7727
rect 5994 -7932 6004 -7732
rect 6204 -7932 6214 -7732
rect 5994 -7937 6214 -7932
rect 6738 -7732 6958 -7727
rect 6738 -7932 6748 -7732
rect 6948 -7932 6958 -7732
rect 6738 -7937 6958 -7932
rect 7482 -7732 7702 -7727
rect 7482 -7932 7492 -7732
rect 7692 -7932 7702 -7732
rect 7482 -7937 7702 -7932
rect 8226 -7732 8446 -7727
rect 8226 -7932 8236 -7732
rect 8436 -7932 8446 -7732
rect 8226 -7937 8446 -7932
rect 8970 -7732 9190 -7727
rect 8970 -7932 8980 -7732
rect 9180 -7932 9190 -7732
rect 8970 -7937 9190 -7932
rect 9714 -7732 9934 -7727
rect 9714 -7932 9724 -7732
rect 9924 -7932 9934 -7732
rect 9714 -7937 9934 -7932
<< via3 >>
rect -322 1314 -122 1514
rect 422 1314 622 1514
rect 1166 1314 1366 1514
rect 1910 1314 2110 1514
rect 2654 1314 2854 1514
rect 3398 1314 3598 1514
rect 4142 1314 4342 1514
rect 4886 1314 5086 1514
rect 5258 1314 5458 1514
rect 6002 1314 6202 1514
rect 6746 1314 6946 1514
rect 7490 1314 7690 1514
rect 8234 1314 8434 1514
rect 8978 1314 9178 1514
rect 9722 1314 9922 1514
rect 10466 1314 10666 1514
rect 11210 1314 11410 1514
rect 6012 -3088 6294 -2816
rect 5686 -3690 5846 -3528
rect 5686 -4090 5846 -3928
rect 5686 -4490 5846 -4328
rect 816 -7932 1016 -7732
rect 1540 -7932 1740 -7732
rect 2284 -7932 2484 -7732
rect 3028 -7932 3228 -7732
rect 3772 -7932 3972 -7732
rect 4516 -7932 4716 -7732
rect 5260 -7932 5460 -7732
rect 6004 -7932 6204 -7732
rect 6748 -7932 6948 -7732
rect 7492 -7932 7692 -7732
rect 8236 -7932 8436 -7732
rect 8980 -7932 9180 -7732
rect 9724 -7932 9924 -7732
<< mimcap >>
rect 6908 -1696 9708 -1656
rect 6908 -4416 6948 -1696
rect 9668 -4416 9708 -1696
rect 6908 -4456 9708 -4416
<< mimcapcontact >>
rect 6948 -4416 9668 -1696
<< metal4 >>
rect -928 1514 11596 2292
rect -928 1314 -322 1514
rect -122 1314 422 1514
rect 622 1314 1166 1514
rect 1366 1314 1910 1514
rect 2110 1314 2654 1514
rect 2854 1314 3398 1514
rect 3598 1314 4142 1514
rect 4342 1314 4886 1514
rect 5086 1314 5258 1514
rect 5458 1314 6002 1514
rect 6202 1314 6746 1514
rect 6946 1314 7490 1514
rect 7690 1314 8234 1514
rect 8434 1314 8978 1514
rect 9178 1314 9722 1514
rect 9922 1314 10466 1514
rect 10666 1314 11210 1514
rect 11410 1314 11596 1514
rect -928 1288 11596 1314
rect 6947 -1696 9669 -1695
rect 6011 -2816 6295 -2815
rect 6011 -3088 6012 -2816
rect 6294 -2844 6295 -2816
rect 6947 -2844 6948 -1696
rect 6294 -3062 6948 -2844
rect 6294 -3088 6295 -3062
rect 6011 -3089 6295 -3088
rect 5638 -3528 5876 -3490
rect 5638 -3690 5686 -3528
rect 5846 -3690 5876 -3528
rect 5638 -3928 5876 -3690
rect 5638 -4090 5686 -3928
rect 5846 -4090 5876 -3928
rect 5638 -4328 5876 -4090
rect 5638 -4490 5686 -4328
rect 5846 -4490 5876 -4328
rect 6947 -4416 6948 -3062
rect 9668 -4416 9669 -1696
rect 6947 -4417 9669 -4416
rect 5638 -7708 5876 -4490
rect -928 -7732 11596 -7708
rect -928 -7932 816 -7732
rect 1016 -7932 1540 -7732
rect 1740 -7932 2284 -7732
rect 2484 -7932 3028 -7732
rect 3228 -7932 3772 -7732
rect 3972 -7932 4516 -7732
rect 4716 -7932 5260 -7732
rect 5460 -7932 6004 -7732
rect 6204 -7932 6748 -7732
rect 6948 -7932 7492 -7732
rect 7692 -7932 8236 -7732
rect 8436 -7932 8980 -7732
rect 9180 -7932 9724 -7732
rect 9924 -7932 11596 -7732
rect -928 -8712 11596 -7932
<< labels >>
flabel metal4 268 1966 268 1966 0 FreeSans 8000 0 0 0 vdd
port 0 nsew
flabel metal4 -166 -8548 -166 -8548 0 FreeSans 8000 0 0 0 vss
port 4 nsew
flabel metal2 546 -1130 546 -1130 0 FreeSans 8000 0 0 0 vn
port 2 nsew
flabel metal2 582 -5530 582 -5530 0 FreeSans 8000 0 0 0 vp
port 1 nsew
flabel metal3 10132 -3112 10132 -3112 0 FreeSans 8000 0 0 0 vout
port 5 nsew
flabel metal1 -542 -130 -542 -130 0 FreeSans 8000 0 0 0 vbias
port 3 nsew
<< end >>
