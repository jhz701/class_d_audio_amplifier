magic
tech sky130A
magscale 1 2
timestamp 1629189331
<< pwell >>
rect -1869 5189 127 7817
rect 25383 4217 25785 7213
rect 25383 1347 25785 3343
<< psubdiff >>
rect -1833 7747 -1737 7781
rect -5 7747 91 7781
rect -1833 7685 -1799 7747
rect 57 7685 91 7747
rect -1833 5259 -1799 5321
rect 57 5259 91 5321
rect -1833 5225 -1737 5259
rect -5 5225 91 5259
rect 25419 7143 25515 7177
rect 25653 7143 25749 7177
rect 25419 7081 25453 7143
rect 25715 7081 25749 7143
rect 25419 4287 25453 4349
rect 25715 4287 25749 4349
rect 25419 4253 25515 4287
rect 25653 4253 25749 4287
rect 25419 3273 25515 3307
rect 25653 3273 25749 3307
rect 25419 3211 25453 3273
rect 25715 3211 25749 3273
rect 25419 1417 25453 1479
rect 25715 1417 25749 1479
rect 25419 1383 25515 1417
rect 25653 1383 25749 1417
<< psubdiffcont >>
rect -1737 7747 -5 7781
rect -1833 5321 -1799 7685
rect 57 5321 91 7685
rect -1737 5225 -5 5259
rect 25515 7143 25653 7177
rect 25419 4349 25453 7081
rect 25715 4349 25749 7081
rect 25515 4253 25653 4287
rect 25515 3273 25653 3307
rect 25419 1479 25453 3211
rect 25715 1479 25749 3211
rect 25515 1383 25653 1417
<< xpolycontact >>
rect -1703 7581 -1271 7651
rect -471 7581 -39 7651
rect -1703 7263 -1271 7333
rect -471 7263 -39 7333
rect -1703 6945 -1271 7015
rect -471 6945 -39 7015
rect -1703 6627 -1271 6697
rect -471 6627 -39 6697
rect -1703 6309 -1271 6379
rect -471 6309 -39 6379
rect -1703 5991 -1271 6061
rect -471 5991 -39 6061
rect -1703 5673 -1271 5743
rect -471 5673 -39 5743
rect -1703 5355 -1271 5425
rect -471 5355 -39 5425
rect 25549 6615 25619 7047
rect 25549 4383 25619 4815
rect 25549 2745 25619 3177
rect 25549 1513 25619 1945
<< xpolyres >>
rect -1271 7581 -471 7651
rect -1271 7263 -471 7333
rect -1271 6945 -471 7015
rect -1271 6627 -471 6697
rect -1271 6309 -471 6379
rect -1271 5991 -471 6061
rect -1271 5673 -471 5743
rect -1271 5355 -471 5425
rect 25549 4815 25619 6615
rect 25549 1945 25619 2745
<< locali >>
rect -1833 7747 -1737 7781
rect -5 7747 91 7781
rect -1833 7685 -1799 7747
rect 57 7685 91 7747
rect 25419 7143 25515 7177
rect 25653 7143 25749 7177
rect 25419 7081 25453 7143
rect -1833 5259 -1799 5321
rect 57 5259 91 5321
rect -1833 5225 -1737 5259
rect -5 5225 91 5259
rect 25715 7081 25749 7143
rect 25419 4287 25453 4349
rect 25715 4287 25749 4349
rect 25419 4253 25515 4287
rect 25653 4253 25749 4287
rect 25419 3273 25515 3307
rect 25653 3273 25749 3307
rect 25419 3211 25453 3273
rect 25715 3211 25749 3273
rect 25419 1417 25453 1479
rect 25715 1417 25749 1479
rect 25419 1383 25515 1417
rect 25653 1383 25749 1417
<< viali >>
rect -1685 7597 -1288 7635
rect -454 7597 -57 7635
rect -1685 7279 -1288 7317
rect -454 7279 -57 7317
rect -1685 6961 -1288 6999
rect 42 7010 57 7068
rect 57 7010 91 7068
rect 91 7010 106 7068
rect -454 6961 -57 6999
rect -1685 6643 -1288 6681
rect -454 6643 -57 6681
rect 42 6610 57 6668
rect 57 6610 91 6668
rect 91 6610 106 6668
rect -1685 6325 -1288 6363
rect -454 6325 -57 6363
rect 42 6210 57 6268
rect 57 6210 91 6268
rect 91 6210 106 6268
rect -1685 6007 -1288 6045
rect -454 6007 -57 6045
rect 42 5810 57 5868
rect 57 5810 91 5868
rect 91 5810 106 5868
rect -1685 5689 -1288 5727
rect -454 5689 -57 5727
rect -1685 5371 -1288 5409
rect -454 5371 -57 5409
rect 25565 6632 25603 7029
rect 25700 5970 25715 6028
rect 25715 5970 25749 6028
rect 25749 5970 25764 6028
rect 25700 5570 25715 5628
rect 25715 5570 25749 5628
rect 25749 5570 25764 5628
rect 25700 5170 25715 5228
rect 25715 5170 25749 5228
rect 25749 5170 25764 5228
rect 25565 4401 25603 4798
rect 25700 4770 25715 4828
rect 25715 4770 25749 4828
rect 25749 4770 25764 4828
rect 25565 2762 25603 3159
rect 25700 2970 25715 3028
rect 25715 2970 25749 3028
rect 25749 2970 25764 3028
rect 25700 2570 25715 2628
rect 25715 2570 25749 2628
rect 25749 2570 25764 2628
rect 25700 2170 25715 2228
rect 25715 2170 25749 2228
rect 25749 2170 25764 2228
rect 25565 1531 25603 1928
rect 25700 1770 25715 1828
rect 25715 1770 25749 1828
rect 25749 1770 25764 1828
<< metal1 >>
rect -1410 11818 -1400 12532
rect -652 11818 -642 12532
rect -1134 11544 -906 11818
rect -1134 11316 -48 11544
rect -276 7654 -48 11316
rect 360 9168 406 9264
rect 13884 9192 13922 9282
rect 344 7654 354 7816
rect -1704 7635 -1270 7652
rect -276 7641 354 7654
rect -1704 7597 -1685 7635
rect -1288 7597 -1270 7635
rect -1704 7317 -1270 7597
rect -466 7635 354 7641
rect -466 7597 -454 7635
rect -57 7597 354 7635
rect -466 7591 354 7597
rect -276 7584 354 7591
rect -262 7582 354 7584
rect 344 7416 354 7582
rect 754 7416 764 7816
rect -1704 7279 -1685 7317
rect -1288 7279 -1270 7317
rect -1704 7262 -1270 7279
rect -472 7317 -38 7334
rect -472 7279 -454 7317
rect -57 7279 -38 7317
rect -1704 6999 -1270 7016
rect -1704 6961 -1685 6999
rect -1288 6961 -1270 6999
rect -1704 6681 -1270 6961
rect -472 6999 -38 7279
rect 380 7074 390 7140
rect 30 7068 390 7074
rect 30 7010 42 7068
rect 106 7010 390 7068
rect 30 7004 390 7010
rect -472 6961 -454 6999
rect -57 6961 -38 6999
rect 380 6970 390 7004
rect 558 6970 568 7140
rect -472 6944 -38 6961
rect -1704 6643 -1685 6681
rect -1288 6643 -1270 6681
rect -1704 6626 -1270 6643
rect -472 6681 -38 6698
rect -472 6643 -454 6681
rect -57 6643 -38 6681
rect 380 6674 390 6740
rect -1704 6363 -1270 6380
rect -1704 6325 -1685 6363
rect -1288 6325 -1270 6363
rect -1704 6045 -1270 6325
rect -472 6363 -38 6643
rect 30 6668 390 6674
rect 30 6610 42 6668
rect 106 6610 390 6668
rect 30 6604 390 6610
rect 380 6570 390 6604
rect 558 6570 568 6740
rect 24362 6718 24372 7106
rect 24754 7048 24764 7106
rect 24754 7029 25620 7048
rect 24754 6850 25565 7029
rect 24754 6718 24764 6850
rect 25559 6632 25565 6850
rect 25603 6850 25620 7029
rect 25603 6632 25609 6850
rect 25559 6620 25609 6632
rect -472 6325 -454 6363
rect -57 6325 -38 6363
rect -472 6308 -38 6325
rect 380 6274 390 6340
rect 30 6268 390 6274
rect 30 6210 42 6268
rect 106 6210 390 6268
rect 30 6204 390 6210
rect 380 6170 390 6204
rect 558 6170 568 6340
rect -1704 6007 -1685 6045
rect -1288 6007 -1270 6045
rect -1704 5990 -1270 6007
rect -472 6045 -38 6062
rect -472 6007 -454 6045
rect -57 6007 -38 6045
rect 25948 6034 25958 6100
rect -1704 5727 -1270 5744
rect -1704 5689 -1685 5727
rect -1288 5689 -1270 5727
rect -1704 5409 -1270 5689
rect -472 5727 -38 6007
rect 25688 6028 25958 6034
rect 25688 5970 25700 6028
rect 25764 5970 25958 6028
rect 25688 5964 25958 5970
rect 380 5874 390 5940
rect 30 5868 390 5874
rect 30 5810 42 5868
rect 106 5810 390 5868
rect 30 5804 390 5810
rect 380 5770 390 5804
rect 558 5770 568 5940
rect 25948 5930 25958 5964
rect 26126 5930 26136 6100
rect -472 5689 -454 5727
rect -57 5689 -38 5727
rect -472 5672 -38 5689
rect 25948 5634 25958 5700
rect 25688 5628 25958 5634
rect 25688 5570 25700 5628
rect 25764 5570 25958 5628
rect 25688 5564 25958 5570
rect 25948 5530 25958 5564
rect 26126 5530 26136 5700
rect -1704 5371 -1685 5409
rect -1288 5371 -1270 5409
rect -1704 5354 -1270 5371
rect -466 5409 -45 5415
rect -466 5371 -454 5409
rect -57 5371 -45 5409
rect -466 5365 -45 5371
rect -420 -286 -100 5365
rect 25948 5234 25958 5300
rect 25688 5228 25958 5234
rect 25688 5170 25700 5228
rect 25764 5170 25958 5228
rect 25688 5164 25958 5170
rect 25948 5130 25958 5164
rect 26126 5130 26136 5300
rect 25948 4834 25958 4900
rect 25688 4828 25958 4834
rect 25548 4798 25620 4816
rect 25548 4401 25565 4798
rect 25603 4401 25620 4798
rect 25688 4770 25700 4828
rect 25764 4770 25958 4828
rect 25688 4764 25958 4770
rect 25948 4730 25958 4764
rect 26126 4730 26136 4900
rect 25548 3928 25620 4401
rect 25402 3570 25412 3928
rect 25748 3570 25758 3928
rect 25548 3159 25620 3570
rect 25548 2762 25565 3159
rect 25603 2762 25620 3159
rect 25948 3034 25958 3100
rect 25688 3028 25958 3034
rect 25688 2970 25700 3028
rect 25764 2970 25958 3028
rect 25688 2964 25958 2970
rect 25948 2930 25958 2964
rect 26126 2930 26136 3100
rect 25548 2744 25620 2762
rect 25948 2634 25958 2700
rect 25688 2628 25958 2634
rect 25688 2570 25700 2628
rect 25764 2570 25958 2628
rect 25688 2564 25958 2570
rect 25948 2530 25958 2564
rect 26126 2530 26136 2700
rect 25948 2234 25958 2300
rect 25688 2228 25958 2234
rect 25688 2170 25700 2228
rect 25764 2170 25958 2228
rect 25688 2164 25958 2170
rect 25948 2130 25958 2164
rect 26126 2130 26136 2300
rect 25548 1928 25620 1946
rect 25548 1531 25565 1928
rect 25603 1531 25620 1928
rect 25948 1834 25958 1900
rect 25688 1828 25958 1834
rect 25688 1770 25700 1828
rect 25764 1770 25958 1828
rect 25688 1764 25958 1770
rect 25948 1730 25958 1764
rect 26126 1730 26136 1900
rect 25548 356 25620 1531
rect 25400 -2 25410 356
rect 25746 -2 25756 356
rect -474 -686 -464 -286
rect -64 -686 -54 -286
<< via1 >>
rect -1400 11818 -652 12532
rect 354 7416 754 7816
rect 390 6970 558 7140
rect 390 6570 558 6740
rect 24372 6718 24754 7106
rect 390 6170 558 6340
rect 390 5770 558 5940
rect 25958 5930 26126 6100
rect 25958 5530 26126 5700
rect 25958 5130 26126 5300
rect 25958 4730 26126 4900
rect 25412 3570 25748 3928
rect 25958 2930 26126 3100
rect 25958 2530 26126 2700
rect 25958 2130 26126 2300
rect 25958 1730 26126 1900
rect 25410 -2 25746 356
rect -464 -686 -64 -286
<< metal2 >>
rect -1400 12532 -652 12542
rect -1400 11808 -652 11818
rect 354 7816 754 7826
rect 754 7562 1556 7660
rect 14382 7562 15028 7660
rect 354 7406 754 7416
rect 390 7140 558 7150
rect 390 6960 558 6970
rect 390 6740 558 6750
rect 390 6560 558 6570
rect 14382 6556 14524 7562
rect 24372 7106 24754 7116
rect 24372 6708 24754 6718
rect 5042 6430 14524 6556
rect 390 6340 558 6350
rect 390 6160 558 6170
rect 390 5940 558 5950
rect 390 5760 558 5770
rect 5042 3798 5176 6430
rect 25958 6100 26126 6110
rect 25958 5920 26126 5930
rect 25958 5700 26126 5710
rect 25958 5520 26126 5530
rect 25958 5300 26126 5310
rect 25958 5120 26126 5130
rect 25958 4900 26126 4910
rect 25958 4720 26126 4730
rect 25412 3928 25748 3938
rect 4854 3694 5176 3798
rect 4854 3264 4950 3694
rect 18312 3652 25412 3822
rect 18312 3264 18476 3652
rect 25412 3560 25748 3570
rect 1382 3160 1548 3258
rect 3754 3160 4956 3264
rect 17274 3160 18476 3264
rect 25958 3100 26126 3110
rect 25958 2920 26126 2930
rect 25958 2700 26126 2710
rect 25958 2520 26126 2530
rect 25958 2300 26126 2310
rect 25958 2120 26126 2130
rect 25958 1900 26126 1910
rect 25958 1720 26126 1730
rect 11872 734 12626 744
rect 25410 356 25746 366
rect 12626 22 25410 332
rect 11872 12 12626 22
rect 25410 -12 25746 -2
rect 24180 -132 24934 -122
rect -464 -286 -64 -276
rect -64 -686 24180 -376
rect -464 -696 -64 -686
rect 24180 -854 24934 -844
<< via2 >>
rect -1400 11818 -652 12532
rect 390 6970 558 7140
rect 390 6570 558 6740
rect 24372 6718 24754 7106
rect 390 6170 558 6340
rect 390 5770 558 5940
rect 25958 5930 26126 6100
rect 25958 5530 26126 5700
rect 25958 5130 26126 5300
rect 25958 4730 26126 4900
rect 25958 2930 26126 3100
rect 25958 2530 26126 2700
rect 25958 2130 26126 2300
rect 25958 1730 26126 1900
rect 11872 22 12626 734
rect 24180 -844 24934 -132
<< metal3 >>
rect -1410 12532 -642 12537
rect -1410 11818 -1400 12532
rect -652 11818 -642 12532
rect -1410 11813 -642 11818
rect -336 11488 26052 14688
rect 380 7140 568 7145
rect 380 6970 390 7140
rect 558 6970 568 7140
rect 380 6965 568 6970
rect 380 6740 568 6745
rect 380 6570 390 6740
rect 558 6570 568 6740
rect 380 6565 568 6570
rect 380 6340 568 6345
rect 380 6170 390 6340
rect 558 6170 568 6340
rect 380 6165 568 6170
rect 380 5940 568 5945
rect 380 5770 390 5940
rect 558 5770 568 5940
rect 380 5765 568 5770
rect 12760 5572 13160 11488
rect 24362 7106 24764 7111
rect 24362 6718 24372 7106
rect 24754 6718 24764 7106
rect 24362 6713 24764 6718
rect 11872 4822 13160 5572
rect 24374 6012 24748 6713
rect 25948 6100 26136 6105
rect 24374 5272 24812 6012
rect 25948 5930 25958 6100
rect 26126 5930 26136 6100
rect 25948 5925 26136 5930
rect 25948 5700 26136 5705
rect 25948 5530 25958 5700
rect 26126 5530 26136 5700
rect 25948 5525 26136 5530
rect 11872 739 12520 4822
rect 11862 734 12636 739
rect 11862 22 11872 734
rect 12626 22 12636 734
rect 11862 17 12636 22
rect 11872 -1600 12520 17
rect 24438 -127 24812 5272
rect 25948 5300 26136 5305
rect 25948 5130 25958 5300
rect 26126 5130 26136 5300
rect 25948 5125 26136 5130
rect 25948 4900 26136 4905
rect 25948 4730 25958 4900
rect 26126 4730 26136 4900
rect 25948 4725 26136 4730
rect 25948 3100 26136 3105
rect 25948 2930 25958 3100
rect 26126 2930 26136 3100
rect 25948 2925 26136 2930
rect 25948 2700 26136 2705
rect 25948 2530 25958 2700
rect 26126 2530 26136 2700
rect 25948 2525 26136 2530
rect 25948 2300 26136 2305
rect 25948 2130 25958 2300
rect 26126 2130 26136 2300
rect 25948 2125 26136 2130
rect 25948 1900 26136 1905
rect 25948 1730 25958 1900
rect 26126 1730 26136 1900
rect 25948 1725 26136 1730
rect 24170 -132 24944 -127
rect 24170 -844 24180 -132
rect 24934 -844 24944 -132
rect 24170 -849 24944 -844
<< via3 >>
rect -1400 11818 -652 12532
rect 390 6970 558 7140
rect 390 6570 558 6740
rect 390 6170 558 6340
rect 390 5770 558 5940
rect 25958 5930 26126 6100
rect 25958 5530 26126 5700
rect 25958 5130 26126 5300
rect 25958 4730 26126 4900
rect 25958 2930 26126 3100
rect 25958 2530 26126 2700
rect 25958 2130 26126 2300
rect 25958 1730 26126 1900
<< mimcap >>
rect -235 14548 2765 14588
rect -235 11628 -195 14548
rect 2725 11628 2765 14548
rect -235 11588 2765 11628
rect 3084 14548 6084 14588
rect 3084 11628 3124 14548
rect 6044 11628 6084 14548
rect 3084 11588 6084 11628
rect 6403 14548 9403 14588
rect 6403 11628 6443 14548
rect 9363 11628 9403 14548
rect 6403 11588 9403 11628
rect 9722 14548 12722 14588
rect 9722 11628 9762 14548
rect 12682 11628 12722 14548
rect 9722 11588 12722 11628
rect 13041 14548 16041 14588
rect 13041 11628 13081 14548
rect 16001 11628 16041 14548
rect 13041 11588 16041 11628
rect 16360 14548 19360 14588
rect 16360 11628 16400 14548
rect 19320 11628 19360 14548
rect 16360 11588 19360 11628
rect 19679 14548 22679 14588
rect 19679 11628 19719 14548
rect 22639 11628 22679 14548
rect 19679 11588 22679 11628
rect 22998 14548 25998 14588
rect 22998 11628 23038 14548
rect 25958 11628 25998 14548
rect 22998 11588 25998 11628
<< mimcapcontact >>
rect -195 11628 2725 14548
rect 3124 11628 6044 14548
rect 6443 11628 9363 14548
rect 9762 11628 12682 14548
rect 13081 11628 16001 14548
rect 16400 11628 19320 14548
rect 19719 11628 22639 14548
rect 23038 11628 25958 14548
<< metal4 >>
rect -336 14548 26052 14688
rect -1401 12532 -651 12533
rect -1401 11818 -1400 12532
rect -652 12456 -651 12532
rect -336 12456 -195 14548
rect -652 11860 -195 12456
rect -652 11818 -651 11860
rect -1401 11817 -651 11818
rect -336 11628 -195 11860
rect 2725 11628 3124 14548
rect 6044 11628 6443 14548
rect 9363 11628 9762 14548
rect 12682 11628 13081 14548
rect 16001 11628 16400 14548
rect 19320 11628 19719 14548
rect 22639 11628 23038 14548
rect 25958 11628 26052 14548
rect -336 11488 26052 11628
rect -8 10010 26040 11014
rect 322 7188 584 7192
rect 322 7140 602 7188
rect 322 6970 390 7140
rect 558 6970 602 7140
rect 322 6740 602 6970
rect 322 6570 390 6740
rect 558 6570 602 6740
rect 322 6340 602 6570
rect 322 6170 390 6340
rect 558 6170 602 6340
rect 322 5940 602 6170
rect 322 5770 390 5940
rect 558 5770 602 5940
rect 322 1014 602 5770
rect 25922 6100 26228 7140
rect 25922 5930 25958 6100
rect 26126 5930 26228 6100
rect 25922 5700 26228 5930
rect 25922 5530 25958 5700
rect 26126 5530 26228 5700
rect 25922 5300 26228 5530
rect 25922 5130 25958 5300
rect 26126 5130 26228 5300
rect 25922 4900 26228 5130
rect 25922 4730 25958 4900
rect 26126 4730 26228 4900
rect 25922 3100 26228 4730
rect 25922 2930 25958 3100
rect 26126 2930 26228 3100
rect 25922 2700 26228 2930
rect 25922 2530 25958 2700
rect 26126 2530 26228 2700
rect 25922 2300 26228 2530
rect 25922 2130 25958 2300
rect 26126 2130 26228 2300
rect 25922 1900 26228 2130
rect 25922 1730 25958 1900
rect 26126 1730 26228 1900
rect 25922 1014 26228 1730
rect -8 834 26228 1014
rect -8 10 26040 834
use OTA_revised  OTA_revised_0 ~/magic/class_d_audio_amplifier/OTA
timestamp 1629189150
transform 1 0 14444 0 1 8722
box -928 -8712 11596 2292
use OTA_tri_revised  OTA_tri_revised_0 ~/magic/class_d_audio_amplifier/OTA
timestamp 1629189117
transform 1 0 -28408 0 1 -2358
box 28400 2368 40924 13372
<< labels >>
flabel metal2 1446 3184 1446 3184 0 FreeSans 8000 0 0 0 vref
port 3 nsew
flabel metal1 376 9212 376 9212 0 FreeSans 8000 0 0 0 vbias1
port 1 nsew
flabel metal1 13896 9236 13896 9236 0 FreeSans 8000 0 0 0 vbias2
port 2 nsew
flabel metal3 12326 -1286 12326 -1286 0 FreeSans 8000 0 0 0 vt
port 6 nsew
flabel metal4 3374 10634 3374 10634 0 FreeSans 8000 0 0 0 vdd
port 0 nsew
flabel metal4 2594 294 2594 294 0 FreeSans 8000 0 0 0 vss
port 4 nsew
flabel metal3 24566 6226 24566 6226 0 FreeSans 8000 0 0 0 vsquare
port 5 nsew
<< end >>
