magic
tech sky130A
magscale 1 2
timestamp 1630379054
<< nwell >>
rect 126416 20570 135414 23100
rect 121544 19144 135414 20570
rect 118942 17718 135414 19144
rect 116132 15836 116646 16348
rect 115706 15552 116646 15554
rect 115704 15042 116646 15552
rect 115704 14990 116026 15042
rect 118942 12246 125984 13672
rect 121544 10820 125984 12246
<< pwell >>
rect 126446 25334 135770 28416
rect 121772 20684 125972 22212
rect 118988 19238 120962 20412
rect 116154 16502 116632 16926
rect 115678 14624 116022 14854
rect 116154 14464 116632 14888
rect 118988 10978 120962 12152
rect 121772 7778 125972 9306
<< nmos >>
rect 126932 26980 126962 27980
rect 127142 26980 127172 27980
rect 127352 26980 127382 27980
rect 127562 26980 127592 27980
rect 127772 26980 127802 27980
rect 127982 26980 128012 27980
rect 128192 26980 128222 27980
rect 128402 26980 128432 27980
rect 128612 26980 128642 27980
rect 128822 26980 128852 27980
rect 129032 26980 129062 27980
rect 129242 26980 129272 27980
rect 129452 26980 129482 27980
rect 129662 26980 129692 27980
rect 129872 26980 129902 27980
rect 130082 26980 130112 27980
rect 130292 26980 130322 27980
rect 130502 26980 130532 27980
rect 130712 26980 130742 27980
rect 130922 26980 130952 27980
rect 131132 26980 131162 27980
rect 131342 26980 131372 27980
rect 131552 26980 131582 27980
rect 131762 26980 131792 27980
rect 131972 26980 132002 27980
rect 132182 26980 132212 27980
rect 132392 26980 132422 27980
rect 132602 26980 132632 27980
rect 132812 26980 132842 27980
rect 133022 26980 133052 27980
rect 133232 26980 133262 27980
rect 133442 26980 133472 27980
rect 133652 26980 133682 27980
rect 133862 26980 133892 27980
rect 134072 26980 134102 27980
rect 134282 26980 134312 27980
rect 134492 26980 134522 27980
rect 134702 26980 134732 27980
rect 134912 26980 134942 27980
rect 135122 26980 135152 27980
rect 126932 25762 126962 26762
rect 127142 25762 127172 26762
rect 127352 25762 127382 26762
rect 127562 25762 127592 26762
rect 127772 25762 127802 26762
rect 127982 25762 128012 26762
rect 128192 25762 128222 26762
rect 128402 25762 128432 26762
rect 128612 25762 128642 26762
rect 128822 25762 128852 26762
rect 129032 25762 129062 26762
rect 129242 25762 129272 26762
rect 129452 25762 129482 26762
rect 129662 25762 129692 26762
rect 129872 25762 129902 26762
rect 130082 25762 130112 26762
rect 130292 25762 130322 26762
rect 130502 25762 130532 26762
rect 130712 25762 130742 26762
rect 130922 25762 130952 26762
rect 131132 25762 131162 26762
rect 131342 25762 131372 26762
rect 131552 25762 131582 26762
rect 131762 25762 131792 26762
rect 131972 25762 132002 26762
rect 132182 25762 132212 26762
rect 132392 25762 132422 26762
rect 132602 25762 132632 26762
rect 132812 25762 132842 26762
rect 133022 25762 133052 26762
rect 133232 25762 133262 26762
rect 133442 25762 133472 26762
rect 133652 25762 133682 26762
rect 133862 25762 133892 26762
rect 134072 25762 134102 26762
rect 134282 25762 134312 26762
rect 134492 25762 134522 26762
rect 134702 25762 134732 26762
rect 134912 25762 134942 26762
rect 135122 25762 135152 26762
rect 122082 20896 122112 21896
rect 122292 20896 122322 21896
rect 122502 20896 122532 21896
rect 122712 20896 122742 21896
rect 122922 20896 122952 21896
rect 123132 20896 123162 21896
rect 123342 20896 123372 21896
rect 123552 20896 123582 21896
rect 123762 20896 123792 21896
rect 123972 20896 124002 21896
rect 124182 20896 124212 21896
rect 124392 20896 124422 21896
rect 124602 20896 124632 21896
rect 124812 20896 124842 21896
rect 125022 20896 125052 21896
rect 125232 20896 125262 21896
rect 125442 20896 125472 21896
rect 125652 20896 125682 21896
rect 119170 19272 119200 20272
rect 120118 19272 120148 20272
rect 120328 19272 120358 20272
rect 120538 19272 120568 20272
rect 120748 19272 120778 20272
rect 116428 16518 116458 16918
rect 116522 16518 116552 16918
rect 115902 14634 115932 14834
rect 116428 14472 116458 14872
rect 116522 14472 116552 14872
rect 119170 11118 119200 12118
rect 120118 11118 120148 12118
rect 120328 11118 120358 12118
rect 120538 11118 120568 12118
rect 120748 11118 120778 12118
rect 122082 8094 122112 9094
rect 122292 8094 122322 9094
rect 122502 8094 122532 9094
rect 122712 8094 122742 9094
rect 122922 8094 122952 9094
rect 123132 8094 123162 9094
rect 123342 8094 123372 9094
rect 123552 8094 123582 9094
rect 123762 8094 123792 9094
rect 123972 8094 124002 9094
rect 124182 8094 124212 9094
rect 124392 8094 124422 9094
rect 124602 8094 124632 9094
rect 124812 8094 124842 9094
rect 125022 8094 125052 9094
rect 125232 8094 125262 9094
rect 125442 8094 125472 9094
rect 125652 8094 125682 9094
<< pmos >>
rect 119170 18044 119200 19044
rect 119266 18044 119296 19044
rect 119908 18044 119938 19044
rect 120118 18044 120148 19044
rect 120328 18044 120358 19044
rect 120538 18044 120568 19044
rect 120748 18044 120778 19044
rect 120958 18044 120988 19044
rect 121168 18044 121198 19044
rect 121378 18044 121408 19044
rect 122082 19280 122112 20280
rect 122292 19280 122322 20280
rect 122502 19280 122532 20280
rect 122712 19280 122742 20280
rect 122922 19280 122952 20280
rect 123132 19280 123162 20280
rect 123342 19280 123372 20280
rect 123552 19280 123582 20280
rect 123762 19280 123792 20280
rect 123972 19280 124002 20280
rect 124182 19280 124212 20280
rect 124392 19280 124422 20280
rect 124602 19280 124632 20280
rect 124812 19280 124842 20280
rect 125022 19280 125052 20280
rect 125232 19280 125262 20280
rect 125442 19280 125472 20280
rect 125652 19280 125682 20280
rect 122082 18044 122112 19044
rect 122292 18044 122322 19044
rect 122502 18044 122532 19044
rect 122712 18044 122742 19044
rect 122922 18044 122952 19044
rect 123132 18044 123162 19044
rect 123342 18044 123372 19044
rect 123552 18044 123582 19044
rect 123762 18044 123792 19044
rect 123972 18044 124002 19044
rect 124182 18044 124212 19044
rect 124392 18044 124422 19044
rect 124602 18044 124632 19044
rect 124812 18044 124842 19044
rect 125022 18044 125052 19044
rect 125232 18044 125262 19044
rect 125442 18044 125472 19044
rect 125652 18044 125682 19044
rect 126932 21752 126962 22752
rect 127142 21752 127172 22752
rect 127352 21752 127382 22752
rect 127562 21752 127592 22752
rect 127772 21752 127802 22752
rect 127982 21752 128012 22752
rect 128192 21752 128222 22752
rect 128402 21752 128432 22752
rect 128612 21752 128642 22752
rect 128822 21752 128852 22752
rect 129032 21752 129062 22752
rect 129242 21752 129272 22752
rect 129452 21752 129482 22752
rect 129662 21752 129692 22752
rect 129872 21752 129902 22752
rect 130082 21752 130112 22752
rect 130292 21752 130322 22752
rect 130502 21752 130532 22752
rect 130712 21752 130742 22752
rect 130922 21752 130952 22752
rect 131132 21752 131162 22752
rect 131342 21752 131372 22752
rect 131552 21752 131582 22752
rect 131762 21752 131792 22752
rect 131972 21752 132002 22752
rect 132182 21752 132212 22752
rect 132392 21752 132422 22752
rect 132602 21752 132632 22752
rect 132812 21752 132842 22752
rect 133022 21752 133052 22752
rect 133232 21752 133262 22752
rect 133442 21752 133472 22752
rect 133652 21752 133682 22752
rect 133862 21752 133892 22752
rect 134072 21752 134102 22752
rect 134282 21752 134312 22752
rect 134492 21752 134522 22752
rect 134702 21752 134732 22752
rect 134912 21752 134942 22752
rect 135122 21752 135152 22752
rect 126932 20516 126962 21516
rect 127142 20516 127172 21516
rect 127352 20516 127382 21516
rect 127562 20516 127592 21516
rect 127772 20516 127802 21516
rect 127982 20516 128012 21516
rect 128192 20516 128222 21516
rect 128402 20516 128432 21516
rect 128612 20516 128642 21516
rect 128822 20516 128852 21516
rect 129032 20516 129062 21516
rect 129242 20516 129272 21516
rect 129452 20516 129482 21516
rect 129662 20516 129692 21516
rect 129872 20516 129902 21516
rect 130082 20516 130112 21516
rect 130292 20516 130322 21516
rect 130502 20516 130532 21516
rect 130712 20516 130742 21516
rect 130922 20516 130952 21516
rect 131132 20516 131162 21516
rect 131342 20516 131372 21516
rect 131552 20516 131582 21516
rect 131762 20516 131792 21516
rect 131972 20516 132002 21516
rect 132182 20516 132212 21516
rect 132392 20516 132422 21516
rect 132602 20516 132632 21516
rect 132812 20516 132842 21516
rect 133022 20516 133052 21516
rect 133232 20516 133262 21516
rect 133442 20516 133472 21516
rect 133652 20516 133682 21516
rect 133862 20516 133892 21516
rect 134072 20516 134102 21516
rect 134282 20516 134312 21516
rect 134492 20516 134522 21516
rect 134702 20516 134732 21516
rect 134912 20516 134942 21516
rect 135122 20516 135152 21516
rect 126932 19280 126962 20280
rect 127142 19280 127172 20280
rect 127352 19280 127382 20280
rect 127562 19280 127592 20280
rect 127772 19280 127802 20280
rect 127982 19280 128012 20280
rect 128192 19280 128222 20280
rect 128402 19280 128432 20280
rect 128612 19280 128642 20280
rect 128822 19280 128852 20280
rect 129032 19280 129062 20280
rect 129242 19280 129272 20280
rect 129452 19280 129482 20280
rect 129662 19280 129692 20280
rect 129872 19280 129902 20280
rect 130082 19280 130112 20280
rect 130292 19280 130322 20280
rect 130502 19280 130532 20280
rect 130712 19280 130742 20280
rect 130922 19280 130952 20280
rect 131132 19280 131162 20280
rect 131342 19280 131372 20280
rect 131552 19280 131582 20280
rect 131762 19280 131792 20280
rect 131972 19280 132002 20280
rect 132182 19280 132212 20280
rect 132392 19280 132422 20280
rect 132602 19280 132632 20280
rect 132812 19280 132842 20280
rect 133022 19280 133052 20280
rect 133232 19280 133262 20280
rect 133442 19280 133472 20280
rect 133652 19280 133682 20280
rect 133862 19280 133892 20280
rect 134072 19280 134102 20280
rect 134282 19280 134312 20280
rect 134492 19280 134522 20280
rect 134702 19280 134732 20280
rect 134912 19280 134942 20280
rect 135122 19280 135152 20280
rect 126932 18044 126962 19044
rect 127142 18044 127172 19044
rect 127352 18044 127382 19044
rect 127562 18044 127592 19044
rect 127772 18044 127802 19044
rect 127982 18044 128012 19044
rect 128192 18044 128222 19044
rect 128402 18044 128432 19044
rect 128612 18044 128642 19044
rect 128822 18044 128852 19044
rect 129032 18044 129062 19044
rect 129242 18044 129272 19044
rect 129452 18044 129482 19044
rect 129662 18044 129692 19044
rect 129872 18044 129902 19044
rect 130082 18044 130112 19044
rect 130292 18044 130322 19044
rect 130502 18044 130532 19044
rect 130712 18044 130742 19044
rect 130922 18044 130952 19044
rect 131132 18044 131162 19044
rect 131342 18044 131372 19044
rect 131552 18044 131582 19044
rect 131762 18044 131792 19044
rect 131972 18044 132002 19044
rect 132182 18044 132212 19044
rect 132392 18044 132422 19044
rect 132602 18044 132632 19044
rect 132812 18044 132842 19044
rect 133022 18044 133052 19044
rect 133232 18044 133262 19044
rect 133442 18044 133472 19044
rect 133652 18044 133682 19044
rect 133862 18044 133892 19044
rect 134072 18044 134102 19044
rect 134282 18044 134312 19044
rect 134492 18044 134522 19044
rect 134702 18044 134732 19044
rect 134912 18044 134942 19044
rect 135122 18044 135152 19044
rect 116428 15898 116458 16298
rect 116522 15898 116552 16298
rect 115902 15090 115932 15490
rect 116428 15092 116458 15492
rect 116522 15092 116552 15492
rect 119170 12346 119200 13346
rect 119266 12346 119296 13346
rect 119908 12346 119938 13346
rect 120118 12346 120148 13346
rect 120328 12346 120358 13346
rect 120538 12346 120568 13346
rect 120748 12346 120778 13346
rect 120958 12346 120988 13346
rect 121168 12346 121198 13346
rect 121378 12346 121408 13346
rect 122082 12346 122112 13346
rect 122292 12346 122322 13346
rect 122502 12346 122532 13346
rect 122712 12346 122742 13346
rect 122922 12346 122952 13346
rect 123132 12346 123162 13346
rect 123342 12346 123372 13346
rect 123552 12346 123582 13346
rect 123762 12346 123792 13346
rect 123972 12346 124002 13346
rect 124182 12346 124212 13346
rect 124392 12346 124422 13346
rect 124602 12346 124632 13346
rect 124812 12346 124842 13346
rect 125022 12346 125052 13346
rect 125232 12346 125262 13346
rect 125442 12346 125472 13346
rect 125652 12346 125682 13346
rect 122082 11110 122112 12110
rect 122292 11110 122322 12110
rect 122502 11110 122532 12110
rect 122712 11110 122742 12110
rect 122922 11110 122952 12110
rect 123132 11110 123162 12110
rect 123342 11110 123372 12110
rect 123552 11110 123582 12110
rect 123762 11110 123792 12110
rect 123972 11110 124002 12110
rect 124182 11110 124212 12110
rect 124392 11110 124422 12110
rect 124602 11110 124632 12110
rect 124812 11110 124842 12110
rect 125022 11110 125052 12110
rect 125232 11110 125262 12110
rect 125442 11110 125472 12110
rect 125652 11110 125682 12110
<< ndiff >>
rect 126870 27968 126932 27980
rect 126870 26992 126882 27968
rect 126916 26992 126932 27968
rect 126870 26980 126932 26992
rect 126962 27968 127024 27980
rect 126962 26992 126978 27968
rect 127012 26992 127024 27968
rect 126962 26980 127024 26992
rect 127080 27968 127142 27980
rect 127080 26992 127092 27968
rect 127126 26992 127142 27968
rect 127080 26980 127142 26992
rect 127172 27968 127234 27980
rect 127172 26992 127188 27968
rect 127222 26992 127234 27968
rect 127172 26980 127234 26992
rect 127290 27968 127352 27980
rect 127290 26992 127302 27968
rect 127336 26992 127352 27968
rect 127290 26980 127352 26992
rect 127382 27968 127444 27980
rect 127382 26992 127398 27968
rect 127432 26992 127444 27968
rect 127382 26980 127444 26992
rect 127500 27968 127562 27980
rect 127500 26992 127512 27968
rect 127546 26992 127562 27968
rect 127500 26980 127562 26992
rect 127592 27968 127654 27980
rect 127592 26992 127608 27968
rect 127642 26992 127654 27968
rect 127592 26980 127654 26992
rect 127710 27968 127772 27980
rect 127710 26992 127722 27968
rect 127756 26992 127772 27968
rect 127710 26980 127772 26992
rect 127802 27968 127864 27980
rect 127802 26992 127818 27968
rect 127852 26992 127864 27968
rect 127802 26980 127864 26992
rect 127920 27968 127982 27980
rect 127920 26992 127932 27968
rect 127966 26992 127982 27968
rect 127920 26980 127982 26992
rect 128012 27968 128074 27980
rect 128012 26992 128028 27968
rect 128062 26992 128074 27968
rect 128012 26980 128074 26992
rect 128130 27968 128192 27980
rect 128130 26992 128142 27968
rect 128176 26992 128192 27968
rect 128130 26980 128192 26992
rect 128222 27968 128284 27980
rect 128222 26992 128238 27968
rect 128272 26992 128284 27968
rect 128222 26980 128284 26992
rect 128340 27968 128402 27980
rect 128340 26992 128352 27968
rect 128386 26992 128402 27968
rect 128340 26980 128402 26992
rect 128432 27968 128494 27980
rect 128432 26992 128448 27968
rect 128482 26992 128494 27968
rect 128432 26980 128494 26992
rect 128550 27968 128612 27980
rect 128550 26992 128562 27968
rect 128596 26992 128612 27968
rect 128550 26980 128612 26992
rect 128642 27968 128704 27980
rect 128642 26992 128658 27968
rect 128692 26992 128704 27968
rect 128642 26980 128704 26992
rect 128760 27968 128822 27980
rect 128760 26992 128772 27968
rect 128806 26992 128822 27968
rect 128760 26980 128822 26992
rect 128852 27968 128914 27980
rect 128852 26992 128868 27968
rect 128902 26992 128914 27968
rect 128852 26980 128914 26992
rect 128970 27968 129032 27980
rect 128970 26992 128982 27968
rect 129016 26992 129032 27968
rect 128970 26980 129032 26992
rect 129062 27968 129124 27980
rect 129062 26992 129078 27968
rect 129112 26992 129124 27968
rect 129062 26980 129124 26992
rect 129180 27968 129242 27980
rect 129180 26992 129192 27968
rect 129226 26992 129242 27968
rect 129180 26980 129242 26992
rect 129272 27968 129334 27980
rect 129272 26992 129288 27968
rect 129322 26992 129334 27968
rect 129272 26980 129334 26992
rect 129390 27968 129452 27980
rect 129390 26992 129402 27968
rect 129436 26992 129452 27968
rect 129390 26980 129452 26992
rect 129482 27968 129544 27980
rect 129482 26992 129498 27968
rect 129532 26992 129544 27968
rect 129482 26980 129544 26992
rect 129600 27968 129662 27980
rect 129600 26992 129612 27968
rect 129646 26992 129662 27968
rect 129600 26980 129662 26992
rect 129692 27968 129754 27980
rect 129692 26992 129708 27968
rect 129742 26992 129754 27968
rect 129692 26980 129754 26992
rect 129810 27968 129872 27980
rect 129810 26992 129822 27968
rect 129856 26992 129872 27968
rect 129810 26980 129872 26992
rect 129902 27968 129964 27980
rect 129902 26992 129918 27968
rect 129952 26992 129964 27968
rect 129902 26980 129964 26992
rect 130020 27968 130082 27980
rect 130020 26992 130032 27968
rect 130066 26992 130082 27968
rect 130020 26980 130082 26992
rect 130112 27968 130174 27980
rect 130112 26992 130128 27968
rect 130162 26992 130174 27968
rect 130112 26980 130174 26992
rect 130230 27968 130292 27980
rect 130230 26992 130242 27968
rect 130276 26992 130292 27968
rect 130230 26980 130292 26992
rect 130322 27968 130384 27980
rect 130322 26992 130338 27968
rect 130372 26992 130384 27968
rect 130322 26980 130384 26992
rect 130440 27968 130502 27980
rect 130440 26992 130452 27968
rect 130486 26992 130502 27968
rect 130440 26980 130502 26992
rect 130532 27968 130594 27980
rect 130532 26992 130548 27968
rect 130582 26992 130594 27968
rect 130532 26980 130594 26992
rect 130650 27968 130712 27980
rect 130650 26992 130662 27968
rect 130696 26992 130712 27968
rect 130650 26980 130712 26992
rect 130742 27968 130804 27980
rect 130742 26992 130758 27968
rect 130792 26992 130804 27968
rect 130742 26980 130804 26992
rect 130860 27968 130922 27980
rect 130860 26992 130872 27968
rect 130906 26992 130922 27968
rect 130860 26980 130922 26992
rect 130952 27968 131014 27980
rect 130952 26992 130968 27968
rect 131002 26992 131014 27968
rect 130952 26980 131014 26992
rect 131070 27968 131132 27980
rect 131070 26992 131082 27968
rect 131116 26992 131132 27968
rect 131070 26980 131132 26992
rect 131162 27968 131224 27980
rect 131162 26992 131178 27968
rect 131212 26992 131224 27968
rect 131162 26980 131224 26992
rect 131280 27968 131342 27980
rect 131280 26992 131292 27968
rect 131326 26992 131342 27968
rect 131280 26980 131342 26992
rect 131372 27968 131434 27980
rect 131372 26992 131388 27968
rect 131422 26992 131434 27968
rect 131372 26980 131434 26992
rect 131490 27968 131552 27980
rect 131490 26992 131502 27968
rect 131536 26992 131552 27968
rect 131490 26980 131552 26992
rect 131582 27968 131644 27980
rect 131582 26992 131598 27968
rect 131632 26992 131644 27968
rect 131582 26980 131644 26992
rect 131700 27968 131762 27980
rect 131700 26992 131712 27968
rect 131746 26992 131762 27968
rect 131700 26980 131762 26992
rect 131792 27968 131854 27980
rect 131792 26992 131808 27968
rect 131842 26992 131854 27968
rect 131792 26980 131854 26992
rect 131910 27968 131972 27980
rect 131910 26992 131922 27968
rect 131956 26992 131972 27968
rect 131910 26980 131972 26992
rect 132002 27968 132064 27980
rect 132002 26992 132018 27968
rect 132052 26992 132064 27968
rect 132002 26980 132064 26992
rect 132120 27968 132182 27980
rect 132120 26992 132132 27968
rect 132166 26992 132182 27968
rect 132120 26980 132182 26992
rect 132212 27968 132274 27980
rect 132212 26992 132228 27968
rect 132262 26992 132274 27968
rect 132212 26980 132274 26992
rect 132330 27968 132392 27980
rect 132330 26992 132342 27968
rect 132376 26992 132392 27968
rect 132330 26980 132392 26992
rect 132422 27968 132484 27980
rect 132422 26992 132438 27968
rect 132472 26992 132484 27968
rect 132422 26980 132484 26992
rect 132540 27968 132602 27980
rect 132540 26992 132552 27968
rect 132586 26992 132602 27968
rect 132540 26980 132602 26992
rect 132632 27968 132694 27980
rect 132632 26992 132648 27968
rect 132682 26992 132694 27968
rect 132632 26980 132694 26992
rect 132750 27968 132812 27980
rect 132750 26992 132762 27968
rect 132796 26992 132812 27968
rect 132750 26980 132812 26992
rect 132842 27968 132904 27980
rect 132842 26992 132858 27968
rect 132892 26992 132904 27968
rect 132842 26980 132904 26992
rect 132960 27968 133022 27980
rect 132960 26992 132972 27968
rect 133006 26992 133022 27968
rect 132960 26980 133022 26992
rect 133052 27968 133114 27980
rect 133052 26992 133068 27968
rect 133102 26992 133114 27968
rect 133052 26980 133114 26992
rect 133170 27968 133232 27980
rect 133170 26992 133182 27968
rect 133216 26992 133232 27968
rect 133170 26980 133232 26992
rect 133262 27968 133324 27980
rect 133262 26992 133278 27968
rect 133312 26992 133324 27968
rect 133262 26980 133324 26992
rect 133380 27968 133442 27980
rect 133380 26992 133392 27968
rect 133426 26992 133442 27968
rect 133380 26980 133442 26992
rect 133472 27968 133534 27980
rect 133472 26992 133488 27968
rect 133522 26992 133534 27968
rect 133472 26980 133534 26992
rect 133590 27968 133652 27980
rect 133590 26992 133602 27968
rect 133636 26992 133652 27968
rect 133590 26980 133652 26992
rect 133682 27968 133744 27980
rect 133682 26992 133698 27968
rect 133732 26992 133744 27968
rect 133682 26980 133744 26992
rect 133800 27968 133862 27980
rect 133800 26992 133812 27968
rect 133846 26992 133862 27968
rect 133800 26980 133862 26992
rect 133892 27968 133954 27980
rect 133892 26992 133908 27968
rect 133942 26992 133954 27968
rect 133892 26980 133954 26992
rect 134010 27968 134072 27980
rect 134010 26992 134022 27968
rect 134056 26992 134072 27968
rect 134010 26980 134072 26992
rect 134102 27968 134164 27980
rect 134102 26992 134118 27968
rect 134152 26992 134164 27968
rect 134102 26980 134164 26992
rect 134220 27968 134282 27980
rect 134220 26992 134232 27968
rect 134266 26992 134282 27968
rect 134220 26980 134282 26992
rect 134312 27968 134374 27980
rect 134312 26992 134328 27968
rect 134362 26992 134374 27968
rect 134312 26980 134374 26992
rect 134430 27968 134492 27980
rect 134430 26992 134442 27968
rect 134476 26992 134492 27968
rect 134430 26980 134492 26992
rect 134522 27968 134584 27980
rect 134522 26992 134538 27968
rect 134572 26992 134584 27968
rect 134522 26980 134584 26992
rect 134640 27968 134702 27980
rect 134640 26992 134652 27968
rect 134686 26992 134702 27968
rect 134640 26980 134702 26992
rect 134732 27968 134794 27980
rect 134732 26992 134748 27968
rect 134782 26992 134794 27968
rect 134732 26980 134794 26992
rect 134850 27968 134912 27980
rect 134850 26992 134862 27968
rect 134896 26992 134912 27968
rect 134850 26980 134912 26992
rect 134942 27968 135004 27980
rect 134942 26992 134958 27968
rect 134992 26992 135004 27968
rect 134942 26980 135004 26992
rect 135060 27968 135122 27980
rect 135060 26992 135072 27968
rect 135106 26992 135122 27968
rect 135060 26980 135122 26992
rect 135152 27968 135214 27980
rect 135152 26992 135168 27968
rect 135202 26992 135214 27968
rect 135152 26980 135214 26992
rect 126870 26750 126932 26762
rect 126870 25774 126882 26750
rect 126916 25774 126932 26750
rect 126870 25762 126932 25774
rect 126962 26750 127024 26762
rect 126962 25774 126978 26750
rect 127012 25774 127024 26750
rect 126962 25762 127024 25774
rect 127080 26750 127142 26762
rect 127080 25774 127092 26750
rect 127126 25774 127142 26750
rect 127080 25762 127142 25774
rect 127172 26750 127234 26762
rect 127172 25774 127188 26750
rect 127222 25774 127234 26750
rect 127172 25762 127234 25774
rect 127290 26750 127352 26762
rect 127290 25774 127302 26750
rect 127336 25774 127352 26750
rect 127290 25762 127352 25774
rect 127382 26750 127444 26762
rect 127382 25774 127398 26750
rect 127432 25774 127444 26750
rect 127382 25762 127444 25774
rect 127500 26750 127562 26762
rect 127500 25774 127512 26750
rect 127546 25774 127562 26750
rect 127500 25762 127562 25774
rect 127592 26750 127654 26762
rect 127592 25774 127608 26750
rect 127642 25774 127654 26750
rect 127592 25762 127654 25774
rect 127710 26750 127772 26762
rect 127710 25774 127722 26750
rect 127756 25774 127772 26750
rect 127710 25762 127772 25774
rect 127802 26750 127864 26762
rect 127802 25774 127818 26750
rect 127852 25774 127864 26750
rect 127802 25762 127864 25774
rect 127920 26750 127982 26762
rect 127920 25774 127932 26750
rect 127966 25774 127982 26750
rect 127920 25762 127982 25774
rect 128012 26750 128074 26762
rect 128012 25774 128028 26750
rect 128062 25774 128074 26750
rect 128012 25762 128074 25774
rect 128130 26750 128192 26762
rect 128130 25774 128142 26750
rect 128176 25774 128192 26750
rect 128130 25762 128192 25774
rect 128222 26750 128284 26762
rect 128222 25774 128238 26750
rect 128272 25774 128284 26750
rect 128222 25762 128284 25774
rect 128340 26750 128402 26762
rect 128340 25774 128352 26750
rect 128386 25774 128402 26750
rect 128340 25762 128402 25774
rect 128432 26750 128494 26762
rect 128432 25774 128448 26750
rect 128482 25774 128494 26750
rect 128432 25762 128494 25774
rect 128550 26750 128612 26762
rect 128550 25774 128562 26750
rect 128596 25774 128612 26750
rect 128550 25762 128612 25774
rect 128642 26750 128704 26762
rect 128642 25774 128658 26750
rect 128692 25774 128704 26750
rect 128642 25762 128704 25774
rect 128760 26750 128822 26762
rect 128760 25774 128772 26750
rect 128806 25774 128822 26750
rect 128760 25762 128822 25774
rect 128852 26750 128914 26762
rect 128852 25774 128868 26750
rect 128902 25774 128914 26750
rect 128852 25762 128914 25774
rect 128970 26750 129032 26762
rect 128970 25774 128982 26750
rect 129016 25774 129032 26750
rect 128970 25762 129032 25774
rect 129062 26750 129124 26762
rect 129062 25774 129078 26750
rect 129112 25774 129124 26750
rect 129062 25762 129124 25774
rect 129180 26750 129242 26762
rect 129180 25774 129192 26750
rect 129226 25774 129242 26750
rect 129180 25762 129242 25774
rect 129272 26750 129334 26762
rect 129272 25774 129288 26750
rect 129322 25774 129334 26750
rect 129272 25762 129334 25774
rect 129390 26750 129452 26762
rect 129390 25774 129402 26750
rect 129436 25774 129452 26750
rect 129390 25762 129452 25774
rect 129482 26750 129544 26762
rect 129482 25774 129498 26750
rect 129532 25774 129544 26750
rect 129482 25762 129544 25774
rect 129600 26750 129662 26762
rect 129600 25774 129612 26750
rect 129646 25774 129662 26750
rect 129600 25762 129662 25774
rect 129692 26750 129754 26762
rect 129692 25774 129708 26750
rect 129742 25774 129754 26750
rect 129692 25762 129754 25774
rect 129810 26750 129872 26762
rect 129810 25774 129822 26750
rect 129856 25774 129872 26750
rect 129810 25762 129872 25774
rect 129902 26750 129964 26762
rect 129902 25774 129918 26750
rect 129952 25774 129964 26750
rect 129902 25762 129964 25774
rect 130020 26750 130082 26762
rect 130020 25774 130032 26750
rect 130066 25774 130082 26750
rect 130020 25762 130082 25774
rect 130112 26750 130174 26762
rect 130112 25774 130128 26750
rect 130162 25774 130174 26750
rect 130112 25762 130174 25774
rect 130230 26750 130292 26762
rect 130230 25774 130242 26750
rect 130276 25774 130292 26750
rect 130230 25762 130292 25774
rect 130322 26750 130384 26762
rect 130322 25774 130338 26750
rect 130372 25774 130384 26750
rect 130322 25762 130384 25774
rect 130440 26750 130502 26762
rect 130440 25774 130452 26750
rect 130486 25774 130502 26750
rect 130440 25762 130502 25774
rect 130532 26750 130594 26762
rect 130532 25774 130548 26750
rect 130582 25774 130594 26750
rect 130532 25762 130594 25774
rect 130650 26750 130712 26762
rect 130650 25774 130662 26750
rect 130696 25774 130712 26750
rect 130650 25762 130712 25774
rect 130742 26750 130804 26762
rect 130742 25774 130758 26750
rect 130792 25774 130804 26750
rect 130742 25762 130804 25774
rect 130860 26750 130922 26762
rect 130860 25774 130872 26750
rect 130906 25774 130922 26750
rect 130860 25762 130922 25774
rect 130952 26750 131014 26762
rect 130952 25774 130968 26750
rect 131002 25774 131014 26750
rect 130952 25762 131014 25774
rect 131070 26750 131132 26762
rect 131070 25774 131082 26750
rect 131116 25774 131132 26750
rect 131070 25762 131132 25774
rect 131162 26750 131224 26762
rect 131162 25774 131178 26750
rect 131212 25774 131224 26750
rect 131162 25762 131224 25774
rect 131280 26750 131342 26762
rect 131280 25774 131292 26750
rect 131326 25774 131342 26750
rect 131280 25762 131342 25774
rect 131372 26750 131434 26762
rect 131372 25774 131388 26750
rect 131422 25774 131434 26750
rect 131372 25762 131434 25774
rect 131490 26750 131552 26762
rect 131490 25774 131502 26750
rect 131536 25774 131552 26750
rect 131490 25762 131552 25774
rect 131582 26750 131644 26762
rect 131582 25774 131598 26750
rect 131632 25774 131644 26750
rect 131582 25762 131644 25774
rect 131700 26750 131762 26762
rect 131700 25774 131712 26750
rect 131746 25774 131762 26750
rect 131700 25762 131762 25774
rect 131792 26750 131854 26762
rect 131792 25774 131808 26750
rect 131842 25774 131854 26750
rect 131792 25762 131854 25774
rect 131910 26750 131972 26762
rect 131910 25774 131922 26750
rect 131956 25774 131972 26750
rect 131910 25762 131972 25774
rect 132002 26750 132064 26762
rect 132002 25774 132018 26750
rect 132052 25774 132064 26750
rect 132002 25762 132064 25774
rect 132120 26750 132182 26762
rect 132120 25774 132132 26750
rect 132166 25774 132182 26750
rect 132120 25762 132182 25774
rect 132212 26750 132274 26762
rect 132212 25774 132228 26750
rect 132262 25774 132274 26750
rect 132212 25762 132274 25774
rect 132330 26750 132392 26762
rect 132330 25774 132342 26750
rect 132376 25774 132392 26750
rect 132330 25762 132392 25774
rect 132422 26750 132484 26762
rect 132422 25774 132438 26750
rect 132472 25774 132484 26750
rect 132422 25762 132484 25774
rect 132540 26750 132602 26762
rect 132540 25774 132552 26750
rect 132586 25774 132602 26750
rect 132540 25762 132602 25774
rect 132632 26750 132694 26762
rect 132632 25774 132648 26750
rect 132682 25774 132694 26750
rect 132632 25762 132694 25774
rect 132750 26750 132812 26762
rect 132750 25774 132762 26750
rect 132796 25774 132812 26750
rect 132750 25762 132812 25774
rect 132842 26750 132904 26762
rect 132842 25774 132858 26750
rect 132892 25774 132904 26750
rect 132842 25762 132904 25774
rect 132960 26750 133022 26762
rect 132960 25774 132972 26750
rect 133006 25774 133022 26750
rect 132960 25762 133022 25774
rect 133052 26750 133114 26762
rect 133052 25774 133068 26750
rect 133102 25774 133114 26750
rect 133052 25762 133114 25774
rect 133170 26750 133232 26762
rect 133170 25774 133182 26750
rect 133216 25774 133232 26750
rect 133170 25762 133232 25774
rect 133262 26750 133324 26762
rect 133262 25774 133278 26750
rect 133312 25774 133324 26750
rect 133262 25762 133324 25774
rect 133380 26750 133442 26762
rect 133380 25774 133392 26750
rect 133426 25774 133442 26750
rect 133380 25762 133442 25774
rect 133472 26750 133534 26762
rect 133472 25774 133488 26750
rect 133522 25774 133534 26750
rect 133472 25762 133534 25774
rect 133590 26750 133652 26762
rect 133590 25774 133602 26750
rect 133636 25774 133652 26750
rect 133590 25762 133652 25774
rect 133682 26750 133744 26762
rect 133682 25774 133698 26750
rect 133732 25774 133744 26750
rect 133682 25762 133744 25774
rect 133800 26750 133862 26762
rect 133800 25774 133812 26750
rect 133846 25774 133862 26750
rect 133800 25762 133862 25774
rect 133892 26750 133954 26762
rect 133892 25774 133908 26750
rect 133942 25774 133954 26750
rect 133892 25762 133954 25774
rect 134010 26750 134072 26762
rect 134010 25774 134022 26750
rect 134056 25774 134072 26750
rect 134010 25762 134072 25774
rect 134102 26750 134164 26762
rect 134102 25774 134118 26750
rect 134152 25774 134164 26750
rect 134102 25762 134164 25774
rect 134220 26750 134282 26762
rect 134220 25774 134232 26750
rect 134266 25774 134282 26750
rect 134220 25762 134282 25774
rect 134312 26750 134374 26762
rect 134312 25774 134328 26750
rect 134362 25774 134374 26750
rect 134312 25762 134374 25774
rect 134430 26750 134492 26762
rect 134430 25774 134442 26750
rect 134476 25774 134492 26750
rect 134430 25762 134492 25774
rect 134522 26750 134584 26762
rect 134522 25774 134538 26750
rect 134572 25774 134584 26750
rect 134522 25762 134584 25774
rect 134640 26750 134702 26762
rect 134640 25774 134652 26750
rect 134686 25774 134702 26750
rect 134640 25762 134702 25774
rect 134732 26750 134794 26762
rect 134732 25774 134748 26750
rect 134782 25774 134794 26750
rect 134732 25762 134794 25774
rect 134850 26750 134912 26762
rect 134850 25774 134862 26750
rect 134896 25774 134912 26750
rect 134850 25762 134912 25774
rect 134942 26750 135004 26762
rect 134942 25774 134958 26750
rect 134992 25774 135004 26750
rect 134942 25762 135004 25774
rect 135060 26750 135122 26762
rect 135060 25774 135072 26750
rect 135106 25774 135122 26750
rect 135060 25762 135122 25774
rect 135152 26750 135214 26762
rect 135152 25774 135168 26750
rect 135202 25774 135214 26750
rect 135152 25762 135214 25774
rect 122020 21884 122082 21896
rect 122020 20908 122032 21884
rect 122066 20908 122082 21884
rect 122020 20896 122082 20908
rect 122112 21884 122174 21896
rect 122112 20908 122128 21884
rect 122162 20908 122174 21884
rect 122112 20896 122174 20908
rect 122230 21884 122292 21896
rect 122230 20908 122242 21884
rect 122276 20908 122292 21884
rect 122230 20896 122292 20908
rect 122322 21884 122384 21896
rect 122322 20908 122338 21884
rect 122372 20908 122384 21884
rect 122322 20896 122384 20908
rect 122440 21884 122502 21896
rect 122440 20908 122452 21884
rect 122486 20908 122502 21884
rect 122440 20896 122502 20908
rect 122532 21884 122594 21896
rect 122532 20908 122548 21884
rect 122582 20908 122594 21884
rect 122532 20896 122594 20908
rect 122650 21884 122712 21896
rect 122650 20908 122662 21884
rect 122696 20908 122712 21884
rect 122650 20896 122712 20908
rect 122742 21884 122804 21896
rect 122742 20908 122758 21884
rect 122792 20908 122804 21884
rect 122742 20896 122804 20908
rect 122860 21884 122922 21896
rect 122860 20908 122872 21884
rect 122906 20908 122922 21884
rect 122860 20896 122922 20908
rect 122952 21884 123014 21896
rect 122952 20908 122968 21884
rect 123002 20908 123014 21884
rect 122952 20896 123014 20908
rect 123070 21884 123132 21896
rect 123070 20908 123082 21884
rect 123116 20908 123132 21884
rect 123070 20896 123132 20908
rect 123162 21884 123224 21896
rect 123162 20908 123178 21884
rect 123212 20908 123224 21884
rect 123162 20896 123224 20908
rect 123280 21884 123342 21896
rect 123280 20908 123292 21884
rect 123326 20908 123342 21884
rect 123280 20896 123342 20908
rect 123372 21884 123434 21896
rect 123372 20908 123388 21884
rect 123422 20908 123434 21884
rect 123372 20896 123434 20908
rect 123490 21884 123552 21896
rect 123490 20908 123502 21884
rect 123536 20908 123552 21884
rect 123490 20896 123552 20908
rect 123582 21884 123644 21896
rect 123582 20908 123598 21884
rect 123632 20908 123644 21884
rect 123582 20896 123644 20908
rect 123700 21884 123762 21896
rect 123700 20908 123712 21884
rect 123746 20908 123762 21884
rect 123700 20896 123762 20908
rect 123792 21884 123854 21896
rect 123792 20908 123808 21884
rect 123842 20908 123854 21884
rect 123792 20896 123854 20908
rect 123910 21884 123972 21896
rect 123910 20908 123922 21884
rect 123956 20908 123972 21884
rect 123910 20896 123972 20908
rect 124002 21884 124064 21896
rect 124002 20908 124018 21884
rect 124052 20908 124064 21884
rect 124002 20896 124064 20908
rect 124120 21884 124182 21896
rect 124120 20908 124132 21884
rect 124166 20908 124182 21884
rect 124120 20896 124182 20908
rect 124212 21884 124274 21896
rect 124212 20908 124228 21884
rect 124262 20908 124274 21884
rect 124212 20896 124274 20908
rect 124330 21884 124392 21896
rect 124330 20908 124342 21884
rect 124376 20908 124392 21884
rect 124330 20896 124392 20908
rect 124422 21884 124484 21896
rect 124422 20908 124438 21884
rect 124472 20908 124484 21884
rect 124422 20896 124484 20908
rect 124540 21884 124602 21896
rect 124540 20908 124552 21884
rect 124586 20908 124602 21884
rect 124540 20896 124602 20908
rect 124632 21884 124694 21896
rect 124632 20908 124648 21884
rect 124682 20908 124694 21884
rect 124632 20896 124694 20908
rect 124750 21884 124812 21896
rect 124750 20908 124762 21884
rect 124796 20908 124812 21884
rect 124750 20896 124812 20908
rect 124842 21884 124904 21896
rect 124842 20908 124858 21884
rect 124892 20908 124904 21884
rect 124842 20896 124904 20908
rect 124960 21884 125022 21896
rect 124960 20908 124972 21884
rect 125006 20908 125022 21884
rect 124960 20896 125022 20908
rect 125052 21884 125114 21896
rect 125052 20908 125068 21884
rect 125102 20908 125114 21884
rect 125052 20896 125114 20908
rect 125170 21884 125232 21896
rect 125170 20908 125182 21884
rect 125216 20908 125232 21884
rect 125170 20896 125232 20908
rect 125262 21884 125324 21896
rect 125262 20908 125278 21884
rect 125312 20908 125324 21884
rect 125262 20896 125324 20908
rect 125380 21884 125442 21896
rect 125380 20908 125392 21884
rect 125426 20908 125442 21884
rect 125380 20896 125442 20908
rect 125472 21884 125534 21896
rect 125472 20908 125488 21884
rect 125522 20908 125534 21884
rect 125472 20896 125534 20908
rect 125590 21884 125652 21896
rect 125590 20908 125602 21884
rect 125636 20908 125652 21884
rect 125590 20896 125652 20908
rect 125682 21884 125744 21896
rect 125682 20908 125698 21884
rect 125732 20908 125744 21884
rect 125682 20896 125744 20908
rect 119112 20260 119170 20272
rect 119112 19284 119124 20260
rect 119158 19284 119170 20260
rect 119112 19272 119170 19284
rect 119200 20260 119258 20272
rect 119200 19284 119212 20260
rect 119246 19284 119258 20260
rect 120056 20260 120118 20272
rect 119200 19272 119258 19284
rect 120056 19284 120068 20260
rect 120102 19284 120118 20260
rect 120056 19272 120118 19284
rect 120148 20260 120210 20272
rect 120148 19284 120164 20260
rect 120198 19284 120210 20260
rect 120148 19272 120210 19284
rect 120266 20260 120328 20272
rect 120266 19284 120278 20260
rect 120312 19284 120328 20260
rect 120266 19272 120328 19284
rect 120358 20260 120420 20272
rect 120358 19284 120374 20260
rect 120408 19284 120420 20260
rect 120358 19272 120420 19284
rect 120476 20260 120538 20272
rect 120476 19284 120488 20260
rect 120522 19284 120538 20260
rect 120476 19272 120538 19284
rect 120568 20260 120630 20272
rect 120568 19284 120584 20260
rect 120618 19284 120630 20260
rect 120568 19272 120630 19284
rect 120686 20260 120748 20272
rect 120686 19284 120698 20260
rect 120732 19284 120748 20260
rect 120686 19272 120748 19284
rect 120778 20260 120840 20272
rect 120778 19284 120794 20260
rect 120828 19284 120840 20260
rect 120778 19272 120840 19284
rect 116370 16906 116428 16918
rect 116370 16530 116382 16906
rect 116416 16530 116428 16906
rect 116370 16518 116428 16530
rect 116458 16906 116522 16918
rect 116458 16530 116476 16906
rect 116510 16530 116522 16906
rect 116458 16518 116522 16530
rect 116552 16906 116610 16918
rect 116552 16530 116564 16906
rect 116598 16530 116610 16906
rect 116552 16518 116610 16530
rect 116370 14860 116428 14872
rect 115844 14822 115902 14834
rect 115844 14646 115856 14822
rect 115890 14646 115902 14822
rect 115844 14634 115902 14646
rect 115932 14822 115990 14834
rect 115932 14646 115944 14822
rect 115978 14646 115990 14822
rect 115932 14634 115990 14646
rect 116370 14484 116382 14860
rect 116416 14484 116428 14860
rect 116370 14472 116428 14484
rect 116458 14860 116522 14872
rect 116458 14484 116476 14860
rect 116510 14484 116522 14860
rect 116458 14472 116522 14484
rect 116552 14860 116610 14872
rect 116552 14484 116564 14860
rect 116598 14484 116610 14860
rect 116552 14472 116610 14484
rect 119112 12106 119170 12118
rect 119112 11130 119124 12106
rect 119158 11130 119170 12106
rect 119112 11118 119170 11130
rect 119200 12106 119258 12118
rect 119200 11130 119212 12106
rect 119246 11130 119258 12106
rect 120056 12106 120118 12118
rect 119200 11118 119258 11130
rect 120056 11130 120068 12106
rect 120102 11130 120118 12106
rect 120056 11118 120118 11130
rect 120148 12106 120210 12118
rect 120148 11130 120164 12106
rect 120198 11130 120210 12106
rect 120148 11118 120210 11130
rect 120266 12106 120328 12118
rect 120266 11130 120278 12106
rect 120312 11130 120328 12106
rect 120266 11118 120328 11130
rect 120358 12106 120420 12118
rect 120358 11130 120374 12106
rect 120408 11130 120420 12106
rect 120358 11118 120420 11130
rect 120476 12106 120538 12118
rect 120476 11130 120488 12106
rect 120522 11130 120538 12106
rect 120476 11118 120538 11130
rect 120568 12106 120630 12118
rect 120568 11130 120584 12106
rect 120618 11130 120630 12106
rect 120568 11118 120630 11130
rect 120686 12106 120748 12118
rect 120686 11130 120698 12106
rect 120732 11130 120748 12106
rect 120686 11118 120748 11130
rect 120778 12106 120840 12118
rect 120778 11130 120794 12106
rect 120828 11130 120840 12106
rect 120778 11118 120840 11130
rect 122020 9082 122082 9094
rect 122020 8106 122032 9082
rect 122066 8106 122082 9082
rect 122020 8094 122082 8106
rect 122112 9082 122174 9094
rect 122112 8106 122128 9082
rect 122162 8106 122174 9082
rect 122112 8094 122174 8106
rect 122230 9082 122292 9094
rect 122230 8106 122242 9082
rect 122276 8106 122292 9082
rect 122230 8094 122292 8106
rect 122322 9082 122384 9094
rect 122322 8106 122338 9082
rect 122372 8106 122384 9082
rect 122322 8094 122384 8106
rect 122440 9082 122502 9094
rect 122440 8106 122452 9082
rect 122486 8106 122502 9082
rect 122440 8094 122502 8106
rect 122532 9082 122594 9094
rect 122532 8106 122548 9082
rect 122582 8106 122594 9082
rect 122532 8094 122594 8106
rect 122650 9082 122712 9094
rect 122650 8106 122662 9082
rect 122696 8106 122712 9082
rect 122650 8094 122712 8106
rect 122742 9082 122804 9094
rect 122742 8106 122758 9082
rect 122792 8106 122804 9082
rect 122742 8094 122804 8106
rect 122860 9082 122922 9094
rect 122860 8106 122872 9082
rect 122906 8106 122922 9082
rect 122860 8094 122922 8106
rect 122952 9082 123014 9094
rect 122952 8106 122968 9082
rect 123002 8106 123014 9082
rect 122952 8094 123014 8106
rect 123070 9082 123132 9094
rect 123070 8106 123082 9082
rect 123116 8106 123132 9082
rect 123070 8094 123132 8106
rect 123162 9082 123224 9094
rect 123162 8106 123178 9082
rect 123212 8106 123224 9082
rect 123162 8094 123224 8106
rect 123280 9082 123342 9094
rect 123280 8106 123292 9082
rect 123326 8106 123342 9082
rect 123280 8094 123342 8106
rect 123372 9082 123434 9094
rect 123372 8106 123388 9082
rect 123422 8106 123434 9082
rect 123372 8094 123434 8106
rect 123490 9082 123552 9094
rect 123490 8106 123502 9082
rect 123536 8106 123552 9082
rect 123490 8094 123552 8106
rect 123582 9082 123644 9094
rect 123582 8106 123598 9082
rect 123632 8106 123644 9082
rect 123582 8094 123644 8106
rect 123700 9082 123762 9094
rect 123700 8106 123712 9082
rect 123746 8106 123762 9082
rect 123700 8094 123762 8106
rect 123792 9082 123854 9094
rect 123792 8106 123808 9082
rect 123842 8106 123854 9082
rect 123792 8094 123854 8106
rect 123910 9082 123972 9094
rect 123910 8106 123922 9082
rect 123956 8106 123972 9082
rect 123910 8094 123972 8106
rect 124002 9082 124064 9094
rect 124002 8106 124018 9082
rect 124052 8106 124064 9082
rect 124002 8094 124064 8106
rect 124120 9082 124182 9094
rect 124120 8106 124132 9082
rect 124166 8106 124182 9082
rect 124120 8094 124182 8106
rect 124212 9082 124274 9094
rect 124212 8106 124228 9082
rect 124262 8106 124274 9082
rect 124212 8094 124274 8106
rect 124330 9082 124392 9094
rect 124330 8106 124342 9082
rect 124376 8106 124392 9082
rect 124330 8094 124392 8106
rect 124422 9082 124484 9094
rect 124422 8106 124438 9082
rect 124472 8106 124484 9082
rect 124422 8094 124484 8106
rect 124540 9082 124602 9094
rect 124540 8106 124552 9082
rect 124586 8106 124602 9082
rect 124540 8094 124602 8106
rect 124632 9082 124694 9094
rect 124632 8106 124648 9082
rect 124682 8106 124694 9082
rect 124632 8094 124694 8106
rect 124750 9082 124812 9094
rect 124750 8106 124762 9082
rect 124796 8106 124812 9082
rect 124750 8094 124812 8106
rect 124842 9082 124904 9094
rect 124842 8106 124858 9082
rect 124892 8106 124904 9082
rect 124842 8094 124904 8106
rect 124960 9082 125022 9094
rect 124960 8106 124972 9082
rect 125006 8106 125022 9082
rect 124960 8094 125022 8106
rect 125052 9082 125114 9094
rect 125052 8106 125068 9082
rect 125102 8106 125114 9082
rect 125052 8094 125114 8106
rect 125170 9082 125232 9094
rect 125170 8106 125182 9082
rect 125216 8106 125232 9082
rect 125170 8094 125232 8106
rect 125262 9082 125324 9094
rect 125262 8106 125278 9082
rect 125312 8106 125324 9082
rect 125262 8094 125324 8106
rect 125380 9082 125442 9094
rect 125380 8106 125392 9082
rect 125426 8106 125442 9082
rect 125380 8094 125442 8106
rect 125472 9082 125534 9094
rect 125472 8106 125488 9082
rect 125522 8106 125534 9082
rect 125472 8094 125534 8106
rect 125590 9082 125652 9094
rect 125590 8106 125602 9082
rect 125636 8106 125652 9082
rect 125590 8094 125652 8106
rect 125682 9082 125744 9094
rect 125682 8106 125698 9082
rect 125732 8106 125744 9082
rect 125682 8094 125744 8106
<< pdiff >>
rect 119108 19032 119170 19044
rect 119108 18056 119120 19032
rect 119154 18056 119170 19032
rect 119108 18044 119170 18056
rect 119200 19032 119266 19044
rect 119200 18056 119216 19032
rect 119250 18056 119266 19032
rect 119200 18044 119266 18056
rect 119296 19032 119358 19044
rect 119296 18056 119312 19032
rect 119346 18056 119358 19032
rect 119846 19032 119908 19044
rect 119296 18044 119358 18056
rect 119846 18056 119858 19032
rect 119892 18056 119908 19032
rect 119846 18044 119908 18056
rect 119938 19032 120000 19044
rect 119938 18056 119954 19032
rect 119988 18056 120000 19032
rect 119938 18044 120000 18056
rect 120056 19032 120118 19044
rect 120056 18056 120068 19032
rect 120102 18056 120118 19032
rect 120056 18044 120118 18056
rect 120148 19032 120210 19044
rect 120148 18056 120164 19032
rect 120198 18056 120210 19032
rect 120148 18044 120210 18056
rect 120266 19032 120328 19044
rect 120266 18056 120278 19032
rect 120312 18056 120328 19032
rect 120266 18044 120328 18056
rect 120358 19032 120420 19044
rect 120358 18056 120374 19032
rect 120408 18056 120420 19032
rect 120358 18044 120420 18056
rect 120476 19032 120538 19044
rect 120476 18056 120488 19032
rect 120522 18056 120538 19032
rect 120476 18044 120538 18056
rect 120568 19032 120630 19044
rect 120568 18056 120584 19032
rect 120618 18056 120630 19032
rect 120568 18044 120630 18056
rect 120686 19032 120748 19044
rect 120686 18056 120698 19032
rect 120732 18056 120748 19032
rect 120686 18044 120748 18056
rect 120778 19032 120840 19044
rect 120778 18056 120794 19032
rect 120828 18056 120840 19032
rect 120778 18044 120840 18056
rect 120896 19032 120958 19044
rect 120896 18056 120908 19032
rect 120942 18056 120958 19032
rect 120896 18044 120958 18056
rect 120988 19032 121050 19044
rect 120988 18056 121004 19032
rect 121038 18056 121050 19032
rect 120988 18044 121050 18056
rect 121106 19032 121168 19044
rect 121106 18056 121118 19032
rect 121152 18056 121168 19032
rect 121106 18044 121168 18056
rect 121198 19032 121260 19044
rect 121198 18056 121214 19032
rect 121248 18056 121260 19032
rect 121198 18044 121260 18056
rect 121316 19032 121378 19044
rect 121316 18056 121328 19032
rect 121362 18056 121378 19032
rect 121316 18044 121378 18056
rect 121408 19032 121470 19044
rect 121408 18056 121424 19032
rect 121458 18056 121470 19032
rect 121408 18044 121470 18056
rect 122020 20268 122082 20280
rect 122020 19292 122032 20268
rect 122066 19292 122082 20268
rect 122020 19280 122082 19292
rect 122112 20268 122174 20280
rect 122112 19292 122128 20268
rect 122162 19292 122174 20268
rect 122112 19280 122174 19292
rect 122230 20268 122292 20280
rect 122230 19292 122242 20268
rect 122276 19292 122292 20268
rect 122230 19280 122292 19292
rect 122322 20268 122384 20280
rect 122322 19292 122338 20268
rect 122372 19292 122384 20268
rect 122322 19280 122384 19292
rect 122440 20268 122502 20280
rect 122440 19292 122452 20268
rect 122486 19292 122502 20268
rect 122440 19280 122502 19292
rect 122532 20268 122594 20280
rect 122532 19292 122548 20268
rect 122582 19292 122594 20268
rect 122532 19280 122594 19292
rect 122650 20268 122712 20280
rect 122650 19292 122662 20268
rect 122696 19292 122712 20268
rect 122650 19280 122712 19292
rect 122742 20268 122804 20280
rect 122742 19292 122758 20268
rect 122792 19292 122804 20268
rect 122742 19280 122804 19292
rect 122860 20268 122922 20280
rect 122860 19292 122872 20268
rect 122906 19292 122922 20268
rect 122860 19280 122922 19292
rect 122952 20268 123014 20280
rect 122952 19292 122968 20268
rect 123002 19292 123014 20268
rect 122952 19280 123014 19292
rect 123070 20268 123132 20280
rect 123070 19292 123082 20268
rect 123116 19292 123132 20268
rect 123070 19280 123132 19292
rect 123162 20268 123224 20280
rect 123162 19292 123178 20268
rect 123212 19292 123224 20268
rect 123162 19280 123224 19292
rect 123280 20268 123342 20280
rect 123280 19292 123292 20268
rect 123326 19292 123342 20268
rect 123280 19280 123342 19292
rect 123372 20268 123434 20280
rect 123372 19292 123388 20268
rect 123422 19292 123434 20268
rect 123372 19280 123434 19292
rect 123490 20268 123552 20280
rect 123490 19292 123502 20268
rect 123536 19292 123552 20268
rect 123490 19280 123552 19292
rect 123582 20268 123644 20280
rect 123582 19292 123598 20268
rect 123632 19292 123644 20268
rect 123582 19280 123644 19292
rect 123700 20268 123762 20280
rect 123700 19292 123712 20268
rect 123746 19292 123762 20268
rect 123700 19280 123762 19292
rect 123792 20268 123854 20280
rect 123792 19292 123808 20268
rect 123842 19292 123854 20268
rect 123792 19280 123854 19292
rect 123910 20268 123972 20280
rect 123910 19292 123922 20268
rect 123956 19292 123972 20268
rect 123910 19280 123972 19292
rect 124002 20268 124064 20280
rect 124002 19292 124018 20268
rect 124052 19292 124064 20268
rect 124002 19280 124064 19292
rect 124120 20268 124182 20280
rect 124120 19292 124132 20268
rect 124166 19292 124182 20268
rect 124120 19280 124182 19292
rect 124212 20268 124274 20280
rect 124212 19292 124228 20268
rect 124262 19292 124274 20268
rect 124212 19280 124274 19292
rect 124330 20268 124392 20280
rect 124330 19292 124342 20268
rect 124376 19292 124392 20268
rect 124330 19280 124392 19292
rect 124422 20268 124484 20280
rect 124422 19292 124438 20268
rect 124472 19292 124484 20268
rect 124422 19280 124484 19292
rect 124540 20268 124602 20280
rect 124540 19292 124552 20268
rect 124586 19292 124602 20268
rect 124540 19280 124602 19292
rect 124632 20268 124694 20280
rect 124632 19292 124648 20268
rect 124682 19292 124694 20268
rect 124632 19280 124694 19292
rect 124750 20268 124812 20280
rect 124750 19292 124762 20268
rect 124796 19292 124812 20268
rect 124750 19280 124812 19292
rect 124842 20268 124904 20280
rect 124842 19292 124858 20268
rect 124892 19292 124904 20268
rect 124842 19280 124904 19292
rect 124960 20268 125022 20280
rect 124960 19292 124972 20268
rect 125006 19292 125022 20268
rect 124960 19280 125022 19292
rect 125052 20268 125114 20280
rect 125052 19292 125068 20268
rect 125102 19292 125114 20268
rect 125052 19280 125114 19292
rect 125170 20268 125232 20280
rect 125170 19292 125182 20268
rect 125216 19292 125232 20268
rect 125170 19280 125232 19292
rect 125262 20268 125324 20280
rect 125262 19292 125278 20268
rect 125312 19292 125324 20268
rect 125262 19280 125324 19292
rect 125380 20268 125442 20280
rect 125380 19292 125392 20268
rect 125426 19292 125442 20268
rect 125380 19280 125442 19292
rect 125472 20268 125534 20280
rect 125472 19292 125488 20268
rect 125522 19292 125534 20268
rect 125472 19280 125534 19292
rect 125590 20268 125652 20280
rect 125590 19292 125602 20268
rect 125636 19292 125652 20268
rect 125590 19280 125652 19292
rect 125682 20268 125744 20280
rect 125682 19292 125698 20268
rect 125732 19292 125744 20268
rect 125682 19280 125744 19292
rect 122020 19032 122082 19044
rect 122020 18056 122032 19032
rect 122066 18056 122082 19032
rect 122020 18044 122082 18056
rect 122112 19032 122174 19044
rect 122112 18056 122128 19032
rect 122162 18056 122174 19032
rect 122112 18044 122174 18056
rect 122230 19032 122292 19044
rect 122230 18056 122242 19032
rect 122276 18056 122292 19032
rect 122230 18044 122292 18056
rect 122322 19032 122384 19044
rect 122322 18056 122338 19032
rect 122372 18056 122384 19032
rect 122322 18044 122384 18056
rect 122440 19032 122502 19044
rect 122440 18056 122452 19032
rect 122486 18056 122502 19032
rect 122440 18044 122502 18056
rect 122532 19032 122594 19044
rect 122532 18056 122548 19032
rect 122582 18056 122594 19032
rect 122532 18044 122594 18056
rect 122650 19032 122712 19044
rect 122650 18056 122662 19032
rect 122696 18056 122712 19032
rect 122650 18044 122712 18056
rect 122742 19032 122804 19044
rect 122742 18056 122758 19032
rect 122792 18056 122804 19032
rect 122742 18044 122804 18056
rect 122860 19032 122922 19044
rect 122860 18056 122872 19032
rect 122906 18056 122922 19032
rect 122860 18044 122922 18056
rect 122952 19032 123014 19044
rect 122952 18056 122968 19032
rect 123002 18056 123014 19032
rect 122952 18044 123014 18056
rect 123070 19032 123132 19044
rect 123070 18056 123082 19032
rect 123116 18056 123132 19032
rect 123070 18044 123132 18056
rect 123162 19032 123224 19044
rect 123162 18056 123178 19032
rect 123212 18056 123224 19032
rect 123162 18044 123224 18056
rect 123280 19032 123342 19044
rect 123280 18056 123292 19032
rect 123326 18056 123342 19032
rect 123280 18044 123342 18056
rect 123372 19032 123434 19044
rect 123372 18056 123388 19032
rect 123422 18056 123434 19032
rect 123372 18044 123434 18056
rect 123490 19032 123552 19044
rect 123490 18056 123502 19032
rect 123536 18056 123552 19032
rect 123490 18044 123552 18056
rect 123582 19032 123644 19044
rect 123582 18056 123598 19032
rect 123632 18056 123644 19032
rect 123582 18044 123644 18056
rect 123700 19032 123762 19044
rect 123700 18056 123712 19032
rect 123746 18056 123762 19032
rect 123700 18044 123762 18056
rect 123792 19032 123854 19044
rect 123792 18056 123808 19032
rect 123842 18056 123854 19032
rect 123792 18044 123854 18056
rect 123910 19032 123972 19044
rect 123910 18056 123922 19032
rect 123956 18056 123972 19032
rect 123910 18044 123972 18056
rect 124002 19032 124064 19044
rect 124002 18056 124018 19032
rect 124052 18056 124064 19032
rect 124002 18044 124064 18056
rect 124120 19032 124182 19044
rect 124120 18056 124132 19032
rect 124166 18056 124182 19032
rect 124120 18044 124182 18056
rect 124212 19032 124274 19044
rect 124212 18056 124228 19032
rect 124262 18056 124274 19032
rect 124212 18044 124274 18056
rect 124330 19032 124392 19044
rect 124330 18056 124342 19032
rect 124376 18056 124392 19032
rect 124330 18044 124392 18056
rect 124422 19032 124484 19044
rect 124422 18056 124438 19032
rect 124472 18056 124484 19032
rect 124422 18044 124484 18056
rect 124540 19032 124602 19044
rect 124540 18056 124552 19032
rect 124586 18056 124602 19032
rect 124540 18044 124602 18056
rect 124632 19032 124694 19044
rect 124632 18056 124648 19032
rect 124682 18056 124694 19032
rect 124632 18044 124694 18056
rect 124750 19032 124812 19044
rect 124750 18056 124762 19032
rect 124796 18056 124812 19032
rect 124750 18044 124812 18056
rect 124842 19032 124904 19044
rect 124842 18056 124858 19032
rect 124892 18056 124904 19032
rect 124842 18044 124904 18056
rect 124960 19032 125022 19044
rect 124960 18056 124972 19032
rect 125006 18056 125022 19032
rect 124960 18044 125022 18056
rect 125052 19032 125114 19044
rect 125052 18056 125068 19032
rect 125102 18056 125114 19032
rect 125052 18044 125114 18056
rect 125170 19032 125232 19044
rect 125170 18056 125182 19032
rect 125216 18056 125232 19032
rect 125170 18044 125232 18056
rect 125262 19032 125324 19044
rect 125262 18056 125278 19032
rect 125312 18056 125324 19032
rect 125262 18044 125324 18056
rect 125380 19032 125442 19044
rect 125380 18056 125392 19032
rect 125426 18056 125442 19032
rect 125380 18044 125442 18056
rect 125472 19032 125534 19044
rect 125472 18056 125488 19032
rect 125522 18056 125534 19032
rect 125472 18044 125534 18056
rect 125590 19032 125652 19044
rect 125590 18056 125602 19032
rect 125636 18056 125652 19032
rect 125590 18044 125652 18056
rect 125682 19032 125744 19044
rect 125682 18056 125698 19032
rect 125732 18056 125744 19032
rect 125682 18044 125744 18056
rect 126870 22740 126932 22752
rect 126870 21764 126882 22740
rect 126916 21764 126932 22740
rect 126870 21752 126932 21764
rect 126962 22740 127024 22752
rect 126962 21764 126978 22740
rect 127012 21764 127024 22740
rect 126962 21752 127024 21764
rect 127080 22740 127142 22752
rect 127080 21764 127092 22740
rect 127126 21764 127142 22740
rect 127080 21752 127142 21764
rect 127172 22740 127234 22752
rect 127172 21764 127188 22740
rect 127222 21764 127234 22740
rect 127172 21752 127234 21764
rect 127290 22740 127352 22752
rect 127290 21764 127302 22740
rect 127336 21764 127352 22740
rect 127290 21752 127352 21764
rect 127382 22740 127444 22752
rect 127382 21764 127398 22740
rect 127432 21764 127444 22740
rect 127382 21752 127444 21764
rect 127500 22740 127562 22752
rect 127500 21764 127512 22740
rect 127546 21764 127562 22740
rect 127500 21752 127562 21764
rect 127592 22740 127654 22752
rect 127592 21764 127608 22740
rect 127642 21764 127654 22740
rect 127592 21752 127654 21764
rect 127710 22740 127772 22752
rect 127710 21764 127722 22740
rect 127756 21764 127772 22740
rect 127710 21752 127772 21764
rect 127802 22740 127864 22752
rect 127802 21764 127818 22740
rect 127852 21764 127864 22740
rect 127802 21752 127864 21764
rect 127920 22740 127982 22752
rect 127920 21764 127932 22740
rect 127966 21764 127982 22740
rect 127920 21752 127982 21764
rect 128012 22740 128074 22752
rect 128012 21764 128028 22740
rect 128062 21764 128074 22740
rect 128012 21752 128074 21764
rect 128130 22740 128192 22752
rect 128130 21764 128142 22740
rect 128176 21764 128192 22740
rect 128130 21752 128192 21764
rect 128222 22740 128284 22752
rect 128222 21764 128238 22740
rect 128272 21764 128284 22740
rect 128222 21752 128284 21764
rect 128340 22740 128402 22752
rect 128340 21764 128352 22740
rect 128386 21764 128402 22740
rect 128340 21752 128402 21764
rect 128432 22740 128494 22752
rect 128432 21764 128448 22740
rect 128482 21764 128494 22740
rect 128432 21752 128494 21764
rect 128550 22740 128612 22752
rect 128550 21764 128562 22740
rect 128596 21764 128612 22740
rect 128550 21752 128612 21764
rect 128642 22740 128704 22752
rect 128642 21764 128658 22740
rect 128692 21764 128704 22740
rect 128642 21752 128704 21764
rect 128760 22740 128822 22752
rect 128760 21764 128772 22740
rect 128806 21764 128822 22740
rect 128760 21752 128822 21764
rect 128852 22740 128914 22752
rect 128852 21764 128868 22740
rect 128902 21764 128914 22740
rect 128852 21752 128914 21764
rect 128970 22740 129032 22752
rect 128970 21764 128982 22740
rect 129016 21764 129032 22740
rect 128970 21752 129032 21764
rect 129062 22740 129124 22752
rect 129062 21764 129078 22740
rect 129112 21764 129124 22740
rect 129062 21752 129124 21764
rect 129180 22740 129242 22752
rect 129180 21764 129192 22740
rect 129226 21764 129242 22740
rect 129180 21752 129242 21764
rect 129272 22740 129334 22752
rect 129272 21764 129288 22740
rect 129322 21764 129334 22740
rect 129272 21752 129334 21764
rect 129390 22740 129452 22752
rect 129390 21764 129402 22740
rect 129436 21764 129452 22740
rect 129390 21752 129452 21764
rect 129482 22740 129544 22752
rect 129482 21764 129498 22740
rect 129532 21764 129544 22740
rect 129482 21752 129544 21764
rect 129600 22740 129662 22752
rect 129600 21764 129612 22740
rect 129646 21764 129662 22740
rect 129600 21752 129662 21764
rect 129692 22740 129754 22752
rect 129692 21764 129708 22740
rect 129742 21764 129754 22740
rect 129692 21752 129754 21764
rect 129810 22740 129872 22752
rect 129810 21764 129822 22740
rect 129856 21764 129872 22740
rect 129810 21752 129872 21764
rect 129902 22740 129964 22752
rect 129902 21764 129918 22740
rect 129952 21764 129964 22740
rect 129902 21752 129964 21764
rect 130020 22740 130082 22752
rect 130020 21764 130032 22740
rect 130066 21764 130082 22740
rect 130020 21752 130082 21764
rect 130112 22740 130174 22752
rect 130112 21764 130128 22740
rect 130162 21764 130174 22740
rect 130112 21752 130174 21764
rect 130230 22740 130292 22752
rect 130230 21764 130242 22740
rect 130276 21764 130292 22740
rect 130230 21752 130292 21764
rect 130322 22740 130384 22752
rect 130322 21764 130338 22740
rect 130372 21764 130384 22740
rect 130322 21752 130384 21764
rect 130440 22740 130502 22752
rect 130440 21764 130452 22740
rect 130486 21764 130502 22740
rect 130440 21752 130502 21764
rect 130532 22740 130594 22752
rect 130532 21764 130548 22740
rect 130582 21764 130594 22740
rect 130532 21752 130594 21764
rect 130650 22740 130712 22752
rect 130650 21764 130662 22740
rect 130696 21764 130712 22740
rect 130650 21752 130712 21764
rect 130742 22740 130804 22752
rect 130742 21764 130758 22740
rect 130792 21764 130804 22740
rect 130742 21752 130804 21764
rect 130860 22740 130922 22752
rect 130860 21764 130872 22740
rect 130906 21764 130922 22740
rect 130860 21752 130922 21764
rect 130952 22740 131014 22752
rect 130952 21764 130968 22740
rect 131002 21764 131014 22740
rect 130952 21752 131014 21764
rect 131070 22740 131132 22752
rect 131070 21764 131082 22740
rect 131116 21764 131132 22740
rect 131070 21752 131132 21764
rect 131162 22740 131224 22752
rect 131162 21764 131178 22740
rect 131212 21764 131224 22740
rect 131162 21752 131224 21764
rect 131280 22740 131342 22752
rect 131280 21764 131292 22740
rect 131326 21764 131342 22740
rect 131280 21752 131342 21764
rect 131372 22740 131434 22752
rect 131372 21764 131388 22740
rect 131422 21764 131434 22740
rect 131372 21752 131434 21764
rect 131490 22740 131552 22752
rect 131490 21764 131502 22740
rect 131536 21764 131552 22740
rect 131490 21752 131552 21764
rect 131582 22740 131644 22752
rect 131582 21764 131598 22740
rect 131632 21764 131644 22740
rect 131582 21752 131644 21764
rect 131700 22740 131762 22752
rect 131700 21764 131712 22740
rect 131746 21764 131762 22740
rect 131700 21752 131762 21764
rect 131792 22740 131854 22752
rect 131792 21764 131808 22740
rect 131842 21764 131854 22740
rect 131792 21752 131854 21764
rect 131910 22740 131972 22752
rect 131910 21764 131922 22740
rect 131956 21764 131972 22740
rect 131910 21752 131972 21764
rect 132002 22740 132064 22752
rect 132002 21764 132018 22740
rect 132052 21764 132064 22740
rect 132002 21752 132064 21764
rect 132120 22740 132182 22752
rect 132120 21764 132132 22740
rect 132166 21764 132182 22740
rect 132120 21752 132182 21764
rect 132212 22740 132274 22752
rect 132212 21764 132228 22740
rect 132262 21764 132274 22740
rect 132212 21752 132274 21764
rect 132330 22740 132392 22752
rect 132330 21764 132342 22740
rect 132376 21764 132392 22740
rect 132330 21752 132392 21764
rect 132422 22740 132484 22752
rect 132422 21764 132438 22740
rect 132472 21764 132484 22740
rect 132422 21752 132484 21764
rect 132540 22740 132602 22752
rect 132540 21764 132552 22740
rect 132586 21764 132602 22740
rect 132540 21752 132602 21764
rect 132632 22740 132694 22752
rect 132632 21764 132648 22740
rect 132682 21764 132694 22740
rect 132632 21752 132694 21764
rect 132750 22740 132812 22752
rect 132750 21764 132762 22740
rect 132796 21764 132812 22740
rect 132750 21752 132812 21764
rect 132842 22740 132904 22752
rect 132842 21764 132858 22740
rect 132892 21764 132904 22740
rect 132842 21752 132904 21764
rect 132960 22740 133022 22752
rect 132960 21764 132972 22740
rect 133006 21764 133022 22740
rect 132960 21752 133022 21764
rect 133052 22740 133114 22752
rect 133052 21764 133068 22740
rect 133102 21764 133114 22740
rect 133052 21752 133114 21764
rect 133170 22740 133232 22752
rect 133170 21764 133182 22740
rect 133216 21764 133232 22740
rect 133170 21752 133232 21764
rect 133262 22740 133324 22752
rect 133262 21764 133278 22740
rect 133312 21764 133324 22740
rect 133262 21752 133324 21764
rect 133380 22740 133442 22752
rect 133380 21764 133392 22740
rect 133426 21764 133442 22740
rect 133380 21752 133442 21764
rect 133472 22740 133534 22752
rect 133472 21764 133488 22740
rect 133522 21764 133534 22740
rect 133472 21752 133534 21764
rect 133590 22740 133652 22752
rect 133590 21764 133602 22740
rect 133636 21764 133652 22740
rect 133590 21752 133652 21764
rect 133682 22740 133744 22752
rect 133682 21764 133698 22740
rect 133732 21764 133744 22740
rect 133682 21752 133744 21764
rect 133800 22740 133862 22752
rect 133800 21764 133812 22740
rect 133846 21764 133862 22740
rect 133800 21752 133862 21764
rect 133892 22740 133954 22752
rect 133892 21764 133908 22740
rect 133942 21764 133954 22740
rect 133892 21752 133954 21764
rect 134010 22740 134072 22752
rect 134010 21764 134022 22740
rect 134056 21764 134072 22740
rect 134010 21752 134072 21764
rect 134102 22740 134164 22752
rect 134102 21764 134118 22740
rect 134152 21764 134164 22740
rect 134102 21752 134164 21764
rect 134220 22740 134282 22752
rect 134220 21764 134232 22740
rect 134266 21764 134282 22740
rect 134220 21752 134282 21764
rect 134312 22740 134374 22752
rect 134312 21764 134328 22740
rect 134362 21764 134374 22740
rect 134312 21752 134374 21764
rect 134430 22740 134492 22752
rect 134430 21764 134442 22740
rect 134476 21764 134492 22740
rect 134430 21752 134492 21764
rect 134522 22740 134584 22752
rect 134522 21764 134538 22740
rect 134572 21764 134584 22740
rect 134522 21752 134584 21764
rect 134640 22740 134702 22752
rect 134640 21764 134652 22740
rect 134686 21764 134702 22740
rect 134640 21752 134702 21764
rect 134732 22740 134794 22752
rect 134732 21764 134748 22740
rect 134782 21764 134794 22740
rect 134732 21752 134794 21764
rect 134850 22740 134912 22752
rect 134850 21764 134862 22740
rect 134896 21764 134912 22740
rect 134850 21752 134912 21764
rect 134942 22740 135004 22752
rect 134942 21764 134958 22740
rect 134992 21764 135004 22740
rect 134942 21752 135004 21764
rect 135060 22740 135122 22752
rect 135060 21764 135072 22740
rect 135106 21764 135122 22740
rect 135060 21752 135122 21764
rect 135152 22740 135214 22752
rect 135152 21764 135168 22740
rect 135202 21764 135214 22740
rect 135152 21752 135214 21764
rect 126870 21504 126932 21516
rect 126870 20528 126882 21504
rect 126916 20528 126932 21504
rect 126870 20516 126932 20528
rect 126962 21504 127024 21516
rect 126962 20528 126978 21504
rect 127012 20528 127024 21504
rect 126962 20516 127024 20528
rect 127080 21504 127142 21516
rect 127080 20528 127092 21504
rect 127126 20528 127142 21504
rect 127080 20516 127142 20528
rect 127172 21504 127234 21516
rect 127172 20528 127188 21504
rect 127222 20528 127234 21504
rect 127172 20516 127234 20528
rect 127290 21504 127352 21516
rect 127290 20528 127302 21504
rect 127336 20528 127352 21504
rect 127290 20516 127352 20528
rect 127382 21504 127444 21516
rect 127382 20528 127398 21504
rect 127432 20528 127444 21504
rect 127382 20516 127444 20528
rect 127500 21504 127562 21516
rect 127500 20528 127512 21504
rect 127546 20528 127562 21504
rect 127500 20516 127562 20528
rect 127592 21504 127654 21516
rect 127592 20528 127608 21504
rect 127642 20528 127654 21504
rect 127592 20516 127654 20528
rect 127710 21504 127772 21516
rect 127710 20528 127722 21504
rect 127756 20528 127772 21504
rect 127710 20516 127772 20528
rect 127802 21504 127864 21516
rect 127802 20528 127818 21504
rect 127852 20528 127864 21504
rect 127802 20516 127864 20528
rect 127920 21504 127982 21516
rect 127920 20528 127932 21504
rect 127966 20528 127982 21504
rect 127920 20516 127982 20528
rect 128012 21504 128074 21516
rect 128012 20528 128028 21504
rect 128062 20528 128074 21504
rect 128012 20516 128074 20528
rect 128130 21504 128192 21516
rect 128130 20528 128142 21504
rect 128176 20528 128192 21504
rect 128130 20516 128192 20528
rect 128222 21504 128284 21516
rect 128222 20528 128238 21504
rect 128272 20528 128284 21504
rect 128222 20516 128284 20528
rect 128340 21504 128402 21516
rect 128340 20528 128352 21504
rect 128386 20528 128402 21504
rect 128340 20516 128402 20528
rect 128432 21504 128494 21516
rect 128432 20528 128448 21504
rect 128482 20528 128494 21504
rect 128432 20516 128494 20528
rect 128550 21504 128612 21516
rect 128550 20528 128562 21504
rect 128596 20528 128612 21504
rect 128550 20516 128612 20528
rect 128642 21504 128704 21516
rect 128642 20528 128658 21504
rect 128692 20528 128704 21504
rect 128642 20516 128704 20528
rect 128760 21504 128822 21516
rect 128760 20528 128772 21504
rect 128806 20528 128822 21504
rect 128760 20516 128822 20528
rect 128852 21504 128914 21516
rect 128852 20528 128868 21504
rect 128902 20528 128914 21504
rect 128852 20516 128914 20528
rect 128970 21504 129032 21516
rect 128970 20528 128982 21504
rect 129016 20528 129032 21504
rect 128970 20516 129032 20528
rect 129062 21504 129124 21516
rect 129062 20528 129078 21504
rect 129112 20528 129124 21504
rect 129062 20516 129124 20528
rect 129180 21504 129242 21516
rect 129180 20528 129192 21504
rect 129226 20528 129242 21504
rect 129180 20516 129242 20528
rect 129272 21504 129334 21516
rect 129272 20528 129288 21504
rect 129322 20528 129334 21504
rect 129272 20516 129334 20528
rect 129390 21504 129452 21516
rect 129390 20528 129402 21504
rect 129436 20528 129452 21504
rect 129390 20516 129452 20528
rect 129482 21504 129544 21516
rect 129482 20528 129498 21504
rect 129532 20528 129544 21504
rect 129482 20516 129544 20528
rect 129600 21504 129662 21516
rect 129600 20528 129612 21504
rect 129646 20528 129662 21504
rect 129600 20516 129662 20528
rect 129692 21504 129754 21516
rect 129692 20528 129708 21504
rect 129742 20528 129754 21504
rect 129692 20516 129754 20528
rect 129810 21504 129872 21516
rect 129810 20528 129822 21504
rect 129856 20528 129872 21504
rect 129810 20516 129872 20528
rect 129902 21504 129964 21516
rect 129902 20528 129918 21504
rect 129952 20528 129964 21504
rect 129902 20516 129964 20528
rect 130020 21504 130082 21516
rect 130020 20528 130032 21504
rect 130066 20528 130082 21504
rect 130020 20516 130082 20528
rect 130112 21504 130174 21516
rect 130112 20528 130128 21504
rect 130162 20528 130174 21504
rect 130112 20516 130174 20528
rect 130230 21504 130292 21516
rect 130230 20528 130242 21504
rect 130276 20528 130292 21504
rect 130230 20516 130292 20528
rect 130322 21504 130384 21516
rect 130322 20528 130338 21504
rect 130372 20528 130384 21504
rect 130322 20516 130384 20528
rect 130440 21504 130502 21516
rect 130440 20528 130452 21504
rect 130486 20528 130502 21504
rect 130440 20516 130502 20528
rect 130532 21504 130594 21516
rect 130532 20528 130548 21504
rect 130582 20528 130594 21504
rect 130532 20516 130594 20528
rect 130650 21504 130712 21516
rect 130650 20528 130662 21504
rect 130696 20528 130712 21504
rect 130650 20516 130712 20528
rect 130742 21504 130804 21516
rect 130742 20528 130758 21504
rect 130792 20528 130804 21504
rect 130742 20516 130804 20528
rect 130860 21504 130922 21516
rect 130860 20528 130872 21504
rect 130906 20528 130922 21504
rect 130860 20516 130922 20528
rect 130952 21504 131014 21516
rect 130952 20528 130968 21504
rect 131002 20528 131014 21504
rect 130952 20516 131014 20528
rect 131070 21504 131132 21516
rect 131070 20528 131082 21504
rect 131116 20528 131132 21504
rect 131070 20516 131132 20528
rect 131162 21504 131224 21516
rect 131162 20528 131178 21504
rect 131212 20528 131224 21504
rect 131162 20516 131224 20528
rect 131280 21504 131342 21516
rect 131280 20528 131292 21504
rect 131326 20528 131342 21504
rect 131280 20516 131342 20528
rect 131372 21504 131434 21516
rect 131372 20528 131388 21504
rect 131422 20528 131434 21504
rect 131372 20516 131434 20528
rect 131490 21504 131552 21516
rect 131490 20528 131502 21504
rect 131536 20528 131552 21504
rect 131490 20516 131552 20528
rect 131582 21504 131644 21516
rect 131582 20528 131598 21504
rect 131632 20528 131644 21504
rect 131582 20516 131644 20528
rect 131700 21504 131762 21516
rect 131700 20528 131712 21504
rect 131746 20528 131762 21504
rect 131700 20516 131762 20528
rect 131792 21504 131854 21516
rect 131792 20528 131808 21504
rect 131842 20528 131854 21504
rect 131792 20516 131854 20528
rect 131910 21504 131972 21516
rect 131910 20528 131922 21504
rect 131956 20528 131972 21504
rect 131910 20516 131972 20528
rect 132002 21504 132064 21516
rect 132002 20528 132018 21504
rect 132052 20528 132064 21504
rect 132002 20516 132064 20528
rect 132120 21504 132182 21516
rect 132120 20528 132132 21504
rect 132166 20528 132182 21504
rect 132120 20516 132182 20528
rect 132212 21504 132274 21516
rect 132212 20528 132228 21504
rect 132262 20528 132274 21504
rect 132212 20516 132274 20528
rect 132330 21504 132392 21516
rect 132330 20528 132342 21504
rect 132376 20528 132392 21504
rect 132330 20516 132392 20528
rect 132422 21504 132484 21516
rect 132422 20528 132438 21504
rect 132472 20528 132484 21504
rect 132422 20516 132484 20528
rect 132540 21504 132602 21516
rect 132540 20528 132552 21504
rect 132586 20528 132602 21504
rect 132540 20516 132602 20528
rect 132632 21504 132694 21516
rect 132632 20528 132648 21504
rect 132682 20528 132694 21504
rect 132632 20516 132694 20528
rect 132750 21504 132812 21516
rect 132750 20528 132762 21504
rect 132796 20528 132812 21504
rect 132750 20516 132812 20528
rect 132842 21504 132904 21516
rect 132842 20528 132858 21504
rect 132892 20528 132904 21504
rect 132842 20516 132904 20528
rect 132960 21504 133022 21516
rect 132960 20528 132972 21504
rect 133006 20528 133022 21504
rect 132960 20516 133022 20528
rect 133052 21504 133114 21516
rect 133052 20528 133068 21504
rect 133102 20528 133114 21504
rect 133052 20516 133114 20528
rect 133170 21504 133232 21516
rect 133170 20528 133182 21504
rect 133216 20528 133232 21504
rect 133170 20516 133232 20528
rect 133262 21504 133324 21516
rect 133262 20528 133278 21504
rect 133312 20528 133324 21504
rect 133262 20516 133324 20528
rect 133380 21504 133442 21516
rect 133380 20528 133392 21504
rect 133426 20528 133442 21504
rect 133380 20516 133442 20528
rect 133472 21504 133534 21516
rect 133472 20528 133488 21504
rect 133522 20528 133534 21504
rect 133472 20516 133534 20528
rect 133590 21504 133652 21516
rect 133590 20528 133602 21504
rect 133636 20528 133652 21504
rect 133590 20516 133652 20528
rect 133682 21504 133744 21516
rect 133682 20528 133698 21504
rect 133732 20528 133744 21504
rect 133682 20516 133744 20528
rect 133800 21504 133862 21516
rect 133800 20528 133812 21504
rect 133846 20528 133862 21504
rect 133800 20516 133862 20528
rect 133892 21504 133954 21516
rect 133892 20528 133908 21504
rect 133942 20528 133954 21504
rect 133892 20516 133954 20528
rect 134010 21504 134072 21516
rect 134010 20528 134022 21504
rect 134056 20528 134072 21504
rect 134010 20516 134072 20528
rect 134102 21504 134164 21516
rect 134102 20528 134118 21504
rect 134152 20528 134164 21504
rect 134102 20516 134164 20528
rect 134220 21504 134282 21516
rect 134220 20528 134232 21504
rect 134266 20528 134282 21504
rect 134220 20516 134282 20528
rect 134312 21504 134374 21516
rect 134312 20528 134328 21504
rect 134362 20528 134374 21504
rect 134312 20516 134374 20528
rect 134430 21504 134492 21516
rect 134430 20528 134442 21504
rect 134476 20528 134492 21504
rect 134430 20516 134492 20528
rect 134522 21504 134584 21516
rect 134522 20528 134538 21504
rect 134572 20528 134584 21504
rect 134522 20516 134584 20528
rect 134640 21504 134702 21516
rect 134640 20528 134652 21504
rect 134686 20528 134702 21504
rect 134640 20516 134702 20528
rect 134732 21504 134794 21516
rect 134732 20528 134748 21504
rect 134782 20528 134794 21504
rect 134732 20516 134794 20528
rect 134850 21504 134912 21516
rect 134850 20528 134862 21504
rect 134896 20528 134912 21504
rect 134850 20516 134912 20528
rect 134942 21504 135004 21516
rect 134942 20528 134958 21504
rect 134992 20528 135004 21504
rect 134942 20516 135004 20528
rect 135060 21504 135122 21516
rect 135060 20528 135072 21504
rect 135106 20528 135122 21504
rect 135060 20516 135122 20528
rect 135152 21504 135214 21516
rect 135152 20528 135168 21504
rect 135202 20528 135214 21504
rect 135152 20516 135214 20528
rect 126870 20268 126932 20280
rect 126870 19292 126882 20268
rect 126916 19292 126932 20268
rect 126870 19280 126932 19292
rect 126962 20268 127024 20280
rect 126962 19292 126978 20268
rect 127012 19292 127024 20268
rect 126962 19280 127024 19292
rect 127080 20268 127142 20280
rect 127080 19292 127092 20268
rect 127126 19292 127142 20268
rect 127080 19280 127142 19292
rect 127172 20268 127234 20280
rect 127172 19292 127188 20268
rect 127222 19292 127234 20268
rect 127172 19280 127234 19292
rect 127290 20268 127352 20280
rect 127290 19292 127302 20268
rect 127336 19292 127352 20268
rect 127290 19280 127352 19292
rect 127382 20268 127444 20280
rect 127382 19292 127398 20268
rect 127432 19292 127444 20268
rect 127382 19280 127444 19292
rect 127500 20268 127562 20280
rect 127500 19292 127512 20268
rect 127546 19292 127562 20268
rect 127500 19280 127562 19292
rect 127592 20268 127654 20280
rect 127592 19292 127608 20268
rect 127642 19292 127654 20268
rect 127592 19280 127654 19292
rect 127710 20268 127772 20280
rect 127710 19292 127722 20268
rect 127756 19292 127772 20268
rect 127710 19280 127772 19292
rect 127802 20268 127864 20280
rect 127802 19292 127818 20268
rect 127852 19292 127864 20268
rect 127802 19280 127864 19292
rect 127920 20268 127982 20280
rect 127920 19292 127932 20268
rect 127966 19292 127982 20268
rect 127920 19280 127982 19292
rect 128012 20268 128074 20280
rect 128012 19292 128028 20268
rect 128062 19292 128074 20268
rect 128012 19280 128074 19292
rect 128130 20268 128192 20280
rect 128130 19292 128142 20268
rect 128176 19292 128192 20268
rect 128130 19280 128192 19292
rect 128222 20268 128284 20280
rect 128222 19292 128238 20268
rect 128272 19292 128284 20268
rect 128222 19280 128284 19292
rect 128340 20268 128402 20280
rect 128340 19292 128352 20268
rect 128386 19292 128402 20268
rect 128340 19280 128402 19292
rect 128432 20268 128494 20280
rect 128432 19292 128448 20268
rect 128482 19292 128494 20268
rect 128432 19280 128494 19292
rect 128550 20268 128612 20280
rect 128550 19292 128562 20268
rect 128596 19292 128612 20268
rect 128550 19280 128612 19292
rect 128642 20268 128704 20280
rect 128642 19292 128658 20268
rect 128692 19292 128704 20268
rect 128642 19280 128704 19292
rect 128760 20268 128822 20280
rect 128760 19292 128772 20268
rect 128806 19292 128822 20268
rect 128760 19280 128822 19292
rect 128852 20268 128914 20280
rect 128852 19292 128868 20268
rect 128902 19292 128914 20268
rect 128852 19280 128914 19292
rect 128970 20268 129032 20280
rect 128970 19292 128982 20268
rect 129016 19292 129032 20268
rect 128970 19280 129032 19292
rect 129062 20268 129124 20280
rect 129062 19292 129078 20268
rect 129112 19292 129124 20268
rect 129062 19280 129124 19292
rect 129180 20268 129242 20280
rect 129180 19292 129192 20268
rect 129226 19292 129242 20268
rect 129180 19280 129242 19292
rect 129272 20268 129334 20280
rect 129272 19292 129288 20268
rect 129322 19292 129334 20268
rect 129272 19280 129334 19292
rect 129390 20268 129452 20280
rect 129390 19292 129402 20268
rect 129436 19292 129452 20268
rect 129390 19280 129452 19292
rect 129482 20268 129544 20280
rect 129482 19292 129498 20268
rect 129532 19292 129544 20268
rect 129482 19280 129544 19292
rect 129600 20268 129662 20280
rect 129600 19292 129612 20268
rect 129646 19292 129662 20268
rect 129600 19280 129662 19292
rect 129692 20268 129754 20280
rect 129692 19292 129708 20268
rect 129742 19292 129754 20268
rect 129692 19280 129754 19292
rect 129810 20268 129872 20280
rect 129810 19292 129822 20268
rect 129856 19292 129872 20268
rect 129810 19280 129872 19292
rect 129902 20268 129964 20280
rect 129902 19292 129918 20268
rect 129952 19292 129964 20268
rect 129902 19280 129964 19292
rect 130020 20268 130082 20280
rect 130020 19292 130032 20268
rect 130066 19292 130082 20268
rect 130020 19280 130082 19292
rect 130112 20268 130174 20280
rect 130112 19292 130128 20268
rect 130162 19292 130174 20268
rect 130112 19280 130174 19292
rect 130230 20268 130292 20280
rect 130230 19292 130242 20268
rect 130276 19292 130292 20268
rect 130230 19280 130292 19292
rect 130322 20268 130384 20280
rect 130322 19292 130338 20268
rect 130372 19292 130384 20268
rect 130322 19280 130384 19292
rect 130440 20268 130502 20280
rect 130440 19292 130452 20268
rect 130486 19292 130502 20268
rect 130440 19280 130502 19292
rect 130532 20268 130594 20280
rect 130532 19292 130548 20268
rect 130582 19292 130594 20268
rect 130532 19280 130594 19292
rect 130650 20268 130712 20280
rect 130650 19292 130662 20268
rect 130696 19292 130712 20268
rect 130650 19280 130712 19292
rect 130742 20268 130804 20280
rect 130742 19292 130758 20268
rect 130792 19292 130804 20268
rect 130742 19280 130804 19292
rect 130860 20268 130922 20280
rect 130860 19292 130872 20268
rect 130906 19292 130922 20268
rect 130860 19280 130922 19292
rect 130952 20268 131014 20280
rect 130952 19292 130968 20268
rect 131002 19292 131014 20268
rect 130952 19280 131014 19292
rect 131070 20268 131132 20280
rect 131070 19292 131082 20268
rect 131116 19292 131132 20268
rect 131070 19280 131132 19292
rect 131162 20268 131224 20280
rect 131162 19292 131178 20268
rect 131212 19292 131224 20268
rect 131162 19280 131224 19292
rect 131280 20268 131342 20280
rect 131280 19292 131292 20268
rect 131326 19292 131342 20268
rect 131280 19280 131342 19292
rect 131372 20268 131434 20280
rect 131372 19292 131388 20268
rect 131422 19292 131434 20268
rect 131372 19280 131434 19292
rect 131490 20268 131552 20280
rect 131490 19292 131502 20268
rect 131536 19292 131552 20268
rect 131490 19280 131552 19292
rect 131582 20268 131644 20280
rect 131582 19292 131598 20268
rect 131632 19292 131644 20268
rect 131582 19280 131644 19292
rect 131700 20268 131762 20280
rect 131700 19292 131712 20268
rect 131746 19292 131762 20268
rect 131700 19280 131762 19292
rect 131792 20268 131854 20280
rect 131792 19292 131808 20268
rect 131842 19292 131854 20268
rect 131792 19280 131854 19292
rect 131910 20268 131972 20280
rect 131910 19292 131922 20268
rect 131956 19292 131972 20268
rect 131910 19280 131972 19292
rect 132002 20268 132064 20280
rect 132002 19292 132018 20268
rect 132052 19292 132064 20268
rect 132002 19280 132064 19292
rect 132120 20268 132182 20280
rect 132120 19292 132132 20268
rect 132166 19292 132182 20268
rect 132120 19280 132182 19292
rect 132212 20268 132274 20280
rect 132212 19292 132228 20268
rect 132262 19292 132274 20268
rect 132212 19280 132274 19292
rect 132330 20268 132392 20280
rect 132330 19292 132342 20268
rect 132376 19292 132392 20268
rect 132330 19280 132392 19292
rect 132422 20268 132484 20280
rect 132422 19292 132438 20268
rect 132472 19292 132484 20268
rect 132422 19280 132484 19292
rect 132540 20268 132602 20280
rect 132540 19292 132552 20268
rect 132586 19292 132602 20268
rect 132540 19280 132602 19292
rect 132632 20268 132694 20280
rect 132632 19292 132648 20268
rect 132682 19292 132694 20268
rect 132632 19280 132694 19292
rect 132750 20268 132812 20280
rect 132750 19292 132762 20268
rect 132796 19292 132812 20268
rect 132750 19280 132812 19292
rect 132842 20268 132904 20280
rect 132842 19292 132858 20268
rect 132892 19292 132904 20268
rect 132842 19280 132904 19292
rect 132960 20268 133022 20280
rect 132960 19292 132972 20268
rect 133006 19292 133022 20268
rect 132960 19280 133022 19292
rect 133052 20268 133114 20280
rect 133052 19292 133068 20268
rect 133102 19292 133114 20268
rect 133052 19280 133114 19292
rect 133170 20268 133232 20280
rect 133170 19292 133182 20268
rect 133216 19292 133232 20268
rect 133170 19280 133232 19292
rect 133262 20268 133324 20280
rect 133262 19292 133278 20268
rect 133312 19292 133324 20268
rect 133262 19280 133324 19292
rect 133380 20268 133442 20280
rect 133380 19292 133392 20268
rect 133426 19292 133442 20268
rect 133380 19280 133442 19292
rect 133472 20268 133534 20280
rect 133472 19292 133488 20268
rect 133522 19292 133534 20268
rect 133472 19280 133534 19292
rect 133590 20268 133652 20280
rect 133590 19292 133602 20268
rect 133636 19292 133652 20268
rect 133590 19280 133652 19292
rect 133682 20268 133744 20280
rect 133682 19292 133698 20268
rect 133732 19292 133744 20268
rect 133682 19280 133744 19292
rect 133800 20268 133862 20280
rect 133800 19292 133812 20268
rect 133846 19292 133862 20268
rect 133800 19280 133862 19292
rect 133892 20268 133954 20280
rect 133892 19292 133908 20268
rect 133942 19292 133954 20268
rect 133892 19280 133954 19292
rect 134010 20268 134072 20280
rect 134010 19292 134022 20268
rect 134056 19292 134072 20268
rect 134010 19280 134072 19292
rect 134102 20268 134164 20280
rect 134102 19292 134118 20268
rect 134152 19292 134164 20268
rect 134102 19280 134164 19292
rect 134220 20268 134282 20280
rect 134220 19292 134232 20268
rect 134266 19292 134282 20268
rect 134220 19280 134282 19292
rect 134312 20268 134374 20280
rect 134312 19292 134328 20268
rect 134362 19292 134374 20268
rect 134312 19280 134374 19292
rect 134430 20268 134492 20280
rect 134430 19292 134442 20268
rect 134476 19292 134492 20268
rect 134430 19280 134492 19292
rect 134522 20268 134584 20280
rect 134522 19292 134538 20268
rect 134572 19292 134584 20268
rect 134522 19280 134584 19292
rect 134640 20268 134702 20280
rect 134640 19292 134652 20268
rect 134686 19292 134702 20268
rect 134640 19280 134702 19292
rect 134732 20268 134794 20280
rect 134732 19292 134748 20268
rect 134782 19292 134794 20268
rect 134732 19280 134794 19292
rect 134850 20268 134912 20280
rect 134850 19292 134862 20268
rect 134896 19292 134912 20268
rect 134850 19280 134912 19292
rect 134942 20268 135004 20280
rect 134942 19292 134958 20268
rect 134992 19292 135004 20268
rect 134942 19280 135004 19292
rect 135060 20268 135122 20280
rect 135060 19292 135072 20268
rect 135106 19292 135122 20268
rect 135060 19280 135122 19292
rect 135152 20268 135214 20280
rect 135152 19292 135168 20268
rect 135202 19292 135214 20268
rect 135152 19280 135214 19292
rect 126870 19032 126932 19044
rect 126870 18056 126882 19032
rect 126916 18056 126932 19032
rect 126870 18044 126932 18056
rect 126962 19032 127024 19044
rect 126962 18056 126978 19032
rect 127012 18056 127024 19032
rect 126962 18044 127024 18056
rect 127080 19032 127142 19044
rect 127080 18056 127092 19032
rect 127126 18056 127142 19032
rect 127080 18044 127142 18056
rect 127172 19032 127234 19044
rect 127172 18056 127188 19032
rect 127222 18056 127234 19032
rect 127172 18044 127234 18056
rect 127290 19032 127352 19044
rect 127290 18056 127302 19032
rect 127336 18056 127352 19032
rect 127290 18044 127352 18056
rect 127382 19032 127444 19044
rect 127382 18056 127398 19032
rect 127432 18056 127444 19032
rect 127382 18044 127444 18056
rect 127500 19032 127562 19044
rect 127500 18056 127512 19032
rect 127546 18056 127562 19032
rect 127500 18044 127562 18056
rect 127592 19032 127654 19044
rect 127592 18056 127608 19032
rect 127642 18056 127654 19032
rect 127592 18044 127654 18056
rect 127710 19032 127772 19044
rect 127710 18056 127722 19032
rect 127756 18056 127772 19032
rect 127710 18044 127772 18056
rect 127802 19032 127864 19044
rect 127802 18056 127818 19032
rect 127852 18056 127864 19032
rect 127802 18044 127864 18056
rect 127920 19032 127982 19044
rect 127920 18056 127932 19032
rect 127966 18056 127982 19032
rect 127920 18044 127982 18056
rect 128012 19032 128074 19044
rect 128012 18056 128028 19032
rect 128062 18056 128074 19032
rect 128012 18044 128074 18056
rect 128130 19032 128192 19044
rect 128130 18056 128142 19032
rect 128176 18056 128192 19032
rect 128130 18044 128192 18056
rect 128222 19032 128284 19044
rect 128222 18056 128238 19032
rect 128272 18056 128284 19032
rect 128222 18044 128284 18056
rect 128340 19032 128402 19044
rect 128340 18056 128352 19032
rect 128386 18056 128402 19032
rect 128340 18044 128402 18056
rect 128432 19032 128494 19044
rect 128432 18056 128448 19032
rect 128482 18056 128494 19032
rect 128432 18044 128494 18056
rect 128550 19032 128612 19044
rect 128550 18056 128562 19032
rect 128596 18056 128612 19032
rect 128550 18044 128612 18056
rect 128642 19032 128704 19044
rect 128642 18056 128658 19032
rect 128692 18056 128704 19032
rect 128642 18044 128704 18056
rect 128760 19032 128822 19044
rect 128760 18056 128772 19032
rect 128806 18056 128822 19032
rect 128760 18044 128822 18056
rect 128852 19032 128914 19044
rect 128852 18056 128868 19032
rect 128902 18056 128914 19032
rect 128852 18044 128914 18056
rect 128970 19032 129032 19044
rect 128970 18056 128982 19032
rect 129016 18056 129032 19032
rect 128970 18044 129032 18056
rect 129062 19032 129124 19044
rect 129062 18056 129078 19032
rect 129112 18056 129124 19032
rect 129062 18044 129124 18056
rect 129180 19032 129242 19044
rect 129180 18056 129192 19032
rect 129226 18056 129242 19032
rect 129180 18044 129242 18056
rect 129272 19032 129334 19044
rect 129272 18056 129288 19032
rect 129322 18056 129334 19032
rect 129272 18044 129334 18056
rect 129390 19032 129452 19044
rect 129390 18056 129402 19032
rect 129436 18056 129452 19032
rect 129390 18044 129452 18056
rect 129482 19032 129544 19044
rect 129482 18056 129498 19032
rect 129532 18056 129544 19032
rect 129482 18044 129544 18056
rect 129600 19032 129662 19044
rect 129600 18056 129612 19032
rect 129646 18056 129662 19032
rect 129600 18044 129662 18056
rect 129692 19032 129754 19044
rect 129692 18056 129708 19032
rect 129742 18056 129754 19032
rect 129692 18044 129754 18056
rect 129810 19032 129872 19044
rect 129810 18056 129822 19032
rect 129856 18056 129872 19032
rect 129810 18044 129872 18056
rect 129902 19032 129964 19044
rect 129902 18056 129918 19032
rect 129952 18056 129964 19032
rect 129902 18044 129964 18056
rect 130020 19032 130082 19044
rect 130020 18056 130032 19032
rect 130066 18056 130082 19032
rect 130020 18044 130082 18056
rect 130112 19032 130174 19044
rect 130112 18056 130128 19032
rect 130162 18056 130174 19032
rect 130112 18044 130174 18056
rect 130230 19032 130292 19044
rect 130230 18056 130242 19032
rect 130276 18056 130292 19032
rect 130230 18044 130292 18056
rect 130322 19032 130384 19044
rect 130322 18056 130338 19032
rect 130372 18056 130384 19032
rect 130322 18044 130384 18056
rect 130440 19032 130502 19044
rect 130440 18056 130452 19032
rect 130486 18056 130502 19032
rect 130440 18044 130502 18056
rect 130532 19032 130594 19044
rect 130532 18056 130548 19032
rect 130582 18056 130594 19032
rect 130532 18044 130594 18056
rect 130650 19032 130712 19044
rect 130650 18056 130662 19032
rect 130696 18056 130712 19032
rect 130650 18044 130712 18056
rect 130742 19032 130804 19044
rect 130742 18056 130758 19032
rect 130792 18056 130804 19032
rect 130742 18044 130804 18056
rect 130860 19032 130922 19044
rect 130860 18056 130872 19032
rect 130906 18056 130922 19032
rect 130860 18044 130922 18056
rect 130952 19032 131014 19044
rect 130952 18056 130968 19032
rect 131002 18056 131014 19032
rect 130952 18044 131014 18056
rect 131070 19032 131132 19044
rect 131070 18056 131082 19032
rect 131116 18056 131132 19032
rect 131070 18044 131132 18056
rect 131162 19032 131224 19044
rect 131162 18056 131178 19032
rect 131212 18056 131224 19032
rect 131162 18044 131224 18056
rect 131280 19032 131342 19044
rect 131280 18056 131292 19032
rect 131326 18056 131342 19032
rect 131280 18044 131342 18056
rect 131372 19032 131434 19044
rect 131372 18056 131388 19032
rect 131422 18056 131434 19032
rect 131372 18044 131434 18056
rect 131490 19032 131552 19044
rect 131490 18056 131502 19032
rect 131536 18056 131552 19032
rect 131490 18044 131552 18056
rect 131582 19032 131644 19044
rect 131582 18056 131598 19032
rect 131632 18056 131644 19032
rect 131582 18044 131644 18056
rect 131700 19032 131762 19044
rect 131700 18056 131712 19032
rect 131746 18056 131762 19032
rect 131700 18044 131762 18056
rect 131792 19032 131854 19044
rect 131792 18056 131808 19032
rect 131842 18056 131854 19032
rect 131792 18044 131854 18056
rect 131910 19032 131972 19044
rect 131910 18056 131922 19032
rect 131956 18056 131972 19032
rect 131910 18044 131972 18056
rect 132002 19032 132064 19044
rect 132002 18056 132018 19032
rect 132052 18056 132064 19032
rect 132002 18044 132064 18056
rect 132120 19032 132182 19044
rect 132120 18056 132132 19032
rect 132166 18056 132182 19032
rect 132120 18044 132182 18056
rect 132212 19032 132274 19044
rect 132212 18056 132228 19032
rect 132262 18056 132274 19032
rect 132212 18044 132274 18056
rect 132330 19032 132392 19044
rect 132330 18056 132342 19032
rect 132376 18056 132392 19032
rect 132330 18044 132392 18056
rect 132422 19032 132484 19044
rect 132422 18056 132438 19032
rect 132472 18056 132484 19032
rect 132422 18044 132484 18056
rect 132540 19032 132602 19044
rect 132540 18056 132552 19032
rect 132586 18056 132602 19032
rect 132540 18044 132602 18056
rect 132632 19032 132694 19044
rect 132632 18056 132648 19032
rect 132682 18056 132694 19032
rect 132632 18044 132694 18056
rect 132750 19032 132812 19044
rect 132750 18056 132762 19032
rect 132796 18056 132812 19032
rect 132750 18044 132812 18056
rect 132842 19032 132904 19044
rect 132842 18056 132858 19032
rect 132892 18056 132904 19032
rect 132842 18044 132904 18056
rect 132960 19032 133022 19044
rect 132960 18056 132972 19032
rect 133006 18056 133022 19032
rect 132960 18044 133022 18056
rect 133052 19032 133114 19044
rect 133052 18056 133068 19032
rect 133102 18056 133114 19032
rect 133052 18044 133114 18056
rect 133170 19032 133232 19044
rect 133170 18056 133182 19032
rect 133216 18056 133232 19032
rect 133170 18044 133232 18056
rect 133262 19032 133324 19044
rect 133262 18056 133278 19032
rect 133312 18056 133324 19032
rect 133262 18044 133324 18056
rect 133380 19032 133442 19044
rect 133380 18056 133392 19032
rect 133426 18056 133442 19032
rect 133380 18044 133442 18056
rect 133472 19032 133534 19044
rect 133472 18056 133488 19032
rect 133522 18056 133534 19032
rect 133472 18044 133534 18056
rect 133590 19032 133652 19044
rect 133590 18056 133602 19032
rect 133636 18056 133652 19032
rect 133590 18044 133652 18056
rect 133682 19032 133744 19044
rect 133682 18056 133698 19032
rect 133732 18056 133744 19032
rect 133682 18044 133744 18056
rect 133800 19032 133862 19044
rect 133800 18056 133812 19032
rect 133846 18056 133862 19032
rect 133800 18044 133862 18056
rect 133892 19032 133954 19044
rect 133892 18056 133908 19032
rect 133942 18056 133954 19032
rect 133892 18044 133954 18056
rect 134010 19032 134072 19044
rect 134010 18056 134022 19032
rect 134056 18056 134072 19032
rect 134010 18044 134072 18056
rect 134102 19032 134164 19044
rect 134102 18056 134118 19032
rect 134152 18056 134164 19032
rect 134102 18044 134164 18056
rect 134220 19032 134282 19044
rect 134220 18056 134232 19032
rect 134266 18056 134282 19032
rect 134220 18044 134282 18056
rect 134312 19032 134374 19044
rect 134312 18056 134328 19032
rect 134362 18056 134374 19032
rect 134312 18044 134374 18056
rect 134430 19032 134492 19044
rect 134430 18056 134442 19032
rect 134476 18056 134492 19032
rect 134430 18044 134492 18056
rect 134522 19032 134584 19044
rect 134522 18056 134538 19032
rect 134572 18056 134584 19032
rect 134522 18044 134584 18056
rect 134640 19032 134702 19044
rect 134640 18056 134652 19032
rect 134686 18056 134702 19032
rect 134640 18044 134702 18056
rect 134732 19032 134794 19044
rect 134732 18056 134748 19032
rect 134782 18056 134794 19032
rect 134732 18044 134794 18056
rect 134850 19032 134912 19044
rect 134850 18056 134862 19032
rect 134896 18056 134912 19032
rect 134850 18044 134912 18056
rect 134942 19032 135004 19044
rect 134942 18056 134958 19032
rect 134992 18056 135004 19032
rect 134942 18044 135004 18056
rect 135060 19032 135122 19044
rect 135060 18056 135072 19032
rect 135106 18056 135122 19032
rect 135060 18044 135122 18056
rect 135152 19032 135214 19044
rect 135152 18056 135168 19032
rect 135202 18056 135214 19032
rect 135152 18044 135214 18056
rect 116370 16286 116428 16298
rect 116370 15910 116382 16286
rect 116416 15910 116428 16286
rect 116370 15898 116428 15910
rect 116458 16286 116522 16298
rect 116458 15910 116476 16286
rect 116510 15910 116522 16286
rect 116458 15898 116522 15910
rect 116552 16286 116610 16298
rect 116552 15910 116564 16286
rect 116598 15910 116610 16286
rect 116552 15898 116610 15910
rect 115844 15478 115902 15490
rect 115844 15102 115856 15478
rect 115890 15102 115902 15478
rect 115844 15090 115902 15102
rect 115932 15478 115990 15490
rect 115932 15102 115944 15478
rect 115978 15102 115990 15478
rect 116370 15480 116428 15492
rect 115932 15090 115990 15102
rect 116370 15104 116382 15480
rect 116416 15104 116428 15480
rect 116370 15092 116428 15104
rect 116458 15480 116522 15492
rect 116458 15104 116476 15480
rect 116510 15104 116522 15480
rect 116458 15092 116522 15104
rect 116552 15480 116610 15492
rect 116552 15104 116564 15480
rect 116598 15104 116610 15480
rect 116552 15092 116610 15104
rect 119108 13334 119170 13346
rect 119108 12358 119120 13334
rect 119154 12358 119170 13334
rect 119108 12346 119170 12358
rect 119200 13334 119266 13346
rect 119200 12358 119216 13334
rect 119250 12358 119266 13334
rect 119200 12346 119266 12358
rect 119296 13334 119358 13346
rect 119296 12358 119312 13334
rect 119346 12358 119358 13334
rect 119846 13334 119908 13346
rect 119296 12346 119358 12358
rect 119846 12358 119858 13334
rect 119892 12358 119908 13334
rect 119846 12346 119908 12358
rect 119938 13334 120000 13346
rect 119938 12358 119954 13334
rect 119988 12358 120000 13334
rect 119938 12346 120000 12358
rect 120056 13334 120118 13346
rect 120056 12358 120068 13334
rect 120102 12358 120118 13334
rect 120056 12346 120118 12358
rect 120148 13334 120210 13346
rect 120148 12358 120164 13334
rect 120198 12358 120210 13334
rect 120148 12346 120210 12358
rect 120266 13334 120328 13346
rect 120266 12358 120278 13334
rect 120312 12358 120328 13334
rect 120266 12346 120328 12358
rect 120358 13334 120420 13346
rect 120358 12358 120374 13334
rect 120408 12358 120420 13334
rect 120358 12346 120420 12358
rect 120476 13334 120538 13346
rect 120476 12358 120488 13334
rect 120522 12358 120538 13334
rect 120476 12346 120538 12358
rect 120568 13334 120630 13346
rect 120568 12358 120584 13334
rect 120618 12358 120630 13334
rect 120568 12346 120630 12358
rect 120686 13334 120748 13346
rect 120686 12358 120698 13334
rect 120732 12358 120748 13334
rect 120686 12346 120748 12358
rect 120778 13334 120840 13346
rect 120778 12358 120794 13334
rect 120828 12358 120840 13334
rect 120778 12346 120840 12358
rect 120896 13334 120958 13346
rect 120896 12358 120908 13334
rect 120942 12358 120958 13334
rect 120896 12346 120958 12358
rect 120988 13334 121050 13346
rect 120988 12358 121004 13334
rect 121038 12358 121050 13334
rect 120988 12346 121050 12358
rect 121106 13334 121168 13346
rect 121106 12358 121118 13334
rect 121152 12358 121168 13334
rect 121106 12346 121168 12358
rect 121198 13334 121260 13346
rect 121198 12358 121214 13334
rect 121248 12358 121260 13334
rect 121198 12346 121260 12358
rect 121316 13334 121378 13346
rect 121316 12358 121328 13334
rect 121362 12358 121378 13334
rect 121316 12346 121378 12358
rect 121408 13334 121470 13346
rect 121408 12358 121424 13334
rect 121458 12358 121470 13334
rect 121408 12346 121470 12358
rect 122020 13334 122082 13346
rect 122020 12358 122032 13334
rect 122066 12358 122082 13334
rect 122020 12346 122082 12358
rect 122112 13334 122174 13346
rect 122112 12358 122128 13334
rect 122162 12358 122174 13334
rect 122112 12346 122174 12358
rect 122230 13334 122292 13346
rect 122230 12358 122242 13334
rect 122276 12358 122292 13334
rect 122230 12346 122292 12358
rect 122322 13334 122384 13346
rect 122322 12358 122338 13334
rect 122372 12358 122384 13334
rect 122322 12346 122384 12358
rect 122440 13334 122502 13346
rect 122440 12358 122452 13334
rect 122486 12358 122502 13334
rect 122440 12346 122502 12358
rect 122532 13334 122594 13346
rect 122532 12358 122548 13334
rect 122582 12358 122594 13334
rect 122532 12346 122594 12358
rect 122650 13334 122712 13346
rect 122650 12358 122662 13334
rect 122696 12358 122712 13334
rect 122650 12346 122712 12358
rect 122742 13334 122804 13346
rect 122742 12358 122758 13334
rect 122792 12358 122804 13334
rect 122742 12346 122804 12358
rect 122860 13334 122922 13346
rect 122860 12358 122872 13334
rect 122906 12358 122922 13334
rect 122860 12346 122922 12358
rect 122952 13334 123014 13346
rect 122952 12358 122968 13334
rect 123002 12358 123014 13334
rect 122952 12346 123014 12358
rect 123070 13334 123132 13346
rect 123070 12358 123082 13334
rect 123116 12358 123132 13334
rect 123070 12346 123132 12358
rect 123162 13334 123224 13346
rect 123162 12358 123178 13334
rect 123212 12358 123224 13334
rect 123162 12346 123224 12358
rect 123280 13334 123342 13346
rect 123280 12358 123292 13334
rect 123326 12358 123342 13334
rect 123280 12346 123342 12358
rect 123372 13334 123434 13346
rect 123372 12358 123388 13334
rect 123422 12358 123434 13334
rect 123372 12346 123434 12358
rect 123490 13334 123552 13346
rect 123490 12358 123502 13334
rect 123536 12358 123552 13334
rect 123490 12346 123552 12358
rect 123582 13334 123644 13346
rect 123582 12358 123598 13334
rect 123632 12358 123644 13334
rect 123582 12346 123644 12358
rect 123700 13334 123762 13346
rect 123700 12358 123712 13334
rect 123746 12358 123762 13334
rect 123700 12346 123762 12358
rect 123792 13334 123854 13346
rect 123792 12358 123808 13334
rect 123842 12358 123854 13334
rect 123792 12346 123854 12358
rect 123910 13334 123972 13346
rect 123910 12358 123922 13334
rect 123956 12358 123972 13334
rect 123910 12346 123972 12358
rect 124002 13334 124064 13346
rect 124002 12358 124018 13334
rect 124052 12358 124064 13334
rect 124002 12346 124064 12358
rect 124120 13334 124182 13346
rect 124120 12358 124132 13334
rect 124166 12358 124182 13334
rect 124120 12346 124182 12358
rect 124212 13334 124274 13346
rect 124212 12358 124228 13334
rect 124262 12358 124274 13334
rect 124212 12346 124274 12358
rect 124330 13334 124392 13346
rect 124330 12358 124342 13334
rect 124376 12358 124392 13334
rect 124330 12346 124392 12358
rect 124422 13334 124484 13346
rect 124422 12358 124438 13334
rect 124472 12358 124484 13334
rect 124422 12346 124484 12358
rect 124540 13334 124602 13346
rect 124540 12358 124552 13334
rect 124586 12358 124602 13334
rect 124540 12346 124602 12358
rect 124632 13334 124694 13346
rect 124632 12358 124648 13334
rect 124682 12358 124694 13334
rect 124632 12346 124694 12358
rect 124750 13334 124812 13346
rect 124750 12358 124762 13334
rect 124796 12358 124812 13334
rect 124750 12346 124812 12358
rect 124842 13334 124904 13346
rect 124842 12358 124858 13334
rect 124892 12358 124904 13334
rect 124842 12346 124904 12358
rect 124960 13334 125022 13346
rect 124960 12358 124972 13334
rect 125006 12358 125022 13334
rect 124960 12346 125022 12358
rect 125052 13334 125114 13346
rect 125052 12358 125068 13334
rect 125102 12358 125114 13334
rect 125052 12346 125114 12358
rect 125170 13334 125232 13346
rect 125170 12358 125182 13334
rect 125216 12358 125232 13334
rect 125170 12346 125232 12358
rect 125262 13334 125324 13346
rect 125262 12358 125278 13334
rect 125312 12358 125324 13334
rect 125262 12346 125324 12358
rect 125380 13334 125442 13346
rect 125380 12358 125392 13334
rect 125426 12358 125442 13334
rect 125380 12346 125442 12358
rect 125472 13334 125534 13346
rect 125472 12358 125488 13334
rect 125522 12358 125534 13334
rect 125472 12346 125534 12358
rect 125590 13334 125652 13346
rect 125590 12358 125602 13334
rect 125636 12358 125652 13334
rect 125590 12346 125652 12358
rect 125682 13334 125744 13346
rect 125682 12358 125698 13334
rect 125732 12358 125744 13334
rect 125682 12346 125744 12358
rect 122020 12098 122082 12110
rect 122020 11122 122032 12098
rect 122066 11122 122082 12098
rect 122020 11110 122082 11122
rect 122112 12098 122174 12110
rect 122112 11122 122128 12098
rect 122162 11122 122174 12098
rect 122112 11110 122174 11122
rect 122230 12098 122292 12110
rect 122230 11122 122242 12098
rect 122276 11122 122292 12098
rect 122230 11110 122292 11122
rect 122322 12098 122384 12110
rect 122322 11122 122338 12098
rect 122372 11122 122384 12098
rect 122322 11110 122384 11122
rect 122440 12098 122502 12110
rect 122440 11122 122452 12098
rect 122486 11122 122502 12098
rect 122440 11110 122502 11122
rect 122532 12098 122594 12110
rect 122532 11122 122548 12098
rect 122582 11122 122594 12098
rect 122532 11110 122594 11122
rect 122650 12098 122712 12110
rect 122650 11122 122662 12098
rect 122696 11122 122712 12098
rect 122650 11110 122712 11122
rect 122742 12098 122804 12110
rect 122742 11122 122758 12098
rect 122792 11122 122804 12098
rect 122742 11110 122804 11122
rect 122860 12098 122922 12110
rect 122860 11122 122872 12098
rect 122906 11122 122922 12098
rect 122860 11110 122922 11122
rect 122952 12098 123014 12110
rect 122952 11122 122968 12098
rect 123002 11122 123014 12098
rect 122952 11110 123014 11122
rect 123070 12098 123132 12110
rect 123070 11122 123082 12098
rect 123116 11122 123132 12098
rect 123070 11110 123132 11122
rect 123162 12098 123224 12110
rect 123162 11122 123178 12098
rect 123212 11122 123224 12098
rect 123162 11110 123224 11122
rect 123280 12098 123342 12110
rect 123280 11122 123292 12098
rect 123326 11122 123342 12098
rect 123280 11110 123342 11122
rect 123372 12098 123434 12110
rect 123372 11122 123388 12098
rect 123422 11122 123434 12098
rect 123372 11110 123434 11122
rect 123490 12098 123552 12110
rect 123490 11122 123502 12098
rect 123536 11122 123552 12098
rect 123490 11110 123552 11122
rect 123582 12098 123644 12110
rect 123582 11122 123598 12098
rect 123632 11122 123644 12098
rect 123582 11110 123644 11122
rect 123700 12098 123762 12110
rect 123700 11122 123712 12098
rect 123746 11122 123762 12098
rect 123700 11110 123762 11122
rect 123792 12098 123854 12110
rect 123792 11122 123808 12098
rect 123842 11122 123854 12098
rect 123792 11110 123854 11122
rect 123910 12098 123972 12110
rect 123910 11122 123922 12098
rect 123956 11122 123972 12098
rect 123910 11110 123972 11122
rect 124002 12098 124064 12110
rect 124002 11122 124018 12098
rect 124052 11122 124064 12098
rect 124002 11110 124064 11122
rect 124120 12098 124182 12110
rect 124120 11122 124132 12098
rect 124166 11122 124182 12098
rect 124120 11110 124182 11122
rect 124212 12098 124274 12110
rect 124212 11122 124228 12098
rect 124262 11122 124274 12098
rect 124212 11110 124274 11122
rect 124330 12098 124392 12110
rect 124330 11122 124342 12098
rect 124376 11122 124392 12098
rect 124330 11110 124392 11122
rect 124422 12098 124484 12110
rect 124422 11122 124438 12098
rect 124472 11122 124484 12098
rect 124422 11110 124484 11122
rect 124540 12098 124602 12110
rect 124540 11122 124552 12098
rect 124586 11122 124602 12098
rect 124540 11110 124602 11122
rect 124632 12098 124694 12110
rect 124632 11122 124648 12098
rect 124682 11122 124694 12098
rect 124632 11110 124694 11122
rect 124750 12098 124812 12110
rect 124750 11122 124762 12098
rect 124796 11122 124812 12098
rect 124750 11110 124812 11122
rect 124842 12098 124904 12110
rect 124842 11122 124858 12098
rect 124892 11122 124904 12098
rect 124842 11110 124904 11122
rect 124960 12098 125022 12110
rect 124960 11122 124972 12098
rect 125006 11122 125022 12098
rect 124960 11110 125022 11122
rect 125052 12098 125114 12110
rect 125052 11122 125068 12098
rect 125102 11122 125114 12098
rect 125052 11110 125114 11122
rect 125170 12098 125232 12110
rect 125170 11122 125182 12098
rect 125216 11122 125232 12098
rect 125170 11110 125232 11122
rect 125262 12098 125324 12110
rect 125262 11122 125278 12098
rect 125312 11122 125324 12098
rect 125262 11110 125324 11122
rect 125380 12098 125442 12110
rect 125380 11122 125392 12098
rect 125426 11122 125442 12098
rect 125380 11110 125442 11122
rect 125472 12098 125534 12110
rect 125472 11122 125488 12098
rect 125522 11122 125534 12098
rect 125472 11110 125534 11122
rect 125590 12098 125652 12110
rect 125590 11122 125602 12098
rect 125636 11122 125652 12098
rect 125590 11110 125652 11122
rect 125682 12098 125744 12110
rect 125682 11122 125698 12098
rect 125732 11122 125744 12098
rect 125682 11110 125744 11122
<< ndiffc >>
rect 126882 26992 126916 27968
rect 126978 26992 127012 27968
rect 127092 26992 127126 27968
rect 127188 26992 127222 27968
rect 127302 26992 127336 27968
rect 127398 26992 127432 27968
rect 127512 26992 127546 27968
rect 127608 26992 127642 27968
rect 127722 26992 127756 27968
rect 127818 26992 127852 27968
rect 127932 26992 127966 27968
rect 128028 26992 128062 27968
rect 128142 26992 128176 27968
rect 128238 26992 128272 27968
rect 128352 26992 128386 27968
rect 128448 26992 128482 27968
rect 128562 26992 128596 27968
rect 128658 26992 128692 27968
rect 128772 26992 128806 27968
rect 128868 26992 128902 27968
rect 128982 26992 129016 27968
rect 129078 26992 129112 27968
rect 129192 26992 129226 27968
rect 129288 26992 129322 27968
rect 129402 26992 129436 27968
rect 129498 26992 129532 27968
rect 129612 26992 129646 27968
rect 129708 26992 129742 27968
rect 129822 26992 129856 27968
rect 129918 26992 129952 27968
rect 130032 26992 130066 27968
rect 130128 26992 130162 27968
rect 130242 26992 130276 27968
rect 130338 26992 130372 27968
rect 130452 26992 130486 27968
rect 130548 26992 130582 27968
rect 130662 26992 130696 27968
rect 130758 26992 130792 27968
rect 130872 26992 130906 27968
rect 130968 26992 131002 27968
rect 131082 26992 131116 27968
rect 131178 26992 131212 27968
rect 131292 26992 131326 27968
rect 131388 26992 131422 27968
rect 131502 26992 131536 27968
rect 131598 26992 131632 27968
rect 131712 26992 131746 27968
rect 131808 26992 131842 27968
rect 131922 26992 131956 27968
rect 132018 26992 132052 27968
rect 132132 26992 132166 27968
rect 132228 26992 132262 27968
rect 132342 26992 132376 27968
rect 132438 26992 132472 27968
rect 132552 26992 132586 27968
rect 132648 26992 132682 27968
rect 132762 26992 132796 27968
rect 132858 26992 132892 27968
rect 132972 26992 133006 27968
rect 133068 26992 133102 27968
rect 133182 26992 133216 27968
rect 133278 26992 133312 27968
rect 133392 26992 133426 27968
rect 133488 26992 133522 27968
rect 133602 26992 133636 27968
rect 133698 26992 133732 27968
rect 133812 26992 133846 27968
rect 133908 26992 133942 27968
rect 134022 26992 134056 27968
rect 134118 26992 134152 27968
rect 134232 26992 134266 27968
rect 134328 26992 134362 27968
rect 134442 26992 134476 27968
rect 134538 26992 134572 27968
rect 134652 26992 134686 27968
rect 134748 26992 134782 27968
rect 134862 26992 134896 27968
rect 134958 26992 134992 27968
rect 135072 26992 135106 27968
rect 135168 26992 135202 27968
rect 126882 25774 126916 26750
rect 126978 25774 127012 26750
rect 127092 25774 127126 26750
rect 127188 25774 127222 26750
rect 127302 25774 127336 26750
rect 127398 25774 127432 26750
rect 127512 25774 127546 26750
rect 127608 25774 127642 26750
rect 127722 25774 127756 26750
rect 127818 25774 127852 26750
rect 127932 25774 127966 26750
rect 128028 25774 128062 26750
rect 128142 25774 128176 26750
rect 128238 25774 128272 26750
rect 128352 25774 128386 26750
rect 128448 25774 128482 26750
rect 128562 25774 128596 26750
rect 128658 25774 128692 26750
rect 128772 25774 128806 26750
rect 128868 25774 128902 26750
rect 128982 25774 129016 26750
rect 129078 25774 129112 26750
rect 129192 25774 129226 26750
rect 129288 25774 129322 26750
rect 129402 25774 129436 26750
rect 129498 25774 129532 26750
rect 129612 25774 129646 26750
rect 129708 25774 129742 26750
rect 129822 25774 129856 26750
rect 129918 25774 129952 26750
rect 130032 25774 130066 26750
rect 130128 25774 130162 26750
rect 130242 25774 130276 26750
rect 130338 25774 130372 26750
rect 130452 25774 130486 26750
rect 130548 25774 130582 26750
rect 130662 25774 130696 26750
rect 130758 25774 130792 26750
rect 130872 25774 130906 26750
rect 130968 25774 131002 26750
rect 131082 25774 131116 26750
rect 131178 25774 131212 26750
rect 131292 25774 131326 26750
rect 131388 25774 131422 26750
rect 131502 25774 131536 26750
rect 131598 25774 131632 26750
rect 131712 25774 131746 26750
rect 131808 25774 131842 26750
rect 131922 25774 131956 26750
rect 132018 25774 132052 26750
rect 132132 25774 132166 26750
rect 132228 25774 132262 26750
rect 132342 25774 132376 26750
rect 132438 25774 132472 26750
rect 132552 25774 132586 26750
rect 132648 25774 132682 26750
rect 132762 25774 132796 26750
rect 132858 25774 132892 26750
rect 132972 25774 133006 26750
rect 133068 25774 133102 26750
rect 133182 25774 133216 26750
rect 133278 25774 133312 26750
rect 133392 25774 133426 26750
rect 133488 25774 133522 26750
rect 133602 25774 133636 26750
rect 133698 25774 133732 26750
rect 133812 25774 133846 26750
rect 133908 25774 133942 26750
rect 134022 25774 134056 26750
rect 134118 25774 134152 26750
rect 134232 25774 134266 26750
rect 134328 25774 134362 26750
rect 134442 25774 134476 26750
rect 134538 25774 134572 26750
rect 134652 25774 134686 26750
rect 134748 25774 134782 26750
rect 134862 25774 134896 26750
rect 134958 25774 134992 26750
rect 135072 25774 135106 26750
rect 135168 25774 135202 26750
rect 122032 20908 122066 21884
rect 122128 20908 122162 21884
rect 122242 20908 122276 21884
rect 122338 20908 122372 21884
rect 122452 20908 122486 21884
rect 122548 20908 122582 21884
rect 122662 20908 122696 21884
rect 122758 20908 122792 21884
rect 122872 20908 122906 21884
rect 122968 20908 123002 21884
rect 123082 20908 123116 21884
rect 123178 20908 123212 21884
rect 123292 20908 123326 21884
rect 123388 20908 123422 21884
rect 123502 20908 123536 21884
rect 123598 20908 123632 21884
rect 123712 20908 123746 21884
rect 123808 20908 123842 21884
rect 123922 20908 123956 21884
rect 124018 20908 124052 21884
rect 124132 20908 124166 21884
rect 124228 20908 124262 21884
rect 124342 20908 124376 21884
rect 124438 20908 124472 21884
rect 124552 20908 124586 21884
rect 124648 20908 124682 21884
rect 124762 20908 124796 21884
rect 124858 20908 124892 21884
rect 124972 20908 125006 21884
rect 125068 20908 125102 21884
rect 125182 20908 125216 21884
rect 125278 20908 125312 21884
rect 125392 20908 125426 21884
rect 125488 20908 125522 21884
rect 125602 20908 125636 21884
rect 125698 20908 125732 21884
rect 119124 19284 119158 20260
rect 119212 19284 119246 20260
rect 120068 19284 120102 20260
rect 120164 19284 120198 20260
rect 120278 19284 120312 20260
rect 120374 19284 120408 20260
rect 120488 19284 120522 20260
rect 120584 19284 120618 20260
rect 120698 19284 120732 20260
rect 120794 19284 120828 20260
rect 116382 16530 116416 16906
rect 116476 16530 116510 16906
rect 116564 16530 116598 16906
rect 115856 14646 115890 14822
rect 115944 14646 115978 14822
rect 116382 14484 116416 14860
rect 116476 14484 116510 14860
rect 116564 14484 116598 14860
rect 119124 11130 119158 12106
rect 119212 11130 119246 12106
rect 120068 11130 120102 12106
rect 120164 11130 120198 12106
rect 120278 11130 120312 12106
rect 120374 11130 120408 12106
rect 120488 11130 120522 12106
rect 120584 11130 120618 12106
rect 120698 11130 120732 12106
rect 120794 11130 120828 12106
rect 122032 8106 122066 9082
rect 122128 8106 122162 9082
rect 122242 8106 122276 9082
rect 122338 8106 122372 9082
rect 122452 8106 122486 9082
rect 122548 8106 122582 9082
rect 122662 8106 122696 9082
rect 122758 8106 122792 9082
rect 122872 8106 122906 9082
rect 122968 8106 123002 9082
rect 123082 8106 123116 9082
rect 123178 8106 123212 9082
rect 123292 8106 123326 9082
rect 123388 8106 123422 9082
rect 123502 8106 123536 9082
rect 123598 8106 123632 9082
rect 123712 8106 123746 9082
rect 123808 8106 123842 9082
rect 123922 8106 123956 9082
rect 124018 8106 124052 9082
rect 124132 8106 124166 9082
rect 124228 8106 124262 9082
rect 124342 8106 124376 9082
rect 124438 8106 124472 9082
rect 124552 8106 124586 9082
rect 124648 8106 124682 9082
rect 124762 8106 124796 9082
rect 124858 8106 124892 9082
rect 124972 8106 125006 9082
rect 125068 8106 125102 9082
rect 125182 8106 125216 9082
rect 125278 8106 125312 9082
rect 125392 8106 125426 9082
rect 125488 8106 125522 9082
rect 125602 8106 125636 9082
rect 125698 8106 125732 9082
<< pdiffc >>
rect 119120 18056 119154 19032
rect 119216 18056 119250 19032
rect 119312 18056 119346 19032
rect 119858 18056 119892 19032
rect 119954 18056 119988 19032
rect 120068 18056 120102 19032
rect 120164 18056 120198 19032
rect 120278 18056 120312 19032
rect 120374 18056 120408 19032
rect 120488 18056 120522 19032
rect 120584 18056 120618 19032
rect 120698 18056 120732 19032
rect 120794 18056 120828 19032
rect 120908 18056 120942 19032
rect 121004 18056 121038 19032
rect 121118 18056 121152 19032
rect 121214 18056 121248 19032
rect 121328 18056 121362 19032
rect 121424 18056 121458 19032
rect 122032 19292 122066 20268
rect 122128 19292 122162 20268
rect 122242 19292 122276 20268
rect 122338 19292 122372 20268
rect 122452 19292 122486 20268
rect 122548 19292 122582 20268
rect 122662 19292 122696 20268
rect 122758 19292 122792 20268
rect 122872 19292 122906 20268
rect 122968 19292 123002 20268
rect 123082 19292 123116 20268
rect 123178 19292 123212 20268
rect 123292 19292 123326 20268
rect 123388 19292 123422 20268
rect 123502 19292 123536 20268
rect 123598 19292 123632 20268
rect 123712 19292 123746 20268
rect 123808 19292 123842 20268
rect 123922 19292 123956 20268
rect 124018 19292 124052 20268
rect 124132 19292 124166 20268
rect 124228 19292 124262 20268
rect 124342 19292 124376 20268
rect 124438 19292 124472 20268
rect 124552 19292 124586 20268
rect 124648 19292 124682 20268
rect 124762 19292 124796 20268
rect 124858 19292 124892 20268
rect 124972 19292 125006 20268
rect 125068 19292 125102 20268
rect 125182 19292 125216 20268
rect 125278 19292 125312 20268
rect 125392 19292 125426 20268
rect 125488 19292 125522 20268
rect 125602 19292 125636 20268
rect 125698 19292 125732 20268
rect 122032 18056 122066 19032
rect 122128 18056 122162 19032
rect 122242 18056 122276 19032
rect 122338 18056 122372 19032
rect 122452 18056 122486 19032
rect 122548 18056 122582 19032
rect 122662 18056 122696 19032
rect 122758 18056 122792 19032
rect 122872 18056 122906 19032
rect 122968 18056 123002 19032
rect 123082 18056 123116 19032
rect 123178 18056 123212 19032
rect 123292 18056 123326 19032
rect 123388 18056 123422 19032
rect 123502 18056 123536 19032
rect 123598 18056 123632 19032
rect 123712 18056 123746 19032
rect 123808 18056 123842 19032
rect 123922 18056 123956 19032
rect 124018 18056 124052 19032
rect 124132 18056 124166 19032
rect 124228 18056 124262 19032
rect 124342 18056 124376 19032
rect 124438 18056 124472 19032
rect 124552 18056 124586 19032
rect 124648 18056 124682 19032
rect 124762 18056 124796 19032
rect 124858 18056 124892 19032
rect 124972 18056 125006 19032
rect 125068 18056 125102 19032
rect 125182 18056 125216 19032
rect 125278 18056 125312 19032
rect 125392 18056 125426 19032
rect 125488 18056 125522 19032
rect 125602 18056 125636 19032
rect 125698 18056 125732 19032
rect 126882 21764 126916 22740
rect 126978 21764 127012 22740
rect 127092 21764 127126 22740
rect 127188 21764 127222 22740
rect 127302 21764 127336 22740
rect 127398 21764 127432 22740
rect 127512 21764 127546 22740
rect 127608 21764 127642 22740
rect 127722 21764 127756 22740
rect 127818 21764 127852 22740
rect 127932 21764 127966 22740
rect 128028 21764 128062 22740
rect 128142 21764 128176 22740
rect 128238 21764 128272 22740
rect 128352 21764 128386 22740
rect 128448 21764 128482 22740
rect 128562 21764 128596 22740
rect 128658 21764 128692 22740
rect 128772 21764 128806 22740
rect 128868 21764 128902 22740
rect 128982 21764 129016 22740
rect 129078 21764 129112 22740
rect 129192 21764 129226 22740
rect 129288 21764 129322 22740
rect 129402 21764 129436 22740
rect 129498 21764 129532 22740
rect 129612 21764 129646 22740
rect 129708 21764 129742 22740
rect 129822 21764 129856 22740
rect 129918 21764 129952 22740
rect 130032 21764 130066 22740
rect 130128 21764 130162 22740
rect 130242 21764 130276 22740
rect 130338 21764 130372 22740
rect 130452 21764 130486 22740
rect 130548 21764 130582 22740
rect 130662 21764 130696 22740
rect 130758 21764 130792 22740
rect 130872 21764 130906 22740
rect 130968 21764 131002 22740
rect 131082 21764 131116 22740
rect 131178 21764 131212 22740
rect 131292 21764 131326 22740
rect 131388 21764 131422 22740
rect 131502 21764 131536 22740
rect 131598 21764 131632 22740
rect 131712 21764 131746 22740
rect 131808 21764 131842 22740
rect 131922 21764 131956 22740
rect 132018 21764 132052 22740
rect 132132 21764 132166 22740
rect 132228 21764 132262 22740
rect 132342 21764 132376 22740
rect 132438 21764 132472 22740
rect 132552 21764 132586 22740
rect 132648 21764 132682 22740
rect 132762 21764 132796 22740
rect 132858 21764 132892 22740
rect 132972 21764 133006 22740
rect 133068 21764 133102 22740
rect 133182 21764 133216 22740
rect 133278 21764 133312 22740
rect 133392 21764 133426 22740
rect 133488 21764 133522 22740
rect 133602 21764 133636 22740
rect 133698 21764 133732 22740
rect 133812 21764 133846 22740
rect 133908 21764 133942 22740
rect 134022 21764 134056 22740
rect 134118 21764 134152 22740
rect 134232 21764 134266 22740
rect 134328 21764 134362 22740
rect 134442 21764 134476 22740
rect 134538 21764 134572 22740
rect 134652 21764 134686 22740
rect 134748 21764 134782 22740
rect 134862 21764 134896 22740
rect 134958 21764 134992 22740
rect 135072 21764 135106 22740
rect 135168 21764 135202 22740
rect 126882 20528 126916 21504
rect 126978 20528 127012 21504
rect 127092 20528 127126 21504
rect 127188 20528 127222 21504
rect 127302 20528 127336 21504
rect 127398 20528 127432 21504
rect 127512 20528 127546 21504
rect 127608 20528 127642 21504
rect 127722 20528 127756 21504
rect 127818 20528 127852 21504
rect 127932 20528 127966 21504
rect 128028 20528 128062 21504
rect 128142 20528 128176 21504
rect 128238 20528 128272 21504
rect 128352 20528 128386 21504
rect 128448 20528 128482 21504
rect 128562 20528 128596 21504
rect 128658 20528 128692 21504
rect 128772 20528 128806 21504
rect 128868 20528 128902 21504
rect 128982 20528 129016 21504
rect 129078 20528 129112 21504
rect 129192 20528 129226 21504
rect 129288 20528 129322 21504
rect 129402 20528 129436 21504
rect 129498 20528 129532 21504
rect 129612 20528 129646 21504
rect 129708 20528 129742 21504
rect 129822 20528 129856 21504
rect 129918 20528 129952 21504
rect 130032 20528 130066 21504
rect 130128 20528 130162 21504
rect 130242 20528 130276 21504
rect 130338 20528 130372 21504
rect 130452 20528 130486 21504
rect 130548 20528 130582 21504
rect 130662 20528 130696 21504
rect 130758 20528 130792 21504
rect 130872 20528 130906 21504
rect 130968 20528 131002 21504
rect 131082 20528 131116 21504
rect 131178 20528 131212 21504
rect 131292 20528 131326 21504
rect 131388 20528 131422 21504
rect 131502 20528 131536 21504
rect 131598 20528 131632 21504
rect 131712 20528 131746 21504
rect 131808 20528 131842 21504
rect 131922 20528 131956 21504
rect 132018 20528 132052 21504
rect 132132 20528 132166 21504
rect 132228 20528 132262 21504
rect 132342 20528 132376 21504
rect 132438 20528 132472 21504
rect 132552 20528 132586 21504
rect 132648 20528 132682 21504
rect 132762 20528 132796 21504
rect 132858 20528 132892 21504
rect 132972 20528 133006 21504
rect 133068 20528 133102 21504
rect 133182 20528 133216 21504
rect 133278 20528 133312 21504
rect 133392 20528 133426 21504
rect 133488 20528 133522 21504
rect 133602 20528 133636 21504
rect 133698 20528 133732 21504
rect 133812 20528 133846 21504
rect 133908 20528 133942 21504
rect 134022 20528 134056 21504
rect 134118 20528 134152 21504
rect 134232 20528 134266 21504
rect 134328 20528 134362 21504
rect 134442 20528 134476 21504
rect 134538 20528 134572 21504
rect 134652 20528 134686 21504
rect 134748 20528 134782 21504
rect 134862 20528 134896 21504
rect 134958 20528 134992 21504
rect 135072 20528 135106 21504
rect 135168 20528 135202 21504
rect 126882 19292 126916 20268
rect 126978 19292 127012 20268
rect 127092 19292 127126 20268
rect 127188 19292 127222 20268
rect 127302 19292 127336 20268
rect 127398 19292 127432 20268
rect 127512 19292 127546 20268
rect 127608 19292 127642 20268
rect 127722 19292 127756 20268
rect 127818 19292 127852 20268
rect 127932 19292 127966 20268
rect 128028 19292 128062 20268
rect 128142 19292 128176 20268
rect 128238 19292 128272 20268
rect 128352 19292 128386 20268
rect 128448 19292 128482 20268
rect 128562 19292 128596 20268
rect 128658 19292 128692 20268
rect 128772 19292 128806 20268
rect 128868 19292 128902 20268
rect 128982 19292 129016 20268
rect 129078 19292 129112 20268
rect 129192 19292 129226 20268
rect 129288 19292 129322 20268
rect 129402 19292 129436 20268
rect 129498 19292 129532 20268
rect 129612 19292 129646 20268
rect 129708 19292 129742 20268
rect 129822 19292 129856 20268
rect 129918 19292 129952 20268
rect 130032 19292 130066 20268
rect 130128 19292 130162 20268
rect 130242 19292 130276 20268
rect 130338 19292 130372 20268
rect 130452 19292 130486 20268
rect 130548 19292 130582 20268
rect 130662 19292 130696 20268
rect 130758 19292 130792 20268
rect 130872 19292 130906 20268
rect 130968 19292 131002 20268
rect 131082 19292 131116 20268
rect 131178 19292 131212 20268
rect 131292 19292 131326 20268
rect 131388 19292 131422 20268
rect 131502 19292 131536 20268
rect 131598 19292 131632 20268
rect 131712 19292 131746 20268
rect 131808 19292 131842 20268
rect 131922 19292 131956 20268
rect 132018 19292 132052 20268
rect 132132 19292 132166 20268
rect 132228 19292 132262 20268
rect 132342 19292 132376 20268
rect 132438 19292 132472 20268
rect 132552 19292 132586 20268
rect 132648 19292 132682 20268
rect 132762 19292 132796 20268
rect 132858 19292 132892 20268
rect 132972 19292 133006 20268
rect 133068 19292 133102 20268
rect 133182 19292 133216 20268
rect 133278 19292 133312 20268
rect 133392 19292 133426 20268
rect 133488 19292 133522 20268
rect 133602 19292 133636 20268
rect 133698 19292 133732 20268
rect 133812 19292 133846 20268
rect 133908 19292 133942 20268
rect 134022 19292 134056 20268
rect 134118 19292 134152 20268
rect 134232 19292 134266 20268
rect 134328 19292 134362 20268
rect 134442 19292 134476 20268
rect 134538 19292 134572 20268
rect 134652 19292 134686 20268
rect 134748 19292 134782 20268
rect 134862 19292 134896 20268
rect 134958 19292 134992 20268
rect 135072 19292 135106 20268
rect 135168 19292 135202 20268
rect 126882 18056 126916 19032
rect 126978 18056 127012 19032
rect 127092 18056 127126 19032
rect 127188 18056 127222 19032
rect 127302 18056 127336 19032
rect 127398 18056 127432 19032
rect 127512 18056 127546 19032
rect 127608 18056 127642 19032
rect 127722 18056 127756 19032
rect 127818 18056 127852 19032
rect 127932 18056 127966 19032
rect 128028 18056 128062 19032
rect 128142 18056 128176 19032
rect 128238 18056 128272 19032
rect 128352 18056 128386 19032
rect 128448 18056 128482 19032
rect 128562 18056 128596 19032
rect 128658 18056 128692 19032
rect 128772 18056 128806 19032
rect 128868 18056 128902 19032
rect 128982 18056 129016 19032
rect 129078 18056 129112 19032
rect 129192 18056 129226 19032
rect 129288 18056 129322 19032
rect 129402 18056 129436 19032
rect 129498 18056 129532 19032
rect 129612 18056 129646 19032
rect 129708 18056 129742 19032
rect 129822 18056 129856 19032
rect 129918 18056 129952 19032
rect 130032 18056 130066 19032
rect 130128 18056 130162 19032
rect 130242 18056 130276 19032
rect 130338 18056 130372 19032
rect 130452 18056 130486 19032
rect 130548 18056 130582 19032
rect 130662 18056 130696 19032
rect 130758 18056 130792 19032
rect 130872 18056 130906 19032
rect 130968 18056 131002 19032
rect 131082 18056 131116 19032
rect 131178 18056 131212 19032
rect 131292 18056 131326 19032
rect 131388 18056 131422 19032
rect 131502 18056 131536 19032
rect 131598 18056 131632 19032
rect 131712 18056 131746 19032
rect 131808 18056 131842 19032
rect 131922 18056 131956 19032
rect 132018 18056 132052 19032
rect 132132 18056 132166 19032
rect 132228 18056 132262 19032
rect 132342 18056 132376 19032
rect 132438 18056 132472 19032
rect 132552 18056 132586 19032
rect 132648 18056 132682 19032
rect 132762 18056 132796 19032
rect 132858 18056 132892 19032
rect 132972 18056 133006 19032
rect 133068 18056 133102 19032
rect 133182 18056 133216 19032
rect 133278 18056 133312 19032
rect 133392 18056 133426 19032
rect 133488 18056 133522 19032
rect 133602 18056 133636 19032
rect 133698 18056 133732 19032
rect 133812 18056 133846 19032
rect 133908 18056 133942 19032
rect 134022 18056 134056 19032
rect 134118 18056 134152 19032
rect 134232 18056 134266 19032
rect 134328 18056 134362 19032
rect 134442 18056 134476 19032
rect 134538 18056 134572 19032
rect 134652 18056 134686 19032
rect 134748 18056 134782 19032
rect 134862 18056 134896 19032
rect 134958 18056 134992 19032
rect 135072 18056 135106 19032
rect 135168 18056 135202 19032
rect 116382 15910 116416 16286
rect 116476 15910 116510 16286
rect 116564 15910 116598 16286
rect 115856 15102 115890 15478
rect 115944 15102 115978 15478
rect 116382 15104 116416 15480
rect 116476 15104 116510 15480
rect 116564 15104 116598 15480
rect 119120 12358 119154 13334
rect 119216 12358 119250 13334
rect 119312 12358 119346 13334
rect 119858 12358 119892 13334
rect 119954 12358 119988 13334
rect 120068 12358 120102 13334
rect 120164 12358 120198 13334
rect 120278 12358 120312 13334
rect 120374 12358 120408 13334
rect 120488 12358 120522 13334
rect 120584 12358 120618 13334
rect 120698 12358 120732 13334
rect 120794 12358 120828 13334
rect 120908 12358 120942 13334
rect 121004 12358 121038 13334
rect 121118 12358 121152 13334
rect 121214 12358 121248 13334
rect 121328 12358 121362 13334
rect 121424 12358 121458 13334
rect 122032 12358 122066 13334
rect 122128 12358 122162 13334
rect 122242 12358 122276 13334
rect 122338 12358 122372 13334
rect 122452 12358 122486 13334
rect 122548 12358 122582 13334
rect 122662 12358 122696 13334
rect 122758 12358 122792 13334
rect 122872 12358 122906 13334
rect 122968 12358 123002 13334
rect 123082 12358 123116 13334
rect 123178 12358 123212 13334
rect 123292 12358 123326 13334
rect 123388 12358 123422 13334
rect 123502 12358 123536 13334
rect 123598 12358 123632 13334
rect 123712 12358 123746 13334
rect 123808 12358 123842 13334
rect 123922 12358 123956 13334
rect 124018 12358 124052 13334
rect 124132 12358 124166 13334
rect 124228 12358 124262 13334
rect 124342 12358 124376 13334
rect 124438 12358 124472 13334
rect 124552 12358 124586 13334
rect 124648 12358 124682 13334
rect 124762 12358 124796 13334
rect 124858 12358 124892 13334
rect 124972 12358 125006 13334
rect 125068 12358 125102 13334
rect 125182 12358 125216 13334
rect 125278 12358 125312 13334
rect 125392 12358 125426 13334
rect 125488 12358 125522 13334
rect 125602 12358 125636 13334
rect 125698 12358 125732 13334
rect 122032 11122 122066 12098
rect 122128 11122 122162 12098
rect 122242 11122 122276 12098
rect 122338 11122 122372 12098
rect 122452 11122 122486 12098
rect 122548 11122 122582 12098
rect 122662 11122 122696 12098
rect 122758 11122 122792 12098
rect 122872 11122 122906 12098
rect 122968 11122 123002 12098
rect 123082 11122 123116 12098
rect 123178 11122 123212 12098
rect 123292 11122 123326 12098
rect 123388 11122 123422 12098
rect 123502 11122 123536 12098
rect 123598 11122 123632 12098
rect 123712 11122 123746 12098
rect 123808 11122 123842 12098
rect 123922 11122 123956 12098
rect 124018 11122 124052 12098
rect 124132 11122 124166 12098
rect 124228 11122 124262 12098
rect 124342 11122 124376 12098
rect 124438 11122 124472 12098
rect 124552 11122 124586 12098
rect 124648 11122 124682 12098
rect 124762 11122 124796 12098
rect 124858 11122 124892 12098
rect 124972 11122 125006 12098
rect 125068 11122 125102 12098
rect 125182 11122 125216 12098
rect 125278 11122 125312 12098
rect 125392 11122 125426 12098
rect 125488 11122 125522 12098
rect 125602 11122 125636 12098
rect 125698 11122 125732 12098
<< psubdiffcont >>
rect 126786 28200 135210 28234
rect 126642 25706 126676 28078
rect 135362 25694 135396 28106
rect 126798 25524 135168 25558
rect 122018 22028 125742 22062
rect 121886 20892 121920 21912
rect 125814 20894 125848 21936
rect 121978 20740 125698 20774
rect 119538 19458 119744 20150
rect 116190 16616 116284 16830
rect 115726 14668 115790 14810
rect 116190 14560 116284 14774
rect 119538 11240 119744 11932
rect 121978 9216 125698 9250
rect 121886 8078 121920 9098
rect 125814 8054 125848 9096
rect 122018 7928 125742 7962
<< nsubdiffcont >>
rect 126896 22928 135218 22962
rect 122052 20468 125754 20502
rect 119462 18256 119668 18948
rect 121922 17958 121956 20426
rect 125836 17996 125870 20284
rect 126670 17978 126704 22776
rect 135300 18040 135334 22758
rect 122024 17836 125796 17870
rect 126860 17820 135182 17854
rect 116208 15998 116284 16204
rect 115750 15322 115790 15438
rect 116208 15186 116284 15392
rect 122024 13520 125796 13554
rect 119462 12442 119668 13134
rect 121922 10964 121956 13432
rect 125836 11106 125870 13394
rect 122052 10888 125754 10922
<< poly >>
rect 126914 28052 127030 28068
rect 126914 28018 126930 28052
rect 127014 28018 127030 28052
rect 126914 28002 127030 28018
rect 127334 28052 127450 28068
rect 127334 28018 127350 28052
rect 127434 28018 127450 28052
rect 126932 27980 126962 28002
rect 127142 27980 127172 28006
rect 127334 28002 127450 28018
rect 127754 28052 127870 28068
rect 127754 28018 127770 28052
rect 127854 28018 127870 28052
rect 127352 27980 127382 28002
rect 127562 27980 127592 28006
rect 127754 28002 127870 28018
rect 128174 28052 128290 28068
rect 128174 28018 128190 28052
rect 128274 28018 128290 28052
rect 127772 27980 127802 28002
rect 127982 27980 128012 28006
rect 128174 28002 128290 28018
rect 128594 28052 128710 28068
rect 128594 28018 128610 28052
rect 128694 28018 128710 28052
rect 128192 27980 128222 28002
rect 128402 27980 128432 28006
rect 128594 28002 128710 28018
rect 129014 28052 129130 28068
rect 129014 28018 129030 28052
rect 129114 28018 129130 28052
rect 128612 27980 128642 28002
rect 128822 27980 128852 28006
rect 129014 28002 129130 28018
rect 129434 28052 129550 28068
rect 129434 28018 129450 28052
rect 129534 28018 129550 28052
rect 129032 27980 129062 28002
rect 129242 27980 129272 28006
rect 129434 28002 129550 28018
rect 129854 28052 129970 28068
rect 129854 28018 129870 28052
rect 129954 28018 129970 28052
rect 129452 27980 129482 28002
rect 129662 27980 129692 28006
rect 129854 28002 129970 28018
rect 130274 28052 130390 28068
rect 130274 28018 130290 28052
rect 130374 28018 130390 28052
rect 129872 27980 129902 28002
rect 130082 27980 130112 28006
rect 130274 28002 130390 28018
rect 130694 28052 130810 28068
rect 130694 28018 130710 28052
rect 130794 28018 130810 28052
rect 130292 27980 130322 28002
rect 130502 27980 130532 28006
rect 130694 28002 130810 28018
rect 131114 28052 131230 28068
rect 131114 28018 131130 28052
rect 131214 28018 131230 28052
rect 130712 27980 130742 28002
rect 130922 27980 130952 28006
rect 131114 28002 131230 28018
rect 131534 28052 131650 28068
rect 131534 28018 131550 28052
rect 131634 28018 131650 28052
rect 131132 27980 131162 28002
rect 131342 27980 131372 28006
rect 131534 28002 131650 28018
rect 131954 28052 132070 28068
rect 131954 28018 131970 28052
rect 132054 28018 132070 28052
rect 131552 27980 131582 28002
rect 131762 27980 131792 28006
rect 131954 28002 132070 28018
rect 132374 28052 132490 28068
rect 132374 28018 132390 28052
rect 132474 28018 132490 28052
rect 131972 27980 132002 28002
rect 132182 27980 132212 28006
rect 132374 28002 132490 28018
rect 132794 28052 132910 28068
rect 132794 28018 132810 28052
rect 132894 28018 132910 28052
rect 132392 27980 132422 28002
rect 132602 27980 132632 28006
rect 132794 28002 132910 28018
rect 133214 28052 133330 28068
rect 133214 28018 133230 28052
rect 133314 28018 133330 28052
rect 132812 27980 132842 28002
rect 133022 27980 133052 28006
rect 133214 28002 133330 28018
rect 133634 28052 133750 28068
rect 133634 28018 133650 28052
rect 133734 28018 133750 28052
rect 133232 27980 133262 28002
rect 133442 27980 133472 28006
rect 133634 28002 133750 28018
rect 134054 28052 134170 28068
rect 134054 28018 134070 28052
rect 134154 28018 134170 28052
rect 133652 27980 133682 28002
rect 133862 27980 133892 28006
rect 134054 28002 134170 28018
rect 134474 28052 134590 28068
rect 134474 28018 134490 28052
rect 134574 28018 134590 28052
rect 134072 27980 134102 28002
rect 134282 27980 134312 28006
rect 134474 28002 134590 28018
rect 134894 28052 135010 28068
rect 134894 28018 134910 28052
rect 134994 28018 135010 28052
rect 134492 27980 134522 28002
rect 134702 27980 134732 28006
rect 134894 28002 135010 28018
rect 134912 27980 134942 28002
rect 135122 27980 135152 28006
rect 126932 26954 126962 26980
rect 127142 26958 127172 26980
rect 127124 26942 127190 26958
rect 127352 26954 127382 26980
rect 127562 26958 127592 26980
rect 127124 26800 127140 26942
rect 127174 26800 127190 26942
rect 126932 26762 126962 26788
rect 127124 26784 127190 26800
rect 127544 26942 127610 26958
rect 127772 26954 127802 26980
rect 127982 26958 128012 26980
rect 127544 26800 127560 26942
rect 127594 26800 127610 26942
rect 127142 26762 127172 26784
rect 127352 26762 127382 26788
rect 127544 26784 127610 26800
rect 127964 26942 128030 26958
rect 128192 26954 128222 26980
rect 128402 26958 128432 26980
rect 127964 26800 127980 26942
rect 128014 26800 128030 26942
rect 127562 26762 127592 26784
rect 127772 26762 127802 26788
rect 127964 26784 128030 26800
rect 128384 26942 128450 26958
rect 128612 26954 128642 26980
rect 128822 26958 128852 26980
rect 128384 26800 128400 26942
rect 128434 26800 128450 26942
rect 127982 26762 128012 26784
rect 128192 26762 128222 26788
rect 128384 26784 128450 26800
rect 128804 26942 128870 26958
rect 129032 26954 129062 26980
rect 129242 26958 129272 26980
rect 128804 26800 128820 26942
rect 128854 26800 128870 26942
rect 128402 26762 128432 26784
rect 128612 26762 128642 26788
rect 128804 26784 128870 26800
rect 129224 26942 129290 26958
rect 129452 26954 129482 26980
rect 129662 26958 129692 26980
rect 129224 26800 129240 26942
rect 129274 26800 129290 26942
rect 128822 26762 128852 26784
rect 129032 26762 129062 26788
rect 129224 26784 129290 26800
rect 129644 26942 129710 26958
rect 129872 26954 129902 26980
rect 130082 26958 130112 26980
rect 129644 26800 129660 26942
rect 129694 26800 129710 26942
rect 129242 26762 129272 26784
rect 129452 26762 129482 26788
rect 129644 26784 129710 26800
rect 130064 26942 130130 26958
rect 130292 26954 130322 26980
rect 130502 26958 130532 26980
rect 130064 26800 130080 26942
rect 130114 26800 130130 26942
rect 129662 26762 129692 26784
rect 129872 26762 129902 26788
rect 130064 26784 130130 26800
rect 130484 26942 130550 26958
rect 130712 26954 130742 26980
rect 130922 26958 130952 26980
rect 130484 26800 130500 26942
rect 130534 26800 130550 26942
rect 130082 26762 130112 26784
rect 130292 26762 130322 26788
rect 130484 26784 130550 26800
rect 130904 26942 130970 26958
rect 131132 26954 131162 26980
rect 131342 26958 131372 26980
rect 130904 26800 130920 26942
rect 130954 26800 130970 26942
rect 130502 26762 130532 26784
rect 130712 26762 130742 26788
rect 130904 26784 130970 26800
rect 131324 26942 131390 26958
rect 131552 26954 131582 26980
rect 131762 26958 131792 26980
rect 131324 26800 131340 26942
rect 131374 26800 131390 26942
rect 130922 26762 130952 26784
rect 131132 26762 131162 26788
rect 131324 26784 131390 26800
rect 131744 26942 131810 26958
rect 131972 26954 132002 26980
rect 132182 26958 132212 26980
rect 131744 26800 131760 26942
rect 131794 26800 131810 26942
rect 131342 26762 131372 26784
rect 131552 26762 131582 26788
rect 131744 26784 131810 26800
rect 132164 26942 132230 26958
rect 132392 26954 132422 26980
rect 132602 26958 132632 26980
rect 132164 26800 132180 26942
rect 132214 26800 132230 26942
rect 131762 26762 131792 26784
rect 131972 26762 132002 26788
rect 132164 26784 132230 26800
rect 132584 26942 132650 26958
rect 132812 26954 132842 26980
rect 133022 26958 133052 26980
rect 132584 26800 132600 26942
rect 132634 26800 132650 26942
rect 132182 26762 132212 26784
rect 132392 26762 132422 26788
rect 132584 26784 132650 26800
rect 133004 26942 133070 26958
rect 133232 26954 133262 26980
rect 133442 26958 133472 26980
rect 133004 26800 133020 26942
rect 133054 26800 133070 26942
rect 132602 26762 132632 26784
rect 132812 26762 132842 26788
rect 133004 26784 133070 26800
rect 133424 26942 133490 26958
rect 133652 26954 133682 26980
rect 133862 26958 133892 26980
rect 133424 26800 133440 26942
rect 133474 26800 133490 26942
rect 133022 26762 133052 26784
rect 133232 26762 133262 26788
rect 133424 26784 133490 26800
rect 133844 26942 133910 26958
rect 134072 26954 134102 26980
rect 134282 26958 134312 26980
rect 133844 26800 133860 26942
rect 133894 26800 133910 26942
rect 133442 26762 133472 26784
rect 133652 26762 133682 26788
rect 133844 26784 133910 26800
rect 134264 26942 134330 26958
rect 134492 26954 134522 26980
rect 134702 26958 134732 26980
rect 134264 26800 134280 26942
rect 134314 26800 134330 26942
rect 133862 26762 133892 26784
rect 134072 26762 134102 26788
rect 134264 26784 134330 26800
rect 134684 26942 134750 26958
rect 134912 26954 134942 26980
rect 135122 26958 135152 26980
rect 134684 26800 134700 26942
rect 134734 26800 134750 26942
rect 134282 26762 134312 26784
rect 134492 26762 134522 26788
rect 134684 26784 134750 26800
rect 135104 26942 135170 26958
rect 135104 26800 135120 26942
rect 135154 26800 135170 26942
rect 134702 26762 134732 26784
rect 134912 26762 134942 26788
rect 135104 26784 135170 26800
rect 135122 26762 135152 26784
rect 126932 25740 126962 25762
rect 126914 25724 127030 25740
rect 127142 25736 127172 25762
rect 127352 25740 127382 25762
rect 126914 25690 126930 25724
rect 127014 25690 127030 25724
rect 126914 25674 127030 25690
rect 127334 25724 127450 25740
rect 127562 25736 127592 25762
rect 127772 25740 127802 25762
rect 127334 25690 127350 25724
rect 127434 25690 127450 25724
rect 127334 25674 127450 25690
rect 127754 25724 127870 25740
rect 127982 25736 128012 25762
rect 128192 25740 128222 25762
rect 127754 25690 127770 25724
rect 127854 25690 127870 25724
rect 127754 25674 127870 25690
rect 128174 25724 128290 25740
rect 128402 25736 128432 25762
rect 128612 25740 128642 25762
rect 128174 25690 128190 25724
rect 128274 25690 128290 25724
rect 128174 25674 128290 25690
rect 128594 25724 128710 25740
rect 128822 25736 128852 25762
rect 129032 25740 129062 25762
rect 128594 25690 128610 25724
rect 128694 25690 128710 25724
rect 128594 25674 128710 25690
rect 129014 25724 129130 25740
rect 129242 25736 129272 25762
rect 129452 25740 129482 25762
rect 129014 25690 129030 25724
rect 129114 25690 129130 25724
rect 129014 25674 129130 25690
rect 129434 25724 129550 25740
rect 129662 25736 129692 25762
rect 129872 25740 129902 25762
rect 129434 25690 129450 25724
rect 129534 25690 129550 25724
rect 129434 25674 129550 25690
rect 129854 25724 129970 25740
rect 130082 25736 130112 25762
rect 130292 25740 130322 25762
rect 129854 25690 129870 25724
rect 129954 25690 129970 25724
rect 129854 25674 129970 25690
rect 130274 25724 130390 25740
rect 130502 25736 130532 25762
rect 130712 25740 130742 25762
rect 130274 25690 130290 25724
rect 130374 25690 130390 25724
rect 130274 25674 130390 25690
rect 130694 25724 130810 25740
rect 130922 25736 130952 25762
rect 131132 25740 131162 25762
rect 130694 25690 130710 25724
rect 130794 25690 130810 25724
rect 130694 25674 130810 25690
rect 131114 25724 131230 25740
rect 131342 25736 131372 25762
rect 131552 25740 131582 25762
rect 131114 25690 131130 25724
rect 131214 25690 131230 25724
rect 131114 25674 131230 25690
rect 131534 25724 131650 25740
rect 131762 25736 131792 25762
rect 131972 25740 132002 25762
rect 131534 25690 131550 25724
rect 131634 25690 131650 25724
rect 131534 25674 131650 25690
rect 131954 25724 132070 25740
rect 132182 25736 132212 25762
rect 132392 25740 132422 25762
rect 131954 25690 131970 25724
rect 132054 25690 132070 25724
rect 131954 25674 132070 25690
rect 132374 25724 132490 25740
rect 132602 25736 132632 25762
rect 132812 25740 132842 25762
rect 132374 25690 132390 25724
rect 132474 25690 132490 25724
rect 132374 25674 132490 25690
rect 132794 25724 132910 25740
rect 133022 25736 133052 25762
rect 133232 25740 133262 25762
rect 132794 25690 132810 25724
rect 132894 25690 132910 25724
rect 132794 25674 132910 25690
rect 133214 25724 133330 25740
rect 133442 25736 133472 25762
rect 133652 25740 133682 25762
rect 133214 25690 133230 25724
rect 133314 25690 133330 25724
rect 133214 25674 133330 25690
rect 133634 25724 133750 25740
rect 133862 25736 133892 25762
rect 134072 25740 134102 25762
rect 133634 25690 133650 25724
rect 133734 25690 133750 25724
rect 133634 25674 133750 25690
rect 134054 25724 134170 25740
rect 134282 25736 134312 25762
rect 134492 25740 134522 25762
rect 134054 25690 134070 25724
rect 134154 25690 134170 25724
rect 134054 25674 134170 25690
rect 134474 25724 134590 25740
rect 134702 25736 134732 25762
rect 134912 25740 134942 25762
rect 134474 25690 134490 25724
rect 134574 25690 134590 25724
rect 134474 25674 134590 25690
rect 134894 25724 135010 25740
rect 135122 25736 135152 25762
rect 134894 25690 134910 25724
rect 134994 25690 135010 25724
rect 134894 25674 135010 25690
rect 126914 22833 127030 22850
rect 126914 22798 126930 22833
rect 126964 22832 127030 22833
rect 127014 22798 127030 22832
rect 126914 22782 127030 22798
rect 127334 22833 127450 22850
rect 127334 22798 127350 22833
rect 127384 22832 127450 22833
rect 127434 22798 127450 22832
rect 127334 22782 127450 22798
rect 127754 22833 127870 22850
rect 127754 22798 127770 22833
rect 127804 22832 127870 22833
rect 127854 22798 127870 22832
rect 127754 22782 127870 22798
rect 128174 22833 128290 22850
rect 128174 22798 128190 22833
rect 128224 22832 128290 22833
rect 128274 22798 128290 22832
rect 128174 22782 128290 22798
rect 128594 22833 128710 22850
rect 128594 22798 128610 22833
rect 128644 22832 128710 22833
rect 128694 22798 128710 22832
rect 128594 22782 128710 22798
rect 129014 22833 129130 22850
rect 129014 22798 129030 22833
rect 129064 22832 129130 22833
rect 129114 22798 129130 22832
rect 129014 22782 129130 22798
rect 129434 22833 129550 22850
rect 129434 22798 129450 22833
rect 129484 22832 129550 22833
rect 129534 22798 129550 22832
rect 129434 22782 129550 22798
rect 129854 22833 129970 22850
rect 129854 22798 129870 22833
rect 129904 22832 129970 22833
rect 129954 22798 129970 22832
rect 129854 22782 129970 22798
rect 130274 22833 130390 22850
rect 130274 22798 130290 22833
rect 130324 22832 130390 22833
rect 130374 22798 130390 22832
rect 130274 22782 130390 22798
rect 130694 22833 130810 22850
rect 130694 22798 130710 22833
rect 130744 22832 130810 22833
rect 130794 22798 130810 22832
rect 130694 22782 130810 22798
rect 131114 22833 131230 22850
rect 131114 22798 131130 22833
rect 131164 22832 131230 22833
rect 131214 22798 131230 22832
rect 131114 22782 131230 22798
rect 131534 22833 131650 22850
rect 131534 22798 131550 22833
rect 131584 22832 131650 22833
rect 131634 22798 131650 22832
rect 131534 22782 131650 22798
rect 131954 22833 132070 22850
rect 131954 22798 131970 22833
rect 132004 22832 132070 22833
rect 132054 22798 132070 22832
rect 131954 22782 132070 22798
rect 132374 22833 132490 22850
rect 132374 22798 132390 22833
rect 132424 22832 132490 22833
rect 132474 22798 132490 22832
rect 132374 22782 132490 22798
rect 132794 22833 132910 22850
rect 132794 22798 132810 22833
rect 132844 22832 132910 22833
rect 132894 22798 132910 22832
rect 132794 22782 132910 22798
rect 133214 22833 133330 22850
rect 133214 22798 133230 22833
rect 133264 22832 133330 22833
rect 133314 22798 133330 22832
rect 133214 22782 133330 22798
rect 133634 22833 133750 22850
rect 133634 22798 133650 22833
rect 133684 22832 133750 22833
rect 133734 22798 133750 22832
rect 133634 22782 133750 22798
rect 134054 22833 134170 22850
rect 134054 22798 134070 22833
rect 134104 22832 134170 22833
rect 134154 22798 134170 22832
rect 134054 22782 134170 22798
rect 134474 22833 134590 22850
rect 134474 22798 134490 22833
rect 134524 22832 134590 22833
rect 134574 22798 134590 22832
rect 134474 22782 134590 22798
rect 134894 22833 135010 22850
rect 134894 22798 134910 22833
rect 134944 22832 135010 22833
rect 134994 22798 135010 22832
rect 134894 22782 135010 22798
rect 122274 21976 122390 21994
rect 122274 21942 122290 21976
rect 122374 21942 122390 21976
rect 122274 21926 122390 21942
rect 122694 21976 122810 21994
rect 122694 21934 122710 21976
rect 122794 21942 122810 21976
rect 122744 21934 122810 21942
rect 122694 21926 122810 21934
rect 123114 21976 123230 21994
rect 123114 21934 123130 21976
rect 123214 21942 123230 21976
rect 123164 21934 123230 21942
rect 123114 21926 123230 21934
rect 123534 21976 123650 21994
rect 123534 21934 123550 21976
rect 123634 21942 123650 21976
rect 123584 21934 123650 21942
rect 123534 21926 123650 21934
rect 123954 21976 124070 21994
rect 123954 21934 123970 21976
rect 124054 21942 124070 21976
rect 124004 21934 124070 21942
rect 123954 21926 124070 21934
rect 124374 21976 124490 21994
rect 124374 21934 124390 21976
rect 124474 21942 124490 21976
rect 124424 21934 124490 21942
rect 124374 21926 124490 21934
rect 124794 21976 124910 21994
rect 124794 21934 124810 21976
rect 124894 21942 124910 21976
rect 124844 21934 124910 21942
rect 124794 21926 124910 21934
rect 125214 21976 125330 21994
rect 125214 21934 125230 21976
rect 125314 21942 125330 21976
rect 125264 21934 125330 21942
rect 125214 21926 125330 21934
rect 125634 21976 125750 21994
rect 125634 21934 125650 21976
rect 125734 21942 125750 21976
rect 125684 21934 125750 21942
rect 125634 21926 125750 21934
rect 122082 21896 122112 21922
rect 122292 21896 122322 21926
rect 122502 21896 122532 21922
rect 122694 21918 122760 21926
rect 122712 21896 122742 21918
rect 122922 21896 122952 21922
rect 123114 21918 123180 21926
rect 123132 21896 123162 21918
rect 123342 21896 123372 21922
rect 123534 21918 123600 21926
rect 123552 21896 123582 21918
rect 123762 21896 123792 21922
rect 123954 21918 124020 21926
rect 123972 21896 124002 21918
rect 124182 21896 124212 21922
rect 124374 21918 124440 21926
rect 124392 21896 124422 21918
rect 124602 21896 124632 21922
rect 124794 21918 124860 21926
rect 124812 21896 124842 21918
rect 125022 21896 125052 21922
rect 125214 21918 125280 21926
rect 125232 21896 125262 21918
rect 125442 21896 125472 21922
rect 125634 21918 125700 21926
rect 125652 21896 125682 21918
rect 122082 20870 122112 20896
rect 122292 20870 122322 20896
rect 122502 20870 122532 20896
rect 122712 20870 122742 20896
rect 122922 20874 122952 20896
rect 122904 20870 122970 20874
rect 123132 20870 123162 20896
rect 123342 20874 123372 20896
rect 123324 20870 123390 20874
rect 123552 20870 123582 20896
rect 123762 20874 123792 20896
rect 123744 20870 123810 20874
rect 123972 20870 124002 20896
rect 124182 20874 124212 20896
rect 124164 20870 124230 20874
rect 124392 20870 124422 20896
rect 124602 20874 124632 20896
rect 124584 20870 124650 20874
rect 124812 20870 124842 20896
rect 125022 20874 125052 20896
rect 125004 20870 125070 20874
rect 125232 20870 125262 20896
rect 125442 20874 125472 20896
rect 125424 20870 125490 20874
rect 125652 20870 125682 20896
rect 122064 20853 122180 20870
rect 122064 20818 122080 20853
rect 122114 20852 122180 20853
rect 122164 20818 122180 20852
rect 122064 20802 122180 20818
rect 122484 20853 122600 20870
rect 122484 20818 122500 20853
rect 122534 20852 122600 20853
rect 122584 20818 122600 20852
rect 122484 20802 122600 20818
rect 122904 20858 123020 20870
rect 122904 20818 122920 20858
rect 122954 20852 123020 20858
rect 123004 20818 123020 20852
rect 122904 20802 123020 20818
rect 123324 20858 123440 20870
rect 123324 20818 123340 20858
rect 123374 20852 123440 20858
rect 123424 20818 123440 20852
rect 123324 20802 123440 20818
rect 123744 20858 123860 20870
rect 123744 20818 123760 20858
rect 123794 20852 123860 20858
rect 123844 20818 123860 20852
rect 123744 20802 123860 20818
rect 124164 20858 124280 20870
rect 124164 20818 124180 20858
rect 124214 20852 124280 20858
rect 124264 20818 124280 20852
rect 124164 20802 124280 20818
rect 124584 20858 124700 20870
rect 124584 20818 124600 20858
rect 124634 20852 124700 20858
rect 124684 20818 124700 20852
rect 124584 20802 124700 20818
rect 125004 20858 125120 20870
rect 125004 20818 125020 20858
rect 125054 20852 125120 20858
rect 125104 20818 125120 20852
rect 125004 20802 125120 20818
rect 125424 20858 125540 20870
rect 125424 20818 125440 20858
rect 125474 20852 125540 20858
rect 125524 20818 125540 20852
rect 125424 20802 125540 20818
rect 120310 20353 120426 20370
rect 120310 20318 120326 20353
rect 120360 20352 120426 20353
rect 120410 20318 120426 20352
rect 120310 20302 120426 20318
rect 120730 20353 120846 20370
rect 120730 20318 120746 20353
rect 120780 20352 120846 20353
rect 120830 20318 120846 20352
rect 120730 20302 120846 20318
rect 119170 20272 119200 20298
rect 120118 20272 120148 20298
rect 120328 20272 120358 20302
rect 120538 20272 120568 20298
rect 120748 20272 120778 20302
rect 119170 19250 119200 19272
rect 120118 19250 120148 19272
rect 119152 19234 119218 19250
rect 119152 19091 119168 19234
rect 119202 19091 119218 19234
rect 119152 19075 119218 19091
rect 120100 19234 120166 19250
rect 120328 19246 120358 19272
rect 120538 19250 120568 19272
rect 120100 19091 120116 19234
rect 120150 19091 120166 19234
rect 120100 19075 120166 19091
rect 120520 19234 120586 19250
rect 120748 19246 120778 19272
rect 120520 19091 120536 19234
rect 120570 19091 120586 19234
rect 120520 19075 120586 19091
rect 120940 19125 121056 19142
rect 120940 19090 120956 19125
rect 120990 19124 121056 19125
rect 121040 19090 121056 19124
rect 119170 19044 119200 19075
rect 119266 19044 119296 19070
rect 119908 19044 119938 19070
rect 120118 19044 120148 19075
rect 120328 19044 120358 19070
rect 120538 19044 120568 19075
rect 120940 19074 121056 19090
rect 121360 19125 121476 19142
rect 121360 19090 121376 19125
rect 121410 19124 121476 19125
rect 121460 19090 121476 19124
rect 121360 19074 121476 19090
rect 120748 19044 120778 19070
rect 120958 19044 120988 19074
rect 121168 19044 121198 19070
rect 121378 19044 121408 19074
rect 119170 18018 119200 18044
rect 119266 18014 119296 18044
rect 119908 18014 119938 18044
rect 120118 18018 120148 18044
rect 120328 18014 120358 18044
rect 120538 18018 120568 18044
rect 120748 18014 120778 18044
rect 120958 18018 120988 18044
rect 121168 18014 121198 18044
rect 121378 18018 121408 18044
rect 119248 17998 119364 18014
rect 119248 17964 119264 17998
rect 119348 17964 119364 17998
rect 119248 17948 119364 17964
rect 119890 17997 120006 18014
rect 119890 17962 119906 17997
rect 119940 17996 120006 17997
rect 119990 17962 120006 17996
rect 119890 17946 120006 17962
rect 120310 17997 120426 18014
rect 120310 17962 120326 17997
rect 120360 17996 120426 17997
rect 120410 17962 120426 17996
rect 120310 17946 120426 17962
rect 120730 17997 120846 18014
rect 120730 17962 120746 17997
rect 120780 17996 120846 17997
rect 120830 17962 120846 17996
rect 120730 17946 120846 17962
rect 121150 17997 121266 18014
rect 121150 17962 121166 17997
rect 121200 17996 121266 17997
rect 121250 17962 121266 17996
rect 121150 17946 121266 17962
rect 122064 20361 122180 20378
rect 122064 20326 122080 20361
rect 122114 20360 122180 20361
rect 122164 20326 122180 20360
rect 122064 20310 122180 20326
rect 122484 20361 122600 20378
rect 122484 20326 122500 20361
rect 122534 20360 122600 20361
rect 122584 20326 122600 20360
rect 122484 20310 122600 20326
rect 122904 20361 123020 20378
rect 122904 20326 122920 20361
rect 122954 20360 123020 20361
rect 123004 20326 123020 20360
rect 122904 20310 123020 20326
rect 123324 20361 123440 20378
rect 123324 20326 123340 20361
rect 123374 20360 123440 20361
rect 123424 20326 123440 20360
rect 123324 20310 123440 20326
rect 123744 20361 123860 20378
rect 123744 20326 123760 20361
rect 123794 20360 123860 20361
rect 123844 20326 123860 20360
rect 123744 20310 123860 20326
rect 124164 20361 124280 20378
rect 124164 20326 124180 20361
rect 124214 20360 124280 20361
rect 124264 20326 124280 20360
rect 124164 20310 124280 20326
rect 124584 20361 124700 20378
rect 124584 20326 124600 20361
rect 124634 20360 124700 20361
rect 124684 20326 124700 20360
rect 124584 20310 124700 20326
rect 125004 20361 125120 20378
rect 125004 20326 125020 20361
rect 125054 20360 125120 20361
rect 125104 20326 125120 20360
rect 125004 20310 125120 20326
rect 125424 20361 125540 20378
rect 125424 20326 125440 20361
rect 125474 20360 125540 20361
rect 125524 20326 125540 20360
rect 125424 20310 125540 20326
rect 122082 20280 122112 20310
rect 122292 20280 122322 20306
rect 122502 20280 122532 20310
rect 122712 20280 122742 20306
rect 122922 20280 122952 20310
rect 123132 20280 123162 20306
rect 123342 20280 123372 20310
rect 123552 20280 123582 20306
rect 123762 20280 123792 20310
rect 123972 20280 124002 20306
rect 124182 20280 124212 20310
rect 124392 20280 124422 20306
rect 124602 20280 124632 20310
rect 124812 20280 124842 20306
rect 125022 20280 125052 20310
rect 125232 20280 125262 20306
rect 125442 20280 125472 20310
rect 125652 20280 125682 20306
rect 122082 19254 122112 19280
rect 122292 19249 122322 19280
rect 122502 19254 122532 19280
rect 122712 19249 122742 19280
rect 122922 19254 122952 19280
rect 123132 19249 123162 19280
rect 123342 19254 123372 19280
rect 123552 19249 123582 19280
rect 123762 19254 123792 19280
rect 123972 19249 124002 19280
rect 124182 19254 124212 19280
rect 124392 19249 124422 19280
rect 124602 19254 124632 19280
rect 124812 19249 124842 19280
rect 125022 19254 125052 19280
rect 125232 19249 125262 19280
rect 125442 19254 125472 19280
rect 125652 19249 125682 19280
rect 122274 19233 122340 19249
rect 122274 19091 122290 19233
rect 122324 19091 122340 19233
rect 122274 19075 122340 19091
rect 122694 19233 122760 19249
rect 122694 19091 122710 19233
rect 122744 19091 122760 19233
rect 122694 19075 122760 19091
rect 123114 19233 123180 19249
rect 123114 19091 123130 19233
rect 123164 19091 123180 19233
rect 123114 19075 123180 19091
rect 123534 19233 123600 19249
rect 123534 19091 123550 19233
rect 123584 19091 123600 19233
rect 123534 19075 123600 19091
rect 123954 19233 124020 19249
rect 123954 19091 123970 19233
rect 124004 19091 124020 19233
rect 123954 19075 124020 19091
rect 124374 19233 124440 19249
rect 124374 19091 124390 19233
rect 124424 19091 124440 19233
rect 124374 19075 124440 19091
rect 124794 19233 124860 19249
rect 124794 19091 124810 19233
rect 124844 19091 124860 19233
rect 124794 19075 124860 19091
rect 125214 19233 125280 19249
rect 125214 19091 125230 19233
rect 125264 19091 125280 19233
rect 125214 19075 125280 19091
rect 125634 19233 125700 19249
rect 125634 19091 125650 19233
rect 125684 19091 125700 19233
rect 125634 19075 125700 19091
rect 122082 19044 122112 19070
rect 122292 19044 122322 19075
rect 122502 19044 122532 19070
rect 122712 19044 122742 19075
rect 122922 19044 122952 19070
rect 123132 19044 123162 19075
rect 123342 19044 123372 19070
rect 123552 19044 123582 19075
rect 123762 19044 123792 19070
rect 123972 19044 124002 19075
rect 124182 19044 124212 19070
rect 124392 19044 124422 19075
rect 124602 19044 124632 19070
rect 124812 19044 124842 19075
rect 125022 19044 125052 19070
rect 125232 19044 125262 19075
rect 125442 19044 125472 19070
rect 125652 19044 125682 19075
rect 122082 18014 122112 18044
rect 122292 18018 122322 18044
rect 122502 18014 122532 18044
rect 122712 18018 122742 18044
rect 122922 18014 122952 18044
rect 123132 18018 123162 18044
rect 123342 18014 123372 18044
rect 123552 18018 123582 18044
rect 123762 18014 123792 18044
rect 123972 18018 124002 18044
rect 124182 18014 124212 18044
rect 124392 18018 124422 18044
rect 124602 18014 124632 18044
rect 124812 18018 124842 18044
rect 125022 18014 125052 18044
rect 125232 18018 125262 18044
rect 125442 18014 125472 18044
rect 125652 18018 125682 18044
rect 122064 17997 122180 18014
rect 122064 17962 122080 17997
rect 122114 17996 122180 17997
rect 122164 17962 122180 17996
rect 122064 17946 122180 17962
rect 122484 17997 122600 18014
rect 122484 17962 122500 17997
rect 122534 17996 122600 17997
rect 122584 17962 122600 17996
rect 122484 17946 122600 17962
rect 122904 17997 123020 18014
rect 122904 17962 122920 17997
rect 122954 17996 123020 17997
rect 123004 17962 123020 17996
rect 122904 17946 123020 17962
rect 123324 17997 123440 18014
rect 123324 17962 123340 17997
rect 123374 17996 123440 17997
rect 123424 17962 123440 17996
rect 123324 17946 123440 17962
rect 123744 17997 123860 18014
rect 123744 17962 123760 17997
rect 123794 17996 123860 17997
rect 123844 17962 123860 17996
rect 123744 17946 123860 17962
rect 124164 17997 124280 18014
rect 124164 17962 124180 17997
rect 124214 17996 124280 17997
rect 124264 17962 124280 17996
rect 124164 17946 124280 17962
rect 124584 17997 124700 18014
rect 124584 17962 124600 17997
rect 124634 17996 124700 17997
rect 124684 17962 124700 17996
rect 124584 17946 124700 17962
rect 125004 17997 125120 18014
rect 125004 17962 125020 17997
rect 125054 17996 125120 17997
rect 125104 17962 125120 17996
rect 125004 17946 125120 17962
rect 125424 17997 125540 18014
rect 125424 17962 125440 17997
rect 125474 17996 125540 17997
rect 125524 17962 125540 17996
rect 126932 22752 126962 22782
rect 127142 22752 127172 22778
rect 127352 22752 127382 22782
rect 127562 22752 127592 22778
rect 127772 22752 127802 22782
rect 127982 22752 128012 22778
rect 128192 22752 128222 22782
rect 128402 22752 128432 22778
rect 128612 22752 128642 22782
rect 128822 22752 128852 22778
rect 129032 22752 129062 22782
rect 129242 22752 129272 22778
rect 129452 22752 129482 22782
rect 129662 22752 129692 22778
rect 129872 22752 129902 22782
rect 130082 22752 130112 22778
rect 130292 22752 130322 22782
rect 130502 22752 130532 22778
rect 130712 22752 130742 22782
rect 130922 22752 130952 22778
rect 131132 22752 131162 22782
rect 131342 22752 131372 22778
rect 131552 22752 131582 22782
rect 131762 22752 131792 22778
rect 131972 22752 132002 22782
rect 132182 22752 132212 22778
rect 132392 22752 132422 22782
rect 132602 22752 132632 22778
rect 132812 22752 132842 22782
rect 133022 22752 133052 22778
rect 133232 22752 133262 22782
rect 133442 22752 133472 22778
rect 133652 22752 133682 22782
rect 133862 22752 133892 22778
rect 134072 22752 134102 22782
rect 134282 22752 134312 22778
rect 134492 22752 134522 22782
rect 134702 22752 134732 22778
rect 134912 22752 134942 22782
rect 135122 22752 135152 22778
rect 126932 21726 126962 21752
rect 127142 21721 127172 21752
rect 127352 21726 127382 21752
rect 127562 21721 127592 21752
rect 127772 21726 127802 21752
rect 127982 21721 128012 21752
rect 128192 21726 128222 21752
rect 128402 21721 128432 21752
rect 128612 21726 128642 21752
rect 128822 21721 128852 21752
rect 129032 21726 129062 21752
rect 129242 21721 129272 21752
rect 129452 21726 129482 21752
rect 129662 21721 129692 21752
rect 129872 21726 129902 21752
rect 130082 21721 130112 21752
rect 130292 21726 130322 21752
rect 130502 21721 130532 21752
rect 130712 21726 130742 21752
rect 130922 21721 130952 21752
rect 131132 21726 131162 21752
rect 131342 21721 131372 21752
rect 131552 21726 131582 21752
rect 131762 21721 131792 21752
rect 131972 21726 132002 21752
rect 132182 21721 132212 21752
rect 132392 21726 132422 21752
rect 132602 21721 132632 21752
rect 132812 21726 132842 21752
rect 133022 21721 133052 21752
rect 133232 21726 133262 21752
rect 133442 21721 133472 21752
rect 133652 21726 133682 21752
rect 133862 21721 133892 21752
rect 134072 21726 134102 21752
rect 134282 21721 134312 21752
rect 134492 21726 134522 21752
rect 134702 21721 134732 21752
rect 134912 21726 134942 21752
rect 135122 21721 135152 21752
rect 127124 21705 127190 21721
rect 127124 21563 127140 21705
rect 127174 21563 127190 21705
rect 127124 21547 127190 21563
rect 127544 21705 127610 21721
rect 127544 21563 127560 21705
rect 127594 21563 127610 21705
rect 127544 21547 127610 21563
rect 127964 21705 128030 21721
rect 127964 21563 127980 21705
rect 128014 21563 128030 21705
rect 127964 21547 128030 21563
rect 128384 21705 128450 21721
rect 128384 21563 128400 21705
rect 128434 21563 128450 21705
rect 128384 21547 128450 21563
rect 128804 21705 128870 21721
rect 128804 21563 128820 21705
rect 128854 21563 128870 21705
rect 128804 21547 128870 21563
rect 129224 21705 129290 21721
rect 129224 21563 129240 21705
rect 129274 21563 129290 21705
rect 129224 21547 129290 21563
rect 129644 21705 129710 21721
rect 129644 21563 129660 21705
rect 129694 21563 129710 21705
rect 129644 21547 129710 21563
rect 130064 21705 130130 21721
rect 130064 21563 130080 21705
rect 130114 21563 130130 21705
rect 130064 21547 130130 21563
rect 130484 21705 130550 21721
rect 130484 21563 130500 21705
rect 130534 21563 130550 21705
rect 130484 21547 130550 21563
rect 130904 21705 130970 21721
rect 130904 21563 130920 21705
rect 130954 21563 130970 21705
rect 130904 21547 130970 21563
rect 131324 21705 131390 21721
rect 131324 21563 131340 21705
rect 131374 21563 131390 21705
rect 131324 21547 131390 21563
rect 131744 21705 131810 21721
rect 131744 21563 131760 21705
rect 131794 21563 131810 21705
rect 131744 21547 131810 21563
rect 132164 21705 132230 21721
rect 132164 21563 132180 21705
rect 132214 21563 132230 21705
rect 132164 21547 132230 21563
rect 132584 21705 132650 21721
rect 132584 21563 132600 21705
rect 132634 21563 132650 21705
rect 132584 21547 132650 21563
rect 133004 21705 133070 21721
rect 133004 21563 133020 21705
rect 133054 21563 133070 21705
rect 133004 21547 133070 21563
rect 133424 21705 133490 21721
rect 133424 21563 133440 21705
rect 133474 21563 133490 21705
rect 133424 21547 133490 21563
rect 133844 21705 133910 21721
rect 133844 21563 133860 21705
rect 133894 21563 133910 21705
rect 133844 21547 133910 21563
rect 134264 21705 134330 21721
rect 134264 21563 134280 21705
rect 134314 21563 134330 21705
rect 134264 21547 134330 21563
rect 134684 21705 134750 21721
rect 134684 21563 134700 21705
rect 134734 21563 134750 21705
rect 134684 21547 134750 21563
rect 135104 21705 135170 21721
rect 135104 21563 135120 21705
rect 135154 21563 135170 21705
rect 135104 21547 135170 21563
rect 126932 21516 126962 21542
rect 127142 21516 127172 21547
rect 127352 21516 127382 21542
rect 127562 21516 127592 21547
rect 127772 21516 127802 21542
rect 127982 21516 128012 21547
rect 128192 21516 128222 21542
rect 128402 21516 128432 21547
rect 128612 21516 128642 21542
rect 128822 21516 128852 21547
rect 129032 21516 129062 21542
rect 129242 21516 129272 21547
rect 129452 21516 129482 21542
rect 129662 21516 129692 21547
rect 129872 21516 129902 21542
rect 130082 21516 130112 21547
rect 130292 21516 130322 21542
rect 130502 21516 130532 21547
rect 130712 21516 130742 21542
rect 130922 21516 130952 21547
rect 131132 21516 131162 21542
rect 131342 21516 131372 21547
rect 131552 21516 131582 21542
rect 131762 21516 131792 21547
rect 131972 21516 132002 21542
rect 132182 21516 132212 21547
rect 132392 21516 132422 21542
rect 132602 21516 132632 21547
rect 132812 21516 132842 21542
rect 133022 21516 133052 21547
rect 133232 21516 133262 21542
rect 133442 21516 133472 21547
rect 133652 21516 133682 21542
rect 133862 21516 133892 21547
rect 134072 21516 134102 21542
rect 134282 21516 134312 21547
rect 134492 21516 134522 21542
rect 134702 21516 134732 21547
rect 134912 21516 134942 21542
rect 135122 21516 135152 21547
rect 126932 20485 126962 20516
rect 127142 20490 127172 20516
rect 127352 20485 127382 20516
rect 127562 20490 127592 20516
rect 127772 20485 127802 20516
rect 127982 20490 128012 20516
rect 128192 20485 128222 20516
rect 128402 20490 128432 20516
rect 128612 20485 128642 20516
rect 128822 20490 128852 20516
rect 129032 20485 129062 20516
rect 129242 20490 129272 20516
rect 129452 20485 129482 20516
rect 129662 20490 129692 20516
rect 129872 20485 129902 20516
rect 130082 20490 130112 20516
rect 130292 20485 130322 20516
rect 130502 20490 130532 20516
rect 130712 20485 130742 20516
rect 130922 20490 130952 20516
rect 131132 20485 131162 20516
rect 131342 20490 131372 20516
rect 131552 20485 131582 20516
rect 131762 20490 131792 20516
rect 131972 20485 132002 20516
rect 132182 20490 132212 20516
rect 132392 20485 132422 20516
rect 132602 20490 132632 20516
rect 132812 20485 132842 20516
rect 133022 20490 133052 20516
rect 133232 20485 133262 20516
rect 133442 20490 133472 20516
rect 133652 20485 133682 20516
rect 133862 20490 133892 20516
rect 134072 20485 134102 20516
rect 134282 20490 134312 20516
rect 134492 20485 134522 20516
rect 134702 20490 134732 20516
rect 134912 20485 134942 20516
rect 135122 20490 135152 20516
rect 126914 20469 126980 20485
rect 126914 20327 126930 20469
rect 126964 20327 126980 20469
rect 126914 20311 126980 20327
rect 127334 20469 127400 20485
rect 127334 20327 127350 20469
rect 127384 20327 127400 20469
rect 127334 20311 127400 20327
rect 127754 20469 127820 20485
rect 127754 20327 127770 20469
rect 127804 20327 127820 20469
rect 127754 20311 127820 20327
rect 128174 20469 128240 20485
rect 128174 20327 128190 20469
rect 128224 20327 128240 20469
rect 128174 20311 128240 20327
rect 128594 20469 128660 20485
rect 128594 20327 128610 20469
rect 128644 20327 128660 20469
rect 128594 20311 128660 20327
rect 129014 20469 129080 20485
rect 129014 20327 129030 20469
rect 129064 20327 129080 20469
rect 129014 20311 129080 20327
rect 129434 20469 129500 20485
rect 129434 20327 129450 20469
rect 129484 20327 129500 20469
rect 129434 20311 129500 20327
rect 129854 20469 129920 20485
rect 129854 20327 129870 20469
rect 129904 20327 129920 20469
rect 129854 20311 129920 20327
rect 130274 20469 130340 20485
rect 130274 20327 130290 20469
rect 130324 20327 130340 20469
rect 130274 20311 130340 20327
rect 130694 20469 130760 20485
rect 130694 20327 130710 20469
rect 130744 20327 130760 20469
rect 130694 20311 130760 20327
rect 131114 20469 131180 20485
rect 131114 20327 131130 20469
rect 131164 20327 131180 20469
rect 131114 20311 131180 20327
rect 131534 20469 131600 20485
rect 131534 20327 131550 20469
rect 131584 20327 131600 20469
rect 131534 20311 131600 20327
rect 131954 20469 132020 20485
rect 131954 20327 131970 20469
rect 132004 20327 132020 20469
rect 131954 20311 132020 20327
rect 132374 20469 132440 20485
rect 132374 20327 132390 20469
rect 132424 20327 132440 20469
rect 132374 20311 132440 20327
rect 132794 20469 132860 20485
rect 132794 20327 132810 20469
rect 132844 20327 132860 20469
rect 132794 20311 132860 20327
rect 133214 20469 133280 20485
rect 133214 20327 133230 20469
rect 133264 20327 133280 20469
rect 133214 20311 133280 20327
rect 133634 20469 133700 20485
rect 133634 20327 133650 20469
rect 133684 20327 133700 20469
rect 133634 20311 133700 20327
rect 134054 20469 134120 20485
rect 134054 20327 134070 20469
rect 134104 20327 134120 20469
rect 134054 20311 134120 20327
rect 134474 20469 134540 20485
rect 134474 20327 134490 20469
rect 134524 20327 134540 20469
rect 134474 20311 134540 20327
rect 134894 20469 134960 20485
rect 134894 20327 134910 20469
rect 134944 20327 134960 20469
rect 134894 20311 134960 20327
rect 126932 20280 126962 20311
rect 127142 20280 127172 20306
rect 127352 20280 127382 20311
rect 127562 20280 127592 20306
rect 127772 20280 127802 20311
rect 127982 20280 128012 20306
rect 128192 20280 128222 20311
rect 128402 20280 128432 20306
rect 128612 20280 128642 20311
rect 128822 20280 128852 20306
rect 129032 20280 129062 20311
rect 129242 20280 129272 20306
rect 129452 20280 129482 20311
rect 129662 20280 129692 20306
rect 129872 20280 129902 20311
rect 130082 20280 130112 20306
rect 130292 20280 130322 20311
rect 130502 20280 130532 20306
rect 130712 20280 130742 20311
rect 130922 20280 130952 20306
rect 131132 20280 131162 20311
rect 131342 20280 131372 20306
rect 131552 20280 131582 20311
rect 131762 20280 131792 20306
rect 131972 20280 132002 20311
rect 132182 20280 132212 20306
rect 132392 20280 132422 20311
rect 132602 20280 132632 20306
rect 132812 20280 132842 20311
rect 133022 20280 133052 20306
rect 133232 20280 133262 20311
rect 133442 20280 133472 20306
rect 133652 20280 133682 20311
rect 133862 20280 133892 20306
rect 134072 20280 134102 20311
rect 134282 20280 134312 20306
rect 134492 20280 134522 20311
rect 134702 20280 134732 20306
rect 134912 20280 134942 20311
rect 135122 20280 135152 20306
rect 126932 19254 126962 19280
rect 127142 19249 127172 19280
rect 127352 19254 127382 19280
rect 127562 19249 127592 19280
rect 127772 19254 127802 19280
rect 127982 19249 128012 19280
rect 128192 19254 128222 19280
rect 128402 19249 128432 19280
rect 128612 19254 128642 19280
rect 128822 19249 128852 19280
rect 129032 19254 129062 19280
rect 129242 19249 129272 19280
rect 129452 19254 129482 19280
rect 129662 19249 129692 19280
rect 129872 19254 129902 19280
rect 130082 19249 130112 19280
rect 130292 19254 130322 19280
rect 130502 19249 130532 19280
rect 130712 19254 130742 19280
rect 130922 19249 130952 19280
rect 131132 19254 131162 19280
rect 131342 19249 131372 19280
rect 131552 19254 131582 19280
rect 131762 19249 131792 19280
rect 131972 19254 132002 19280
rect 132182 19249 132212 19280
rect 132392 19254 132422 19280
rect 132602 19249 132632 19280
rect 132812 19254 132842 19280
rect 133022 19249 133052 19280
rect 133232 19254 133262 19280
rect 133442 19249 133472 19280
rect 133652 19254 133682 19280
rect 133862 19249 133892 19280
rect 134072 19254 134102 19280
rect 134282 19249 134312 19280
rect 134492 19254 134522 19280
rect 134702 19249 134732 19280
rect 134912 19254 134942 19280
rect 135122 19249 135152 19280
rect 127124 19233 127190 19249
rect 127124 19091 127140 19233
rect 127174 19091 127190 19233
rect 127124 19075 127190 19091
rect 127544 19233 127610 19249
rect 127544 19091 127560 19233
rect 127594 19091 127610 19233
rect 127544 19075 127610 19091
rect 127964 19233 128030 19249
rect 127964 19091 127980 19233
rect 128014 19091 128030 19233
rect 127964 19075 128030 19091
rect 128384 19233 128450 19249
rect 128384 19091 128400 19233
rect 128434 19091 128450 19233
rect 128384 19075 128450 19091
rect 128804 19233 128870 19249
rect 128804 19091 128820 19233
rect 128854 19091 128870 19233
rect 128804 19075 128870 19091
rect 129224 19233 129290 19249
rect 129224 19091 129240 19233
rect 129274 19091 129290 19233
rect 129224 19075 129290 19091
rect 129644 19233 129710 19249
rect 129644 19091 129660 19233
rect 129694 19091 129710 19233
rect 129644 19075 129710 19091
rect 130064 19233 130130 19249
rect 130064 19091 130080 19233
rect 130114 19091 130130 19233
rect 130064 19075 130130 19091
rect 130484 19233 130550 19249
rect 130484 19091 130500 19233
rect 130534 19091 130550 19233
rect 130484 19075 130550 19091
rect 130904 19233 130970 19249
rect 130904 19091 130920 19233
rect 130954 19091 130970 19233
rect 130904 19075 130970 19091
rect 131324 19233 131390 19249
rect 131324 19091 131340 19233
rect 131374 19091 131390 19233
rect 131324 19075 131390 19091
rect 131744 19233 131810 19249
rect 131744 19091 131760 19233
rect 131794 19091 131810 19233
rect 131744 19075 131810 19091
rect 132164 19233 132230 19249
rect 132164 19091 132180 19233
rect 132214 19091 132230 19233
rect 132164 19075 132230 19091
rect 132584 19233 132650 19249
rect 132584 19091 132600 19233
rect 132634 19091 132650 19233
rect 132584 19075 132650 19091
rect 133004 19233 133070 19249
rect 133004 19091 133020 19233
rect 133054 19091 133070 19233
rect 133004 19075 133070 19091
rect 133424 19233 133490 19249
rect 133424 19091 133440 19233
rect 133474 19091 133490 19233
rect 133424 19075 133490 19091
rect 133844 19233 133910 19249
rect 133844 19091 133860 19233
rect 133894 19091 133910 19233
rect 133844 19075 133910 19091
rect 134264 19233 134330 19249
rect 134264 19091 134280 19233
rect 134314 19091 134330 19233
rect 134264 19075 134330 19091
rect 134684 19233 134750 19249
rect 134684 19091 134700 19233
rect 134734 19091 134750 19233
rect 134684 19075 134750 19091
rect 135104 19233 135170 19249
rect 135104 19091 135120 19233
rect 135154 19091 135170 19233
rect 135104 19075 135170 19091
rect 126932 19044 126962 19070
rect 127142 19044 127172 19075
rect 127352 19044 127382 19070
rect 127562 19044 127592 19075
rect 127772 19044 127802 19070
rect 127982 19044 128012 19075
rect 128192 19044 128222 19070
rect 128402 19044 128432 19075
rect 128612 19044 128642 19070
rect 128822 19044 128852 19075
rect 129032 19044 129062 19070
rect 129242 19044 129272 19075
rect 129452 19044 129482 19070
rect 129662 19044 129692 19075
rect 129872 19044 129902 19070
rect 130082 19044 130112 19075
rect 130292 19044 130322 19070
rect 130502 19044 130532 19075
rect 130712 19044 130742 19070
rect 130922 19044 130952 19075
rect 131132 19044 131162 19070
rect 131342 19044 131372 19075
rect 131552 19044 131582 19070
rect 131762 19044 131792 19075
rect 131972 19044 132002 19070
rect 132182 19044 132212 19075
rect 132392 19044 132422 19070
rect 132602 19044 132632 19075
rect 132812 19044 132842 19070
rect 133022 19044 133052 19075
rect 133232 19044 133262 19070
rect 133442 19044 133472 19075
rect 133652 19044 133682 19070
rect 133862 19044 133892 19075
rect 134072 19044 134102 19070
rect 134282 19044 134312 19075
rect 134492 19044 134522 19070
rect 134702 19044 134732 19075
rect 134912 19044 134942 19070
rect 135122 19044 135152 19075
rect 126932 18014 126962 18044
rect 127142 18018 127172 18044
rect 127352 18014 127382 18044
rect 127562 18018 127592 18044
rect 127772 18014 127802 18044
rect 127982 18018 128012 18044
rect 128192 18014 128222 18044
rect 128402 18018 128432 18044
rect 128612 18014 128642 18044
rect 128822 18018 128852 18044
rect 129032 18014 129062 18044
rect 129242 18018 129272 18044
rect 129452 18014 129482 18044
rect 129662 18018 129692 18044
rect 129872 18014 129902 18044
rect 130082 18018 130112 18044
rect 130292 18014 130322 18044
rect 130502 18018 130532 18044
rect 130712 18014 130742 18044
rect 130922 18018 130952 18044
rect 131132 18014 131162 18044
rect 131342 18018 131372 18044
rect 131552 18014 131582 18044
rect 131762 18018 131792 18044
rect 131972 18014 132002 18044
rect 132182 18018 132212 18044
rect 132392 18014 132422 18044
rect 132602 18018 132632 18044
rect 132812 18014 132842 18044
rect 133022 18018 133052 18044
rect 133232 18014 133262 18044
rect 133442 18018 133472 18044
rect 133652 18014 133682 18044
rect 133862 18018 133892 18044
rect 134072 18014 134102 18044
rect 134282 18018 134312 18044
rect 134492 18014 134522 18044
rect 134702 18018 134732 18044
rect 134912 18014 134942 18044
rect 135122 18018 135152 18044
rect 126914 17997 127030 18014
rect 125424 17946 125540 17962
rect 126914 17962 126930 17997
rect 126964 17996 127030 17997
rect 127014 17962 127030 17996
rect 126914 17946 127030 17962
rect 127334 17997 127450 18014
rect 127334 17962 127350 17997
rect 127384 17996 127450 17997
rect 127434 17962 127450 17996
rect 127334 17946 127450 17962
rect 127754 17997 127870 18014
rect 127754 17962 127770 17997
rect 127804 17996 127870 17997
rect 127854 17962 127870 17996
rect 127754 17946 127870 17962
rect 128174 17997 128290 18014
rect 128174 17962 128190 17997
rect 128224 17996 128290 17997
rect 128274 17962 128290 17996
rect 128174 17946 128290 17962
rect 128594 17997 128710 18014
rect 128594 17962 128610 17997
rect 128644 17996 128710 17997
rect 128694 17962 128710 17996
rect 128594 17946 128710 17962
rect 129014 17997 129130 18014
rect 129014 17962 129030 17997
rect 129064 17996 129130 17997
rect 129114 17962 129130 17996
rect 129014 17946 129130 17962
rect 129434 17997 129550 18014
rect 129434 17962 129450 17997
rect 129484 17996 129550 17997
rect 129534 17962 129550 17996
rect 129434 17946 129550 17962
rect 129854 17997 129970 18014
rect 129854 17962 129870 17997
rect 129904 17996 129970 17997
rect 129954 17962 129970 17996
rect 129854 17946 129970 17962
rect 130274 17997 130390 18014
rect 130274 17962 130290 17997
rect 130324 17996 130390 17997
rect 130374 17962 130390 17996
rect 130274 17946 130390 17962
rect 130694 17997 130810 18014
rect 130694 17962 130710 17997
rect 130744 17996 130810 17997
rect 130794 17962 130810 17996
rect 130694 17946 130810 17962
rect 131114 17997 131230 18014
rect 131114 17962 131130 17997
rect 131164 17996 131230 17997
rect 131214 17962 131230 17996
rect 131114 17946 131230 17962
rect 131534 17997 131650 18014
rect 131534 17962 131550 17997
rect 131584 17996 131650 17997
rect 131634 17962 131650 17996
rect 131534 17946 131650 17962
rect 131954 17997 132070 18014
rect 131954 17962 131970 17997
rect 132004 17996 132070 17997
rect 132054 17962 132070 17996
rect 131954 17946 132070 17962
rect 132374 17997 132490 18014
rect 132374 17962 132390 17997
rect 132424 17996 132490 17997
rect 132474 17962 132490 17996
rect 132374 17946 132490 17962
rect 132794 17997 132910 18014
rect 132794 17962 132810 17997
rect 132844 17996 132910 17997
rect 132894 17962 132910 17996
rect 132794 17946 132910 17962
rect 133214 17997 133330 18014
rect 133214 17962 133230 17997
rect 133264 17996 133330 17997
rect 133314 17962 133330 17996
rect 133214 17946 133330 17962
rect 133634 17997 133750 18014
rect 133634 17962 133650 17997
rect 133684 17996 133750 17997
rect 133734 17962 133750 17996
rect 133634 17946 133750 17962
rect 134054 17997 134170 18014
rect 134054 17962 134070 17997
rect 134104 17996 134170 17997
rect 134154 17962 134170 17996
rect 134054 17946 134170 17962
rect 134474 17997 134590 18014
rect 134474 17962 134490 17997
rect 134524 17996 134590 17997
rect 134574 17962 134590 17996
rect 134474 17946 134590 17962
rect 134894 17997 135010 18014
rect 134894 17962 134910 17997
rect 134944 17996 135010 17997
rect 134994 17962 135010 17996
rect 134894 17946 135010 17962
rect 116428 16918 116458 16944
rect 116522 16918 116552 16944
rect 116428 16390 116458 16518
rect 116522 16476 116552 16518
rect 116500 16464 116594 16476
rect 116500 16432 116518 16464
rect 116576 16432 116594 16464
rect 116500 16418 116594 16432
rect 116342 16378 116458 16390
rect 116342 16346 116360 16378
rect 116418 16346 116458 16378
rect 116342 16332 116458 16346
rect 116428 16298 116458 16332
rect 116522 16298 116552 16418
rect 116428 15872 116458 15898
rect 116522 15872 116552 15898
rect 115902 15490 115932 15516
rect 116428 15492 116458 15518
rect 116522 15492 116552 15518
rect 115902 15059 115932 15090
rect 115884 15043 115950 15059
rect 116428 15058 116458 15092
rect 115884 15009 115900 15043
rect 115934 15009 115950 15043
rect 115884 14906 115950 15009
rect 116342 15044 116458 15058
rect 116342 15012 116360 15044
rect 116418 15012 116458 15044
rect 116342 15000 116458 15012
rect 115884 14872 115900 14906
rect 115934 14872 115950 14906
rect 116428 14872 116458 15000
rect 116522 14972 116552 15092
rect 116500 14958 116594 14972
rect 116500 14926 116518 14958
rect 116576 14926 116594 14958
rect 116500 14914 116594 14926
rect 116522 14872 116552 14914
rect 115884 14856 115950 14872
rect 115902 14834 115932 14856
rect 115902 14608 115932 14634
rect 116428 14446 116458 14472
rect 116522 14446 116552 14472
rect 119248 13426 119364 13442
rect 119248 13392 119264 13426
rect 119348 13392 119364 13426
rect 119248 13376 119364 13392
rect 119890 13428 120006 13444
rect 119890 13393 119906 13428
rect 119990 13394 120006 13428
rect 119940 13393 120006 13394
rect 119890 13376 120006 13393
rect 120310 13428 120426 13444
rect 120310 13393 120326 13428
rect 120410 13394 120426 13428
rect 120360 13393 120426 13394
rect 120310 13376 120426 13393
rect 120730 13428 120846 13444
rect 120730 13393 120746 13428
rect 120830 13394 120846 13428
rect 120780 13393 120846 13394
rect 120730 13376 120846 13393
rect 121150 13428 121266 13444
rect 121150 13393 121166 13428
rect 121250 13394 121266 13428
rect 121200 13393 121266 13394
rect 121150 13376 121266 13393
rect 119170 13346 119200 13372
rect 119266 13346 119296 13376
rect 119908 13346 119938 13376
rect 120118 13346 120148 13372
rect 120328 13346 120358 13376
rect 120538 13346 120568 13372
rect 120748 13346 120778 13376
rect 120958 13346 120988 13372
rect 121168 13346 121198 13376
rect 121378 13346 121408 13372
rect 119170 12315 119200 12346
rect 119266 12320 119296 12346
rect 119908 12320 119938 12346
rect 120118 12315 120148 12346
rect 120328 12320 120358 12346
rect 120538 12315 120568 12346
rect 120748 12320 120778 12346
rect 120958 12316 120988 12346
rect 121168 12320 121198 12346
rect 121378 12316 121408 12346
rect 119152 12299 119218 12315
rect 119152 12156 119168 12299
rect 119202 12156 119218 12299
rect 119152 12140 119218 12156
rect 120100 12299 120166 12315
rect 120100 12156 120116 12299
rect 120150 12156 120166 12299
rect 120100 12140 120166 12156
rect 120520 12299 120586 12315
rect 120520 12156 120536 12299
rect 120570 12156 120586 12299
rect 120940 12300 121056 12316
rect 120940 12265 120956 12300
rect 121040 12266 121056 12300
rect 120990 12265 121056 12266
rect 120940 12248 121056 12265
rect 121360 12300 121476 12316
rect 121360 12265 121376 12300
rect 121460 12266 121476 12300
rect 121410 12265 121476 12266
rect 121360 12248 121476 12265
rect 119170 12118 119200 12140
rect 120118 12118 120148 12140
rect 120328 12118 120358 12144
rect 120520 12140 120586 12156
rect 120538 12118 120568 12140
rect 120748 12118 120778 12144
rect 119170 11092 119200 11118
rect 120118 11092 120148 11118
rect 120328 11088 120358 11118
rect 120538 11092 120568 11118
rect 120748 11088 120778 11118
rect 120310 11072 120426 11088
rect 120310 11037 120326 11072
rect 120410 11038 120426 11072
rect 120360 11037 120426 11038
rect 120310 11020 120426 11037
rect 120730 11072 120846 11088
rect 120730 11037 120746 11072
rect 120830 11038 120846 11072
rect 120780 11037 120846 11038
rect 120730 11020 120846 11037
rect 122064 13428 122180 13444
rect 122064 13393 122080 13428
rect 122164 13394 122180 13428
rect 122114 13393 122180 13394
rect 122064 13376 122180 13393
rect 122484 13428 122600 13444
rect 122484 13393 122500 13428
rect 122584 13394 122600 13428
rect 122534 13393 122600 13394
rect 122484 13376 122600 13393
rect 122904 13428 123020 13444
rect 122904 13393 122920 13428
rect 123004 13394 123020 13428
rect 122954 13393 123020 13394
rect 122904 13376 123020 13393
rect 123324 13428 123440 13444
rect 123324 13393 123340 13428
rect 123424 13394 123440 13428
rect 123374 13393 123440 13394
rect 123324 13376 123440 13393
rect 123744 13428 123860 13444
rect 123744 13393 123760 13428
rect 123844 13394 123860 13428
rect 123794 13393 123860 13394
rect 123744 13376 123860 13393
rect 124164 13428 124280 13444
rect 124164 13393 124180 13428
rect 124264 13394 124280 13428
rect 124214 13393 124280 13394
rect 124164 13376 124280 13393
rect 124584 13428 124700 13444
rect 124584 13393 124600 13428
rect 124684 13394 124700 13428
rect 124634 13393 124700 13394
rect 124584 13376 124700 13393
rect 125004 13428 125120 13444
rect 125004 13393 125020 13428
rect 125104 13394 125120 13428
rect 125054 13393 125120 13394
rect 125004 13376 125120 13393
rect 125424 13428 125540 13444
rect 125424 13393 125440 13428
rect 125524 13394 125540 13428
rect 125474 13393 125540 13394
rect 125424 13376 125540 13393
rect 122082 13346 122112 13376
rect 122292 13346 122322 13372
rect 122502 13346 122532 13376
rect 122712 13346 122742 13372
rect 122922 13346 122952 13376
rect 123132 13346 123162 13372
rect 123342 13346 123372 13376
rect 123552 13346 123582 13372
rect 123762 13346 123792 13376
rect 123972 13346 124002 13372
rect 124182 13346 124212 13376
rect 124392 13346 124422 13372
rect 124602 13346 124632 13376
rect 124812 13346 124842 13372
rect 125022 13346 125052 13376
rect 125232 13346 125262 13372
rect 125442 13346 125472 13376
rect 125652 13346 125682 13372
rect 122082 12320 122112 12346
rect 122292 12315 122322 12346
rect 122502 12320 122532 12346
rect 122712 12315 122742 12346
rect 122922 12320 122952 12346
rect 123132 12315 123162 12346
rect 123342 12320 123372 12346
rect 123552 12315 123582 12346
rect 123762 12320 123792 12346
rect 123972 12315 124002 12346
rect 124182 12320 124212 12346
rect 124392 12315 124422 12346
rect 124602 12320 124632 12346
rect 124812 12315 124842 12346
rect 125022 12320 125052 12346
rect 125232 12315 125262 12346
rect 125442 12320 125472 12346
rect 125652 12315 125682 12346
rect 122274 12299 122340 12315
rect 122274 12157 122290 12299
rect 122324 12157 122340 12299
rect 122274 12141 122340 12157
rect 122694 12299 122760 12315
rect 122694 12157 122710 12299
rect 122744 12157 122760 12299
rect 122694 12141 122760 12157
rect 123114 12299 123180 12315
rect 123114 12157 123130 12299
rect 123164 12157 123180 12299
rect 123114 12141 123180 12157
rect 123534 12299 123600 12315
rect 123534 12157 123550 12299
rect 123584 12157 123600 12299
rect 123534 12141 123600 12157
rect 123954 12299 124020 12315
rect 123954 12157 123970 12299
rect 124004 12157 124020 12299
rect 123954 12141 124020 12157
rect 124374 12299 124440 12315
rect 124374 12157 124390 12299
rect 124424 12157 124440 12299
rect 124374 12141 124440 12157
rect 124794 12299 124860 12315
rect 124794 12157 124810 12299
rect 124844 12157 124860 12299
rect 124794 12141 124860 12157
rect 125214 12299 125280 12315
rect 125214 12157 125230 12299
rect 125264 12157 125280 12299
rect 125214 12141 125280 12157
rect 125634 12299 125700 12315
rect 125634 12157 125650 12299
rect 125684 12157 125700 12299
rect 125634 12141 125700 12157
rect 122082 12110 122112 12136
rect 122292 12110 122322 12141
rect 122502 12110 122532 12136
rect 122712 12110 122742 12141
rect 122922 12110 122952 12136
rect 123132 12110 123162 12141
rect 123342 12110 123372 12136
rect 123552 12110 123582 12141
rect 123762 12110 123792 12136
rect 123972 12110 124002 12141
rect 124182 12110 124212 12136
rect 124392 12110 124422 12141
rect 124602 12110 124632 12136
rect 124812 12110 124842 12141
rect 125022 12110 125052 12136
rect 125232 12110 125262 12141
rect 125442 12110 125472 12136
rect 125652 12110 125682 12141
rect 122082 11080 122112 11110
rect 122292 11084 122322 11110
rect 122502 11080 122532 11110
rect 122712 11084 122742 11110
rect 122922 11080 122952 11110
rect 123132 11084 123162 11110
rect 123342 11080 123372 11110
rect 123552 11084 123582 11110
rect 123762 11080 123792 11110
rect 123972 11084 124002 11110
rect 124182 11080 124212 11110
rect 124392 11084 124422 11110
rect 124602 11080 124632 11110
rect 124812 11084 124842 11110
rect 125022 11080 125052 11110
rect 125232 11084 125262 11110
rect 125442 11080 125472 11110
rect 125652 11084 125682 11110
rect 122064 11064 122180 11080
rect 122064 11029 122080 11064
rect 122164 11030 122180 11064
rect 122114 11029 122180 11030
rect 122064 11012 122180 11029
rect 122484 11064 122600 11080
rect 122484 11029 122500 11064
rect 122584 11030 122600 11064
rect 122534 11029 122600 11030
rect 122484 11012 122600 11029
rect 122904 11064 123020 11080
rect 122904 11029 122920 11064
rect 123004 11030 123020 11064
rect 122954 11029 123020 11030
rect 122904 11012 123020 11029
rect 123324 11064 123440 11080
rect 123324 11029 123340 11064
rect 123424 11030 123440 11064
rect 123374 11029 123440 11030
rect 123324 11012 123440 11029
rect 123744 11064 123860 11080
rect 123744 11029 123760 11064
rect 123844 11030 123860 11064
rect 123794 11029 123860 11030
rect 123744 11012 123860 11029
rect 124164 11064 124280 11080
rect 124164 11029 124180 11064
rect 124264 11030 124280 11064
rect 124214 11029 124280 11030
rect 124164 11012 124280 11029
rect 124584 11064 124700 11080
rect 124584 11029 124600 11064
rect 124684 11030 124700 11064
rect 124634 11029 124700 11030
rect 124584 11012 124700 11029
rect 125004 11064 125120 11080
rect 125004 11029 125020 11064
rect 125104 11030 125120 11064
rect 125054 11029 125120 11030
rect 125004 11012 125120 11029
rect 125424 11064 125540 11080
rect 125424 11029 125440 11064
rect 125524 11030 125540 11064
rect 125474 11029 125540 11030
rect 125424 11012 125540 11029
rect 122064 9172 122180 9188
rect 122064 9137 122080 9172
rect 122164 9138 122180 9172
rect 122114 9137 122180 9138
rect 122064 9120 122180 9137
rect 122484 9172 122600 9188
rect 122484 9137 122500 9172
rect 122584 9138 122600 9172
rect 122534 9137 122600 9138
rect 122484 9120 122600 9137
rect 122904 9172 123020 9188
rect 122904 9132 122920 9172
rect 123004 9138 123020 9172
rect 122954 9132 123020 9138
rect 122904 9120 123020 9132
rect 123324 9172 123440 9188
rect 123324 9132 123340 9172
rect 123424 9138 123440 9172
rect 123374 9132 123440 9138
rect 123324 9120 123440 9132
rect 123744 9172 123860 9188
rect 123744 9132 123760 9172
rect 123844 9138 123860 9172
rect 123794 9132 123860 9138
rect 123744 9120 123860 9132
rect 124164 9172 124280 9188
rect 124164 9132 124180 9172
rect 124264 9138 124280 9172
rect 124214 9132 124280 9138
rect 124164 9120 124280 9132
rect 124584 9172 124700 9188
rect 124584 9132 124600 9172
rect 124684 9138 124700 9172
rect 124634 9132 124700 9138
rect 124584 9120 124700 9132
rect 125004 9172 125120 9188
rect 125004 9132 125020 9172
rect 125104 9138 125120 9172
rect 125054 9132 125120 9138
rect 125004 9120 125120 9132
rect 125424 9172 125540 9188
rect 125424 9132 125440 9172
rect 125524 9138 125540 9172
rect 125474 9132 125540 9138
rect 125424 9120 125540 9132
rect 122082 9094 122112 9120
rect 122292 9094 122322 9120
rect 122502 9094 122532 9120
rect 122712 9094 122742 9120
rect 122904 9116 122970 9120
rect 122922 9094 122952 9116
rect 123132 9094 123162 9120
rect 123324 9116 123390 9120
rect 123342 9094 123372 9116
rect 123552 9094 123582 9120
rect 123744 9116 123810 9120
rect 123762 9094 123792 9116
rect 123972 9094 124002 9120
rect 124164 9116 124230 9120
rect 124182 9094 124212 9116
rect 124392 9094 124422 9120
rect 124584 9116 124650 9120
rect 124602 9094 124632 9116
rect 124812 9094 124842 9120
rect 125004 9116 125070 9120
rect 125022 9094 125052 9116
rect 125232 9094 125262 9120
rect 125424 9116 125490 9120
rect 125442 9094 125472 9116
rect 125652 9094 125682 9120
rect 122082 8068 122112 8094
rect 122292 8064 122322 8094
rect 122502 8068 122532 8094
rect 122712 8072 122742 8094
rect 122694 8064 122760 8072
rect 122922 8068 122952 8094
rect 123132 8072 123162 8094
rect 123114 8064 123180 8072
rect 123342 8068 123372 8094
rect 123552 8072 123582 8094
rect 123534 8064 123600 8072
rect 123762 8068 123792 8094
rect 123972 8072 124002 8094
rect 123954 8064 124020 8072
rect 124182 8068 124212 8094
rect 124392 8072 124422 8094
rect 124374 8064 124440 8072
rect 124602 8068 124632 8094
rect 124812 8072 124842 8094
rect 124794 8064 124860 8072
rect 125022 8068 125052 8094
rect 125232 8072 125262 8094
rect 125214 8064 125280 8072
rect 125442 8068 125472 8094
rect 125652 8072 125682 8094
rect 125634 8064 125700 8072
rect 122274 8048 122390 8064
rect 122274 8014 122290 8048
rect 122374 8014 122390 8048
rect 122274 7996 122390 8014
rect 122694 8056 122810 8064
rect 122694 8014 122710 8056
rect 122744 8048 122810 8056
rect 122794 8014 122810 8048
rect 122694 7996 122810 8014
rect 123114 8056 123230 8064
rect 123114 8014 123130 8056
rect 123164 8048 123230 8056
rect 123214 8014 123230 8048
rect 123114 7996 123230 8014
rect 123534 8056 123650 8064
rect 123534 8014 123550 8056
rect 123584 8048 123650 8056
rect 123634 8014 123650 8048
rect 123534 7996 123650 8014
rect 123954 8056 124070 8064
rect 123954 8014 123970 8056
rect 124004 8048 124070 8056
rect 124054 8014 124070 8048
rect 123954 7996 124070 8014
rect 124374 8056 124490 8064
rect 124374 8014 124390 8056
rect 124424 8048 124490 8056
rect 124474 8014 124490 8048
rect 124374 7996 124490 8014
rect 124794 8056 124910 8064
rect 124794 8014 124810 8056
rect 124844 8048 124910 8056
rect 124894 8014 124910 8048
rect 124794 7996 124910 8014
rect 125214 8056 125330 8064
rect 125214 8014 125230 8056
rect 125264 8048 125330 8056
rect 125314 8014 125330 8048
rect 125214 7996 125330 8014
rect 125634 8056 125750 8064
rect 125634 8014 125650 8056
rect 125684 8048 125750 8056
rect 125734 8014 125750 8048
rect 125634 7996 125750 8014
<< polycont >>
rect 126930 28018 127014 28052
rect 127350 28018 127434 28052
rect 127770 28018 127854 28052
rect 128190 28018 128274 28052
rect 128610 28018 128694 28052
rect 129030 28018 129114 28052
rect 129450 28018 129534 28052
rect 129870 28018 129954 28052
rect 130290 28018 130374 28052
rect 130710 28018 130794 28052
rect 131130 28018 131214 28052
rect 131550 28018 131634 28052
rect 131970 28018 132054 28052
rect 132390 28018 132474 28052
rect 132810 28018 132894 28052
rect 133230 28018 133314 28052
rect 133650 28018 133734 28052
rect 134070 28018 134154 28052
rect 134490 28018 134574 28052
rect 134910 28018 134994 28052
rect 127140 26800 127174 26942
rect 127560 26800 127594 26942
rect 127980 26800 128014 26942
rect 128400 26800 128434 26942
rect 128820 26800 128854 26942
rect 129240 26800 129274 26942
rect 129660 26800 129694 26942
rect 130080 26800 130114 26942
rect 130500 26800 130534 26942
rect 130920 26800 130954 26942
rect 131340 26800 131374 26942
rect 131760 26800 131794 26942
rect 132180 26800 132214 26942
rect 132600 26800 132634 26942
rect 133020 26800 133054 26942
rect 133440 26800 133474 26942
rect 133860 26800 133894 26942
rect 134280 26800 134314 26942
rect 134700 26800 134734 26942
rect 135120 26800 135154 26942
rect 126930 25690 127014 25724
rect 127350 25690 127434 25724
rect 127770 25690 127854 25724
rect 128190 25690 128274 25724
rect 128610 25690 128694 25724
rect 129030 25690 129114 25724
rect 129450 25690 129534 25724
rect 129870 25690 129954 25724
rect 130290 25690 130374 25724
rect 130710 25690 130794 25724
rect 131130 25690 131214 25724
rect 131550 25690 131634 25724
rect 131970 25690 132054 25724
rect 132390 25690 132474 25724
rect 132810 25690 132894 25724
rect 133230 25690 133314 25724
rect 133650 25690 133734 25724
rect 134070 25690 134154 25724
rect 134490 25690 134574 25724
rect 134910 25690 134994 25724
rect 126930 22832 126964 22833
rect 126930 22798 127014 22832
rect 127350 22832 127384 22833
rect 127350 22798 127434 22832
rect 127770 22832 127804 22833
rect 127770 22798 127854 22832
rect 128190 22832 128224 22833
rect 128190 22798 128274 22832
rect 128610 22832 128644 22833
rect 128610 22798 128694 22832
rect 129030 22832 129064 22833
rect 129030 22798 129114 22832
rect 129450 22832 129484 22833
rect 129450 22798 129534 22832
rect 129870 22832 129904 22833
rect 129870 22798 129954 22832
rect 130290 22832 130324 22833
rect 130290 22798 130374 22832
rect 130710 22832 130744 22833
rect 130710 22798 130794 22832
rect 131130 22832 131164 22833
rect 131130 22798 131214 22832
rect 131550 22832 131584 22833
rect 131550 22798 131634 22832
rect 131970 22832 132004 22833
rect 131970 22798 132054 22832
rect 132390 22832 132424 22833
rect 132390 22798 132474 22832
rect 132810 22832 132844 22833
rect 132810 22798 132894 22832
rect 133230 22832 133264 22833
rect 133230 22798 133314 22832
rect 133650 22832 133684 22833
rect 133650 22798 133734 22832
rect 134070 22832 134104 22833
rect 134070 22798 134154 22832
rect 134490 22832 134524 22833
rect 134490 22798 134574 22832
rect 134910 22832 134944 22833
rect 134910 22798 134994 22832
rect 122290 21942 122374 21976
rect 122710 21942 122794 21976
rect 122710 21934 122744 21942
rect 123130 21942 123214 21976
rect 123130 21934 123164 21942
rect 123550 21942 123634 21976
rect 123550 21934 123584 21942
rect 123970 21942 124054 21976
rect 123970 21934 124004 21942
rect 124390 21942 124474 21976
rect 124390 21934 124424 21942
rect 124810 21942 124894 21976
rect 124810 21934 124844 21942
rect 125230 21942 125314 21976
rect 125230 21934 125264 21942
rect 125650 21942 125734 21976
rect 125650 21934 125684 21942
rect 122080 20852 122114 20853
rect 122080 20818 122164 20852
rect 122500 20852 122534 20853
rect 122500 20818 122584 20852
rect 122920 20852 122954 20858
rect 122920 20818 123004 20852
rect 123340 20852 123374 20858
rect 123340 20818 123424 20852
rect 123760 20852 123794 20858
rect 123760 20818 123844 20852
rect 124180 20852 124214 20858
rect 124180 20818 124264 20852
rect 124600 20852 124634 20858
rect 124600 20818 124684 20852
rect 125020 20852 125054 20858
rect 125020 20818 125104 20852
rect 125440 20852 125474 20858
rect 125440 20818 125524 20852
rect 120326 20352 120360 20353
rect 120326 20318 120410 20352
rect 120746 20352 120780 20353
rect 120746 20318 120830 20352
rect 119168 19091 119202 19234
rect 120116 19091 120150 19234
rect 120536 19091 120570 19234
rect 120956 19124 120990 19125
rect 120956 19090 121040 19124
rect 121376 19124 121410 19125
rect 121376 19090 121460 19124
rect 119264 17964 119348 17998
rect 119906 17996 119940 17997
rect 119906 17962 119990 17996
rect 120326 17996 120360 17997
rect 120326 17962 120410 17996
rect 120746 17996 120780 17997
rect 120746 17962 120830 17996
rect 121166 17996 121200 17997
rect 121166 17962 121250 17996
rect 122080 20360 122114 20361
rect 122080 20326 122164 20360
rect 122500 20360 122534 20361
rect 122500 20326 122584 20360
rect 122920 20360 122954 20361
rect 122920 20326 123004 20360
rect 123340 20360 123374 20361
rect 123340 20326 123424 20360
rect 123760 20360 123794 20361
rect 123760 20326 123844 20360
rect 124180 20360 124214 20361
rect 124180 20326 124264 20360
rect 124600 20360 124634 20361
rect 124600 20326 124684 20360
rect 125020 20360 125054 20361
rect 125020 20326 125104 20360
rect 125440 20360 125474 20361
rect 125440 20326 125524 20360
rect 122290 19091 122324 19233
rect 122710 19091 122744 19233
rect 123130 19091 123164 19233
rect 123550 19091 123584 19233
rect 123970 19091 124004 19233
rect 124390 19091 124424 19233
rect 124810 19091 124844 19233
rect 125230 19091 125264 19233
rect 125650 19091 125684 19233
rect 122080 17996 122114 17997
rect 122080 17962 122164 17996
rect 122500 17996 122534 17997
rect 122500 17962 122584 17996
rect 122920 17996 122954 17997
rect 122920 17962 123004 17996
rect 123340 17996 123374 17997
rect 123340 17962 123424 17996
rect 123760 17996 123794 17997
rect 123760 17962 123844 17996
rect 124180 17996 124214 17997
rect 124180 17962 124264 17996
rect 124600 17996 124634 17997
rect 124600 17962 124684 17996
rect 125020 17996 125054 17997
rect 125020 17962 125104 17996
rect 125440 17996 125474 17997
rect 125440 17962 125524 17996
rect 127140 21563 127174 21705
rect 127560 21563 127594 21705
rect 127980 21563 128014 21705
rect 128400 21563 128434 21705
rect 128820 21563 128854 21705
rect 129240 21563 129274 21705
rect 129660 21563 129694 21705
rect 130080 21563 130114 21705
rect 130500 21563 130534 21705
rect 130920 21563 130954 21705
rect 131340 21563 131374 21705
rect 131760 21563 131794 21705
rect 132180 21563 132214 21705
rect 132600 21563 132634 21705
rect 133020 21563 133054 21705
rect 133440 21563 133474 21705
rect 133860 21563 133894 21705
rect 134280 21563 134314 21705
rect 134700 21563 134734 21705
rect 135120 21563 135154 21705
rect 126930 20327 126964 20469
rect 127350 20327 127384 20469
rect 127770 20327 127804 20469
rect 128190 20327 128224 20469
rect 128610 20327 128644 20469
rect 129030 20327 129064 20469
rect 129450 20327 129484 20469
rect 129870 20327 129904 20469
rect 130290 20327 130324 20469
rect 130710 20327 130744 20469
rect 131130 20327 131164 20469
rect 131550 20327 131584 20469
rect 131970 20327 132004 20469
rect 132390 20327 132424 20469
rect 132810 20327 132844 20469
rect 133230 20327 133264 20469
rect 133650 20327 133684 20469
rect 134070 20327 134104 20469
rect 134490 20327 134524 20469
rect 134910 20327 134944 20469
rect 127140 19091 127174 19233
rect 127560 19091 127594 19233
rect 127980 19091 128014 19233
rect 128400 19091 128434 19233
rect 128820 19091 128854 19233
rect 129240 19091 129274 19233
rect 129660 19091 129694 19233
rect 130080 19091 130114 19233
rect 130500 19091 130534 19233
rect 130920 19091 130954 19233
rect 131340 19091 131374 19233
rect 131760 19091 131794 19233
rect 132180 19091 132214 19233
rect 132600 19091 132634 19233
rect 133020 19091 133054 19233
rect 133440 19091 133474 19233
rect 133860 19091 133894 19233
rect 134280 19091 134314 19233
rect 134700 19091 134734 19233
rect 135120 19091 135154 19233
rect 126930 17996 126964 17997
rect 126930 17962 127014 17996
rect 127350 17996 127384 17997
rect 127350 17962 127434 17996
rect 127770 17996 127804 17997
rect 127770 17962 127854 17996
rect 128190 17996 128224 17997
rect 128190 17962 128274 17996
rect 128610 17996 128644 17997
rect 128610 17962 128694 17996
rect 129030 17996 129064 17997
rect 129030 17962 129114 17996
rect 129450 17996 129484 17997
rect 129450 17962 129534 17996
rect 129870 17996 129904 17997
rect 129870 17962 129954 17996
rect 130290 17996 130324 17997
rect 130290 17962 130374 17996
rect 130710 17996 130744 17997
rect 130710 17962 130794 17996
rect 131130 17996 131164 17997
rect 131130 17962 131214 17996
rect 131550 17996 131584 17997
rect 131550 17962 131634 17996
rect 131970 17996 132004 17997
rect 131970 17962 132054 17996
rect 132390 17996 132424 17997
rect 132390 17962 132474 17996
rect 132810 17996 132844 17997
rect 132810 17962 132894 17996
rect 133230 17996 133264 17997
rect 133230 17962 133314 17996
rect 133650 17996 133684 17997
rect 133650 17962 133734 17996
rect 134070 17996 134104 17997
rect 134070 17962 134154 17996
rect 134490 17996 134524 17997
rect 134490 17962 134574 17996
rect 134910 17996 134944 17997
rect 134910 17962 134994 17996
rect 116518 16432 116576 16464
rect 116360 16346 116418 16378
rect 115900 15009 115934 15043
rect 116360 15012 116418 15044
rect 115900 14872 115934 14906
rect 116518 14926 116576 14958
rect 119264 13392 119348 13426
rect 119906 13394 119990 13428
rect 119906 13393 119940 13394
rect 120326 13394 120410 13428
rect 120326 13393 120360 13394
rect 120746 13394 120830 13428
rect 120746 13393 120780 13394
rect 121166 13394 121250 13428
rect 121166 13393 121200 13394
rect 119168 12156 119202 12299
rect 120116 12156 120150 12299
rect 120536 12156 120570 12299
rect 120956 12266 121040 12300
rect 120956 12265 120990 12266
rect 121376 12266 121460 12300
rect 121376 12265 121410 12266
rect 120326 11038 120410 11072
rect 120326 11037 120360 11038
rect 120746 11038 120830 11072
rect 120746 11037 120780 11038
rect 122080 13394 122164 13428
rect 122080 13393 122114 13394
rect 122500 13394 122584 13428
rect 122500 13393 122534 13394
rect 122920 13394 123004 13428
rect 122920 13393 122954 13394
rect 123340 13394 123424 13428
rect 123340 13393 123374 13394
rect 123760 13394 123844 13428
rect 123760 13393 123794 13394
rect 124180 13394 124264 13428
rect 124180 13393 124214 13394
rect 124600 13394 124684 13428
rect 124600 13393 124634 13394
rect 125020 13394 125104 13428
rect 125020 13393 125054 13394
rect 125440 13394 125524 13428
rect 125440 13393 125474 13394
rect 122290 12157 122324 12299
rect 122710 12157 122744 12299
rect 123130 12157 123164 12299
rect 123550 12157 123584 12299
rect 123970 12157 124004 12299
rect 124390 12157 124424 12299
rect 124810 12157 124844 12299
rect 125230 12157 125264 12299
rect 125650 12157 125684 12299
rect 122080 11030 122164 11064
rect 122080 11029 122114 11030
rect 122500 11030 122584 11064
rect 122500 11029 122534 11030
rect 122920 11030 123004 11064
rect 122920 11029 122954 11030
rect 123340 11030 123424 11064
rect 123340 11029 123374 11030
rect 123760 11030 123844 11064
rect 123760 11029 123794 11030
rect 124180 11030 124264 11064
rect 124180 11029 124214 11030
rect 124600 11030 124684 11064
rect 124600 11029 124634 11030
rect 125020 11030 125104 11064
rect 125020 11029 125054 11030
rect 125440 11030 125524 11064
rect 125440 11029 125474 11030
rect 122080 9138 122164 9172
rect 122080 9137 122114 9138
rect 122500 9138 122584 9172
rect 122500 9137 122534 9138
rect 122920 9138 123004 9172
rect 122920 9132 122954 9138
rect 123340 9138 123424 9172
rect 123340 9132 123374 9138
rect 123760 9138 123844 9172
rect 123760 9132 123794 9138
rect 124180 9138 124264 9172
rect 124180 9132 124214 9138
rect 124600 9138 124684 9172
rect 124600 9132 124634 9138
rect 125020 9138 125104 9172
rect 125020 9132 125054 9138
rect 125440 9138 125524 9172
rect 125440 9132 125474 9138
rect 122290 8014 122374 8048
rect 122710 8048 122744 8056
rect 122710 8014 122794 8048
rect 123130 8048 123164 8056
rect 123130 8014 123214 8048
rect 123550 8048 123584 8056
rect 123550 8014 123634 8048
rect 123970 8048 124004 8056
rect 123970 8014 124054 8048
rect 124390 8048 124424 8056
rect 124390 8014 124474 8048
rect 124810 8048 124844 8056
rect 124810 8014 124894 8048
rect 125230 8048 125264 8056
rect 125230 8014 125314 8048
rect 125650 8048 125684 8056
rect 125650 8014 125734 8048
<< locali >>
rect 126642 28200 126786 28234
rect 135266 28200 135396 28234
rect 126642 28078 126676 28200
rect 135362 28106 135396 28200
rect 126914 28018 126930 28052
rect 127014 28018 127030 28052
rect 127334 28018 127350 28052
rect 127434 28018 127450 28052
rect 127754 28018 127770 28052
rect 127854 28018 127870 28052
rect 128174 28018 128190 28052
rect 128274 28018 128290 28052
rect 128594 28018 128610 28052
rect 128694 28018 128710 28052
rect 129014 28018 129030 28052
rect 129114 28018 129130 28052
rect 129434 28018 129450 28052
rect 129534 28018 129550 28052
rect 129854 28018 129870 28052
rect 129954 28018 129970 28052
rect 130274 28018 130290 28052
rect 130374 28018 130390 28052
rect 130694 28018 130710 28052
rect 130794 28018 130810 28052
rect 131114 28018 131130 28052
rect 131214 28018 131230 28052
rect 131534 28018 131550 28052
rect 131634 28018 131650 28052
rect 131954 28018 131970 28052
rect 132054 28018 132070 28052
rect 132374 28018 132390 28052
rect 132474 28018 132490 28052
rect 132794 28018 132810 28052
rect 132894 28018 132910 28052
rect 133214 28018 133230 28052
rect 133314 28018 133330 28052
rect 133634 28018 133650 28052
rect 133734 28018 133750 28052
rect 134054 28018 134070 28052
rect 134154 28018 134170 28052
rect 134474 28018 134490 28052
rect 134574 28018 134590 28052
rect 134894 28018 134910 28052
rect 134994 28018 135010 28052
rect 126882 27968 126916 27984
rect 126882 26976 126916 26992
rect 126978 27968 127012 27984
rect 126978 26976 127012 26992
rect 127092 27968 127126 27984
rect 127092 26976 127126 26992
rect 127188 27968 127222 27984
rect 127188 26976 127222 26992
rect 127302 27968 127336 27984
rect 127302 26976 127336 26992
rect 127398 27968 127432 27984
rect 127398 26976 127432 26992
rect 127512 27968 127546 27984
rect 127512 26976 127546 26992
rect 127608 27968 127642 27984
rect 127608 26976 127642 26992
rect 127722 27968 127756 27984
rect 127722 26976 127756 26992
rect 127818 27968 127852 27984
rect 127818 26976 127852 26992
rect 127932 27968 127966 27984
rect 127932 26976 127966 26992
rect 128028 27968 128062 27984
rect 128028 26976 128062 26992
rect 128142 27968 128176 27984
rect 128142 26976 128176 26992
rect 128238 27968 128272 27984
rect 128238 26976 128272 26992
rect 128352 27968 128386 27984
rect 128352 26976 128386 26992
rect 128448 27968 128482 27984
rect 128448 26976 128482 26992
rect 128562 27968 128596 27984
rect 128562 26976 128596 26992
rect 128658 27968 128692 27984
rect 128658 26976 128692 26992
rect 128772 27968 128806 27984
rect 128772 26976 128806 26992
rect 128868 27968 128902 27984
rect 128868 26976 128902 26992
rect 128982 27968 129016 27984
rect 128982 26976 129016 26992
rect 129078 27968 129112 27984
rect 129078 26976 129112 26992
rect 129192 27968 129226 27984
rect 129192 26976 129226 26992
rect 129288 27968 129322 27984
rect 129288 26976 129322 26992
rect 129402 27968 129436 27984
rect 129402 26976 129436 26992
rect 129498 27968 129532 27984
rect 129498 26976 129532 26992
rect 129612 27968 129646 27984
rect 129612 26976 129646 26992
rect 129708 27968 129742 27984
rect 129708 26976 129742 26992
rect 129822 27968 129856 27984
rect 129822 26976 129856 26992
rect 129918 27968 129952 27984
rect 129918 26976 129952 26992
rect 130032 27968 130066 27984
rect 130032 26976 130066 26992
rect 130128 27968 130162 27984
rect 130128 26976 130162 26992
rect 130242 27968 130276 27984
rect 130242 26976 130276 26992
rect 130338 27968 130372 27984
rect 130338 26976 130372 26992
rect 130452 27968 130486 27984
rect 130452 26976 130486 26992
rect 130548 27968 130582 27984
rect 130548 26976 130582 26992
rect 130662 27968 130696 27984
rect 130662 26976 130696 26992
rect 130758 27968 130792 27984
rect 130758 26976 130792 26992
rect 130872 27968 130906 27984
rect 130872 26976 130906 26992
rect 130968 27968 131002 27984
rect 130968 26976 131002 26992
rect 131082 27968 131116 27984
rect 131082 26976 131116 26992
rect 131178 27968 131212 27984
rect 131178 26976 131212 26992
rect 131292 27968 131326 27984
rect 131292 26976 131326 26992
rect 131388 27968 131422 27984
rect 131388 26976 131422 26992
rect 131502 27968 131536 27984
rect 131502 26976 131536 26992
rect 131598 27968 131632 27984
rect 131598 26976 131632 26992
rect 131712 27968 131746 27984
rect 131712 26976 131746 26992
rect 131808 27968 131842 27984
rect 131808 26976 131842 26992
rect 131922 27968 131956 27984
rect 131922 26976 131956 26992
rect 132018 27968 132052 27984
rect 132018 26976 132052 26992
rect 132132 27968 132166 27984
rect 132132 26976 132166 26992
rect 132228 27968 132262 27984
rect 132228 26976 132262 26992
rect 132342 27968 132376 27984
rect 132342 26976 132376 26992
rect 132438 27968 132472 27984
rect 132438 26976 132472 26992
rect 132552 27968 132586 27984
rect 132552 26976 132586 26992
rect 132648 27968 132682 27984
rect 132648 26976 132682 26992
rect 132762 27968 132796 27984
rect 132762 26976 132796 26992
rect 132858 27968 132892 27984
rect 132858 26976 132892 26992
rect 132972 27968 133006 27984
rect 132972 26976 133006 26992
rect 133068 27968 133102 27984
rect 133068 26976 133102 26992
rect 133182 27968 133216 27984
rect 133182 26976 133216 26992
rect 133278 27968 133312 27984
rect 133278 26976 133312 26992
rect 133392 27968 133426 27984
rect 133392 26976 133426 26992
rect 133488 27968 133522 27984
rect 133488 26976 133522 26992
rect 133602 27968 133636 27984
rect 133602 26976 133636 26992
rect 133698 27968 133732 27984
rect 133698 26976 133732 26992
rect 133812 27968 133846 27984
rect 133812 26976 133846 26992
rect 133908 27968 133942 27984
rect 133908 26976 133942 26992
rect 134022 27968 134056 27984
rect 134022 26976 134056 26992
rect 134118 27968 134152 27984
rect 134118 26976 134152 26992
rect 134232 27968 134266 27984
rect 134232 26976 134266 26992
rect 134328 27968 134362 27984
rect 134328 26976 134362 26992
rect 134442 27968 134476 27984
rect 134442 26976 134476 26992
rect 134538 27968 134572 27984
rect 134538 26976 134572 26992
rect 134652 27968 134686 27984
rect 134652 26976 134686 26992
rect 134748 27968 134782 27984
rect 134748 26976 134782 26992
rect 134862 27968 134896 27984
rect 134862 26976 134896 26992
rect 134958 27968 134992 27984
rect 134958 26976 134992 26992
rect 135072 27968 135106 27984
rect 135072 26976 135106 26992
rect 135168 27968 135202 27984
rect 135168 26976 135202 26992
rect 127124 26908 127140 26942
rect 127124 26800 127140 26834
rect 127174 26908 127190 26942
rect 127544 26908 127560 26942
rect 127174 26800 127190 26834
rect 127544 26800 127560 26834
rect 127594 26908 127610 26942
rect 127964 26908 127980 26942
rect 127594 26800 127610 26834
rect 127964 26800 127980 26834
rect 128014 26908 128030 26942
rect 128384 26908 128400 26942
rect 128014 26800 128030 26834
rect 128384 26800 128400 26834
rect 128434 26908 128450 26942
rect 128804 26908 128820 26942
rect 128434 26800 128450 26834
rect 128804 26800 128820 26834
rect 128854 26908 128870 26942
rect 129224 26908 129240 26942
rect 128854 26800 128870 26834
rect 129224 26800 129240 26834
rect 129274 26908 129290 26942
rect 129644 26908 129660 26942
rect 129274 26800 129290 26834
rect 129644 26800 129660 26834
rect 129694 26908 129710 26942
rect 130064 26908 130080 26942
rect 129694 26800 129710 26834
rect 130064 26800 130080 26834
rect 130114 26908 130130 26942
rect 130484 26908 130500 26942
rect 130114 26800 130130 26834
rect 130484 26800 130500 26834
rect 130534 26908 130550 26942
rect 130904 26908 130920 26942
rect 130534 26800 130550 26834
rect 130904 26800 130920 26834
rect 130954 26908 130970 26942
rect 131324 26908 131340 26942
rect 130954 26800 130970 26834
rect 131324 26800 131340 26834
rect 131374 26908 131390 26942
rect 131744 26908 131760 26942
rect 131374 26800 131390 26834
rect 131744 26800 131760 26834
rect 131794 26908 131810 26942
rect 132164 26908 132180 26942
rect 131794 26800 131810 26834
rect 132164 26800 132180 26834
rect 132214 26908 132230 26942
rect 132584 26908 132600 26942
rect 132214 26800 132230 26834
rect 132584 26800 132600 26834
rect 132634 26908 132650 26942
rect 133004 26908 133020 26942
rect 132634 26800 132650 26834
rect 133004 26800 133020 26834
rect 133054 26908 133070 26942
rect 133424 26908 133440 26942
rect 133054 26800 133070 26834
rect 133424 26800 133440 26834
rect 133474 26908 133490 26942
rect 133844 26908 133860 26942
rect 133474 26800 133490 26834
rect 133844 26800 133860 26834
rect 133894 26908 133910 26942
rect 134264 26908 134280 26942
rect 133894 26800 133910 26834
rect 134264 26800 134280 26834
rect 134314 26908 134330 26942
rect 134684 26908 134700 26942
rect 134314 26800 134330 26834
rect 134684 26800 134700 26834
rect 134734 26908 134750 26942
rect 135104 26908 135120 26942
rect 134734 26800 134750 26834
rect 135104 26800 135120 26834
rect 135154 26908 135170 26942
rect 135154 26800 135170 26834
rect 126882 26750 126916 26766
rect 126882 25758 126916 25774
rect 126978 26750 127012 26766
rect 126978 25758 127012 25774
rect 127092 26750 127126 26766
rect 127092 25758 127126 25774
rect 127188 26750 127222 26766
rect 127188 25758 127222 25774
rect 127302 26750 127336 26766
rect 127302 25758 127336 25774
rect 127398 26750 127432 26766
rect 127398 25758 127432 25774
rect 127512 26750 127546 26766
rect 127512 25758 127546 25774
rect 127608 26750 127642 26766
rect 127608 25758 127642 25774
rect 127722 26750 127756 26766
rect 127722 25758 127756 25774
rect 127818 26750 127852 26766
rect 127818 25758 127852 25774
rect 127932 26750 127966 26766
rect 127932 25758 127966 25774
rect 128028 26750 128062 26766
rect 128028 25758 128062 25774
rect 128142 26750 128176 26766
rect 128142 25758 128176 25774
rect 128238 26750 128272 26766
rect 128238 25758 128272 25774
rect 128352 26750 128386 26766
rect 128352 25758 128386 25774
rect 128448 26750 128482 26766
rect 128448 25758 128482 25774
rect 128562 26750 128596 26766
rect 128562 25758 128596 25774
rect 128658 26750 128692 26766
rect 128658 25758 128692 25774
rect 128772 26750 128806 26766
rect 128772 25758 128806 25774
rect 128868 26750 128902 26766
rect 128868 25758 128902 25774
rect 128982 26750 129016 26766
rect 128982 25758 129016 25774
rect 129078 26750 129112 26766
rect 129078 25758 129112 25774
rect 129192 26750 129226 26766
rect 129192 25758 129226 25774
rect 129288 26750 129322 26766
rect 129288 25758 129322 25774
rect 129402 26750 129436 26766
rect 129402 25758 129436 25774
rect 129498 26750 129532 26766
rect 129498 25758 129532 25774
rect 129612 26750 129646 26766
rect 129612 25758 129646 25774
rect 129708 26750 129742 26766
rect 129708 25758 129742 25774
rect 129822 26750 129856 26766
rect 129822 25758 129856 25774
rect 129918 26750 129952 26766
rect 129918 25758 129952 25774
rect 130032 26750 130066 26766
rect 130032 25758 130066 25774
rect 130128 26750 130162 26766
rect 130128 25758 130162 25774
rect 130242 26750 130276 26766
rect 130242 25758 130276 25774
rect 130338 26750 130372 26766
rect 130338 25758 130372 25774
rect 130452 26750 130486 26766
rect 130452 25758 130486 25774
rect 130548 26750 130582 26766
rect 130548 25758 130582 25774
rect 130662 26750 130696 26766
rect 130662 25758 130696 25774
rect 130758 26750 130792 26766
rect 130758 25758 130792 25774
rect 130872 26750 130906 26766
rect 130872 25758 130906 25774
rect 130968 26750 131002 26766
rect 130968 25758 131002 25774
rect 131082 26750 131116 26766
rect 131082 25758 131116 25774
rect 131178 26750 131212 26766
rect 131178 25758 131212 25774
rect 131292 26750 131326 26766
rect 131292 25758 131326 25774
rect 131388 26750 131422 26766
rect 131388 25758 131422 25774
rect 131502 26750 131536 26766
rect 131502 25758 131536 25774
rect 131598 26750 131632 26766
rect 131598 25758 131632 25774
rect 131712 26750 131746 26766
rect 131712 25758 131746 25774
rect 131808 26750 131842 26766
rect 131808 25758 131842 25774
rect 131922 26750 131956 26766
rect 131922 25758 131956 25774
rect 132018 26750 132052 26766
rect 132018 25758 132052 25774
rect 132132 26750 132166 26766
rect 132132 25758 132166 25774
rect 132228 26750 132262 26766
rect 132228 25758 132262 25774
rect 132342 26750 132376 26766
rect 132342 25758 132376 25774
rect 132438 26750 132472 26766
rect 132438 25758 132472 25774
rect 132552 26750 132586 26766
rect 132552 25758 132586 25774
rect 132648 26750 132682 26766
rect 132648 25758 132682 25774
rect 132762 26750 132796 26766
rect 132762 25758 132796 25774
rect 132858 26750 132892 26766
rect 132858 25758 132892 25774
rect 132972 26750 133006 26766
rect 132972 25758 133006 25774
rect 133068 26750 133102 26766
rect 133068 25758 133102 25774
rect 133182 26750 133216 26766
rect 133182 25758 133216 25774
rect 133278 26750 133312 26766
rect 133278 25758 133312 25774
rect 133392 26750 133426 26766
rect 133392 25758 133426 25774
rect 133488 26750 133522 26766
rect 133488 25758 133522 25774
rect 133602 26750 133636 26766
rect 133602 25758 133636 25774
rect 133698 26750 133732 26766
rect 133698 25758 133732 25774
rect 133812 26750 133846 26766
rect 133812 25758 133846 25774
rect 133908 26750 133942 26766
rect 133908 25758 133942 25774
rect 134022 26750 134056 26766
rect 134022 25758 134056 25774
rect 134118 26750 134152 26766
rect 134118 25758 134152 25774
rect 134232 26750 134266 26766
rect 134232 25758 134266 25774
rect 134328 26750 134362 26766
rect 134328 25758 134362 25774
rect 134442 26750 134476 26766
rect 134442 25758 134476 25774
rect 134538 26750 134572 26766
rect 134538 25758 134572 25774
rect 134652 26750 134686 26766
rect 134652 25758 134686 25774
rect 134748 26750 134782 26766
rect 134748 25758 134782 25774
rect 134862 26750 134896 26766
rect 134862 25758 134896 25774
rect 134958 26750 134992 26766
rect 134958 25758 134992 25774
rect 135072 26750 135106 26766
rect 135072 25758 135106 25774
rect 135168 26750 135202 26766
rect 135168 25758 135202 25774
rect 126642 25558 126676 25706
rect 126914 25690 126930 25724
rect 127014 25690 127030 25724
rect 127334 25690 127350 25724
rect 127434 25690 127450 25724
rect 127754 25690 127770 25724
rect 127854 25690 127870 25724
rect 128174 25690 128190 25724
rect 128274 25690 128290 25724
rect 128594 25690 128610 25724
rect 128694 25690 128710 25724
rect 129014 25690 129030 25724
rect 129114 25690 129130 25724
rect 129434 25690 129450 25724
rect 129534 25690 129550 25724
rect 129854 25690 129870 25724
rect 129954 25690 129970 25724
rect 130274 25690 130290 25724
rect 130374 25690 130390 25724
rect 130694 25690 130710 25724
rect 130794 25690 130810 25724
rect 131114 25690 131130 25724
rect 131214 25690 131230 25724
rect 131534 25690 131550 25724
rect 131634 25690 131650 25724
rect 131954 25690 131970 25724
rect 132054 25690 132070 25724
rect 132374 25690 132390 25724
rect 132474 25690 132490 25724
rect 132794 25690 132810 25724
rect 132894 25690 132910 25724
rect 133214 25690 133230 25724
rect 133314 25690 133330 25724
rect 133634 25690 133650 25724
rect 133734 25690 133750 25724
rect 134054 25690 134070 25724
rect 134154 25690 134170 25724
rect 134474 25690 134490 25724
rect 134574 25690 134590 25724
rect 134894 25690 134910 25724
rect 134994 25690 135010 25724
rect 135362 25558 135396 25694
rect 126642 25524 126798 25558
rect 135168 25524 135396 25558
rect 126670 22928 126896 22962
rect 135218 22928 135334 22962
rect 126670 22776 126704 22928
rect 126914 22833 126965 22838
rect 127334 22833 127385 22838
rect 127754 22833 127805 22838
rect 128174 22833 128225 22838
rect 128594 22833 128645 22838
rect 129014 22833 129065 22838
rect 129434 22833 129485 22838
rect 129854 22833 129905 22838
rect 130274 22833 130325 22838
rect 130694 22833 130745 22838
rect 131114 22833 131165 22838
rect 131534 22833 131585 22838
rect 131954 22833 132005 22838
rect 132374 22833 132425 22838
rect 132794 22833 132845 22838
rect 133214 22833 133265 22838
rect 133634 22833 133685 22838
rect 134054 22833 134105 22838
rect 134474 22833 134525 22838
rect 134894 22833 134945 22838
rect 126914 22798 126930 22833
rect 126964 22832 126980 22833
rect 127014 22798 127030 22832
rect 127334 22798 127350 22833
rect 127384 22832 127400 22833
rect 127434 22798 127450 22832
rect 127754 22798 127770 22833
rect 127804 22832 127820 22833
rect 127854 22798 127870 22832
rect 128174 22798 128190 22833
rect 128224 22832 128240 22833
rect 128274 22798 128290 22832
rect 128594 22798 128610 22833
rect 128644 22832 128660 22833
rect 128694 22798 128710 22832
rect 129014 22798 129030 22833
rect 129064 22832 129080 22833
rect 129114 22798 129130 22832
rect 129434 22798 129450 22833
rect 129484 22832 129500 22833
rect 129534 22798 129550 22832
rect 129854 22798 129870 22833
rect 129904 22832 129920 22833
rect 129954 22798 129970 22832
rect 130274 22798 130290 22833
rect 130324 22832 130340 22833
rect 130374 22798 130390 22832
rect 130694 22798 130710 22833
rect 130744 22832 130760 22833
rect 130794 22798 130810 22832
rect 131114 22798 131130 22833
rect 131164 22832 131180 22833
rect 131214 22798 131230 22832
rect 131534 22798 131550 22833
rect 131584 22832 131600 22833
rect 131634 22798 131650 22832
rect 131954 22798 131970 22833
rect 132004 22832 132020 22833
rect 132054 22798 132070 22832
rect 132374 22798 132390 22833
rect 132424 22832 132440 22833
rect 132474 22798 132490 22832
rect 132794 22798 132810 22833
rect 132844 22832 132860 22833
rect 132894 22798 132910 22832
rect 133214 22798 133230 22833
rect 133264 22832 133280 22833
rect 133314 22798 133330 22832
rect 133634 22798 133650 22833
rect 133684 22832 133700 22833
rect 133734 22798 133750 22832
rect 134054 22798 134070 22833
rect 134104 22832 134120 22833
rect 134154 22798 134170 22832
rect 134474 22798 134490 22833
rect 134524 22832 134540 22833
rect 134574 22798 134590 22832
rect 134894 22798 134910 22833
rect 134944 22832 134960 22833
rect 134994 22798 135010 22832
rect 126914 22790 126965 22798
rect 127334 22790 127385 22798
rect 127754 22790 127805 22798
rect 128174 22790 128225 22798
rect 128594 22790 128645 22798
rect 129014 22790 129065 22798
rect 129434 22790 129485 22798
rect 129854 22790 129905 22798
rect 130274 22790 130325 22798
rect 130694 22790 130745 22798
rect 131114 22790 131165 22798
rect 131534 22790 131585 22798
rect 131954 22790 132005 22798
rect 132374 22790 132425 22798
rect 132794 22790 132845 22798
rect 133214 22790 133265 22798
rect 133634 22790 133685 22798
rect 134054 22790 134105 22798
rect 134474 22790 134525 22798
rect 134894 22790 134945 22798
rect 121886 22028 122018 22062
rect 125742 22028 125848 22062
rect 121886 21912 121920 22028
rect 122274 21977 122325 21982
rect 122694 21977 122745 21982
rect 123114 21977 123165 21982
rect 123534 21977 123585 21982
rect 123954 21977 124005 21982
rect 124374 21977 124425 21982
rect 124794 21977 124845 21982
rect 125214 21977 125265 21982
rect 125634 21977 125685 21982
rect 122274 21976 122340 21977
rect 122694 21976 122760 21977
rect 123114 21976 123180 21977
rect 123534 21976 123600 21977
rect 123954 21976 124020 21977
rect 124374 21976 124440 21977
rect 124794 21976 124860 21977
rect 125214 21976 125280 21977
rect 125634 21976 125700 21977
rect 122274 21942 122290 21976
rect 122374 21942 122390 21976
rect 122274 21934 122325 21942
rect 122694 21934 122710 21976
rect 122794 21942 122810 21976
rect 122744 21934 122760 21942
rect 123114 21934 123130 21976
rect 123214 21942 123230 21976
rect 123164 21934 123180 21942
rect 123534 21934 123550 21976
rect 123634 21942 123650 21976
rect 123584 21934 123600 21942
rect 123954 21934 123970 21976
rect 124054 21942 124070 21976
rect 124004 21934 124020 21942
rect 124374 21934 124390 21976
rect 124474 21942 124490 21976
rect 124424 21934 124440 21942
rect 124794 21934 124810 21976
rect 124894 21942 124910 21976
rect 124844 21934 124860 21942
rect 125214 21934 125230 21976
rect 125314 21942 125330 21976
rect 125264 21934 125280 21942
rect 125634 21934 125650 21976
rect 125734 21942 125750 21976
rect 125684 21934 125700 21942
rect 125814 21936 125848 22028
rect 122032 21884 122066 21900
rect 122032 20892 122066 20908
rect 122128 21884 122162 21900
rect 122128 20892 122162 20908
rect 122242 21884 122276 21900
rect 122242 20892 122276 20908
rect 122338 21884 122372 21900
rect 122338 20892 122372 20908
rect 122452 21884 122486 21900
rect 122452 20892 122486 20908
rect 122548 21884 122582 21900
rect 122548 20892 122582 20908
rect 122662 21884 122696 21900
rect 122662 20892 122696 20908
rect 122758 21884 122792 21900
rect 122758 20892 122792 20908
rect 122872 21884 122906 21900
rect 122872 20892 122906 20908
rect 122968 21884 123002 21900
rect 122968 20892 123002 20908
rect 123082 21884 123116 21900
rect 123082 20892 123116 20908
rect 123178 21884 123212 21900
rect 123178 20892 123212 20908
rect 123292 21884 123326 21900
rect 123292 20892 123326 20908
rect 123388 21884 123422 21900
rect 123388 20892 123422 20908
rect 123502 21884 123536 21900
rect 123502 20892 123536 20908
rect 123598 21884 123632 21900
rect 123598 20892 123632 20908
rect 123712 21884 123746 21900
rect 123712 20892 123746 20908
rect 123808 21884 123842 21900
rect 123808 20892 123842 20908
rect 123922 21884 123956 21900
rect 123922 20892 123956 20908
rect 124018 21884 124052 21900
rect 124018 20892 124052 20908
rect 124132 21884 124166 21900
rect 124132 20892 124166 20908
rect 124228 21884 124262 21900
rect 124228 20892 124262 20908
rect 124342 21884 124376 21900
rect 124342 20892 124376 20908
rect 124438 21884 124472 21900
rect 124438 20892 124472 20908
rect 124552 21884 124586 21900
rect 124552 20892 124586 20908
rect 124648 21884 124682 21900
rect 124648 20892 124682 20908
rect 124762 21884 124796 21900
rect 124762 20892 124796 20908
rect 124858 21884 124892 21900
rect 124858 20892 124892 20908
rect 124972 21884 125006 21900
rect 124972 20892 125006 20908
rect 125068 21884 125102 21900
rect 125068 20892 125102 20908
rect 125182 21884 125216 21900
rect 125182 20892 125216 20908
rect 125278 21884 125312 21900
rect 125278 20892 125312 20908
rect 125392 21884 125426 21900
rect 125392 20892 125426 20908
rect 125488 21884 125522 21900
rect 125488 20892 125522 20908
rect 125602 21884 125636 21900
rect 125602 20892 125636 20908
rect 125698 21884 125732 21900
rect 125698 20892 125732 20908
rect 121886 20774 121920 20892
rect 122064 20853 122115 20858
rect 122484 20853 122535 20858
rect 122064 20818 122080 20853
rect 122114 20852 122130 20853
rect 122164 20818 122180 20852
rect 122484 20818 122500 20853
rect 122534 20852 122550 20853
rect 122584 20818 122600 20852
rect 122904 20818 122920 20858
rect 122954 20852 122970 20858
rect 123004 20818 123020 20852
rect 123324 20818 123340 20858
rect 123374 20852 123390 20858
rect 123424 20818 123440 20852
rect 123744 20818 123760 20858
rect 123794 20852 123810 20858
rect 123844 20818 123860 20852
rect 124164 20818 124180 20858
rect 124214 20852 124230 20858
rect 124264 20818 124280 20852
rect 124584 20818 124600 20858
rect 124634 20852 124650 20858
rect 124684 20818 124700 20852
rect 125004 20818 125020 20858
rect 125054 20852 125070 20858
rect 125104 20818 125120 20852
rect 125424 20818 125440 20858
rect 125474 20852 125490 20858
rect 125524 20818 125540 20852
rect 122064 20810 122115 20818
rect 122484 20810 122535 20818
rect 122904 20810 122955 20818
rect 123324 20810 123375 20818
rect 123744 20810 123795 20818
rect 124164 20810 124215 20818
rect 124584 20810 124635 20818
rect 125004 20810 125055 20818
rect 125424 20810 125475 20818
rect 125814 20774 125848 20894
rect 121886 20740 121978 20774
rect 125698 20740 125848 20774
rect 121922 20468 122052 20502
rect 125754 20468 125870 20502
rect 119124 20260 119158 20276
rect 119124 19268 119158 19284
rect 119212 20260 119246 20276
rect 119602 20166 119698 20448
rect 121922 20426 121956 20468
rect 120310 20353 120361 20358
rect 120730 20353 120781 20358
rect 120310 20318 120326 20353
rect 120360 20352 120376 20353
rect 120410 20318 120426 20352
rect 120730 20318 120746 20353
rect 120780 20352 120796 20353
rect 120830 20318 120846 20352
rect 120310 20310 120361 20318
rect 120730 20310 120781 20318
rect 120068 20260 120102 20276
rect 119538 20150 119744 20166
rect 119538 19442 119744 19458
rect 119212 19268 119246 19284
rect 120068 19268 120102 19284
rect 120164 20260 120198 20276
rect 120164 19268 120198 19284
rect 120278 20260 120312 20276
rect 120278 19268 120312 19284
rect 120374 20260 120408 20276
rect 120374 19268 120408 19284
rect 120488 20260 120522 20276
rect 120488 19268 120522 19284
rect 120584 20260 120618 20276
rect 120584 19268 120618 19284
rect 120698 20260 120732 20276
rect 120698 19268 120732 19284
rect 120794 20260 120828 20276
rect 120794 19268 120828 19284
rect 119152 19200 119168 19234
rect 119152 19091 119168 19125
rect 119202 19200 119218 19234
rect 120100 19200 120116 19234
rect 119202 19091 119218 19125
rect 120100 19091 120116 19125
rect 120150 19200 120166 19234
rect 120520 19200 120536 19234
rect 120150 19091 120166 19125
rect 120520 19091 120536 19125
rect 120570 19200 120586 19234
rect 120940 19125 120991 19130
rect 121360 19125 121411 19130
rect 120570 19091 120586 19125
rect 120940 19090 120956 19125
rect 120990 19124 121006 19125
rect 121040 19090 121056 19124
rect 121360 19090 121376 19125
rect 121410 19124 121426 19125
rect 121460 19090 121476 19124
rect 120940 19082 120991 19090
rect 121360 19082 121411 19090
rect 119120 19032 119154 19048
rect 119120 18040 119154 18056
rect 119216 19032 119250 19048
rect 119216 18040 119250 18056
rect 119312 19032 119346 19048
rect 119858 19032 119892 19048
rect 119462 18948 119668 18964
rect 119462 18240 119668 18256
rect 119312 18040 119346 18056
rect 119248 17998 119299 18004
rect 119248 17964 119264 17998
rect 119348 17964 119364 17998
rect 119248 17956 119299 17964
rect 119548 17770 119642 18240
rect 119858 18040 119892 18056
rect 119954 19032 119988 19048
rect 119954 18040 119988 18056
rect 120068 19032 120102 19048
rect 120068 18040 120102 18056
rect 120164 19032 120198 19048
rect 120164 18040 120198 18056
rect 120278 19032 120312 19048
rect 120278 18040 120312 18056
rect 120374 19032 120408 19048
rect 120374 18040 120408 18056
rect 120488 19032 120522 19048
rect 120488 18040 120522 18056
rect 120584 19032 120618 19048
rect 120584 18040 120618 18056
rect 120698 19032 120732 19048
rect 120698 18040 120732 18056
rect 120794 19032 120828 19048
rect 120794 18040 120828 18056
rect 120908 19032 120942 19048
rect 120908 18040 120942 18056
rect 121004 19032 121038 19048
rect 121004 18040 121038 18056
rect 121118 19032 121152 19048
rect 121118 18040 121152 18056
rect 121214 19032 121248 19048
rect 121214 18040 121248 18056
rect 121328 19032 121362 19048
rect 121328 18040 121362 18056
rect 121424 19032 121458 19048
rect 121424 18040 121458 18056
rect 119890 17997 119941 18002
rect 120310 17997 120361 18002
rect 120730 17997 120781 18002
rect 121150 17997 121201 18002
rect 119890 17962 119906 17997
rect 119940 17996 119956 17997
rect 119990 17962 120006 17996
rect 120310 17962 120326 17997
rect 120360 17996 120376 17997
rect 120410 17962 120426 17996
rect 120730 17962 120746 17997
rect 120780 17996 120796 17997
rect 120830 17962 120846 17996
rect 121150 17962 121166 17997
rect 121200 17996 121216 17997
rect 121250 17962 121266 17996
rect 119890 17954 119941 17962
rect 120310 17954 120361 17962
rect 120730 17954 120781 17962
rect 121150 17954 121201 17962
rect 122064 20361 122115 20366
rect 122484 20361 122535 20366
rect 122904 20361 122955 20366
rect 123324 20361 123375 20366
rect 123744 20361 123795 20366
rect 124164 20361 124215 20366
rect 124584 20361 124635 20366
rect 125004 20361 125055 20366
rect 125424 20361 125475 20366
rect 122064 20326 122080 20361
rect 122114 20360 122130 20361
rect 122164 20326 122180 20360
rect 122484 20326 122500 20361
rect 122534 20360 122550 20361
rect 122584 20326 122600 20360
rect 122904 20326 122920 20361
rect 122954 20360 122970 20361
rect 123004 20326 123020 20360
rect 123324 20326 123340 20361
rect 123374 20360 123390 20361
rect 123424 20326 123440 20360
rect 123744 20326 123760 20361
rect 123794 20360 123810 20361
rect 123844 20326 123860 20360
rect 124164 20326 124180 20361
rect 124214 20360 124230 20361
rect 124264 20326 124280 20360
rect 124584 20326 124600 20361
rect 124634 20360 124650 20361
rect 124684 20326 124700 20360
rect 125004 20326 125020 20361
rect 125054 20360 125070 20361
rect 125104 20326 125120 20360
rect 125424 20326 125440 20361
rect 125474 20360 125490 20361
rect 125524 20326 125540 20360
rect 122064 20318 122115 20326
rect 122484 20318 122535 20326
rect 122904 20318 122955 20326
rect 123324 20318 123375 20326
rect 123744 20318 123795 20326
rect 124164 20318 124215 20326
rect 124584 20318 124635 20326
rect 125004 20318 125055 20326
rect 125424 20318 125475 20326
rect 125836 20284 125870 20468
rect 122032 20268 122066 20284
rect 122032 19276 122066 19292
rect 122128 20268 122162 20284
rect 122128 19276 122162 19292
rect 122242 20268 122276 20284
rect 122242 19276 122276 19292
rect 122338 20268 122372 20284
rect 122338 19276 122372 19292
rect 122452 20268 122486 20284
rect 122452 19276 122486 19292
rect 122548 20268 122582 20284
rect 122548 19276 122582 19292
rect 122662 20268 122696 20284
rect 122662 19276 122696 19292
rect 122758 20268 122792 20284
rect 122758 19276 122792 19292
rect 122872 20268 122906 20284
rect 122872 19276 122906 19292
rect 122968 20268 123002 20284
rect 122968 19276 123002 19292
rect 123082 20268 123116 20284
rect 123082 19276 123116 19292
rect 123178 20268 123212 20284
rect 123178 19276 123212 19292
rect 123292 20268 123326 20284
rect 123292 19276 123326 19292
rect 123388 20268 123422 20284
rect 123388 19276 123422 19292
rect 123502 20268 123536 20284
rect 123502 19276 123536 19292
rect 123598 20268 123632 20284
rect 123598 19276 123632 19292
rect 123712 20268 123746 20284
rect 123712 19276 123746 19292
rect 123808 20268 123842 20284
rect 123808 19276 123842 19292
rect 123922 20268 123956 20284
rect 123922 19276 123956 19292
rect 124018 20268 124052 20284
rect 124018 19276 124052 19292
rect 124132 20268 124166 20284
rect 124132 19276 124166 19292
rect 124228 20268 124262 20284
rect 124228 19276 124262 19292
rect 124342 20268 124376 20284
rect 124342 19276 124376 19292
rect 124438 20268 124472 20284
rect 124438 19276 124472 19292
rect 124552 20268 124586 20284
rect 124552 19276 124586 19292
rect 124648 20268 124682 20284
rect 124648 19276 124682 19292
rect 124762 20268 124796 20284
rect 124762 19276 124796 19292
rect 124858 20268 124892 20284
rect 124858 19276 124892 19292
rect 124972 20268 125006 20284
rect 124972 19276 125006 19292
rect 125068 20268 125102 20284
rect 125068 19276 125102 19292
rect 125182 20268 125216 20284
rect 125182 19276 125216 19292
rect 125278 20268 125312 20284
rect 125278 19276 125312 19292
rect 125392 20268 125426 20284
rect 125392 19276 125426 19292
rect 125488 20268 125522 20284
rect 125488 19276 125522 19292
rect 125602 20268 125636 20284
rect 125602 19276 125636 19292
rect 125698 20268 125732 20284
rect 125698 19276 125732 19292
rect 122274 19199 122290 19233
rect 122274 19091 122290 19125
rect 122324 19199 122340 19233
rect 122694 19199 122710 19233
rect 122324 19091 122340 19125
rect 122694 19091 122710 19125
rect 122744 19199 122760 19233
rect 123114 19199 123130 19233
rect 122744 19091 122760 19125
rect 123114 19091 123130 19125
rect 123164 19199 123180 19233
rect 123534 19199 123550 19233
rect 123164 19091 123180 19125
rect 123534 19091 123550 19125
rect 123584 19199 123600 19233
rect 123954 19199 123970 19233
rect 123584 19091 123600 19125
rect 123954 19091 123970 19125
rect 124004 19199 124020 19233
rect 124374 19199 124390 19233
rect 124004 19091 124020 19125
rect 124374 19091 124390 19125
rect 124424 19199 124440 19233
rect 124794 19199 124810 19233
rect 124424 19091 124440 19125
rect 124794 19091 124810 19125
rect 124844 19199 124860 19233
rect 125214 19199 125230 19233
rect 124844 19091 124860 19125
rect 125214 19091 125230 19125
rect 125264 19199 125280 19233
rect 125634 19199 125650 19233
rect 125264 19091 125280 19125
rect 125634 19091 125650 19125
rect 125684 19199 125700 19233
rect 125684 19091 125700 19125
rect 122032 19032 122066 19048
rect 122032 18040 122066 18056
rect 122128 19032 122162 19048
rect 122128 18040 122162 18056
rect 122242 19032 122276 19048
rect 122242 18040 122276 18056
rect 122338 19032 122372 19048
rect 122338 18040 122372 18056
rect 122452 19032 122486 19048
rect 122452 18040 122486 18056
rect 122548 19032 122582 19048
rect 122548 18040 122582 18056
rect 122662 19032 122696 19048
rect 122662 18040 122696 18056
rect 122758 19032 122792 19048
rect 122758 18040 122792 18056
rect 122872 19032 122906 19048
rect 122872 18040 122906 18056
rect 122968 19032 123002 19048
rect 122968 18040 123002 18056
rect 123082 19032 123116 19048
rect 123082 18040 123116 18056
rect 123178 19032 123212 19048
rect 123178 18040 123212 18056
rect 123292 19032 123326 19048
rect 123292 18040 123326 18056
rect 123388 19032 123422 19048
rect 123388 18040 123422 18056
rect 123502 19032 123536 19048
rect 123502 18040 123536 18056
rect 123598 19032 123632 19048
rect 123598 18040 123632 18056
rect 123712 19032 123746 19048
rect 123712 18040 123746 18056
rect 123808 19032 123842 19048
rect 123808 18040 123842 18056
rect 123922 19032 123956 19048
rect 123922 18040 123956 18056
rect 124018 19032 124052 19048
rect 124018 18040 124052 18056
rect 124132 19032 124166 19048
rect 124132 18040 124166 18056
rect 124228 19032 124262 19048
rect 124228 18040 124262 18056
rect 124342 19032 124376 19048
rect 124342 18040 124376 18056
rect 124438 19032 124472 19048
rect 124438 18040 124472 18056
rect 124552 19032 124586 19048
rect 124552 18040 124586 18056
rect 124648 19032 124682 19048
rect 124648 18040 124682 18056
rect 124762 19032 124796 19048
rect 124762 18040 124796 18056
rect 124858 19032 124892 19048
rect 124858 18040 124892 18056
rect 124972 19032 125006 19048
rect 124972 18040 125006 18056
rect 125068 19032 125102 19048
rect 125068 18040 125102 18056
rect 125182 19032 125216 19048
rect 125182 18040 125216 18056
rect 125278 19032 125312 19048
rect 125278 18040 125312 18056
rect 125392 19032 125426 19048
rect 125392 18040 125426 18056
rect 125488 19032 125522 19048
rect 125488 18040 125522 18056
rect 125602 19032 125636 19048
rect 125602 18040 125636 18056
rect 125698 19032 125732 19048
rect 125698 18040 125732 18056
rect 121922 17902 121956 17958
rect 122064 17997 122115 18002
rect 122484 17997 122535 18002
rect 122904 17997 122955 18002
rect 123324 17997 123375 18002
rect 123744 17997 123795 18002
rect 124164 17997 124215 18002
rect 124584 17997 124635 18002
rect 125004 17997 125055 18002
rect 125424 17997 125475 18002
rect 122064 17962 122080 17997
rect 122114 17996 122130 17997
rect 122164 17962 122180 17996
rect 122484 17962 122500 17997
rect 122534 17996 122550 17997
rect 122584 17962 122600 17996
rect 122904 17962 122920 17997
rect 122954 17996 122970 17997
rect 123004 17962 123020 17996
rect 123324 17962 123340 17997
rect 123374 17996 123390 17997
rect 123424 17962 123440 17996
rect 123744 17962 123760 17997
rect 123794 17996 123810 17997
rect 123844 17962 123860 17996
rect 124164 17962 124180 17997
rect 124214 17996 124230 17997
rect 124264 17962 124280 17996
rect 124584 17962 124600 17997
rect 124634 17996 124650 17997
rect 124684 17962 124700 17996
rect 125004 17962 125020 17997
rect 125054 17996 125070 17997
rect 125104 17962 125120 17996
rect 125424 17962 125440 17997
rect 125474 17996 125490 17997
rect 125524 17962 125540 17996
rect 122064 17954 122115 17962
rect 122484 17954 122535 17962
rect 122904 17954 122955 17962
rect 123324 17954 123375 17962
rect 123744 17954 123795 17962
rect 124164 17954 124215 17962
rect 124584 17954 124635 17962
rect 125004 17954 125055 17962
rect 125424 17954 125475 17962
rect 125836 17870 125870 17996
rect 122004 17836 122024 17870
rect 125796 17836 125870 17870
rect 135300 22758 135334 22928
rect 126882 22740 126916 22756
rect 126882 21748 126916 21764
rect 126978 22740 127012 22756
rect 126978 21748 127012 21764
rect 127092 22740 127126 22756
rect 127092 21748 127126 21764
rect 127188 22740 127222 22756
rect 127188 21748 127222 21764
rect 127302 22740 127336 22756
rect 127302 21748 127336 21764
rect 127398 22740 127432 22756
rect 127398 21748 127432 21764
rect 127512 22740 127546 22756
rect 127512 21748 127546 21764
rect 127608 22740 127642 22756
rect 127608 21748 127642 21764
rect 127722 22740 127756 22756
rect 127722 21748 127756 21764
rect 127818 22740 127852 22756
rect 127818 21748 127852 21764
rect 127932 22740 127966 22756
rect 127932 21748 127966 21764
rect 128028 22740 128062 22756
rect 128028 21748 128062 21764
rect 128142 22740 128176 22756
rect 128142 21748 128176 21764
rect 128238 22740 128272 22756
rect 128238 21748 128272 21764
rect 128352 22740 128386 22756
rect 128352 21748 128386 21764
rect 128448 22740 128482 22756
rect 128448 21748 128482 21764
rect 128562 22740 128596 22756
rect 128562 21748 128596 21764
rect 128658 22740 128692 22756
rect 128658 21748 128692 21764
rect 128772 22740 128806 22756
rect 128772 21748 128806 21764
rect 128868 22740 128902 22756
rect 128868 21748 128902 21764
rect 128982 22740 129016 22756
rect 128982 21748 129016 21764
rect 129078 22740 129112 22756
rect 129078 21748 129112 21764
rect 129192 22740 129226 22756
rect 129192 21748 129226 21764
rect 129288 22740 129322 22756
rect 129288 21748 129322 21764
rect 129402 22740 129436 22756
rect 129402 21748 129436 21764
rect 129498 22740 129532 22756
rect 129498 21748 129532 21764
rect 129612 22740 129646 22756
rect 129612 21748 129646 21764
rect 129708 22740 129742 22756
rect 129708 21748 129742 21764
rect 129822 22740 129856 22756
rect 129822 21748 129856 21764
rect 129918 22740 129952 22756
rect 129918 21748 129952 21764
rect 130032 22740 130066 22756
rect 130032 21748 130066 21764
rect 130128 22740 130162 22756
rect 130128 21748 130162 21764
rect 130242 22740 130276 22756
rect 130242 21748 130276 21764
rect 130338 22740 130372 22756
rect 130338 21748 130372 21764
rect 130452 22740 130486 22756
rect 130452 21748 130486 21764
rect 130548 22740 130582 22756
rect 130548 21748 130582 21764
rect 130662 22740 130696 22756
rect 130662 21748 130696 21764
rect 130758 22740 130792 22756
rect 130758 21748 130792 21764
rect 130872 22740 130906 22756
rect 130872 21748 130906 21764
rect 130968 22740 131002 22756
rect 130968 21748 131002 21764
rect 131082 22740 131116 22756
rect 131082 21748 131116 21764
rect 131178 22740 131212 22756
rect 131178 21748 131212 21764
rect 131292 22740 131326 22756
rect 131292 21748 131326 21764
rect 131388 22740 131422 22756
rect 131388 21748 131422 21764
rect 131502 22740 131536 22756
rect 131502 21748 131536 21764
rect 131598 22740 131632 22756
rect 131598 21748 131632 21764
rect 131712 22740 131746 22756
rect 131712 21748 131746 21764
rect 131808 22740 131842 22756
rect 131808 21748 131842 21764
rect 131922 22740 131956 22756
rect 131922 21748 131956 21764
rect 132018 22740 132052 22756
rect 132018 21748 132052 21764
rect 132132 22740 132166 22756
rect 132132 21748 132166 21764
rect 132228 22740 132262 22756
rect 132228 21748 132262 21764
rect 132342 22740 132376 22756
rect 132342 21748 132376 21764
rect 132438 22740 132472 22756
rect 132438 21748 132472 21764
rect 132552 22740 132586 22756
rect 132552 21748 132586 21764
rect 132648 22740 132682 22756
rect 132648 21748 132682 21764
rect 132762 22740 132796 22756
rect 132762 21748 132796 21764
rect 132858 22740 132892 22756
rect 132858 21748 132892 21764
rect 132972 22740 133006 22756
rect 132972 21748 133006 21764
rect 133068 22740 133102 22756
rect 133068 21748 133102 21764
rect 133182 22740 133216 22756
rect 133182 21748 133216 21764
rect 133278 22740 133312 22756
rect 133278 21748 133312 21764
rect 133392 22740 133426 22756
rect 133392 21748 133426 21764
rect 133488 22740 133522 22756
rect 133488 21748 133522 21764
rect 133602 22740 133636 22756
rect 133602 21748 133636 21764
rect 133698 22740 133732 22756
rect 133698 21748 133732 21764
rect 133812 22740 133846 22756
rect 133812 21748 133846 21764
rect 133908 22740 133942 22756
rect 133908 21748 133942 21764
rect 134022 22740 134056 22756
rect 134022 21748 134056 21764
rect 134118 22740 134152 22756
rect 134118 21748 134152 21764
rect 134232 22740 134266 22756
rect 134232 21748 134266 21764
rect 134328 22740 134362 22756
rect 134328 21748 134362 21764
rect 134442 22740 134476 22756
rect 134442 21748 134476 21764
rect 134538 22740 134572 22756
rect 134538 21748 134572 21764
rect 134652 22740 134686 22756
rect 134652 21748 134686 21764
rect 134748 22740 134782 22756
rect 134748 21748 134782 21764
rect 134862 22740 134896 22756
rect 134862 21748 134896 21764
rect 134958 22740 134992 22756
rect 134958 21748 134992 21764
rect 135072 22740 135106 22756
rect 135072 21748 135106 21764
rect 135168 22740 135202 22756
rect 135168 21748 135202 21764
rect 127124 21671 127140 21705
rect 127124 21563 127140 21597
rect 127174 21671 127190 21705
rect 127544 21671 127560 21705
rect 127174 21563 127190 21597
rect 127544 21563 127560 21597
rect 127594 21671 127610 21705
rect 127964 21671 127980 21705
rect 127594 21563 127610 21597
rect 127964 21563 127980 21597
rect 128014 21671 128030 21705
rect 128384 21671 128400 21705
rect 128014 21563 128030 21597
rect 128384 21563 128400 21597
rect 128434 21671 128450 21705
rect 128804 21671 128820 21705
rect 128434 21563 128450 21597
rect 128804 21563 128820 21597
rect 128854 21671 128870 21705
rect 129224 21671 129240 21705
rect 128854 21563 128870 21597
rect 129224 21563 129240 21597
rect 129274 21671 129290 21705
rect 129644 21671 129660 21705
rect 129274 21563 129290 21597
rect 129644 21563 129660 21597
rect 129694 21671 129710 21705
rect 130064 21671 130080 21705
rect 129694 21563 129710 21597
rect 130064 21563 130080 21597
rect 130114 21671 130130 21705
rect 130484 21671 130500 21705
rect 130114 21563 130130 21597
rect 130484 21563 130500 21597
rect 130534 21671 130550 21705
rect 130904 21671 130920 21705
rect 130534 21563 130550 21597
rect 130904 21563 130920 21597
rect 130954 21671 130970 21705
rect 131324 21671 131340 21705
rect 130954 21563 130970 21597
rect 131324 21563 131340 21597
rect 131374 21671 131390 21705
rect 131744 21671 131760 21705
rect 131374 21563 131390 21597
rect 131744 21563 131760 21597
rect 131794 21671 131810 21705
rect 132164 21671 132180 21705
rect 131794 21563 131810 21597
rect 132164 21563 132180 21597
rect 132214 21671 132230 21705
rect 132584 21671 132600 21705
rect 132214 21563 132230 21597
rect 132584 21563 132600 21597
rect 132634 21671 132650 21705
rect 133004 21671 133020 21705
rect 132634 21563 132650 21597
rect 133004 21563 133020 21597
rect 133054 21671 133070 21705
rect 133424 21671 133440 21705
rect 133054 21563 133070 21597
rect 133424 21563 133440 21597
rect 133474 21671 133490 21705
rect 133844 21671 133860 21705
rect 133474 21563 133490 21597
rect 133844 21563 133860 21597
rect 133894 21671 133910 21705
rect 134264 21671 134280 21705
rect 133894 21563 133910 21597
rect 134264 21563 134280 21597
rect 134314 21671 134330 21705
rect 134684 21671 134700 21705
rect 134314 21563 134330 21597
rect 134684 21563 134700 21597
rect 134734 21671 134750 21705
rect 135104 21671 135120 21705
rect 134734 21563 134750 21597
rect 135104 21563 135120 21597
rect 135154 21671 135170 21705
rect 135154 21563 135170 21597
rect 126882 21504 126916 21520
rect 126882 20512 126916 20528
rect 126978 21504 127012 21520
rect 126978 20512 127012 20528
rect 127092 21504 127126 21520
rect 127092 20512 127126 20528
rect 127188 21504 127222 21520
rect 127188 20512 127222 20528
rect 127302 21504 127336 21520
rect 127302 20512 127336 20528
rect 127398 21504 127432 21520
rect 127398 20512 127432 20528
rect 127512 21504 127546 21520
rect 127512 20512 127546 20528
rect 127608 21504 127642 21520
rect 127608 20512 127642 20528
rect 127722 21504 127756 21520
rect 127722 20512 127756 20528
rect 127818 21504 127852 21520
rect 127818 20512 127852 20528
rect 127932 21504 127966 21520
rect 127932 20512 127966 20528
rect 128028 21504 128062 21520
rect 128028 20512 128062 20528
rect 128142 21504 128176 21520
rect 128142 20512 128176 20528
rect 128238 21504 128272 21520
rect 128238 20512 128272 20528
rect 128352 21504 128386 21520
rect 128352 20512 128386 20528
rect 128448 21504 128482 21520
rect 128448 20512 128482 20528
rect 128562 21504 128596 21520
rect 128562 20512 128596 20528
rect 128658 21504 128692 21520
rect 128658 20512 128692 20528
rect 128772 21504 128806 21520
rect 128772 20512 128806 20528
rect 128868 21504 128902 21520
rect 128868 20512 128902 20528
rect 128982 21504 129016 21520
rect 128982 20512 129016 20528
rect 129078 21504 129112 21520
rect 129078 20512 129112 20528
rect 129192 21504 129226 21520
rect 129192 20512 129226 20528
rect 129288 21504 129322 21520
rect 129288 20512 129322 20528
rect 129402 21504 129436 21520
rect 129402 20512 129436 20528
rect 129498 21504 129532 21520
rect 129498 20512 129532 20528
rect 129612 21504 129646 21520
rect 129612 20512 129646 20528
rect 129708 21504 129742 21520
rect 129708 20512 129742 20528
rect 129822 21504 129856 21520
rect 129822 20512 129856 20528
rect 129918 21504 129952 21520
rect 129918 20512 129952 20528
rect 130032 21504 130066 21520
rect 130032 20512 130066 20528
rect 130128 21504 130162 21520
rect 130128 20512 130162 20528
rect 130242 21504 130276 21520
rect 130242 20512 130276 20528
rect 130338 21504 130372 21520
rect 130338 20512 130372 20528
rect 130452 21504 130486 21520
rect 130452 20512 130486 20528
rect 130548 21504 130582 21520
rect 130548 20512 130582 20528
rect 130662 21504 130696 21520
rect 130662 20512 130696 20528
rect 130758 21504 130792 21520
rect 130758 20512 130792 20528
rect 130872 21504 130906 21520
rect 130872 20512 130906 20528
rect 130968 21504 131002 21520
rect 130968 20512 131002 20528
rect 131082 21504 131116 21520
rect 131082 20512 131116 20528
rect 131178 21504 131212 21520
rect 131178 20512 131212 20528
rect 131292 21504 131326 21520
rect 131292 20512 131326 20528
rect 131388 21504 131422 21520
rect 131388 20512 131422 20528
rect 131502 21504 131536 21520
rect 131502 20512 131536 20528
rect 131598 21504 131632 21520
rect 131598 20512 131632 20528
rect 131712 21504 131746 21520
rect 131712 20512 131746 20528
rect 131808 21504 131842 21520
rect 131808 20512 131842 20528
rect 131922 21504 131956 21520
rect 131922 20512 131956 20528
rect 132018 21504 132052 21520
rect 132018 20512 132052 20528
rect 132132 21504 132166 21520
rect 132132 20512 132166 20528
rect 132228 21504 132262 21520
rect 132228 20512 132262 20528
rect 132342 21504 132376 21520
rect 132342 20512 132376 20528
rect 132438 21504 132472 21520
rect 132438 20512 132472 20528
rect 132552 21504 132586 21520
rect 132552 20512 132586 20528
rect 132648 21504 132682 21520
rect 132648 20512 132682 20528
rect 132762 21504 132796 21520
rect 132762 20512 132796 20528
rect 132858 21504 132892 21520
rect 132858 20512 132892 20528
rect 132972 21504 133006 21520
rect 132972 20512 133006 20528
rect 133068 21504 133102 21520
rect 133068 20512 133102 20528
rect 133182 21504 133216 21520
rect 133182 20512 133216 20528
rect 133278 21504 133312 21520
rect 133278 20512 133312 20528
rect 133392 21504 133426 21520
rect 133392 20512 133426 20528
rect 133488 21504 133522 21520
rect 133488 20512 133522 20528
rect 133602 21504 133636 21520
rect 133602 20512 133636 20528
rect 133698 21504 133732 21520
rect 133698 20512 133732 20528
rect 133812 21504 133846 21520
rect 133812 20512 133846 20528
rect 133908 21504 133942 21520
rect 133908 20512 133942 20528
rect 134022 21504 134056 21520
rect 134022 20512 134056 20528
rect 134118 21504 134152 21520
rect 134118 20512 134152 20528
rect 134232 21504 134266 21520
rect 134232 20512 134266 20528
rect 134328 21504 134362 21520
rect 134328 20512 134362 20528
rect 134442 21504 134476 21520
rect 134442 20512 134476 20528
rect 134538 21504 134572 21520
rect 134538 20512 134572 20528
rect 134652 21504 134686 21520
rect 134652 20512 134686 20528
rect 134748 21504 134782 21520
rect 134748 20512 134782 20528
rect 134862 21504 134896 21520
rect 134862 20512 134896 20528
rect 134958 21504 134992 21520
rect 134958 20512 134992 20528
rect 135072 21504 135106 21520
rect 135072 20512 135106 20528
rect 135168 21504 135202 21520
rect 135168 20512 135202 20528
rect 126914 20435 126930 20469
rect 126914 20327 126930 20361
rect 126964 20435 126980 20469
rect 127334 20435 127350 20469
rect 126964 20327 126980 20361
rect 127334 20327 127350 20361
rect 127384 20435 127400 20469
rect 127754 20435 127770 20469
rect 127384 20327 127400 20361
rect 127754 20327 127770 20361
rect 127804 20435 127820 20469
rect 128174 20435 128190 20469
rect 127804 20327 127820 20361
rect 128174 20327 128190 20361
rect 128224 20435 128240 20469
rect 128594 20435 128610 20469
rect 128224 20327 128240 20361
rect 128594 20327 128610 20361
rect 128644 20435 128660 20469
rect 129014 20435 129030 20469
rect 128644 20327 128660 20361
rect 129014 20327 129030 20361
rect 129064 20435 129080 20469
rect 129434 20435 129450 20469
rect 129064 20327 129080 20361
rect 129434 20327 129450 20361
rect 129484 20435 129500 20469
rect 129854 20435 129870 20469
rect 129484 20327 129500 20361
rect 129854 20327 129870 20361
rect 129904 20435 129920 20469
rect 130274 20435 130290 20469
rect 129904 20327 129920 20361
rect 130274 20327 130290 20361
rect 130324 20435 130340 20469
rect 130694 20435 130710 20469
rect 130324 20327 130340 20361
rect 130694 20327 130710 20361
rect 130744 20435 130760 20469
rect 131114 20435 131130 20469
rect 130744 20327 130760 20361
rect 131114 20327 131130 20361
rect 131164 20435 131180 20469
rect 131534 20435 131550 20469
rect 131164 20327 131180 20361
rect 131534 20327 131550 20361
rect 131584 20435 131600 20469
rect 131954 20435 131970 20469
rect 131584 20327 131600 20361
rect 131954 20327 131970 20361
rect 132004 20435 132020 20469
rect 132374 20435 132390 20469
rect 132004 20327 132020 20361
rect 132374 20327 132390 20361
rect 132424 20435 132440 20469
rect 132794 20435 132810 20469
rect 132424 20327 132440 20361
rect 132794 20327 132810 20361
rect 132844 20435 132860 20469
rect 133214 20435 133230 20469
rect 132844 20327 132860 20361
rect 133214 20327 133230 20361
rect 133264 20435 133280 20469
rect 133634 20435 133650 20469
rect 133264 20327 133280 20361
rect 133634 20327 133650 20361
rect 133684 20435 133700 20469
rect 134054 20435 134070 20469
rect 133684 20327 133700 20361
rect 134054 20327 134070 20361
rect 134104 20435 134120 20469
rect 134474 20435 134490 20469
rect 134104 20327 134120 20361
rect 134474 20327 134490 20361
rect 134524 20435 134540 20469
rect 134894 20435 134910 20469
rect 134524 20327 134540 20361
rect 134894 20327 134910 20361
rect 134944 20435 134960 20469
rect 134944 20327 134960 20361
rect 126882 20268 126916 20284
rect 126882 19276 126916 19292
rect 126978 20268 127012 20284
rect 126978 19276 127012 19292
rect 127092 20268 127126 20284
rect 127092 19276 127126 19292
rect 127188 20268 127222 20284
rect 127188 19276 127222 19292
rect 127302 20268 127336 20284
rect 127302 19276 127336 19292
rect 127398 20268 127432 20284
rect 127398 19276 127432 19292
rect 127512 20268 127546 20284
rect 127512 19276 127546 19292
rect 127608 20268 127642 20284
rect 127608 19276 127642 19292
rect 127722 20268 127756 20284
rect 127722 19276 127756 19292
rect 127818 20268 127852 20284
rect 127818 19276 127852 19292
rect 127932 20268 127966 20284
rect 127932 19276 127966 19292
rect 128028 20268 128062 20284
rect 128028 19276 128062 19292
rect 128142 20268 128176 20284
rect 128142 19276 128176 19292
rect 128238 20268 128272 20284
rect 128238 19276 128272 19292
rect 128352 20268 128386 20284
rect 128352 19276 128386 19292
rect 128448 20268 128482 20284
rect 128448 19276 128482 19292
rect 128562 20268 128596 20284
rect 128562 19276 128596 19292
rect 128658 20268 128692 20284
rect 128658 19276 128692 19292
rect 128772 20268 128806 20284
rect 128772 19276 128806 19292
rect 128868 20268 128902 20284
rect 128868 19276 128902 19292
rect 128982 20268 129016 20284
rect 128982 19276 129016 19292
rect 129078 20268 129112 20284
rect 129078 19276 129112 19292
rect 129192 20268 129226 20284
rect 129192 19276 129226 19292
rect 129288 20268 129322 20284
rect 129288 19276 129322 19292
rect 129402 20268 129436 20284
rect 129402 19276 129436 19292
rect 129498 20268 129532 20284
rect 129498 19276 129532 19292
rect 129612 20268 129646 20284
rect 129612 19276 129646 19292
rect 129708 20268 129742 20284
rect 129708 19276 129742 19292
rect 129822 20268 129856 20284
rect 129822 19276 129856 19292
rect 129918 20268 129952 20284
rect 129918 19276 129952 19292
rect 130032 20268 130066 20284
rect 130032 19276 130066 19292
rect 130128 20268 130162 20284
rect 130128 19276 130162 19292
rect 130242 20268 130276 20284
rect 130242 19276 130276 19292
rect 130338 20268 130372 20284
rect 130338 19276 130372 19292
rect 130452 20268 130486 20284
rect 130452 19276 130486 19292
rect 130548 20268 130582 20284
rect 130548 19276 130582 19292
rect 130662 20268 130696 20284
rect 130662 19276 130696 19292
rect 130758 20268 130792 20284
rect 130758 19276 130792 19292
rect 130872 20268 130906 20284
rect 130872 19276 130906 19292
rect 130968 20268 131002 20284
rect 130968 19276 131002 19292
rect 131082 20268 131116 20284
rect 131082 19276 131116 19292
rect 131178 20268 131212 20284
rect 131178 19276 131212 19292
rect 131292 20268 131326 20284
rect 131292 19276 131326 19292
rect 131388 20268 131422 20284
rect 131388 19276 131422 19292
rect 131502 20268 131536 20284
rect 131502 19276 131536 19292
rect 131598 20268 131632 20284
rect 131598 19276 131632 19292
rect 131712 20268 131746 20284
rect 131712 19276 131746 19292
rect 131808 20268 131842 20284
rect 131808 19276 131842 19292
rect 131922 20268 131956 20284
rect 131922 19276 131956 19292
rect 132018 20268 132052 20284
rect 132018 19276 132052 19292
rect 132132 20268 132166 20284
rect 132132 19276 132166 19292
rect 132228 20268 132262 20284
rect 132228 19276 132262 19292
rect 132342 20268 132376 20284
rect 132342 19276 132376 19292
rect 132438 20268 132472 20284
rect 132438 19276 132472 19292
rect 132552 20268 132586 20284
rect 132552 19276 132586 19292
rect 132648 20268 132682 20284
rect 132648 19276 132682 19292
rect 132762 20268 132796 20284
rect 132762 19276 132796 19292
rect 132858 20268 132892 20284
rect 132858 19276 132892 19292
rect 132972 20268 133006 20284
rect 132972 19276 133006 19292
rect 133068 20268 133102 20284
rect 133068 19276 133102 19292
rect 133182 20268 133216 20284
rect 133182 19276 133216 19292
rect 133278 20268 133312 20284
rect 133278 19276 133312 19292
rect 133392 20268 133426 20284
rect 133392 19276 133426 19292
rect 133488 20268 133522 20284
rect 133488 19276 133522 19292
rect 133602 20268 133636 20284
rect 133602 19276 133636 19292
rect 133698 20268 133732 20284
rect 133698 19276 133732 19292
rect 133812 20268 133846 20284
rect 133812 19276 133846 19292
rect 133908 20268 133942 20284
rect 133908 19276 133942 19292
rect 134022 20268 134056 20284
rect 134022 19276 134056 19292
rect 134118 20268 134152 20284
rect 134118 19276 134152 19292
rect 134232 20268 134266 20284
rect 134232 19276 134266 19292
rect 134328 20268 134362 20284
rect 134328 19276 134362 19292
rect 134442 20268 134476 20284
rect 134442 19276 134476 19292
rect 134538 20268 134572 20284
rect 134538 19276 134572 19292
rect 134652 20268 134686 20284
rect 134652 19276 134686 19292
rect 134748 20268 134782 20284
rect 134748 19276 134782 19292
rect 134862 20268 134896 20284
rect 134862 19276 134896 19292
rect 134958 20268 134992 20284
rect 134958 19276 134992 19292
rect 135072 20268 135106 20284
rect 135072 19276 135106 19292
rect 135168 20268 135202 20284
rect 135168 19276 135202 19292
rect 127124 19199 127140 19233
rect 127124 19091 127140 19125
rect 127174 19199 127190 19233
rect 127544 19199 127560 19233
rect 127174 19091 127190 19125
rect 127544 19091 127560 19125
rect 127594 19199 127610 19233
rect 127964 19199 127980 19233
rect 127594 19091 127610 19125
rect 127964 19091 127980 19125
rect 128014 19199 128030 19233
rect 128384 19199 128400 19233
rect 128014 19091 128030 19125
rect 128384 19091 128400 19125
rect 128434 19199 128450 19233
rect 128804 19199 128820 19233
rect 128434 19091 128450 19125
rect 128804 19091 128820 19125
rect 128854 19199 128870 19233
rect 129224 19199 129240 19233
rect 128854 19091 128870 19125
rect 129224 19091 129240 19125
rect 129274 19199 129290 19233
rect 129644 19199 129660 19233
rect 129274 19091 129290 19125
rect 129644 19091 129660 19125
rect 129694 19199 129710 19233
rect 130064 19199 130080 19233
rect 129694 19091 129710 19125
rect 130064 19091 130080 19125
rect 130114 19199 130130 19233
rect 130484 19199 130500 19233
rect 130114 19091 130130 19125
rect 130484 19091 130500 19125
rect 130534 19199 130550 19233
rect 130904 19199 130920 19233
rect 130534 19091 130550 19125
rect 130904 19091 130920 19125
rect 130954 19199 130970 19233
rect 131324 19199 131340 19233
rect 130954 19091 130970 19125
rect 131324 19091 131340 19125
rect 131374 19199 131390 19233
rect 131744 19199 131760 19233
rect 131374 19091 131390 19125
rect 131744 19091 131760 19125
rect 131794 19199 131810 19233
rect 132164 19199 132180 19233
rect 131794 19091 131810 19125
rect 132164 19091 132180 19125
rect 132214 19199 132230 19233
rect 132584 19199 132600 19233
rect 132214 19091 132230 19125
rect 132584 19091 132600 19125
rect 132634 19199 132650 19233
rect 133004 19199 133020 19233
rect 132634 19091 132650 19125
rect 133004 19091 133020 19125
rect 133054 19199 133070 19233
rect 133424 19199 133440 19233
rect 133054 19091 133070 19125
rect 133424 19091 133440 19125
rect 133474 19199 133490 19233
rect 133844 19199 133860 19233
rect 133474 19091 133490 19125
rect 133844 19091 133860 19125
rect 133894 19199 133910 19233
rect 134264 19199 134280 19233
rect 133894 19091 133910 19125
rect 134264 19091 134280 19125
rect 134314 19199 134330 19233
rect 134684 19199 134700 19233
rect 134314 19091 134330 19125
rect 134684 19091 134700 19125
rect 134734 19199 134750 19233
rect 135104 19199 135120 19233
rect 134734 19091 134750 19125
rect 135104 19091 135120 19125
rect 135154 19199 135170 19233
rect 135154 19091 135170 19125
rect 126882 19032 126916 19048
rect 126882 18040 126916 18056
rect 126978 19032 127012 19048
rect 126978 18040 127012 18056
rect 127092 19032 127126 19048
rect 127092 18040 127126 18056
rect 127188 19032 127222 19048
rect 127188 18040 127222 18056
rect 127302 19032 127336 19048
rect 127302 18040 127336 18056
rect 127398 19032 127432 19048
rect 127398 18040 127432 18056
rect 127512 19032 127546 19048
rect 127512 18040 127546 18056
rect 127608 19032 127642 19048
rect 127608 18040 127642 18056
rect 127722 19032 127756 19048
rect 127722 18040 127756 18056
rect 127818 19032 127852 19048
rect 127818 18040 127852 18056
rect 127932 19032 127966 19048
rect 127932 18040 127966 18056
rect 128028 19032 128062 19048
rect 128028 18040 128062 18056
rect 128142 19032 128176 19048
rect 128142 18040 128176 18056
rect 128238 19032 128272 19048
rect 128238 18040 128272 18056
rect 128352 19032 128386 19048
rect 128352 18040 128386 18056
rect 128448 19032 128482 19048
rect 128448 18040 128482 18056
rect 128562 19032 128596 19048
rect 128562 18040 128596 18056
rect 128658 19032 128692 19048
rect 128658 18040 128692 18056
rect 128772 19032 128806 19048
rect 128772 18040 128806 18056
rect 128868 19032 128902 19048
rect 128868 18040 128902 18056
rect 128982 19032 129016 19048
rect 128982 18040 129016 18056
rect 129078 19032 129112 19048
rect 129078 18040 129112 18056
rect 129192 19032 129226 19048
rect 129192 18040 129226 18056
rect 129288 19032 129322 19048
rect 129288 18040 129322 18056
rect 129402 19032 129436 19048
rect 129402 18040 129436 18056
rect 129498 19032 129532 19048
rect 129498 18040 129532 18056
rect 129612 19032 129646 19048
rect 129612 18040 129646 18056
rect 129708 19032 129742 19048
rect 129708 18040 129742 18056
rect 129822 19032 129856 19048
rect 129822 18040 129856 18056
rect 129918 19032 129952 19048
rect 129918 18040 129952 18056
rect 130032 19032 130066 19048
rect 130032 18040 130066 18056
rect 130128 19032 130162 19048
rect 130128 18040 130162 18056
rect 130242 19032 130276 19048
rect 130242 18040 130276 18056
rect 130338 19032 130372 19048
rect 130338 18040 130372 18056
rect 130452 19032 130486 19048
rect 130452 18040 130486 18056
rect 130548 19032 130582 19048
rect 130548 18040 130582 18056
rect 130662 19032 130696 19048
rect 130662 18040 130696 18056
rect 130758 19032 130792 19048
rect 130758 18040 130792 18056
rect 130872 19032 130906 19048
rect 130872 18040 130906 18056
rect 130968 19032 131002 19048
rect 130968 18040 131002 18056
rect 131082 19032 131116 19048
rect 131082 18040 131116 18056
rect 131178 19032 131212 19048
rect 131178 18040 131212 18056
rect 131292 19032 131326 19048
rect 131292 18040 131326 18056
rect 131388 19032 131422 19048
rect 131388 18040 131422 18056
rect 131502 19032 131536 19048
rect 131502 18040 131536 18056
rect 131598 19032 131632 19048
rect 131598 18040 131632 18056
rect 131712 19032 131746 19048
rect 131712 18040 131746 18056
rect 131808 19032 131842 19048
rect 131808 18040 131842 18056
rect 131922 19032 131956 19048
rect 131922 18040 131956 18056
rect 132018 19032 132052 19048
rect 132018 18040 132052 18056
rect 132132 19032 132166 19048
rect 132132 18040 132166 18056
rect 132228 19032 132262 19048
rect 132228 18040 132262 18056
rect 132342 19032 132376 19048
rect 132342 18040 132376 18056
rect 132438 19032 132472 19048
rect 132438 18040 132472 18056
rect 132552 19032 132586 19048
rect 132552 18040 132586 18056
rect 132648 19032 132682 19048
rect 132648 18040 132682 18056
rect 132762 19032 132796 19048
rect 132762 18040 132796 18056
rect 132858 19032 132892 19048
rect 132858 18040 132892 18056
rect 132972 19032 133006 19048
rect 132972 18040 133006 18056
rect 133068 19032 133102 19048
rect 133068 18040 133102 18056
rect 133182 19032 133216 19048
rect 133182 18040 133216 18056
rect 133278 19032 133312 19048
rect 133278 18040 133312 18056
rect 133392 19032 133426 19048
rect 133392 18040 133426 18056
rect 133488 19032 133522 19048
rect 133488 18040 133522 18056
rect 133602 19032 133636 19048
rect 133602 18040 133636 18056
rect 133698 19032 133732 19048
rect 133698 18040 133732 18056
rect 133812 19032 133846 19048
rect 133812 18040 133846 18056
rect 133908 19032 133942 19048
rect 133908 18040 133942 18056
rect 134022 19032 134056 19048
rect 134022 18040 134056 18056
rect 134118 19032 134152 19048
rect 134118 18040 134152 18056
rect 134232 19032 134266 19048
rect 134232 18040 134266 18056
rect 134328 19032 134362 19048
rect 134328 18040 134362 18056
rect 134442 19032 134476 19048
rect 134442 18040 134476 18056
rect 134538 19032 134572 19048
rect 134538 18040 134572 18056
rect 134652 19032 134686 19048
rect 134652 18040 134686 18056
rect 134748 19032 134782 19048
rect 134748 18040 134782 18056
rect 134862 19032 134896 19048
rect 134862 18040 134896 18056
rect 134958 19032 134992 19048
rect 134958 18040 134992 18056
rect 135072 19032 135106 19048
rect 135072 18040 135106 18056
rect 135168 19032 135202 19048
rect 135168 18040 135202 18056
rect 126670 17854 126704 17978
rect 126914 17997 126965 18002
rect 127334 17997 127385 18002
rect 127754 17997 127805 18002
rect 128174 17997 128225 18002
rect 128594 17997 128645 18002
rect 129014 17997 129065 18002
rect 129434 17997 129485 18002
rect 129854 17997 129905 18002
rect 130274 17997 130325 18002
rect 130694 17997 130745 18002
rect 131114 17997 131165 18002
rect 131534 17997 131585 18002
rect 131954 17997 132005 18002
rect 132374 17997 132425 18002
rect 132794 17997 132845 18002
rect 133214 17997 133265 18002
rect 133634 17997 133685 18002
rect 134054 17997 134105 18002
rect 134474 17997 134525 18002
rect 134894 17997 134945 18002
rect 126914 17962 126930 17997
rect 126964 17996 126980 17997
rect 127014 17962 127030 17996
rect 127334 17962 127350 17997
rect 127384 17996 127400 17997
rect 127434 17962 127450 17996
rect 127754 17962 127770 17997
rect 127804 17996 127820 17997
rect 127854 17962 127870 17996
rect 128174 17962 128190 17997
rect 128224 17996 128240 17997
rect 128274 17962 128290 17996
rect 128594 17962 128610 17997
rect 128644 17996 128660 17997
rect 128694 17962 128710 17996
rect 129014 17962 129030 17997
rect 129064 17996 129080 17997
rect 129114 17962 129130 17996
rect 129434 17962 129450 17997
rect 129484 17996 129500 17997
rect 129534 17962 129550 17996
rect 129854 17962 129870 17997
rect 129904 17996 129920 17997
rect 129954 17962 129970 17996
rect 130274 17962 130290 17997
rect 130324 17996 130340 17997
rect 130374 17962 130390 17996
rect 130694 17962 130710 17997
rect 130744 17996 130760 17997
rect 130794 17962 130810 17996
rect 131114 17962 131130 17997
rect 131164 17996 131180 17997
rect 131214 17962 131230 17996
rect 131534 17962 131550 17997
rect 131584 17996 131600 17997
rect 131634 17962 131650 17996
rect 131954 17962 131970 17997
rect 132004 17996 132020 17997
rect 132054 17962 132070 17996
rect 132374 17962 132390 17997
rect 132424 17996 132440 17997
rect 132474 17962 132490 17996
rect 132794 17962 132810 17997
rect 132844 17996 132860 17997
rect 132894 17962 132910 17996
rect 133214 17962 133230 17997
rect 133264 17996 133280 17997
rect 133314 17962 133330 17996
rect 133634 17962 133650 17997
rect 133684 17996 133700 17997
rect 133734 17962 133750 17996
rect 134054 17962 134070 17997
rect 134104 17996 134120 17997
rect 134154 17962 134170 17996
rect 134474 17962 134490 17997
rect 134524 17996 134540 17997
rect 134574 17962 134590 17996
rect 134894 17962 134910 17997
rect 134944 17996 134960 17997
rect 134994 17962 135010 17996
rect 126914 17954 126965 17962
rect 127334 17954 127385 17962
rect 127754 17954 127805 17962
rect 128174 17954 128225 17962
rect 128594 17954 128645 17962
rect 129014 17954 129065 17962
rect 129434 17954 129485 17962
rect 129854 17954 129905 17962
rect 130274 17954 130325 17962
rect 130694 17954 130745 17962
rect 131114 17954 131165 17962
rect 131534 17954 131585 17962
rect 131954 17954 132005 17962
rect 132374 17954 132425 17962
rect 132794 17954 132845 17962
rect 133214 17954 133265 17962
rect 133634 17954 133685 17962
rect 134054 17954 134105 17962
rect 134474 17954 134525 17962
rect 134894 17954 134945 17962
rect 126670 17820 126746 17854
rect 135300 17854 135334 18040
rect 126846 17820 126860 17854
rect 135246 17820 135334 17854
rect 116382 16906 116416 16922
rect 116172 16830 116300 16846
rect 116172 16616 116190 16830
rect 116284 16616 116300 16830
rect 116172 16594 116300 16616
rect 116382 16514 116416 16530
rect 116470 16906 116510 16922
rect 116470 16530 116476 16906
rect 116470 16514 116510 16530
rect 116564 16906 116598 16922
rect 116564 16514 116598 16530
rect 116502 16430 116512 16464
rect 116586 16430 116592 16464
rect 116344 16344 116350 16378
rect 116424 16344 116434 16378
rect 116382 16286 116416 16302
rect 116190 16204 116304 16222
rect 116190 15998 116208 16204
rect 116284 15998 116304 16204
rect 116190 15976 116304 15998
rect 116382 15894 116416 15910
rect 116470 16286 116510 16302
rect 116470 15910 116476 16286
rect 116470 15894 116510 15910
rect 116564 16286 116598 16302
rect 116564 15894 116598 15910
rect 115856 15478 115890 15494
rect 115730 15438 115808 15458
rect 115730 15322 115750 15438
rect 115790 15322 115808 15438
rect 115730 15302 115808 15322
rect 115856 15086 115890 15102
rect 115944 15478 115978 15494
rect 116382 15480 116416 15496
rect 116190 15392 116304 15414
rect 116190 15186 116208 15392
rect 116284 15186 116304 15392
rect 116190 15168 116304 15186
rect 115944 15086 115978 15102
rect 116382 15088 116416 15104
rect 116470 15480 116510 15496
rect 116470 15104 116476 15480
rect 116470 15088 116510 15104
rect 116564 15480 116598 15496
rect 116564 15088 116598 15104
rect 115884 15009 115900 15043
rect 115934 15009 115950 15043
rect 116344 15012 116350 15046
rect 116424 15012 116434 15046
rect 116502 14926 116512 14960
rect 116586 14926 116592 14960
rect 115884 14872 115900 14906
rect 115934 14872 115950 14906
rect 116382 14860 116416 14876
rect 115708 14810 115806 14826
rect 115708 14668 115726 14810
rect 115790 14668 115806 14810
rect 115708 14652 115806 14668
rect 115856 14822 115890 14838
rect 115856 14630 115890 14646
rect 115944 14822 115978 14838
rect 115944 14630 115978 14646
rect 116172 14774 116300 14796
rect 116172 14560 116190 14774
rect 116284 14560 116300 14774
rect 116172 14544 116300 14560
rect 116382 14468 116416 14484
rect 116470 14860 116510 14876
rect 116470 14484 116476 14860
rect 116470 14468 116510 14484
rect 116564 14860 116598 14876
rect 116564 14468 116598 14484
rect 119248 13426 119299 13434
rect 119248 13392 119264 13426
rect 119348 13392 119364 13426
rect 119248 13386 119299 13392
rect 119120 13334 119154 13350
rect 119120 12342 119154 12358
rect 119216 13334 119250 13350
rect 119216 12342 119250 12358
rect 119312 13334 119346 13350
rect 119548 13150 119642 13620
rect 122004 13520 122024 13554
rect 125796 13520 125870 13554
rect 119890 13428 119941 13436
rect 120310 13428 120361 13436
rect 120730 13428 120781 13436
rect 121150 13428 121201 13436
rect 121922 13432 121956 13488
rect 119890 13393 119906 13428
rect 119990 13394 120006 13428
rect 119940 13393 119956 13394
rect 120310 13393 120326 13428
rect 120410 13394 120426 13428
rect 120360 13393 120376 13394
rect 120730 13393 120746 13428
rect 120830 13394 120846 13428
rect 120780 13393 120796 13394
rect 121150 13393 121166 13428
rect 121250 13394 121266 13428
rect 121200 13393 121216 13394
rect 119890 13388 119941 13393
rect 120310 13388 120361 13393
rect 120730 13388 120781 13393
rect 121150 13388 121201 13393
rect 119858 13334 119892 13350
rect 119462 13134 119668 13150
rect 119462 12426 119668 12442
rect 119312 12342 119346 12358
rect 119858 12342 119892 12358
rect 119954 13334 119988 13350
rect 119954 12342 119988 12358
rect 120068 13334 120102 13350
rect 120068 12342 120102 12358
rect 120164 13334 120198 13350
rect 120164 12342 120198 12358
rect 120278 13334 120312 13350
rect 120278 12342 120312 12358
rect 120374 13334 120408 13350
rect 120374 12342 120408 12358
rect 120488 13334 120522 13350
rect 120488 12342 120522 12358
rect 120584 13334 120618 13350
rect 120584 12342 120618 12358
rect 120698 13334 120732 13350
rect 120698 12342 120732 12358
rect 120794 13334 120828 13350
rect 120794 12342 120828 12358
rect 120908 13334 120942 13350
rect 120908 12342 120942 12358
rect 121004 13334 121038 13350
rect 121004 12342 121038 12358
rect 121118 13334 121152 13350
rect 121118 12342 121152 12358
rect 121214 13334 121248 13350
rect 121214 12342 121248 12358
rect 121328 13334 121362 13350
rect 121328 12342 121362 12358
rect 121424 13334 121458 13350
rect 121424 12342 121458 12358
rect 120940 12300 120991 12308
rect 121360 12300 121411 12308
rect 119152 12265 119168 12299
rect 119152 12156 119168 12190
rect 119202 12265 119218 12299
rect 120100 12265 120116 12299
rect 119202 12156 119218 12190
rect 120100 12156 120116 12190
rect 120150 12265 120166 12299
rect 120520 12265 120536 12299
rect 120150 12156 120166 12190
rect 120520 12156 120536 12190
rect 120570 12265 120586 12299
rect 120940 12265 120956 12300
rect 121040 12266 121056 12300
rect 120990 12265 121006 12266
rect 121360 12265 121376 12300
rect 121460 12266 121476 12300
rect 121410 12265 121426 12266
rect 120940 12260 120991 12265
rect 121360 12260 121411 12265
rect 120570 12156 120586 12190
rect 119124 12106 119158 12122
rect 119124 11114 119158 11130
rect 119212 12106 119246 12122
rect 120068 12106 120102 12122
rect 119538 11932 119744 11948
rect 119538 11224 119744 11240
rect 119212 11114 119246 11130
rect 119602 10942 119698 11224
rect 120068 11114 120102 11130
rect 120164 12106 120198 12122
rect 120164 11114 120198 11130
rect 120278 12106 120312 12122
rect 120278 11114 120312 11130
rect 120374 12106 120408 12122
rect 120374 11114 120408 11130
rect 120488 12106 120522 12122
rect 120488 11114 120522 11130
rect 120584 12106 120618 12122
rect 120584 11114 120618 11130
rect 120698 12106 120732 12122
rect 120698 11114 120732 11130
rect 120794 12106 120828 12122
rect 120794 11114 120828 11130
rect 120310 11072 120361 11080
rect 120730 11072 120781 11080
rect 120310 11037 120326 11072
rect 120410 11038 120426 11072
rect 120360 11037 120376 11038
rect 120730 11037 120746 11072
rect 120830 11038 120846 11072
rect 120780 11037 120796 11038
rect 120310 11032 120361 11037
rect 120730 11032 120781 11037
rect 122064 13428 122115 13436
rect 122484 13428 122535 13436
rect 122904 13428 122955 13436
rect 123324 13428 123375 13436
rect 123744 13428 123795 13436
rect 124164 13428 124215 13436
rect 124584 13428 124635 13436
rect 125004 13428 125055 13436
rect 125424 13428 125475 13436
rect 122064 13393 122080 13428
rect 122164 13394 122180 13428
rect 122114 13393 122130 13394
rect 122484 13393 122500 13428
rect 122584 13394 122600 13428
rect 122534 13393 122550 13394
rect 122904 13393 122920 13428
rect 123004 13394 123020 13428
rect 122954 13393 122970 13394
rect 123324 13393 123340 13428
rect 123424 13394 123440 13428
rect 123374 13393 123390 13394
rect 123744 13393 123760 13428
rect 123844 13394 123860 13428
rect 123794 13393 123810 13394
rect 124164 13393 124180 13428
rect 124264 13394 124280 13428
rect 124214 13393 124230 13394
rect 124584 13393 124600 13428
rect 124684 13394 124700 13428
rect 124634 13393 124650 13394
rect 125004 13393 125020 13428
rect 125104 13394 125120 13428
rect 125054 13393 125070 13394
rect 125424 13393 125440 13428
rect 125524 13394 125540 13428
rect 125836 13394 125870 13520
rect 125474 13393 125490 13394
rect 122064 13388 122115 13393
rect 122484 13388 122535 13393
rect 122904 13388 122955 13393
rect 123324 13388 123375 13393
rect 123744 13388 123795 13393
rect 124164 13388 124215 13393
rect 124584 13388 124635 13393
rect 125004 13388 125055 13393
rect 125424 13388 125475 13393
rect 122032 13334 122066 13350
rect 122032 12342 122066 12358
rect 122128 13334 122162 13350
rect 122128 12342 122162 12358
rect 122242 13334 122276 13350
rect 122242 12342 122276 12358
rect 122338 13334 122372 13350
rect 122338 12342 122372 12358
rect 122452 13334 122486 13350
rect 122452 12342 122486 12358
rect 122548 13334 122582 13350
rect 122548 12342 122582 12358
rect 122662 13334 122696 13350
rect 122662 12342 122696 12358
rect 122758 13334 122792 13350
rect 122758 12342 122792 12358
rect 122872 13334 122906 13350
rect 122872 12342 122906 12358
rect 122968 13334 123002 13350
rect 122968 12342 123002 12358
rect 123082 13334 123116 13350
rect 123082 12342 123116 12358
rect 123178 13334 123212 13350
rect 123178 12342 123212 12358
rect 123292 13334 123326 13350
rect 123292 12342 123326 12358
rect 123388 13334 123422 13350
rect 123388 12342 123422 12358
rect 123502 13334 123536 13350
rect 123502 12342 123536 12358
rect 123598 13334 123632 13350
rect 123598 12342 123632 12358
rect 123712 13334 123746 13350
rect 123712 12342 123746 12358
rect 123808 13334 123842 13350
rect 123808 12342 123842 12358
rect 123922 13334 123956 13350
rect 123922 12342 123956 12358
rect 124018 13334 124052 13350
rect 124018 12342 124052 12358
rect 124132 13334 124166 13350
rect 124132 12342 124166 12358
rect 124228 13334 124262 13350
rect 124228 12342 124262 12358
rect 124342 13334 124376 13350
rect 124342 12342 124376 12358
rect 124438 13334 124472 13350
rect 124438 12342 124472 12358
rect 124552 13334 124586 13350
rect 124552 12342 124586 12358
rect 124648 13334 124682 13350
rect 124648 12342 124682 12358
rect 124762 13334 124796 13350
rect 124762 12342 124796 12358
rect 124858 13334 124892 13350
rect 124858 12342 124892 12358
rect 124972 13334 125006 13350
rect 124972 12342 125006 12358
rect 125068 13334 125102 13350
rect 125068 12342 125102 12358
rect 125182 13334 125216 13350
rect 125182 12342 125216 12358
rect 125278 13334 125312 13350
rect 125278 12342 125312 12358
rect 125392 13334 125426 13350
rect 125392 12342 125426 12358
rect 125488 13334 125522 13350
rect 125488 12342 125522 12358
rect 125602 13334 125636 13350
rect 125602 12342 125636 12358
rect 125698 13334 125732 13350
rect 125698 12342 125732 12358
rect 122274 12265 122290 12299
rect 122274 12157 122290 12191
rect 122324 12265 122340 12299
rect 122694 12265 122710 12299
rect 122324 12157 122340 12191
rect 122694 12157 122710 12191
rect 122744 12265 122760 12299
rect 123114 12265 123130 12299
rect 122744 12157 122760 12191
rect 123114 12157 123130 12191
rect 123164 12265 123180 12299
rect 123534 12265 123550 12299
rect 123164 12157 123180 12191
rect 123534 12157 123550 12191
rect 123584 12265 123600 12299
rect 123954 12265 123970 12299
rect 123584 12157 123600 12191
rect 123954 12157 123970 12191
rect 124004 12265 124020 12299
rect 124374 12265 124390 12299
rect 124004 12157 124020 12191
rect 124374 12157 124390 12191
rect 124424 12265 124440 12299
rect 124794 12265 124810 12299
rect 124424 12157 124440 12191
rect 124794 12157 124810 12191
rect 124844 12265 124860 12299
rect 125214 12265 125230 12299
rect 124844 12157 124860 12191
rect 125214 12157 125230 12191
rect 125264 12265 125280 12299
rect 125634 12265 125650 12299
rect 125264 12157 125280 12191
rect 125634 12157 125650 12191
rect 125684 12265 125700 12299
rect 125684 12157 125700 12191
rect 122032 12098 122066 12114
rect 122032 11106 122066 11122
rect 122128 12098 122162 12114
rect 122128 11106 122162 11122
rect 122242 12098 122276 12114
rect 122242 11106 122276 11122
rect 122338 12098 122372 12114
rect 122338 11106 122372 11122
rect 122452 12098 122486 12114
rect 122452 11106 122486 11122
rect 122548 12098 122582 12114
rect 122548 11106 122582 11122
rect 122662 12098 122696 12114
rect 122662 11106 122696 11122
rect 122758 12098 122792 12114
rect 122758 11106 122792 11122
rect 122872 12098 122906 12114
rect 122872 11106 122906 11122
rect 122968 12098 123002 12114
rect 122968 11106 123002 11122
rect 123082 12098 123116 12114
rect 123082 11106 123116 11122
rect 123178 12098 123212 12114
rect 123178 11106 123212 11122
rect 123292 12098 123326 12114
rect 123292 11106 123326 11122
rect 123388 12098 123422 12114
rect 123388 11106 123422 11122
rect 123502 12098 123536 12114
rect 123502 11106 123536 11122
rect 123598 12098 123632 12114
rect 123598 11106 123632 11122
rect 123712 12098 123746 12114
rect 123712 11106 123746 11122
rect 123808 12098 123842 12114
rect 123808 11106 123842 11122
rect 123922 12098 123956 12114
rect 123922 11106 123956 11122
rect 124018 12098 124052 12114
rect 124018 11106 124052 11122
rect 124132 12098 124166 12114
rect 124132 11106 124166 11122
rect 124228 12098 124262 12114
rect 124228 11106 124262 11122
rect 124342 12098 124376 12114
rect 124342 11106 124376 11122
rect 124438 12098 124472 12114
rect 124438 11106 124472 11122
rect 124552 12098 124586 12114
rect 124552 11106 124586 11122
rect 124648 12098 124682 12114
rect 124648 11106 124682 11122
rect 124762 12098 124796 12114
rect 124762 11106 124796 11122
rect 124858 12098 124892 12114
rect 124858 11106 124892 11122
rect 124972 12098 125006 12114
rect 124972 11106 125006 11122
rect 125068 12098 125102 12114
rect 125068 11106 125102 11122
rect 125182 12098 125216 12114
rect 125182 11106 125216 11122
rect 125278 12098 125312 12114
rect 125278 11106 125312 11122
rect 125392 12098 125426 12114
rect 125392 11106 125426 11122
rect 125488 12098 125522 12114
rect 125488 11106 125522 11122
rect 125602 12098 125636 12114
rect 125602 11106 125636 11122
rect 125698 12098 125732 12114
rect 125698 11106 125732 11122
rect 122064 11064 122115 11072
rect 122484 11064 122535 11072
rect 122904 11064 122955 11072
rect 123324 11064 123375 11072
rect 123744 11064 123795 11072
rect 124164 11064 124215 11072
rect 124584 11064 124635 11072
rect 125004 11064 125055 11072
rect 125424 11064 125475 11072
rect 122064 11029 122080 11064
rect 122164 11030 122180 11064
rect 122114 11029 122130 11030
rect 122484 11029 122500 11064
rect 122584 11030 122600 11064
rect 122534 11029 122550 11030
rect 122904 11029 122920 11064
rect 123004 11030 123020 11064
rect 122954 11029 122970 11030
rect 123324 11029 123340 11064
rect 123424 11030 123440 11064
rect 123374 11029 123390 11030
rect 123744 11029 123760 11064
rect 123844 11030 123860 11064
rect 123794 11029 123810 11030
rect 124164 11029 124180 11064
rect 124264 11030 124280 11064
rect 124214 11029 124230 11030
rect 124584 11029 124600 11064
rect 124684 11030 124700 11064
rect 124634 11029 124650 11030
rect 125004 11029 125020 11064
rect 125104 11030 125120 11064
rect 125054 11029 125070 11030
rect 125424 11029 125440 11064
rect 125524 11030 125540 11064
rect 125474 11029 125490 11030
rect 122064 11024 122115 11029
rect 122484 11024 122535 11029
rect 122904 11024 122955 11029
rect 123324 11024 123375 11029
rect 123744 11024 123795 11029
rect 124164 11024 124215 11029
rect 124584 11024 124635 11029
rect 125004 11024 125055 11029
rect 125424 11024 125475 11029
rect 121922 10922 121956 10964
rect 125836 10922 125870 11106
rect 121922 10888 122052 10922
rect 125754 10888 125870 10922
rect 121886 9216 121978 9250
rect 125698 9216 125848 9250
rect 121886 9098 121920 9216
rect 122064 9172 122115 9180
rect 122484 9172 122535 9180
rect 122904 9172 122955 9180
rect 123324 9172 123375 9180
rect 123744 9172 123795 9180
rect 124164 9172 124215 9180
rect 124584 9172 124635 9180
rect 125004 9172 125055 9180
rect 125424 9172 125475 9180
rect 122064 9137 122080 9172
rect 122164 9138 122180 9172
rect 122114 9137 122130 9138
rect 122484 9137 122500 9172
rect 122584 9138 122600 9172
rect 122534 9137 122550 9138
rect 122064 9132 122115 9137
rect 122484 9132 122535 9137
rect 122904 9132 122920 9172
rect 123004 9138 123020 9172
rect 122954 9132 122970 9138
rect 123324 9132 123340 9172
rect 123424 9138 123440 9172
rect 123374 9132 123390 9138
rect 123744 9132 123760 9172
rect 123844 9138 123860 9172
rect 123794 9132 123810 9138
rect 124164 9132 124180 9172
rect 124264 9138 124280 9172
rect 124214 9132 124230 9138
rect 124584 9132 124600 9172
rect 124684 9138 124700 9172
rect 124634 9132 124650 9138
rect 125004 9132 125020 9172
rect 125104 9138 125120 9172
rect 125054 9132 125070 9138
rect 125424 9132 125440 9172
rect 125524 9138 125540 9172
rect 125474 9132 125490 9138
rect 122032 9082 122066 9098
rect 122032 8090 122066 8106
rect 122128 9082 122162 9098
rect 122128 8090 122162 8106
rect 122242 9082 122276 9098
rect 122242 8090 122276 8106
rect 122338 9082 122372 9098
rect 122338 8090 122372 8106
rect 122452 9082 122486 9098
rect 122452 8090 122486 8106
rect 122548 9082 122582 9098
rect 122548 8090 122582 8106
rect 122662 9082 122696 9098
rect 122662 8090 122696 8106
rect 122758 9082 122792 9098
rect 122758 8090 122792 8106
rect 122872 9082 122906 9098
rect 122872 8090 122906 8106
rect 122968 9082 123002 9098
rect 122968 8090 123002 8106
rect 123082 9082 123116 9098
rect 123082 8090 123116 8106
rect 123178 9082 123212 9098
rect 123178 8090 123212 8106
rect 123292 9082 123326 9098
rect 123292 8090 123326 8106
rect 123388 9082 123422 9098
rect 123388 8090 123422 8106
rect 123502 9082 123536 9098
rect 123502 8090 123536 8106
rect 123598 9082 123632 9098
rect 123598 8090 123632 8106
rect 123712 9082 123746 9098
rect 123712 8090 123746 8106
rect 123808 9082 123842 9098
rect 123808 8090 123842 8106
rect 123922 9082 123956 9098
rect 123922 8090 123956 8106
rect 124018 9082 124052 9098
rect 124018 8090 124052 8106
rect 124132 9082 124166 9098
rect 124132 8090 124166 8106
rect 124228 9082 124262 9098
rect 124228 8090 124262 8106
rect 124342 9082 124376 9098
rect 124342 8090 124376 8106
rect 124438 9082 124472 9098
rect 124438 8090 124472 8106
rect 124552 9082 124586 9098
rect 124552 8090 124586 8106
rect 124648 9082 124682 9098
rect 124648 8090 124682 8106
rect 124762 9082 124796 9098
rect 124762 8090 124796 8106
rect 124858 9082 124892 9098
rect 124858 8090 124892 8106
rect 124972 9082 125006 9098
rect 124972 8090 125006 8106
rect 125068 9082 125102 9098
rect 125068 8090 125102 8106
rect 125182 9082 125216 9098
rect 125182 8090 125216 8106
rect 125278 9082 125312 9098
rect 125278 8090 125312 8106
rect 125392 9082 125426 9098
rect 125392 8090 125426 8106
rect 125488 9082 125522 9098
rect 125488 8090 125522 8106
rect 125602 9082 125636 9098
rect 125602 8090 125636 8106
rect 125698 9082 125732 9098
rect 125698 8090 125732 8106
rect 125814 9096 125848 9216
rect 121886 7962 121920 8078
rect 122274 8048 122325 8056
rect 122274 8014 122290 8048
rect 122374 8014 122390 8048
rect 122694 8014 122710 8056
rect 122744 8048 122760 8056
rect 122794 8014 122810 8048
rect 123114 8014 123130 8056
rect 123164 8048 123180 8056
rect 123214 8014 123230 8048
rect 123534 8014 123550 8056
rect 123584 8048 123600 8056
rect 123634 8014 123650 8048
rect 123954 8014 123970 8056
rect 124004 8048 124020 8056
rect 124054 8014 124070 8048
rect 124374 8014 124390 8056
rect 124424 8048 124440 8056
rect 124474 8014 124490 8048
rect 124794 8014 124810 8056
rect 124844 8048 124860 8056
rect 124894 8014 124910 8048
rect 125214 8014 125230 8056
rect 125264 8048 125280 8056
rect 125314 8014 125330 8048
rect 125634 8014 125650 8056
rect 125684 8048 125700 8056
rect 125734 8014 125750 8048
rect 122274 8013 122340 8014
rect 122694 8013 122760 8014
rect 123114 8013 123180 8014
rect 123534 8013 123600 8014
rect 123954 8013 124020 8014
rect 124374 8013 124440 8014
rect 124794 8013 124860 8014
rect 125214 8013 125280 8014
rect 125634 8013 125700 8014
rect 122274 8008 122325 8013
rect 122694 8008 122745 8013
rect 123114 8008 123165 8013
rect 123534 8008 123585 8013
rect 123954 8008 124005 8013
rect 124374 8008 124425 8013
rect 124794 8008 124845 8013
rect 125214 8008 125265 8013
rect 125634 8008 125685 8013
rect 125814 7962 125848 8054
rect 121886 7928 122018 7962
rect 125742 7928 125848 7962
<< viali >>
rect 126840 28234 126938 28304
rect 127260 28234 127358 28304
rect 127680 28234 127778 28304
rect 128100 28234 128198 28304
rect 128520 28234 128618 28304
rect 128940 28234 129038 28304
rect 129360 28234 129458 28304
rect 129780 28234 129878 28304
rect 130200 28234 130298 28304
rect 130620 28234 130718 28304
rect 131040 28234 131138 28304
rect 131460 28234 131558 28304
rect 131880 28234 131978 28304
rect 132300 28234 132398 28304
rect 132720 28234 132818 28304
rect 133140 28234 133238 28304
rect 133560 28234 133658 28304
rect 133980 28234 134078 28304
rect 134400 28234 134498 28304
rect 134820 28234 134918 28304
rect 135168 28234 135266 28304
rect 126840 28200 126938 28234
rect 127260 28200 127358 28234
rect 127680 28200 127778 28234
rect 128100 28200 128198 28234
rect 128520 28200 128618 28234
rect 128940 28200 129038 28234
rect 129360 28200 129458 28234
rect 129780 28200 129878 28234
rect 130200 28200 130298 28234
rect 130620 28200 130718 28234
rect 131040 28200 131138 28234
rect 131460 28200 131558 28234
rect 131880 28200 131978 28234
rect 132300 28200 132398 28234
rect 132720 28200 132818 28234
rect 133140 28200 133238 28234
rect 133560 28200 133658 28234
rect 133980 28200 134078 28234
rect 134400 28200 134498 28234
rect 134820 28200 134918 28234
rect 135168 28200 135210 28234
rect 135210 28200 135266 28234
rect 126930 28018 127014 28052
rect 127350 28018 127434 28052
rect 127770 28018 127854 28052
rect 128190 28018 128274 28052
rect 128610 28018 128694 28052
rect 129030 28018 129114 28052
rect 129450 28018 129534 28052
rect 129870 28018 129954 28052
rect 130290 28018 130374 28052
rect 130710 28018 130794 28052
rect 131130 28018 131214 28052
rect 131550 28018 131634 28052
rect 131970 28018 132054 28052
rect 132390 28018 132474 28052
rect 132810 28018 132894 28052
rect 133230 28018 133314 28052
rect 133650 28018 133734 28052
rect 134070 28018 134154 28052
rect 134490 28018 134574 28052
rect 134910 28018 134994 28052
rect 126882 26992 126916 27968
rect 126978 26992 127012 27968
rect 127092 26992 127126 27968
rect 127188 26992 127222 27968
rect 127302 26992 127336 27968
rect 127398 26992 127432 27968
rect 127512 26992 127546 27968
rect 127608 26992 127642 27968
rect 127722 26992 127756 27968
rect 127818 26992 127852 27968
rect 127932 26992 127966 27968
rect 128028 26992 128062 27968
rect 128142 26992 128176 27968
rect 128238 26992 128272 27968
rect 128352 26992 128386 27968
rect 128448 26992 128482 27968
rect 128562 26992 128596 27968
rect 128658 26992 128692 27968
rect 128772 26992 128806 27968
rect 128868 26992 128902 27968
rect 128982 26992 129016 27968
rect 129078 26992 129112 27968
rect 129192 26992 129226 27968
rect 129288 26992 129322 27968
rect 129402 26992 129436 27968
rect 129498 26992 129532 27968
rect 129612 26992 129646 27968
rect 129708 26992 129742 27968
rect 129822 26992 129856 27968
rect 129918 26992 129952 27968
rect 130032 26992 130066 27968
rect 130128 26992 130162 27968
rect 130242 26992 130276 27968
rect 130338 26992 130372 27968
rect 130452 26992 130486 27968
rect 130548 26992 130582 27968
rect 130662 26992 130696 27968
rect 130758 26992 130792 27968
rect 130872 26992 130906 27968
rect 130968 26992 131002 27968
rect 131082 26992 131116 27968
rect 131178 26992 131212 27968
rect 131292 26992 131326 27968
rect 131388 26992 131422 27968
rect 131502 26992 131536 27968
rect 131598 26992 131632 27968
rect 131712 26992 131746 27968
rect 131808 26992 131842 27968
rect 131922 26992 131956 27968
rect 132018 26992 132052 27968
rect 132132 26992 132166 27968
rect 132228 26992 132262 27968
rect 132342 26992 132376 27968
rect 132438 26992 132472 27968
rect 132552 26992 132586 27968
rect 132648 26992 132682 27968
rect 132762 26992 132796 27968
rect 132858 26992 132892 27968
rect 132972 26992 133006 27968
rect 133068 26992 133102 27968
rect 133182 26992 133216 27968
rect 133278 26992 133312 27968
rect 133392 26992 133426 27968
rect 133488 26992 133522 27968
rect 133602 26992 133636 27968
rect 133698 26992 133732 27968
rect 133812 26992 133846 27968
rect 133908 26992 133942 27968
rect 134022 26992 134056 27968
rect 134118 26992 134152 27968
rect 134232 26992 134266 27968
rect 134328 26992 134362 27968
rect 134442 26992 134476 27968
rect 134538 26992 134572 27968
rect 134652 26992 134686 27968
rect 134748 26992 134782 27968
rect 134862 26992 134896 27968
rect 134958 26992 134992 27968
rect 135072 26992 135106 27968
rect 135168 26992 135202 27968
rect 127140 26800 127174 26942
rect 127560 26800 127594 26942
rect 127980 26800 128014 26942
rect 128400 26800 128434 26942
rect 128820 26800 128854 26942
rect 129240 26800 129274 26942
rect 129660 26800 129694 26942
rect 130080 26800 130114 26942
rect 130500 26800 130534 26942
rect 130920 26800 130954 26942
rect 131340 26800 131374 26942
rect 131760 26800 131794 26942
rect 132180 26800 132214 26942
rect 132600 26800 132634 26942
rect 133020 26800 133054 26942
rect 133440 26800 133474 26942
rect 133860 26800 133894 26942
rect 134280 26800 134314 26942
rect 134700 26800 134734 26942
rect 135120 26800 135154 26942
rect 126882 25774 126916 26750
rect 126978 25774 127012 26750
rect 127092 25774 127126 26750
rect 127188 25774 127222 26750
rect 127302 25774 127336 26750
rect 127398 25774 127432 26750
rect 127512 25774 127546 26750
rect 127608 25774 127642 26750
rect 127722 25774 127756 26750
rect 127818 25774 127852 26750
rect 127932 25774 127966 26750
rect 128028 25774 128062 26750
rect 128142 25774 128176 26750
rect 128238 25774 128272 26750
rect 128352 25774 128386 26750
rect 128448 25774 128482 26750
rect 128562 25774 128596 26750
rect 128658 25774 128692 26750
rect 128772 25774 128806 26750
rect 128868 25774 128902 26750
rect 128982 25774 129016 26750
rect 129078 25774 129112 26750
rect 129192 25774 129226 26750
rect 129288 25774 129322 26750
rect 129402 25774 129436 26750
rect 129498 25774 129532 26750
rect 129612 25774 129646 26750
rect 129708 25774 129742 26750
rect 129822 25774 129856 26750
rect 129918 25774 129952 26750
rect 130032 25774 130066 26750
rect 130128 25774 130162 26750
rect 130242 25774 130276 26750
rect 130338 25774 130372 26750
rect 130452 25774 130486 26750
rect 130548 25774 130582 26750
rect 130662 25774 130696 26750
rect 130758 25774 130792 26750
rect 130872 25774 130906 26750
rect 130968 25774 131002 26750
rect 131082 25774 131116 26750
rect 131178 25774 131212 26750
rect 131292 25774 131326 26750
rect 131388 25774 131422 26750
rect 131502 25774 131536 26750
rect 131598 25774 131632 26750
rect 131712 25774 131746 26750
rect 131808 25774 131842 26750
rect 131922 25774 131956 26750
rect 132018 25774 132052 26750
rect 132132 25774 132166 26750
rect 132228 25774 132262 26750
rect 132342 25774 132376 26750
rect 132438 25774 132472 26750
rect 132552 25774 132586 26750
rect 132648 25774 132682 26750
rect 132762 25774 132796 26750
rect 132858 25774 132892 26750
rect 132972 25774 133006 26750
rect 133068 25774 133102 26750
rect 133182 25774 133216 26750
rect 133278 25774 133312 26750
rect 133392 25774 133426 26750
rect 133488 25774 133522 26750
rect 133602 25774 133636 26750
rect 133698 25774 133732 26750
rect 133812 25774 133846 26750
rect 133908 25774 133942 26750
rect 134022 25774 134056 26750
rect 134118 25774 134152 26750
rect 134232 25774 134266 26750
rect 134328 25774 134362 26750
rect 134442 25774 134476 26750
rect 134538 25774 134572 26750
rect 134652 25774 134686 26750
rect 134748 25774 134782 26750
rect 134862 25774 134896 26750
rect 134958 25774 134992 26750
rect 135072 25774 135106 26750
rect 135168 25774 135202 26750
rect 126930 25690 127014 25724
rect 127350 25690 127434 25724
rect 127770 25690 127854 25724
rect 128190 25690 128274 25724
rect 128610 25690 128694 25724
rect 129030 25690 129114 25724
rect 129450 25690 129534 25724
rect 129870 25690 129954 25724
rect 130290 25690 130374 25724
rect 130710 25690 130794 25724
rect 131130 25690 131214 25724
rect 131550 25690 131634 25724
rect 131970 25690 132054 25724
rect 132390 25690 132474 25724
rect 132810 25690 132894 25724
rect 133230 25690 133314 25724
rect 133650 25690 133734 25724
rect 134070 25690 134154 25724
rect 134490 25690 134574 25724
rect 134910 25690 134994 25724
rect 126930 22832 126964 22833
rect 126930 22798 127014 22832
rect 127350 22832 127384 22833
rect 127350 22798 127434 22832
rect 127770 22832 127804 22833
rect 127770 22798 127854 22832
rect 128190 22832 128224 22833
rect 128190 22798 128274 22832
rect 128610 22832 128644 22833
rect 128610 22798 128694 22832
rect 129030 22832 129064 22833
rect 129030 22798 129114 22832
rect 129450 22832 129484 22833
rect 129450 22798 129534 22832
rect 129870 22832 129904 22833
rect 129870 22798 129954 22832
rect 130290 22832 130324 22833
rect 130290 22798 130374 22832
rect 130710 22832 130744 22833
rect 130710 22798 130794 22832
rect 131130 22832 131164 22833
rect 131130 22798 131214 22832
rect 131550 22832 131584 22833
rect 131550 22798 131634 22832
rect 131970 22832 132004 22833
rect 131970 22798 132054 22832
rect 132390 22832 132424 22833
rect 132390 22798 132474 22832
rect 132810 22832 132844 22833
rect 132810 22798 132894 22832
rect 133230 22832 133264 22833
rect 133230 22798 133314 22832
rect 133650 22832 133684 22833
rect 133650 22798 133734 22832
rect 134070 22832 134104 22833
rect 134070 22798 134154 22832
rect 134490 22832 134524 22833
rect 134490 22798 134574 22832
rect 134910 22832 134944 22833
rect 134910 22798 134994 22832
rect 122028 22062 122128 22162
rect 122448 22062 122548 22162
rect 122868 22062 122968 22162
rect 123288 22062 123388 22162
rect 123708 22062 123808 22162
rect 124128 22062 124228 22162
rect 124548 22062 124648 22162
rect 124968 22062 125068 22162
rect 125388 22062 125488 22162
rect 125714 22062 125814 22162
rect 122290 21942 122374 21976
rect 122710 21942 122794 21976
rect 122710 21934 122744 21942
rect 123130 21942 123214 21976
rect 123130 21934 123164 21942
rect 123550 21942 123634 21976
rect 123550 21934 123584 21942
rect 123970 21942 124054 21976
rect 123970 21934 124004 21942
rect 124390 21942 124474 21976
rect 124390 21934 124424 21942
rect 124810 21942 124894 21976
rect 124810 21934 124844 21942
rect 125230 21942 125314 21976
rect 125230 21934 125264 21942
rect 125650 21942 125734 21976
rect 125650 21934 125684 21942
rect 122032 20908 122066 21884
rect 122128 20908 122162 21884
rect 122242 20908 122276 21884
rect 122338 20908 122372 21884
rect 122452 20908 122486 21884
rect 122548 20908 122582 21884
rect 122662 20908 122696 21884
rect 122758 20908 122792 21884
rect 122872 20908 122906 21884
rect 122968 20908 123002 21884
rect 123082 20908 123116 21884
rect 123178 20908 123212 21884
rect 123292 20908 123326 21884
rect 123388 20908 123422 21884
rect 123502 20908 123536 21884
rect 123598 20908 123632 21884
rect 123712 20908 123746 21884
rect 123808 20908 123842 21884
rect 123922 20908 123956 21884
rect 124018 20908 124052 21884
rect 124132 20908 124166 21884
rect 124228 20908 124262 21884
rect 124342 20908 124376 21884
rect 124438 20908 124472 21884
rect 124552 20908 124586 21884
rect 124648 20908 124682 21884
rect 124762 20908 124796 21884
rect 124858 20908 124892 21884
rect 124972 20908 125006 21884
rect 125068 20908 125102 21884
rect 125182 20908 125216 21884
rect 125278 20908 125312 21884
rect 125392 20908 125426 21884
rect 125488 20908 125522 21884
rect 125602 20908 125636 21884
rect 125698 20908 125732 21884
rect 122080 20852 122114 20853
rect 122080 20818 122164 20852
rect 122500 20852 122534 20853
rect 122500 20818 122584 20852
rect 122920 20852 122954 20858
rect 122920 20818 123004 20852
rect 123340 20852 123374 20858
rect 123340 20818 123424 20852
rect 123760 20852 123794 20858
rect 123760 20818 123844 20852
rect 124180 20852 124214 20858
rect 124180 20818 124264 20852
rect 124600 20852 124634 20858
rect 124600 20818 124684 20852
rect 125020 20852 125054 20858
rect 125020 20818 125104 20852
rect 125440 20852 125474 20858
rect 125440 20818 125524 20852
rect 119488 20448 119786 20730
rect 119124 19284 119158 20260
rect 119212 19284 119246 20260
rect 120326 20352 120360 20353
rect 120326 20318 120410 20352
rect 120746 20352 120780 20353
rect 120746 20318 120830 20352
rect 120068 19284 120102 20260
rect 120164 19284 120198 20260
rect 120278 19284 120312 20260
rect 120374 19284 120408 20260
rect 120488 19284 120522 20260
rect 120584 19284 120618 20260
rect 120698 19284 120732 20260
rect 120794 19284 120828 20260
rect 119168 19091 119202 19234
rect 120116 19091 120150 19234
rect 120536 19091 120570 19234
rect 120956 19124 120990 19125
rect 120956 19090 121040 19124
rect 121376 19124 121410 19125
rect 121376 19090 121460 19124
rect 119120 18056 119154 19032
rect 119216 18056 119250 19032
rect 119312 18056 119346 19032
rect 119264 17964 119348 17998
rect 119858 18056 119892 19032
rect 119954 18056 119988 19032
rect 120068 18056 120102 19032
rect 120164 18056 120198 19032
rect 120278 18056 120312 19032
rect 120374 18056 120408 19032
rect 120488 18056 120522 19032
rect 120584 18056 120618 19032
rect 120698 18056 120732 19032
rect 120794 18056 120828 19032
rect 120908 18056 120942 19032
rect 121004 18056 121038 19032
rect 121118 18056 121152 19032
rect 121214 18056 121248 19032
rect 121328 18056 121362 19032
rect 121424 18056 121458 19032
rect 119906 17996 119940 17997
rect 119906 17962 119990 17996
rect 120326 17996 120360 17997
rect 120326 17962 120410 17996
rect 120746 17996 120780 17997
rect 120746 17962 120830 17996
rect 121166 17996 121200 17997
rect 121166 17962 121250 17996
rect 122080 20360 122114 20361
rect 122080 20326 122164 20360
rect 122500 20360 122534 20361
rect 122500 20326 122584 20360
rect 122920 20360 122954 20361
rect 122920 20326 123004 20360
rect 123340 20360 123374 20361
rect 123340 20326 123424 20360
rect 123760 20360 123794 20361
rect 123760 20326 123844 20360
rect 124180 20360 124214 20361
rect 124180 20326 124264 20360
rect 124600 20360 124634 20361
rect 124600 20326 124684 20360
rect 125020 20360 125054 20361
rect 125020 20326 125104 20360
rect 125440 20360 125474 20361
rect 125440 20326 125524 20360
rect 122032 19292 122066 20268
rect 122128 19292 122162 20268
rect 122242 19292 122276 20268
rect 122338 19292 122372 20268
rect 122452 19292 122486 20268
rect 122548 19292 122582 20268
rect 122662 19292 122696 20268
rect 122758 19292 122792 20268
rect 122872 19292 122906 20268
rect 122968 19292 123002 20268
rect 123082 19292 123116 20268
rect 123178 19292 123212 20268
rect 123292 19292 123326 20268
rect 123388 19292 123422 20268
rect 123502 19292 123536 20268
rect 123598 19292 123632 20268
rect 123712 19292 123746 20268
rect 123808 19292 123842 20268
rect 123922 19292 123956 20268
rect 124018 19292 124052 20268
rect 124132 19292 124166 20268
rect 124228 19292 124262 20268
rect 124342 19292 124376 20268
rect 124438 19292 124472 20268
rect 124552 19292 124586 20268
rect 124648 19292 124682 20268
rect 124762 19292 124796 20268
rect 124858 19292 124892 20268
rect 124972 19292 125006 20268
rect 125068 19292 125102 20268
rect 125182 19292 125216 20268
rect 125278 19292 125312 20268
rect 125392 19292 125426 20268
rect 125488 19292 125522 20268
rect 125602 19292 125636 20268
rect 125698 19292 125732 20268
rect 122290 19091 122324 19233
rect 122710 19091 122744 19233
rect 123130 19091 123164 19233
rect 123550 19091 123584 19233
rect 123970 19091 124004 19233
rect 124390 19091 124424 19233
rect 124810 19091 124844 19233
rect 125230 19091 125264 19233
rect 125650 19091 125684 19233
rect 122032 18056 122066 19032
rect 122128 18056 122162 19032
rect 122242 18056 122276 19032
rect 122338 18056 122372 19032
rect 122452 18056 122486 19032
rect 122548 18056 122582 19032
rect 122662 18056 122696 19032
rect 122758 18056 122792 19032
rect 122872 18056 122906 19032
rect 122968 18056 123002 19032
rect 123082 18056 123116 19032
rect 123178 18056 123212 19032
rect 123292 18056 123326 19032
rect 123388 18056 123422 19032
rect 123502 18056 123536 19032
rect 123598 18056 123632 19032
rect 123712 18056 123746 19032
rect 123808 18056 123842 19032
rect 123922 18056 123956 19032
rect 124018 18056 124052 19032
rect 124132 18056 124166 19032
rect 124228 18056 124262 19032
rect 124342 18056 124376 19032
rect 124438 18056 124472 19032
rect 124552 18056 124586 19032
rect 124648 18056 124682 19032
rect 124762 18056 124796 19032
rect 124858 18056 124892 19032
rect 124972 18056 125006 19032
rect 125068 18056 125102 19032
rect 125182 18056 125216 19032
rect 125278 18056 125312 19032
rect 125392 18056 125426 19032
rect 125488 18056 125522 19032
rect 125602 18056 125636 19032
rect 125698 18056 125732 19032
rect 122080 17996 122114 17997
rect 122080 17962 122164 17996
rect 122500 17996 122534 17997
rect 122500 17962 122584 17996
rect 122920 17996 122954 17997
rect 122920 17962 123004 17996
rect 123340 17996 123374 17997
rect 123340 17962 123424 17996
rect 123760 17996 123794 17997
rect 123760 17962 123844 17996
rect 124180 17996 124214 17997
rect 124180 17962 124264 17996
rect 124600 17996 124634 17997
rect 124600 17962 124684 17996
rect 125020 17996 125054 17997
rect 125020 17962 125104 17996
rect 125440 17996 125474 17997
rect 125440 17962 125524 17996
rect 121904 17802 122004 17902
rect 122324 17870 122424 17902
rect 122744 17870 122844 17902
rect 123164 17870 123264 17902
rect 123584 17870 123684 17902
rect 124004 17870 124104 17902
rect 124424 17870 124524 17902
rect 124844 17870 124944 17902
rect 125264 17870 125364 17902
rect 125684 17870 125784 17902
rect 122324 17836 122424 17870
rect 122744 17836 122844 17870
rect 123164 17836 123264 17870
rect 123584 17836 123684 17870
rect 124004 17836 124104 17870
rect 124424 17836 124524 17870
rect 124844 17836 124944 17870
rect 125264 17836 125364 17870
rect 125684 17836 125784 17870
rect 126882 21764 126916 22740
rect 126978 21764 127012 22740
rect 127092 21764 127126 22740
rect 127188 21764 127222 22740
rect 127302 21764 127336 22740
rect 127398 21764 127432 22740
rect 127512 21764 127546 22740
rect 127608 21764 127642 22740
rect 127722 21764 127756 22740
rect 127818 21764 127852 22740
rect 127932 21764 127966 22740
rect 128028 21764 128062 22740
rect 128142 21764 128176 22740
rect 128238 21764 128272 22740
rect 128352 21764 128386 22740
rect 128448 21764 128482 22740
rect 128562 21764 128596 22740
rect 128658 21764 128692 22740
rect 128772 21764 128806 22740
rect 128868 21764 128902 22740
rect 128982 21764 129016 22740
rect 129078 21764 129112 22740
rect 129192 21764 129226 22740
rect 129288 21764 129322 22740
rect 129402 21764 129436 22740
rect 129498 21764 129532 22740
rect 129612 21764 129646 22740
rect 129708 21764 129742 22740
rect 129822 21764 129856 22740
rect 129918 21764 129952 22740
rect 130032 21764 130066 22740
rect 130128 21764 130162 22740
rect 130242 21764 130276 22740
rect 130338 21764 130372 22740
rect 130452 21764 130486 22740
rect 130548 21764 130582 22740
rect 130662 21764 130696 22740
rect 130758 21764 130792 22740
rect 130872 21764 130906 22740
rect 130968 21764 131002 22740
rect 131082 21764 131116 22740
rect 131178 21764 131212 22740
rect 131292 21764 131326 22740
rect 131388 21764 131422 22740
rect 131502 21764 131536 22740
rect 131598 21764 131632 22740
rect 131712 21764 131746 22740
rect 131808 21764 131842 22740
rect 131922 21764 131956 22740
rect 132018 21764 132052 22740
rect 132132 21764 132166 22740
rect 132228 21764 132262 22740
rect 132342 21764 132376 22740
rect 132438 21764 132472 22740
rect 132552 21764 132586 22740
rect 132648 21764 132682 22740
rect 132762 21764 132796 22740
rect 132858 21764 132892 22740
rect 132972 21764 133006 22740
rect 133068 21764 133102 22740
rect 133182 21764 133216 22740
rect 133278 21764 133312 22740
rect 133392 21764 133426 22740
rect 133488 21764 133522 22740
rect 133602 21764 133636 22740
rect 133698 21764 133732 22740
rect 133812 21764 133846 22740
rect 133908 21764 133942 22740
rect 134022 21764 134056 22740
rect 134118 21764 134152 22740
rect 134232 21764 134266 22740
rect 134328 21764 134362 22740
rect 134442 21764 134476 22740
rect 134538 21764 134572 22740
rect 134652 21764 134686 22740
rect 134748 21764 134782 22740
rect 134862 21764 134896 22740
rect 134958 21764 134992 22740
rect 135072 21764 135106 22740
rect 135168 21764 135202 22740
rect 127140 21563 127174 21705
rect 127560 21563 127594 21705
rect 127980 21563 128014 21705
rect 128400 21563 128434 21705
rect 128820 21563 128854 21705
rect 129240 21563 129274 21705
rect 129660 21563 129694 21705
rect 130080 21563 130114 21705
rect 130500 21563 130534 21705
rect 130920 21563 130954 21705
rect 131340 21563 131374 21705
rect 131760 21563 131794 21705
rect 132180 21563 132214 21705
rect 132600 21563 132634 21705
rect 133020 21563 133054 21705
rect 133440 21563 133474 21705
rect 133860 21563 133894 21705
rect 134280 21563 134314 21705
rect 134700 21563 134734 21705
rect 135120 21563 135154 21705
rect 126882 20528 126916 21504
rect 126978 20528 127012 21504
rect 127092 20528 127126 21504
rect 127188 20528 127222 21504
rect 127302 20528 127336 21504
rect 127398 20528 127432 21504
rect 127512 20528 127546 21504
rect 127608 20528 127642 21504
rect 127722 20528 127756 21504
rect 127818 20528 127852 21504
rect 127932 20528 127966 21504
rect 128028 20528 128062 21504
rect 128142 20528 128176 21504
rect 128238 20528 128272 21504
rect 128352 20528 128386 21504
rect 128448 20528 128482 21504
rect 128562 20528 128596 21504
rect 128658 20528 128692 21504
rect 128772 20528 128806 21504
rect 128868 20528 128902 21504
rect 128982 20528 129016 21504
rect 129078 20528 129112 21504
rect 129192 20528 129226 21504
rect 129288 20528 129322 21504
rect 129402 20528 129436 21504
rect 129498 20528 129532 21504
rect 129612 20528 129646 21504
rect 129708 20528 129742 21504
rect 129822 20528 129856 21504
rect 129918 20528 129952 21504
rect 130032 20528 130066 21504
rect 130128 20528 130162 21504
rect 130242 20528 130276 21504
rect 130338 20528 130372 21504
rect 130452 20528 130486 21504
rect 130548 20528 130582 21504
rect 130662 20528 130696 21504
rect 130758 20528 130792 21504
rect 130872 20528 130906 21504
rect 130968 20528 131002 21504
rect 131082 20528 131116 21504
rect 131178 20528 131212 21504
rect 131292 20528 131326 21504
rect 131388 20528 131422 21504
rect 131502 20528 131536 21504
rect 131598 20528 131632 21504
rect 131712 20528 131746 21504
rect 131808 20528 131842 21504
rect 131922 20528 131956 21504
rect 132018 20528 132052 21504
rect 132132 20528 132166 21504
rect 132228 20528 132262 21504
rect 132342 20528 132376 21504
rect 132438 20528 132472 21504
rect 132552 20528 132586 21504
rect 132648 20528 132682 21504
rect 132762 20528 132796 21504
rect 132858 20528 132892 21504
rect 132972 20528 133006 21504
rect 133068 20528 133102 21504
rect 133182 20528 133216 21504
rect 133278 20528 133312 21504
rect 133392 20528 133426 21504
rect 133488 20528 133522 21504
rect 133602 20528 133636 21504
rect 133698 20528 133732 21504
rect 133812 20528 133846 21504
rect 133908 20528 133942 21504
rect 134022 20528 134056 21504
rect 134118 20528 134152 21504
rect 134232 20528 134266 21504
rect 134328 20528 134362 21504
rect 134442 20528 134476 21504
rect 134538 20528 134572 21504
rect 134652 20528 134686 21504
rect 134748 20528 134782 21504
rect 134862 20528 134896 21504
rect 134958 20528 134992 21504
rect 135072 20528 135106 21504
rect 135168 20528 135202 21504
rect 126930 20327 126964 20469
rect 127350 20327 127384 20469
rect 127770 20327 127804 20469
rect 128190 20327 128224 20469
rect 128610 20327 128644 20469
rect 129030 20327 129064 20469
rect 129450 20327 129484 20469
rect 129870 20327 129904 20469
rect 130290 20327 130324 20469
rect 130710 20327 130744 20469
rect 131130 20327 131164 20469
rect 131550 20327 131584 20469
rect 131970 20327 132004 20469
rect 132390 20327 132424 20469
rect 132810 20327 132844 20469
rect 133230 20327 133264 20469
rect 133650 20327 133684 20469
rect 134070 20327 134104 20469
rect 134490 20327 134524 20469
rect 134910 20327 134944 20469
rect 126882 19292 126916 20268
rect 126978 19292 127012 20268
rect 127092 19292 127126 20268
rect 127188 19292 127222 20268
rect 127302 19292 127336 20268
rect 127398 19292 127432 20268
rect 127512 19292 127546 20268
rect 127608 19292 127642 20268
rect 127722 19292 127756 20268
rect 127818 19292 127852 20268
rect 127932 19292 127966 20268
rect 128028 19292 128062 20268
rect 128142 19292 128176 20268
rect 128238 19292 128272 20268
rect 128352 19292 128386 20268
rect 128448 19292 128482 20268
rect 128562 19292 128596 20268
rect 128658 19292 128692 20268
rect 128772 19292 128806 20268
rect 128868 19292 128902 20268
rect 128982 19292 129016 20268
rect 129078 19292 129112 20268
rect 129192 19292 129226 20268
rect 129288 19292 129322 20268
rect 129402 19292 129436 20268
rect 129498 19292 129532 20268
rect 129612 19292 129646 20268
rect 129708 19292 129742 20268
rect 129822 19292 129856 20268
rect 129918 19292 129952 20268
rect 130032 19292 130066 20268
rect 130128 19292 130162 20268
rect 130242 19292 130276 20268
rect 130338 19292 130372 20268
rect 130452 19292 130486 20268
rect 130548 19292 130582 20268
rect 130662 19292 130696 20268
rect 130758 19292 130792 20268
rect 130872 19292 130906 20268
rect 130968 19292 131002 20268
rect 131082 19292 131116 20268
rect 131178 19292 131212 20268
rect 131292 19292 131326 20268
rect 131388 19292 131422 20268
rect 131502 19292 131536 20268
rect 131598 19292 131632 20268
rect 131712 19292 131746 20268
rect 131808 19292 131842 20268
rect 131922 19292 131956 20268
rect 132018 19292 132052 20268
rect 132132 19292 132166 20268
rect 132228 19292 132262 20268
rect 132342 19292 132376 20268
rect 132438 19292 132472 20268
rect 132552 19292 132586 20268
rect 132648 19292 132682 20268
rect 132762 19292 132796 20268
rect 132858 19292 132892 20268
rect 132972 19292 133006 20268
rect 133068 19292 133102 20268
rect 133182 19292 133216 20268
rect 133278 19292 133312 20268
rect 133392 19292 133426 20268
rect 133488 19292 133522 20268
rect 133602 19292 133636 20268
rect 133698 19292 133732 20268
rect 133812 19292 133846 20268
rect 133908 19292 133942 20268
rect 134022 19292 134056 20268
rect 134118 19292 134152 20268
rect 134232 19292 134266 20268
rect 134328 19292 134362 20268
rect 134442 19292 134476 20268
rect 134538 19292 134572 20268
rect 134652 19292 134686 20268
rect 134748 19292 134782 20268
rect 134862 19292 134896 20268
rect 134958 19292 134992 20268
rect 135072 19292 135106 20268
rect 135168 19292 135202 20268
rect 127140 19091 127174 19233
rect 127560 19091 127594 19233
rect 127980 19091 128014 19233
rect 128400 19091 128434 19233
rect 128820 19091 128854 19233
rect 129240 19091 129274 19233
rect 129660 19091 129694 19233
rect 130080 19091 130114 19233
rect 130500 19091 130534 19233
rect 130920 19091 130954 19233
rect 131340 19091 131374 19233
rect 131760 19091 131794 19233
rect 132180 19091 132214 19233
rect 132600 19091 132634 19233
rect 133020 19091 133054 19233
rect 133440 19091 133474 19233
rect 133860 19091 133894 19233
rect 134280 19091 134314 19233
rect 134700 19091 134734 19233
rect 135120 19091 135154 19233
rect 126882 18056 126916 19032
rect 126978 18056 127012 19032
rect 127092 18056 127126 19032
rect 127188 18056 127222 19032
rect 127302 18056 127336 19032
rect 127398 18056 127432 19032
rect 127512 18056 127546 19032
rect 127608 18056 127642 19032
rect 127722 18056 127756 19032
rect 127818 18056 127852 19032
rect 127932 18056 127966 19032
rect 128028 18056 128062 19032
rect 128142 18056 128176 19032
rect 128238 18056 128272 19032
rect 128352 18056 128386 19032
rect 128448 18056 128482 19032
rect 128562 18056 128596 19032
rect 128658 18056 128692 19032
rect 128772 18056 128806 19032
rect 128868 18056 128902 19032
rect 128982 18056 129016 19032
rect 129078 18056 129112 19032
rect 129192 18056 129226 19032
rect 129288 18056 129322 19032
rect 129402 18056 129436 19032
rect 129498 18056 129532 19032
rect 129612 18056 129646 19032
rect 129708 18056 129742 19032
rect 129822 18056 129856 19032
rect 129918 18056 129952 19032
rect 130032 18056 130066 19032
rect 130128 18056 130162 19032
rect 130242 18056 130276 19032
rect 130338 18056 130372 19032
rect 130452 18056 130486 19032
rect 130548 18056 130582 19032
rect 130662 18056 130696 19032
rect 130758 18056 130792 19032
rect 130872 18056 130906 19032
rect 130968 18056 131002 19032
rect 131082 18056 131116 19032
rect 131178 18056 131212 19032
rect 131292 18056 131326 19032
rect 131388 18056 131422 19032
rect 131502 18056 131536 19032
rect 131598 18056 131632 19032
rect 131712 18056 131746 19032
rect 131808 18056 131842 19032
rect 131922 18056 131956 19032
rect 132018 18056 132052 19032
rect 132132 18056 132166 19032
rect 132228 18056 132262 19032
rect 132342 18056 132376 19032
rect 132438 18056 132472 19032
rect 132552 18056 132586 19032
rect 132648 18056 132682 19032
rect 132762 18056 132796 19032
rect 132858 18056 132892 19032
rect 132972 18056 133006 19032
rect 133068 18056 133102 19032
rect 133182 18056 133216 19032
rect 133278 18056 133312 19032
rect 133392 18056 133426 19032
rect 133488 18056 133522 19032
rect 133602 18056 133636 19032
rect 133698 18056 133732 19032
rect 133812 18056 133846 19032
rect 133908 18056 133942 19032
rect 134022 18056 134056 19032
rect 134118 18056 134152 19032
rect 134232 18056 134266 19032
rect 134328 18056 134362 19032
rect 134442 18056 134476 19032
rect 134538 18056 134572 19032
rect 134652 18056 134686 19032
rect 134748 18056 134782 19032
rect 134862 18056 134896 19032
rect 134958 18056 134992 19032
rect 135072 18056 135106 19032
rect 135168 18056 135202 19032
rect 126930 17996 126964 17997
rect 126930 17962 127014 17996
rect 127350 17996 127384 17997
rect 127350 17962 127434 17996
rect 127770 17996 127804 17997
rect 127770 17962 127854 17996
rect 128190 17996 128224 17997
rect 128190 17962 128274 17996
rect 128610 17996 128644 17997
rect 128610 17962 128694 17996
rect 129030 17996 129064 17997
rect 129030 17962 129114 17996
rect 129450 17996 129484 17997
rect 129450 17962 129534 17996
rect 129870 17996 129904 17997
rect 129870 17962 129954 17996
rect 130290 17996 130324 17997
rect 130290 17962 130374 17996
rect 130710 17996 130744 17997
rect 130710 17962 130794 17996
rect 131130 17996 131164 17997
rect 131130 17962 131214 17996
rect 131550 17996 131584 17997
rect 131550 17962 131634 17996
rect 131970 17996 132004 17997
rect 131970 17962 132054 17996
rect 132390 17996 132424 17997
rect 132390 17962 132474 17996
rect 132810 17996 132844 17997
rect 132810 17962 132894 17996
rect 133230 17996 133264 17997
rect 133230 17962 133314 17996
rect 133650 17996 133684 17997
rect 133650 17962 133734 17996
rect 134070 17996 134104 17997
rect 134070 17962 134154 17996
rect 134490 17996 134524 17997
rect 134490 17962 134574 17996
rect 134910 17996 134944 17997
rect 134910 17962 134994 17996
rect 122324 17802 122424 17836
rect 122744 17802 122844 17836
rect 123164 17802 123264 17836
rect 123584 17802 123684 17836
rect 124004 17802 124104 17836
rect 124424 17802 124524 17836
rect 124844 17802 124944 17836
rect 125264 17802 125364 17836
rect 125684 17802 125784 17836
rect 126746 17786 126846 17886
rect 127166 17854 127266 17886
rect 127586 17854 127686 17886
rect 128006 17854 128106 17886
rect 128426 17854 128526 17886
rect 128846 17854 128946 17886
rect 129266 17854 129366 17886
rect 129686 17854 129786 17886
rect 130106 17854 130206 17886
rect 130526 17854 130626 17886
rect 130946 17854 131046 17886
rect 131366 17854 131466 17886
rect 131786 17854 131886 17886
rect 132206 17854 132306 17886
rect 132626 17854 132726 17886
rect 133046 17854 133146 17886
rect 133466 17854 133566 17886
rect 133886 17854 133986 17886
rect 134306 17854 134406 17886
rect 134726 17854 134826 17886
rect 135146 17854 135246 17886
rect 127166 17820 127266 17854
rect 127586 17820 127686 17854
rect 128006 17820 128106 17854
rect 128426 17820 128526 17854
rect 128846 17820 128946 17854
rect 129266 17820 129366 17854
rect 129686 17820 129786 17854
rect 130106 17820 130206 17854
rect 130526 17820 130626 17854
rect 130946 17820 131046 17854
rect 131366 17820 131466 17854
rect 131786 17820 131886 17854
rect 132206 17820 132306 17854
rect 132626 17820 132726 17854
rect 133046 17820 133146 17854
rect 133466 17820 133566 17854
rect 133886 17820 133986 17854
rect 134306 17820 134406 17854
rect 134726 17820 134826 17854
rect 135146 17820 135182 17854
rect 135182 17820 135246 17854
rect 127166 17786 127266 17820
rect 127586 17786 127686 17820
rect 128006 17786 128106 17820
rect 128426 17786 128526 17820
rect 128846 17786 128946 17820
rect 129266 17786 129366 17820
rect 129686 17786 129786 17820
rect 130106 17786 130206 17820
rect 130526 17786 130626 17820
rect 130946 17786 131046 17820
rect 131366 17786 131466 17820
rect 131786 17786 131886 17820
rect 132206 17786 132306 17820
rect 132626 17786 132726 17820
rect 133046 17786 133146 17820
rect 133466 17786 133566 17820
rect 133886 17786 133986 17820
rect 134306 17786 134406 17820
rect 134726 17786 134826 17820
rect 135146 17786 135246 17820
rect 119522 17622 119666 17770
rect 116190 16616 116284 16830
rect 116382 16530 116416 16906
rect 116476 16530 116510 16906
rect 116564 16530 116598 16906
rect 116512 16464 116586 16470
rect 116512 16432 116518 16464
rect 116518 16432 116576 16464
rect 116576 16432 116586 16464
rect 116512 16424 116586 16432
rect 116350 16378 116424 16384
rect 116350 16346 116360 16378
rect 116360 16346 116418 16378
rect 116418 16346 116424 16378
rect 116350 16338 116424 16346
rect 116208 15998 116284 16204
rect 116382 15910 116416 16286
rect 116476 15910 116510 16286
rect 116564 15910 116598 16286
rect 115750 15322 115790 15438
rect 115856 15102 115890 15478
rect 115944 15102 115978 15478
rect 116208 15186 116284 15392
rect 116382 15104 116416 15480
rect 116476 15104 116510 15480
rect 116564 15104 116598 15480
rect 115900 15043 115934 15044
rect 115900 15009 115934 15043
rect 116350 15044 116424 15052
rect 116350 15012 116360 15044
rect 116360 15012 116418 15044
rect 116418 15012 116424 15044
rect 115900 14906 115934 15009
rect 116350 15006 116424 15012
rect 116512 14958 116586 14966
rect 116512 14926 116518 14958
rect 116518 14926 116576 14958
rect 116576 14926 116586 14958
rect 116512 14920 116586 14926
rect 115900 14872 115934 14906
rect 115726 14668 115790 14810
rect 115856 14646 115890 14822
rect 115944 14646 115978 14822
rect 116190 14560 116284 14774
rect 116382 14484 116416 14860
rect 116476 14484 116510 14860
rect 116564 14484 116598 14860
rect 119522 13620 119666 13768
rect 119264 13392 119348 13426
rect 119120 12358 119154 13334
rect 119216 12358 119250 13334
rect 119312 12358 119346 13334
rect 121904 13488 122004 13588
rect 122324 13554 122424 13588
rect 122744 13554 122844 13588
rect 123164 13554 123264 13588
rect 123584 13554 123684 13588
rect 124004 13554 124104 13588
rect 124424 13554 124524 13588
rect 124844 13554 124944 13588
rect 125264 13554 125364 13588
rect 125684 13554 125784 13588
rect 122324 13520 122424 13554
rect 122744 13520 122844 13554
rect 123164 13520 123264 13554
rect 123584 13520 123684 13554
rect 124004 13520 124104 13554
rect 124424 13520 124524 13554
rect 124844 13520 124944 13554
rect 125264 13520 125364 13554
rect 125684 13520 125784 13554
rect 122324 13488 122424 13520
rect 122744 13488 122844 13520
rect 123164 13488 123264 13520
rect 123584 13488 123684 13520
rect 124004 13488 124104 13520
rect 124424 13488 124524 13520
rect 124844 13488 124944 13520
rect 125264 13488 125364 13520
rect 125684 13488 125784 13520
rect 119906 13394 119990 13428
rect 119906 13393 119940 13394
rect 120326 13394 120410 13428
rect 120326 13393 120360 13394
rect 120746 13394 120830 13428
rect 120746 13393 120780 13394
rect 121166 13394 121250 13428
rect 121166 13393 121200 13394
rect 119858 12358 119892 13334
rect 119954 12358 119988 13334
rect 120068 12358 120102 13334
rect 120164 12358 120198 13334
rect 120278 12358 120312 13334
rect 120374 12358 120408 13334
rect 120488 12358 120522 13334
rect 120584 12358 120618 13334
rect 120698 12358 120732 13334
rect 120794 12358 120828 13334
rect 120908 12358 120942 13334
rect 121004 12358 121038 13334
rect 121118 12358 121152 13334
rect 121214 12358 121248 13334
rect 121328 12358 121362 13334
rect 121424 12358 121458 13334
rect 119168 12156 119202 12299
rect 120116 12156 120150 12299
rect 120536 12156 120570 12299
rect 120956 12266 121040 12300
rect 120956 12265 120990 12266
rect 121376 12266 121460 12300
rect 121376 12265 121410 12266
rect 119124 11130 119158 12106
rect 119212 11130 119246 12106
rect 120068 11130 120102 12106
rect 120164 11130 120198 12106
rect 120278 11130 120312 12106
rect 120374 11130 120408 12106
rect 120488 11130 120522 12106
rect 120584 11130 120618 12106
rect 120698 11130 120732 12106
rect 120794 11130 120828 12106
rect 120326 11038 120410 11072
rect 120326 11037 120360 11038
rect 120746 11038 120830 11072
rect 120746 11037 120780 11038
rect 122080 13394 122164 13428
rect 122080 13393 122114 13394
rect 122500 13394 122584 13428
rect 122500 13393 122534 13394
rect 122920 13394 123004 13428
rect 122920 13393 122954 13394
rect 123340 13394 123424 13428
rect 123340 13393 123374 13394
rect 123760 13394 123844 13428
rect 123760 13393 123794 13394
rect 124180 13394 124264 13428
rect 124180 13393 124214 13394
rect 124600 13394 124684 13428
rect 124600 13393 124634 13394
rect 125020 13394 125104 13428
rect 125020 13393 125054 13394
rect 125440 13394 125524 13428
rect 125440 13393 125474 13394
rect 122032 12358 122066 13334
rect 122128 12358 122162 13334
rect 122242 12358 122276 13334
rect 122338 12358 122372 13334
rect 122452 12358 122486 13334
rect 122548 12358 122582 13334
rect 122662 12358 122696 13334
rect 122758 12358 122792 13334
rect 122872 12358 122906 13334
rect 122968 12358 123002 13334
rect 123082 12358 123116 13334
rect 123178 12358 123212 13334
rect 123292 12358 123326 13334
rect 123388 12358 123422 13334
rect 123502 12358 123536 13334
rect 123598 12358 123632 13334
rect 123712 12358 123746 13334
rect 123808 12358 123842 13334
rect 123922 12358 123956 13334
rect 124018 12358 124052 13334
rect 124132 12358 124166 13334
rect 124228 12358 124262 13334
rect 124342 12358 124376 13334
rect 124438 12358 124472 13334
rect 124552 12358 124586 13334
rect 124648 12358 124682 13334
rect 124762 12358 124796 13334
rect 124858 12358 124892 13334
rect 124972 12358 125006 13334
rect 125068 12358 125102 13334
rect 125182 12358 125216 13334
rect 125278 12358 125312 13334
rect 125392 12358 125426 13334
rect 125488 12358 125522 13334
rect 125602 12358 125636 13334
rect 125698 12358 125732 13334
rect 122290 12157 122324 12299
rect 122710 12157 122744 12299
rect 123130 12157 123164 12299
rect 123550 12157 123584 12299
rect 123970 12157 124004 12299
rect 124390 12157 124424 12299
rect 124810 12157 124844 12299
rect 125230 12157 125264 12299
rect 125650 12157 125684 12299
rect 122032 11122 122066 12098
rect 122128 11122 122162 12098
rect 122242 11122 122276 12098
rect 122338 11122 122372 12098
rect 122452 11122 122486 12098
rect 122548 11122 122582 12098
rect 122662 11122 122696 12098
rect 122758 11122 122792 12098
rect 122872 11122 122906 12098
rect 122968 11122 123002 12098
rect 123082 11122 123116 12098
rect 123178 11122 123212 12098
rect 123292 11122 123326 12098
rect 123388 11122 123422 12098
rect 123502 11122 123536 12098
rect 123598 11122 123632 12098
rect 123712 11122 123746 12098
rect 123808 11122 123842 12098
rect 123922 11122 123956 12098
rect 124018 11122 124052 12098
rect 124132 11122 124166 12098
rect 124228 11122 124262 12098
rect 124342 11122 124376 12098
rect 124438 11122 124472 12098
rect 124552 11122 124586 12098
rect 124648 11122 124682 12098
rect 124762 11122 124796 12098
rect 124858 11122 124892 12098
rect 124972 11122 125006 12098
rect 125068 11122 125102 12098
rect 125182 11122 125216 12098
rect 125278 11122 125312 12098
rect 125392 11122 125426 12098
rect 125488 11122 125522 12098
rect 125602 11122 125636 12098
rect 125698 11122 125732 12098
rect 122080 11030 122164 11064
rect 122080 11029 122114 11030
rect 122500 11030 122584 11064
rect 122500 11029 122534 11030
rect 122920 11030 123004 11064
rect 122920 11029 122954 11030
rect 123340 11030 123424 11064
rect 123340 11029 123374 11030
rect 123760 11030 123844 11064
rect 123760 11029 123794 11030
rect 124180 11030 124264 11064
rect 124180 11029 124214 11030
rect 124600 11030 124684 11064
rect 124600 11029 124634 11030
rect 125020 11030 125104 11064
rect 125020 11029 125054 11030
rect 125440 11030 125524 11064
rect 125440 11029 125474 11030
rect 119488 10660 119786 10942
rect 122080 9138 122164 9172
rect 122080 9137 122114 9138
rect 122500 9138 122584 9172
rect 122500 9137 122534 9138
rect 122920 9138 123004 9172
rect 122920 9132 122954 9138
rect 123340 9138 123424 9172
rect 123340 9132 123374 9138
rect 123760 9138 123844 9172
rect 123760 9132 123794 9138
rect 124180 9138 124264 9172
rect 124180 9132 124214 9138
rect 124600 9138 124684 9172
rect 124600 9132 124634 9138
rect 125020 9138 125104 9172
rect 125020 9132 125054 9138
rect 125440 9138 125524 9172
rect 125440 9132 125474 9138
rect 122032 8106 122066 9082
rect 122128 8106 122162 9082
rect 122242 8106 122276 9082
rect 122338 8106 122372 9082
rect 122452 8106 122486 9082
rect 122548 8106 122582 9082
rect 122662 8106 122696 9082
rect 122758 8106 122792 9082
rect 122872 8106 122906 9082
rect 122968 8106 123002 9082
rect 123082 8106 123116 9082
rect 123178 8106 123212 9082
rect 123292 8106 123326 9082
rect 123388 8106 123422 9082
rect 123502 8106 123536 9082
rect 123598 8106 123632 9082
rect 123712 8106 123746 9082
rect 123808 8106 123842 9082
rect 123922 8106 123956 9082
rect 124018 8106 124052 9082
rect 124132 8106 124166 9082
rect 124228 8106 124262 9082
rect 124342 8106 124376 9082
rect 124438 8106 124472 9082
rect 124552 8106 124586 9082
rect 124648 8106 124682 9082
rect 124762 8106 124796 9082
rect 124858 8106 124892 9082
rect 124972 8106 125006 9082
rect 125068 8106 125102 9082
rect 125182 8106 125216 9082
rect 125278 8106 125312 9082
rect 125392 8106 125426 9082
rect 125488 8106 125522 9082
rect 125602 8106 125636 9082
rect 125698 8106 125732 9082
rect 122290 8014 122374 8048
rect 122710 8048 122744 8056
rect 122710 8014 122794 8048
rect 123130 8048 123164 8056
rect 123130 8014 123214 8048
rect 123550 8048 123584 8056
rect 123550 8014 123634 8048
rect 123970 8048 124004 8056
rect 123970 8014 124054 8048
rect 124390 8048 124424 8056
rect 124390 8014 124474 8048
rect 124810 8048 124844 8056
rect 124810 8014 124894 8048
rect 125230 8048 125264 8056
rect 125230 8014 125314 8048
rect 125650 8048 125684 8056
rect 125650 8014 125734 8048
rect 122028 7828 122128 7928
rect 122448 7828 122548 7928
rect 122868 7828 122968 7928
rect 123288 7828 123388 7928
rect 123708 7828 123808 7928
rect 124128 7828 124228 7928
rect 124548 7828 124648 7928
rect 124968 7828 125068 7928
rect 125388 7828 125488 7928
rect 125714 7828 125814 7928
<< metal1 >>
rect 126834 28304 126944 28316
rect 127254 28304 127364 28316
rect 127674 28304 127784 28316
rect 128094 28304 128204 28316
rect 128514 28304 128624 28316
rect 128934 28304 129044 28316
rect 129354 28304 129464 28316
rect 129774 28304 129884 28316
rect 130194 28304 130304 28316
rect 130614 28304 130724 28316
rect 131034 28304 131144 28316
rect 131454 28304 131564 28316
rect 131874 28304 131984 28316
rect 132294 28304 132404 28316
rect 132714 28304 132824 28316
rect 133134 28304 133244 28316
rect 133554 28304 133664 28316
rect 133974 28304 134084 28316
rect 134394 28304 134504 28316
rect 134814 28304 134924 28316
rect 135162 28304 135272 28316
rect 126830 28200 126840 28304
rect 126938 28200 126948 28304
rect 127250 28200 127260 28304
rect 127358 28200 127368 28304
rect 127670 28200 127680 28304
rect 127778 28200 127788 28304
rect 128090 28200 128100 28304
rect 128198 28200 128208 28304
rect 128510 28200 128520 28304
rect 128618 28200 128628 28304
rect 128930 28200 128940 28304
rect 129038 28200 129048 28304
rect 129350 28200 129360 28304
rect 129458 28200 129468 28304
rect 129770 28200 129780 28304
rect 129878 28200 129888 28304
rect 130190 28200 130200 28304
rect 130298 28200 130308 28304
rect 130610 28200 130620 28304
rect 130718 28200 130728 28304
rect 131030 28200 131040 28304
rect 131138 28200 131148 28304
rect 131450 28200 131460 28304
rect 131558 28200 131568 28304
rect 131870 28200 131880 28304
rect 131978 28200 131988 28304
rect 132290 28200 132300 28304
rect 132398 28200 132408 28304
rect 132710 28200 132720 28304
rect 132818 28200 132828 28304
rect 133130 28200 133140 28304
rect 133238 28200 133248 28304
rect 133550 28200 133560 28304
rect 133658 28200 133668 28304
rect 133970 28200 133980 28304
rect 134078 28200 134088 28304
rect 134390 28200 134400 28304
rect 134498 28200 134508 28304
rect 134810 28200 134820 28304
rect 134918 28200 134928 28304
rect 135158 28200 135168 28304
rect 135266 28200 135276 28304
rect 126834 28188 126944 28200
rect 127254 28188 127364 28200
rect 127674 28188 127784 28200
rect 128094 28188 128204 28200
rect 128514 28188 128624 28200
rect 128934 28188 129044 28200
rect 129354 28188 129464 28200
rect 129774 28188 129884 28200
rect 130194 28188 130304 28200
rect 130614 28188 130724 28200
rect 131034 28188 131144 28200
rect 131454 28188 131564 28200
rect 131874 28188 131984 28200
rect 132294 28188 132404 28200
rect 132714 28188 132824 28200
rect 133134 28188 133244 28200
rect 133554 28188 133664 28200
rect 133974 28188 134084 28200
rect 134394 28188 134504 28200
rect 134814 28188 134924 28200
rect 135162 28188 135272 28200
rect 125964 28052 135006 28058
rect 125964 28018 126930 28052
rect 127014 28018 127350 28052
rect 127434 28018 127770 28052
rect 127854 28018 128190 28052
rect 128274 28018 128610 28052
rect 128694 28018 129030 28052
rect 129114 28018 129450 28052
rect 129534 28018 129870 28052
rect 129954 28018 130290 28052
rect 130374 28018 130710 28052
rect 130794 28018 131130 28052
rect 131214 28018 131550 28052
rect 131634 28018 131970 28052
rect 132054 28018 132390 28052
rect 132474 28018 132810 28052
rect 132894 28018 133230 28052
rect 133314 28018 133650 28052
rect 133734 28018 134070 28052
rect 134154 28018 134490 28052
rect 134574 28018 134910 28052
rect 134994 28018 135006 28052
rect 125964 28012 135006 28018
rect 125964 26952 126436 28012
rect 126876 27968 126922 27980
rect 126972 27968 127018 27980
rect 127086 27968 127132 27980
rect 127182 27968 127228 27980
rect 127296 27968 127342 27980
rect 127392 27968 127438 27980
rect 127506 27968 127552 27980
rect 127602 27968 127648 27980
rect 127716 27968 127762 27980
rect 127812 27968 127858 27980
rect 127926 27968 127972 27980
rect 128022 27968 128068 27980
rect 128136 27968 128182 27980
rect 128232 27968 128278 27980
rect 128346 27968 128392 27980
rect 128442 27968 128488 27980
rect 128556 27968 128602 27980
rect 128652 27968 128698 27980
rect 128766 27968 128812 27980
rect 128862 27968 128908 27980
rect 128976 27968 129022 27980
rect 129072 27968 129118 27980
rect 129186 27968 129232 27980
rect 129282 27968 129328 27980
rect 129396 27968 129442 27980
rect 129492 27968 129538 27980
rect 129606 27968 129652 27980
rect 129702 27968 129748 27980
rect 129816 27968 129862 27980
rect 129912 27968 129958 27980
rect 130026 27968 130072 27980
rect 130122 27968 130168 27980
rect 130236 27968 130282 27980
rect 130332 27968 130378 27980
rect 130446 27968 130492 27980
rect 130542 27968 130588 27980
rect 130656 27968 130702 27980
rect 130752 27968 130798 27980
rect 130866 27968 130912 27980
rect 130962 27968 131008 27980
rect 131076 27968 131122 27980
rect 131172 27968 131218 27980
rect 131286 27968 131332 27980
rect 131382 27968 131428 27980
rect 131496 27968 131542 27980
rect 131592 27968 131638 27980
rect 131706 27968 131752 27980
rect 131802 27968 131848 27980
rect 131916 27968 131962 27980
rect 132012 27968 132058 27980
rect 132126 27968 132172 27980
rect 132222 27968 132268 27980
rect 132336 27968 132382 27980
rect 132432 27968 132478 27980
rect 132546 27968 132592 27980
rect 132642 27968 132688 27980
rect 132756 27968 132802 27980
rect 132852 27968 132898 27980
rect 132966 27968 133012 27980
rect 133062 27968 133108 27980
rect 133176 27968 133222 27980
rect 133272 27968 133318 27980
rect 133386 27968 133432 27980
rect 133482 27968 133528 27980
rect 133596 27968 133642 27980
rect 133692 27968 133738 27980
rect 133806 27968 133852 27980
rect 133902 27968 133948 27980
rect 134016 27968 134062 27980
rect 134112 27968 134158 27980
rect 134226 27968 134272 27980
rect 134322 27968 134368 27980
rect 134436 27968 134482 27980
rect 134532 27968 134578 27980
rect 134646 27968 134692 27980
rect 134742 27968 134788 27980
rect 134856 27968 134902 27980
rect 134952 27968 134998 27980
rect 135066 27968 135112 27980
rect 135162 27968 135208 27980
rect 126848 26992 126858 27968
rect 126916 26992 126926 27968
rect 126968 26992 126978 27968
rect 127126 26992 127136 27968
rect 127178 26992 127188 27968
rect 127336 26992 127346 27968
rect 127388 26992 127398 27968
rect 127546 26992 127556 27968
rect 127598 26992 127608 27968
rect 127756 26992 127766 27968
rect 127808 26992 127818 27968
rect 127966 26992 127976 27968
rect 128018 26992 128028 27968
rect 128176 26992 128186 27968
rect 128228 26992 128238 27968
rect 128386 26992 128396 27968
rect 128438 26992 128448 27968
rect 128596 26992 128606 27968
rect 128648 26992 128658 27968
rect 128806 26992 128816 27968
rect 128858 26992 128868 27968
rect 129016 26992 129026 27968
rect 129068 26992 129078 27968
rect 129226 26992 129236 27968
rect 129278 26992 129288 27968
rect 129436 26992 129446 27968
rect 129488 26992 129498 27968
rect 129646 26992 129656 27968
rect 129698 26992 129708 27968
rect 129856 26992 129866 27968
rect 129908 26992 129918 27968
rect 130066 26992 130076 27968
rect 130118 26992 130128 27968
rect 130276 26992 130286 27968
rect 130328 26992 130338 27968
rect 130486 26992 130496 27968
rect 130538 26992 130548 27968
rect 130696 26992 130706 27968
rect 130748 26992 130758 27968
rect 130906 26992 130916 27968
rect 130958 26992 130968 27968
rect 131116 26992 131126 27968
rect 131168 26992 131178 27968
rect 131326 26992 131336 27968
rect 131378 26992 131388 27968
rect 131536 26992 131546 27968
rect 131588 26992 131598 27968
rect 131746 26992 131756 27968
rect 131798 26992 131808 27968
rect 131956 26992 131966 27968
rect 132008 26992 132018 27968
rect 132166 26992 132176 27968
rect 132218 26992 132228 27968
rect 132376 26992 132386 27968
rect 132428 26992 132438 27968
rect 132586 26992 132596 27968
rect 132638 26992 132648 27968
rect 132796 26992 132806 27968
rect 132848 26992 132858 27968
rect 133006 26992 133016 27968
rect 133058 26992 133068 27968
rect 133216 26992 133226 27968
rect 133268 26992 133278 27968
rect 133426 26992 133436 27968
rect 133478 26992 133488 27968
rect 133636 26992 133646 27968
rect 133688 26992 133698 27968
rect 133846 26992 133856 27968
rect 133898 26992 133908 27968
rect 134056 26992 134066 27968
rect 134108 26992 134118 27968
rect 134266 26992 134276 27968
rect 134318 26992 134328 27968
rect 134476 26992 134486 27968
rect 134528 26992 134538 27968
rect 134686 26992 134696 27968
rect 134738 26992 134748 27968
rect 134896 26992 134906 27968
rect 134948 26992 134958 27968
rect 135106 26992 135116 27968
rect 135158 26992 135168 27968
rect 135226 26992 135236 27968
rect 126876 26980 126922 26992
rect 126972 26980 127018 26992
rect 127086 26980 127132 26992
rect 127182 26980 127228 26992
rect 127296 26980 127342 26992
rect 127392 26980 127438 26992
rect 127506 26980 127552 26992
rect 127602 26980 127648 26992
rect 127716 26980 127762 26992
rect 127812 26980 127858 26992
rect 127926 26980 127972 26992
rect 128022 26980 128068 26992
rect 128136 26980 128182 26992
rect 128232 26980 128278 26992
rect 128346 26980 128392 26992
rect 128442 26980 128488 26992
rect 128556 26980 128602 26992
rect 128652 26980 128698 26992
rect 128766 26980 128812 26992
rect 128862 26980 128908 26992
rect 128976 26980 129022 26992
rect 129072 26980 129118 26992
rect 129186 26980 129232 26992
rect 129282 26980 129328 26992
rect 129396 26980 129442 26992
rect 129492 26980 129538 26992
rect 129606 26980 129652 26992
rect 129702 26980 129748 26992
rect 129816 26980 129862 26992
rect 129912 26980 129958 26992
rect 130026 26980 130072 26992
rect 130122 26980 130168 26992
rect 130236 26980 130282 26992
rect 130332 26980 130378 26992
rect 130446 26980 130492 26992
rect 130542 26980 130588 26992
rect 130656 26980 130702 26992
rect 130752 26980 130798 26992
rect 130866 26980 130912 26992
rect 130962 26980 131008 26992
rect 131076 26980 131122 26992
rect 131172 26980 131218 26992
rect 131286 26980 131332 26992
rect 131382 26980 131428 26992
rect 131496 26980 131542 26992
rect 131592 26980 131638 26992
rect 131706 26980 131752 26992
rect 131802 26980 131848 26992
rect 131916 26980 131962 26992
rect 132012 26980 132058 26992
rect 132126 26980 132172 26992
rect 132222 26980 132268 26992
rect 132336 26980 132382 26992
rect 132432 26980 132478 26992
rect 132546 26980 132592 26992
rect 132642 26980 132688 26992
rect 132756 26980 132802 26992
rect 132852 26980 132898 26992
rect 132966 26980 133012 26992
rect 133062 26980 133108 26992
rect 133176 26980 133222 26992
rect 133272 26980 133318 26992
rect 133386 26980 133432 26992
rect 133482 26980 133528 26992
rect 133596 26980 133642 26992
rect 133692 26980 133738 26992
rect 133806 26980 133852 26992
rect 133902 26980 133948 26992
rect 134016 26980 134062 26992
rect 134112 26980 134158 26992
rect 134226 26980 134272 26992
rect 134322 26980 134368 26992
rect 134436 26980 134482 26992
rect 134532 26980 134578 26992
rect 134646 26980 134692 26992
rect 134742 26980 134788 26992
rect 134856 26980 134902 26992
rect 134952 26980 134998 26992
rect 135066 26980 135112 26992
rect 135162 26980 135208 26992
rect 125964 26942 135166 26952
rect 125964 26800 127140 26942
rect 127174 26800 127560 26942
rect 127594 26800 127980 26942
rect 128014 26800 128400 26942
rect 128434 26800 128820 26942
rect 128854 26800 129240 26942
rect 129274 26800 129660 26942
rect 129694 26800 130080 26942
rect 130114 26800 130500 26942
rect 130534 26800 130920 26942
rect 130954 26800 131340 26942
rect 131374 26800 131760 26942
rect 131794 26800 132180 26942
rect 132214 26800 132600 26942
rect 132634 26800 133020 26942
rect 133054 26800 133440 26942
rect 133474 26800 133860 26942
rect 133894 26800 134280 26942
rect 134314 26800 134700 26942
rect 134734 26800 135120 26942
rect 135154 26800 135166 26942
rect 125964 26790 135166 26800
rect 125964 25730 126436 26790
rect 126876 26750 126922 26762
rect 126972 26750 127018 26762
rect 127086 26750 127132 26762
rect 127182 26750 127228 26762
rect 127296 26750 127342 26762
rect 127392 26750 127438 26762
rect 127506 26750 127552 26762
rect 127602 26750 127648 26762
rect 127716 26750 127762 26762
rect 127812 26750 127858 26762
rect 127926 26750 127972 26762
rect 128022 26750 128068 26762
rect 128136 26750 128182 26762
rect 128232 26750 128278 26762
rect 128346 26750 128392 26762
rect 128442 26750 128488 26762
rect 128556 26750 128602 26762
rect 128652 26750 128698 26762
rect 128766 26750 128812 26762
rect 128862 26750 128908 26762
rect 128976 26750 129022 26762
rect 129072 26750 129118 26762
rect 129186 26750 129232 26762
rect 129282 26750 129328 26762
rect 129396 26750 129442 26762
rect 129492 26750 129538 26762
rect 129606 26750 129652 26762
rect 129702 26750 129748 26762
rect 129816 26750 129862 26762
rect 129912 26750 129958 26762
rect 130026 26750 130072 26762
rect 130122 26750 130168 26762
rect 130236 26750 130282 26762
rect 130332 26750 130378 26762
rect 130446 26750 130492 26762
rect 130542 26750 130588 26762
rect 130656 26750 130702 26762
rect 130752 26750 130798 26762
rect 130866 26750 130912 26762
rect 130962 26750 131008 26762
rect 131076 26750 131122 26762
rect 131172 26750 131218 26762
rect 131286 26750 131332 26762
rect 131382 26750 131428 26762
rect 131496 26750 131542 26762
rect 131592 26750 131638 26762
rect 131706 26750 131752 26762
rect 131802 26750 131848 26762
rect 131916 26750 131962 26762
rect 132012 26750 132058 26762
rect 132126 26750 132172 26762
rect 132222 26750 132268 26762
rect 132336 26750 132382 26762
rect 132432 26750 132478 26762
rect 132546 26750 132592 26762
rect 132642 26750 132688 26762
rect 132756 26750 132802 26762
rect 132852 26750 132898 26762
rect 132966 26750 133012 26762
rect 133062 26750 133108 26762
rect 133176 26750 133222 26762
rect 133272 26750 133318 26762
rect 133386 26750 133432 26762
rect 133482 26750 133528 26762
rect 133596 26750 133642 26762
rect 133692 26750 133738 26762
rect 133806 26750 133852 26762
rect 133902 26750 133948 26762
rect 134016 26750 134062 26762
rect 134112 26750 134158 26762
rect 134226 26750 134272 26762
rect 134322 26750 134368 26762
rect 134436 26750 134482 26762
rect 134532 26750 134578 26762
rect 134646 26750 134692 26762
rect 134742 26750 134788 26762
rect 134856 26750 134902 26762
rect 134952 26750 134998 26762
rect 135066 26750 135112 26762
rect 135162 26750 135208 26762
rect 126848 25774 126858 26750
rect 126916 25774 126926 26750
rect 126968 25774 126978 26750
rect 127126 25774 127136 26750
rect 127178 25774 127188 26750
rect 127336 25774 127346 26750
rect 127388 25774 127398 26750
rect 127546 25774 127556 26750
rect 127598 25774 127608 26750
rect 127756 25774 127766 26750
rect 127808 25774 127818 26750
rect 127966 25774 127976 26750
rect 128018 25774 128028 26750
rect 128176 25774 128186 26750
rect 128228 25774 128238 26750
rect 128386 25774 128396 26750
rect 128438 25774 128448 26750
rect 128596 25774 128606 26750
rect 128648 25774 128658 26750
rect 128806 25774 128816 26750
rect 128858 25774 128868 26750
rect 129016 25774 129026 26750
rect 129068 25774 129078 26750
rect 129226 25774 129236 26750
rect 129278 25774 129288 26750
rect 129436 25774 129446 26750
rect 129488 25774 129498 26750
rect 129646 25774 129656 26750
rect 129698 25774 129708 26750
rect 129856 25774 129866 26750
rect 129908 25774 129918 26750
rect 130066 25774 130076 26750
rect 130118 25774 130128 26750
rect 130276 25774 130286 26750
rect 130328 25774 130338 26750
rect 130486 25774 130496 26750
rect 130538 25774 130548 26750
rect 130696 25774 130706 26750
rect 130748 25774 130758 26750
rect 130906 25774 130916 26750
rect 130958 25774 130968 26750
rect 131116 25774 131126 26750
rect 131168 25774 131178 26750
rect 131326 25774 131336 26750
rect 131378 25774 131388 26750
rect 131536 25774 131546 26750
rect 131588 25774 131598 26750
rect 131746 25774 131756 26750
rect 131798 25774 131808 26750
rect 131956 25774 131966 26750
rect 132008 25774 132018 26750
rect 132166 25774 132176 26750
rect 132218 25774 132228 26750
rect 132376 25774 132386 26750
rect 132428 25774 132438 26750
rect 132586 25774 132596 26750
rect 132638 25774 132648 26750
rect 132796 25774 132806 26750
rect 132848 25774 132858 26750
rect 133006 25774 133016 26750
rect 133058 25774 133068 26750
rect 133216 25774 133226 26750
rect 133268 25774 133278 26750
rect 133426 25774 133436 26750
rect 133478 25774 133488 26750
rect 133636 25774 133646 26750
rect 133688 25774 133698 26750
rect 133846 25774 133856 26750
rect 133898 25774 133908 26750
rect 134056 25774 134066 26750
rect 134108 25774 134118 26750
rect 134266 25774 134276 26750
rect 134318 25774 134328 26750
rect 134476 25774 134486 26750
rect 134528 25774 134538 26750
rect 134686 25774 134696 26750
rect 134738 25774 134748 26750
rect 134896 25774 134906 26750
rect 134948 25774 134958 26750
rect 135106 25774 135116 26750
rect 135158 25774 135168 26750
rect 135226 25774 135236 26750
rect 126876 25762 126922 25774
rect 126972 25762 127018 25774
rect 127086 25762 127132 25774
rect 127182 25762 127228 25774
rect 127296 25762 127342 25774
rect 127392 25762 127438 25774
rect 127506 25762 127552 25774
rect 127602 25762 127648 25774
rect 127716 25762 127762 25774
rect 127812 25762 127858 25774
rect 127926 25762 127972 25774
rect 128022 25762 128068 25774
rect 128136 25762 128182 25774
rect 128232 25762 128278 25774
rect 128346 25762 128392 25774
rect 128442 25762 128488 25774
rect 128556 25762 128602 25774
rect 128652 25762 128698 25774
rect 128766 25762 128812 25774
rect 128862 25762 128908 25774
rect 128976 25762 129022 25774
rect 129072 25762 129118 25774
rect 129186 25762 129232 25774
rect 129282 25762 129328 25774
rect 129396 25762 129442 25774
rect 129492 25762 129538 25774
rect 129606 25762 129652 25774
rect 129702 25762 129748 25774
rect 129816 25762 129862 25774
rect 129912 25762 129958 25774
rect 130026 25762 130072 25774
rect 130122 25762 130168 25774
rect 130236 25762 130282 25774
rect 130332 25762 130378 25774
rect 130446 25762 130492 25774
rect 130542 25762 130588 25774
rect 130656 25762 130702 25774
rect 130752 25762 130798 25774
rect 130866 25762 130912 25774
rect 130962 25762 131008 25774
rect 131076 25762 131122 25774
rect 131172 25762 131218 25774
rect 131286 25762 131332 25774
rect 131382 25762 131428 25774
rect 131496 25762 131542 25774
rect 131592 25762 131638 25774
rect 131706 25762 131752 25774
rect 131802 25762 131848 25774
rect 131916 25762 131962 25774
rect 132012 25762 132058 25774
rect 132126 25762 132172 25774
rect 132222 25762 132268 25774
rect 132336 25762 132382 25774
rect 132432 25762 132478 25774
rect 132546 25762 132592 25774
rect 132642 25762 132688 25774
rect 132756 25762 132802 25774
rect 132852 25762 132898 25774
rect 132966 25762 133012 25774
rect 133062 25762 133108 25774
rect 133176 25762 133222 25774
rect 133272 25762 133318 25774
rect 133386 25762 133432 25774
rect 133482 25762 133528 25774
rect 133596 25762 133642 25774
rect 133692 25762 133738 25774
rect 133806 25762 133852 25774
rect 133902 25762 133948 25774
rect 134016 25762 134062 25774
rect 134112 25762 134158 25774
rect 134226 25762 134272 25774
rect 134322 25762 134368 25774
rect 134436 25762 134482 25774
rect 134532 25762 134578 25774
rect 134646 25762 134692 25774
rect 134742 25762 134788 25774
rect 134856 25762 134902 25774
rect 134952 25762 134998 25774
rect 135066 25762 135112 25774
rect 135162 25762 135208 25774
rect 125964 25724 135006 25730
rect 125964 25690 126930 25724
rect 127014 25690 127350 25724
rect 127434 25690 127770 25724
rect 127854 25690 128190 25724
rect 128274 25690 128610 25724
rect 128694 25690 129030 25724
rect 129114 25690 129450 25724
rect 129534 25690 129870 25724
rect 129954 25690 130290 25724
rect 130374 25690 130710 25724
rect 130794 25690 131130 25724
rect 131214 25690 131550 25724
rect 131634 25690 131970 25724
rect 132054 25690 132390 25724
rect 132474 25690 132810 25724
rect 132894 25690 133230 25724
rect 133314 25690 133650 25724
rect 133734 25690 134070 25724
rect 134154 25690 134490 25724
rect 134574 25690 134910 25724
rect 134994 25690 135006 25724
rect 125964 25684 135006 25690
rect 125964 22840 126436 25684
rect 125964 22833 135006 22840
rect 125964 22798 126930 22833
rect 126964 22832 127350 22833
rect 127384 22832 127770 22833
rect 127804 22832 128190 22833
rect 128224 22832 128610 22833
rect 128644 22832 129030 22833
rect 129064 22832 129450 22833
rect 129484 22832 129870 22833
rect 129904 22832 130290 22833
rect 130324 22832 130710 22833
rect 130744 22832 131130 22833
rect 131164 22832 131550 22833
rect 131584 22832 131970 22833
rect 132004 22832 132390 22833
rect 132424 22832 132810 22833
rect 132844 22832 133230 22833
rect 133264 22832 133650 22833
rect 133684 22832 134070 22833
rect 134104 22832 134490 22833
rect 134524 22832 134910 22833
rect 134944 22832 135006 22833
rect 127014 22798 127350 22832
rect 127434 22798 127770 22832
rect 127854 22798 128190 22832
rect 128274 22798 128610 22832
rect 128694 22798 129030 22832
rect 129114 22798 129450 22832
rect 129534 22798 129870 22832
rect 129954 22798 130290 22832
rect 130374 22798 130710 22832
rect 130794 22798 131130 22832
rect 131214 22798 131550 22832
rect 131634 22798 131970 22832
rect 132054 22798 132390 22832
rect 132474 22798 132810 22832
rect 132894 22798 133230 22832
rect 133314 22798 133650 22832
rect 133734 22798 134070 22832
rect 134154 22798 134490 22832
rect 134574 22798 134910 22832
rect 134994 22798 135006 22832
rect 125964 22790 135006 22798
rect 122016 22162 122140 22168
rect 122016 22062 122028 22162
rect 122128 22062 122140 22162
rect 122016 22056 122140 22062
rect 122436 22162 122560 22168
rect 122436 22062 122448 22162
rect 122548 22062 122560 22162
rect 122436 22056 122560 22062
rect 122856 22162 122980 22168
rect 122856 22062 122868 22162
rect 122968 22062 122980 22162
rect 122856 22056 122980 22062
rect 123276 22162 123400 22168
rect 123276 22062 123288 22162
rect 123388 22062 123400 22162
rect 123276 22056 123400 22062
rect 123696 22162 123820 22168
rect 123696 22062 123708 22162
rect 123808 22062 123820 22162
rect 123696 22056 123820 22062
rect 124116 22162 124240 22168
rect 124116 22062 124128 22162
rect 124228 22062 124240 22162
rect 124116 22056 124240 22062
rect 124536 22162 124660 22168
rect 124536 22062 124548 22162
rect 124648 22062 124660 22162
rect 124536 22056 124660 22062
rect 124956 22162 125080 22168
rect 124956 22062 124968 22162
rect 125068 22062 125080 22162
rect 124956 22056 125080 22062
rect 125376 22162 125500 22168
rect 125376 22062 125388 22162
rect 125488 22062 125500 22162
rect 125376 22056 125500 22062
rect 125702 22162 125826 22168
rect 125702 22062 125714 22162
rect 125814 22062 125826 22162
rect 125702 22056 125826 22062
rect 121590 21976 125750 21984
rect 121590 21942 122290 21976
rect 122374 21942 122710 21976
rect 122794 21942 123130 21976
rect 123214 21942 123550 21976
rect 123634 21942 123970 21976
rect 124054 21942 124390 21976
rect 124474 21942 124810 21976
rect 124894 21942 125230 21976
rect 125314 21942 125650 21976
rect 125734 21942 125750 21976
rect 121590 21934 122710 21942
rect 122744 21934 123130 21942
rect 123164 21934 123550 21942
rect 123584 21934 123970 21942
rect 124004 21934 124390 21942
rect 124424 21934 124810 21942
rect 124844 21934 125230 21942
rect 125264 21934 125650 21942
rect 125684 21934 125750 21942
rect 121590 21928 125750 21934
rect 121590 20864 121776 21928
rect 122026 21884 122072 21896
rect 122122 21884 122168 21896
rect 122236 21884 122282 21896
rect 122332 21884 122378 21896
rect 122446 21884 122492 21896
rect 122542 21884 122588 21896
rect 122656 21884 122702 21896
rect 122752 21884 122798 21896
rect 122866 21884 122912 21896
rect 122962 21884 123008 21896
rect 123076 21884 123122 21896
rect 123172 21884 123218 21896
rect 123286 21884 123332 21896
rect 123382 21884 123428 21896
rect 123496 21884 123542 21896
rect 123592 21884 123638 21896
rect 123706 21884 123752 21896
rect 123802 21884 123848 21896
rect 123916 21884 123962 21896
rect 124012 21884 124058 21896
rect 124126 21884 124172 21896
rect 124222 21884 124268 21896
rect 124336 21884 124382 21896
rect 124432 21884 124478 21896
rect 124546 21884 124592 21896
rect 124642 21884 124688 21896
rect 124756 21884 124802 21896
rect 124852 21884 124898 21896
rect 124966 21884 125012 21896
rect 125062 21884 125108 21896
rect 125176 21884 125222 21896
rect 125272 21884 125318 21896
rect 125386 21884 125432 21896
rect 125482 21884 125528 21896
rect 125596 21884 125642 21896
rect 125692 21884 125738 21896
rect 121998 20908 122008 21884
rect 122066 20908 122076 21884
rect 122118 20908 122128 21884
rect 122276 20908 122286 21884
rect 122328 20908 122338 21884
rect 122486 20908 122496 21884
rect 122538 20908 122548 21884
rect 122696 20908 122706 21884
rect 122748 20908 122758 21884
rect 122906 20908 122916 21884
rect 122958 20908 122968 21884
rect 123116 20908 123126 21884
rect 123168 20908 123178 21884
rect 123326 20908 123336 21884
rect 123378 20908 123388 21884
rect 123536 20908 123546 21884
rect 123588 20908 123598 21884
rect 123746 20908 123756 21884
rect 123798 20908 123808 21884
rect 123956 20908 123966 21884
rect 124008 20908 124018 21884
rect 124166 20908 124176 21884
rect 124218 20908 124228 21884
rect 124376 20908 124386 21884
rect 124428 20908 124438 21884
rect 124586 20908 124596 21884
rect 124638 20908 124648 21884
rect 124796 20908 124806 21884
rect 124848 20908 124858 21884
rect 125006 20908 125016 21884
rect 125058 20908 125068 21884
rect 125216 20908 125226 21884
rect 125268 20908 125278 21884
rect 125426 20908 125436 21884
rect 125478 20908 125488 21884
rect 125636 20908 125646 21884
rect 125688 20908 125698 21884
rect 125756 20908 125766 21884
rect 125964 21712 126436 22790
rect 126876 22740 126922 22752
rect 126972 22740 127018 22752
rect 127086 22740 127132 22752
rect 127182 22740 127228 22752
rect 127296 22740 127342 22752
rect 127392 22740 127438 22752
rect 127506 22740 127552 22752
rect 127602 22740 127648 22752
rect 127716 22740 127762 22752
rect 127812 22740 127858 22752
rect 127926 22740 127972 22752
rect 128022 22740 128068 22752
rect 128136 22740 128182 22752
rect 128232 22740 128278 22752
rect 128346 22740 128392 22752
rect 128442 22740 128488 22752
rect 128556 22740 128602 22752
rect 128652 22740 128698 22752
rect 128766 22740 128812 22752
rect 128862 22740 128908 22752
rect 128976 22740 129022 22752
rect 129072 22740 129118 22752
rect 129186 22740 129232 22752
rect 129282 22740 129328 22752
rect 129396 22740 129442 22752
rect 129492 22740 129538 22752
rect 129606 22740 129652 22752
rect 129702 22740 129748 22752
rect 129816 22740 129862 22752
rect 129912 22740 129958 22752
rect 130026 22740 130072 22752
rect 130122 22740 130168 22752
rect 130236 22740 130282 22752
rect 130332 22740 130378 22752
rect 130446 22740 130492 22752
rect 130542 22740 130588 22752
rect 130656 22740 130702 22752
rect 130752 22740 130798 22752
rect 130866 22740 130912 22752
rect 130962 22740 131008 22752
rect 131076 22740 131122 22752
rect 131172 22740 131218 22752
rect 131286 22740 131332 22752
rect 131382 22740 131428 22752
rect 131496 22740 131542 22752
rect 131592 22740 131638 22752
rect 131706 22740 131752 22752
rect 131802 22740 131848 22752
rect 131916 22740 131962 22752
rect 132012 22740 132058 22752
rect 132126 22740 132172 22752
rect 132222 22740 132268 22752
rect 132336 22740 132382 22752
rect 132432 22740 132478 22752
rect 132546 22740 132592 22752
rect 132642 22740 132688 22752
rect 132756 22740 132802 22752
rect 132852 22740 132898 22752
rect 132966 22740 133012 22752
rect 133062 22740 133108 22752
rect 133176 22740 133222 22752
rect 133272 22740 133318 22752
rect 133386 22740 133432 22752
rect 133482 22740 133528 22752
rect 133596 22740 133642 22752
rect 133692 22740 133738 22752
rect 133806 22740 133852 22752
rect 133902 22740 133948 22752
rect 134016 22740 134062 22752
rect 134112 22740 134158 22752
rect 134226 22740 134272 22752
rect 134322 22740 134368 22752
rect 134436 22740 134482 22752
rect 134532 22740 134578 22752
rect 134646 22740 134692 22752
rect 134742 22740 134788 22752
rect 134856 22740 134902 22752
rect 134952 22740 134998 22752
rect 135066 22740 135112 22752
rect 135162 22740 135208 22752
rect 126848 21764 126858 22740
rect 126916 21764 126926 22740
rect 126968 21764 126978 22740
rect 127126 21764 127136 22740
rect 127178 21764 127188 22740
rect 127336 21764 127346 22740
rect 127388 21764 127398 22740
rect 127546 21764 127556 22740
rect 127598 21764 127608 22740
rect 127756 21764 127766 22740
rect 127808 21764 127818 22740
rect 127966 21764 127976 22740
rect 128018 21764 128028 22740
rect 128176 21764 128186 22740
rect 128228 21764 128238 22740
rect 128386 21764 128396 22740
rect 128438 21764 128448 22740
rect 128596 21764 128606 22740
rect 128648 21764 128658 22740
rect 128806 21764 128816 22740
rect 128858 21764 128868 22740
rect 129016 21764 129026 22740
rect 129068 21764 129078 22740
rect 129226 21764 129236 22740
rect 129278 21764 129288 22740
rect 129436 21764 129446 22740
rect 129488 21764 129498 22740
rect 129646 21764 129656 22740
rect 129698 21764 129708 22740
rect 129856 21764 129866 22740
rect 129908 21764 129918 22740
rect 130066 21764 130076 22740
rect 130118 21764 130128 22740
rect 130276 21764 130286 22740
rect 130328 21764 130338 22740
rect 130486 21764 130496 22740
rect 130538 21764 130548 22740
rect 130696 21764 130706 22740
rect 130748 21764 130758 22740
rect 130906 21764 130916 22740
rect 130958 21764 130968 22740
rect 131116 21764 131126 22740
rect 131168 21764 131178 22740
rect 131326 21764 131336 22740
rect 131378 21764 131388 22740
rect 131536 21764 131546 22740
rect 131588 21764 131598 22740
rect 131746 21764 131756 22740
rect 131798 21764 131808 22740
rect 131956 21764 131966 22740
rect 132008 21764 132018 22740
rect 132166 21764 132176 22740
rect 132218 21764 132228 22740
rect 132376 21764 132386 22740
rect 132428 21764 132438 22740
rect 132586 21764 132596 22740
rect 132638 21764 132648 22740
rect 132796 21764 132806 22740
rect 132848 21764 132858 22740
rect 133006 21764 133016 22740
rect 133058 21764 133068 22740
rect 133216 21764 133226 22740
rect 133268 21764 133278 22740
rect 133426 21764 133436 22740
rect 133478 21764 133488 22740
rect 133636 21764 133646 22740
rect 133688 21764 133698 22740
rect 133846 21764 133856 22740
rect 133898 21764 133908 22740
rect 134056 21764 134066 22740
rect 134108 21764 134118 22740
rect 134266 21764 134276 22740
rect 134318 21764 134328 22740
rect 134476 21764 134486 22740
rect 134528 21764 134538 22740
rect 134686 21764 134696 22740
rect 134738 21764 134748 22740
rect 134896 21764 134906 22740
rect 134948 21764 134958 22740
rect 135106 21764 135116 22740
rect 135158 21764 135168 22740
rect 135226 21764 135236 22740
rect 126876 21752 126922 21764
rect 126972 21752 127018 21764
rect 127086 21752 127132 21764
rect 127182 21752 127228 21764
rect 127296 21752 127342 21764
rect 127392 21752 127438 21764
rect 127506 21752 127552 21764
rect 127602 21752 127648 21764
rect 127716 21752 127762 21764
rect 127812 21752 127858 21764
rect 127926 21752 127972 21764
rect 128022 21752 128068 21764
rect 128136 21752 128182 21764
rect 128232 21752 128278 21764
rect 128346 21752 128392 21764
rect 128442 21752 128488 21764
rect 128556 21752 128602 21764
rect 128652 21752 128698 21764
rect 128766 21752 128812 21764
rect 128862 21752 128908 21764
rect 128976 21752 129022 21764
rect 129072 21752 129118 21764
rect 129186 21752 129232 21764
rect 129282 21752 129328 21764
rect 129396 21752 129442 21764
rect 129492 21752 129538 21764
rect 129606 21752 129652 21764
rect 129702 21752 129748 21764
rect 129816 21752 129862 21764
rect 129912 21752 129958 21764
rect 130026 21752 130072 21764
rect 130122 21752 130168 21764
rect 130236 21752 130282 21764
rect 130332 21752 130378 21764
rect 130446 21752 130492 21764
rect 130542 21752 130588 21764
rect 130656 21752 130702 21764
rect 130752 21752 130798 21764
rect 130866 21752 130912 21764
rect 130962 21752 131008 21764
rect 131076 21752 131122 21764
rect 131172 21752 131218 21764
rect 131286 21752 131332 21764
rect 131382 21752 131428 21764
rect 131496 21752 131542 21764
rect 131592 21752 131638 21764
rect 131706 21752 131752 21764
rect 131802 21752 131848 21764
rect 131916 21752 131962 21764
rect 132012 21752 132058 21764
rect 132126 21752 132172 21764
rect 132222 21752 132268 21764
rect 132336 21752 132382 21764
rect 132432 21752 132478 21764
rect 132546 21752 132592 21764
rect 132642 21752 132688 21764
rect 132756 21752 132802 21764
rect 132852 21752 132898 21764
rect 132966 21752 133012 21764
rect 133062 21752 133108 21764
rect 133176 21752 133222 21764
rect 133272 21752 133318 21764
rect 133386 21752 133432 21764
rect 133482 21752 133528 21764
rect 133596 21752 133642 21764
rect 133692 21752 133738 21764
rect 133806 21752 133852 21764
rect 133902 21752 133948 21764
rect 134016 21752 134062 21764
rect 134112 21752 134158 21764
rect 134226 21752 134272 21764
rect 134322 21752 134368 21764
rect 134436 21752 134482 21764
rect 134532 21752 134578 21764
rect 134646 21752 134692 21764
rect 134742 21752 134788 21764
rect 134856 21752 134902 21764
rect 134952 21752 134998 21764
rect 135066 21752 135112 21764
rect 135162 21752 135208 21764
rect 125964 21705 135166 21712
rect 125964 21563 127140 21705
rect 127174 21563 127560 21705
rect 127594 21563 127980 21705
rect 128014 21563 128400 21705
rect 128434 21563 128820 21705
rect 128854 21563 129240 21705
rect 129274 21563 129660 21705
rect 129694 21563 130080 21705
rect 130114 21563 130500 21705
rect 130534 21563 130920 21705
rect 130954 21563 131340 21705
rect 131374 21563 131760 21705
rect 131794 21563 132180 21705
rect 132214 21563 132600 21705
rect 132634 21563 133020 21705
rect 133054 21563 133440 21705
rect 133474 21563 133860 21705
rect 133894 21563 134280 21705
rect 134314 21563 134700 21705
rect 134734 21563 135120 21705
rect 135154 21563 135166 21705
rect 125964 21556 135166 21563
rect 125964 20928 126436 21556
rect 126876 21504 126922 21516
rect 126972 21504 127018 21516
rect 127086 21504 127132 21516
rect 127182 21504 127228 21516
rect 127296 21504 127342 21516
rect 127392 21504 127438 21516
rect 127506 21504 127552 21516
rect 127602 21504 127648 21516
rect 127716 21504 127762 21516
rect 127812 21504 127858 21516
rect 127926 21504 127972 21516
rect 128022 21504 128068 21516
rect 128136 21504 128182 21516
rect 128232 21504 128278 21516
rect 128346 21504 128392 21516
rect 128442 21504 128488 21516
rect 128556 21504 128602 21516
rect 128652 21504 128698 21516
rect 128766 21504 128812 21516
rect 128862 21504 128908 21516
rect 128976 21504 129022 21516
rect 129072 21504 129118 21516
rect 129186 21504 129232 21516
rect 129282 21504 129328 21516
rect 129396 21504 129442 21516
rect 129492 21504 129538 21516
rect 129606 21504 129652 21516
rect 129702 21504 129748 21516
rect 129816 21504 129862 21516
rect 129912 21504 129958 21516
rect 130026 21504 130072 21516
rect 130122 21504 130168 21516
rect 130236 21504 130282 21516
rect 130332 21504 130378 21516
rect 130446 21504 130492 21516
rect 130542 21504 130588 21516
rect 130656 21504 130702 21516
rect 130752 21504 130798 21516
rect 130866 21504 130912 21516
rect 130962 21504 131008 21516
rect 131076 21504 131122 21516
rect 131172 21504 131218 21516
rect 131286 21504 131332 21516
rect 131382 21504 131428 21516
rect 131496 21504 131542 21516
rect 131592 21504 131638 21516
rect 131706 21504 131752 21516
rect 131802 21504 131848 21516
rect 131916 21504 131962 21516
rect 132012 21504 132058 21516
rect 132126 21504 132172 21516
rect 132222 21504 132268 21516
rect 132336 21504 132382 21516
rect 132432 21504 132478 21516
rect 132546 21504 132592 21516
rect 132642 21504 132688 21516
rect 132756 21504 132802 21516
rect 132852 21504 132898 21516
rect 132966 21504 133012 21516
rect 133062 21504 133108 21516
rect 133176 21504 133222 21516
rect 133272 21504 133318 21516
rect 133386 21504 133432 21516
rect 133482 21504 133528 21516
rect 133596 21504 133642 21516
rect 133692 21504 133738 21516
rect 133806 21504 133852 21516
rect 133902 21504 133948 21516
rect 134016 21504 134062 21516
rect 134112 21504 134158 21516
rect 134226 21504 134272 21516
rect 134322 21504 134368 21516
rect 134436 21504 134482 21516
rect 134532 21504 134578 21516
rect 134646 21504 134692 21516
rect 134742 21504 134788 21516
rect 134856 21504 134902 21516
rect 134952 21504 134998 21516
rect 135066 21504 135112 21516
rect 135162 21504 135208 21516
rect 122026 20896 122072 20908
rect 122122 20896 122168 20908
rect 122236 20896 122282 20908
rect 122332 20896 122378 20908
rect 122446 20896 122492 20908
rect 122542 20896 122588 20908
rect 122656 20896 122702 20908
rect 122752 20896 122798 20908
rect 122866 20896 122912 20908
rect 122962 20896 123008 20908
rect 123076 20896 123122 20908
rect 123172 20896 123218 20908
rect 123286 20896 123332 20908
rect 123382 20896 123428 20908
rect 123496 20896 123542 20908
rect 123592 20896 123638 20908
rect 123706 20896 123752 20908
rect 123802 20896 123848 20908
rect 123916 20896 123962 20908
rect 124012 20896 124058 20908
rect 124126 20896 124172 20908
rect 124222 20896 124268 20908
rect 124336 20896 124382 20908
rect 124432 20896 124478 20908
rect 124546 20896 124592 20908
rect 124642 20896 124688 20908
rect 124756 20896 124802 20908
rect 124852 20896 124898 20908
rect 124966 20896 125012 20908
rect 125062 20896 125108 20908
rect 125176 20896 125222 20908
rect 125272 20896 125318 20908
rect 125386 20896 125432 20908
rect 125482 20896 125528 20908
rect 125596 20896 125642 20908
rect 125692 20896 125738 20908
rect 121590 20858 125636 20864
rect 121590 20853 122920 20858
rect 121590 20818 122080 20853
rect 122114 20852 122500 20853
rect 122534 20852 122920 20853
rect 122954 20852 123340 20858
rect 123374 20852 123760 20858
rect 123794 20852 124180 20858
rect 124214 20852 124600 20858
rect 124634 20852 125020 20858
rect 125054 20852 125440 20858
rect 125474 20852 125636 20858
rect 122164 20818 122500 20852
rect 122584 20818 122920 20852
rect 123004 20818 123340 20852
rect 123424 20818 123760 20852
rect 123844 20818 124180 20852
rect 124264 20818 124600 20852
rect 124684 20818 125020 20852
rect 125104 20818 125440 20852
rect 125524 20818 125636 20852
rect 121590 20804 125636 20818
rect 119476 20730 119798 20736
rect 119476 20448 119488 20730
rect 119786 20448 119798 20730
rect 119476 20442 119798 20448
rect 121590 20368 121776 20804
rect 121590 20361 125636 20368
rect 119322 20353 120842 20360
rect 119322 20318 120326 20353
rect 120360 20352 120746 20353
rect 120780 20352 120842 20353
rect 120410 20318 120746 20352
rect 120830 20318 120842 20352
rect 119322 20304 120842 20318
rect 121590 20326 122080 20361
rect 122114 20360 122500 20361
rect 122534 20360 122920 20361
rect 122954 20360 123340 20361
rect 123374 20360 123760 20361
rect 123794 20360 124180 20361
rect 124214 20360 124600 20361
rect 124634 20360 125020 20361
rect 125054 20360 125440 20361
rect 125474 20360 125636 20361
rect 122164 20326 122500 20360
rect 122584 20326 122920 20360
rect 123004 20326 123340 20360
rect 123424 20326 123760 20360
rect 123844 20326 124180 20360
rect 124264 20326 124600 20360
rect 124684 20326 125020 20360
rect 125104 20326 125440 20360
rect 125524 20326 125636 20360
rect 121590 20318 125636 20326
rect 119118 20260 119164 20272
rect 119206 20260 119252 20272
rect 119094 19284 119104 20260
rect 119158 19284 119168 20260
rect 119202 19284 119212 20260
rect 119266 19284 119276 20260
rect 119322 19336 119436 20304
rect 120062 20260 120108 20272
rect 120158 20260 120204 20272
rect 120272 20260 120318 20272
rect 120368 20260 120414 20272
rect 120482 20260 120528 20272
rect 120578 20260 120624 20272
rect 120692 20260 120738 20272
rect 120788 20260 120834 20272
rect 119118 19272 119164 19284
rect 119206 19272 119252 19284
rect 119156 19234 119214 19240
rect 119156 19182 119168 19234
rect 118766 19134 119168 19182
rect 118766 18004 118860 19134
rect 119156 19091 119168 19134
rect 119202 19091 119214 19234
rect 119322 19188 119332 19336
rect 119474 19206 119484 19336
rect 120038 19284 120048 20260
rect 120102 19284 120112 20260
rect 120154 19284 120164 20260
rect 120312 19284 120322 20260
rect 120364 19284 120374 20260
rect 120522 19284 120532 20260
rect 120574 19284 120584 20260
rect 120732 19284 120742 20260
rect 120784 19284 120794 20260
rect 120848 19284 120858 20260
rect 121254 19432 121264 19696
rect 121546 19668 121556 19696
rect 121590 19668 121776 20318
rect 125854 20310 125864 20928
rect 126474 20476 126484 20928
rect 126848 20528 126858 21504
rect 126916 20528 126926 21504
rect 126968 20528 126978 21504
rect 127126 20528 127136 21504
rect 127178 20528 127188 21504
rect 127336 20528 127346 21504
rect 127388 20528 127398 21504
rect 127546 20528 127556 21504
rect 127598 20528 127608 21504
rect 127756 20528 127766 21504
rect 127808 20528 127818 21504
rect 127966 20528 127976 21504
rect 128018 20528 128028 21504
rect 128176 20528 128186 21504
rect 128228 20528 128238 21504
rect 128386 20528 128396 21504
rect 128438 20528 128448 21504
rect 128596 20528 128606 21504
rect 128648 20528 128658 21504
rect 128806 20528 128816 21504
rect 128858 20528 128868 21504
rect 129016 20528 129026 21504
rect 129068 20528 129078 21504
rect 129226 20528 129236 21504
rect 129278 20528 129288 21504
rect 129436 20528 129446 21504
rect 129488 20528 129498 21504
rect 129646 20528 129656 21504
rect 129698 20528 129708 21504
rect 129856 20528 129866 21504
rect 129908 20528 129918 21504
rect 130066 20528 130076 21504
rect 130118 20528 130128 21504
rect 130276 20528 130286 21504
rect 130328 20528 130338 21504
rect 130486 20528 130496 21504
rect 130538 20528 130548 21504
rect 130696 20528 130706 21504
rect 130748 20528 130758 21504
rect 130906 20528 130916 21504
rect 130958 20528 130968 21504
rect 131116 20528 131126 21504
rect 131168 20528 131178 21504
rect 131326 20528 131336 21504
rect 131378 20528 131388 21504
rect 131536 20528 131546 21504
rect 131588 20528 131598 21504
rect 131746 20528 131756 21504
rect 131798 20528 131808 21504
rect 131956 20528 131966 21504
rect 132008 20528 132018 21504
rect 132166 20528 132176 21504
rect 132218 20528 132228 21504
rect 132376 20528 132386 21504
rect 132428 20528 132438 21504
rect 132586 20528 132596 21504
rect 132638 20528 132648 21504
rect 132796 20528 132806 21504
rect 132848 20528 132858 21504
rect 133006 20528 133016 21504
rect 133058 20528 133068 21504
rect 133216 20528 133226 21504
rect 133268 20528 133278 21504
rect 133426 20528 133436 21504
rect 133478 20528 133488 21504
rect 133636 20528 133646 21504
rect 133688 20528 133698 21504
rect 133846 20528 133856 21504
rect 133898 20528 133908 21504
rect 134056 20528 134066 21504
rect 134108 20528 134118 21504
rect 134266 20528 134276 21504
rect 134318 20528 134328 21504
rect 134476 20528 134486 21504
rect 134528 20528 134538 21504
rect 134686 20528 134696 21504
rect 134738 20528 134748 21504
rect 134896 20528 134906 21504
rect 134948 20528 134958 21504
rect 135106 20528 135116 21504
rect 135158 20528 135168 21504
rect 135226 20528 135236 21504
rect 126876 20516 126922 20528
rect 126972 20516 127018 20528
rect 127086 20516 127132 20528
rect 127182 20516 127228 20528
rect 127296 20516 127342 20528
rect 127392 20516 127438 20528
rect 127506 20516 127552 20528
rect 127602 20516 127648 20528
rect 127716 20516 127762 20528
rect 127812 20516 127858 20528
rect 127926 20516 127972 20528
rect 128022 20516 128068 20528
rect 128136 20516 128182 20528
rect 128232 20516 128278 20528
rect 128346 20516 128392 20528
rect 128442 20516 128488 20528
rect 128556 20516 128602 20528
rect 128652 20516 128698 20528
rect 128766 20516 128812 20528
rect 128862 20516 128908 20528
rect 128976 20516 129022 20528
rect 129072 20516 129118 20528
rect 129186 20516 129232 20528
rect 129282 20516 129328 20528
rect 129396 20516 129442 20528
rect 129492 20516 129538 20528
rect 129606 20516 129652 20528
rect 129702 20516 129748 20528
rect 129816 20516 129862 20528
rect 129912 20516 129958 20528
rect 130026 20516 130072 20528
rect 130122 20516 130168 20528
rect 130236 20516 130282 20528
rect 130332 20516 130378 20528
rect 130446 20516 130492 20528
rect 130542 20516 130588 20528
rect 130656 20516 130702 20528
rect 130752 20516 130798 20528
rect 130866 20516 130912 20528
rect 130962 20516 131008 20528
rect 131076 20516 131122 20528
rect 131172 20516 131218 20528
rect 131286 20516 131332 20528
rect 131382 20516 131428 20528
rect 131496 20516 131542 20528
rect 131592 20516 131638 20528
rect 131706 20516 131752 20528
rect 131802 20516 131848 20528
rect 131916 20516 131962 20528
rect 132012 20516 132058 20528
rect 132126 20516 132172 20528
rect 132222 20516 132268 20528
rect 132336 20516 132382 20528
rect 132432 20516 132478 20528
rect 132546 20516 132592 20528
rect 132642 20516 132688 20528
rect 132756 20516 132802 20528
rect 132852 20516 132898 20528
rect 132966 20516 133012 20528
rect 133062 20516 133108 20528
rect 133176 20516 133222 20528
rect 133272 20516 133318 20528
rect 133386 20516 133432 20528
rect 133482 20516 133528 20528
rect 133596 20516 133642 20528
rect 133692 20516 133738 20528
rect 133806 20516 133852 20528
rect 133902 20516 133948 20528
rect 134016 20516 134062 20528
rect 134112 20516 134158 20528
rect 134226 20516 134272 20528
rect 134322 20516 134368 20528
rect 134436 20516 134482 20528
rect 134532 20516 134578 20528
rect 134646 20516 134692 20528
rect 134742 20516 134788 20528
rect 134856 20516 134902 20528
rect 134952 20516 134998 20528
rect 135066 20516 135112 20528
rect 135162 20516 135208 20528
rect 126474 20469 134956 20476
rect 126474 20327 126930 20469
rect 126964 20327 127350 20469
rect 127384 20327 127770 20469
rect 127804 20327 128190 20469
rect 128224 20327 128610 20469
rect 128644 20327 129030 20469
rect 129064 20327 129450 20469
rect 129484 20327 129870 20469
rect 129904 20327 130290 20469
rect 130324 20327 130710 20469
rect 130744 20327 131130 20469
rect 131164 20327 131550 20469
rect 131584 20327 131970 20469
rect 132004 20327 132390 20469
rect 132424 20327 132810 20469
rect 132844 20327 133230 20469
rect 133264 20327 133650 20469
rect 133684 20327 134070 20469
rect 134104 20327 134490 20469
rect 134524 20327 134910 20469
rect 134944 20327 134956 20469
rect 126474 20320 134956 20327
rect 126474 20310 126484 20320
rect 122026 20268 122072 20280
rect 122122 20268 122168 20280
rect 122236 20268 122282 20280
rect 122332 20268 122378 20280
rect 122446 20268 122492 20280
rect 122542 20268 122588 20280
rect 122656 20268 122702 20280
rect 122752 20268 122798 20280
rect 122866 20268 122912 20280
rect 122962 20268 123008 20280
rect 123076 20268 123122 20280
rect 123172 20268 123218 20280
rect 123286 20268 123332 20280
rect 123382 20268 123428 20280
rect 123496 20268 123542 20280
rect 123592 20268 123638 20280
rect 123706 20268 123752 20280
rect 123802 20268 123848 20280
rect 123916 20268 123962 20280
rect 124012 20268 124058 20280
rect 124126 20268 124172 20280
rect 124222 20268 124268 20280
rect 124336 20268 124382 20280
rect 124432 20268 124478 20280
rect 124546 20268 124592 20280
rect 124642 20268 124688 20280
rect 124756 20268 124802 20280
rect 124852 20268 124898 20280
rect 124966 20268 125012 20280
rect 125062 20268 125108 20280
rect 125176 20268 125222 20280
rect 125272 20268 125318 20280
rect 125386 20268 125432 20280
rect 125482 20268 125528 20280
rect 125596 20268 125642 20280
rect 125692 20268 125738 20280
rect 121546 19452 121776 19668
rect 121546 19432 121556 19452
rect 120062 19272 120108 19284
rect 120158 19272 120204 19284
rect 120272 19272 120318 19284
rect 120368 19272 120414 19284
rect 120482 19272 120528 19284
rect 120578 19272 120624 19284
rect 120692 19272 120738 19284
rect 120788 19272 120834 19284
rect 120104 19234 120162 19240
rect 120104 19206 120116 19234
rect 119474 19188 120116 19206
rect 119322 19128 120116 19188
rect 119156 19084 119214 19091
rect 119114 19032 119160 19044
rect 119210 19032 119256 19044
rect 119306 19032 119352 19044
rect 119072 18056 119082 19032
rect 119154 18056 119164 19032
rect 119196 18056 119206 19032
rect 119260 18056 119270 19032
rect 119302 18056 119312 19032
rect 119384 18056 119394 19032
rect 119114 18044 119160 18056
rect 119210 18044 119256 18056
rect 119306 18044 119352 18056
rect 119534 18004 119648 19128
rect 120104 19091 120116 19128
rect 120150 19206 120162 19234
rect 120524 19234 120582 19240
rect 120524 19206 120536 19234
rect 120150 19128 120536 19206
rect 120150 19091 120162 19128
rect 120104 19085 120162 19091
rect 120524 19091 120536 19128
rect 120570 19194 120582 19234
rect 121590 19234 121776 19452
rect 121998 19292 122008 20268
rect 122066 19292 122076 20268
rect 122118 19292 122128 20268
rect 122276 19292 122286 20268
rect 122328 19292 122338 20268
rect 122486 19292 122496 20268
rect 122538 19292 122548 20268
rect 122696 19292 122706 20268
rect 122748 19292 122758 20268
rect 122906 19292 122916 20268
rect 122958 19292 122968 20268
rect 123116 19292 123126 20268
rect 123168 19292 123178 20268
rect 123326 19292 123336 20268
rect 123378 19292 123388 20268
rect 123536 19292 123546 20268
rect 123588 19292 123598 20268
rect 123746 19292 123756 20268
rect 123798 19292 123808 20268
rect 123956 19292 123966 20268
rect 124008 19292 124018 20268
rect 124166 19292 124176 20268
rect 124218 19292 124228 20268
rect 124376 19292 124386 20268
rect 124428 19292 124438 20268
rect 124586 19292 124596 20268
rect 124638 19292 124648 20268
rect 124796 19292 124806 20268
rect 124848 19292 124858 20268
rect 125006 19292 125016 20268
rect 125058 19292 125068 20268
rect 125216 19292 125226 20268
rect 125268 19292 125278 20268
rect 125426 19292 125436 20268
rect 125478 19292 125488 20268
rect 125636 19292 125646 20268
rect 125688 19292 125698 20268
rect 125756 19292 125766 20268
rect 122026 19280 122072 19292
rect 122122 19280 122168 19292
rect 122236 19280 122282 19292
rect 122332 19280 122378 19292
rect 122446 19280 122492 19292
rect 122542 19280 122588 19292
rect 122656 19280 122702 19292
rect 122752 19280 122798 19292
rect 122866 19280 122912 19292
rect 122962 19280 123008 19292
rect 123076 19280 123122 19292
rect 123172 19280 123218 19292
rect 123286 19280 123332 19292
rect 123382 19280 123428 19292
rect 123496 19280 123542 19292
rect 123592 19280 123638 19292
rect 123706 19280 123752 19292
rect 123802 19280 123848 19292
rect 123916 19280 123962 19292
rect 124012 19280 124058 19292
rect 124126 19280 124172 19292
rect 124222 19280 124268 19292
rect 124336 19280 124382 19292
rect 124432 19280 124478 19292
rect 124546 19280 124592 19292
rect 124642 19280 124688 19292
rect 124756 19280 124802 19292
rect 124852 19280 124898 19292
rect 124966 19280 125012 19292
rect 125062 19280 125108 19292
rect 125176 19280 125222 19292
rect 125272 19280 125318 19292
rect 125386 19280 125432 19292
rect 125482 19280 125528 19292
rect 125596 19280 125642 19292
rect 125692 19280 125738 19292
rect 125964 19240 126436 20310
rect 126876 20268 126922 20280
rect 126972 20268 127018 20280
rect 127086 20268 127132 20280
rect 127182 20268 127228 20280
rect 127296 20268 127342 20280
rect 127392 20268 127438 20280
rect 127506 20268 127552 20280
rect 127602 20268 127648 20280
rect 127716 20268 127762 20280
rect 127812 20268 127858 20280
rect 127926 20268 127972 20280
rect 128022 20268 128068 20280
rect 128136 20268 128182 20280
rect 128232 20268 128278 20280
rect 128346 20268 128392 20280
rect 128442 20268 128488 20280
rect 128556 20268 128602 20280
rect 128652 20268 128698 20280
rect 128766 20268 128812 20280
rect 128862 20268 128908 20280
rect 128976 20268 129022 20280
rect 129072 20268 129118 20280
rect 129186 20268 129232 20280
rect 129282 20268 129328 20280
rect 129396 20268 129442 20280
rect 129492 20268 129538 20280
rect 129606 20268 129652 20280
rect 129702 20268 129748 20280
rect 129816 20268 129862 20280
rect 129912 20268 129958 20280
rect 130026 20268 130072 20280
rect 130122 20268 130168 20280
rect 130236 20268 130282 20280
rect 130332 20268 130378 20280
rect 130446 20268 130492 20280
rect 130542 20268 130588 20280
rect 130656 20268 130702 20280
rect 130752 20268 130798 20280
rect 130866 20268 130912 20280
rect 130962 20268 131008 20280
rect 131076 20268 131122 20280
rect 131172 20268 131218 20280
rect 131286 20268 131332 20280
rect 131382 20268 131428 20280
rect 131496 20268 131542 20280
rect 131592 20268 131638 20280
rect 131706 20268 131752 20280
rect 131802 20268 131848 20280
rect 131916 20268 131962 20280
rect 132012 20268 132058 20280
rect 132126 20268 132172 20280
rect 132222 20268 132268 20280
rect 132336 20268 132382 20280
rect 132432 20268 132478 20280
rect 132546 20268 132592 20280
rect 132642 20268 132688 20280
rect 132756 20268 132802 20280
rect 132852 20268 132898 20280
rect 132966 20268 133012 20280
rect 133062 20268 133108 20280
rect 133176 20268 133222 20280
rect 133272 20268 133318 20280
rect 133386 20268 133432 20280
rect 133482 20268 133528 20280
rect 133596 20268 133642 20280
rect 133692 20268 133738 20280
rect 133806 20268 133852 20280
rect 133902 20268 133948 20280
rect 134016 20268 134062 20280
rect 134112 20268 134158 20280
rect 134226 20268 134272 20280
rect 134322 20268 134368 20280
rect 134436 20268 134482 20280
rect 134532 20268 134578 20280
rect 134646 20268 134692 20280
rect 134742 20268 134788 20280
rect 134856 20268 134902 20280
rect 134952 20268 134998 20280
rect 135066 20268 135112 20280
rect 135162 20268 135208 20280
rect 126848 19292 126858 20268
rect 126916 19292 126926 20268
rect 126968 19292 126978 20268
rect 127126 19292 127136 20268
rect 127178 19292 127188 20268
rect 127336 19292 127346 20268
rect 127388 19292 127398 20268
rect 127546 19292 127556 20268
rect 127598 19292 127608 20268
rect 127756 19292 127766 20268
rect 127808 19292 127818 20268
rect 127966 19292 127976 20268
rect 128018 19292 128028 20268
rect 128176 19292 128186 20268
rect 128228 19292 128238 20268
rect 128386 19292 128396 20268
rect 128438 19292 128448 20268
rect 128596 19292 128606 20268
rect 128648 19292 128658 20268
rect 128806 19292 128816 20268
rect 128858 19292 128868 20268
rect 129016 19292 129026 20268
rect 129068 19292 129078 20268
rect 129226 19292 129236 20268
rect 129278 19292 129288 20268
rect 129436 19292 129446 20268
rect 129488 19292 129498 20268
rect 129646 19292 129656 20268
rect 129698 19292 129708 20268
rect 129856 19292 129866 20268
rect 129908 19292 129918 20268
rect 130066 19292 130076 20268
rect 130118 19292 130128 20268
rect 130276 19292 130286 20268
rect 130328 19292 130338 20268
rect 130486 19292 130496 20268
rect 130538 19292 130548 20268
rect 130696 19292 130706 20268
rect 130748 19292 130758 20268
rect 130906 19292 130916 20268
rect 130958 19292 130968 20268
rect 131116 19292 131126 20268
rect 131168 19292 131178 20268
rect 131326 19292 131336 20268
rect 131378 19292 131388 20268
rect 131536 19292 131546 20268
rect 131588 19292 131598 20268
rect 131746 19292 131756 20268
rect 131798 19292 131808 20268
rect 131956 19292 131966 20268
rect 132008 19292 132018 20268
rect 132166 19292 132176 20268
rect 132218 19292 132228 20268
rect 132376 19292 132386 20268
rect 132428 19292 132438 20268
rect 132586 19292 132596 20268
rect 132638 19292 132648 20268
rect 132796 19292 132806 20268
rect 132848 19292 132858 20268
rect 133006 19292 133016 20268
rect 133058 19292 133068 20268
rect 133216 19292 133226 20268
rect 133268 19292 133278 20268
rect 133426 19292 133436 20268
rect 133478 19292 133488 20268
rect 133636 19292 133646 20268
rect 133688 19292 133698 20268
rect 133846 19292 133856 20268
rect 133898 19292 133908 20268
rect 134056 19292 134066 20268
rect 134108 19292 134118 20268
rect 134266 19292 134276 20268
rect 134318 19292 134328 20268
rect 134476 19292 134486 20268
rect 134528 19292 134538 20268
rect 134686 19292 134696 20268
rect 134738 19292 134748 20268
rect 134896 19292 134906 20268
rect 134948 19292 134958 20268
rect 135106 19292 135116 20268
rect 135158 19292 135168 20268
rect 135226 19292 135236 20268
rect 126876 19280 126922 19292
rect 126972 19280 127018 19292
rect 127086 19280 127132 19292
rect 127182 19280 127228 19292
rect 127296 19280 127342 19292
rect 127392 19280 127438 19292
rect 127506 19280 127552 19292
rect 127602 19280 127648 19292
rect 127716 19280 127762 19292
rect 127812 19280 127858 19292
rect 127926 19280 127972 19292
rect 128022 19280 128068 19292
rect 128136 19280 128182 19292
rect 128232 19280 128278 19292
rect 128346 19280 128392 19292
rect 128442 19280 128488 19292
rect 128556 19280 128602 19292
rect 128652 19280 128698 19292
rect 128766 19280 128812 19292
rect 128862 19280 128908 19292
rect 128976 19280 129022 19292
rect 129072 19280 129118 19292
rect 129186 19280 129232 19292
rect 129282 19280 129328 19292
rect 129396 19280 129442 19292
rect 129492 19280 129538 19292
rect 129606 19280 129652 19292
rect 129702 19280 129748 19292
rect 129816 19280 129862 19292
rect 129912 19280 129958 19292
rect 130026 19280 130072 19292
rect 130122 19280 130168 19292
rect 130236 19280 130282 19292
rect 130332 19280 130378 19292
rect 130446 19280 130492 19292
rect 130542 19280 130588 19292
rect 130656 19280 130702 19292
rect 130752 19280 130798 19292
rect 130866 19280 130912 19292
rect 130962 19280 131008 19292
rect 131076 19280 131122 19292
rect 131172 19280 131218 19292
rect 131286 19280 131332 19292
rect 131382 19280 131428 19292
rect 131496 19280 131542 19292
rect 131592 19280 131638 19292
rect 131706 19280 131752 19292
rect 131802 19280 131848 19292
rect 131916 19280 131962 19292
rect 132012 19280 132058 19292
rect 132126 19280 132172 19292
rect 132222 19280 132268 19292
rect 132336 19280 132382 19292
rect 132432 19280 132478 19292
rect 132546 19280 132592 19292
rect 132642 19280 132688 19292
rect 132756 19280 132802 19292
rect 132852 19280 132898 19292
rect 132966 19280 133012 19292
rect 133062 19280 133108 19292
rect 133176 19280 133222 19292
rect 133272 19280 133318 19292
rect 133386 19280 133432 19292
rect 133482 19280 133528 19292
rect 133596 19280 133642 19292
rect 133692 19280 133738 19292
rect 133806 19280 133852 19292
rect 133902 19280 133948 19292
rect 134016 19280 134062 19292
rect 134112 19280 134158 19292
rect 134226 19280 134272 19292
rect 134322 19280 134368 19292
rect 134436 19280 134482 19292
rect 134532 19280 134578 19292
rect 134646 19280 134692 19292
rect 134742 19280 134788 19292
rect 134856 19280 134902 19292
rect 134952 19280 134998 19292
rect 135066 19280 135112 19292
rect 135162 19280 135208 19292
rect 122278 19234 122336 19239
rect 122698 19234 122756 19239
rect 123118 19234 123176 19239
rect 123538 19234 123596 19239
rect 123958 19234 124016 19239
rect 124378 19234 124436 19239
rect 124798 19234 124856 19239
rect 125218 19234 125276 19239
rect 125638 19234 125696 19239
rect 121590 19233 125696 19234
rect 120570 19132 120576 19194
rect 120570 19125 121472 19132
rect 120570 19091 120956 19125
rect 120990 19124 121376 19125
rect 121410 19124 121472 19125
rect 120524 19090 120956 19091
rect 121040 19090 121376 19124
rect 121460 19090 121472 19124
rect 120524 19085 121472 19090
rect 120574 19082 121472 19085
rect 121590 19091 122290 19233
rect 122324 19091 122710 19233
rect 122744 19091 123130 19233
rect 123164 19091 123550 19233
rect 123584 19091 123970 19233
rect 124004 19091 124390 19233
rect 124424 19091 124810 19233
rect 124844 19091 125230 19233
rect 125264 19091 125650 19233
rect 125684 19091 125696 19233
rect 121590 19084 125696 19091
rect 125964 19233 135166 19240
rect 125964 19091 127140 19233
rect 127174 19091 127560 19233
rect 127594 19091 127980 19233
rect 128014 19091 128400 19233
rect 128434 19091 128820 19233
rect 128854 19091 129240 19233
rect 129274 19091 129660 19233
rect 129694 19091 130080 19233
rect 130114 19091 130500 19233
rect 130534 19091 130920 19233
rect 130954 19091 131340 19233
rect 131374 19091 131760 19233
rect 131794 19091 132180 19233
rect 132214 19091 132600 19233
rect 132634 19091 133020 19233
rect 133054 19091 133440 19233
rect 133474 19091 133860 19233
rect 133894 19091 134280 19233
rect 134314 19091 134700 19233
rect 134734 19091 135120 19233
rect 135154 19091 135166 19233
rect 125964 19084 135166 19091
rect 119852 19032 119898 19044
rect 119948 19032 119994 19044
rect 120062 19032 120108 19044
rect 120158 19032 120204 19044
rect 120272 19032 120318 19044
rect 120368 19032 120414 19044
rect 120482 19032 120528 19044
rect 120578 19032 120624 19044
rect 120692 19032 120738 19044
rect 120788 19032 120834 19044
rect 120902 19032 120948 19044
rect 120998 19032 121044 19044
rect 121112 19032 121158 19044
rect 121208 19032 121254 19044
rect 121322 19032 121368 19044
rect 121418 19032 121464 19044
rect 119824 18056 119834 19032
rect 119892 18056 119902 19032
rect 119944 18056 119954 19032
rect 120102 18056 120112 19032
rect 120154 18056 120164 19032
rect 120312 18056 120322 19032
rect 120364 18056 120374 19032
rect 120522 18056 120532 19032
rect 120574 18056 120584 19032
rect 120732 18056 120742 19032
rect 120784 18056 120794 19032
rect 120942 18056 120952 19032
rect 120994 18056 121004 19032
rect 121152 18056 121162 19032
rect 121204 18056 121214 19032
rect 121362 18056 121372 19032
rect 121414 18056 121424 19032
rect 121482 18056 121492 19032
rect 119852 18044 119898 18056
rect 119948 18044 119994 18056
rect 120062 18044 120108 18056
rect 120158 18044 120204 18056
rect 120272 18044 120318 18056
rect 120368 18044 120414 18056
rect 120482 18044 120528 18056
rect 120578 18044 120624 18056
rect 120692 18044 120738 18056
rect 120788 18044 120834 18056
rect 120902 18044 120948 18056
rect 120998 18044 121044 18056
rect 121112 18044 121158 18056
rect 121208 18044 121254 18056
rect 121322 18044 121368 18056
rect 121418 18044 121464 18056
rect 121590 18004 121776 19084
rect 122026 19032 122072 19044
rect 122122 19032 122168 19044
rect 122236 19032 122282 19044
rect 122332 19032 122378 19044
rect 122446 19032 122492 19044
rect 122542 19032 122588 19044
rect 122656 19032 122702 19044
rect 122752 19032 122798 19044
rect 122866 19032 122912 19044
rect 122962 19032 123008 19044
rect 123076 19032 123122 19044
rect 123172 19032 123218 19044
rect 123286 19032 123332 19044
rect 123382 19032 123428 19044
rect 123496 19032 123542 19044
rect 123592 19032 123638 19044
rect 123706 19032 123752 19044
rect 123802 19032 123848 19044
rect 123916 19032 123962 19044
rect 124012 19032 124058 19044
rect 124126 19032 124172 19044
rect 124222 19032 124268 19044
rect 124336 19032 124382 19044
rect 124432 19032 124478 19044
rect 124546 19032 124592 19044
rect 124642 19032 124688 19044
rect 124756 19032 124802 19044
rect 124852 19032 124898 19044
rect 124966 19032 125012 19044
rect 125062 19032 125108 19044
rect 125176 19032 125222 19044
rect 125272 19032 125318 19044
rect 125386 19032 125432 19044
rect 125482 19032 125528 19044
rect 125596 19032 125642 19044
rect 125692 19032 125738 19044
rect 121998 18056 122008 19032
rect 122066 18056 122076 19032
rect 122118 18056 122128 19032
rect 122276 18056 122286 19032
rect 122328 18056 122338 19032
rect 122486 18056 122496 19032
rect 122538 18056 122548 19032
rect 122696 18056 122706 19032
rect 122748 18056 122758 19032
rect 122906 18056 122916 19032
rect 122958 18056 122968 19032
rect 123116 18056 123126 19032
rect 123168 18056 123178 19032
rect 123326 18056 123336 19032
rect 123378 18056 123388 19032
rect 123536 18056 123546 19032
rect 123588 18056 123598 19032
rect 123746 18056 123756 19032
rect 123798 18056 123808 19032
rect 123956 18056 123966 19032
rect 124008 18056 124018 19032
rect 124166 18056 124176 19032
rect 124218 18056 124228 19032
rect 124376 18056 124386 19032
rect 124428 18056 124438 19032
rect 124586 18056 124596 19032
rect 124638 18056 124648 19032
rect 124796 18056 124806 19032
rect 124848 18056 124858 19032
rect 125006 18056 125016 19032
rect 125058 18056 125068 19032
rect 125216 18056 125226 19032
rect 125268 18056 125278 19032
rect 125426 18056 125436 19032
rect 125478 18056 125488 19032
rect 125636 18056 125646 19032
rect 125688 18056 125698 19032
rect 125756 18056 125766 19032
rect 122026 18044 122072 18056
rect 122122 18044 122168 18056
rect 122236 18044 122282 18056
rect 122332 18044 122378 18056
rect 122446 18044 122492 18056
rect 122542 18044 122588 18056
rect 122656 18044 122702 18056
rect 122752 18044 122798 18056
rect 122866 18044 122912 18056
rect 122962 18044 123008 18056
rect 123076 18044 123122 18056
rect 123172 18044 123218 18056
rect 123286 18044 123332 18056
rect 123382 18044 123428 18056
rect 123496 18044 123542 18056
rect 123592 18044 123638 18056
rect 123706 18044 123752 18056
rect 123802 18044 123848 18056
rect 123916 18044 123962 18056
rect 124012 18044 124058 18056
rect 124126 18044 124172 18056
rect 124222 18044 124268 18056
rect 124336 18044 124382 18056
rect 124432 18044 124478 18056
rect 124546 18044 124592 18056
rect 124642 18044 124688 18056
rect 124756 18044 124802 18056
rect 124852 18044 124898 18056
rect 124966 18044 125012 18056
rect 125062 18044 125108 18056
rect 125176 18044 125222 18056
rect 125272 18044 125318 18056
rect 125386 18044 125432 18056
rect 125482 18044 125528 18056
rect 125596 18044 125642 18056
rect 125692 18044 125738 18056
rect 125964 18004 126436 19084
rect 126876 19032 126922 19044
rect 126972 19032 127018 19044
rect 127086 19032 127132 19044
rect 127182 19032 127228 19044
rect 127296 19032 127342 19044
rect 127392 19032 127438 19044
rect 127506 19032 127552 19044
rect 127602 19032 127648 19044
rect 127716 19032 127762 19044
rect 127812 19032 127858 19044
rect 127926 19032 127972 19044
rect 128022 19032 128068 19044
rect 128136 19032 128182 19044
rect 128232 19032 128278 19044
rect 128346 19032 128392 19044
rect 128442 19032 128488 19044
rect 128556 19032 128602 19044
rect 128652 19032 128698 19044
rect 128766 19032 128812 19044
rect 128862 19032 128908 19044
rect 128976 19032 129022 19044
rect 129072 19032 129118 19044
rect 129186 19032 129232 19044
rect 129282 19032 129328 19044
rect 129396 19032 129442 19044
rect 129492 19032 129538 19044
rect 129606 19032 129652 19044
rect 129702 19032 129748 19044
rect 129816 19032 129862 19044
rect 129912 19032 129958 19044
rect 130026 19032 130072 19044
rect 130122 19032 130168 19044
rect 130236 19032 130282 19044
rect 130332 19032 130378 19044
rect 130446 19032 130492 19044
rect 130542 19032 130588 19044
rect 130656 19032 130702 19044
rect 130752 19032 130798 19044
rect 130866 19032 130912 19044
rect 130962 19032 131008 19044
rect 131076 19032 131122 19044
rect 131172 19032 131218 19044
rect 131286 19032 131332 19044
rect 131382 19032 131428 19044
rect 131496 19032 131542 19044
rect 131592 19032 131638 19044
rect 131706 19032 131752 19044
rect 131802 19032 131848 19044
rect 131916 19032 131962 19044
rect 132012 19032 132058 19044
rect 132126 19032 132172 19044
rect 132222 19032 132268 19044
rect 132336 19032 132382 19044
rect 132432 19032 132478 19044
rect 132546 19032 132592 19044
rect 132642 19032 132688 19044
rect 132756 19032 132802 19044
rect 132852 19032 132898 19044
rect 132966 19032 133012 19044
rect 133062 19032 133108 19044
rect 133176 19032 133222 19044
rect 133272 19032 133318 19044
rect 133386 19032 133432 19044
rect 133482 19032 133528 19044
rect 133596 19032 133642 19044
rect 133692 19032 133738 19044
rect 133806 19032 133852 19044
rect 133902 19032 133948 19044
rect 134016 19032 134062 19044
rect 134112 19032 134158 19044
rect 134226 19032 134272 19044
rect 134322 19032 134368 19044
rect 134436 19032 134482 19044
rect 134532 19032 134578 19044
rect 134646 19032 134692 19044
rect 134742 19032 134788 19044
rect 134856 19032 134902 19044
rect 134952 19032 134998 19044
rect 135066 19032 135112 19044
rect 135162 19032 135208 19044
rect 126848 18056 126858 19032
rect 126916 18056 126926 19032
rect 126968 18056 126978 19032
rect 127126 18056 127136 19032
rect 127178 18056 127188 19032
rect 127336 18056 127346 19032
rect 127388 18056 127398 19032
rect 127546 18056 127556 19032
rect 127598 18056 127608 19032
rect 127756 18056 127766 19032
rect 127808 18056 127818 19032
rect 127966 18056 127976 19032
rect 128018 18056 128028 19032
rect 128176 18056 128186 19032
rect 128228 18056 128238 19032
rect 128386 18056 128396 19032
rect 128438 18056 128448 19032
rect 128596 18056 128606 19032
rect 128648 18056 128658 19032
rect 128806 18056 128816 19032
rect 128858 18056 128868 19032
rect 129016 18056 129026 19032
rect 129068 18056 129078 19032
rect 129226 18056 129236 19032
rect 129278 18056 129288 19032
rect 129436 18056 129446 19032
rect 129488 18056 129498 19032
rect 129646 18056 129656 19032
rect 129698 18056 129708 19032
rect 129856 18056 129866 19032
rect 129908 18056 129918 19032
rect 130066 18056 130076 19032
rect 130118 18056 130128 19032
rect 130276 18056 130286 19032
rect 130328 18056 130338 19032
rect 130486 18056 130496 19032
rect 130538 18056 130548 19032
rect 130696 18056 130706 19032
rect 130748 18056 130758 19032
rect 130906 18056 130916 19032
rect 130958 18056 130968 19032
rect 131116 18056 131126 19032
rect 131168 18056 131178 19032
rect 131326 18056 131336 19032
rect 131378 18056 131388 19032
rect 131536 18056 131546 19032
rect 131588 18056 131598 19032
rect 131746 18056 131756 19032
rect 131798 18056 131808 19032
rect 131956 18056 131966 19032
rect 132008 18056 132018 19032
rect 132166 18056 132176 19032
rect 132218 18056 132228 19032
rect 132376 18056 132386 19032
rect 132428 18056 132438 19032
rect 132586 18056 132596 19032
rect 132638 18056 132648 19032
rect 132796 18056 132806 19032
rect 132848 18056 132858 19032
rect 133006 18056 133016 19032
rect 133058 18056 133068 19032
rect 133216 18056 133226 19032
rect 133268 18056 133278 19032
rect 133426 18056 133436 19032
rect 133478 18056 133488 19032
rect 133636 18056 133646 19032
rect 133688 18056 133698 19032
rect 133846 18056 133856 19032
rect 133898 18056 133908 19032
rect 134056 18056 134066 19032
rect 134108 18056 134118 19032
rect 134266 18056 134276 19032
rect 134318 18056 134328 19032
rect 134476 18056 134486 19032
rect 134528 18056 134538 19032
rect 134686 18056 134696 19032
rect 134738 18056 134748 19032
rect 134896 18056 134906 19032
rect 134948 18056 134958 19032
rect 135106 18056 135116 19032
rect 135158 18056 135168 19032
rect 135226 18056 135236 19032
rect 126876 18044 126922 18056
rect 126972 18044 127018 18056
rect 127086 18044 127132 18056
rect 127182 18044 127228 18056
rect 127296 18044 127342 18056
rect 127392 18044 127438 18056
rect 127506 18044 127552 18056
rect 127602 18044 127648 18056
rect 127716 18044 127762 18056
rect 127812 18044 127858 18056
rect 127926 18044 127972 18056
rect 128022 18044 128068 18056
rect 128136 18044 128182 18056
rect 128232 18044 128278 18056
rect 128346 18044 128392 18056
rect 128442 18044 128488 18056
rect 128556 18044 128602 18056
rect 128652 18044 128698 18056
rect 128766 18044 128812 18056
rect 128862 18044 128908 18056
rect 128976 18044 129022 18056
rect 129072 18044 129118 18056
rect 129186 18044 129232 18056
rect 129282 18044 129328 18056
rect 129396 18044 129442 18056
rect 129492 18044 129538 18056
rect 129606 18044 129652 18056
rect 129702 18044 129748 18056
rect 129816 18044 129862 18056
rect 129912 18044 129958 18056
rect 130026 18044 130072 18056
rect 130122 18044 130168 18056
rect 130236 18044 130282 18056
rect 130332 18044 130378 18056
rect 130446 18044 130492 18056
rect 130542 18044 130588 18056
rect 130656 18044 130702 18056
rect 130752 18044 130798 18056
rect 130866 18044 130912 18056
rect 130962 18044 131008 18056
rect 131076 18044 131122 18056
rect 131172 18044 131218 18056
rect 131286 18044 131332 18056
rect 131382 18044 131428 18056
rect 131496 18044 131542 18056
rect 131592 18044 131638 18056
rect 131706 18044 131752 18056
rect 131802 18044 131848 18056
rect 131916 18044 131962 18056
rect 132012 18044 132058 18056
rect 132126 18044 132172 18056
rect 132222 18044 132268 18056
rect 132336 18044 132382 18056
rect 132432 18044 132478 18056
rect 132546 18044 132592 18056
rect 132642 18044 132688 18056
rect 132756 18044 132802 18056
rect 132852 18044 132898 18056
rect 132966 18044 133012 18056
rect 133062 18044 133108 18056
rect 133176 18044 133222 18056
rect 133272 18044 133318 18056
rect 133386 18044 133432 18056
rect 133482 18044 133528 18056
rect 133596 18044 133642 18056
rect 133692 18044 133738 18056
rect 133806 18044 133852 18056
rect 133902 18044 133948 18056
rect 134016 18044 134062 18056
rect 134112 18044 134158 18056
rect 134226 18044 134272 18056
rect 134322 18044 134368 18056
rect 134436 18044 134482 18056
rect 134532 18044 134578 18056
rect 134646 18044 134692 18056
rect 134742 18044 134788 18056
rect 134856 18044 134902 18056
rect 134952 18044 134998 18056
rect 135066 18044 135112 18056
rect 135162 18044 135208 18056
rect 118766 17998 119360 18004
rect 118766 17964 119264 17998
rect 119348 17964 119360 17998
rect 118766 17958 119360 17964
rect 119534 18002 119688 18004
rect 119894 18002 119952 18003
rect 120314 18002 120372 18003
rect 120734 18002 120792 18003
rect 121154 18002 121212 18003
rect 119534 17997 121262 18002
rect 119534 17962 119906 17997
rect 119940 17996 120326 17997
rect 120360 17996 120746 17997
rect 120780 17996 121166 17997
rect 121200 17996 121262 17997
rect 119990 17962 120326 17996
rect 120410 17962 120746 17996
rect 120830 17962 121166 17996
rect 121250 17962 121262 17996
rect 118766 17956 119306 17958
rect 119534 17956 121262 17962
rect 121590 17997 125536 18004
rect 121590 17962 122080 17997
rect 122114 17996 122500 17997
rect 122534 17996 122920 17997
rect 122954 17996 123340 17997
rect 123374 17996 123760 17997
rect 123794 17996 124180 17997
rect 124214 17996 124600 17997
rect 124634 17996 125020 17997
rect 125054 17996 125440 17997
rect 125474 17996 125536 17997
rect 122164 17962 122500 17996
rect 122584 17962 122920 17996
rect 123004 17962 123340 17996
rect 123424 17962 123760 17996
rect 123844 17962 124180 17996
rect 124264 17962 124600 17996
rect 124684 17962 125020 17996
rect 125104 17962 125440 17996
rect 125524 17962 125536 17996
rect 116724 17152 116734 17414
rect 117062 17152 117072 17414
rect 116842 17054 116954 17152
rect 118766 17054 118860 17956
rect 119890 17954 119948 17956
rect 120310 17954 120368 17956
rect 120730 17954 120788 17956
rect 121150 17954 121208 17956
rect 121590 17954 125536 17962
rect 125964 17997 135006 18004
rect 125964 17962 126930 17997
rect 126964 17996 127350 17997
rect 127384 17996 127770 17997
rect 127804 17996 128190 17997
rect 128224 17996 128610 17997
rect 128644 17996 129030 17997
rect 129064 17996 129450 17997
rect 129484 17996 129870 17997
rect 129904 17996 130290 17997
rect 130324 17996 130710 17997
rect 130744 17996 131130 17997
rect 131164 17996 131550 17997
rect 131584 17996 131970 17997
rect 132004 17996 132390 17997
rect 132424 17996 132810 17997
rect 132844 17996 133230 17997
rect 133264 17996 133650 17997
rect 133684 17996 134070 17997
rect 134104 17996 134490 17997
rect 134524 17996 134910 17997
rect 134944 17996 135006 17997
rect 127014 17962 127350 17996
rect 127434 17962 127770 17996
rect 127854 17962 128190 17996
rect 128274 17962 128610 17996
rect 128694 17962 129030 17996
rect 129114 17962 129450 17996
rect 129534 17962 129870 17996
rect 129954 17962 130290 17996
rect 130374 17962 130710 17996
rect 130794 17962 131130 17996
rect 131214 17962 131550 17996
rect 131634 17962 131970 17996
rect 132054 17962 132390 17996
rect 132474 17962 132810 17996
rect 132894 17962 133230 17996
rect 133314 17962 133650 17996
rect 133734 17962 134070 17996
rect 134154 17962 134490 17996
rect 134574 17962 134910 17996
rect 134994 17962 135006 17996
rect 125964 17954 135006 17962
rect 119516 17770 119672 17782
rect 119512 17622 119522 17770
rect 119666 17622 119676 17770
rect 119516 17610 119672 17622
rect 116356 17026 116366 17044
rect 116212 16962 116366 17026
rect 116212 16842 116272 16962
rect 116356 16958 116366 16962
rect 116450 16958 116460 17044
rect 116842 16976 118860 17054
rect 116376 16906 116422 16958
rect 116184 16830 116290 16842
rect 116184 16616 116190 16830
rect 116284 16616 116290 16830
rect 116184 16604 116290 16616
rect 116376 16530 116382 16906
rect 116416 16530 116422 16906
rect 116376 16518 116422 16530
rect 116464 16906 116516 16918
rect 116464 16530 116476 16906
rect 116510 16530 116516 16906
rect 116464 16518 116516 16530
rect 116558 16906 116604 16918
rect 116558 16530 116564 16906
rect 116598 16558 116604 16906
rect 116598 16530 116662 16558
rect 116558 16518 116662 16530
rect 115580 16470 116598 16476
rect 115580 16424 116512 16470
rect 116586 16424 116598 16470
rect 115580 16418 116598 16424
rect 115580 14980 115652 16418
rect 116338 16332 116350 16390
rect 116424 16332 116436 16390
rect 116626 16378 116662 16518
rect 116842 16378 116954 16976
rect 116464 16338 116954 16378
rect 116376 16286 116422 16298
rect 116202 16204 116290 16216
rect 116202 15998 116208 16204
rect 116284 15998 116290 16204
rect 116202 15986 116290 15998
rect 116230 15806 116270 15986
rect 116376 15910 116382 16286
rect 116416 15910 116422 16286
rect 116376 15806 116422 15910
rect 116464 16286 116516 16338
rect 116464 15910 116476 16286
rect 116510 15910 116516 16286
rect 116464 15898 116516 15910
rect 116558 16286 116604 16298
rect 116558 15910 116564 16286
rect 116598 15910 116604 16286
rect 120914 16218 120924 16466
rect 121168 16218 121178 16466
rect 116558 15806 116604 15910
rect 116230 15804 116422 15806
rect 116542 15804 116604 15806
rect 116230 15754 116370 15804
rect 116360 15730 116370 15754
rect 116440 15730 116450 15804
rect 116542 15730 116552 15804
rect 116622 15730 116632 15804
rect 116360 15636 116370 15660
rect 115834 15594 115844 15620
rect 115744 15556 115844 15594
rect 115744 15438 115806 15556
rect 115834 15554 115844 15556
rect 115908 15554 115918 15620
rect 116230 15586 116370 15636
rect 116440 15586 116450 15660
rect 116542 15586 116552 15660
rect 116622 15586 116632 15660
rect 116230 15584 116422 15586
rect 116542 15584 116604 15586
rect 115744 15322 115750 15438
rect 115790 15322 115806 15438
rect 115744 15310 115806 15322
rect 115850 15478 115896 15554
rect 115850 15102 115856 15478
rect 115890 15102 115896 15478
rect 115850 15090 115896 15102
rect 115938 15478 115984 15490
rect 115938 15102 115944 15478
rect 115978 15118 115984 15478
rect 116230 15404 116270 15584
rect 116376 15480 116422 15584
rect 116202 15392 116290 15404
rect 116202 15186 116208 15392
rect 116284 15186 116290 15392
rect 116202 15174 116290 15186
rect 115978 15102 116020 15118
rect 115938 15090 116020 15102
rect 116376 15104 116382 15480
rect 116416 15104 116422 15480
rect 116376 15092 116422 15104
rect 116464 15480 116516 15492
rect 116464 15104 116476 15480
rect 116510 15104 116516 15480
rect 115990 15058 116020 15090
rect 115894 15049 115940 15056
rect 115990 15052 116436 15058
rect 115888 15044 115946 15049
rect 115888 14980 115900 15044
rect 115580 14934 115900 14980
rect 115888 14872 115900 14934
rect 115934 15003 115946 15044
rect 115990 15006 116350 15052
rect 116424 15006 116436 15052
rect 116464 15052 116516 15104
rect 116558 15480 116604 15584
rect 116558 15104 116564 15480
rect 116598 15104 116604 15480
rect 116558 15092 116604 15104
rect 116464 15012 116662 15052
rect 115934 14912 115940 15003
rect 115990 15000 116436 15006
rect 115934 14872 115946 14912
rect 115888 14866 115946 14872
rect 115990 14834 116020 15000
rect 116626 14982 116662 15012
rect 116500 14918 116512 14972
rect 116574 14966 116598 14972
rect 116586 14920 116598 14966
rect 116574 14918 116598 14920
rect 116500 14914 116598 14918
rect 116626 14942 116954 14982
rect 116626 14872 116662 14942
rect 115850 14822 115896 14834
rect 115720 14810 115796 14822
rect 115720 14668 115726 14810
rect 115790 14668 115796 14810
rect 115720 14656 115796 14668
rect 115744 14600 115788 14656
rect 115850 14646 115856 14822
rect 115890 14646 115896 14822
rect 115850 14600 115896 14646
rect 115938 14822 116020 14834
rect 115938 14646 115944 14822
rect 115978 14794 116020 14822
rect 116376 14860 116422 14872
rect 115978 14646 115984 14794
rect 115938 14634 115984 14646
rect 116184 14774 116290 14786
rect 115744 14586 115896 14600
rect 115744 14542 115842 14586
rect 115832 14522 115842 14542
rect 115906 14522 115916 14586
rect 116184 14560 116190 14774
rect 116284 14560 116290 14774
rect 116184 14548 116290 14560
rect 116212 14428 116272 14548
rect 116376 14484 116382 14860
rect 116416 14484 116422 14860
rect 116376 14432 116422 14484
rect 116464 14860 116516 14872
rect 116464 14484 116476 14860
rect 116510 14484 116516 14860
rect 116464 14472 116516 14484
rect 116558 14860 116662 14872
rect 116558 14484 116564 14860
rect 116598 14832 116662 14860
rect 116598 14484 116604 14832
rect 116558 14472 116604 14484
rect 116356 14428 116366 14432
rect 116212 14364 116366 14428
rect 116356 14346 116366 14364
rect 116450 14346 116460 14432
rect 116842 14414 116954 14942
rect 120954 14464 121138 16218
rect 121592 15154 121776 17954
rect 121892 17902 122016 17908
rect 121892 17802 121904 17902
rect 122004 17802 122016 17902
rect 121892 17796 122016 17802
rect 122312 17902 122436 17908
rect 122312 17802 122324 17902
rect 122424 17802 122436 17902
rect 122312 17796 122436 17802
rect 122732 17902 122856 17908
rect 122732 17802 122744 17902
rect 122844 17802 122856 17902
rect 122732 17796 122856 17802
rect 123152 17902 123276 17908
rect 123152 17802 123164 17902
rect 123264 17802 123276 17902
rect 123152 17796 123276 17802
rect 123572 17902 123696 17908
rect 123572 17802 123584 17902
rect 123684 17802 123696 17902
rect 123572 17796 123696 17802
rect 123992 17902 124116 17908
rect 123992 17802 124004 17902
rect 124104 17802 124116 17902
rect 123992 17796 124116 17802
rect 124412 17902 124536 17908
rect 124412 17802 124424 17902
rect 124524 17802 124536 17902
rect 124412 17796 124536 17802
rect 124832 17902 124956 17908
rect 124832 17802 124844 17902
rect 124944 17802 124956 17902
rect 124832 17796 124956 17802
rect 125252 17902 125376 17908
rect 125252 17802 125264 17902
rect 125364 17802 125376 17902
rect 125252 17796 125376 17802
rect 125672 17902 125796 17908
rect 125672 17802 125684 17902
rect 125784 17802 125796 17902
rect 125672 17796 125796 17802
rect 126734 17886 126858 17892
rect 126734 17786 126746 17886
rect 126846 17786 126858 17886
rect 126734 17780 126858 17786
rect 127154 17886 127278 17892
rect 127154 17786 127166 17886
rect 127266 17786 127278 17886
rect 127154 17780 127278 17786
rect 127574 17886 127698 17892
rect 127574 17786 127586 17886
rect 127686 17786 127698 17886
rect 127574 17780 127698 17786
rect 127994 17886 128118 17892
rect 127994 17786 128006 17886
rect 128106 17786 128118 17886
rect 127994 17780 128118 17786
rect 128414 17886 128538 17892
rect 128414 17786 128426 17886
rect 128526 17786 128538 17886
rect 128414 17780 128538 17786
rect 128834 17886 128958 17892
rect 128834 17786 128846 17886
rect 128946 17786 128958 17886
rect 128834 17780 128958 17786
rect 129254 17886 129378 17892
rect 129254 17786 129266 17886
rect 129366 17786 129378 17886
rect 129254 17780 129378 17786
rect 129674 17886 129798 17892
rect 129674 17786 129686 17886
rect 129786 17786 129798 17886
rect 129674 17780 129798 17786
rect 130094 17886 130218 17892
rect 130094 17786 130106 17886
rect 130206 17786 130218 17886
rect 130094 17780 130218 17786
rect 130514 17886 130638 17892
rect 130514 17786 130526 17886
rect 130626 17786 130638 17886
rect 130514 17780 130638 17786
rect 130934 17886 131058 17892
rect 130934 17786 130946 17886
rect 131046 17786 131058 17886
rect 130934 17780 131058 17786
rect 131354 17886 131478 17892
rect 131354 17786 131366 17886
rect 131466 17786 131478 17886
rect 131354 17780 131478 17786
rect 131774 17886 131898 17892
rect 131774 17786 131786 17886
rect 131886 17786 131898 17886
rect 131774 17780 131898 17786
rect 132194 17886 132318 17892
rect 132194 17786 132206 17886
rect 132306 17786 132318 17886
rect 132194 17780 132318 17786
rect 132614 17886 132738 17892
rect 132614 17786 132626 17886
rect 132726 17786 132738 17886
rect 132614 17780 132738 17786
rect 133034 17886 133158 17892
rect 133034 17786 133046 17886
rect 133146 17786 133158 17886
rect 133034 17780 133158 17786
rect 133454 17886 133578 17892
rect 133454 17786 133466 17886
rect 133566 17786 133578 17886
rect 133454 17780 133578 17786
rect 133874 17886 133998 17892
rect 133874 17786 133886 17886
rect 133986 17786 133998 17886
rect 133874 17780 133998 17786
rect 134294 17886 134418 17892
rect 134294 17786 134306 17886
rect 134406 17786 134418 17886
rect 134294 17780 134418 17786
rect 134714 17886 134838 17892
rect 134714 17786 134726 17886
rect 134826 17786 134838 17886
rect 134714 17780 134838 17786
rect 135134 17886 135258 17892
rect 135134 17786 135146 17886
rect 135246 17786 135258 17886
rect 135134 17780 135258 17786
rect 121548 14906 121558 15154
rect 121802 14906 121812 15154
rect 116842 14336 118860 14414
rect 116842 14238 116954 14336
rect 116724 13976 116734 14238
rect 117062 13976 117072 14238
rect 118766 13434 118860 14336
rect 120954 14296 121776 14464
rect 119516 13768 119672 13780
rect 119512 13620 119522 13768
rect 119666 13620 119676 13768
rect 119516 13608 119672 13620
rect 121590 13436 121776 14296
rect 121892 13588 122016 13594
rect 121892 13488 121904 13588
rect 122004 13488 122016 13588
rect 121892 13482 122016 13488
rect 122312 13588 122436 13594
rect 122312 13488 122324 13588
rect 122424 13488 122436 13588
rect 122312 13482 122436 13488
rect 122732 13588 122856 13594
rect 122732 13488 122744 13588
rect 122844 13488 122856 13588
rect 122732 13482 122856 13488
rect 123152 13588 123276 13594
rect 123152 13488 123164 13588
rect 123264 13488 123276 13588
rect 123152 13482 123276 13488
rect 123572 13588 123696 13594
rect 123572 13488 123584 13588
rect 123684 13488 123696 13588
rect 123572 13482 123696 13488
rect 123992 13588 124116 13594
rect 123992 13488 124004 13588
rect 124104 13488 124116 13588
rect 123992 13482 124116 13488
rect 124412 13588 124536 13594
rect 124412 13488 124424 13588
rect 124524 13488 124536 13588
rect 124412 13482 124536 13488
rect 124832 13588 124956 13594
rect 124832 13488 124844 13588
rect 124944 13488 124956 13588
rect 124832 13482 124956 13488
rect 125252 13588 125376 13594
rect 125252 13488 125264 13588
rect 125364 13488 125376 13588
rect 125252 13482 125376 13488
rect 125672 13588 125796 13594
rect 125672 13488 125684 13588
rect 125784 13488 125796 13588
rect 125672 13482 125796 13488
rect 119890 13434 119948 13436
rect 120310 13434 120368 13436
rect 120730 13434 120788 13436
rect 121150 13434 121208 13436
rect 118766 13432 119306 13434
rect 118766 13426 119360 13432
rect 118766 13392 119264 13426
rect 119348 13392 119360 13426
rect 118766 13386 119360 13392
rect 119534 13428 121262 13434
rect 119534 13393 119906 13428
rect 119990 13394 120326 13428
rect 120410 13394 120746 13428
rect 120830 13394 121166 13428
rect 121250 13394 121262 13428
rect 119940 13393 120326 13394
rect 120360 13393 120746 13394
rect 120780 13393 121166 13394
rect 121200 13393 121262 13394
rect 119534 13388 121262 13393
rect 121590 13428 125536 13436
rect 121590 13393 122080 13428
rect 122164 13394 122500 13428
rect 122584 13394 122920 13428
rect 123004 13394 123340 13428
rect 123424 13394 123760 13428
rect 123844 13394 124180 13428
rect 124264 13394 124600 13428
rect 124684 13394 125020 13428
rect 125104 13394 125440 13428
rect 125524 13394 125536 13428
rect 122114 13393 122500 13394
rect 122534 13393 122920 13394
rect 122954 13393 123340 13394
rect 123374 13393 123760 13394
rect 123794 13393 124180 13394
rect 124214 13393 124600 13394
rect 124634 13393 125020 13394
rect 125054 13393 125440 13394
rect 125474 13393 125536 13394
rect 119534 13386 119688 13388
rect 119894 13387 119952 13388
rect 120314 13387 120372 13388
rect 120734 13387 120792 13388
rect 121154 13387 121212 13388
rect 121590 13386 125536 13393
rect 118766 12256 118860 13386
rect 119114 13334 119160 13346
rect 119210 13334 119256 13346
rect 119306 13334 119352 13346
rect 119072 12358 119082 13334
rect 119154 12358 119164 13334
rect 119196 12358 119206 13334
rect 119260 12358 119270 13334
rect 119302 12358 119312 13334
rect 119384 12358 119394 13334
rect 119114 12346 119160 12358
rect 119210 12346 119256 12358
rect 119306 12346 119352 12358
rect 119156 12299 119214 12306
rect 119156 12256 119168 12299
rect 118766 12208 119168 12256
rect 119156 12156 119168 12208
rect 119202 12156 119214 12299
rect 119534 12262 119648 13386
rect 119852 13334 119898 13346
rect 119948 13334 119994 13346
rect 120062 13334 120108 13346
rect 120158 13334 120204 13346
rect 120272 13334 120318 13346
rect 120368 13334 120414 13346
rect 120482 13334 120528 13346
rect 120578 13334 120624 13346
rect 120692 13334 120738 13346
rect 120788 13334 120834 13346
rect 120902 13334 120948 13346
rect 120998 13334 121044 13346
rect 121112 13334 121158 13346
rect 121208 13334 121254 13346
rect 121322 13334 121368 13346
rect 121418 13334 121464 13346
rect 119824 12358 119834 13334
rect 119892 12358 119902 13334
rect 119944 12358 119954 13334
rect 120102 12358 120112 13334
rect 120154 12358 120164 13334
rect 120312 12358 120322 13334
rect 120364 12358 120374 13334
rect 120522 12358 120532 13334
rect 120574 12358 120584 13334
rect 120732 12358 120742 13334
rect 120784 12358 120794 13334
rect 120942 12358 120952 13334
rect 120994 12358 121004 13334
rect 121152 12358 121162 13334
rect 121204 12358 121214 13334
rect 121362 12358 121372 13334
rect 121414 12358 121424 13334
rect 121482 12358 121492 13334
rect 119852 12346 119898 12358
rect 119948 12346 119994 12358
rect 120062 12346 120108 12358
rect 120158 12346 120204 12358
rect 120272 12346 120318 12358
rect 120368 12346 120414 12358
rect 120482 12346 120528 12358
rect 120578 12346 120624 12358
rect 120692 12346 120738 12358
rect 120788 12346 120834 12358
rect 120902 12346 120948 12358
rect 120998 12346 121044 12358
rect 121112 12346 121158 12358
rect 121208 12346 121254 12358
rect 121322 12346 121368 12358
rect 121418 12346 121464 12358
rect 120574 12305 121472 12308
rect 120104 12299 120162 12305
rect 120104 12262 120116 12299
rect 119156 12150 119214 12156
rect 119322 12202 120116 12262
rect 119118 12106 119164 12118
rect 119206 12106 119252 12118
rect 119094 11130 119104 12106
rect 119158 11130 119168 12106
rect 119202 11130 119212 12106
rect 119266 11130 119276 12106
rect 119322 12054 119332 12202
rect 119474 12184 120116 12202
rect 119474 12054 119484 12184
rect 120104 12156 120116 12184
rect 120150 12262 120162 12299
rect 120524 12300 121472 12305
rect 120524 12299 120956 12300
rect 120524 12262 120536 12299
rect 120150 12184 120536 12262
rect 120150 12156 120162 12184
rect 120104 12150 120162 12156
rect 120524 12156 120536 12184
rect 120570 12265 120956 12299
rect 121040 12266 121376 12300
rect 121460 12266 121472 12300
rect 120990 12265 121376 12266
rect 121410 12265 121472 12266
rect 120570 12258 121472 12265
rect 121590 12306 121776 13386
rect 122026 13334 122072 13346
rect 122122 13334 122168 13346
rect 122236 13334 122282 13346
rect 122332 13334 122378 13346
rect 122446 13334 122492 13346
rect 122542 13334 122588 13346
rect 122656 13334 122702 13346
rect 122752 13334 122798 13346
rect 122866 13334 122912 13346
rect 122962 13334 123008 13346
rect 123076 13334 123122 13346
rect 123172 13334 123218 13346
rect 123286 13334 123332 13346
rect 123382 13334 123428 13346
rect 123496 13334 123542 13346
rect 123592 13334 123638 13346
rect 123706 13334 123752 13346
rect 123802 13334 123848 13346
rect 123916 13334 123962 13346
rect 124012 13334 124058 13346
rect 124126 13334 124172 13346
rect 124222 13334 124268 13346
rect 124336 13334 124382 13346
rect 124432 13334 124478 13346
rect 124546 13334 124592 13346
rect 124642 13334 124688 13346
rect 124756 13334 124802 13346
rect 124852 13334 124898 13346
rect 124966 13334 125012 13346
rect 125062 13334 125108 13346
rect 125176 13334 125222 13346
rect 125272 13334 125318 13346
rect 125386 13334 125432 13346
rect 125482 13334 125528 13346
rect 125596 13334 125642 13346
rect 125692 13334 125738 13346
rect 121998 12358 122008 13334
rect 122066 12358 122076 13334
rect 122118 12358 122128 13334
rect 122276 12358 122286 13334
rect 122328 12358 122338 13334
rect 122486 12358 122496 13334
rect 122538 12358 122548 13334
rect 122696 12358 122706 13334
rect 122748 12358 122758 13334
rect 122906 12358 122916 13334
rect 122958 12358 122968 13334
rect 123116 12358 123126 13334
rect 123168 12358 123178 13334
rect 123326 12358 123336 13334
rect 123378 12358 123388 13334
rect 123536 12358 123546 13334
rect 123588 12358 123598 13334
rect 123746 12358 123756 13334
rect 123798 12358 123808 13334
rect 123956 12358 123966 13334
rect 124008 12358 124018 13334
rect 124166 12358 124176 13334
rect 124218 12358 124228 13334
rect 124376 12358 124386 13334
rect 124428 12358 124438 13334
rect 124586 12358 124596 13334
rect 124638 12358 124648 13334
rect 124796 12358 124806 13334
rect 124848 12358 124858 13334
rect 125006 12358 125016 13334
rect 125058 12358 125068 13334
rect 125216 12358 125226 13334
rect 125268 12358 125278 13334
rect 125426 12358 125436 13334
rect 125478 12358 125488 13334
rect 125636 12358 125646 13334
rect 125688 12358 125698 13334
rect 125756 12358 125766 13334
rect 122026 12346 122072 12358
rect 122122 12346 122168 12358
rect 122236 12346 122282 12358
rect 122332 12346 122378 12358
rect 122446 12346 122492 12358
rect 122542 12346 122588 12358
rect 122656 12346 122702 12358
rect 122752 12346 122798 12358
rect 122866 12346 122912 12358
rect 122962 12346 123008 12358
rect 123076 12346 123122 12358
rect 123172 12346 123218 12358
rect 123286 12346 123332 12358
rect 123382 12346 123428 12358
rect 123496 12346 123542 12358
rect 123592 12346 123638 12358
rect 123706 12346 123752 12358
rect 123802 12346 123848 12358
rect 123916 12346 123962 12358
rect 124012 12346 124058 12358
rect 124126 12346 124172 12358
rect 124222 12346 124268 12358
rect 124336 12346 124382 12358
rect 124432 12346 124478 12358
rect 124546 12346 124592 12358
rect 124642 12346 124688 12358
rect 124756 12346 124802 12358
rect 124852 12346 124898 12358
rect 124966 12346 125012 12358
rect 125062 12346 125108 12358
rect 125176 12346 125222 12358
rect 125272 12346 125318 12358
rect 125386 12346 125432 12358
rect 125482 12346 125528 12358
rect 125596 12346 125642 12358
rect 125692 12346 125738 12358
rect 121590 12299 125696 12306
rect 120570 12196 120576 12258
rect 120570 12156 120582 12196
rect 120524 12150 120582 12156
rect 121590 12157 122290 12299
rect 122324 12157 122710 12299
rect 122744 12157 123130 12299
rect 123164 12157 123550 12299
rect 123584 12157 123970 12299
rect 124004 12157 124390 12299
rect 124424 12157 124810 12299
rect 124844 12157 125230 12299
rect 125264 12157 125650 12299
rect 125684 12157 125696 12299
rect 121590 12156 125696 12157
rect 120062 12106 120108 12118
rect 120158 12106 120204 12118
rect 120272 12106 120318 12118
rect 120368 12106 120414 12118
rect 120482 12106 120528 12118
rect 120578 12106 120624 12118
rect 120692 12106 120738 12118
rect 120788 12106 120834 12118
rect 119118 11118 119164 11130
rect 119206 11118 119252 11130
rect 119322 11086 119436 12054
rect 120038 11130 120048 12106
rect 120102 11130 120112 12106
rect 120154 11130 120164 12106
rect 120312 11130 120322 12106
rect 120364 11130 120374 12106
rect 120522 11130 120532 12106
rect 120574 11130 120584 12106
rect 120732 11130 120742 12106
rect 120784 11130 120794 12106
rect 120848 11130 120858 12106
rect 121254 11694 121264 11958
rect 121546 11938 121556 11958
rect 121590 11938 121776 12156
rect 122278 12151 122336 12156
rect 122698 12151 122756 12156
rect 123118 12151 123176 12156
rect 123538 12151 123596 12156
rect 123958 12151 124016 12156
rect 124378 12151 124436 12156
rect 124798 12151 124856 12156
rect 125218 12151 125276 12156
rect 125638 12151 125696 12156
rect 122026 12098 122072 12110
rect 122122 12098 122168 12110
rect 122236 12098 122282 12110
rect 122332 12098 122378 12110
rect 122446 12098 122492 12110
rect 122542 12098 122588 12110
rect 122656 12098 122702 12110
rect 122752 12098 122798 12110
rect 122866 12098 122912 12110
rect 122962 12098 123008 12110
rect 123076 12098 123122 12110
rect 123172 12098 123218 12110
rect 123286 12098 123332 12110
rect 123382 12098 123428 12110
rect 123496 12098 123542 12110
rect 123592 12098 123638 12110
rect 123706 12098 123752 12110
rect 123802 12098 123848 12110
rect 123916 12098 123962 12110
rect 124012 12098 124058 12110
rect 124126 12098 124172 12110
rect 124222 12098 124268 12110
rect 124336 12098 124382 12110
rect 124432 12098 124478 12110
rect 124546 12098 124592 12110
rect 124642 12098 124688 12110
rect 124756 12098 124802 12110
rect 124852 12098 124898 12110
rect 124966 12098 125012 12110
rect 125062 12098 125108 12110
rect 125176 12098 125222 12110
rect 125272 12098 125318 12110
rect 125386 12098 125432 12110
rect 125482 12098 125528 12110
rect 125596 12098 125642 12110
rect 125692 12098 125738 12110
rect 121546 11722 121776 11938
rect 121546 11694 121556 11722
rect 120062 11118 120108 11130
rect 120158 11118 120204 11130
rect 120272 11118 120318 11130
rect 120368 11118 120414 11130
rect 120482 11118 120528 11130
rect 120578 11118 120624 11130
rect 120692 11118 120738 11130
rect 120788 11118 120834 11130
rect 119322 11072 120842 11086
rect 119322 11037 120326 11072
rect 120410 11038 120746 11072
rect 120830 11038 120842 11072
rect 120360 11037 120746 11038
rect 120780 11037 120842 11038
rect 119322 11030 120842 11037
rect 121590 11072 121776 11722
rect 121998 11122 122008 12098
rect 122066 11122 122076 12098
rect 122118 11122 122128 12098
rect 122276 11122 122286 12098
rect 122328 11122 122338 12098
rect 122486 11122 122496 12098
rect 122538 11122 122548 12098
rect 122696 11122 122706 12098
rect 122748 11122 122758 12098
rect 122906 11122 122916 12098
rect 122958 11122 122968 12098
rect 123116 11122 123126 12098
rect 123168 11122 123178 12098
rect 123326 11122 123336 12098
rect 123378 11122 123388 12098
rect 123536 11122 123546 12098
rect 123588 11122 123598 12098
rect 123746 11122 123756 12098
rect 123798 11122 123808 12098
rect 123956 11122 123966 12098
rect 124008 11122 124018 12098
rect 124166 11122 124176 12098
rect 124218 11122 124228 12098
rect 124376 11122 124386 12098
rect 124428 11122 124438 12098
rect 124586 11122 124596 12098
rect 124638 11122 124648 12098
rect 124796 11122 124806 12098
rect 124848 11122 124858 12098
rect 125006 11122 125016 12098
rect 125058 11122 125068 12098
rect 125216 11122 125226 12098
rect 125268 11122 125278 12098
rect 125426 11122 125436 12098
rect 125478 11122 125488 12098
rect 125636 11122 125646 12098
rect 125688 11122 125698 12098
rect 125756 11122 125766 12098
rect 122026 11110 122072 11122
rect 122122 11110 122168 11122
rect 122236 11110 122282 11122
rect 122332 11110 122378 11122
rect 122446 11110 122492 11122
rect 122542 11110 122588 11122
rect 122656 11110 122702 11122
rect 122752 11110 122798 11122
rect 122866 11110 122912 11122
rect 122962 11110 123008 11122
rect 123076 11110 123122 11122
rect 123172 11110 123218 11122
rect 123286 11110 123332 11122
rect 123382 11110 123428 11122
rect 123496 11110 123542 11122
rect 123592 11110 123638 11122
rect 123706 11110 123752 11122
rect 123802 11110 123848 11122
rect 123916 11110 123962 11122
rect 124012 11110 124058 11122
rect 124126 11110 124172 11122
rect 124222 11110 124268 11122
rect 124336 11110 124382 11122
rect 124432 11110 124478 11122
rect 124546 11110 124592 11122
rect 124642 11110 124688 11122
rect 124756 11110 124802 11122
rect 124852 11110 124898 11122
rect 124966 11110 125012 11122
rect 125062 11110 125108 11122
rect 125176 11110 125222 11122
rect 125272 11110 125318 11122
rect 125386 11110 125432 11122
rect 125482 11110 125528 11122
rect 125596 11110 125642 11122
rect 125692 11110 125738 11122
rect 121590 11064 125636 11072
rect 121590 11029 122080 11064
rect 122164 11030 122500 11064
rect 122584 11030 122920 11064
rect 123004 11030 123340 11064
rect 123424 11030 123760 11064
rect 123844 11030 124180 11064
rect 124264 11030 124600 11064
rect 124684 11030 125020 11064
rect 125104 11030 125440 11064
rect 125524 11030 125636 11064
rect 122114 11029 122500 11030
rect 122534 11029 122920 11030
rect 122954 11029 123340 11030
rect 123374 11029 123760 11030
rect 123794 11029 124180 11030
rect 124214 11029 124600 11030
rect 124634 11029 125020 11030
rect 125054 11029 125440 11030
rect 125474 11029 125636 11030
rect 121590 11022 125636 11029
rect 119476 10942 119798 10948
rect 119476 10660 119488 10942
rect 119786 10660 119798 10942
rect 119476 10654 119798 10660
rect 121590 9186 121776 11022
rect 121590 9172 125636 9186
rect 121590 9137 122080 9172
rect 122164 9138 122500 9172
rect 122584 9138 122920 9172
rect 123004 9138 123340 9172
rect 123424 9138 123760 9172
rect 123844 9138 124180 9172
rect 124264 9138 124600 9172
rect 124684 9138 125020 9172
rect 125104 9138 125440 9172
rect 125524 9138 125636 9172
rect 122114 9137 122500 9138
rect 122534 9137 122920 9138
rect 121590 9132 122920 9137
rect 122954 9132 123340 9138
rect 123374 9132 123760 9138
rect 123794 9132 124180 9138
rect 124214 9132 124600 9138
rect 124634 9132 125020 9138
rect 125054 9132 125440 9138
rect 125474 9132 125636 9138
rect 121590 9126 125636 9132
rect 121590 8062 121776 9126
rect 122026 9082 122072 9094
rect 122122 9082 122168 9094
rect 122236 9082 122282 9094
rect 122332 9082 122378 9094
rect 122446 9082 122492 9094
rect 122542 9082 122588 9094
rect 122656 9082 122702 9094
rect 122752 9082 122798 9094
rect 122866 9082 122912 9094
rect 122962 9082 123008 9094
rect 123076 9082 123122 9094
rect 123172 9082 123218 9094
rect 123286 9082 123332 9094
rect 123382 9082 123428 9094
rect 123496 9082 123542 9094
rect 123592 9082 123638 9094
rect 123706 9082 123752 9094
rect 123802 9082 123848 9094
rect 123916 9082 123962 9094
rect 124012 9082 124058 9094
rect 124126 9082 124172 9094
rect 124222 9082 124268 9094
rect 124336 9082 124382 9094
rect 124432 9082 124478 9094
rect 124546 9082 124592 9094
rect 124642 9082 124688 9094
rect 124756 9082 124802 9094
rect 124852 9082 124898 9094
rect 124966 9082 125012 9094
rect 125062 9082 125108 9094
rect 125176 9082 125222 9094
rect 125272 9082 125318 9094
rect 125386 9082 125432 9094
rect 125482 9082 125528 9094
rect 125596 9082 125642 9094
rect 125692 9082 125738 9094
rect 121998 8106 122008 9082
rect 122066 8106 122076 9082
rect 122118 8106 122128 9082
rect 122276 8106 122286 9082
rect 122328 8106 122338 9082
rect 122486 8106 122496 9082
rect 122538 8106 122548 9082
rect 122696 8106 122706 9082
rect 122748 8106 122758 9082
rect 122906 8106 122916 9082
rect 122958 8106 122968 9082
rect 123116 8106 123126 9082
rect 123168 8106 123178 9082
rect 123326 8106 123336 9082
rect 123378 8106 123388 9082
rect 123536 8106 123546 9082
rect 123588 8106 123598 9082
rect 123746 8106 123756 9082
rect 123798 8106 123808 9082
rect 123956 8106 123966 9082
rect 124008 8106 124018 9082
rect 124166 8106 124176 9082
rect 124218 8106 124228 9082
rect 124376 8106 124386 9082
rect 124428 8106 124438 9082
rect 124586 8106 124596 9082
rect 124638 8106 124648 9082
rect 124796 8106 124806 9082
rect 124848 8106 124858 9082
rect 125006 8106 125016 9082
rect 125058 8106 125068 9082
rect 125216 8106 125226 9082
rect 125268 8106 125278 9082
rect 125426 8106 125436 9082
rect 125478 8106 125488 9082
rect 125636 8106 125646 9082
rect 125688 8106 125698 9082
rect 125756 8106 125766 9082
rect 122026 8094 122072 8106
rect 122122 8094 122168 8106
rect 122236 8094 122282 8106
rect 122332 8094 122378 8106
rect 122446 8094 122492 8106
rect 122542 8094 122588 8106
rect 122656 8094 122702 8106
rect 122752 8094 122798 8106
rect 122866 8094 122912 8106
rect 122962 8094 123008 8106
rect 123076 8094 123122 8106
rect 123172 8094 123218 8106
rect 123286 8094 123332 8106
rect 123382 8094 123428 8106
rect 123496 8094 123542 8106
rect 123592 8094 123638 8106
rect 123706 8094 123752 8106
rect 123802 8094 123848 8106
rect 123916 8094 123962 8106
rect 124012 8094 124058 8106
rect 124126 8094 124172 8106
rect 124222 8094 124268 8106
rect 124336 8094 124382 8106
rect 124432 8094 124478 8106
rect 124546 8094 124592 8106
rect 124642 8094 124688 8106
rect 124756 8094 124802 8106
rect 124852 8094 124898 8106
rect 124966 8094 125012 8106
rect 125062 8094 125108 8106
rect 125176 8094 125222 8106
rect 125272 8094 125318 8106
rect 125386 8094 125432 8106
rect 125482 8094 125528 8106
rect 125596 8094 125642 8106
rect 125692 8094 125738 8106
rect 121590 8056 125750 8062
rect 121590 8048 122710 8056
rect 122744 8048 123130 8056
rect 123164 8048 123550 8056
rect 123584 8048 123970 8056
rect 124004 8048 124390 8056
rect 124424 8048 124810 8056
rect 124844 8048 125230 8056
rect 125264 8048 125650 8056
rect 125684 8048 125750 8056
rect 121590 8014 122290 8048
rect 122374 8014 122710 8048
rect 122794 8014 123130 8048
rect 123214 8014 123550 8048
rect 123634 8014 123970 8048
rect 124054 8014 124390 8048
rect 124474 8014 124810 8048
rect 124894 8014 125230 8048
rect 125314 8014 125650 8048
rect 125734 8014 125750 8048
rect 121590 8006 125750 8014
rect 122016 7928 122140 7934
rect 122016 7828 122028 7928
rect 122128 7828 122140 7928
rect 122016 7822 122140 7828
rect 122436 7928 122560 7934
rect 122436 7828 122448 7928
rect 122548 7828 122560 7928
rect 122436 7822 122560 7828
rect 122856 7928 122980 7934
rect 122856 7828 122868 7928
rect 122968 7828 122980 7928
rect 122856 7822 122980 7828
rect 123276 7928 123400 7934
rect 123276 7828 123288 7928
rect 123388 7828 123400 7928
rect 123276 7822 123400 7828
rect 123696 7928 123820 7934
rect 123696 7828 123708 7928
rect 123808 7828 123820 7928
rect 123696 7822 123820 7828
rect 124116 7928 124240 7934
rect 124116 7828 124128 7928
rect 124228 7828 124240 7928
rect 124116 7822 124240 7828
rect 124536 7928 124660 7934
rect 124536 7828 124548 7928
rect 124648 7828 124660 7928
rect 124536 7822 124660 7828
rect 124956 7928 125080 7934
rect 124956 7828 124968 7928
rect 125068 7828 125080 7928
rect 124956 7822 125080 7828
rect 125376 7928 125500 7934
rect 125376 7828 125388 7928
rect 125488 7828 125500 7928
rect 125376 7822 125500 7828
rect 125702 7928 125826 7934
rect 125702 7828 125714 7928
rect 125814 7828 125826 7928
rect 125702 7822 125826 7828
<< via1 >>
rect 126840 28200 126938 28304
rect 127260 28200 127358 28304
rect 127680 28200 127778 28304
rect 128100 28200 128198 28304
rect 128520 28200 128618 28304
rect 128940 28200 129038 28304
rect 129360 28200 129458 28304
rect 129780 28200 129878 28304
rect 130200 28200 130298 28304
rect 130620 28200 130718 28304
rect 131040 28200 131138 28304
rect 131460 28200 131558 28304
rect 131880 28200 131978 28304
rect 132300 28200 132398 28304
rect 132720 28200 132818 28304
rect 133140 28200 133238 28304
rect 133560 28200 133658 28304
rect 133980 28200 134078 28304
rect 134400 28200 134498 28304
rect 134820 28200 134918 28304
rect 135168 28200 135266 28304
rect 126858 26992 126882 27968
rect 126882 26992 126916 27968
rect 126978 26992 127012 27968
rect 127012 26992 127092 27968
rect 127092 26992 127126 27968
rect 127188 26992 127222 27968
rect 127222 26992 127302 27968
rect 127302 26992 127336 27968
rect 127398 26992 127432 27968
rect 127432 26992 127512 27968
rect 127512 26992 127546 27968
rect 127608 26992 127642 27968
rect 127642 26992 127722 27968
rect 127722 26992 127756 27968
rect 127818 26992 127852 27968
rect 127852 26992 127932 27968
rect 127932 26992 127966 27968
rect 128028 26992 128062 27968
rect 128062 26992 128142 27968
rect 128142 26992 128176 27968
rect 128238 26992 128272 27968
rect 128272 26992 128352 27968
rect 128352 26992 128386 27968
rect 128448 26992 128482 27968
rect 128482 26992 128562 27968
rect 128562 26992 128596 27968
rect 128658 26992 128692 27968
rect 128692 26992 128772 27968
rect 128772 26992 128806 27968
rect 128868 26992 128902 27968
rect 128902 26992 128982 27968
rect 128982 26992 129016 27968
rect 129078 26992 129112 27968
rect 129112 26992 129192 27968
rect 129192 26992 129226 27968
rect 129288 26992 129322 27968
rect 129322 26992 129402 27968
rect 129402 26992 129436 27968
rect 129498 26992 129532 27968
rect 129532 26992 129612 27968
rect 129612 26992 129646 27968
rect 129708 26992 129742 27968
rect 129742 26992 129822 27968
rect 129822 26992 129856 27968
rect 129918 26992 129952 27968
rect 129952 26992 130032 27968
rect 130032 26992 130066 27968
rect 130128 26992 130162 27968
rect 130162 26992 130242 27968
rect 130242 26992 130276 27968
rect 130338 26992 130372 27968
rect 130372 26992 130452 27968
rect 130452 26992 130486 27968
rect 130548 26992 130582 27968
rect 130582 26992 130662 27968
rect 130662 26992 130696 27968
rect 130758 26992 130792 27968
rect 130792 26992 130872 27968
rect 130872 26992 130906 27968
rect 130968 26992 131002 27968
rect 131002 26992 131082 27968
rect 131082 26992 131116 27968
rect 131178 26992 131212 27968
rect 131212 26992 131292 27968
rect 131292 26992 131326 27968
rect 131388 26992 131422 27968
rect 131422 26992 131502 27968
rect 131502 26992 131536 27968
rect 131598 26992 131632 27968
rect 131632 26992 131712 27968
rect 131712 26992 131746 27968
rect 131808 26992 131842 27968
rect 131842 26992 131922 27968
rect 131922 26992 131956 27968
rect 132018 26992 132052 27968
rect 132052 26992 132132 27968
rect 132132 26992 132166 27968
rect 132228 26992 132262 27968
rect 132262 26992 132342 27968
rect 132342 26992 132376 27968
rect 132438 26992 132472 27968
rect 132472 26992 132552 27968
rect 132552 26992 132586 27968
rect 132648 26992 132682 27968
rect 132682 26992 132762 27968
rect 132762 26992 132796 27968
rect 132858 26992 132892 27968
rect 132892 26992 132972 27968
rect 132972 26992 133006 27968
rect 133068 26992 133102 27968
rect 133102 26992 133182 27968
rect 133182 26992 133216 27968
rect 133278 26992 133312 27968
rect 133312 26992 133392 27968
rect 133392 26992 133426 27968
rect 133488 26992 133522 27968
rect 133522 26992 133602 27968
rect 133602 26992 133636 27968
rect 133698 26992 133732 27968
rect 133732 26992 133812 27968
rect 133812 26992 133846 27968
rect 133908 26992 133942 27968
rect 133942 26992 134022 27968
rect 134022 26992 134056 27968
rect 134118 26992 134152 27968
rect 134152 26992 134232 27968
rect 134232 26992 134266 27968
rect 134328 26992 134362 27968
rect 134362 26992 134442 27968
rect 134442 26992 134476 27968
rect 134538 26992 134572 27968
rect 134572 26992 134652 27968
rect 134652 26992 134686 27968
rect 134748 26992 134782 27968
rect 134782 26992 134862 27968
rect 134862 26992 134896 27968
rect 134958 26992 134992 27968
rect 134992 26992 135072 27968
rect 135072 26992 135106 27968
rect 135168 26992 135202 27968
rect 135202 26992 135226 27968
rect 126858 25774 126882 26750
rect 126882 25774 126916 26750
rect 126978 25774 127012 26750
rect 127012 25774 127092 26750
rect 127092 25774 127126 26750
rect 127188 25774 127222 26750
rect 127222 25774 127302 26750
rect 127302 25774 127336 26750
rect 127398 25774 127432 26750
rect 127432 25774 127512 26750
rect 127512 25774 127546 26750
rect 127608 25774 127642 26750
rect 127642 25774 127722 26750
rect 127722 25774 127756 26750
rect 127818 25774 127852 26750
rect 127852 25774 127932 26750
rect 127932 25774 127966 26750
rect 128028 25774 128062 26750
rect 128062 25774 128142 26750
rect 128142 25774 128176 26750
rect 128238 25774 128272 26750
rect 128272 25774 128352 26750
rect 128352 25774 128386 26750
rect 128448 25774 128482 26750
rect 128482 25774 128562 26750
rect 128562 25774 128596 26750
rect 128658 25774 128692 26750
rect 128692 25774 128772 26750
rect 128772 25774 128806 26750
rect 128868 25774 128902 26750
rect 128902 25774 128982 26750
rect 128982 25774 129016 26750
rect 129078 25774 129112 26750
rect 129112 25774 129192 26750
rect 129192 25774 129226 26750
rect 129288 25774 129322 26750
rect 129322 25774 129402 26750
rect 129402 25774 129436 26750
rect 129498 25774 129532 26750
rect 129532 25774 129612 26750
rect 129612 25774 129646 26750
rect 129708 25774 129742 26750
rect 129742 25774 129822 26750
rect 129822 25774 129856 26750
rect 129918 25774 129952 26750
rect 129952 25774 130032 26750
rect 130032 25774 130066 26750
rect 130128 25774 130162 26750
rect 130162 25774 130242 26750
rect 130242 25774 130276 26750
rect 130338 25774 130372 26750
rect 130372 25774 130452 26750
rect 130452 25774 130486 26750
rect 130548 25774 130582 26750
rect 130582 25774 130662 26750
rect 130662 25774 130696 26750
rect 130758 25774 130792 26750
rect 130792 25774 130872 26750
rect 130872 25774 130906 26750
rect 130968 25774 131002 26750
rect 131002 25774 131082 26750
rect 131082 25774 131116 26750
rect 131178 25774 131212 26750
rect 131212 25774 131292 26750
rect 131292 25774 131326 26750
rect 131388 25774 131422 26750
rect 131422 25774 131502 26750
rect 131502 25774 131536 26750
rect 131598 25774 131632 26750
rect 131632 25774 131712 26750
rect 131712 25774 131746 26750
rect 131808 25774 131842 26750
rect 131842 25774 131922 26750
rect 131922 25774 131956 26750
rect 132018 25774 132052 26750
rect 132052 25774 132132 26750
rect 132132 25774 132166 26750
rect 132228 25774 132262 26750
rect 132262 25774 132342 26750
rect 132342 25774 132376 26750
rect 132438 25774 132472 26750
rect 132472 25774 132552 26750
rect 132552 25774 132586 26750
rect 132648 25774 132682 26750
rect 132682 25774 132762 26750
rect 132762 25774 132796 26750
rect 132858 25774 132892 26750
rect 132892 25774 132972 26750
rect 132972 25774 133006 26750
rect 133068 25774 133102 26750
rect 133102 25774 133182 26750
rect 133182 25774 133216 26750
rect 133278 25774 133312 26750
rect 133312 25774 133392 26750
rect 133392 25774 133426 26750
rect 133488 25774 133522 26750
rect 133522 25774 133602 26750
rect 133602 25774 133636 26750
rect 133698 25774 133732 26750
rect 133732 25774 133812 26750
rect 133812 25774 133846 26750
rect 133908 25774 133942 26750
rect 133942 25774 134022 26750
rect 134022 25774 134056 26750
rect 134118 25774 134152 26750
rect 134152 25774 134232 26750
rect 134232 25774 134266 26750
rect 134328 25774 134362 26750
rect 134362 25774 134442 26750
rect 134442 25774 134476 26750
rect 134538 25774 134572 26750
rect 134572 25774 134652 26750
rect 134652 25774 134686 26750
rect 134748 25774 134782 26750
rect 134782 25774 134862 26750
rect 134862 25774 134896 26750
rect 134958 25774 134992 26750
rect 134992 25774 135072 26750
rect 135072 25774 135106 26750
rect 135168 25774 135202 26750
rect 135202 25774 135226 26750
rect 122028 22062 122128 22162
rect 122448 22062 122548 22162
rect 122868 22062 122968 22162
rect 123288 22062 123388 22162
rect 123708 22062 123808 22162
rect 124128 22062 124228 22162
rect 124548 22062 124648 22162
rect 124968 22062 125068 22162
rect 125388 22062 125488 22162
rect 125714 22062 125814 22162
rect 122008 20908 122032 21884
rect 122032 20908 122066 21884
rect 122128 20908 122162 21884
rect 122162 20908 122242 21884
rect 122242 20908 122276 21884
rect 122338 20908 122372 21884
rect 122372 20908 122452 21884
rect 122452 20908 122486 21884
rect 122548 20908 122582 21884
rect 122582 20908 122662 21884
rect 122662 20908 122696 21884
rect 122758 20908 122792 21884
rect 122792 20908 122872 21884
rect 122872 20908 122906 21884
rect 122968 20908 123002 21884
rect 123002 20908 123082 21884
rect 123082 20908 123116 21884
rect 123178 20908 123212 21884
rect 123212 20908 123292 21884
rect 123292 20908 123326 21884
rect 123388 20908 123422 21884
rect 123422 20908 123502 21884
rect 123502 20908 123536 21884
rect 123598 20908 123632 21884
rect 123632 20908 123712 21884
rect 123712 20908 123746 21884
rect 123808 20908 123842 21884
rect 123842 20908 123922 21884
rect 123922 20908 123956 21884
rect 124018 20908 124052 21884
rect 124052 20908 124132 21884
rect 124132 20908 124166 21884
rect 124228 20908 124262 21884
rect 124262 20908 124342 21884
rect 124342 20908 124376 21884
rect 124438 20908 124472 21884
rect 124472 20908 124552 21884
rect 124552 20908 124586 21884
rect 124648 20908 124682 21884
rect 124682 20908 124762 21884
rect 124762 20908 124796 21884
rect 124858 20908 124892 21884
rect 124892 20908 124972 21884
rect 124972 20908 125006 21884
rect 125068 20908 125102 21884
rect 125102 20908 125182 21884
rect 125182 20908 125216 21884
rect 125278 20908 125312 21884
rect 125312 20908 125392 21884
rect 125392 20908 125426 21884
rect 125488 20908 125522 21884
rect 125522 20908 125602 21884
rect 125602 20908 125636 21884
rect 125698 20908 125732 21884
rect 125732 20908 125756 21884
rect 126858 21764 126882 22740
rect 126882 21764 126916 22740
rect 126978 21764 127012 22740
rect 127012 21764 127092 22740
rect 127092 21764 127126 22740
rect 127188 21764 127222 22740
rect 127222 21764 127302 22740
rect 127302 21764 127336 22740
rect 127398 21764 127432 22740
rect 127432 21764 127512 22740
rect 127512 21764 127546 22740
rect 127608 21764 127642 22740
rect 127642 21764 127722 22740
rect 127722 21764 127756 22740
rect 127818 21764 127852 22740
rect 127852 21764 127932 22740
rect 127932 21764 127966 22740
rect 128028 21764 128062 22740
rect 128062 21764 128142 22740
rect 128142 21764 128176 22740
rect 128238 21764 128272 22740
rect 128272 21764 128352 22740
rect 128352 21764 128386 22740
rect 128448 21764 128482 22740
rect 128482 21764 128562 22740
rect 128562 21764 128596 22740
rect 128658 21764 128692 22740
rect 128692 21764 128772 22740
rect 128772 21764 128806 22740
rect 128868 21764 128902 22740
rect 128902 21764 128982 22740
rect 128982 21764 129016 22740
rect 129078 21764 129112 22740
rect 129112 21764 129192 22740
rect 129192 21764 129226 22740
rect 129288 21764 129322 22740
rect 129322 21764 129402 22740
rect 129402 21764 129436 22740
rect 129498 21764 129532 22740
rect 129532 21764 129612 22740
rect 129612 21764 129646 22740
rect 129708 21764 129742 22740
rect 129742 21764 129822 22740
rect 129822 21764 129856 22740
rect 129918 21764 129952 22740
rect 129952 21764 130032 22740
rect 130032 21764 130066 22740
rect 130128 21764 130162 22740
rect 130162 21764 130242 22740
rect 130242 21764 130276 22740
rect 130338 21764 130372 22740
rect 130372 21764 130452 22740
rect 130452 21764 130486 22740
rect 130548 21764 130582 22740
rect 130582 21764 130662 22740
rect 130662 21764 130696 22740
rect 130758 21764 130792 22740
rect 130792 21764 130872 22740
rect 130872 21764 130906 22740
rect 130968 21764 131002 22740
rect 131002 21764 131082 22740
rect 131082 21764 131116 22740
rect 131178 21764 131212 22740
rect 131212 21764 131292 22740
rect 131292 21764 131326 22740
rect 131388 21764 131422 22740
rect 131422 21764 131502 22740
rect 131502 21764 131536 22740
rect 131598 21764 131632 22740
rect 131632 21764 131712 22740
rect 131712 21764 131746 22740
rect 131808 21764 131842 22740
rect 131842 21764 131922 22740
rect 131922 21764 131956 22740
rect 132018 21764 132052 22740
rect 132052 21764 132132 22740
rect 132132 21764 132166 22740
rect 132228 21764 132262 22740
rect 132262 21764 132342 22740
rect 132342 21764 132376 22740
rect 132438 21764 132472 22740
rect 132472 21764 132552 22740
rect 132552 21764 132586 22740
rect 132648 21764 132682 22740
rect 132682 21764 132762 22740
rect 132762 21764 132796 22740
rect 132858 21764 132892 22740
rect 132892 21764 132972 22740
rect 132972 21764 133006 22740
rect 133068 21764 133102 22740
rect 133102 21764 133182 22740
rect 133182 21764 133216 22740
rect 133278 21764 133312 22740
rect 133312 21764 133392 22740
rect 133392 21764 133426 22740
rect 133488 21764 133522 22740
rect 133522 21764 133602 22740
rect 133602 21764 133636 22740
rect 133698 21764 133732 22740
rect 133732 21764 133812 22740
rect 133812 21764 133846 22740
rect 133908 21764 133942 22740
rect 133942 21764 134022 22740
rect 134022 21764 134056 22740
rect 134118 21764 134152 22740
rect 134152 21764 134232 22740
rect 134232 21764 134266 22740
rect 134328 21764 134362 22740
rect 134362 21764 134442 22740
rect 134442 21764 134476 22740
rect 134538 21764 134572 22740
rect 134572 21764 134652 22740
rect 134652 21764 134686 22740
rect 134748 21764 134782 22740
rect 134782 21764 134862 22740
rect 134862 21764 134896 22740
rect 134958 21764 134992 22740
rect 134992 21764 135072 22740
rect 135072 21764 135106 22740
rect 135168 21764 135202 22740
rect 135202 21764 135226 22740
rect 119488 20448 119786 20730
rect 119104 19284 119124 20260
rect 119124 19284 119158 20260
rect 119212 19284 119246 20260
rect 119246 19284 119266 20260
rect 119332 19188 119474 19336
rect 120048 19284 120068 20260
rect 120068 19284 120102 20260
rect 120164 19284 120198 20260
rect 120198 19284 120278 20260
rect 120278 19284 120312 20260
rect 120374 19284 120408 20260
rect 120408 19284 120488 20260
rect 120488 19284 120522 20260
rect 120584 19284 120618 20260
rect 120618 19284 120698 20260
rect 120698 19284 120732 20260
rect 120794 19284 120828 20260
rect 120828 19284 120848 20260
rect 121264 19432 121546 19696
rect 125864 20310 126474 20928
rect 126858 20528 126882 21504
rect 126882 20528 126916 21504
rect 126978 20528 127012 21504
rect 127012 20528 127092 21504
rect 127092 20528 127126 21504
rect 127188 20528 127222 21504
rect 127222 20528 127302 21504
rect 127302 20528 127336 21504
rect 127398 20528 127432 21504
rect 127432 20528 127512 21504
rect 127512 20528 127546 21504
rect 127608 20528 127642 21504
rect 127642 20528 127722 21504
rect 127722 20528 127756 21504
rect 127818 20528 127852 21504
rect 127852 20528 127932 21504
rect 127932 20528 127966 21504
rect 128028 20528 128062 21504
rect 128062 20528 128142 21504
rect 128142 20528 128176 21504
rect 128238 20528 128272 21504
rect 128272 20528 128352 21504
rect 128352 20528 128386 21504
rect 128448 20528 128482 21504
rect 128482 20528 128562 21504
rect 128562 20528 128596 21504
rect 128658 20528 128692 21504
rect 128692 20528 128772 21504
rect 128772 20528 128806 21504
rect 128868 20528 128902 21504
rect 128902 20528 128982 21504
rect 128982 20528 129016 21504
rect 129078 20528 129112 21504
rect 129112 20528 129192 21504
rect 129192 20528 129226 21504
rect 129288 20528 129322 21504
rect 129322 20528 129402 21504
rect 129402 20528 129436 21504
rect 129498 20528 129532 21504
rect 129532 20528 129612 21504
rect 129612 20528 129646 21504
rect 129708 20528 129742 21504
rect 129742 20528 129822 21504
rect 129822 20528 129856 21504
rect 129918 20528 129952 21504
rect 129952 20528 130032 21504
rect 130032 20528 130066 21504
rect 130128 20528 130162 21504
rect 130162 20528 130242 21504
rect 130242 20528 130276 21504
rect 130338 20528 130372 21504
rect 130372 20528 130452 21504
rect 130452 20528 130486 21504
rect 130548 20528 130582 21504
rect 130582 20528 130662 21504
rect 130662 20528 130696 21504
rect 130758 20528 130792 21504
rect 130792 20528 130872 21504
rect 130872 20528 130906 21504
rect 130968 20528 131002 21504
rect 131002 20528 131082 21504
rect 131082 20528 131116 21504
rect 131178 20528 131212 21504
rect 131212 20528 131292 21504
rect 131292 20528 131326 21504
rect 131388 20528 131422 21504
rect 131422 20528 131502 21504
rect 131502 20528 131536 21504
rect 131598 20528 131632 21504
rect 131632 20528 131712 21504
rect 131712 20528 131746 21504
rect 131808 20528 131842 21504
rect 131842 20528 131922 21504
rect 131922 20528 131956 21504
rect 132018 20528 132052 21504
rect 132052 20528 132132 21504
rect 132132 20528 132166 21504
rect 132228 20528 132262 21504
rect 132262 20528 132342 21504
rect 132342 20528 132376 21504
rect 132438 20528 132472 21504
rect 132472 20528 132552 21504
rect 132552 20528 132586 21504
rect 132648 20528 132682 21504
rect 132682 20528 132762 21504
rect 132762 20528 132796 21504
rect 132858 20528 132892 21504
rect 132892 20528 132972 21504
rect 132972 20528 133006 21504
rect 133068 20528 133102 21504
rect 133102 20528 133182 21504
rect 133182 20528 133216 21504
rect 133278 20528 133312 21504
rect 133312 20528 133392 21504
rect 133392 20528 133426 21504
rect 133488 20528 133522 21504
rect 133522 20528 133602 21504
rect 133602 20528 133636 21504
rect 133698 20528 133732 21504
rect 133732 20528 133812 21504
rect 133812 20528 133846 21504
rect 133908 20528 133942 21504
rect 133942 20528 134022 21504
rect 134022 20528 134056 21504
rect 134118 20528 134152 21504
rect 134152 20528 134232 21504
rect 134232 20528 134266 21504
rect 134328 20528 134362 21504
rect 134362 20528 134442 21504
rect 134442 20528 134476 21504
rect 134538 20528 134572 21504
rect 134572 20528 134652 21504
rect 134652 20528 134686 21504
rect 134748 20528 134782 21504
rect 134782 20528 134862 21504
rect 134862 20528 134896 21504
rect 134958 20528 134992 21504
rect 134992 20528 135072 21504
rect 135072 20528 135106 21504
rect 135168 20528 135202 21504
rect 135202 20528 135226 21504
rect 119082 18056 119120 19032
rect 119120 18056 119154 19032
rect 119206 18056 119216 19032
rect 119216 18056 119250 19032
rect 119250 18056 119260 19032
rect 119312 18056 119346 19032
rect 119346 18056 119384 19032
rect 122008 19292 122032 20268
rect 122032 19292 122066 20268
rect 122128 19292 122162 20268
rect 122162 19292 122242 20268
rect 122242 19292 122276 20268
rect 122338 19292 122372 20268
rect 122372 19292 122452 20268
rect 122452 19292 122486 20268
rect 122548 19292 122582 20268
rect 122582 19292 122662 20268
rect 122662 19292 122696 20268
rect 122758 19292 122792 20268
rect 122792 19292 122872 20268
rect 122872 19292 122906 20268
rect 122968 19292 123002 20268
rect 123002 19292 123082 20268
rect 123082 19292 123116 20268
rect 123178 19292 123212 20268
rect 123212 19292 123292 20268
rect 123292 19292 123326 20268
rect 123388 19292 123422 20268
rect 123422 19292 123502 20268
rect 123502 19292 123536 20268
rect 123598 19292 123632 20268
rect 123632 19292 123712 20268
rect 123712 19292 123746 20268
rect 123808 19292 123842 20268
rect 123842 19292 123922 20268
rect 123922 19292 123956 20268
rect 124018 19292 124052 20268
rect 124052 19292 124132 20268
rect 124132 19292 124166 20268
rect 124228 19292 124262 20268
rect 124262 19292 124342 20268
rect 124342 19292 124376 20268
rect 124438 19292 124472 20268
rect 124472 19292 124552 20268
rect 124552 19292 124586 20268
rect 124648 19292 124682 20268
rect 124682 19292 124762 20268
rect 124762 19292 124796 20268
rect 124858 19292 124892 20268
rect 124892 19292 124972 20268
rect 124972 19292 125006 20268
rect 125068 19292 125102 20268
rect 125102 19292 125182 20268
rect 125182 19292 125216 20268
rect 125278 19292 125312 20268
rect 125312 19292 125392 20268
rect 125392 19292 125426 20268
rect 125488 19292 125522 20268
rect 125522 19292 125602 20268
rect 125602 19292 125636 20268
rect 125698 19292 125732 20268
rect 125732 19292 125756 20268
rect 126858 19292 126882 20268
rect 126882 19292 126916 20268
rect 126978 19292 127012 20268
rect 127012 19292 127092 20268
rect 127092 19292 127126 20268
rect 127188 19292 127222 20268
rect 127222 19292 127302 20268
rect 127302 19292 127336 20268
rect 127398 19292 127432 20268
rect 127432 19292 127512 20268
rect 127512 19292 127546 20268
rect 127608 19292 127642 20268
rect 127642 19292 127722 20268
rect 127722 19292 127756 20268
rect 127818 19292 127852 20268
rect 127852 19292 127932 20268
rect 127932 19292 127966 20268
rect 128028 19292 128062 20268
rect 128062 19292 128142 20268
rect 128142 19292 128176 20268
rect 128238 19292 128272 20268
rect 128272 19292 128352 20268
rect 128352 19292 128386 20268
rect 128448 19292 128482 20268
rect 128482 19292 128562 20268
rect 128562 19292 128596 20268
rect 128658 19292 128692 20268
rect 128692 19292 128772 20268
rect 128772 19292 128806 20268
rect 128868 19292 128902 20268
rect 128902 19292 128982 20268
rect 128982 19292 129016 20268
rect 129078 19292 129112 20268
rect 129112 19292 129192 20268
rect 129192 19292 129226 20268
rect 129288 19292 129322 20268
rect 129322 19292 129402 20268
rect 129402 19292 129436 20268
rect 129498 19292 129532 20268
rect 129532 19292 129612 20268
rect 129612 19292 129646 20268
rect 129708 19292 129742 20268
rect 129742 19292 129822 20268
rect 129822 19292 129856 20268
rect 129918 19292 129952 20268
rect 129952 19292 130032 20268
rect 130032 19292 130066 20268
rect 130128 19292 130162 20268
rect 130162 19292 130242 20268
rect 130242 19292 130276 20268
rect 130338 19292 130372 20268
rect 130372 19292 130452 20268
rect 130452 19292 130486 20268
rect 130548 19292 130582 20268
rect 130582 19292 130662 20268
rect 130662 19292 130696 20268
rect 130758 19292 130792 20268
rect 130792 19292 130872 20268
rect 130872 19292 130906 20268
rect 130968 19292 131002 20268
rect 131002 19292 131082 20268
rect 131082 19292 131116 20268
rect 131178 19292 131212 20268
rect 131212 19292 131292 20268
rect 131292 19292 131326 20268
rect 131388 19292 131422 20268
rect 131422 19292 131502 20268
rect 131502 19292 131536 20268
rect 131598 19292 131632 20268
rect 131632 19292 131712 20268
rect 131712 19292 131746 20268
rect 131808 19292 131842 20268
rect 131842 19292 131922 20268
rect 131922 19292 131956 20268
rect 132018 19292 132052 20268
rect 132052 19292 132132 20268
rect 132132 19292 132166 20268
rect 132228 19292 132262 20268
rect 132262 19292 132342 20268
rect 132342 19292 132376 20268
rect 132438 19292 132472 20268
rect 132472 19292 132552 20268
rect 132552 19292 132586 20268
rect 132648 19292 132682 20268
rect 132682 19292 132762 20268
rect 132762 19292 132796 20268
rect 132858 19292 132892 20268
rect 132892 19292 132972 20268
rect 132972 19292 133006 20268
rect 133068 19292 133102 20268
rect 133102 19292 133182 20268
rect 133182 19292 133216 20268
rect 133278 19292 133312 20268
rect 133312 19292 133392 20268
rect 133392 19292 133426 20268
rect 133488 19292 133522 20268
rect 133522 19292 133602 20268
rect 133602 19292 133636 20268
rect 133698 19292 133732 20268
rect 133732 19292 133812 20268
rect 133812 19292 133846 20268
rect 133908 19292 133942 20268
rect 133942 19292 134022 20268
rect 134022 19292 134056 20268
rect 134118 19292 134152 20268
rect 134152 19292 134232 20268
rect 134232 19292 134266 20268
rect 134328 19292 134362 20268
rect 134362 19292 134442 20268
rect 134442 19292 134476 20268
rect 134538 19292 134572 20268
rect 134572 19292 134652 20268
rect 134652 19292 134686 20268
rect 134748 19292 134782 20268
rect 134782 19292 134862 20268
rect 134862 19292 134896 20268
rect 134958 19292 134992 20268
rect 134992 19292 135072 20268
rect 135072 19292 135106 20268
rect 135168 19292 135202 20268
rect 135202 19292 135226 20268
rect 119834 18056 119858 19032
rect 119858 18056 119892 19032
rect 119954 18056 119988 19032
rect 119988 18056 120068 19032
rect 120068 18056 120102 19032
rect 120164 18056 120198 19032
rect 120198 18056 120278 19032
rect 120278 18056 120312 19032
rect 120374 18056 120408 19032
rect 120408 18056 120488 19032
rect 120488 18056 120522 19032
rect 120584 18056 120618 19032
rect 120618 18056 120698 19032
rect 120698 18056 120732 19032
rect 120794 18056 120828 19032
rect 120828 18056 120908 19032
rect 120908 18056 120942 19032
rect 121004 18056 121038 19032
rect 121038 18056 121118 19032
rect 121118 18056 121152 19032
rect 121214 18056 121248 19032
rect 121248 18056 121328 19032
rect 121328 18056 121362 19032
rect 121424 18056 121458 19032
rect 121458 18056 121482 19032
rect 122008 18056 122032 19032
rect 122032 18056 122066 19032
rect 122128 18056 122162 19032
rect 122162 18056 122242 19032
rect 122242 18056 122276 19032
rect 122338 18056 122372 19032
rect 122372 18056 122452 19032
rect 122452 18056 122486 19032
rect 122548 18056 122582 19032
rect 122582 18056 122662 19032
rect 122662 18056 122696 19032
rect 122758 18056 122792 19032
rect 122792 18056 122872 19032
rect 122872 18056 122906 19032
rect 122968 18056 123002 19032
rect 123002 18056 123082 19032
rect 123082 18056 123116 19032
rect 123178 18056 123212 19032
rect 123212 18056 123292 19032
rect 123292 18056 123326 19032
rect 123388 18056 123422 19032
rect 123422 18056 123502 19032
rect 123502 18056 123536 19032
rect 123598 18056 123632 19032
rect 123632 18056 123712 19032
rect 123712 18056 123746 19032
rect 123808 18056 123842 19032
rect 123842 18056 123922 19032
rect 123922 18056 123956 19032
rect 124018 18056 124052 19032
rect 124052 18056 124132 19032
rect 124132 18056 124166 19032
rect 124228 18056 124262 19032
rect 124262 18056 124342 19032
rect 124342 18056 124376 19032
rect 124438 18056 124472 19032
rect 124472 18056 124552 19032
rect 124552 18056 124586 19032
rect 124648 18056 124682 19032
rect 124682 18056 124762 19032
rect 124762 18056 124796 19032
rect 124858 18056 124892 19032
rect 124892 18056 124972 19032
rect 124972 18056 125006 19032
rect 125068 18056 125102 19032
rect 125102 18056 125182 19032
rect 125182 18056 125216 19032
rect 125278 18056 125312 19032
rect 125312 18056 125392 19032
rect 125392 18056 125426 19032
rect 125488 18056 125522 19032
rect 125522 18056 125602 19032
rect 125602 18056 125636 19032
rect 125698 18056 125732 19032
rect 125732 18056 125756 19032
rect 126858 18056 126882 19032
rect 126882 18056 126916 19032
rect 126978 18056 127012 19032
rect 127012 18056 127092 19032
rect 127092 18056 127126 19032
rect 127188 18056 127222 19032
rect 127222 18056 127302 19032
rect 127302 18056 127336 19032
rect 127398 18056 127432 19032
rect 127432 18056 127512 19032
rect 127512 18056 127546 19032
rect 127608 18056 127642 19032
rect 127642 18056 127722 19032
rect 127722 18056 127756 19032
rect 127818 18056 127852 19032
rect 127852 18056 127932 19032
rect 127932 18056 127966 19032
rect 128028 18056 128062 19032
rect 128062 18056 128142 19032
rect 128142 18056 128176 19032
rect 128238 18056 128272 19032
rect 128272 18056 128352 19032
rect 128352 18056 128386 19032
rect 128448 18056 128482 19032
rect 128482 18056 128562 19032
rect 128562 18056 128596 19032
rect 128658 18056 128692 19032
rect 128692 18056 128772 19032
rect 128772 18056 128806 19032
rect 128868 18056 128902 19032
rect 128902 18056 128982 19032
rect 128982 18056 129016 19032
rect 129078 18056 129112 19032
rect 129112 18056 129192 19032
rect 129192 18056 129226 19032
rect 129288 18056 129322 19032
rect 129322 18056 129402 19032
rect 129402 18056 129436 19032
rect 129498 18056 129532 19032
rect 129532 18056 129612 19032
rect 129612 18056 129646 19032
rect 129708 18056 129742 19032
rect 129742 18056 129822 19032
rect 129822 18056 129856 19032
rect 129918 18056 129952 19032
rect 129952 18056 130032 19032
rect 130032 18056 130066 19032
rect 130128 18056 130162 19032
rect 130162 18056 130242 19032
rect 130242 18056 130276 19032
rect 130338 18056 130372 19032
rect 130372 18056 130452 19032
rect 130452 18056 130486 19032
rect 130548 18056 130582 19032
rect 130582 18056 130662 19032
rect 130662 18056 130696 19032
rect 130758 18056 130792 19032
rect 130792 18056 130872 19032
rect 130872 18056 130906 19032
rect 130968 18056 131002 19032
rect 131002 18056 131082 19032
rect 131082 18056 131116 19032
rect 131178 18056 131212 19032
rect 131212 18056 131292 19032
rect 131292 18056 131326 19032
rect 131388 18056 131422 19032
rect 131422 18056 131502 19032
rect 131502 18056 131536 19032
rect 131598 18056 131632 19032
rect 131632 18056 131712 19032
rect 131712 18056 131746 19032
rect 131808 18056 131842 19032
rect 131842 18056 131922 19032
rect 131922 18056 131956 19032
rect 132018 18056 132052 19032
rect 132052 18056 132132 19032
rect 132132 18056 132166 19032
rect 132228 18056 132262 19032
rect 132262 18056 132342 19032
rect 132342 18056 132376 19032
rect 132438 18056 132472 19032
rect 132472 18056 132552 19032
rect 132552 18056 132586 19032
rect 132648 18056 132682 19032
rect 132682 18056 132762 19032
rect 132762 18056 132796 19032
rect 132858 18056 132892 19032
rect 132892 18056 132972 19032
rect 132972 18056 133006 19032
rect 133068 18056 133102 19032
rect 133102 18056 133182 19032
rect 133182 18056 133216 19032
rect 133278 18056 133312 19032
rect 133312 18056 133392 19032
rect 133392 18056 133426 19032
rect 133488 18056 133522 19032
rect 133522 18056 133602 19032
rect 133602 18056 133636 19032
rect 133698 18056 133732 19032
rect 133732 18056 133812 19032
rect 133812 18056 133846 19032
rect 133908 18056 133942 19032
rect 133942 18056 134022 19032
rect 134022 18056 134056 19032
rect 134118 18056 134152 19032
rect 134152 18056 134232 19032
rect 134232 18056 134266 19032
rect 134328 18056 134362 19032
rect 134362 18056 134442 19032
rect 134442 18056 134476 19032
rect 134538 18056 134572 19032
rect 134572 18056 134652 19032
rect 134652 18056 134686 19032
rect 134748 18056 134782 19032
rect 134782 18056 134862 19032
rect 134862 18056 134896 19032
rect 134958 18056 134992 19032
rect 134992 18056 135072 19032
rect 135072 18056 135106 19032
rect 135168 18056 135202 19032
rect 135202 18056 135226 19032
rect 116734 17152 117062 17414
rect 119522 17622 119666 17770
rect 116366 16958 116450 17044
rect 116350 16384 116424 16390
rect 116350 16338 116424 16384
rect 116350 16332 116424 16338
rect 120924 16218 121168 16466
rect 116370 15730 116440 15804
rect 116552 15730 116622 15804
rect 115844 15554 115908 15620
rect 116370 15586 116440 15660
rect 116552 15586 116622 15660
rect 116512 14966 116574 14972
rect 116512 14920 116574 14966
rect 116512 14918 116574 14920
rect 115842 14522 115906 14586
rect 116366 14346 116450 14432
rect 121904 17802 122004 17902
rect 122324 17802 122424 17902
rect 122744 17802 122844 17902
rect 123164 17802 123264 17902
rect 123584 17802 123684 17902
rect 124004 17802 124104 17902
rect 124424 17802 124524 17902
rect 124844 17802 124944 17902
rect 125264 17802 125364 17902
rect 125684 17802 125784 17902
rect 126746 17786 126846 17886
rect 127166 17786 127266 17886
rect 127586 17786 127686 17886
rect 128006 17786 128106 17886
rect 128426 17786 128526 17886
rect 128846 17786 128946 17886
rect 129266 17786 129366 17886
rect 129686 17786 129786 17886
rect 130106 17786 130206 17886
rect 130526 17786 130626 17886
rect 130946 17786 131046 17886
rect 131366 17786 131466 17886
rect 131786 17786 131886 17886
rect 132206 17786 132306 17886
rect 132626 17786 132726 17886
rect 133046 17786 133146 17886
rect 133466 17786 133566 17886
rect 133886 17786 133986 17886
rect 134306 17786 134406 17886
rect 134726 17786 134826 17886
rect 135146 17786 135246 17886
rect 121558 14906 121802 15154
rect 116734 13976 117062 14238
rect 119522 13620 119666 13768
rect 121904 13488 122004 13588
rect 122324 13488 122424 13588
rect 122744 13488 122844 13588
rect 123164 13488 123264 13588
rect 123584 13488 123684 13588
rect 124004 13488 124104 13588
rect 124424 13488 124524 13588
rect 124844 13488 124944 13588
rect 125264 13488 125364 13588
rect 125684 13488 125784 13588
rect 119082 12358 119120 13334
rect 119120 12358 119154 13334
rect 119206 12358 119216 13334
rect 119216 12358 119250 13334
rect 119250 12358 119260 13334
rect 119312 12358 119346 13334
rect 119346 12358 119384 13334
rect 119834 12358 119858 13334
rect 119858 12358 119892 13334
rect 119954 12358 119988 13334
rect 119988 12358 120068 13334
rect 120068 12358 120102 13334
rect 120164 12358 120198 13334
rect 120198 12358 120278 13334
rect 120278 12358 120312 13334
rect 120374 12358 120408 13334
rect 120408 12358 120488 13334
rect 120488 12358 120522 13334
rect 120584 12358 120618 13334
rect 120618 12358 120698 13334
rect 120698 12358 120732 13334
rect 120794 12358 120828 13334
rect 120828 12358 120908 13334
rect 120908 12358 120942 13334
rect 121004 12358 121038 13334
rect 121038 12358 121118 13334
rect 121118 12358 121152 13334
rect 121214 12358 121248 13334
rect 121248 12358 121328 13334
rect 121328 12358 121362 13334
rect 121424 12358 121458 13334
rect 121458 12358 121482 13334
rect 119104 11130 119124 12106
rect 119124 11130 119158 12106
rect 119212 11130 119246 12106
rect 119246 11130 119266 12106
rect 119332 12054 119474 12202
rect 122008 12358 122032 13334
rect 122032 12358 122066 13334
rect 122128 12358 122162 13334
rect 122162 12358 122242 13334
rect 122242 12358 122276 13334
rect 122338 12358 122372 13334
rect 122372 12358 122452 13334
rect 122452 12358 122486 13334
rect 122548 12358 122582 13334
rect 122582 12358 122662 13334
rect 122662 12358 122696 13334
rect 122758 12358 122792 13334
rect 122792 12358 122872 13334
rect 122872 12358 122906 13334
rect 122968 12358 123002 13334
rect 123002 12358 123082 13334
rect 123082 12358 123116 13334
rect 123178 12358 123212 13334
rect 123212 12358 123292 13334
rect 123292 12358 123326 13334
rect 123388 12358 123422 13334
rect 123422 12358 123502 13334
rect 123502 12358 123536 13334
rect 123598 12358 123632 13334
rect 123632 12358 123712 13334
rect 123712 12358 123746 13334
rect 123808 12358 123842 13334
rect 123842 12358 123922 13334
rect 123922 12358 123956 13334
rect 124018 12358 124052 13334
rect 124052 12358 124132 13334
rect 124132 12358 124166 13334
rect 124228 12358 124262 13334
rect 124262 12358 124342 13334
rect 124342 12358 124376 13334
rect 124438 12358 124472 13334
rect 124472 12358 124552 13334
rect 124552 12358 124586 13334
rect 124648 12358 124682 13334
rect 124682 12358 124762 13334
rect 124762 12358 124796 13334
rect 124858 12358 124892 13334
rect 124892 12358 124972 13334
rect 124972 12358 125006 13334
rect 125068 12358 125102 13334
rect 125102 12358 125182 13334
rect 125182 12358 125216 13334
rect 125278 12358 125312 13334
rect 125312 12358 125392 13334
rect 125392 12358 125426 13334
rect 125488 12358 125522 13334
rect 125522 12358 125602 13334
rect 125602 12358 125636 13334
rect 125698 12358 125732 13334
rect 125732 12358 125756 13334
rect 120048 11130 120068 12106
rect 120068 11130 120102 12106
rect 120164 11130 120198 12106
rect 120198 11130 120278 12106
rect 120278 11130 120312 12106
rect 120374 11130 120408 12106
rect 120408 11130 120488 12106
rect 120488 11130 120522 12106
rect 120584 11130 120618 12106
rect 120618 11130 120698 12106
rect 120698 11130 120732 12106
rect 120794 11130 120828 12106
rect 120828 11130 120848 12106
rect 121264 11694 121546 11958
rect 122008 11122 122032 12098
rect 122032 11122 122066 12098
rect 122128 11122 122162 12098
rect 122162 11122 122242 12098
rect 122242 11122 122276 12098
rect 122338 11122 122372 12098
rect 122372 11122 122452 12098
rect 122452 11122 122486 12098
rect 122548 11122 122582 12098
rect 122582 11122 122662 12098
rect 122662 11122 122696 12098
rect 122758 11122 122792 12098
rect 122792 11122 122872 12098
rect 122872 11122 122906 12098
rect 122968 11122 123002 12098
rect 123002 11122 123082 12098
rect 123082 11122 123116 12098
rect 123178 11122 123212 12098
rect 123212 11122 123292 12098
rect 123292 11122 123326 12098
rect 123388 11122 123422 12098
rect 123422 11122 123502 12098
rect 123502 11122 123536 12098
rect 123598 11122 123632 12098
rect 123632 11122 123712 12098
rect 123712 11122 123746 12098
rect 123808 11122 123842 12098
rect 123842 11122 123922 12098
rect 123922 11122 123956 12098
rect 124018 11122 124052 12098
rect 124052 11122 124132 12098
rect 124132 11122 124166 12098
rect 124228 11122 124262 12098
rect 124262 11122 124342 12098
rect 124342 11122 124376 12098
rect 124438 11122 124472 12098
rect 124472 11122 124552 12098
rect 124552 11122 124586 12098
rect 124648 11122 124682 12098
rect 124682 11122 124762 12098
rect 124762 11122 124796 12098
rect 124858 11122 124892 12098
rect 124892 11122 124972 12098
rect 124972 11122 125006 12098
rect 125068 11122 125102 12098
rect 125102 11122 125182 12098
rect 125182 11122 125216 12098
rect 125278 11122 125312 12098
rect 125312 11122 125392 12098
rect 125392 11122 125426 12098
rect 125488 11122 125522 12098
rect 125522 11122 125602 12098
rect 125602 11122 125636 12098
rect 125698 11122 125732 12098
rect 125732 11122 125756 12098
rect 119488 10660 119786 10942
rect 122008 8106 122032 9082
rect 122032 8106 122066 9082
rect 122128 8106 122162 9082
rect 122162 8106 122242 9082
rect 122242 8106 122276 9082
rect 122338 8106 122372 9082
rect 122372 8106 122452 9082
rect 122452 8106 122486 9082
rect 122548 8106 122582 9082
rect 122582 8106 122662 9082
rect 122662 8106 122696 9082
rect 122758 8106 122792 9082
rect 122792 8106 122872 9082
rect 122872 8106 122906 9082
rect 122968 8106 123002 9082
rect 123002 8106 123082 9082
rect 123082 8106 123116 9082
rect 123178 8106 123212 9082
rect 123212 8106 123292 9082
rect 123292 8106 123326 9082
rect 123388 8106 123422 9082
rect 123422 8106 123502 9082
rect 123502 8106 123536 9082
rect 123598 8106 123632 9082
rect 123632 8106 123712 9082
rect 123712 8106 123746 9082
rect 123808 8106 123842 9082
rect 123842 8106 123922 9082
rect 123922 8106 123956 9082
rect 124018 8106 124052 9082
rect 124052 8106 124132 9082
rect 124132 8106 124166 9082
rect 124228 8106 124262 9082
rect 124262 8106 124342 9082
rect 124342 8106 124376 9082
rect 124438 8106 124472 9082
rect 124472 8106 124552 9082
rect 124552 8106 124586 9082
rect 124648 8106 124682 9082
rect 124682 8106 124762 9082
rect 124762 8106 124796 9082
rect 124858 8106 124892 9082
rect 124892 8106 124972 9082
rect 124972 8106 125006 9082
rect 125068 8106 125102 9082
rect 125102 8106 125182 9082
rect 125182 8106 125216 9082
rect 125278 8106 125312 9082
rect 125312 8106 125392 9082
rect 125392 8106 125426 9082
rect 125488 8106 125522 9082
rect 125522 8106 125602 9082
rect 125602 8106 125636 9082
rect 125698 8106 125732 9082
rect 125732 8106 125756 9082
rect 122028 7828 122128 7928
rect 122448 7828 122548 7928
rect 122868 7828 122968 7928
rect 123288 7828 123388 7928
rect 123708 7828 123808 7928
rect 124128 7828 124228 7928
rect 124548 7828 124648 7928
rect 124968 7828 125068 7928
rect 125388 7828 125488 7928
rect 125714 7828 125814 7928
<< metal2 >>
rect 126668 28550 126966 28560
rect 126668 28258 126840 28268
rect 126938 28258 126966 28268
rect 127118 28550 127416 28560
rect 127118 28258 127260 28268
rect 126840 28190 126938 28200
rect 127188 28200 127260 28258
rect 127358 28258 127416 28268
rect 127538 28550 127836 28560
rect 127538 28258 127680 28268
rect 127188 28190 127358 28200
rect 127608 28200 127680 28258
rect 127778 28258 127836 28268
rect 127958 28550 128256 28560
rect 127958 28258 128100 28268
rect 127608 28190 127778 28200
rect 128028 28200 128100 28258
rect 128198 28258 128256 28268
rect 128378 28550 128676 28560
rect 128378 28258 128520 28268
rect 128028 28190 128198 28200
rect 128448 28200 128520 28258
rect 128618 28258 128676 28268
rect 128798 28550 129096 28560
rect 128798 28258 128940 28268
rect 128448 28190 128618 28200
rect 128868 28200 128940 28258
rect 129038 28258 129096 28268
rect 129218 28550 129516 28560
rect 129218 28258 129360 28268
rect 128868 28190 129038 28200
rect 129288 28200 129360 28258
rect 129458 28258 129516 28268
rect 129638 28550 129936 28560
rect 129638 28258 129780 28268
rect 129288 28190 129458 28200
rect 129708 28200 129780 28258
rect 129878 28258 129936 28268
rect 130058 28550 130356 28560
rect 130058 28258 130200 28268
rect 129708 28190 129878 28200
rect 130128 28200 130200 28258
rect 130298 28258 130356 28268
rect 130478 28550 130776 28560
rect 130478 28258 130620 28268
rect 130128 28190 130298 28200
rect 130548 28200 130620 28258
rect 130718 28258 130776 28268
rect 130898 28550 131196 28560
rect 130898 28258 131040 28268
rect 130548 28190 130718 28200
rect 130968 28200 131040 28258
rect 131138 28258 131196 28268
rect 131318 28550 131616 28560
rect 131318 28258 131460 28268
rect 130968 28190 131138 28200
rect 131388 28200 131460 28258
rect 131558 28258 131616 28268
rect 131738 28550 132036 28560
rect 131738 28258 131880 28268
rect 131388 28190 131558 28200
rect 131808 28200 131880 28258
rect 131978 28258 132036 28268
rect 132158 28550 132456 28560
rect 132158 28258 132300 28268
rect 131808 28190 131978 28200
rect 132228 28200 132300 28258
rect 132398 28258 132456 28268
rect 132578 28550 132876 28560
rect 132578 28258 132720 28268
rect 132228 28190 132398 28200
rect 132648 28200 132720 28258
rect 132818 28258 132876 28268
rect 132998 28550 133296 28560
rect 132998 28258 133140 28268
rect 132648 28190 132818 28200
rect 133068 28200 133140 28258
rect 133238 28258 133296 28268
rect 133418 28550 133716 28560
rect 133418 28258 133560 28268
rect 133068 28190 133238 28200
rect 133488 28200 133560 28258
rect 133658 28258 133716 28268
rect 133838 28550 134136 28560
rect 133838 28258 133980 28268
rect 133488 28190 133658 28200
rect 133908 28200 133980 28258
rect 134078 28258 134136 28268
rect 134258 28550 134556 28560
rect 134258 28258 134400 28268
rect 133908 28190 134078 28200
rect 134328 28200 134400 28258
rect 134498 28258 134556 28268
rect 134678 28550 134976 28560
rect 134678 28258 134820 28268
rect 134328 28190 134498 28200
rect 134748 28200 134820 28258
rect 134918 28258 134976 28268
rect 135098 28550 135396 28560
rect 135098 28258 135168 28268
rect 134748 28190 134918 28200
rect 135266 28258 135396 28268
rect 135168 28190 135266 28200
rect 126858 27968 126916 28190
rect 126858 26750 126916 26992
rect 126858 25764 126916 25774
rect 126978 27968 127126 27978
rect 126978 26750 127126 26992
rect 126978 25636 127126 25774
rect 127188 27968 127336 28190
rect 127188 26750 127336 26992
rect 127188 25764 127336 25774
rect 127398 27968 127546 27978
rect 127398 26750 127546 26992
rect 127398 25636 127546 25774
rect 127608 27968 127756 28190
rect 127608 26750 127756 26992
rect 127608 25764 127756 25774
rect 127818 27968 127966 27978
rect 127818 26750 127966 26992
rect 127818 25636 127966 25774
rect 128028 27968 128176 28190
rect 128028 26750 128176 26992
rect 128028 25764 128176 25774
rect 128238 27968 128386 27978
rect 128238 26750 128386 26992
rect 128238 25636 128386 25774
rect 128448 27968 128596 28190
rect 128448 26750 128596 26992
rect 128448 25764 128596 25774
rect 128658 27968 128806 27978
rect 128658 26750 128806 26992
rect 128658 25636 128806 25774
rect 128868 27968 129016 28190
rect 128868 26750 129016 26992
rect 128868 25764 129016 25774
rect 129078 27968 129226 27978
rect 129078 26750 129226 26992
rect 129078 25636 129226 25774
rect 129288 27968 129436 28190
rect 129288 26750 129436 26992
rect 129288 25764 129436 25774
rect 129498 27968 129646 27978
rect 129498 26750 129646 26992
rect 129498 25636 129646 25774
rect 129708 27968 129856 28190
rect 129708 26750 129856 26992
rect 129708 25764 129856 25774
rect 129918 27968 130066 27978
rect 129918 26750 130066 26992
rect 129918 25636 130066 25774
rect 130128 27968 130276 28190
rect 130128 26750 130276 26992
rect 130128 25764 130276 25774
rect 130338 27968 130486 27978
rect 130338 26750 130486 26992
rect 130338 25636 130486 25774
rect 130548 27968 130696 28190
rect 130548 26750 130696 26992
rect 130548 25764 130696 25774
rect 130758 27968 130906 27978
rect 130758 26750 130906 26992
rect 130758 25636 130906 25774
rect 130968 27968 131116 28190
rect 130968 26750 131116 26992
rect 130968 25764 131116 25774
rect 131178 27968 131326 27978
rect 131178 26750 131326 26992
rect 131178 25636 131326 25774
rect 131388 27968 131536 28190
rect 131388 26750 131536 26992
rect 131388 25764 131536 25774
rect 131598 27968 131746 27978
rect 131598 26750 131746 26992
rect 131598 25636 131746 25774
rect 131808 27968 131956 28190
rect 131808 26750 131956 26992
rect 131808 25764 131956 25774
rect 132018 27968 132166 27978
rect 132018 26750 132166 26992
rect 132018 25636 132166 25774
rect 132228 27968 132376 28190
rect 132228 26750 132376 26992
rect 132228 25764 132376 25774
rect 132438 27968 132586 27978
rect 132438 26750 132586 26992
rect 132438 25636 132586 25774
rect 132648 27968 132796 28190
rect 132648 26750 132796 26992
rect 132648 25764 132796 25774
rect 132858 27968 133006 27978
rect 132858 26750 133006 26992
rect 132858 25636 133006 25774
rect 133068 27968 133216 28190
rect 133068 26750 133216 26992
rect 133068 25764 133216 25774
rect 133278 27968 133426 27978
rect 133278 26750 133426 26992
rect 133278 25636 133426 25774
rect 133488 27968 133636 28190
rect 133488 26750 133636 26992
rect 133488 25764 133636 25774
rect 133698 27968 133846 27978
rect 133698 26750 133846 26992
rect 133698 25636 133846 25774
rect 133908 27968 134056 28190
rect 133908 26750 134056 26992
rect 133908 25764 134056 25774
rect 134118 27968 134266 27978
rect 134118 26750 134266 26992
rect 134118 25636 134266 25774
rect 134328 27968 134476 28190
rect 134328 26750 134476 26992
rect 134328 25764 134476 25774
rect 134538 27968 134686 27978
rect 134538 26750 134686 26992
rect 134538 25636 134686 25774
rect 134748 27968 134896 28190
rect 134748 26750 134896 26992
rect 134748 25764 134896 25774
rect 134958 27968 135106 27978
rect 134958 26750 135106 26992
rect 134958 25636 135106 25774
rect 135168 27968 135226 28190
rect 135168 26750 135226 26992
rect 135168 25764 135226 25774
rect 126978 22938 135106 25636
rect 126858 22740 126916 22750
rect 121830 22372 122128 22382
rect 121830 22080 122028 22090
rect 122008 22062 122028 22080
rect 122250 22372 122548 22382
rect 122250 22080 122448 22090
rect 122008 22052 122128 22062
rect 122338 22062 122448 22080
rect 122670 22372 122968 22382
rect 122670 22080 122868 22090
rect 122338 22056 122548 22062
rect 122758 22062 122868 22080
rect 123090 22372 123388 22382
rect 123090 22080 123288 22090
rect 122758 22056 122968 22062
rect 123178 22062 123288 22080
rect 123510 22372 123808 22382
rect 123510 22080 123708 22090
rect 123178 22056 123388 22062
rect 123598 22062 123708 22080
rect 123930 22372 124228 22382
rect 123930 22080 124128 22090
rect 123598 22056 123808 22062
rect 124018 22062 124128 22080
rect 124350 22372 124648 22382
rect 124350 22080 124548 22090
rect 124018 22056 124228 22062
rect 124438 22062 124548 22080
rect 124770 22372 125068 22382
rect 124770 22080 124968 22090
rect 124438 22056 124648 22062
rect 124858 22062 124968 22080
rect 125190 22372 125488 22382
rect 125190 22080 125388 22090
rect 124858 22056 125068 22062
rect 125278 22062 125388 22080
rect 125610 22372 125908 22382
rect 125610 22080 125714 22090
rect 125278 22056 125488 22062
rect 125698 22062 125714 22080
rect 125814 22080 125908 22090
rect 122008 21884 122066 22052
rect 122008 20898 122066 20908
rect 122128 21884 122276 21894
rect 122128 20782 122276 20908
rect 122338 21884 122486 22056
rect 122338 20898 122486 20908
rect 122548 21884 122696 21894
rect 122548 20782 122696 20908
rect 122758 21884 122906 22056
rect 122758 20898 122906 20908
rect 122968 21884 123116 21894
rect 122968 20782 123116 20908
rect 123178 21884 123326 22056
rect 123178 20898 123326 20908
rect 123388 21884 123536 21894
rect 123388 20782 123536 20908
rect 123598 21884 123746 22056
rect 123598 20898 123746 20908
rect 123808 21884 123956 21894
rect 123808 20782 123956 20908
rect 124018 21884 124166 22056
rect 124018 20898 124166 20908
rect 124228 21884 124376 21894
rect 124228 20782 124376 20908
rect 124438 21884 124586 22056
rect 124438 20898 124586 20908
rect 124648 21884 124796 21894
rect 124648 20782 124796 20908
rect 124858 21884 125006 22056
rect 124858 20898 125006 20908
rect 125068 21884 125216 21894
rect 125068 20782 125216 20908
rect 125278 21884 125426 22056
rect 125698 22052 125814 22062
rect 125278 20898 125426 20908
rect 125488 21884 125636 21894
rect 125488 20782 125636 20908
rect 125698 21884 125756 22052
rect 126858 21504 126916 21764
rect 125698 20898 125756 20908
rect 125864 20928 126474 20938
rect 119028 20730 119326 20740
rect 119028 20438 119326 20448
rect 119488 20730 119786 20740
rect 119488 20438 119786 20448
rect 119888 20730 120186 20740
rect 119888 20438 120186 20448
rect 120308 20730 120606 20740
rect 120308 20438 120606 20448
rect 120728 20730 121026 20740
rect 120728 20438 121026 20448
rect 119104 20260 119158 20438
rect 119104 19274 119158 19284
rect 119206 20260 119266 20270
rect 119206 19284 119212 20260
rect 120048 20260 120102 20438
rect 119206 19274 119266 19284
rect 119332 19336 119474 19346
rect 119206 19204 119332 19274
rect 119082 19032 119154 19042
rect 119082 17944 119154 18056
rect 119206 19032 119260 19204
rect 120048 19274 120102 19284
rect 120164 20260 120312 20270
rect 120164 19220 120312 19284
rect 120374 20260 120522 20438
rect 120374 19274 120522 19284
rect 120584 20260 120732 20270
rect 120584 19220 120732 19284
rect 120794 20260 120848 20438
rect 120888 20436 120942 20438
rect 122128 20402 125864 20782
rect 122008 20268 122066 20278
rect 121264 19696 121546 19706
rect 121264 19422 121546 19432
rect 120794 19274 120848 19284
rect 121328 19220 121482 19422
rect 119332 19178 119474 19188
rect 119834 19100 121482 19220
rect 119206 18046 119260 18056
rect 119312 19032 119384 19042
rect 119312 17944 119384 18056
rect 119834 19032 119892 19100
rect 119834 18046 119892 18056
rect 119954 19032 120102 19042
rect 119030 17934 119424 17944
rect 119954 17902 120102 18056
rect 120164 19032 120312 19100
rect 120164 18046 120312 18056
rect 120374 19032 120522 19042
rect 120374 17902 120522 18056
rect 120584 19032 120732 19100
rect 120584 18046 120732 18056
rect 120794 19032 120942 19042
rect 120794 17902 120942 18056
rect 121004 19032 121152 19100
rect 121004 18046 121152 18056
rect 121214 19032 121362 19042
rect 121214 17902 121362 18056
rect 121424 19032 121482 19100
rect 121424 18046 121482 18056
rect 122008 19032 122066 19292
rect 122008 17912 122066 18056
rect 122128 20268 122276 20402
rect 122128 19032 122276 19292
rect 122128 18046 122276 18056
rect 122338 20268 122486 20278
rect 122338 19032 122486 19292
rect 122338 17912 122486 18056
rect 122548 20268 122696 20402
rect 122548 19032 122696 19292
rect 122548 18046 122696 18056
rect 122758 20268 122906 20278
rect 122758 19032 122906 19292
rect 121904 17902 122066 17912
rect 122324 17902 122486 17912
rect 122758 17908 122906 18056
rect 122968 20268 123116 20402
rect 122968 19032 123116 19292
rect 122968 18046 123116 18056
rect 123178 20268 123326 20278
rect 123178 19032 123326 19292
rect 123178 17908 123326 18056
rect 123388 20268 123536 20402
rect 123388 19032 123536 19292
rect 123388 18046 123536 18056
rect 123598 20268 123746 20278
rect 123598 19032 123746 19292
rect 123598 17908 123746 18056
rect 123808 20268 123956 20402
rect 123808 19032 123956 19292
rect 123808 18046 123956 18056
rect 124018 20268 124166 20278
rect 124018 19032 124166 19292
rect 124018 17908 124166 18056
rect 124228 20268 124376 20402
rect 124228 19032 124376 19292
rect 124228 18046 124376 18056
rect 124438 20268 124586 20278
rect 124438 19032 124586 19292
rect 124438 17908 124586 18056
rect 124648 20268 124796 20402
rect 124648 19032 124796 19292
rect 124648 18046 124796 18056
rect 124858 20268 125006 20278
rect 124858 19032 125006 19292
rect 124858 17908 125006 18056
rect 125068 20268 125216 20402
rect 125068 19032 125216 19292
rect 125068 18046 125216 18056
rect 125278 20268 125426 20278
rect 125278 19032 125426 19292
rect 125278 17908 125426 18056
rect 125488 20268 125636 20402
rect 125864 20300 126474 20310
rect 125488 19032 125636 19292
rect 125488 18046 125636 18056
rect 125698 20268 125756 20278
rect 125698 19032 125756 19292
rect 125698 17908 125756 18056
rect 126858 20268 126916 20528
rect 126858 19032 126916 19292
rect 122744 17902 122906 17908
rect 123164 17902 123326 17908
rect 123584 17902 123746 17908
rect 124004 17902 124166 17908
rect 124424 17902 124586 17908
rect 124844 17902 125006 17908
rect 125264 17902 125426 17908
rect 125684 17902 125796 17908
rect 126858 17902 126916 18056
rect 126978 22740 127126 22938
rect 126978 21504 127126 21764
rect 126978 20268 127126 20528
rect 126978 19032 127126 19292
rect 126978 18046 127126 18056
rect 127188 22740 127336 22750
rect 127188 21504 127336 21764
rect 127188 20268 127336 20528
rect 127188 19032 127336 19292
rect 127188 17902 127336 18056
rect 127398 22740 127546 22938
rect 127398 21504 127546 21764
rect 127398 20268 127546 20528
rect 127398 19032 127546 19292
rect 127398 18046 127546 18056
rect 127608 22740 127756 22750
rect 127608 21504 127756 21764
rect 127608 20268 127756 20528
rect 127608 19032 127756 19292
rect 127608 17902 127756 18056
rect 127818 22740 127966 22938
rect 127818 21504 127966 21764
rect 127818 20268 127966 20528
rect 127818 19032 127966 19292
rect 127818 18046 127966 18056
rect 128028 22740 128176 22750
rect 128028 21504 128176 21764
rect 128028 20268 128176 20528
rect 128028 19032 128176 19292
rect 128028 17902 128176 18056
rect 128238 22740 128386 22938
rect 128238 21504 128386 21764
rect 128238 20268 128386 20528
rect 128238 19032 128386 19292
rect 128238 18046 128386 18056
rect 128448 22740 128596 22750
rect 128448 21504 128596 21764
rect 128448 20268 128596 20528
rect 128448 19032 128596 19292
rect 128448 17902 128596 18056
rect 128658 22740 128806 22938
rect 128658 21504 128806 21764
rect 128658 20268 128806 20528
rect 128658 19032 128806 19292
rect 128658 18046 128806 18056
rect 128868 22740 129016 22750
rect 128868 21504 129016 21764
rect 128868 20268 129016 20528
rect 128868 19032 129016 19292
rect 128868 17902 129016 18056
rect 129078 22740 129226 22938
rect 129078 21504 129226 21764
rect 129078 20268 129226 20528
rect 129078 19032 129226 19292
rect 129078 18046 129226 18056
rect 129288 22740 129436 22750
rect 129288 21504 129436 21764
rect 129288 20268 129436 20528
rect 129288 19032 129436 19292
rect 129288 17902 129436 18056
rect 129498 22740 129646 22938
rect 129498 21504 129646 21764
rect 129498 20268 129646 20528
rect 129498 19032 129646 19292
rect 129498 18046 129646 18056
rect 129708 22740 129856 22750
rect 129708 21504 129856 21764
rect 129708 20268 129856 20528
rect 129708 19032 129856 19292
rect 129708 17902 129856 18056
rect 129918 22740 130066 22938
rect 129918 21504 130066 21764
rect 129918 20268 130066 20528
rect 129918 19032 130066 19292
rect 129918 18046 130066 18056
rect 130128 22740 130276 22750
rect 130128 21504 130276 21764
rect 130128 20268 130276 20528
rect 130128 19032 130276 19292
rect 130128 17902 130276 18056
rect 130338 22740 130486 22938
rect 130338 21504 130486 21764
rect 130338 20268 130486 20528
rect 130338 19032 130486 19292
rect 130338 18046 130486 18056
rect 130548 22740 130696 22750
rect 130548 21504 130696 21764
rect 130548 20268 130696 20528
rect 130548 19032 130696 19292
rect 130548 17902 130696 18056
rect 130758 22740 130906 22938
rect 130758 21504 130906 21764
rect 130758 20268 130906 20528
rect 130758 19032 130906 19292
rect 130758 18046 130906 18056
rect 130968 22740 131116 22750
rect 130968 21504 131116 21764
rect 130968 20268 131116 20528
rect 130968 19032 131116 19292
rect 130968 17902 131116 18056
rect 131178 22740 131326 22938
rect 131178 21504 131326 21764
rect 131178 20268 131326 20528
rect 131178 19032 131326 19292
rect 131178 18046 131326 18056
rect 131388 22740 131536 22750
rect 131388 21504 131536 21764
rect 131388 20268 131536 20528
rect 131388 19032 131536 19292
rect 131388 17902 131536 18056
rect 131598 22740 131746 22938
rect 131598 21504 131746 21764
rect 131598 20268 131746 20528
rect 131598 19032 131746 19292
rect 131598 18046 131746 18056
rect 131808 22740 131956 22750
rect 131808 21504 131956 21764
rect 131808 20268 131956 20528
rect 131808 19032 131956 19292
rect 131808 17902 131956 18056
rect 132018 22740 132166 22938
rect 132018 21504 132166 21764
rect 132018 20268 132166 20528
rect 132018 19032 132166 19292
rect 132018 18046 132166 18056
rect 132228 22740 132376 22750
rect 132228 21504 132376 21764
rect 132228 20268 132376 20528
rect 132228 19032 132376 19292
rect 132228 17902 132376 18056
rect 132438 22740 132586 22938
rect 132438 21504 132586 21764
rect 132438 20268 132586 20528
rect 132438 19032 132586 19292
rect 132438 18046 132586 18056
rect 132648 22740 132796 22750
rect 132648 21504 132796 21764
rect 132648 20268 132796 20528
rect 132648 19032 132796 19292
rect 132648 17902 132796 18056
rect 132858 22740 133006 22938
rect 132858 21504 133006 21764
rect 132858 20268 133006 20528
rect 132858 19032 133006 19292
rect 132858 18046 133006 18056
rect 133068 22740 133216 22750
rect 133068 21504 133216 21764
rect 133068 20268 133216 20528
rect 133068 19032 133216 19292
rect 133068 17902 133216 18056
rect 133278 22740 133426 22938
rect 133278 21504 133426 21764
rect 133278 20268 133426 20528
rect 133278 19032 133426 19292
rect 133278 18046 133426 18056
rect 133488 22740 133636 22750
rect 133488 21504 133636 21764
rect 133488 20268 133636 20528
rect 133488 19032 133636 19292
rect 133488 17902 133636 18056
rect 133698 22740 133846 22938
rect 133698 21504 133846 21764
rect 133698 20268 133846 20528
rect 133698 19032 133846 19292
rect 133698 18046 133846 18056
rect 133908 22740 134056 22750
rect 133908 21504 134056 21764
rect 133908 20268 134056 20528
rect 133908 19032 134056 19292
rect 133908 17902 134056 18056
rect 134118 22740 134266 22938
rect 134118 21504 134266 21764
rect 134118 20268 134266 20528
rect 134118 19032 134266 19292
rect 134118 18046 134266 18056
rect 134328 22740 134476 22750
rect 134328 21504 134476 21764
rect 134328 20268 134476 20528
rect 134328 19032 134476 19292
rect 134328 17902 134476 18056
rect 134538 22740 134686 22938
rect 134538 21504 134686 21764
rect 134538 20268 134686 20528
rect 134538 19032 134686 19292
rect 134538 18046 134686 18056
rect 134748 22740 134896 22750
rect 134748 21504 134896 21764
rect 134748 20268 134896 20528
rect 134748 19032 134896 19292
rect 134748 17902 134896 18056
rect 134958 22740 135106 22938
rect 134958 21504 135106 21764
rect 134958 20268 135106 20528
rect 134958 19032 135106 19292
rect 134958 18046 135106 18056
rect 135168 22740 135226 22750
rect 135168 21504 135226 21764
rect 135168 20268 135226 20528
rect 135168 19032 135226 19292
rect 135168 17902 135226 18056
rect 119876 17892 120174 17902
rect 119030 17760 119424 17770
rect 119522 17770 119666 17780
rect 119522 17612 119666 17622
rect 119876 17600 120174 17610
rect 120296 17892 120594 17902
rect 120296 17600 120594 17610
rect 120716 17892 121014 17902
rect 120716 17600 121014 17610
rect 121136 17892 121434 17902
rect 121136 17600 121434 17610
rect 121836 17892 121904 17902
rect 122004 17892 122134 17902
rect 121836 17600 122134 17610
rect 122266 17892 122324 17902
rect 122424 17892 122564 17902
rect 122266 17600 122564 17610
rect 122686 17892 122744 17902
rect 122844 17892 122984 17902
rect 122686 17600 122984 17610
rect 123106 17892 123164 17902
rect 123264 17892 123404 17902
rect 123106 17600 123404 17610
rect 123526 17892 123584 17902
rect 123684 17892 123824 17902
rect 123526 17600 123824 17610
rect 123946 17892 124004 17902
rect 124104 17892 124244 17902
rect 123946 17600 124244 17610
rect 124366 17892 124424 17902
rect 124524 17892 124664 17902
rect 124366 17600 124664 17610
rect 124786 17892 124844 17902
rect 124944 17892 125084 17902
rect 124786 17600 125084 17610
rect 125206 17892 125264 17902
rect 125364 17892 125504 17902
rect 125206 17600 125504 17610
rect 125626 17892 125684 17902
rect 125784 17892 125924 17902
rect 125626 17600 125924 17610
rect 126666 17892 126964 17902
rect 126666 17600 126964 17610
rect 127116 17892 127414 17902
rect 127116 17600 127414 17610
rect 127536 17892 127834 17902
rect 127536 17600 127834 17610
rect 127956 17892 128254 17902
rect 127956 17600 128254 17610
rect 128376 17892 128674 17902
rect 128376 17600 128674 17610
rect 128796 17892 129094 17902
rect 128796 17600 129094 17610
rect 129216 17892 129514 17902
rect 129216 17600 129514 17610
rect 129636 17892 129934 17902
rect 129636 17600 129934 17610
rect 130056 17892 130354 17902
rect 130056 17600 130354 17610
rect 130476 17892 130774 17902
rect 130476 17600 130774 17610
rect 130896 17892 131194 17902
rect 130896 17600 131194 17610
rect 131316 17892 131614 17902
rect 131316 17600 131614 17610
rect 131736 17892 132034 17902
rect 131736 17600 132034 17610
rect 132156 17892 132454 17902
rect 132156 17600 132454 17610
rect 132576 17892 132874 17902
rect 132576 17600 132874 17610
rect 132996 17892 133294 17902
rect 132996 17600 133294 17610
rect 133416 17892 133714 17902
rect 133416 17600 133714 17610
rect 133836 17892 134134 17902
rect 133836 17600 134134 17610
rect 134256 17892 134554 17902
rect 134256 17600 134554 17610
rect 134676 17892 134974 17902
rect 134676 17600 134974 17610
rect 135096 17892 135394 17902
rect 135096 17600 135394 17610
rect 116734 17414 117062 17424
rect 116734 17142 117062 17152
rect 116366 17044 116450 17054
rect 116366 16948 116450 16958
rect 120924 16466 121168 16476
rect 116350 16390 120924 16400
rect 116424 16332 120924 16390
rect 116350 16322 120924 16332
rect 120924 16208 121168 16218
rect 116364 15810 116448 15820
rect 116364 15714 116448 15724
rect 116546 15810 116630 15820
rect 116546 15714 116630 15724
rect 116364 15666 116448 15676
rect 115838 15626 115920 15636
rect 116364 15570 116448 15580
rect 116546 15666 116630 15676
rect 116546 15570 116630 15580
rect 115838 15532 115920 15542
rect 121558 15154 121802 15164
rect 116512 14972 121558 14984
rect 116574 14918 121558 14972
rect 116512 14906 121558 14918
rect 121558 14896 121802 14906
rect 115838 14594 115914 14604
rect 115838 14508 115914 14518
rect 116366 14432 116450 14442
rect 116366 14336 116450 14346
rect 116734 14238 117062 14248
rect 116734 13966 117062 13976
rect 119876 13780 120174 13790
rect 119522 13768 119666 13778
rect 119030 13620 119424 13630
rect 119522 13610 119666 13620
rect 119876 13488 120174 13498
rect 120296 13780 120594 13790
rect 120296 13488 120594 13498
rect 120716 13780 121014 13790
rect 120716 13488 121014 13498
rect 121136 13780 121434 13790
rect 121136 13488 121434 13498
rect 121836 13780 122134 13790
rect 121836 13488 121904 13498
rect 122004 13488 122134 13498
rect 122266 13780 122564 13790
rect 122266 13488 122324 13498
rect 122424 13488 122564 13498
rect 122686 13780 122984 13790
rect 122686 13488 122744 13498
rect 122844 13488 122984 13498
rect 123106 13780 123404 13790
rect 123106 13488 123164 13498
rect 123264 13488 123404 13498
rect 123526 13780 123824 13790
rect 123526 13488 123584 13498
rect 123684 13488 123824 13498
rect 123946 13780 124244 13790
rect 123946 13488 124004 13498
rect 124104 13488 124244 13498
rect 124366 13780 124664 13790
rect 124366 13488 124424 13498
rect 124524 13488 124664 13498
rect 124786 13780 125084 13790
rect 124786 13488 124844 13498
rect 124944 13488 125084 13498
rect 125206 13780 125504 13790
rect 125206 13488 125264 13498
rect 125364 13488 125504 13498
rect 125626 13780 125924 13790
rect 125626 13488 125684 13498
rect 125784 13488 125924 13498
rect 119030 13446 119424 13456
rect 119082 13334 119154 13446
rect 119082 12348 119154 12358
rect 119206 13334 119260 13344
rect 119206 12186 119260 12358
rect 119312 13334 119384 13446
rect 119312 12348 119384 12358
rect 119834 13334 119892 13344
rect 119834 12290 119892 12358
rect 119954 13334 120102 13488
rect 119954 12348 120102 12358
rect 120164 13334 120312 13344
rect 120164 12290 120312 12358
rect 120374 13334 120522 13488
rect 120374 12348 120522 12358
rect 120584 13334 120732 13344
rect 120584 12290 120732 12358
rect 120794 13334 120942 13488
rect 120794 12348 120942 12358
rect 121004 13334 121152 13344
rect 121004 12290 121152 12358
rect 121214 13334 121362 13488
rect 121904 13478 122066 13488
rect 122324 13478 122486 13488
rect 122744 13482 122906 13488
rect 123164 13482 123326 13488
rect 123584 13482 123746 13488
rect 124004 13482 124166 13488
rect 124424 13482 124586 13488
rect 124844 13482 125006 13488
rect 125264 13482 125426 13488
rect 125684 13482 125796 13488
rect 121214 12348 121362 12358
rect 121424 13334 121482 13344
rect 121424 12290 121482 12358
rect 119332 12202 119474 12212
rect 119206 12116 119332 12186
rect 119104 12106 119158 12116
rect 119104 10952 119158 11130
rect 119206 12106 119266 12116
rect 119206 11130 119212 12106
rect 119834 12170 121482 12290
rect 119332 12044 119474 12054
rect 120048 12106 120102 12116
rect 119206 11120 119266 11130
rect 120048 10952 120102 11130
rect 120164 12106 120312 12170
rect 120164 11120 120312 11130
rect 120374 12106 120522 12116
rect 120374 10952 120522 11130
rect 120584 12106 120732 12170
rect 120584 11120 120732 11130
rect 120794 12106 120848 12116
rect 121328 11968 121482 12170
rect 122008 13334 122066 13478
rect 122008 12098 122066 12358
rect 121264 11958 121546 11968
rect 121264 11684 121546 11694
rect 120794 10952 120848 11130
rect 122008 11112 122066 11122
rect 122128 13334 122276 13344
rect 122128 12098 122276 12358
rect 122128 10988 122276 11122
rect 122338 13334 122486 13478
rect 122338 12098 122486 12358
rect 122338 11112 122486 11122
rect 122548 13334 122696 13344
rect 122548 12098 122696 12358
rect 122548 10988 122696 11122
rect 122758 13334 122906 13482
rect 122758 12098 122906 12358
rect 122758 11112 122906 11122
rect 122968 13334 123116 13344
rect 122968 12098 123116 12358
rect 122968 10988 123116 11122
rect 123178 13334 123326 13482
rect 123178 12098 123326 12358
rect 123178 11112 123326 11122
rect 123388 13334 123536 13344
rect 123388 12098 123536 12358
rect 123388 10988 123536 11122
rect 123598 13334 123746 13482
rect 123598 12098 123746 12358
rect 123598 11112 123746 11122
rect 123808 13334 123956 13344
rect 123808 12098 123956 12358
rect 123808 10988 123956 11122
rect 124018 13334 124166 13482
rect 124018 12098 124166 12358
rect 124018 11112 124166 11122
rect 124228 13334 124376 13344
rect 124228 12098 124376 12358
rect 124228 10988 124376 11122
rect 124438 13334 124586 13482
rect 124438 12098 124586 12358
rect 124438 11112 124586 11122
rect 124648 13334 124796 13344
rect 124648 12098 124796 12358
rect 124648 10988 124796 11122
rect 124858 13334 125006 13482
rect 124858 12098 125006 12358
rect 124858 11112 125006 11122
rect 125068 13334 125216 13344
rect 125068 12098 125216 12358
rect 125068 10988 125216 11122
rect 125278 13334 125426 13482
rect 125278 12098 125426 12358
rect 125278 11112 125426 11122
rect 125488 13334 125636 13344
rect 125488 12098 125636 12358
rect 125488 10988 125636 11122
rect 125698 13334 125756 13482
rect 125698 12098 125756 12358
rect 125698 11112 125756 11122
rect 120888 10952 120942 10954
rect 119028 10942 119326 10952
rect 119028 10650 119326 10660
rect 119488 10942 119786 10952
rect 119488 10650 119786 10660
rect 119888 10942 120186 10952
rect 119888 10650 120186 10660
rect 120308 10942 120606 10952
rect 120308 10650 120606 10660
rect 120728 10942 121026 10952
rect 120728 10650 121026 10660
rect 122128 9208 125852 10988
rect 122008 9082 122066 9092
rect 122008 7938 122066 8106
rect 122128 9082 122276 9208
rect 122128 8096 122276 8106
rect 122338 9082 122486 9092
rect 122008 7928 122128 7938
rect 122008 7910 122028 7928
rect 121830 7900 122028 7910
rect 122338 7934 122486 8106
rect 122548 9082 122696 9208
rect 122548 8096 122696 8106
rect 122758 9082 122906 9092
rect 122758 7934 122906 8106
rect 122968 9082 123116 9208
rect 122968 8096 123116 8106
rect 123178 9082 123326 9092
rect 123178 7934 123326 8106
rect 123388 9082 123536 9208
rect 123388 8096 123536 8106
rect 123598 9082 123746 9092
rect 123598 7934 123746 8106
rect 123808 9082 123956 9208
rect 123808 8096 123956 8106
rect 124018 9082 124166 9092
rect 124018 7934 124166 8106
rect 124228 9082 124376 9208
rect 124228 8096 124376 8106
rect 124438 9082 124586 9092
rect 124438 7934 124586 8106
rect 124648 9082 124796 9208
rect 124648 8096 124796 8106
rect 124858 9082 125006 9092
rect 124858 7934 125006 8106
rect 125068 9082 125216 9208
rect 125068 8096 125216 8106
rect 125278 9082 125426 9092
rect 125278 7934 125426 8106
rect 125488 9082 125636 9208
rect 125488 8096 125636 8106
rect 125698 9082 125756 9092
rect 125698 7938 125756 8106
rect 122338 7928 122548 7934
rect 122338 7910 122448 7928
rect 121830 7608 122128 7618
rect 122250 7900 122448 7910
rect 122758 7928 122968 7934
rect 122758 7910 122868 7928
rect 122250 7608 122548 7618
rect 122670 7900 122868 7910
rect 123178 7928 123388 7934
rect 123178 7910 123288 7928
rect 122670 7608 122968 7618
rect 123090 7900 123288 7910
rect 123598 7928 123808 7934
rect 123598 7910 123708 7928
rect 123090 7608 123388 7618
rect 123510 7900 123708 7910
rect 124018 7928 124228 7934
rect 124018 7910 124128 7928
rect 123510 7608 123808 7618
rect 123930 7900 124128 7910
rect 124438 7928 124648 7934
rect 124438 7910 124548 7928
rect 123930 7608 124228 7618
rect 124350 7900 124548 7910
rect 124858 7928 125068 7934
rect 124858 7910 124968 7928
rect 124350 7608 124648 7618
rect 124770 7900 124968 7910
rect 125278 7928 125488 7934
rect 125278 7910 125388 7928
rect 124770 7608 125068 7618
rect 125190 7900 125388 7910
rect 125698 7928 125814 7938
rect 125698 7910 125714 7928
rect 125190 7608 125488 7618
rect 125610 7900 125714 7910
rect 125814 7900 125908 7910
rect 125610 7608 125908 7618
<< via2 >>
rect 126668 28304 126966 28550
rect 126668 28268 126840 28304
rect 126840 28268 126938 28304
rect 126938 28268 126966 28304
rect 127118 28304 127416 28550
rect 127118 28268 127260 28304
rect 127260 28268 127358 28304
rect 127358 28268 127416 28304
rect 127538 28304 127836 28550
rect 127538 28268 127680 28304
rect 127680 28268 127778 28304
rect 127778 28268 127836 28304
rect 127958 28304 128256 28550
rect 127958 28268 128100 28304
rect 128100 28268 128198 28304
rect 128198 28268 128256 28304
rect 128378 28304 128676 28550
rect 128378 28268 128520 28304
rect 128520 28268 128618 28304
rect 128618 28268 128676 28304
rect 128798 28304 129096 28550
rect 128798 28268 128940 28304
rect 128940 28268 129038 28304
rect 129038 28268 129096 28304
rect 129218 28304 129516 28550
rect 129218 28268 129360 28304
rect 129360 28268 129458 28304
rect 129458 28268 129516 28304
rect 129638 28304 129936 28550
rect 129638 28268 129780 28304
rect 129780 28268 129878 28304
rect 129878 28268 129936 28304
rect 130058 28304 130356 28550
rect 130058 28268 130200 28304
rect 130200 28268 130298 28304
rect 130298 28268 130356 28304
rect 130478 28304 130776 28550
rect 130478 28268 130620 28304
rect 130620 28268 130718 28304
rect 130718 28268 130776 28304
rect 130898 28304 131196 28550
rect 130898 28268 131040 28304
rect 131040 28268 131138 28304
rect 131138 28268 131196 28304
rect 131318 28304 131616 28550
rect 131318 28268 131460 28304
rect 131460 28268 131558 28304
rect 131558 28268 131616 28304
rect 131738 28304 132036 28550
rect 131738 28268 131880 28304
rect 131880 28268 131978 28304
rect 131978 28268 132036 28304
rect 132158 28304 132456 28550
rect 132158 28268 132300 28304
rect 132300 28268 132398 28304
rect 132398 28268 132456 28304
rect 132578 28304 132876 28550
rect 132578 28268 132720 28304
rect 132720 28268 132818 28304
rect 132818 28268 132876 28304
rect 132998 28304 133296 28550
rect 132998 28268 133140 28304
rect 133140 28268 133238 28304
rect 133238 28268 133296 28304
rect 133418 28304 133716 28550
rect 133418 28268 133560 28304
rect 133560 28268 133658 28304
rect 133658 28268 133716 28304
rect 133838 28304 134136 28550
rect 133838 28268 133980 28304
rect 133980 28268 134078 28304
rect 134078 28268 134136 28304
rect 134258 28304 134556 28550
rect 134258 28268 134400 28304
rect 134400 28268 134498 28304
rect 134498 28268 134556 28304
rect 134678 28304 134976 28550
rect 134678 28268 134820 28304
rect 134820 28268 134918 28304
rect 134918 28268 134976 28304
rect 135098 28304 135396 28550
rect 135098 28268 135168 28304
rect 135168 28268 135266 28304
rect 135266 28268 135396 28304
rect 121830 22162 122128 22372
rect 121830 22090 122028 22162
rect 122028 22090 122128 22162
rect 122250 22162 122548 22372
rect 122250 22090 122448 22162
rect 122448 22090 122548 22162
rect 122670 22162 122968 22372
rect 122670 22090 122868 22162
rect 122868 22090 122968 22162
rect 123090 22162 123388 22372
rect 123090 22090 123288 22162
rect 123288 22090 123388 22162
rect 123510 22162 123808 22372
rect 123510 22090 123708 22162
rect 123708 22090 123808 22162
rect 123930 22162 124228 22372
rect 123930 22090 124128 22162
rect 124128 22090 124228 22162
rect 124350 22162 124648 22372
rect 124350 22090 124548 22162
rect 124548 22090 124648 22162
rect 124770 22162 125068 22372
rect 124770 22090 124968 22162
rect 124968 22090 125068 22162
rect 125190 22162 125488 22372
rect 125190 22090 125388 22162
rect 125388 22090 125488 22162
rect 125610 22162 125908 22372
rect 125610 22090 125714 22162
rect 125714 22090 125814 22162
rect 125814 22090 125908 22162
rect 119028 20448 119326 20730
rect 119488 20448 119786 20730
rect 119888 20448 120186 20730
rect 120308 20448 120606 20730
rect 120728 20448 121026 20730
rect 119030 17770 119424 17934
rect 119522 17622 119666 17770
rect 119876 17610 120174 17892
rect 120296 17610 120594 17892
rect 120716 17610 121014 17892
rect 121136 17610 121434 17892
rect 121836 17802 121904 17892
rect 121904 17802 122004 17892
rect 122004 17802 122134 17892
rect 121836 17610 122134 17802
rect 122266 17802 122324 17892
rect 122324 17802 122424 17892
rect 122424 17802 122564 17892
rect 122266 17610 122564 17802
rect 122686 17802 122744 17892
rect 122744 17802 122844 17892
rect 122844 17802 122984 17892
rect 122686 17610 122984 17802
rect 123106 17802 123164 17892
rect 123164 17802 123264 17892
rect 123264 17802 123404 17892
rect 123106 17610 123404 17802
rect 123526 17802 123584 17892
rect 123584 17802 123684 17892
rect 123684 17802 123824 17892
rect 123526 17610 123824 17802
rect 123946 17802 124004 17892
rect 124004 17802 124104 17892
rect 124104 17802 124244 17892
rect 123946 17610 124244 17802
rect 124366 17802 124424 17892
rect 124424 17802 124524 17892
rect 124524 17802 124664 17892
rect 124366 17610 124664 17802
rect 124786 17802 124844 17892
rect 124844 17802 124944 17892
rect 124944 17802 125084 17892
rect 124786 17610 125084 17802
rect 125206 17802 125264 17892
rect 125264 17802 125364 17892
rect 125364 17802 125504 17892
rect 125206 17610 125504 17802
rect 125626 17802 125684 17892
rect 125684 17802 125784 17892
rect 125784 17802 125924 17892
rect 125626 17610 125924 17802
rect 126666 17886 126964 17892
rect 126666 17786 126746 17886
rect 126746 17786 126846 17886
rect 126846 17786 126964 17886
rect 126666 17610 126964 17786
rect 127116 17886 127414 17892
rect 127116 17786 127166 17886
rect 127166 17786 127266 17886
rect 127266 17786 127414 17886
rect 127116 17610 127414 17786
rect 127536 17886 127834 17892
rect 127536 17786 127586 17886
rect 127586 17786 127686 17886
rect 127686 17786 127834 17886
rect 127536 17610 127834 17786
rect 127956 17886 128254 17892
rect 127956 17786 128006 17886
rect 128006 17786 128106 17886
rect 128106 17786 128254 17886
rect 127956 17610 128254 17786
rect 128376 17886 128674 17892
rect 128376 17786 128426 17886
rect 128426 17786 128526 17886
rect 128526 17786 128674 17886
rect 128376 17610 128674 17786
rect 128796 17886 129094 17892
rect 128796 17786 128846 17886
rect 128846 17786 128946 17886
rect 128946 17786 129094 17886
rect 128796 17610 129094 17786
rect 129216 17886 129514 17892
rect 129216 17786 129266 17886
rect 129266 17786 129366 17886
rect 129366 17786 129514 17886
rect 129216 17610 129514 17786
rect 129636 17886 129934 17892
rect 129636 17786 129686 17886
rect 129686 17786 129786 17886
rect 129786 17786 129934 17886
rect 129636 17610 129934 17786
rect 130056 17886 130354 17892
rect 130056 17786 130106 17886
rect 130106 17786 130206 17886
rect 130206 17786 130354 17886
rect 130056 17610 130354 17786
rect 130476 17886 130774 17892
rect 130476 17786 130526 17886
rect 130526 17786 130626 17886
rect 130626 17786 130774 17886
rect 130476 17610 130774 17786
rect 130896 17886 131194 17892
rect 130896 17786 130946 17886
rect 130946 17786 131046 17886
rect 131046 17786 131194 17886
rect 130896 17610 131194 17786
rect 131316 17886 131614 17892
rect 131316 17786 131366 17886
rect 131366 17786 131466 17886
rect 131466 17786 131614 17886
rect 131316 17610 131614 17786
rect 131736 17886 132034 17892
rect 131736 17786 131786 17886
rect 131786 17786 131886 17886
rect 131886 17786 132034 17886
rect 131736 17610 132034 17786
rect 132156 17886 132454 17892
rect 132156 17786 132206 17886
rect 132206 17786 132306 17886
rect 132306 17786 132454 17886
rect 132156 17610 132454 17786
rect 132576 17886 132874 17892
rect 132576 17786 132626 17886
rect 132626 17786 132726 17886
rect 132726 17786 132874 17886
rect 132576 17610 132874 17786
rect 132996 17886 133294 17892
rect 132996 17786 133046 17886
rect 133046 17786 133146 17886
rect 133146 17786 133294 17886
rect 132996 17610 133294 17786
rect 133416 17886 133714 17892
rect 133416 17786 133466 17886
rect 133466 17786 133566 17886
rect 133566 17786 133714 17886
rect 133416 17610 133714 17786
rect 133836 17886 134134 17892
rect 133836 17786 133886 17886
rect 133886 17786 133986 17886
rect 133986 17786 134134 17886
rect 133836 17610 134134 17786
rect 134256 17886 134554 17892
rect 134256 17786 134306 17886
rect 134306 17786 134406 17886
rect 134406 17786 134554 17886
rect 134256 17610 134554 17786
rect 134676 17886 134974 17892
rect 134676 17786 134726 17886
rect 134726 17786 134826 17886
rect 134826 17786 134974 17886
rect 134676 17610 134974 17786
rect 135096 17886 135394 17892
rect 135096 17786 135146 17886
rect 135146 17786 135246 17886
rect 135246 17786 135394 17886
rect 135096 17610 135394 17786
rect 116734 17152 117062 17414
rect 116366 16958 116450 17044
rect 116364 15804 116448 15810
rect 116364 15730 116370 15804
rect 116370 15730 116440 15804
rect 116440 15730 116448 15804
rect 116364 15724 116448 15730
rect 116546 15804 116630 15810
rect 116546 15730 116552 15804
rect 116552 15730 116622 15804
rect 116622 15730 116630 15804
rect 116546 15724 116630 15730
rect 116364 15660 116448 15666
rect 115838 15620 115920 15626
rect 115838 15554 115844 15620
rect 115844 15554 115908 15620
rect 115908 15554 115920 15620
rect 116364 15586 116370 15660
rect 116370 15586 116440 15660
rect 116440 15586 116448 15660
rect 116364 15580 116448 15586
rect 116546 15660 116630 15666
rect 116546 15586 116552 15660
rect 116552 15586 116622 15660
rect 116622 15586 116630 15660
rect 116546 15580 116630 15586
rect 115838 15542 115920 15554
rect 115838 14586 115914 14594
rect 115838 14522 115842 14586
rect 115842 14522 115906 14586
rect 115906 14522 115914 14586
rect 115838 14518 115914 14522
rect 116366 14346 116450 14432
rect 116734 13976 117062 14238
rect 119030 13456 119424 13620
rect 119522 13620 119666 13768
rect 119876 13498 120174 13780
rect 120296 13498 120594 13780
rect 120716 13498 121014 13780
rect 121136 13498 121434 13780
rect 121836 13588 122134 13780
rect 121836 13498 121904 13588
rect 121904 13498 122004 13588
rect 122004 13498 122134 13588
rect 122266 13588 122564 13780
rect 122266 13498 122324 13588
rect 122324 13498 122424 13588
rect 122424 13498 122564 13588
rect 122686 13588 122984 13780
rect 122686 13498 122744 13588
rect 122744 13498 122844 13588
rect 122844 13498 122984 13588
rect 123106 13588 123404 13780
rect 123106 13498 123164 13588
rect 123164 13498 123264 13588
rect 123264 13498 123404 13588
rect 123526 13588 123824 13780
rect 123526 13498 123584 13588
rect 123584 13498 123684 13588
rect 123684 13498 123824 13588
rect 123946 13588 124244 13780
rect 123946 13498 124004 13588
rect 124004 13498 124104 13588
rect 124104 13498 124244 13588
rect 124366 13588 124664 13780
rect 124366 13498 124424 13588
rect 124424 13498 124524 13588
rect 124524 13498 124664 13588
rect 124786 13588 125084 13780
rect 124786 13498 124844 13588
rect 124844 13498 124944 13588
rect 124944 13498 125084 13588
rect 125206 13588 125504 13780
rect 125206 13498 125264 13588
rect 125264 13498 125364 13588
rect 125364 13498 125504 13588
rect 125626 13588 125924 13780
rect 125626 13498 125684 13588
rect 125684 13498 125784 13588
rect 125784 13498 125924 13588
rect 119028 10660 119326 10942
rect 119488 10660 119786 10942
rect 119888 10660 120186 10942
rect 120308 10660 120606 10942
rect 120728 10660 121026 10942
rect 121830 7828 122028 7900
rect 122028 7828 122128 7900
rect 121830 7618 122128 7828
rect 122250 7828 122448 7900
rect 122448 7828 122548 7900
rect 122250 7618 122548 7828
rect 122670 7828 122868 7900
rect 122868 7828 122968 7900
rect 122670 7618 122968 7828
rect 123090 7828 123288 7900
rect 123288 7828 123388 7900
rect 123090 7618 123388 7828
rect 123510 7828 123708 7900
rect 123708 7828 123808 7900
rect 123510 7618 123808 7828
rect 123930 7828 124128 7900
rect 124128 7828 124228 7900
rect 123930 7618 124228 7828
rect 124350 7828 124548 7900
rect 124548 7828 124648 7900
rect 124350 7618 124648 7828
rect 124770 7828 124968 7900
rect 124968 7828 125068 7900
rect 124770 7618 125068 7828
rect 125190 7828 125388 7900
rect 125388 7828 125488 7900
rect 125190 7618 125488 7828
rect 125610 7828 125714 7900
rect 125714 7828 125814 7900
rect 125814 7828 125908 7900
rect 125610 7618 125908 7828
<< metal3 >>
rect 101824 21608 117150 32954
rect 126658 28550 126976 28555
rect 126658 28268 126668 28550
rect 126966 28268 126976 28550
rect 126658 28263 126976 28268
rect 127108 28550 127426 28555
rect 127108 28268 127118 28550
rect 127416 28268 127426 28550
rect 127108 28263 127426 28268
rect 127528 28550 127846 28555
rect 127528 28268 127538 28550
rect 127836 28268 127846 28550
rect 127528 28263 127846 28268
rect 127948 28550 128266 28555
rect 127948 28268 127958 28550
rect 128256 28268 128266 28550
rect 127948 28263 128266 28268
rect 128368 28550 128686 28555
rect 128368 28268 128378 28550
rect 128676 28268 128686 28550
rect 128368 28263 128686 28268
rect 128788 28550 129106 28555
rect 128788 28268 128798 28550
rect 129096 28268 129106 28550
rect 128788 28263 129106 28268
rect 129208 28550 129526 28555
rect 129208 28268 129218 28550
rect 129516 28268 129526 28550
rect 129208 28263 129526 28268
rect 129628 28550 129946 28555
rect 129628 28268 129638 28550
rect 129936 28268 129946 28550
rect 129628 28263 129946 28268
rect 130048 28550 130366 28555
rect 130048 28268 130058 28550
rect 130356 28268 130366 28550
rect 130048 28263 130366 28268
rect 130468 28550 130786 28555
rect 130468 28268 130478 28550
rect 130776 28268 130786 28550
rect 130468 28263 130786 28268
rect 130888 28550 131206 28555
rect 130888 28268 130898 28550
rect 131196 28268 131206 28550
rect 130888 28263 131206 28268
rect 131308 28550 131626 28555
rect 131308 28268 131318 28550
rect 131616 28268 131626 28550
rect 131308 28263 131626 28268
rect 131728 28550 132046 28555
rect 131728 28268 131738 28550
rect 132036 28268 132046 28550
rect 131728 28263 132046 28268
rect 132148 28550 132466 28555
rect 132148 28268 132158 28550
rect 132456 28268 132466 28550
rect 132148 28263 132466 28268
rect 132568 28550 132886 28555
rect 132568 28268 132578 28550
rect 132876 28268 132886 28550
rect 132568 28263 132886 28268
rect 132988 28550 133306 28555
rect 132988 28268 132998 28550
rect 133296 28268 133306 28550
rect 132988 28263 133306 28268
rect 133408 28550 133726 28555
rect 133408 28268 133418 28550
rect 133716 28268 133726 28550
rect 133408 28263 133726 28268
rect 133828 28550 134146 28555
rect 133828 28268 133838 28550
rect 134136 28268 134146 28550
rect 133828 28263 134146 28268
rect 134248 28550 134566 28555
rect 134248 28268 134258 28550
rect 134556 28268 134566 28550
rect 134248 28263 134566 28268
rect 134668 28550 134986 28555
rect 134668 28268 134678 28550
rect 134976 28268 134986 28550
rect 134668 28263 134986 28268
rect 135088 28550 135406 28555
rect 135088 28268 135098 28550
rect 135396 28268 135406 28550
rect 135088 28263 135406 28268
rect 118988 27720 120998 27778
rect 121814 27720 125890 27848
rect 118988 27438 119692 27720
rect 119990 27438 120112 27720
rect 120410 27438 120532 27720
rect 120830 27438 120952 27720
rect 121250 27438 121260 27720
rect 121362 27438 121372 27720
rect 121670 27438 121680 27720
rect 121782 27438 121792 27720
rect 122090 27438 122212 27720
rect 122510 27438 122632 27720
rect 122930 27438 123052 27720
rect 123350 27438 123472 27720
rect 123770 27438 123892 27720
rect 124190 27438 124312 27720
rect 124610 27438 124732 27720
rect 125030 27438 125152 27720
rect 125450 27438 125890 27720
rect 118988 27300 120998 27438
rect 121814 27300 125890 27438
rect 118988 27018 119692 27300
rect 119990 27018 120112 27300
rect 120410 27018 120532 27300
rect 120830 27018 120952 27300
rect 121250 27018 121260 27300
rect 121362 27018 121372 27300
rect 121670 27018 121680 27300
rect 121782 27018 121792 27300
rect 122090 27018 122212 27300
rect 122510 27018 122632 27300
rect 122930 27018 123052 27300
rect 123350 27018 123472 27300
rect 123770 27018 123892 27300
rect 124190 27018 124312 27300
rect 124610 27018 124732 27300
rect 125030 27018 125152 27300
rect 125450 27018 125890 27300
rect 118988 21608 120998 27018
rect 121814 22377 125890 27018
rect 121814 22372 125918 22377
rect 121814 22090 121830 22372
rect 122128 22090 122250 22372
rect 122548 22090 122670 22372
rect 122968 22090 123090 22372
rect 123388 22090 123510 22372
rect 123808 22090 123930 22372
rect 124228 22090 124350 22372
rect 124648 22090 124770 22372
rect 125068 22090 125190 22372
rect 125488 22090 125610 22372
rect 125908 22090 125918 22372
rect 121814 22085 125918 22090
rect 121814 21826 125890 22085
rect 101824 21246 120998 21608
rect 101824 17654 117150 21246
rect 118988 20744 120998 21246
rect 118988 20730 121032 20744
rect 118988 20448 119028 20730
rect 119326 20448 119488 20730
rect 119786 20448 119888 20730
rect 120186 20448 120308 20730
rect 120606 20448 120728 20730
rect 121026 20448 121032 20730
rect 118988 20436 121032 20448
rect 118988 20192 120998 20436
rect 119020 17934 119434 17939
rect 119020 17770 119030 17934
rect 119424 17770 119434 17934
rect 119866 17892 120184 17897
rect 119020 17765 119434 17770
rect 119512 17770 119676 17775
rect 119512 17622 119522 17770
rect 119666 17622 119676 17770
rect 119512 17617 119676 17622
rect 119866 17610 119876 17892
rect 120174 17610 120184 17892
rect 119866 17605 120184 17610
rect 120286 17892 120604 17897
rect 120286 17610 120296 17892
rect 120594 17610 120604 17892
rect 120286 17605 120604 17610
rect 120706 17892 121024 17897
rect 120706 17610 120716 17892
rect 121014 17610 121024 17892
rect 120706 17605 121024 17610
rect 121126 17892 121444 17897
rect 121126 17610 121136 17892
rect 121434 17610 121444 17892
rect 121126 17605 121444 17610
rect 121826 17892 122144 17897
rect 121826 17610 121836 17892
rect 122134 17610 122144 17892
rect 121826 17605 122144 17610
rect 122256 17892 122574 17897
rect 122256 17610 122266 17892
rect 122564 17610 122574 17892
rect 122256 17605 122574 17610
rect 122676 17892 122994 17897
rect 122676 17610 122686 17892
rect 122984 17610 122994 17892
rect 122676 17605 122994 17610
rect 123096 17892 123414 17897
rect 123096 17610 123106 17892
rect 123404 17610 123414 17892
rect 123096 17605 123414 17610
rect 123516 17892 123834 17897
rect 123516 17610 123526 17892
rect 123824 17610 123834 17892
rect 123516 17605 123834 17610
rect 123936 17892 124254 17897
rect 123936 17610 123946 17892
rect 124244 17610 124254 17892
rect 123936 17605 124254 17610
rect 124356 17892 124674 17897
rect 124356 17610 124366 17892
rect 124664 17610 124674 17892
rect 124356 17605 124674 17610
rect 124776 17892 125094 17897
rect 124776 17610 124786 17892
rect 125084 17610 125094 17892
rect 124776 17605 125094 17610
rect 125196 17892 125514 17897
rect 125196 17610 125206 17892
rect 125504 17610 125514 17892
rect 125196 17605 125514 17610
rect 125616 17892 125934 17897
rect 125616 17610 125626 17892
rect 125924 17610 125934 17892
rect 125616 17605 125934 17610
rect 126656 17892 126974 17897
rect 126656 17610 126666 17892
rect 126964 17610 126974 17892
rect 126656 17605 126974 17610
rect 127106 17892 127424 17897
rect 127106 17610 127116 17892
rect 127414 17610 127424 17892
rect 127106 17605 127424 17610
rect 127526 17892 127844 17897
rect 127526 17610 127536 17892
rect 127834 17610 127844 17892
rect 127526 17605 127844 17610
rect 127946 17892 128264 17897
rect 127946 17610 127956 17892
rect 128254 17610 128264 17892
rect 127946 17605 128264 17610
rect 128366 17892 128684 17897
rect 128366 17610 128376 17892
rect 128674 17610 128684 17892
rect 128366 17605 128684 17610
rect 128786 17892 129104 17897
rect 128786 17610 128796 17892
rect 129094 17610 129104 17892
rect 128786 17605 129104 17610
rect 129206 17892 129524 17897
rect 129206 17610 129216 17892
rect 129514 17610 129524 17892
rect 129206 17605 129524 17610
rect 129626 17892 129944 17897
rect 129626 17610 129636 17892
rect 129934 17610 129944 17892
rect 129626 17605 129944 17610
rect 130046 17892 130364 17897
rect 130046 17610 130056 17892
rect 130354 17610 130364 17892
rect 130046 17605 130364 17610
rect 130466 17892 130784 17897
rect 130466 17610 130476 17892
rect 130774 17610 130784 17892
rect 130466 17605 130784 17610
rect 130886 17892 131204 17897
rect 130886 17610 130896 17892
rect 131194 17610 131204 17892
rect 130886 17605 131204 17610
rect 131306 17892 131624 17897
rect 131306 17610 131316 17892
rect 131614 17610 131624 17892
rect 131306 17605 131624 17610
rect 131726 17892 132044 17897
rect 131726 17610 131736 17892
rect 132034 17610 132044 17892
rect 131726 17605 132044 17610
rect 132146 17892 132464 17897
rect 132146 17610 132156 17892
rect 132454 17610 132464 17892
rect 132146 17605 132464 17610
rect 132566 17892 132884 17897
rect 132566 17610 132576 17892
rect 132874 17610 132884 17892
rect 132566 17605 132884 17610
rect 132986 17892 133304 17897
rect 132986 17610 132996 17892
rect 133294 17610 133304 17892
rect 132986 17605 133304 17610
rect 133406 17892 133724 17897
rect 133406 17610 133416 17892
rect 133714 17610 133724 17892
rect 133406 17605 133724 17610
rect 133826 17892 134144 17897
rect 133826 17610 133836 17892
rect 134134 17610 134144 17892
rect 133826 17605 134144 17610
rect 134246 17892 134564 17897
rect 134246 17610 134256 17892
rect 134554 17610 134564 17892
rect 134246 17605 134564 17610
rect 134666 17892 134984 17897
rect 134666 17610 134676 17892
rect 134974 17610 134984 17892
rect 134666 17605 134984 17610
rect 135086 17892 135404 17897
rect 135086 17610 135096 17892
rect 135394 17610 135404 17892
rect 135086 17605 135404 17610
rect 116724 17414 117072 17419
rect 116724 17152 116734 17414
rect 117062 17152 117072 17414
rect 116724 17147 117072 17152
rect 116356 17044 116460 17049
rect 116356 16958 116366 17044
rect 116450 16958 116460 17044
rect 116356 16953 116460 16958
rect 116354 15810 116458 15815
rect 116354 15724 116364 15810
rect 116448 15724 116458 15810
rect 116536 15810 116640 15815
rect 116536 15734 116546 15810
rect 116354 15666 116458 15724
rect 115828 15628 115930 15632
rect 115828 15536 115838 15628
rect 115920 15536 115930 15628
rect 116354 15580 116364 15666
rect 116448 15580 116458 15666
rect 116520 15724 116546 15734
rect 116630 15724 116640 15810
rect 116520 15666 116640 15724
rect 116520 15656 116546 15666
rect 116354 15575 116458 15580
rect 116536 15580 116546 15656
rect 116630 15580 116640 15666
rect 116536 15575 116640 15580
rect 115826 14600 115928 14606
rect 115824 14512 115834 14600
rect 115922 14512 115932 14600
rect 115826 14506 115928 14512
rect 116356 14432 116460 14437
rect 116356 14346 116366 14432
rect 116450 14346 116460 14432
rect 116356 14341 116460 14346
rect 116724 14238 117072 14243
rect 116724 13976 116734 14238
rect 117062 13976 117072 14238
rect 116724 13971 117072 13976
rect 119866 13780 120184 13785
rect 119512 13768 119676 13773
rect 101824 10144 117150 13736
rect 119020 13620 119434 13625
rect 119020 13456 119030 13620
rect 119424 13456 119434 13620
rect 119512 13620 119522 13768
rect 119666 13620 119676 13768
rect 119512 13615 119676 13620
rect 119866 13498 119876 13780
rect 120174 13498 120184 13780
rect 119866 13493 120184 13498
rect 120286 13780 120604 13785
rect 120286 13498 120296 13780
rect 120594 13498 120604 13780
rect 120286 13493 120604 13498
rect 120706 13780 121024 13785
rect 120706 13498 120716 13780
rect 121014 13498 121024 13780
rect 120706 13493 121024 13498
rect 121126 13780 121444 13785
rect 121126 13498 121136 13780
rect 121434 13498 121444 13780
rect 121126 13493 121444 13498
rect 121826 13780 122144 13785
rect 121826 13498 121836 13780
rect 122134 13498 122144 13780
rect 121826 13493 122144 13498
rect 122256 13780 122574 13785
rect 122256 13498 122266 13780
rect 122564 13498 122574 13780
rect 122256 13493 122574 13498
rect 122676 13780 122994 13785
rect 122676 13498 122686 13780
rect 122984 13498 122994 13780
rect 122676 13493 122994 13498
rect 123096 13780 123414 13785
rect 123096 13498 123106 13780
rect 123404 13498 123414 13780
rect 123096 13493 123414 13498
rect 123516 13780 123834 13785
rect 123516 13498 123526 13780
rect 123824 13498 123834 13780
rect 123516 13493 123834 13498
rect 123936 13780 124254 13785
rect 123936 13498 123946 13780
rect 124244 13498 124254 13780
rect 123936 13493 124254 13498
rect 124356 13780 124674 13785
rect 124356 13498 124366 13780
rect 124664 13498 124674 13780
rect 124356 13493 124674 13498
rect 124776 13780 125094 13785
rect 124776 13498 124786 13780
rect 125084 13498 125094 13780
rect 124776 13493 125094 13498
rect 125196 13780 125514 13785
rect 125196 13498 125206 13780
rect 125504 13498 125514 13780
rect 125196 13493 125514 13498
rect 125616 13780 125934 13785
rect 125616 13498 125626 13780
rect 125924 13498 125934 13780
rect 125616 13493 125934 13498
rect 119020 13451 119434 13456
rect 118988 10954 120998 11198
rect 118988 10942 121032 10954
rect 118988 10660 119028 10942
rect 119326 10660 119488 10942
rect 119786 10660 119888 10942
rect 120186 10660 120308 10942
rect 120606 10660 120728 10942
rect 121026 10660 121032 10942
rect 118988 10646 121032 10660
rect 118988 10144 120998 10646
rect 101824 9782 120998 10144
rect 101824 -1564 117150 9782
rect 118988 4372 120998 9782
rect 121814 7905 125890 8164
rect 121814 7900 125918 7905
rect 121814 7618 121830 7900
rect 122128 7618 122250 7900
rect 122548 7618 122670 7900
rect 122968 7618 123090 7900
rect 123388 7618 123510 7900
rect 123808 7618 123930 7900
rect 124228 7618 124350 7900
rect 124648 7618 124770 7900
rect 125068 7618 125190 7900
rect 125488 7618 125610 7900
rect 125908 7618 125918 7900
rect 121814 7613 125918 7618
rect 121814 4372 125890 7613
rect 118988 4090 119692 4372
rect 119990 4090 120112 4372
rect 120410 4090 120532 4372
rect 120830 4090 120952 4372
rect 121250 4090 121260 4372
rect 121362 4090 121372 4372
rect 121670 4090 121680 4372
rect 121782 4090 121792 4372
rect 122090 4090 122212 4372
rect 122510 4090 122632 4372
rect 122930 4090 123052 4372
rect 123350 4090 123472 4372
rect 123770 4090 123892 4372
rect 124190 4090 124312 4372
rect 124610 4090 124732 4372
rect 125030 4090 125152 4372
rect 125450 4090 125890 4372
rect 118988 3952 120998 4090
rect 121814 3952 125890 4090
rect 118988 3670 119692 3952
rect 119990 3670 120112 3952
rect 120410 3670 120532 3952
rect 120830 3670 120952 3952
rect 121250 3670 121260 3952
rect 121362 3670 121372 3952
rect 121670 3670 121680 3952
rect 121782 3670 121792 3952
rect 122090 3670 122212 3952
rect 122510 3670 122632 3952
rect 122930 3670 123052 3952
rect 123350 3670 123472 3952
rect 123770 3670 123892 3952
rect 124190 3670 124312 3952
rect 124610 3670 124732 3952
rect 125030 3670 125152 3952
rect 125450 3670 125890 3952
rect 118988 3612 120998 3670
rect 121814 3542 125890 3670
<< via3 >>
rect 126668 28268 126966 28550
rect 127118 28268 127416 28550
rect 127538 28268 127836 28550
rect 127958 28268 128256 28550
rect 128378 28268 128676 28550
rect 128798 28268 129096 28550
rect 129218 28268 129516 28550
rect 129638 28268 129936 28550
rect 130058 28268 130356 28550
rect 130478 28268 130776 28550
rect 130898 28268 131196 28550
rect 131318 28268 131616 28550
rect 131738 28268 132036 28550
rect 132158 28268 132456 28550
rect 132578 28268 132876 28550
rect 132998 28268 133296 28550
rect 133418 28268 133716 28550
rect 133838 28268 134136 28550
rect 134258 28268 134556 28550
rect 134678 28268 134976 28550
rect 135098 28268 135396 28550
rect 119692 27438 119990 27720
rect 120112 27438 120410 27720
rect 120532 27438 120830 27720
rect 120952 27438 121250 27720
rect 121372 27438 121670 27720
rect 121792 27438 122090 27720
rect 122212 27438 122510 27720
rect 122632 27438 122930 27720
rect 123052 27438 123350 27720
rect 123472 27438 123770 27720
rect 123892 27438 124190 27720
rect 124312 27438 124610 27720
rect 124732 27438 125030 27720
rect 125152 27438 125450 27720
rect 119692 27018 119990 27300
rect 120112 27018 120410 27300
rect 120532 27018 120830 27300
rect 120952 27018 121250 27300
rect 121372 27018 121670 27300
rect 121792 27018 122090 27300
rect 122212 27018 122510 27300
rect 122632 27018 122930 27300
rect 123052 27018 123350 27300
rect 123472 27018 123770 27300
rect 123892 27018 124190 27300
rect 124312 27018 124610 27300
rect 124732 27018 125030 27300
rect 125152 27018 125450 27300
rect 119030 17770 119424 17934
rect 119522 17622 119666 17770
rect 119876 17610 120174 17892
rect 120296 17610 120594 17892
rect 120716 17610 121014 17892
rect 121136 17610 121434 17892
rect 121836 17610 122134 17892
rect 122266 17610 122564 17892
rect 122686 17610 122984 17892
rect 123106 17610 123404 17892
rect 123526 17610 123824 17892
rect 123946 17610 124244 17892
rect 124366 17610 124664 17892
rect 124786 17610 125084 17892
rect 125206 17610 125504 17892
rect 125626 17610 125924 17892
rect 126666 17610 126964 17892
rect 127116 17610 127414 17892
rect 127536 17610 127834 17892
rect 127956 17610 128254 17892
rect 128376 17610 128674 17892
rect 128796 17610 129094 17892
rect 129216 17610 129514 17892
rect 129636 17610 129934 17892
rect 130056 17610 130354 17892
rect 130476 17610 130774 17892
rect 130896 17610 131194 17892
rect 131316 17610 131614 17892
rect 131736 17610 132034 17892
rect 132156 17610 132454 17892
rect 132576 17610 132874 17892
rect 132996 17610 133294 17892
rect 133416 17610 133714 17892
rect 133836 17610 134134 17892
rect 134256 17610 134554 17892
rect 134676 17610 134974 17892
rect 135096 17610 135394 17892
rect 116734 17152 117062 17414
rect 116366 16958 116450 17044
rect 116364 15724 116448 15810
rect 115838 15626 115920 15628
rect 115838 15542 115920 15626
rect 115838 15536 115920 15542
rect 116364 15580 116448 15666
rect 116546 15724 116630 15810
rect 116546 15580 116630 15666
rect 115834 14594 115922 14600
rect 115834 14518 115838 14594
rect 115838 14518 115914 14594
rect 115914 14518 115922 14594
rect 115834 14512 115922 14518
rect 116366 14346 116450 14432
rect 116734 13976 117062 14238
rect 119030 13456 119424 13620
rect 119522 13620 119666 13768
rect 119876 13498 120174 13780
rect 120296 13498 120594 13780
rect 120716 13498 121014 13780
rect 121136 13498 121434 13780
rect 121836 13498 122134 13780
rect 122266 13498 122564 13780
rect 122686 13498 122984 13780
rect 123106 13498 123404 13780
rect 123526 13498 123824 13780
rect 123946 13498 124244 13780
rect 124366 13498 124664 13780
rect 124786 13498 125084 13780
rect 125206 13498 125504 13780
rect 125626 13498 125924 13780
rect 119692 4090 119990 4372
rect 120112 4090 120410 4372
rect 120532 4090 120830 4372
rect 120952 4090 121250 4372
rect 121372 4090 121670 4372
rect 121792 4090 122090 4372
rect 122212 4090 122510 4372
rect 122632 4090 122930 4372
rect 123052 4090 123350 4372
rect 123472 4090 123770 4372
rect 123892 4090 124190 4372
rect 124312 4090 124610 4372
rect 124732 4090 125030 4372
rect 125152 4090 125450 4372
rect 119692 3670 119990 3952
rect 120112 3670 120410 3952
rect 120532 3670 120830 3952
rect 120952 3670 121250 3952
rect 121372 3670 121670 3952
rect 121792 3670 122090 3952
rect 122212 3670 122510 3952
rect 122632 3670 122930 3952
rect 123052 3670 123350 3952
rect 123472 3670 123770 3952
rect 123892 3670 124190 3952
rect 124312 3670 124610 3952
rect 124732 3670 125030 3952
rect 125152 3670 125450 3952
<< mimcap >>
rect 101925 32814 105475 32854
rect 101925 29344 101965 32814
rect 105435 29344 105475 32814
rect 101925 29304 105475 29344
rect 105794 32814 109344 32854
rect 105794 29344 105834 32814
rect 109304 29344 109344 32814
rect 105794 29304 109344 29344
rect 109663 32814 113213 32854
rect 109663 29344 109703 32814
rect 113173 29344 113213 32814
rect 109663 29304 113213 29344
rect 113532 32814 117082 32854
rect 113532 29344 113572 32814
rect 117042 29344 117082 32814
rect 113532 29304 117082 29344
rect 101925 28964 105475 29004
rect 101925 25494 101965 28964
rect 105435 25494 105475 28964
rect 101925 25454 105475 25494
rect 105794 28964 109344 29004
rect 105794 25494 105834 28964
rect 109304 25494 109344 28964
rect 105794 25454 109344 25494
rect 109663 28964 113213 29004
rect 109663 25494 109703 28964
rect 113173 25494 113213 28964
rect 109663 25454 113213 25494
rect 113532 28964 117082 29004
rect 113532 25494 113572 28964
rect 117042 25494 117082 28964
rect 113532 25454 117082 25494
rect 101925 25114 105475 25154
rect 101925 21644 101965 25114
rect 105435 21644 105475 25114
rect 101925 21604 105475 21644
rect 105794 25114 109344 25154
rect 105794 21644 105834 25114
rect 109304 21644 109344 25114
rect 105794 21604 109344 21644
rect 109663 25114 113213 25154
rect 109663 21644 109703 25114
rect 113173 21644 113213 25114
rect 109663 21604 113213 21644
rect 113532 25114 117082 25154
rect 113532 21644 113572 25114
rect 117042 21644 117082 25114
rect 113532 21604 117082 21644
rect 101925 21264 105475 21304
rect 101925 17794 101965 21264
rect 105435 17794 105475 21264
rect 101925 17754 105475 17794
rect 105794 21264 109344 21304
rect 105794 17794 105834 21264
rect 109304 17794 109344 21264
rect 105794 17754 109344 17794
rect 109663 21264 113213 21304
rect 109663 17794 109703 21264
rect 113173 17794 113213 21264
rect 109663 17754 113213 17794
rect 113532 21264 117082 21304
rect 113532 17794 113572 21264
rect 117042 17794 117082 21264
rect 113532 17754 117082 17794
rect 101925 13596 105475 13636
rect 101925 10126 101965 13596
rect 105435 10126 105475 13596
rect 101925 10086 105475 10126
rect 105794 13596 109344 13636
rect 105794 10126 105834 13596
rect 109304 10126 109344 13596
rect 105794 10086 109344 10126
rect 109663 13596 113213 13636
rect 109663 10126 109703 13596
rect 113173 10126 113213 13596
rect 109663 10086 113213 10126
rect 113532 13596 117082 13636
rect 113532 10126 113572 13596
rect 117042 10126 117082 13596
rect 113532 10086 117082 10126
rect 101925 9746 105475 9786
rect 101925 6276 101965 9746
rect 105435 6276 105475 9746
rect 101925 6236 105475 6276
rect 105794 9746 109344 9786
rect 105794 6276 105834 9746
rect 109304 6276 109344 9746
rect 105794 6236 109344 6276
rect 109663 9746 113213 9786
rect 109663 6276 109703 9746
rect 113173 6276 113213 9746
rect 109663 6236 113213 6276
rect 113532 9746 117082 9786
rect 113532 6276 113572 9746
rect 117042 6276 117082 9746
rect 113532 6236 117082 6276
rect 101925 5896 105475 5936
rect 101925 2426 101965 5896
rect 105435 2426 105475 5896
rect 101925 2386 105475 2426
rect 105794 5896 109344 5936
rect 105794 2426 105834 5896
rect 109304 2426 109344 5896
rect 105794 2386 109344 2426
rect 109663 5896 113213 5936
rect 109663 2426 109703 5896
rect 113173 2426 113213 5896
rect 109663 2386 113213 2426
rect 113532 5896 117082 5936
rect 113532 2426 113572 5896
rect 117042 2426 117082 5896
rect 113532 2386 117082 2426
rect 101925 2046 105475 2086
rect 101925 -1424 101965 2046
rect 105435 -1424 105475 2046
rect 101925 -1464 105475 -1424
rect 105794 2046 109344 2086
rect 105794 -1424 105834 2046
rect 109304 -1424 109344 2046
rect 105794 -1464 109344 -1424
rect 109663 2046 113213 2086
rect 109663 -1424 109703 2046
rect 113173 -1424 113213 2046
rect 109663 -1464 113213 -1424
rect 113532 2046 117082 2086
rect 113532 -1424 113572 2046
rect 117042 -1424 117082 2046
rect 113532 -1464 117082 -1424
<< mimcapcontact >>
rect 101965 29344 105435 32814
rect 105834 29344 109304 32814
rect 109703 29344 113173 32814
rect 113572 29344 117042 32814
rect 101965 25494 105435 28964
rect 105834 25494 109304 28964
rect 109703 25494 113173 28964
rect 113572 25494 117042 28964
rect 101965 21644 105435 25114
rect 105834 21644 109304 25114
rect 109703 21644 113173 25114
rect 113572 21644 117042 25114
rect 101965 17794 105435 21264
rect 105834 17794 109304 21264
rect 109703 17794 113173 21264
rect 113572 17794 117042 21264
rect 101965 10126 105435 13596
rect 105834 10126 109304 13596
rect 109703 10126 113173 13596
rect 113572 10126 117042 13596
rect 101965 6276 105435 9746
rect 105834 6276 109304 9746
rect 109703 6276 113173 9746
rect 113572 6276 117042 9746
rect 101965 2426 105435 5896
rect 105834 2426 109304 5896
rect 109703 2426 113173 5896
rect 113572 2426 117042 5896
rect 101965 -1424 105435 2046
rect 105834 -1424 109304 2046
rect 109703 -1424 113173 2046
rect 113572 -1424 117042 2046
<< metal4 >>
rect 103648 32954 103752 33004
rect 107517 32954 107621 33004
rect 111386 32954 111490 33004
rect 115255 32954 115359 33004
rect 101824 32814 117150 32954
rect 101824 29344 101965 32814
rect 105435 29344 105834 32814
rect 109304 29344 109703 32814
rect 113173 29344 113572 32814
rect 117042 29344 117150 32814
rect 101824 28964 117150 29344
rect 125914 29132 136482 29142
rect 101824 25494 101965 28964
rect 105435 25494 105834 28964
rect 109304 25494 109703 28964
rect 113173 25494 113572 28964
rect 117042 25494 117150 28964
rect 119338 28550 136626 29132
rect 119338 28474 126668 28550
rect 119312 28268 126668 28474
rect 126966 28268 127118 28550
rect 127416 28268 127538 28550
rect 127836 28268 127958 28550
rect 128256 28268 128378 28550
rect 128676 28268 128798 28550
rect 129096 28268 129218 28550
rect 129516 28268 129638 28550
rect 129936 28268 130058 28550
rect 130356 28268 130478 28550
rect 130776 28268 130898 28550
rect 131196 28268 131318 28550
rect 131616 28268 131738 28550
rect 132036 28268 132158 28550
rect 132456 28268 132578 28550
rect 132876 28268 132998 28550
rect 133296 28268 133418 28550
rect 133716 28268 133838 28550
rect 134136 28268 134258 28550
rect 134556 28268 134678 28550
rect 134976 28268 135098 28550
rect 135396 28268 136626 28550
rect 119312 27720 136626 28268
rect 119312 27648 119692 27720
rect 101824 25114 117150 25494
rect 101824 21644 101965 25114
rect 105435 21644 105834 25114
rect 109304 21644 109703 25114
rect 113173 21644 113572 25114
rect 117042 21644 117150 25114
rect 119310 27438 119692 27648
rect 119990 27438 120112 27720
rect 120410 27438 120532 27720
rect 120830 27438 120952 27720
rect 121250 27438 121372 27720
rect 121670 27438 121792 27720
rect 122090 27438 122212 27720
rect 122510 27438 122632 27720
rect 122930 27438 123052 27720
rect 123350 27438 123472 27720
rect 123770 27438 123892 27720
rect 124190 27438 124312 27720
rect 124610 27438 124732 27720
rect 125030 27438 125152 27720
rect 125450 27438 136626 27720
rect 119310 27300 136626 27438
rect 119310 27018 119692 27300
rect 119990 27018 120112 27300
rect 120410 27018 120532 27300
rect 120830 27018 120952 27300
rect 121250 27018 121372 27300
rect 121670 27018 121792 27300
rect 122090 27018 122212 27300
rect 122510 27018 122632 27300
rect 122930 27018 123052 27300
rect 123350 27018 123472 27300
rect 123770 27018 123892 27300
rect 124190 27018 124312 27300
rect 124610 27018 124732 27300
rect 125030 27018 125152 27300
rect 125450 27018 136626 27300
rect 119310 26832 136626 27018
rect 119310 22648 119668 26832
rect 101824 21264 117150 21644
rect 101824 17794 101965 21264
rect 105435 17794 105834 21264
rect 109304 17794 109703 21264
rect 113173 17794 113572 21264
rect 117042 17794 117150 21264
rect 101824 17654 117150 17794
rect 117396 22392 119668 22648
rect 116812 17415 116984 17654
rect 117396 17582 117636 22392
rect 116733 17414 117063 17415
rect 116733 17152 116734 17414
rect 117062 17152 117063 17414
rect 116733 17151 117063 17152
rect 117394 17054 117636 17582
rect 118618 17934 135602 17956
rect 118618 17770 119030 17934
rect 119424 17892 135602 17934
rect 119424 17770 119876 17892
rect 118618 17622 119522 17770
rect 119666 17622 119876 17770
rect 118618 17610 119876 17622
rect 120174 17610 120296 17892
rect 120594 17610 120716 17892
rect 121014 17610 121136 17892
rect 121434 17610 121836 17892
rect 122134 17610 122266 17892
rect 122564 17610 122686 17892
rect 122984 17610 123106 17892
rect 123404 17610 123526 17892
rect 123824 17610 123946 17892
rect 124244 17610 124366 17892
rect 124664 17610 124786 17892
rect 125084 17610 125206 17892
rect 125504 17610 125626 17892
rect 125924 17610 126666 17892
rect 126964 17610 127116 17892
rect 127414 17610 127536 17892
rect 127834 17610 127956 17892
rect 128254 17610 128376 17892
rect 128674 17610 128796 17892
rect 129094 17610 129216 17892
rect 129514 17610 129636 17892
rect 129934 17610 130056 17892
rect 130354 17610 130476 17892
rect 130774 17610 130896 17892
rect 131194 17610 131316 17892
rect 131614 17610 131736 17892
rect 132034 17610 132156 17892
rect 132454 17610 132576 17892
rect 132874 17610 132996 17892
rect 133294 17610 133416 17892
rect 133714 17610 133836 17892
rect 134134 17610 134256 17892
rect 134554 17610 134676 17892
rect 134974 17610 135096 17892
rect 135394 17610 135602 17892
rect 116356 17044 117646 17054
rect 116356 16958 116366 17044
rect 116450 16958 117646 17044
rect 116356 16948 117646 16958
rect 118618 16360 135602 17610
rect 115366 15810 135602 16360
rect 115366 15724 116364 15810
rect 116448 15724 116546 15810
rect 116630 15724 135602 15810
rect 115366 15666 135602 15724
rect 115366 15628 116364 15666
rect 115366 15536 115838 15628
rect 115920 15580 116364 15628
rect 116448 15580 116546 15666
rect 116630 15580 135602 15666
rect 115920 15536 135602 15580
rect 115366 15186 135602 15536
rect 115830 14600 116000 14606
rect 115830 14512 115834 14600
rect 115922 14512 116000 14600
rect 115830 14442 116000 14512
rect 115830 14432 117636 14442
rect 115830 14346 116366 14432
rect 116450 14346 117636 14432
rect 115830 14338 117636 14346
rect 116733 14238 117063 14239
rect 116733 13976 116734 14238
rect 117062 13976 117063 14238
rect 116733 13975 117063 13976
rect 116812 13736 116984 13975
rect 101824 13596 117150 13736
rect 101824 10126 101965 13596
rect 105435 10126 105834 13596
rect 109304 10126 109703 13596
rect 113173 10126 113572 13596
rect 117042 10126 117150 13596
rect 101824 9746 117150 10126
rect 101824 6276 101965 9746
rect 105435 6276 105834 9746
rect 109304 6276 109703 9746
rect 113173 6276 113572 9746
rect 117042 6276 117150 9746
rect 117396 8998 117636 14338
rect 118618 13780 135602 15186
rect 118618 13768 119876 13780
rect 118618 13620 119522 13768
rect 119666 13620 119876 13768
rect 118618 13456 119030 13620
rect 119424 13498 119876 13620
rect 120174 13498 120296 13780
rect 120594 13498 120716 13780
rect 121014 13498 121136 13780
rect 121434 13498 121836 13780
rect 122134 13498 122266 13780
rect 122564 13498 122686 13780
rect 122984 13498 123106 13780
rect 123404 13498 123526 13780
rect 123824 13498 123946 13780
rect 124244 13498 124366 13780
rect 124664 13498 124786 13780
rect 125084 13498 125206 13780
rect 125504 13498 125626 13780
rect 125924 13498 135602 13780
rect 119424 13456 135602 13498
rect 118618 13434 135602 13456
rect 117396 8742 119668 8998
rect 101824 5896 117150 6276
rect 101824 2426 101965 5896
rect 105435 2426 105834 5896
rect 109304 2426 109703 5896
rect 113173 2426 113572 5896
rect 117042 2426 117150 5896
rect 119310 4468 119668 8742
rect 119310 4372 125984 4468
rect 119310 4090 119692 4372
rect 119990 4090 120112 4372
rect 120410 4090 120532 4372
rect 120830 4090 120952 4372
rect 121250 4090 121372 4372
rect 121670 4090 121792 4372
rect 122090 4090 122212 4372
rect 122510 4090 122632 4372
rect 122930 4090 123052 4372
rect 123350 4090 123472 4372
rect 123770 4090 123892 4372
rect 124190 4090 124312 4372
rect 124610 4090 124732 4372
rect 125030 4090 125152 4372
rect 125450 4290 125984 4372
rect 125450 4090 126550 4290
rect 119310 3952 126550 4090
rect 119310 3670 119692 3952
rect 119990 3670 120112 3952
rect 120410 3670 120532 3952
rect 120830 3670 120952 3952
rect 121250 3670 121372 3952
rect 121670 3670 121792 3952
rect 122090 3670 122212 3952
rect 122510 3670 122632 3952
rect 122930 3670 123052 3952
rect 123350 3670 123472 3952
rect 123770 3670 123892 3952
rect 124190 3670 124312 3952
rect 124610 3670 124732 3952
rect 125030 3670 125152 3952
rect 125450 3670 126550 3952
rect 119310 2940 126550 3670
rect 119310 2916 125984 2940
rect 101824 2046 117150 2426
rect 101824 -1424 101965 2046
rect 105435 -1424 105834 2046
rect 109304 -1424 109703 2046
rect 113173 -1424 113572 2046
rect 117042 -1424 117150 2046
rect 101824 -1564 117150 -1424
<< labels >>
flabel metal4 128386 15178 128386 15178 0 FreeSans 8000 0 0 0 vdd
port 0 nsew
flabel metal2 124872 10760 124872 10760 0 FreeSans 8000 0 0 0 vn
port 3 nsew
flabel metal1 119362 19408 119362 19408 0 FreeSans 8000 0 0 0 vp1
flabel metal1 119352 11882 119352 11882 0 FreeSans 8000 0 0 0 vn1
flabel metal1 121712 20842 121712 20842 0 FreeSans 1600 0 0 0 vp2
flabel metal1 115624 15076 115624 15076 0 FreeSans 8000 0 0 0 vin
port 1 nsew
flabel metal1 126170 22210 126170 22210 0 FreeSans 8000 0 0 0 vp3
flabel metal2 133964 23632 133964 23632 0 FreeSans 8000 0 0 0 vp
port 2 nsew
flabel metal1 121666 9178 121666 9178 0 FreeSans 8000 0 0 0 vn2
flabel metal4 116478 15632 116478 15632 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal4 116556 14364 116556 14364 0 FreeSans 1600 0 0 0 vss
port 4 nsew
flabel metal1 116648 14968 116648 14968 0 FreeSans 1600 0 0 0 out
port 3 nsew
flabel via1 116532 14940 116532 14940 0 FreeSans 1600 0 0 0 A
port 2 nsew
flabel viali 116374 15020 116374 15020 0 FreeSans 1600 0 0 0 B
port 1 nsew
flabel metal4 116478 15758 116478 15758 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal4 116556 17026 116556 17026 0 FreeSans 1600 0 0 0 vss
port 4 nsew
flabel metal1 116648 16422 116648 16422 0 FreeSans 1600 0 0 0 out
port 3 nsew
flabel viali 116532 16450 116532 16450 0 FreeSans 1600 0 0 0 A
port 2 nsew
flabel via1 116374 16370 116374 16370 0 FreeSans 1600 0 0 0 B
port 1 nsew
flabel metal4 115972 15582 115972 15582 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal1 115828 14954 115828 14954 0 FreeSans 1600 0 0 0 A
port 1 nsew
flabel metal1 116004 14932 116004 14932 0 FreeSans 1600 0 0 0 B
port 2 nsew
flabel metal4 115970 14514 115970 14514 0 FreeSans 1600 0 0 0 vss
port 3 nsew
<< end >>
