* NGSPICE file created from half_driver.ext - technology: sky130A

.subckt half_driver vdd vp_p vp_n vss out_p
X0 vdd.t1499 vp_p.t0 out_p.t461 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1 out_p.t460 vp_p.t1 vdd.t1498 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2 vdd.t1497 vp_p.t2 out_p.t1213 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3 out_p.t1212 vp_p.t3 vdd.t1496 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4 out_p.t1033 vp_p.t4 vdd.t1495 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5 vss.t299 vp_n.t0 out_p.t112 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X6 out_p.t1032 vp_p.t5 vdd.t1494 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7 vss.t298 vp_n.t1 out_p.t113 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8 vdd.t1493 vp_p.t6 out_p.t1045 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9 vdd.t1492 vp_p.t7 out_p.t1044 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10 out_p.t1489 vp_p.t8 vdd.t1491 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X11 vdd.t1490 vp_p.t9 out_p.t1488 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X12 vdd.t1489 vp_p.t10 out_p.t263 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 vdd.t1488 vp_p.t11 out_p.t262 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X14 vdd.t1487 vp_p.t12 out_p.t1241 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X15 out_p.t1240 vp_p.t13 vdd.t1486 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X16 vss.t297 vp_n.t2 out_p.t106 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X17 out_p.t639 vp_p.t14 vdd.t1485 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 out_p.t638 vp_p.t15 vdd.t1484 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 out_p.t297 vp_p.t16 vdd.t1483 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X20 vdd.t1482 vp_p.t17 out_p.t296 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X21 out_p.t207 vp_p.t18 vdd.t1481 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X22 vdd.t1480 vp_p.t19 out_p.t206 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X23 vdd.t1479 vp_p.t20 out_p.t581 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X24 out_p.t580 vp_p.t21 vdd.t1478 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X25 vdd.t1477 vp_p.t22 out_p.t383 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X26 vdd.t1476 vp_p.t23 out_p.t382 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X27 out_p.t657 vp_p.t24 vdd.t1475 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X28 out_p.t107 vp_n.t3 vss.t296 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X29 vdd.t1474 vp_p.t25 out_p.t656 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X30 out_p.t1307 vp_p.t26 vdd.t1473 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X31 vss.t295 vp_n.t4 out_p.t1772 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X32 out_p.t1773 vp_n.t5 vss.t294 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X33 vdd.t1472 vp_p.t27 out_p.t1306 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X34 out_p.t42 vp_n.t6 vss.t293 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X35 vdd.t1471 vp_p.t28 out_p.t931 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X36 vdd.t1470 vp_p.t29 out_p.t930 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X37 vdd.t1469 vp_p.t30 out_p.t1075 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X38 out_p.t1074 vp_p.t31 vdd.t1468 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X39 vdd.t1467 vp_p.t32 out_p.t1451 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X40 vdd.t1466 vp_p.t33 out_p.t1450 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X41 vdd.t1465 vp_p.t34 out_p.t437 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X42 out_p.t436 vp_p.t35 vdd.t1464 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X43 out_p.t43 vp_n.t7 vss.t292 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X44 out_p.t1051 vp_p.t36 vdd.t1463 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X45 out_p.t1050 vp_p.t37 vdd.t1462 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X46 vdd.t1461 vp_p.t38 out_p.t1551 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X47 vdd.t1460 vp_p.t39 out_p.t1550 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X48 out_p.t457 vp_p.t40 vdd.t1459 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X49 out_p.t1748 vp_n.t8 vss.t291 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X50 vdd.t1458 vp_p.t41 out_p.t456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X51 vdd.t1457 vp_p.t42 out_p.t1593 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X52 out_p.t1592 vp_p.t43 vdd.t1456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X53 out_p.t1601 vp_p.t44 vdd.t1455 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X54 out_p.t1600 vp_p.t45 vdd.t1454 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X55 out_p.t239 vp_p.t46 vdd.t1453 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X56 vdd.t1452 vp_p.t47 out_p.t238 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X57 vdd.t1451 vp_p.t48 out_p.t1357 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X58 vss.t290 vp_n.t9 out_p.t1749 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X59 vdd.t1450 vp_p.t49 out_p.t1356 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X60 vdd.t1449 vp_p.t50 out_p.t745 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X61 vdd.t1448 vp_p.t51 out_p.t744 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X62 vss.t289 vp_n.t10 out_p.t22 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X63 out_p.t367 vp_p.t52 vdd.t1447 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X64 vdd.t1446 vp_p.t53 out_p.t366 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X65 out_p.t23 vp_n.t11 vss.t288 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X66 out_p.t1760 vp_n.t12 vss.t287 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X67 vdd.t1445 vp_p.t54 out_p.t223 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X68 out_p.t222 vp_p.t55 vdd.t1444 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X69 out_p.t1231 vp_p.t56 vdd.t1443 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X70 out_p.t1230 vp_p.t57 vdd.t1442 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X71 vdd.t1441 vp_p.t58 out_p.t1091 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X72 vdd.t1440 vp_p.t59 out_p.t1090 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X73 vdd.t1439 vp_p.t60 out_p.t933 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X74 vdd.t1438 vp_p.t61 out_p.t932 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X75 vdd.t1437 vp_p.t62 out_p.t1405 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X76 out_p.t1404 vp_p.t63 vdd.t1436 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X77 vss.t286 vp_n.t13 out_p.t1761 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X78 out_p.t1035 vp_p.t64 vdd.t1435 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X79 vdd.t1434 vp_p.t65 out_p.t1034 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X80 vdd.t1433 vp_p.t66 out_p.t1073 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X81 vdd.t1432 vp_p.t67 out_p.t1072 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X82 vdd.t1431 vp_p.t68 out_p.t1185 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X83 out_p.t1184 vp_p.t69 vdd.t1430 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X84 out_p.t1752 vp_n.t14 vss.t285 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X85 out_p.t375 vp_p.t70 vdd.t1429 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X86 out_p.t374 vp_p.t71 vdd.t1428 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X87 out_p.t1383 vp_p.t72 vdd.t1427 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X88 out_p.t1753 vp_n.t15 vss.t284 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X89 vss.t283 vp_n.t16 out_p.t36 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X90 vdd.t1426 vp_p.t73 out_p.t1382 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X91 out_p.t483 vp_p.t74 vdd.t1425 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X92 vdd.t1424 vp_p.t75 out_p.t482 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X93 vdd.t1423 vp_p.t76 out_p.t1303 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X94 out_p.t1302 vp_p.t77 vdd.t1422 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X95 vss.t282 vp_n.t17 out_p.t37 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X96 out_p.t1505 vp_p.t78 vdd.t1421 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X97 vdd.t1420 vp_p.t79 out_p.t1504 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X98 out_p.t547 vp_p.t80 vdd.t1419 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X99 vdd.t1418 vp_p.t81 out_p.t546 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X100 vss.t281 vp_n.t18 out_p.t122 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X101 vdd.t1417 vp_p.t82 out_p.t181 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X102 out_p.t180 vp_p.t83 vdd.t1416 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X103 out_p.t185 vp_p.t84 vdd.t1415 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X104 out_p.t123 vp_n.t19 vss.t280 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X105 out_p.t184 vp_p.t85 vdd.t1414 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X106 out_p.t963 vp_p.t86 vdd.t1413 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X107 vdd.t1412 vp_p.t87 out_p.t962 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X108 vdd.t1411 vp_p.t88 out_p.t395 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X109 out_p.t130 vp_n.t20 vss.t279 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X110 out_p.t131 vp_n.t21 vss.t278 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X111 out_p.t394 vp_p.t89 vdd.t1410 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X112 out_p.t435 vp_p.t90 vdd.t1409 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X113 vdd.t1408 vp_p.t91 out_p.t434 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X114 vdd.t1407 vp_p.t92 out_p.t937 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X115 out_p.t936 vp_p.t93 vdd.t1406 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X116 out_p.t1455 vp_p.t94 vdd.t1405 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X117 vdd.t1404 vp_p.t95 out_p.t1454 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X118 vdd.t1403 vp_p.t96 out_p.t535 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X119 vdd.t1402 vp_p.t97 out_p.t534 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X120 out_p.t631 vp_p.t98 vdd.t1401 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X121 vss.t277 vp_n.t22 out_p.t134 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X122 out_p.t135 vp_n.t23 vss.t276 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X123 out_p.t630 vp_p.t99 vdd.t1400 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X124 out_p.t241 vp_p.t100 vdd.t1399 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X125 vss.t275 vp_n.t24 out_p.t138 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X126 out_p.t240 vp_p.t101 vdd.t1398 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X127 vdd.t1397 vp_p.t102 out_p.t1107 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X128 out_p.t1106 vp_p.t103 vdd.t1396 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X129 vdd.t1395 vp_p.t104 out_p.t189 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X130 out_p.t188 vp_p.t105 vdd.t1394 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X131 out_p.t139 vp_n.t25 vss.t274 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X132 vdd.t1393 vp_p.t106 out_p.t625 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X133 vdd.t1392 vp_p.t107 out_p.t624 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X134 vdd.t1391 vp_p.t108 out_p.t343 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X135 out_p.t342 vp_p.t109 vdd.t1390 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X136 out_p.t311 vp_p.t110 vdd.t1389 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X137 out_p.t310 vp_p.t111 vdd.t1388 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X138 out_p.t1481 vp_p.t112 vdd.t1387 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X139 out_p.t1480 vp_p.t113 vdd.t1386 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X140 vdd.t1385 vp_p.t114 out_p.t1577 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X141 vdd.t1384 vp_p.t115 out_p.t1576 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X142 out_p.t753 vp_p.t116 vdd.t1383 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X143 vdd.t1382 vp_p.t117 out_p.t752 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X144 vdd.t1381 vp_p.t118 out_p.t1459 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X145 vdd.t1380 vp_p.t119 out_p.t1458 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X146 vdd.t1379 vp_p.t120 out_p.t725 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X147 out_p.t724 vp_p.t121 vdd.t1378 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X148 vdd.t1377 vp_p.t122 out_p.t583 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X149 vss.t273 vp_n.t26 out_p.t128 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X150 out_p.t582 vp_p.t123 vdd.t1376 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X151 vdd.t1375 vp_p.t124 out_p.t299 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X152 vdd.t1374 vp_p.t125 out_p.t298 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X153 vdd.t1373 vp_p.t126 out_p.t1579 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X154 vdd.t1372 vp_p.t127 out_p.t1578 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X155 vss.t272 vp_n.t27 out_p.t129 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X156 vdd.t1371 vp_p.t128 out_p.t681 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X157 out_p.t680 vp_p.t129 vdd.t1370 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X158 vss.t271 vp_n.t28 out_p.t108 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X159 vdd.t1369 vp_p.t130 out_p.t979 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X160 out_p.t978 vp_p.t131 vdd.t1368 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X161 out_p.t109 vp_n.t29 vss.t270 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X162 out_p.t847 vp_p.t132 vdd.t1367 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X163 vdd.t1366 vp_p.t133 out_p.t846 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X164 out_p.t523 vp_p.t134 vdd.t1365 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X165 out_p.t522 vp_p.t135 vdd.t1364 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X166 out_p.t1347 vp_p.t136 vdd.t1363 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X167 vdd.t1362 vp_p.t137 out_p.t1346 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X168 vdd.t1361 vp_p.t138 out_p.t209 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X169 vdd.t1360 vp_p.t139 out_p.t208 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X170 out_p.t84 vp_n.t30 vss.t269 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X171 vdd.t1359 vp_p.t140 out_p.t407 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X172 out_p.t406 vp_p.t141 vdd.t1358 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X173 out_p.t777 vp_p.t142 vdd.t1357 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X174 vdd.t1356 vp_p.t143 out_p.t776 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X175 vdd.t1355 vp_p.t144 out_p.t1201 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X176 vss.t268 vp_n.t31 out_p.t85 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X177 out_p.t1200 vp_p.t145 vdd.t1354 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X178 out_p.t469 vp_p.t146 vdd.t1353 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X179 out_p.t468 vp_p.t147 vdd.t1352 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X180 vdd.t1351 vp_p.t148 out_p.t173 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X181 vdd.t1350 vp_p.t149 out_p.t172 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X182 vdd.t1349 vp_p.t150 out_p.t565 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X183 vdd.t1348 vp_p.t151 out_p.t564 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X184 out_p.t1155 vp_p.t152 vdd.t1347 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X185 out_p.t1722 vp_n.t32 vss.t267 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X186 out_p.t1154 vp_p.t153 vdd.t1346 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X187 out_p.t1437 vp_p.t154 vdd.t1345 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X188 vdd.t1344 vp_p.t155 out_p.t1436 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X189 vdd.t1343 vp_p.t156 out_p.t793 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X190 vdd.t1342 vp_p.t157 out_p.t792 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X191 out_p.t425 vp_p.t158 vdd.t1341 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X192 out_p.t1723 vp_n.t33 vss.t266 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X193 vss.t265 vp_n.t34 out_p.t1684 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X194 out_p.t424 vp_p.t159 vdd.t1340 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X195 out_p.t1541 vp_p.t160 vdd.t1339 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X196 out_p.t1540 vp_p.t161 vdd.t1338 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X197 out_p.t1685 vp_n.t35 vss.t264 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X198 vdd.t1337 vp_p.t162 out_p.t957 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X199 vdd.t1336 vp_p.t163 out_p.t956 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X200 out_p.t213 vp_p.t164 vdd.t1335 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X201 out_p.t212 vp_p.t165 vdd.t1334 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X202 vdd.t1333 vp_p.t166 out_p.t763 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X203 out_p.t762 vp_p.t167 vdd.t1332 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X204 out_p.t1561 vp_p.t168 vdd.t1331 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X205 vdd.t1330 vp_p.t169 out_p.t1560 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X206 vdd.t1329 vp_p.t170 out_p.t389 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X207 out_p.t388 vp_p.t171 vdd.t1328 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X208 out_p.t475 vp_p.t172 vdd.t1327 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X209 vss.t263 vp_n.t36 out_p.t1724 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X210 vdd.t1326 vp_p.t173 out_p.t474 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X211 out_p.t969 vp_p.t174 vdd.t1325 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X212 vss.t262 vp_n.t37 out_p.t1725 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X213 out_p.t968 vp_p.t175 vdd.t1324 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X214 vdd.t1323 vp_p.t176 out_p.t1413 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X215 out_p.t1412 vp_p.t177 vdd.t1322 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X216 vdd.t1321 vp_p.t178 out_p.t233 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X217 vdd.t1320 vp_p.t179 out_p.t232 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X218 vdd.t1319 vp_p.t180 out_p.t545 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X219 vdd.t1318 vp_p.t181 out_p.t544 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X220 out_p.t1053 vp_p.t182 vdd.t1317 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X221 vss.t261 vp_n.t38 out_p.t46 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X222 out_p.t1052 vp_p.t183 vdd.t1316 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X223 out_p.t493 vp_p.t184 vdd.t1315 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X224 out_p.t492 vp_p.t185 vdd.t1314 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X225 vdd.t1313 vp_p.t186 out_p.t1227 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X226 out_p.t1226 vp_p.t187 vdd.t1312 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X227 vdd.t1311 vp_p.t188 out_p.t653 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X228 vdd.t1310 vp_p.t189 out_p.t652 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X229 out_p.t985 vp_p.t190 vdd.t1309 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X230 vdd.t1308 vp_p.t191 out_p.t984 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X231 out_p.t1093 vp_p.t192 vdd.t1307 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X232 out_p.t47 vp_n.t39 vss.t260 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X233 out_p.t1092 vp_p.t193 vdd.t1306 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X234 vdd.t1305 vp_p.t194 out_p.t1159 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X235 out_p.t1158 vp_p.t195 vdd.t1304 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X236 vss.t259 vp_n.t40 out_p.t68 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X237 out_p.t381 vp_p.t196 vdd.t1303 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X238 vdd.t1302 vp_p.t197 out_p.t380 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X239 out_p.t69 vp_n.t41 vss.t258 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X240 out_p.t1401 vp_p.t198 vdd.t1301 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X241 vdd.t1300 vp_p.t199 out_p.t1400 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X242 out_p.t1617 vp_p.t200 vdd.t1299 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X243 vdd.t1298 vp_p.t201 out_p.t1616 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X244 vdd.t1297 vp_p.t202 out_p.t877 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X245 vdd.t1296 vp_p.t203 out_p.t876 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X246 out_p.t167 vp_p.t204 vdd.t1295 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X247 out_p.t32 vp_n.t42 vss.t257 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X248 out_p.t166 vp_p.t205 vdd.t1294 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X249 vdd.t1293 vp_p.t206 out_p.t1149 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X250 out_p.t1148 vp_p.t207 vdd.t1292 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X251 out_p.t667 vp_p.t208 vdd.t1291 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X252 out_p.t666 vp_p.t209 vdd.t1290 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X253 out_p.t481 vp_p.t210 vdd.t1289 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X254 vdd.t1288 vp_p.t211 out_p.t480 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X255 out_p.t33 vp_n.t43 vss.t256 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X256 vdd.t1287 vp_p.t212 out_p.t1061 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X257 out_p.t1060 vp_p.t213 vdd.t1286 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X258 vdd.t1285 vp_p.t214 out_p.t943 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X259 vdd.t1284 vp_p.t215 out_p.t942 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X260 out_p.t539 vp_p.t216 vdd.t1283 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X261 out_p.t538 vp_p.t217 vdd.t1282 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X262 out_p.t369 vp_p.t218 vdd.t1281 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X263 out_p.t368 vp_p.t219 vdd.t1280 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X264 vdd.t1279 vp_p.t220 out_p.t1529 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X265 vdd.t1278 vp_p.t221 out_p.t1528 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X266 vss.t255 vp_n.t44 out_p.t1730 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X267 out_p.t513 vp_p.t222 vdd.t1277 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X268 vss.t254 vp_n.t45 out_p.t1731 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X269 vdd.t1276 vp_p.t223 out_p.t512 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X270 vdd.t1275 vp_p.t224 out_p.t1643 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X271 vss.t253 vp_n.t46 out_p.t116 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X272 out_p.t1642 vp_p.t225 vdd.t1274 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X273 out_p.t371 vp_p.t226 vdd.t1273 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X274 out_p.t370 vp_p.t227 vdd.t1272 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X275 vdd.t1271 vp_p.t228 out_p.t357 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X276 out_p.t356 vp_p.t229 vdd.t1270 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X277 vdd.t1269 vp_p.t230 out_p.t1031 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X278 out_p.t1030 vp_p.t231 vdd.t1268 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X279 out_p.t721 vp_p.t232 vdd.t1267 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X280 out_p.t720 vp_p.t233 vdd.t1266 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X281 vss.t252 vp_n.t47 out_p.t117 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X282 out_p.t1023 vp_p.t234 vdd.t1265 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X283 vdd.t1264 vp_p.t235 out_p.t1022 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X284 vdd.t1263 vp_p.t236 out_p.t703 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X285 vdd.t1262 vp_p.t237 out_p.t702 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X286 out_p.t1407 vp_p.t238 vdd.t1261 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X287 vdd.t1260 vp_p.t239 out_p.t1406 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X288 vdd.t1259 vp_p.t240 out_p.t621 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X289 out_p.t620 vp_p.t241 vdd.t1258 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X290 vdd.t1257 vp_p.t242 out_p.t1301 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X291 vdd.t1256 vp_p.t243 out_p.t1300 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X292 vdd.t1255 vp_p.t244 out_p.t859 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X293 out_p.t858 vp_p.t245 vdd.t1254 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X294 vdd.t1253 vp_p.t246 out_p.t559 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X295 out_p.t558 vp_p.t247 vdd.t1252 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X296 out_p.t94 vp_n.t48 vss.t251 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X297 out_p.t413 vp_p.t248 vdd.t1251 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X298 out_p.t412 vp_p.t249 vdd.t1250 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X299 out_p.t393 vp_p.t250 vdd.t1249 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X300 vdd.t1248 vp_p.t251 out_p.t392 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X301 out_p.t95 vp_n.t49 vss.t250 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X302 vss.t249 vp_n.t50 out_p.t1740 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X303 vdd.t1247 vp_p.t252 out_p.t1445 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X304 vdd.t1246 vp_p.t253 out_p.t1444 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X305 out_p.t285 vp_p.t254 vdd.t1245 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X306 vdd.t1244 vp_p.t255 out_p.t284 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X307 vss.t248 vp_n.t51 out_p.t1741 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X308 vdd.t1243 vp_p.t256 out_p.t1639 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X309 out_p.t1638 vp_p.t257 vdd.t1242 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X310 out_p.t567 vp_p.t258 vdd.t1241 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X311 vdd.t1240 vp_p.t259 out_p.t566 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X312 vdd.t1239 vp_p.t260 out_p.t569 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X313 vdd.t1238 vp_p.t261 out_p.t568 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X314 vdd.t1237 vp_p.t262 out_p.t1511 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X315 out_p.t1736 vp_n.t52 vss.t247 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X316 vdd.t1236 vp_p.t263 out_p.t1510 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X317 out_p.t1359 vp_p.t264 vdd.t1235 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X318 out_p.t1358 vp_p.t265 vdd.t1234 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X319 out_p.t1253 vp_p.t266 vdd.t1233 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X320 vdd.t1232 vp_p.t267 out_p.t1252 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X321 out_p.t1175 vp_p.t268 vdd.t1231 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X322 out_p.t1174 vp_p.t269 vdd.t1230 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X323 out_p.t1067 vp_p.t270 vdd.t1229 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X324 vdd.t1228 vp_p.t271 out_p.t1066 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X325 vdd.t1227 vp_p.t272 out_p.t865 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X326 vdd.t1226 vp_p.t273 out_p.t864 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X327 out_p.t291 vp_p.t274 vdd.t1225 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X328 out_p.t290 vp_p.t275 vdd.t1224 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X329 vdd.t1223 vp_p.t276 out_p.t809 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X330 vdd.t1222 vp_p.t277 out_p.t808 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X331 vss.t246 vp_n.t53 out_p.t1737 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X332 vdd.t1221 vp_p.t278 out_p.t273 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X333 vdd.t1220 vp_p.t279 out_p.t272 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X334 vdd.t1219 vp_p.t280 out_p.t1497 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X335 out_p.t1496 vp_p.t281 vdd.t1218 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X336 vdd.t1217 vp_p.t282 out_p.t363 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X337 vdd.t1216 vp_p.t283 out_p.t362 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X338 out_p.t150 vp_n.t54 vss.t245 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X339 out_p.t691 vp_p.t284 vdd.t1215 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X340 vss.t244 vp_n.t55 out_p.t151 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X341 vdd.t1214 vp_p.t285 out_p.t690 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X342 out_p.t439 vp_p.t286 vdd.t1213 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X343 out_p.t438 vp_p.t287 vdd.t1212 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X344 vdd.t1211 vp_p.t288 out_p.t527 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X345 out_p.t1744 vp_n.t56 vss.t243 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X346 vdd.t1210 vp_p.t289 out_p.t526 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X347 vdd.t1209 vp_p.t290 out_p.t799 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X348 out_p.t798 vp_p.t291 vdd.t1208 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X349 vdd.t1207 vp_p.t292 out_p.t805 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X350 out_p.t804 vp_p.t293 vdd.t1206 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X351 out_p.t1745 vp_n.t57 vss.t242 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X352 out_p.t281 vp_p.t294 vdd.t1205 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X353 vdd.t1204 vp_p.t295 out_p.t280 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X354 vdd.t1203 vp_p.t296 out_p.t1069 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X355 vdd.t1202 vp_p.t297 out_p.t1068 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X356 vss.t241 vp_n.t58 out_p.t48 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X357 vss.t240 vp_n.t59 out_p.t49 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X358 out_p.t491 vp_p.t298 vdd.t1201 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X359 vdd.t1200 vp_p.t299 out_p.t490 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X360 vdd.t1199 vp_p.t300 out_p.t1211 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X361 vss.t239 vp_n.t60 out_p.t78 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X362 out_p.t1210 vp_p.t301 vdd.t1198 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X363 out_p.t543 vp_p.t302 vdd.t1197 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X364 out_p.t542 vp_p.t303 vdd.t1196 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X365 out_p.t79 vp_n.t61 vss.t238 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X366 vdd.t1195 vp_p.t304 out_p.t1555 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X367 out_p.t1554 vp_p.t305 vdd.t1194 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X368 out_p.t1589 vp_p.t306 vdd.t1193 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X369 out_p.t1588 vp_p.t307 vdd.t1192 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X370 vdd.t1191 vp_p.t308 out_p.t231 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X371 out_p.t230 vp_p.t309 vdd.t1190 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X372 vss.t237 vp_n.t62 out_p.t1728 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X373 vdd.t1189 vp_p.t310 out_p.t623 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X374 vdd.t1188 vp_p.t311 out_p.t622 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X375 out_p.t1729 vp_n.t63 vss.t236 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X376 out_p.t1563 vp_p.t312 vdd.t1187 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X377 out_p.t102 vp_n.t64 vss.t235 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X378 vdd.t1186 vp_p.t313 out_p.t1562 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X379 vdd.t1185 vp_p.t314 out_p.t1495 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X380 vdd.t1184 vp_p.t315 out_p.t1494 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X381 out_p.t339 vp_p.t316 vdd.t1183 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X382 out_p.t338 vp_p.t317 vdd.t1182 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X383 out_p.t1647 vp_p.t318 vdd.t1181 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X384 vdd.t1180 vp_p.t319 out_p.t1646 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X385 vdd.t1179 vp_p.t320 out_p.t175 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X386 vdd.t1178 vp_p.t321 out_p.t174 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X387 out_p.t853 vp_p.t322 vdd.t1177 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X388 vdd.t1176 vp_p.t323 out_p.t852 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X389 out_p.t1017 vp_p.t324 vdd.t1175 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X390 out_p.t1016 vp_p.t325 vdd.t1174 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X391 vdd.t1173 vp_p.t326 out_p.t797 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X392 out_p.t796 vp_p.t327 vdd.t1172 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X393 out_p.t1571 vp_p.t328 vdd.t1171 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X394 out_p.t1570 vp_p.t329 vdd.t1170 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X395 out_p.t821 vp_p.t330 vdd.t1169 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X396 vdd.t1168 vp_p.t331 out_p.t820 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X397 out_p.t911 vp_p.t332 vdd.t1167 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X398 out_p.t103 vp_n.t65 vss.t234 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X399 vss.t233 vp_n.t66 out_p.t1786 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X400 out_p.t910 vp_p.t333 vdd.t1166 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X401 out_p.t345 vp_p.t334 vdd.t1165 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X402 out_p.t344 vp_p.t335 vdd.t1164 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X403 out_p.t1787 vp_n.t67 vss.t232 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X404 out_p.t541 vp_p.t336 vdd.t1163 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X405 vdd.t1162 vp_p.t337 out_p.t540 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X406 out_p.t1766 vp_n.t68 vss.t231 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X407 out_p.t1475 vp_p.t338 vdd.t1161 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X408 vdd.t1160 vp_p.t339 out_p.t1474 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X409 vdd.t1159 vp_p.t340 out_p.t1363 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X410 vss.t230 vp_n.t69 out_p.t1767 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X411 out_p.t1362 vp_p.t341 vdd.t1158 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X412 vdd.t1157 vp_p.t342 out_p.t1575 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X413 vdd.t1156 vp_p.t343 out_p.t1574 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X414 vdd.t1155 vp_p.t344 out_p.t1473 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X415 out_p.t1472 vp_p.t345 vdd.t1154 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X416 vdd.t1153 vp_p.t346 out_p.t1341 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X417 vdd.t1152 vp_p.t347 out_p.t1340 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X418 out_p.t1373 vp_p.t348 vdd.t1151 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X419 vss.t229 vp_n.t70 out_p.t28 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X420 vss.t228 vp_n.t71 out_p.t29 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X421 out_p.t1372 vp_p.t349 vdd.t1150 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X422 vdd.t1149 vp_p.t350 out_p.t1243 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X423 out_p.t1242 vp_p.t351 vdd.t1148 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X424 out_p.t1299 vp_p.t352 vdd.t1147 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X425 out_p.t1784 vp_n.t72 vss.t227 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X426 vdd.t1146 vp_p.t353 out_p.t1298 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X427 vdd.t1145 vp_p.t354 out_p.t265 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X428 vdd.t1144 vp_p.t355 out_p.t264 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X429 vdd.t1143 vp_p.t356 out_p.t1047 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X430 vdd.t1142 vp_p.t357 out_p.t1046 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X431 out_p.t669 vp_p.t358 vdd.t1141 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X432 out_p.t668 vp_p.t359 vdd.t1140 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X433 out_p.t293 vp_p.t360 vdd.t1139 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X434 vdd.t1138 vp_p.t361 out_p.t292 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X435 vdd.t1137 vp_p.t362 out_p.t1651 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X436 vdd.t1136 vp_p.t363 out_p.t1650 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X437 out_p.t1599 vp_p.t364 vdd.t1135 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X438 out_p.t1598 vp_p.t365 vdd.t1134 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X439 vdd.t1133 vp_p.t366 out_p.t683 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X440 vdd.t1132 vp_p.t367 out_p.t682 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X441 out_p.t179 vp_p.t368 vdd.t1131 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X442 vss.t226 vp_n.t73 out_p.t1785 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X443 out_p.t1782 vp_n.t74 vss.t225 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X444 vdd.t1130 vp_p.t369 out_p.t178 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X445 out_p.t1783 vp_n.t75 vss.t224 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X446 vdd.t1129 vp_p.t370 out_p.t1085 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X447 out_p.t1084 vp_p.t371 vdd.t1128 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X448 vdd.t1127 vp_p.t372 out_p.t1251 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X449 vdd.t1126 vp_p.t373 out_p.t1250 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X450 out_p.t693 vp_p.t374 vdd.t1125 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X451 out_p.t692 vp_p.t375 vdd.t1124 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X452 out_p.t701 vp_p.t376 vdd.t1123 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X453 vdd.t1122 vp_p.t377 out_p.t700 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X454 vdd.t1121 vp_p.t378 out_p.t1369 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X455 out_p.t1368 vp_p.t379 vdd.t1120 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X456 vdd.t1119 vp_p.t380 out_p.t451 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X457 out_p.t100 vp_n.t76 vss.t223 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X458 vdd.t1118 vp_p.t381 out_p.t450 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X459 out_p.t101 vp_n.t77 vss.t222 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X460 vdd.t1117 vp_p.t382 out_p.t1573 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X461 out_p.t1572 vp_p.t383 vdd.t1116 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X462 out_p.t261 vp_p.t384 vdd.t1115 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X463 out_p.t260 vp_p.t385 vdd.t1114 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X464 out_p.t627 vp_p.t386 vdd.t1113 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X465 out_p.t626 vp_p.t387 vdd.t1112 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X466 out_p.t1788 vp_n.t78 vss.t221 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X467 vdd.t1111 vp_p.t388 out_p.t801 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X468 out_p.t800 vp_p.t389 vdd.t1110 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X469 vdd.t1109 vp_p.t390 out_p.t817 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X470 vdd.t1108 vp_p.t391 out_p.t816 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X471 out_p.t1449 vp_p.t392 vdd.t1107 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X472 vdd.t1106 vp_p.t393 out_p.t1448 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X473 vss.t220 vp_n.t79 out_p.t1789 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X474 vss.t219 vp_n.t80 out_p.t34 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X475 vdd.t1105 vp_p.t394 out_p.t1057 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X476 out_p.t1056 vp_p.t395 vdd.t1104 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X477 out_p.t35 vp_n.t81 vss.t218 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X478 out_p.t1708 vp_n.t82 vss.t217 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X479 vdd.t1103 vp_p.t396 out_p.t1077 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X480 out_p.t1076 vp_p.t397 vdd.t1102 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X481 vdd.t1101 vp_p.t398 out_p.t1465 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X482 out_p.t1464 vp_p.t399 vdd.t1100 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X483 vdd.t1099 vp_p.t400 out_p.t643 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X484 out_p.t642 vp_p.t401 vdd.t1098 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X485 out_p.t983 vp_p.t402 vdd.t1097 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X486 vdd.t1096 vp_p.t403 out_p.t982 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X487 out_p.t783 vp_p.t404 vdd.t1095 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X488 vss.t216 vp_n.t83 out_p.t1709 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X489 out_p.t782 vp_p.t405 vdd.t1094 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X490 vss.t215 vp_n.t84 out_p.t1674 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X491 vdd.t1093 vp_p.t406 out_p.t1127 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X492 vdd.t1092 vp_p.t407 out_p.t1126 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X493 vdd.t1091 vp_p.t408 out_p.t1327 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X494 vdd.t1090 vp_p.t409 out_p.t1326 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X495 out_p.t401 vp_p.t410 vdd.t1089 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X496 out_p.t400 vp_p.t411 vdd.t1088 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X497 out_p.t1101 vp_p.t412 vdd.t1087 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X498 out_p.t1100 vp_p.t413 vdd.t1086 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X499 vdd.t1085 vp_p.t414 out_p.t1319 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X500 out_p.t1318 vp_p.t415 vdd.t1084 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X501 out_p.t741 vp_p.t416 vdd.t1083 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X502 out_p.t1675 vp_n.t85 vss.t214 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X503 vdd.t1082 vp_p.t417 out_p.t740 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X504 out_p.t387 vp_p.t418 vdd.t1081 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X505 out_p.t1796 vp_n.t86 vss.t213 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X506 out_p.t386 vp_p.t419 vdd.t1080 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X507 vdd.t1079 vp_p.t420 out_p.t953 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X508 out_p.t1797 vp_n.t87 vss.t212 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X509 vss.t211 vp_n.t88 out_p.t1656 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X510 vdd.t1078 vp_p.t421 out_p.t952 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X511 vdd.t1077 vp_p.t422 out_p.t1321 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X512 vdd.t1076 vp_p.t423 out_p.t1320 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X513 out_p.t253 vp_p.t424 vdd.t1075 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X514 out_p.t252 vp_p.t425 vdd.t1074 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X515 out_p.t645 vp_p.t426 vdd.t1073 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X516 vdd.t1072 vp_p.t427 out_p.t644 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X517 vdd.t1071 vp_p.t428 out_p.t431 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X518 out_p.t1657 vp_n.t89 vss.t210 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X519 out_p.t430 vp_p.t429 vdd.t1070 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X520 vdd.t1069 vp_p.t430 out_p.t1605 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X521 out_p.t74 vp_n.t90 vss.t209 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X522 out_p.t1604 vp_p.t431 vdd.t1068 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X523 out_p.t839 vp_p.t432 vdd.t1067 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X524 out_p.t838 vp_p.t433 vdd.t1066 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X525 vdd.t1065 vp_p.t434 out_p.t1263 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X526 out_p.t1262 vp_p.t435 vdd.t1064 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X527 out_p.t1011 vp_p.t436 vdd.t1063 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X528 vdd.t1062 vp_p.t437 out_p.t1010 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X529 vdd.t1061 vp_p.t438 out_p.t1535 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X530 vss.t208 vp_n.t91 out_p.t75 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X531 vss.t207 vp_n.t92 out_p.t16 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X532 vdd.t1060 vp_p.t439 out_p.t1534 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X533 out_p.t517 vp_p.t440 vdd.t1059 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X534 vdd.t1058 vp_p.t441 out_p.t516 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X535 vdd.t1057 vp_p.t442 out_p.t697 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X536 out_p.t17 vp_n.t93 vss.t206 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X537 out_p.t696 vp_p.t443 vdd.t1056 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X538 vdd.t1055 vp_p.t444 out_p.t1391 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X539 out_p.t1390 vp_p.t445 vdd.t1054 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X540 out_p.t665 vp_p.t446 vdd.t1053 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X541 out_p.t664 vp_p.t447 vdd.t1052 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X542 out_p.t965 vp_p.t448 vdd.t1051 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X543 vdd.t1050 vp_p.t449 out_p.t964 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X544 out_p.t1339 vp_p.t450 vdd.t1049 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X545 out_p.t1338 vp_p.t451 vdd.t1048 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X546 vdd.t1047 vp_p.t452 out_p.t895 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X547 out_p.t894 vp_p.t453 vdd.t1046 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X548 vdd.t1045 vp_p.t454 out_p.t195 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X549 vdd.t1044 vp_p.t455 out_p.t194 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X550 out_p.t967 vp_p.t456 vdd.t1043 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X551 vdd.t1042 vp_p.t457 out_p.t966 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X552 vss.t205 vp_n.t94 out_p.t1702 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X553 out_p.t257 vp_p.t458 vdd.t1041 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X554 out_p.t256 vp_p.t459 vdd.t1040 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X555 vdd.t1039 vp_p.t460 out_p.t1533 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X556 vdd.t1038 vp_p.t461 out_p.t1532 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X557 out_p.t1581 vp_p.t462 vdd.t1037 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X558 vdd.t1036 vp_p.t463 out_p.t1580 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X559 vdd.t1035 vp_p.t464 out_p.t1615 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X560 vss.t204 vp_n.t95 out_p.t1703 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X561 vdd.t1034 vp_p.t465 out_p.t1614 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X562 vdd.t1033 vp_p.t466 out_p.t731 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X563 out_p.t730 vp_p.t467 vdd.t1032 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X564 vdd.t1031 vp_p.t468 out_p.t1491 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X565 vdd.t1030 vp_p.t469 out_p.t1490 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X566 out_p.t1635 vp_p.t470 vdd.t1029 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X567 out_p.t1634 vp_p.t471 vdd.t1028 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X568 out_p.t126 vp_n.t96 vss.t203 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X569 vdd.t1027 vp_p.t472 out_p.t463 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X570 out_p.t462 vp_p.t473 vdd.t1026 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X571 out_p.t127 vp_n.t97 vss.t202 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X572 out_p.t229 vp_p.t474 vdd.t1025 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X573 vdd.t1024 vp_p.t475 out_p.t228 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X574 out_p.t675 vp_p.t476 vdd.t1023 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X575 out_p.t674 vp_p.t477 vdd.t1022 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X576 out_p.t1525 vp_p.t478 vdd.t1021 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X577 vss.t201 vp_n.t98 out_p.t142 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X578 vdd.t1020 vp_p.t479 out_p.t1524 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X579 out_p.t1281 vp_p.t480 vdd.t1019 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X580 out_p.t1280 vp_p.t481 vdd.t1018 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X581 out_p.t143 vp_n.t99 vss.t200 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X582 vdd.t1017 vp_p.t482 out_p.t1295 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X583 vdd.t1016 vp_p.t483 out_p.t1294 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X584 out_p.t1567 vp_p.t484 vdd.t1015 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X585 vdd.t1014 vp_p.t485 out_p.t1566 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X586 vss.t199 vp_n.t100 out_p.t1710 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X587 out_p.t1409 vp_p.t486 vdd.t1013 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X588 out_p.t1408 vp_p.t487 vdd.t1012 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X589 vdd.t1011 vp_p.t488 out_p.t749 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X590 out_p.t748 vp_p.t489 vdd.t1010 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X591 vdd.t1009 vp_p.t490 out_p.t199 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X592 out_p.t198 vp_p.t491 vdd.t1008 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X593 vss.t198 vp_n.t101 out_p.t1711 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X594 out_p.t455 vp_p.t492 vdd.t1007 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X595 out_p.t454 vp_p.t493 vdd.t1006 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X596 out_p.t211 vp_p.t494 vdd.t1005 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X597 out_p.t1706 vp_n.t102 vss.t197 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X598 out_p.t1707 vp_n.t103 vss.t196 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X599 vdd.t1004 vp_p.t495 out_p.t210 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X600 out_p.t359 vp_p.t496 vdd.t1003 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X601 out_p.t358 vp_p.t497 vdd.t1002 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X602 out_p.t687 vp_p.t498 vdd.t1001 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X603 vdd.t1000 vp_p.t499 out_p.t686 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X604 vdd.t999 vp_p.t500 out_p.t1603 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X605 vss.t195 vp_n.t104 out_p.t18 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X606 out_p.t1602 vp_p.t501 vdd.t998 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X607 out_p.t879 vp_p.t502 vdd.t997 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X608 vdd.t996 vp_p.t503 out_p.t878 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X609 vdd.t995 vp_p.t504 out_p.t419 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X610 vdd.t994 vp_p.t505 out_p.t418 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X611 vdd.t993 vp_p.t506 out_p.t1545 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X612 out_p.t1544 vp_p.t507 vdd.t992 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X613 vdd.t991 vp_p.t508 out_p.t1283 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X614 out_p.t19 vp_n.t105 vss.t194 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X615 out_p.t1282 vp_p.t509 vdd.t990 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X616 vss.t193 vp_n.t106 out_p.t1718 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X617 vdd.t989 vp_p.t510 out_p.t377 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X618 vss.t192 vp_n.t107 out_p.t1719 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X619 out_p.t376 vp_p.t511 vdd.t988 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X620 out_p.t579 vp_p.t512 vdd.t987 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X621 out_p.t578 vp_p.t513 vdd.t986 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X622 out_p.t515 vp_p.t514 vdd.t985 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X623 vdd.t984 vp_p.t515 out_p.t514 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X624 vdd.t983 vp_p.t516 out_p.t573 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X625 out_p.t572 vp_p.t517 vdd.t982 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X626 vdd.t981 vp_p.t518 out_p.t1109 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X627 out_p.t1108 vp_p.t519 vdd.t980 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X628 out_p.t921 vp_p.t520 vdd.t979 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X629 vdd.t978 vp_p.t521 out_p.t920 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X630 vdd.t977 vp_p.t522 out_p.t1493 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X631 out_p.t1492 vp_p.t523 vdd.t976 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X632 out_p.t1523 vp_p.t524 vdd.t975 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X633 vdd.t974 vp_p.t525 out_p.t1522 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X634 vdd.t973 vp_p.t526 out_p.t655 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X635 out_p.t1714 vp_n.t108 vss.t191 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X636 out_p.t654 vp_p.t527 vdd.t972 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X637 vdd.t971 vp_p.t528 out_p.t1333 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X638 vdd.t970 vp_p.t529 out_p.t1332 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X639 vdd.t969 vp_p.t530 out_p.t637 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X640 out_p.t636 vp_p.t531 vdd.t968 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X641 vss.t190 vp_n.t109 out_p.t1715 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X642 out_p.t146 vp_n.t110 vss.t189 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X643 vdd.t967 vp_p.t532 out_p.t609 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X644 vdd.t966 vp_p.t533 out_p.t608 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X645 vdd.t965 vp_p.t534 out_p.t1417 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X646 vss.t188 vp_n.t111 out_p.t147 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X647 vdd.t964 vp_p.t535 out_p.t1416 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X648 vdd.t963 vp_p.t536 out_p.t1039 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X649 out_p.t1038 vp_p.t537 vdd.t962 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X650 vss.t187 vp_n.t112 out_p.t1682 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X651 vdd.t961 vp_p.t538 out_p.t1223 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X652 out_p.t1222 vp_p.t539 vdd.t960 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X653 vdd.t959 vp_p.t540 out_p.t869 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X654 vdd.t958 vp_p.t541 out_p.t868 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X655 out_p.t1683 vp_n.t113 vss.t186 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X656 vdd.t957 vp_p.t542 out_p.t449 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X657 out_p.t448 vp_p.t543 vdd.t956 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X658 out_p.t651 vp_p.t544 vdd.t955 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X659 out_p.t650 vp_p.t545 vdd.t954 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X660 vdd.t953 vp_p.t546 out_p.t337 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X661 out_p.t336 vp_p.t547 vdd.t952 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X662 out_p.t991 vp_p.t548 vdd.t951 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X663 vdd.t950 vp_p.t549 out_p.t990 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X664 vdd.t949 vp_p.t550 out_p.t571 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X665 out_p.t1778 vp_n.t114 vss.t185 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X666 vdd.t948 vp_p.t551 out_p.t570 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X667 out_p.t1779 vp_n.t115 vss.t184 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X668 vdd.t947 vp_p.t552 out_p.t1337 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X669 vdd.t946 vp_p.t553 out_p.t1336 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X670 vdd.t945 vp_p.t554 out_p.t275 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X671 out_p.t274 vp_p.t555 vdd.t944 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X672 out_p.t473 vp_p.t556 vdd.t943 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X673 out_p.t472 vp_p.t557 vdd.t942 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X674 out_p.t1439 vp_p.t558 vdd.t941 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X675 out_p.t1438 vp_p.t559 vdd.t940 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X676 vdd.t939 vp_p.t560 out_p.t1125 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X677 vdd.t938 vp_p.t561 out_p.t1124 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X678 vdd.t937 vp_p.t562 out_p.t587 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X679 out_p.t586 vp_p.t563 vdd.t936 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X680 out_p.t737 vp_p.t564 vdd.t935 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X681 out_p.t736 vp_p.t565 vdd.t934 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X682 out_p.t1371 vp_p.t566 vdd.t933 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X683 out_p.t1370 vp_p.t567 vdd.t932 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X684 vdd.t931 vp_p.t568 out_p.t1331 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X685 out_p.t1764 vp_n.t116 vss.t183 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X686 vss.t182 vp_n.t117 out_p.t1765 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X687 out_p.t1330 vp_p.t569 vdd.t930 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X688 vss.t181 vp_n.t118 out_p.t1658 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X689 out_p.t1293 vp_p.t570 vdd.t929 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X690 out_p.t1292 vp_p.t571 vdd.t928 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X691 out_p.t485 vp_p.t572 vdd.t927 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X692 out_p.t484 vp_p.t573 vdd.t926 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X693 vdd.t925 vp_p.t574 out_p.t1065 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X694 vdd.t924 vp_p.t575 out_p.t1064 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X695 vdd.t923 vp_p.t576 out_p.t1165 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X696 out_p.t1164 vp_p.t577 vdd.t922 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X697 out_p.t1531 vp_p.t578 vdd.t921 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X698 vdd.t920 vp_p.t579 out_p.t1530 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X699 vdd.t919 vp_p.t580 out_p.t1487 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X700 out_p.t1486 vp_p.t581 vdd.t918 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X701 vss.t180 vp_n.t119 out_p.t1659 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X702 out_p.t1527 vp_p.t582 vdd.t917 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X703 vss.t179 vp_n.t120 out_p.t62 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X704 out_p.t1526 vp_p.t583 vdd.t916 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X705 vdd.t915 vp_p.t584 out_p.t219 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X706 vdd.t914 vp_p.t585 out_p.t218 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X707 vdd.t913 vp_p.t586 out_p.t341 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X708 out_p.t340 vp_p.t587 vdd.t912 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X709 out_p.t919 vp_p.t588 vdd.t911 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X710 vdd.t910 vp_p.t589 out_p.t918 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X711 out_p.t781 vp_p.t590 vdd.t909 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X712 vdd.t908 vp_p.t591 out_p.t780 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X713 out_p.t599 vp_p.t592 vdd.t907 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X714 out_p.t598 vp_p.t593 vdd.t906 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X715 out_p.t63 vp_n.t121 vss.t178 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X716 vdd.t905 vp_p.t594 out_p.t1257 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X717 out_p.t1726 vp_n.t122 vss.t177 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X718 vdd.t904 vp_p.t595 out_p.t1256 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X719 vss.t176 vp_n.t123 out_p.t1727 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X720 out_p.t1119 vp_p.t596 vdd.t903 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X721 out_p.t1118 vp_p.t597 vdd.t902 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X722 vdd.t901 vp_p.t598 out_p.t1099 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X723 vdd.t900 vp_p.t599 out_p.t1098 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X724 vdd.t899 vp_p.t600 out_p.t1083 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X725 out_p.t1082 vp_p.t601 vdd.t898 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X726 out_p.t989 vp_p.t602 vdd.t897 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X727 vdd.t896 vp_p.t603 out_p.t988 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X728 out_p.t409 vp_p.t604 vdd.t895 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X729 out_p.t408 vp_p.t605 vdd.t894 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X730 vdd.t893 vp_p.t606 out_p.t557 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X731 vdd.t892 vp_p.t607 out_p.t556 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X732 out_p.t1662 vp_n.t124 vss.t175 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X733 out_p.t1663 vp_n.t125 vss.t174 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X734 out_p.t951 vp_p.t608 vdd.t891 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X735 vdd.t890 vp_p.t609 out_p.t950 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X736 vdd.t889 vp_p.t610 out_p.t941 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X737 out_p.t940 vp_p.t611 vdd.t888 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X738 out_p.t1181 vp_p.t612 vdd.t887 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X739 vdd.t886 vp_p.t613 out_p.t1180 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X740 out_p.t611 vp_p.t614 vdd.t885 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X741 vdd.t884 vp_p.t615 out_p.t610 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X742 vdd.t883 vp_p.t616 out_p.t1353 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X743 vdd.t882 vp_p.t617 out_p.t1352 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X744 vdd.t881 vp_p.t618 out_p.t1517 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X745 vss.t173 vp_n.t126 out_p.t1768 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X746 vss.t172 vp_n.t127 out_p.t1769 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X747 vdd.t880 vp_p.t619 out_p.t1516 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X748 vss.t171 vp_n.t128 out_p.t1690 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X749 out_p.t601 vp_p.t620 vdd.t879 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X750 vdd.t878 vp_p.t621 out_p.t600 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X751 out_p.t1691 vp_n.t129 vss.t170 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X752 out_p.t1692 vp_n.t130 vss.t169 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X753 vdd.t877 vp_p.t622 out_p.t511 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X754 out_p.t510 vp_p.t623 vdd.t876 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X755 out_p.t1591 vp_p.t624 vdd.t875 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X756 out_p.t1590 vp_p.t625 vdd.t874 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X757 out_p.t505 vp_p.t626 vdd.t873 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X758 vdd.t872 vp_p.t627 out_p.t504 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X759 vdd.t871 vp_p.t628 out_p.t1457 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X760 vdd.t870 vp_p.t629 out_p.t1456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X761 vss.t168 vp_n.t131 out_p.t1693 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X762 vdd.t869 vp_p.t630 out_p.t305 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X763 out_p.t304 vp_p.t631 vdd.t868 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X764 vss.t167 vp_n.t132 out_p.t1694 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X765 out_p.t751 vp_p.t632 vdd.t867 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X766 vdd.t866 vp_p.t633 out_p.t750 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X767 vss.t166 vp_n.t133 out_p.t1695 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X768 vdd.t865 vp_p.t634 out_p.t575 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X769 vdd.t864 vp_p.t635 out_p.t574 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X770 vdd.t863 vp_p.t636 out_p.t661 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X771 out_p.t660 vp_p.t637 vdd.t862 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X772 out_p.t629 vp_p.t638 vdd.t861 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X773 out_p.t628 vp_p.t639 vdd.t860 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X774 out_p.t863 vp_p.t640 vdd.t859 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X775 out_p.t0 vp_n.t134 vss.t165 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X776 out_p.t1 vp_n.t135 vss.t164 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X777 vss.t163 vp_n.t136 out_p.t2 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X778 vdd.t858 vp_p.t641 out_p.t862 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X779 out_p.t1193 vp_p.t642 vdd.t857 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X780 vdd.t856 vp_p.t643 out_p.t1192 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X781 out_p.t771 vp_p.t644 vdd.t855 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X782 out_p.t770 vp_p.t645 vdd.t854 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X783 vdd.t853 vp_p.t646 out_p.t1269 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X784 vss.t162 vp_n.t137 out_p.t3 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X785 out_p.t1268 vp_p.t647 vdd.t852 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X786 vdd.t851 vp_p.t648 out_p.t945 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X787 vdd.t850 vp_p.t649 out_p.t944 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X788 vdd.t849 vp_p.t650 out_p.t237 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X789 vdd.t848 vp_p.t651 out_p.t236 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X790 out_p.t1311 vp_p.t652 vdd.t847 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X791 vdd.t846 vp_p.t653 out_p.t1310 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X792 out_p.t1275 vp_p.t654 vdd.t845 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X793 out_p.t1274 vp_p.t655 vdd.t844 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X794 vdd.t843 vp_p.t656 out_p.t267 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X795 vdd.t842 vp_p.t657 out_p.t266 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X796 vdd.t841 vp_p.t658 out_p.t1343 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X797 out_p.t26 vp_n.t138 vss.t161 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X798 out_p.t1342 vp_p.t659 vdd.t840 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X799 vdd.t839 vp_p.t660 out_p.t813 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X800 vdd.t838 vp_p.t661 out_p.t812 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X801 vss.t160 vp_n.t139 out_p.t27 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X802 out_p.t423 vp_p.t662 vdd.t837 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X803 vdd.t836 vp_p.t663 out_p.t422 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X804 out_p.t1217 vp_p.t664 vdd.t835 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X805 out_p.t1216 vp_p.t665 vdd.t834 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X806 out_p.t38 vp_n.t140 vss.t159 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X807 out_p.t39 vp_n.t141 vss.t158 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X808 out_p.t1029 vp_p.t666 vdd.t833 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X809 vdd.t832 vp_p.t667 out_p.t1028 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X810 vdd.t831 vp_p.t668 out_p.t1105 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X811 out_p.t1104 vp_p.t669 vdd.t830 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X812 out_p.t1133 vp_p.t670 vdd.t829 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X813 vdd.t828 vp_p.t671 out_p.t1132 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X814 vss.t157 vp_n.t142 out_p.t30 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X815 vdd.t827 vp_p.t672 out_p.t1089 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X816 vss.t156 vp_n.t143 out_p.t31 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X817 out_p.t1088 vp_p.t673 vdd.t826 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X818 out_p.t999 vp_p.t674 vdd.t825 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X819 vss.t155 vp_n.t144 out_p.t24 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X820 out_p.t998 vp_p.t675 vdd.t824 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X821 out_p.t923 vp_p.t676 vdd.t823 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X822 vdd.t822 vp_p.t677 out_p.t922 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X823 vdd.t821 vp_p.t678 out_p.t1229 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X824 vdd.t820 vp_p.t679 out_p.t1228 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X825 out_p.t833 vp_p.t680 vdd.t819 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X826 out_p.t25 vp_n.t145 vss.t154 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X827 vdd.t818 vp_p.t681 out_p.t832 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X828 out_p.t1597 vp_p.t682 vdd.t817 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X829 vdd.t816 vp_p.t683 out_p.t1596 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X830 vss.t153 vp_n.t146 out_p.t82 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X831 out_p.t871 vp_p.t684 vdd.t815 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X832 out_p.t870 vp_p.t685 vdd.t814 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X833 out_p.t595 vp_p.t686 vdd.t813 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X834 vdd.t812 vp_p.t687 out_p.t594 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X835 out_p.t215 vp_p.t688 vdd.t811 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X836 out_p.t214 vp_p.t689 vdd.t810 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X837 vdd.t809 vp_p.t690 out_p.t747 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X838 vdd.t808 vp_p.t691 out_p.t746 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X839 out_p.t1037 vp_p.t692 vdd.t807 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X840 vdd.t806 vp_p.t693 out_p.t1036 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X841 out_p.t83 vp_n.t147 vss.t152 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X842 vss.t151 vp_n.t148 out_p.t86 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X843 vdd.t805 vp_p.t694 out_p.t1189 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X844 vdd.t804 vp_p.t695 out_p.t1188 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X845 vdd.t803 vp_p.t696 out_p.t899 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X846 vss.t150 vp_n.t149 out_p.t87 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X847 out_p.t898 vp_p.t697 vdd.t802 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X848 vdd.t801 vp_p.t698 out_p.t827 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X849 vdd.t800 vp_p.t699 out_p.t826 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X850 out_p.t1637 vp_p.t700 vdd.t799 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X851 out_p.t1636 vp_p.t701 vdd.t798 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X852 out_p.t939 vp_p.t702 vdd.t797 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X853 out_p.t1700 vp_n.t150 vss.t149 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X854 vdd.t796 vp_p.t703 out_p.t938 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X855 vdd.t795 vp_p.t704 out_p.t221 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X856 out_p.t220 vp_p.t705 vdd.t794 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X857 out_p.t1585 vp_p.t706 vdd.t793 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X858 out_p.t1584 vp_p.t707 vdd.t792 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X859 vdd.t791 vp_p.t708 out_p.t1335 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X860 out_p.t1334 vp_p.t709 vdd.t790 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X861 vdd.t789 vp_p.t710 out_p.t355 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X862 vss.t148 vp_n.t151 out_p.t1701 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X863 out_p.t354 vp_p.t711 vdd.t788 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X864 out_p.t1774 vp_n.t152 vss.t147 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X865 out_p.t1623 vp_p.t712 vdd.t787 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X866 out_p.t1775 vp_n.t153 vss.t146 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X867 vdd.t786 vp_p.t713 out_p.t1622 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X868 vdd.t785 vp_p.t714 out_p.t471 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X869 vdd.t784 vp_p.t715 out_p.t470 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X870 vdd.t783 vp_p.t716 out_p.t815 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X871 out_p.t814 vp_p.t717 vdd.t782 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X872 out_p.t857 vp_p.t718 vdd.t781 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X873 vdd.t780 vp_p.t719 out_p.t856 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X874 vdd.t779 vp_p.t720 out_p.t917 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X875 vdd.t778 vp_p.t721 out_p.t916 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X876 out_p.t689 vp_p.t722 vdd.t777 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X877 out_p.t688 vp_p.t723 vdd.t776 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X878 vdd.t775 vp_p.t724 out_p.t1015 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X879 out_p.t1014 vp_p.t725 vdd.t774 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X880 out_p.t591 vp_p.t726 vdd.t773 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X881 out_p.t590 vp_p.t727 vdd.t772 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X882 vss.t145 vp_n.t154 out_p.t1666 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X883 out_p.t1477 vp_p.t728 vdd.t771 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X884 out_p.t1476 vp_p.t729 vdd.t770 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X885 vdd.t769 vp_p.t730 out_p.t1183 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X886 vdd.t768 vp_p.t731 out_p.t1182 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X887 out_p.t1667 vp_n.t155 vss.t144 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X888 vss.t143 vp_n.t156 out_p.t1720 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X889 out_p.t1163 vp_p.t732 vdd.t767 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X890 out_p.t1162 vp_p.t733 vdd.t766 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X891 out_p.t443 vp_p.t734 vdd.t765 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X892 out_p.t442 vp_p.t735 vdd.t764 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X893 vdd.t763 vp_p.t736 out_p.t1225 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X894 out_p.t1721 vp_n.t157 vss.t142 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X895 out_p.t1224 vp_p.t737 vdd.t762 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X896 vdd.t761 vp_p.t738 out_p.t1361 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X897 vdd.t760 vp_p.t739 out_p.t1360 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X898 out_p.t521 vp_p.t740 vdd.t759 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X899 out_p.t520 vp_p.t741 vdd.t758 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X900 out_p.t1325 vp_p.t742 vdd.t757 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X901 vdd.t756 vp_p.t743 out_p.t1324 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X902 vss.t141 vp_n.t158 out_p.t1668 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X903 vdd.t755 vp_p.t744 out_p.t807 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X904 vdd.t754 vp_p.t745 out_p.t806 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X905 vdd.t753 vp_p.t746 out_p.t1207 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X906 vdd.t752 vp_p.t747 out_p.t1206 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X907 vdd.t751 vp_p.t748 out_p.t421 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X908 out_p.t420 vp_p.t749 vdd.t750 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X909 vdd.t749 vp_p.t750 out_p.t761 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X910 vdd.t748 vp_p.t751 out_p.t760 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X911 out_p.t459 vp_p.t752 vdd.t747 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X912 vss.t140 vp_n.t159 out_p.t1669 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X913 vss.t139 vp_n.t160 out_p.t1672 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X914 out_p.t458 vp_p.t753 vdd.t746 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X915 out_p.t1187 vp_p.t754 vdd.t745 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X916 out_p.t1186 vp_p.t755 vdd.t744 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X917 vdd.t743 vp_p.t756 out_p.t767 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X918 vdd.t742 vp_p.t757 out_p.t766 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X919 vdd.t741 vp_p.t758 out_p.t1547 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X920 out_p.t1546 vp_p.t759 vdd.t740 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X921 vdd.t739 vp_p.t760 out_p.t997 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X922 out_p.t996 vp_p.t761 vdd.t738 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X923 vdd.t737 vp_p.t762 out_p.t441 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X924 out_p.t440 vp_p.t763 vdd.t736 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X925 out_p.t913 vp_p.t764 vdd.t735 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X926 vss.t138 vp_n.t161 out_p.t1673 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X927 out_p.t1670 vp_n.t162 vss.t137 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X928 out_p.t1671 vp_n.t163 vss.t136 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X929 vdd.t734 vp_p.t765 out_p.t912 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X930 vdd.t733 vp_p.t766 out_p.t779 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X931 vss.t135 vp_n.t164 out_p.t1680 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X932 vdd.t732 vp_p.t767 out_p.t778 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X933 vdd.t731 vp_p.t768 out_p.t283 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X934 vdd.t730 vp_p.t769 out_p.t282 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X935 out_p.t717 vp_p.t770 vdd.t729 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X936 out_p.t716 vp_p.t771 vdd.t728 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X937 out_p.t295 vp_p.t772 vdd.t727 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X938 out_p.t294 vp_p.t773 vdd.t726 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X939 out_p.t1385 vp_p.t774 vdd.t725 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X940 vdd.t724 vp_p.t775 out_p.t1384 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X941 vdd.t723 vp_p.t776 out_p.t1003 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X942 out_p.t1681 vp_n.t165 vss.t134 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X943 vdd.t722 vp_p.t777 out_p.t1002 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X944 out_p.t1509 vp_p.t778 vdd.t721 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X945 out_p.t1508 vp_p.t779 vdd.t720 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X946 out_p.t1287 vp_p.t780 vdd.t719 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X947 out_p.t1286 vp_p.t781 vdd.t718 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X948 vdd.t717 vp_p.t782 out_p.t243 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X949 out_p.t242 vp_p.t783 vdd.t716 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X950 vdd.t715 vp_p.t784 out_p.t1485 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X951 vdd.t714 vp_p.t785 out_p.t1484 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X952 vdd.t713 vp_p.t786 out_p.t955 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X953 vss.t133 vp_n.t166 out_p.t1678 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X954 vdd.t712 vp_p.t787 out_p.t954 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X955 vdd.t711 vp_p.t788 out_p.t685 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X956 out_p.t684 vp_p.t789 vdd.t710 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X957 vss.t132 vp_n.t167 out_p.t1679 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X958 vss.t131 vp_n.t168 out_p.t118 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X959 out_p.t995 vp_p.t790 vdd.t709 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X960 out_p.t994 vp_p.t791 vdd.t708 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X961 out_p.t119 vp_n.t169 vss.t130 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X962 out_p.t255 vp_p.t792 vdd.t707 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X963 vdd.t706 vp_p.t793 out_p.t254 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X964 out_p.t1553 vp_p.t794 vdd.t705 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X965 out_p.t1552 vp_p.t795 vdd.t704 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X966 vdd.t703 vp_p.t796 out_p.t713 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X967 vdd.t702 vp_p.t797 out_p.t712 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X968 out_p.t519 vp_p.t798 vdd.t701 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X969 vdd.t700 vp_p.t799 out_p.t518 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X970 vdd.t699 vp_p.t800 out_p.t323 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X971 out_p.t322 vp_p.t801 vdd.t698 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X972 vdd.t697 vp_p.t802 out_p.t217 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X973 out_p.t216 vp_p.t803 vdd.t696 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X974 vdd.t695 vp_p.t804 out_p.t1367 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X975 out_p.t1366 vp_p.t805 vdd.t694 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X976 out_p.t1379 vp_p.t806 vdd.t693 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X977 vss.t129 vp_n.t170 out_p.t1798 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X978 vdd.t692 vp_p.t807 out_p.t1378 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X979 vdd.t691 vp_p.t808 out_p.t1059 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X980 out_p.t1058 vp_p.t809 vdd.t690 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X981 out_p.t1245 vp_p.t810 vdd.t689 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X982 out_p.t1244 vp_p.t811 vdd.t688 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X983 out_p.t1025 vp_p.t812 vdd.t687 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X984 out_p.t1024 vp_p.t813 vdd.t686 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X985 out_p.t489 vp_p.t814 vdd.t685 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X986 vdd.t684 vp_p.t815 out_p.t488 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X987 out_p.t1799 vp_n.t171 vss.t128 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X988 vdd.t683 vp_p.t816 out_p.t881 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X989 out_p.t1794 vp_n.t172 vss.t127 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X990 out_p.t880 vp_p.t817 vdd.t682 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X991 vdd.t681 vp_p.t818 out_p.t427 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X992 vdd.t680 vp_p.t819 out_p.t426 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X993 vdd.t679 vp_p.t820 out_p.t171 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X994 out_p.t170 vp_p.t821 vdd.t678 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X995 out_p.t1005 vp_p.t822 vdd.t677 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X996 vss.t126 vp_n.t173 out_p.t1795 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X997 out_p.t1004 vp_p.t823 vdd.t676 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X998 out_p.t679 vp_p.t824 vdd.t675 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X999 vdd.t674 vp_p.t825 out_p.t678 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1000 vdd.t673 vp_p.t826 out_p.t433 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1001 vdd.t672 vp_p.t827 out_p.t432 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1002 vdd.t671 vp_p.t828 out_p.t1019 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1003 out_p.t1018 vp_p.t829 vdd.t670 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1004 vdd.t669 vp_p.t830 out_p.t663 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1005 out_p.t662 vp_p.t831 vdd.t668 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1006 out_p.t615 vp_p.t832 vdd.t667 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1007 out_p.t614 vp_p.t833 vdd.t666 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1008 out_p.t1607 vp_p.t834 vdd.t665 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1009 out_p.t1606 vp_p.t835 vdd.t664 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1010 out_p.t152 vp_n.t174 vss.t125 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1011 vdd.t663 vp_p.t836 out_p.t929 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1012 out_p.t928 vp_p.t837 vdd.t662 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1013 vdd.t661 vp_p.t838 out_p.t251 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1014 out_p.t153 vp_n.t175 vss.t124 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1015 vdd.t660 vp_p.t839 out_p.t250 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1016 out_p.t1239 vp_p.t840 vdd.t659 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1017 out_p.t4 vp_n.t176 vss.t123 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1018 out_p.t1238 vp_p.t841 vdd.t658 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1019 vdd.t657 vp_p.t842 out_p.t1645 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1020 vdd.t656 vp_p.t843 out_p.t1644 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1021 vdd.t655 vp_p.t844 out_p.t709 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1022 out_p.t708 vp_p.t845 vdd.t654 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1023 vdd.t653 vp_p.t846 out_p.t1427 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1024 vdd.t652 vp_p.t847 out_p.t1426 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1025 vdd.t651 vp_p.t848 out_p.t1387 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1026 vdd.t650 vp_p.t849 out_p.t1386 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1027 vdd.t649 vp_p.t850 out_p.t1097 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1028 out_p.t5 vp_n.t177 vss.t122 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1029 out_p.t1096 vp_p.t851 vdd.t648 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1030 vss.t121 vp_n.t178 out_p.t10 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1031 vdd.t647 vp_p.t852 out_p.t819 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1032 out_p.t818 vp_p.t853 vdd.t646 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1033 vdd.t645 vp_p.t854 out_p.t1215 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1034 vdd.t644 vp_p.t855 out_p.t1214 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1035 out_p.t835 vp_p.t856 vdd.t643 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1036 vdd.t642 vp_p.t857 out_p.t834 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1037 out_p.t11 vp_n.t179 vss.t120 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1038 vdd.t641 vp_p.t858 out_p.t785 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1039 vdd.t640 vp_p.t859 out_p.t784 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1040 out_p.t971 vp_p.t860 vdd.t639 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1041 out_p.t970 vp_p.t861 vdd.t638 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1042 out_p.t1461 vp_p.t862 vdd.t637 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1043 vdd.t636 vp_p.t863 out_p.t1460 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1044 vdd.t635 vp_p.t864 out_p.t349 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1045 vdd.t634 vp_p.t865 out_p.t348 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1046 vdd.t633 vp_p.t866 out_p.t915 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1047 out_p.t914 vp_p.t867 vdd.t632 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1048 vdd.t631 vp_p.t868 out_p.t729 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1049 vdd.t630 vp_p.t869 out_p.t728 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1050 out_p.t1469 vp_p.t870 vdd.t629 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1051 out_p.t1468 vp_p.t871 vdd.t628 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1052 vdd.t627 vp_p.t872 out_p.t633 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1053 out_p.t632 vp_p.t873 vdd.t626 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1054 vss.t119 vp_n.t180 out_p.t120 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1055 out_p.t121 vp_n.t181 vss.t118 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1056 out_p.t1095 vp_p.t874 vdd.t625 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1057 vdd.t624 vp_p.t875 out_p.t1094 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1058 vdd.t623 vp_p.t876 out_p.t271 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1059 vdd.t622 vp_p.t877 out_p.t270 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1060 vss.t117 vp_n.t182 out_p.t8 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1061 out_p.t867 vp_p.t878 vdd.t621 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1062 out_p.t866 vp_p.t879 vdd.t620 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1063 vdd.t619 vp_p.t880 out_p.t765 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1064 out_p.t764 vp_p.t881 vdd.t618 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1065 out_p.t9 vp_n.t183 vss.t116 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1066 out_p.t1519 vp_p.t882 vdd.t617 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1067 out_p.t1518 vp_p.t883 vdd.t616 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1068 out_p.t619 vp_p.t884 vdd.t615 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1069 out_p.t12 vp_n.t184 vss.t115 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1070 vdd.t614 vp_p.t885 out_p.t618 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1071 vdd.t613 vp_p.t886 out_p.t1349 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1072 out_p.t13 vp_n.t185 vss.t114 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1073 vdd.t612 vp_p.t887 out_p.t1348 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1074 vdd.t611 vp_p.t888 out_p.t719 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1075 out_p.t40 vp_n.t186 vss.t113 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1076 out_p.t718 vp_p.t889 vdd.t610 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1077 out_p.t1135 vp_p.t890 vdd.t609 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1078 vdd.t608 vp_p.t891 out_p.t1134 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1079 out_p.t1209 vp_p.t892 vdd.t607 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1080 out_p.t1208 vp_p.t893 vdd.t606 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1081 out_p.t247 vp_p.t894 vdd.t605 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1082 out_p.t246 vp_p.t895 vdd.t604 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1083 out_p.t41 vp_n.t187 vss.t112 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1084 vdd.t603 vp_p.t896 out_p.t885 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1085 out_p.t884 vp_p.t897 vdd.t602 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1086 vdd.t601 vp_p.t898 out_p.t1195 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1087 vdd.t600 vp_p.t899 out_p.t1194 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1088 out_p.t1027 vp_p.t900 vdd.t599 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1089 out_p.t1026 vp_p.t901 vdd.t598 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1090 vdd.t597 vp_p.t902 out_p.t165 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1091 out_p.t164 vp_p.t903 vdd.t596 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1092 out_p.t148 vp_n.t188 vss.t111 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1093 vss.t110 vp_n.t189 out_p.t149 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1094 out_p.t501 vp_p.t904 vdd.t595 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1095 out_p.t500 vp_p.t905 vdd.t594 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1096 out_p.t50 vp_n.t190 vss.t109 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1097 out_p.t1297 vp_p.t906 vdd.t593 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1098 out_p.t1296 vp_p.t907 vdd.t592 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1099 vdd.t591 vp_p.t908 out_p.t1415 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1100 vss.t108 vp_n.t191 out_p.t51 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1101 vdd.t590 vp_p.t909 out_p.t1414 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1102 out_p.t1123 vp_p.t910 vdd.t589 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1103 out_p.t1122 vp_p.t911 vdd.t588 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1104 vdd.t587 vp_p.t912 out_p.t1503 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1105 vss.t107 vp_n.t192 out_p.t54 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1106 vdd.t586 vp_p.t913 out_p.t1502 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1107 vdd.t585 vp_p.t914 out_p.t823 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1108 out_p.t822 vp_p.t915 vdd.t584 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1109 vdd.t583 vp_p.t916 out_p.t1453 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1110 out_p.t55 vp_n.t193 vss.t106 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1111 vdd.t582 vp_p.t917 out_p.t1452 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1112 vdd.t581 vp_p.t918 out_p.t831 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1113 vdd.t580 vp_p.t919 out_p.t830 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1114 vdd.t579 vp_p.t920 out_p.t1309 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1115 vss.t105 vp_n.t194 out_p.t1770 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1116 out_p.t1308 vp_p.t921 vdd.t578 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1117 out_p.t907 vp_p.t922 vdd.t577 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1118 out_p.t906 vp_p.t923 vdd.t576 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1119 out_p.t259 vp_p.t924 vdd.t575 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1120 vdd.t574 vp_p.t925 out_p.t258 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1121 vdd.t573 vp_p.t926 out_p.t1565 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1122 out_p.t1564 vp_p.t927 vdd.t572 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1123 out_p.t1655 vp_p.t928 vdd.t571 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1124 vdd.t570 vp_p.t929 out_p.t1654 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1125 vdd.t569 vp_p.t930 out_p.t1431 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1126 out_p.t1430 vp_p.t931 vdd.t568 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1127 vdd.t567 vp_p.t932 out_p.t1317 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1128 out_p.t1316 vp_p.t933 vdd.t566 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1129 vdd.t565 vp_p.t934 out_p.t525 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1130 vdd.t564 vp_p.t935 out_p.t524 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1131 out_p.t1771 vp_n.t195 vss.t104 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1132 vdd.t563 vp_p.t936 out_p.t649 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1133 out_p.t648 vp_p.t937 vdd.t562 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1134 out_p.t1716 vp_n.t196 vss.t103 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1135 out_p.t1717 vp_n.t197 vss.t102 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1136 vdd.t561 vp_p.t938 out_p.t1537 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1137 vdd.t560 vp_p.t939 out_p.t1536 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1138 vdd.t559 vp_p.t940 out_p.t1219 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1139 vdd.t558 vp_p.t941 out_p.t1218 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1140 vdd.t557 vp_p.t942 out_p.t1007 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1141 vdd.t556 vp_p.t943 out_p.t1006 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1142 out_p.t465 vp_p.t944 vdd.t555 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1143 out_p.t464 vp_p.t945 vdd.t554 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1144 vdd.t553 vp_p.t946 out_p.t1521 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1145 vdd.t552 vp_p.t947 out_p.t1520 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1146 vdd.t551 vp_p.t948 out_p.t1001 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1147 vdd.t550 vp_p.t949 out_p.t1000 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1148 out_p.t903 vp_p.t950 vdd.t549 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1149 vdd.t548 vp_p.t951 out_p.t902 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1150 out_p.t110 vp_n.t198 vss.t101 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1151 out_p.t1169 vp_p.t952 vdd.t547 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1152 vdd.t546 vp_p.t953 out_p.t1168 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1153 out_p.t705 vp_p.t954 vdd.t545 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1154 out_p.t704 vp_p.t955 vdd.t544 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1155 out_p.t1633 vp_p.t956 vdd.t543 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1156 out_p.t1632 vp_p.t957 vdd.t542 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1157 vdd.t541 vp_p.t958 out_p.t977 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1158 out_p.t111 vp_n.t199 vss.t100 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1159 vdd.t540 vp_p.t959 out_p.t976 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1160 vdd.t539 vp_p.t960 out_p.t1271 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1161 vdd.t538 vp_p.t961 out_p.t1270 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1162 out_p.t1549 vp_p.t962 vdd.t537 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1163 out_p.t1548 vp_p.t963 vdd.t536 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1164 vdd.t535 vp_p.t964 out_p.t1355 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1165 out_p.t1354 vp_p.t965 vdd.t534 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1166 out_p.t447 vp_p.t966 vdd.t533 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1167 vdd.t532 vp_p.t967 out_p.t446 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1168 vdd.t531 vp_p.t968 out_p.t1203 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1169 vss.t99 vp_n.t200 out_p.t1686 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1170 out_p.t1202 vp_p.t969 vdd.t530 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1171 vdd.t529 vp_p.t970 out_p.t1619 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1172 vdd.t528 vp_p.t971 out_p.t1618 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1173 out_p.t1687 vp_n.t201 vss.t98 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1174 vss.t97 vp_n.t202 out_p.t114 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1175 out_p.t1081 vp_p.t972 vdd.t527 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1176 out_p.t1080 vp_p.t973 vdd.t526 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1177 out_p.t115 vp_n.t203 vss.t96 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1178 out_p.t1137 vp_p.t974 vdd.t525 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1179 vdd.t524 vp_p.t975 out_p.t1136 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1180 vdd.t523 vp_p.t976 out_p.t1199 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1181 out_p.t1198 vp_p.t977 vdd.t522 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1182 out_p.t1259 vp_p.t978 vdd.t521 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1183 out_p.t1258 vp_p.t979 vdd.t520 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1184 vdd.t519 vp_p.t980 out_p.t1079 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1185 vss.t95 vp_n.t204 out_p.t72 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1186 vdd.t518 vp_p.t981 out_p.t1078 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1187 vdd.t517 vp_p.t982 out_p.t845 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1188 out_p.t844 vp_p.t983 vdd.t516 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1189 vdd.t515 vp_p.t984 out_p.t603 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1190 vdd.t514 vp_p.t985 out_p.t602 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1191 vss.t94 vp_n.t205 out_p.t73 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1192 out_p.t329 vp_p.t986 vdd.t513 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1193 vdd.t512 vp_p.t987 out_p.t328 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1194 vdd.t511 vp_p.t988 out_p.t1377 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1195 out_p.t1376 vp_p.t989 vdd.t510 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1196 out_p.t56 vp_n.t206 vss.t93 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1197 out_p.t597 vp_p.t990 vdd.t509 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1198 out_p.t596 vp_p.t991 vdd.t508 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1199 out_p.t373 vp_p.t992 vdd.t507 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1200 out_p.t57 vp_n.t207 vss.t92 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1201 vss.t91 vp_n.t208 out_p.t104 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1202 vdd.t506 vp_p.t993 out_p.t372 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1203 vdd.t505 vp_p.t994 out_p.t1403 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1204 vss.t90 vp_n.t209 out_p.t105 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1205 out_p.t1402 vp_p.t995 vdd.t504 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1206 vdd.t503 vp_p.t996 out_p.t851 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1207 out_p.t850 vp_p.t997 vdd.t502 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1208 out_p.t1441 vp_p.t998 vdd.t501 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1209 vdd.t500 vp_p.t999 out_p.t1440 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1210 out_p.t1055 vp_p.t1000 vdd.t499 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1211 out_p.t1054 vp_p.t1001 vdd.t498 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1212 vdd.t497 vp_p.t1002 out_p.t1191 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1213 out_p.t1190 vp_p.t1003 vdd.t496 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1214 out_p.t1375 vp_p.t1004 vdd.t495 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1215 out_p.t1374 vp_p.t1005 vdd.t494 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1216 out_p.t1323 vp_p.t1006 vdd.t493 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1217 out_p.t1756 vp_n.t210 vss.t89 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1218 out_p.t1322 vp_p.t1007 vdd.t492 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1219 vdd.t491 vp_p.t1008 out_p.t1131 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1220 vdd.t490 vp_p.t1009 out_p.t1130 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1221 vss.t88 vp_n.t211 out_p.t1757 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1222 vdd.t489 vp_p.t1010 out_p.t577 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1223 vdd.t488 vp_p.t1011 out_p.t576 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1224 out_p.t1291 vp_p.t1012 vdd.t487 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1225 vdd.t486 vp_p.t1013 out_p.t1290 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1226 vdd.t485 vp_p.t1014 out_p.t1103 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1227 vss.t87 vp_n.t212 out_p.t1750 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1228 out_p.t1751 vp_n.t213 vss.t86 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1229 out_p.t1102 vp_p.t1015 vdd.t484 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1230 vss.t85 vp_n.t214 out_p.t1780 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1231 out_p.t307 vp_p.t1016 vdd.t483 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1232 out_p.t306 vp_p.t1017 vdd.t482 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1233 out_p.t509 vp_p.t1018 vdd.t481 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1234 out_p.t508 vp_p.t1019 vdd.t480 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1235 vdd.t479 vp_p.t1020 out_p.t791 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1236 out_p.t790 vp_p.t1021 vdd.t478 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1237 vdd.t477 vp_p.t1022 out_p.t429 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1238 out_p.t428 vp_p.t1023 vdd.t476 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1239 out_p.t205 vp_p.t1024 vdd.t475 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1240 vss.t84 vp_n.t215 out_p.t1781 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1241 out_p.t204 vp_p.t1025 vdd.t474 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1242 out_p.t1365 vp_p.t1026 vdd.t473 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1243 vdd.t472 vp_p.t1027 out_p.t1364 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1244 out_p.t837 vp_p.t1028 vdd.t471 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1245 vdd.t470 vp_p.t1029 out_p.t836 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1246 vdd.t469 vp_p.t1030 out_p.t549 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1247 vdd.t468 vp_p.t1031 out_p.t548 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1248 vdd.t467 vp_p.t1032 out_p.t1515 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1249 vss.t83 vp_n.t216 out_p.t124 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1250 vss.t82 vp_n.t217 out_p.t125 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1251 out_p.t1514 vp_p.t1033 vdd.t466 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1252 vdd.t465 vp_p.t1034 out_p.t183 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1253 out_p.t182 vp_p.t1035 vdd.t464 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1254 vss.t81 vp_n.t218 out_p.t132 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1255 vdd.t463 vp_p.t1036 out_p.t1463 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1256 vdd.t462 vp_p.t1037 out_p.t1462 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1257 out_p.t503 vp_p.t1038 vdd.t461 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1258 out_p.t502 vp_p.t1039 vdd.t460 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1259 out_p.t361 vp_p.t1040 vdd.t459 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1260 vdd.t458 vp_p.t1041 out_p.t360 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1261 vdd.t457 vp_p.t1042 out_p.t415 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1262 out_p.t414 vp_p.t1043 vdd.t456 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1263 vdd.t455 vp_p.t1044 out_p.t1177 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1264 out_p.t1176 vp_p.t1045 vdd.t454 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1265 out_p.t1609 vp_p.t1046 vdd.t453 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1266 out_p.t1608 vp_p.t1047 vdd.t452 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1267 out_p.t589 vp_p.t1048 vdd.t451 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1268 vss.t80 vp_n.t219 out_p.t133 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1269 out_p.t588 vp_p.t1049 vdd.t450 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1270 out_p.t1277 vp_p.t1050 vdd.t449 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1271 vdd.t448 vp_p.t1051 out_p.t1276 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1272 vdd.t447 vp_p.t1052 out_p.t673 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1273 out_p.t136 vp_n.t220 vss.t79 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1274 out_p.t672 vp_p.t1053 vdd.t446 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1275 out_p.t417 vp_p.t1054 vdd.t445 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1276 vdd.t444 vp_p.t1055 out_p.t416 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1277 out_p.t841 vp_p.t1056 vdd.t443 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1278 vdd.t442 vp_p.t1057 out_p.t840 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1279 out_p.t1221 vp_p.t1058 vdd.t441 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1280 vdd.t440 vp_p.t1059 out_p.t1220 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1281 vss.t78 vp_n.t221 out_p.t137 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1282 out_p.t187 vp_p.t1060 vdd.t439 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1283 out_p.t186 vp_p.t1061 vdd.t438 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1284 vdd.t437 vp_p.t1062 out_p.t1129 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1285 vdd.t436 vp_p.t1063 out_p.t1128 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1286 vdd.t435 vp_p.t1064 out_p.t245 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1287 out_p.t244 vp_p.t1065 vdd.t434 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1288 out_p.t1433 vp_p.t1066 vdd.t433 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1289 vdd.t432 vp_p.t1067 out_p.t1432 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1290 vdd.t431 vp_p.t1068 out_p.t803 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1291 out_p.t802 vp_p.t1069 vdd.t430 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1292 out_p.t843 vp_p.t1070 vdd.t429 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1293 vdd.t428 vp_p.t1071 out_p.t842 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1294 out_p.t315 vp_p.t1072 vdd.t427 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1295 out_p.t314 vp_p.t1073 vdd.t426 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1296 out_p.t303 vp_p.t1074 vdd.t425 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1297 vdd.t424 vp_p.t1075 out_p.t302 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1298 vdd.t423 vp_p.t1076 out_p.t1629 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1299 vdd.t422 vp_p.t1077 out_p.t1628 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1300 out_p.t140 vp_n.t222 vss.t77 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1301 vdd.t421 vp_p.t1078 out_p.t755 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1302 out_p.t141 vp_n.t223 vss.t76 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1303 vss.t75 vp_n.t224 out_p.t76 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1304 vdd.t420 vp_p.t1079 out_p.t754 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1305 out_p.t677 vp_p.t1080 vdd.t419 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1306 out_p.t676 vp_p.t1081 vdd.t418 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1307 out_p.t235 vp_p.t1082 vdd.t417 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1308 out_p.t234 vp_p.t1083 vdd.t416 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1309 vdd.t415 vp_p.t1084 out_p.t1313 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1310 vss.t74 vp_n.t225 out_p.t77 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1311 vdd.t414 vp_p.t1085 out_p.t1312 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1312 out_p.t959 vp_p.t1086 vdd.t413 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1313 vdd.t412 vp_p.t1087 out_p.t958 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1314 out_p.t993 vp_p.t1088 vdd.t411 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1315 vss.t73 vp_n.t226 out_p.t14 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1316 out_p.t992 vp_p.t1089 vdd.t410 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1317 vdd.t409 vp_p.t1090 out_p.t301 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1318 vdd.t408 vp_p.t1091 out_p.t300 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1319 vdd.t407 vp_p.t1092 out_p.t1507 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1320 vdd.t406 vp_p.t1093 out_p.t1506 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1321 out_p.t225 vp_p.t1094 vdd.t405 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1322 out_p.t224 vp_p.t1095 vdd.t404 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1323 out_p.t1167 vp_p.t1096 vdd.t403 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1324 vss.t72 vp_n.t227 out_p.t15 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1325 out_p.t1166 vp_p.t1097 vdd.t402 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1326 vss.t71 vp_n.t228 out_p.t80 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1327 out_p.t227 vp_p.t1098 vdd.t401 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1328 out_p.t226 vp_p.t1099 vdd.t400 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1329 out_p.t607 vp_p.t1100 vdd.t399 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1330 out_p.t606 vp_p.t1101 vdd.t398 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1331 vdd.t397 vp_p.t1102 out_p.t385 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1332 vdd.t396 vp_p.t1103 out_p.t384 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1333 vdd.t395 vp_p.t1104 out_p.t735 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1334 out_p.t734 vp_p.t1105 vdd.t394 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1335 vdd.t393 vp_p.t1106 out_p.t351 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1336 out_p.t350 vp_p.t1107 vdd.t392 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1337 vdd.t391 vp_p.t1108 out_p.t533 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1338 out_p.t532 vp_p.t1109 vdd.t390 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1339 out_p.t873 vp_p.t1110 vdd.t389 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1340 vdd.t388 vp_p.t1111 out_p.t872 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1341 out_p.t249 vp_p.t1112 vdd.t387 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1342 vdd.t386 vp_p.t1113 out_p.t248 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1343 vss.t70 vp_n.t229 out_p.t81 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1344 out_p.t1792 vp_n.t230 vss.t69 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1345 vdd.t385 vp_p.t1114 out_p.t695 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1346 vss.t68 vp_n.t231 out_p.t1793 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1347 vdd.t384 vp_p.t1115 out_p.t694 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1348 vdd.t383 vp_p.t1116 out_p.t1329 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1349 out_p.t1328 vp_p.t1117 vdd.t382 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1350 out_p.t1746 vp_n.t232 vss.t67 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1351 out_p.t981 vp_p.t1118 vdd.t381 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1352 out_p.t980 vp_p.t1119 vdd.t380 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1353 vdd.t379 vp_p.t1120 out_p.t1279 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1354 vdd.t378 vp_p.t1121 out_p.t1278 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1355 out_p.t1087 vp_p.t1122 vdd.t377 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1356 vdd.t376 vp_p.t1123 out_p.t1086 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1357 vdd.t375 vp_p.t1124 out_p.t497 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1358 out_p.t1747 vp_n.t233 vss.t66 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1359 out_p.t496 vp_p.t1125 vdd.t374 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1360 out_p.t1071 vp_p.t1126 vdd.t373 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1361 out_p.t1070 vp_p.t1127 vdd.t372 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1362 out_p.t1587 vp_p.t1128 vdd.t371 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1363 out_p.t1586 vp_p.t1129 vdd.t370 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1364 out_p.t1197 vp_p.t1130 vdd.t369 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1365 out_p.t1762 vp_n.t234 vss.t65 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1366 vdd.t368 vp_p.t1131 out_p.t1196 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1367 vdd.t367 vp_p.t1132 out_p.t1049 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1368 vdd.t366 vp_p.t1133 out_p.t1048 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1369 out_p.t711 vp_p.t1134 vdd.t365 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1370 out_p.t710 vp_p.t1135 vdd.t364 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1371 out_p.t707 vp_p.t1136 vdd.t363 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1372 vdd.t362 vp_p.t1137 out_p.t706 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1373 out_p.t1513 vp_p.t1138 vdd.t361 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1374 vdd.t360 vp_p.t1139 out_p.t1512 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1375 out_p.t1247 vp_p.t1140 vdd.t359 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1376 vss.t64 vp_n.t235 out_p.t1763 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1377 out_p.t1246 vp_p.t1141 vdd.t358 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1378 vss.t63 vp_n.t236 out_p.t58 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1379 vdd.t357 vp_p.t1142 out_p.t453 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1380 out_p.t452 vp_p.t1143 vdd.t356 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1381 out_p.t551 vp_p.t1144 vdd.t355 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1382 out_p.t550 vp_p.t1145 vdd.t354 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1383 out_p.t891 vp_p.t1146 vdd.t353 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1384 vdd.t352 vp_p.t1147 out_p.t890 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1385 out_p.t1351 vp_p.t1148 vdd.t351 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1386 vdd.t350 vp_p.t1149 out_p.t1350 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1387 out_p.t1151 vp_p.t1150 vdd.t349 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1388 out_p.t1150 vp_p.t1151 vdd.t348 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1389 out_p.t507 vp_p.t1152 vdd.t347 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1390 vdd.t346 vp_p.t1153 out_p.t506 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1391 out_p.t201 vp_p.t1154 vdd.t345 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1392 vss.t62 vp_n.t237 out_p.t59 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1393 vdd.t344 vp_p.t1155 out_p.t200 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1394 out_p.t309 vp_p.t1156 vdd.t343 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1395 vdd.t342 vp_p.t1157 out_p.t308 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1396 vdd.t341 vp_p.t1158 out_p.t1501 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1397 vdd.t340 vp_p.t1159 out_p.t1500 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1398 vdd.t339 vp_p.t1160 out_p.t397 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1399 out_p.t396 vp_p.t1161 vdd.t338 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1400 vdd.t337 vp_p.t1162 out_p.t193 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1401 out_p.t192 vp_p.t1163 vdd.t336 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1402 out_p.t1583 vp_p.t1164 vdd.t335 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1403 vdd.t334 vp_p.t1165 out_p.t1582 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1404 vdd.t333 vp_p.t1166 out_p.t269 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1405 out_p.t268 vp_p.t1167 vdd.t332 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1406 out_p.t1649 vp_p.t1168 vdd.t331 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1407 vdd.t330 vp_p.t1169 out_p.t1648 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1408 out_p.t1395 vp_p.t1170 vdd.t329 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1409 out_p.t52 vp_n.t238 vss.t61 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1410 out_p.t1394 vp_p.t1171 vdd.t328 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1411 vdd.t327 vp_p.t1172 out_p.t347 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1412 out_p.t346 vp_p.t1173 vdd.t326 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1413 out_p.t53 vp_n.t239 vss.t60 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1414 vss.t59 vp_n.t240 out_p.t1660 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1415 vdd.t325 vp_p.t1174 out_p.t531 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1416 vdd.t324 vp_p.t1175 out_p.t530 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1417 vdd.t323 vp_p.t1176 out_p.t773 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1418 vdd.t322 vp_p.t1177 out_p.t772 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1419 out_p.t1265 vp_p.t1178 vdd.t321 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1420 vdd.t320 vp_p.t1179 out_p.t1264 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1421 out_p.t319 vp_p.t1180 vdd.t319 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1422 out_p.t1661 vp_n.t241 vss.t58 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1423 vdd.t318 vp_p.t1181 out_p.t318 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1424 out_p.t775 vp_p.t1182 vdd.t317 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1425 vdd.t316 vp_p.t1183 out_p.t774 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1426 vdd.t315 vp_p.t1184 out_p.t975 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1427 out_p.t1732 vp_n.t242 vss.t57 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1428 vdd.t314 vp_p.t1185 out_p.t974 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1429 out_p.t825 vp_p.t1186 vdd.t313 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1430 out_p.t824 vp_p.t1187 vdd.t312 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1431 vss.t56 vp_n.t243 out_p.t1733 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1432 out_p.t529 vp_p.t1188 vdd.t311 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1433 out_p.t528 vp_p.t1189 vdd.t310 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1434 vdd.t309 vp_p.t1190 out_p.t961 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1435 vdd.t308 vp_p.t1191 out_p.t960 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1436 out_p.t613 vp_p.t1192 vdd.t307 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1437 out_p.t612 vp_p.t1193 vdd.t306 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1438 vdd.t305 vp_p.t1194 out_p.t1111 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1439 vdd.t304 vp_p.t1195 out_p.t1110 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1440 vdd.t303 vp_p.t1196 out_p.t1043 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1441 vdd.t302 vp_p.t1197 out_p.t1042 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1442 vss.t55 vp_n.t244 out_p.t144 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1443 vdd.t301 vp_p.t1198 out_p.t405 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1444 vdd.t300 vp_p.t1199 out_p.t404 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1445 out_p.t287 vp_p.t1200 vdd.t299 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1446 vdd.t298 vp_p.t1201 out_p.t286 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1447 vdd.t297 vp_p.t1202 out_p.t1381 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1448 out_p.t145 vp_n.t245 vss.t54 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1449 vdd.t296 vp_p.t1203 out_p.t1380 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1450 vdd.t295 vp_p.t1204 out_p.t1411 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1451 out_p.t1410 vp_p.t1205 vdd.t294 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1452 out_p.t1147 vp_p.t1206 vdd.t293 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1453 out_p.t92 vp_n.t246 vss.t53 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1454 vdd.t292 vp_p.t1207 out_p.t1146 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1455 out_p.t1621 vp_p.t1208 vdd.t291 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1456 vdd.t290 vp_p.t1209 out_p.t1620 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1457 out_p.t1115 vp_p.t1210 vdd.t289 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1458 vdd.t288 vp_p.t1211 out_p.t1114 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1459 vdd.t287 vp_p.t1212 out_p.t1157 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1460 vdd.t286 vp_p.t1213 out_p.t1156 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1461 out_p.t537 vp_p.t1214 vdd.t285 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1462 vdd.t284 vp_p.t1215 out_p.t536 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1463 vdd.t283 vp_p.t1216 out_p.t947 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1464 out_p.t946 vp_p.t1217 vdd.t282 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1465 vdd.t281 vp_p.t1218 out_p.t1255 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1466 vss.t52 vp_n.t247 out_p.t93 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1467 vdd.t280 vp_p.t1219 out_p.t1254 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1468 vdd.t279 vp_p.t1220 out_p.t949 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1469 vdd.t278 vp_p.t1221 out_p.t948 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1470 out_p.t1738 vp_n.t248 vss.t51 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1471 out_p.t849 vp_p.t1222 vdd.t277 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1472 out_p.t1739 vp_n.t249 vss.t50 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1473 vdd.t276 vp_p.t1223 out_p.t848 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1474 out_p.t1153 vp_p.t1224 vdd.t275 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1475 vdd.t274 vp_p.t1225 out_p.t1152 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1476 vss.t49 vp_n.t250 out_p.t1734 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1477 out_p.t203 vp_p.t1226 vdd.t273 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1478 vdd.t272 vp_p.t1227 out_p.t202 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1479 out_p.t1315 vp_p.t1228 vdd.t271 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1480 vss.t48 vp_n.t251 out_p.t1735 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1481 vdd.t270 vp_p.t1229 out_p.t1314 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1482 out_p.t88 vp_n.t252 vss.t47 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1483 out_p.t1289 vp_p.t1230 vdd.t269 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1484 vdd.t268 vp_p.t1231 out_p.t1288 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1485 vdd.t267 vp_p.t1232 out_p.t889 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1486 vdd.t266 vp_p.t1233 out_p.t888 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1487 vdd.t265 vp_p.t1234 out_p.t561 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1488 vdd.t264 vp_p.t1235 out_p.t560 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1489 out_p.t445 vp_p.t1236 vdd.t263 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1490 vdd.t262 vp_p.t1237 out_p.t444 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1491 out_p.t89 vp_n.t253 vss.t46 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1492 out_p.t935 vp_p.t1238 vdd.t261 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1493 vdd.t260 vp_p.t1239 out_p.t934 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1494 out_p.t743 vp_p.t1240 vdd.t259 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1495 vdd.t258 vp_p.t1241 out_p.t742 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1496 vdd.t257 vp_p.t1242 out_p.t795 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1497 vdd.t256 vp_p.t1243 out_p.t794 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1498 out_p.t757 vp_p.t1244 vdd.t255 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1499 out_p.t756 vp_p.t1245 vdd.t254 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1500 out_p.t671 vp_p.t1246 vdd.t253 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1501 out_p.t1742 vp_n.t254 vss.t45 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1502 out_p.t1743 vp_n.t255 vss.t44 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1503 vdd.t252 vp_p.t1247 out_p.t670 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1504 vdd.t251 vp_p.t1248 out_p.t1625 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1505 out_p.t1624 vp_p.t1249 vdd.t250 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1506 out_p.t64 vp_n.t256 vss.t43 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1507 out_p.t769 vp_p.t1250 vdd.t249 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1508 out_p.t768 vp_p.t1251 vdd.t248 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1509 vdd.t247 vp_p.t1252 out_p.t1471 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1510 vdd.t246 vp_p.t1253 out_p.t1470 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1511 out_p.t593 vp_p.t1254 vdd.t245 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1512 out_p.t592 vp_p.t1255 vdd.t244 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1513 vdd.t243 vp_p.t1256 out_p.t1041 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1514 out_p.t1040 vp_p.t1257 vdd.t242 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1515 vss.t42 vp_n.t257 out_p.t65 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1516 vdd.t241 vp_p.t1258 out_p.t759 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1517 vdd.t240 vp_p.t1259 out_p.t758 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1518 vdd.t239 vp_p.t1260 out_p.t365 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1519 out_p.t90 vp_n.t258 vss.t41 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1520 vdd.t238 vp_p.t1261 out_p.t364 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1521 out_p.t875 vp_p.t1262 vdd.t237 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1522 out_p.t874 vp_p.t1263 vdd.t236 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1523 vdd.t235 vp_p.t1264 out_p.t909 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1524 vss.t40 vp_n.t259 out_p.t91 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1525 vdd.t234 vp_p.t1265 out_p.t908 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1526 vss.t39 vp_n.t260 out_p.t96 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1527 vdd.t233 vp_p.t1266 out_p.t1483 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1528 out_p.t1482 vp_p.t1267 vdd.t232 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1529 out_p.t313 vp_p.t1268 vdd.t231 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1530 vdd.t230 vp_p.t1269 out_p.t312 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1531 vdd.t229 vp_p.t1270 out_p.t1627 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1532 out_p.t1626 vp_p.t1271 vdd.t228 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1533 vdd.t227 vp_p.t1272 out_p.t1393 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1534 vdd.t226 vp_p.t1273 out_p.t1392 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1535 out_p.t1237 vp_p.t1274 vdd.t225 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1536 out_p.t1236 vp_p.t1275 vdd.t224 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1537 vdd.t223 vp_p.t1276 out_p.t327 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1538 vdd.t222 vp_p.t1277 out_p.t326 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1539 out_p.t1205 vp_p.t1278 vdd.t221 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1540 out_p.t1204 vp_p.t1279 vdd.t220 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1541 vdd.t219 vp_p.t1280 out_p.t1389 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1542 vdd.t218 vp_p.t1281 out_p.t1388 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1543 vdd.t217 vp_p.t1282 out_p.t1267 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1544 vdd.t216 vp_p.t1283 out_p.t1266 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1545 vdd.t215 vp_p.t1284 out_p.t391 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1546 out_p.t390 vp_p.t1285 vdd.t214 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1547 out_p.t1595 vp_p.t1286 vdd.t213 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1548 out_p.t1594 vp_p.t1287 vdd.t212 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1549 out_p.t893 vp_p.t1288 vdd.t211 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1550 vss.t38 vp_n.t261 out_p.t97 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1551 out_p.t1758 vp_n.t262 vss.t37 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1552 out_p.t892 vp_p.t1289 vdd.t210 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1553 vdd.t209 vp_p.t1290 out_p.t901 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1554 vdd.t208 vp_p.t1291 out_p.t900 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1555 out_p.t1249 vp_p.t1292 vdd.t207 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1556 out_p.t1759 vp_n.t263 vss.t36 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1557 out_p.t1248 vp_p.t1293 vdd.t206 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1558 vdd.t205 vp_p.t1294 out_p.t1397 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1559 out_p.t1396 vp_p.t1295 vdd.t204 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1560 vdd.t203 vp_p.t1296 out_p.t1653 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1561 out_p.t1790 vp_n.t264 vss.t35 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1562 vdd.t202 vp_p.t1297 out_p.t1652 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1563 out_p.t887 vp_p.t1298 vdd.t201 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1564 out_p.t886 vp_p.t1299 vdd.t200 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1565 out_p.t353 vp_p.t1300 vdd.t199 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1566 vdd.t198 vp_p.t1301 out_p.t352 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1567 out_p.t829 vp_p.t1302 vdd.t197 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1568 out_p.t828 vp_p.t1303 vdd.t196 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1569 vdd.t195 vp_p.t1304 out_p.t317 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1570 out_p.t1791 vp_n.t265 vss.t34 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1571 vdd.t194 vp_p.t1305 out_p.t316 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1572 out_p.t1754 vp_n.t266 vss.t33 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1573 vdd.t193 vp_p.t1306 out_p.t641 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1574 vdd.t192 vp_p.t1307 out_p.t640 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1575 out_p.t699 vp_p.t1308 vdd.t191 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1576 out_p.t698 vp_p.t1309 vdd.t190 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1577 out_p.t197 vp_p.t1310 vdd.t189 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1578 vdd.t188 vp_p.t1311 out_p.t196 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1579 out_p.t1285 vp_p.t1312 vdd.t187 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1580 out_p.t1284 vp_p.t1313 vdd.t186 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1581 out_p.t605 vp_p.t1314 vdd.t185 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1582 vdd.t184 vp_p.t1315 out_p.t604 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1583 vdd.t183 vp_p.t1316 out_p.t1467 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1584 vss.t32 vp_n.t267 out_p.t1755 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1585 out_p.t1466 vp_p.t1317 vdd.t182 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1586 out_p.t495 vp_p.t1318 vdd.t181 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1587 vdd.t180 vp_p.t1319 out_p.t494 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1588 out_p.t20 vp_n.t268 vss.t31 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1589 vss.t30 vp_n.t269 out_p.t21 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1590 out_p.t331 vp_p.t1320 vdd.t179 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1591 vss.t29 vp_n.t270 out_p.t98 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1592 out_p.t330 vp_p.t1321 vdd.t178 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1593 vdd.t177 vp_p.t1322 out_p.t1305 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1594 out_p.t1304 vp_p.t1323 vdd.t176 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1595 vdd.t175 vp_p.t1324 out_p.t905 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1596 vdd.t174 vp_p.t1325 out_p.t904 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1597 out_p.t1613 vp_p.t1326 vdd.t173 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1598 vdd.t172 vp_p.t1327 out_p.t1612 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1599 out_p.t335 vp_p.t1328 vdd.t171 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1600 out_p.t334 vp_p.t1329 vdd.t170 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1601 vdd.t169 vp_p.t1330 out_p.t379 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1602 vss.t28 vp_n.t271 out_p.t99 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1603 vss.t27 vp_n.t272 out_p.t1696 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1604 out_p.t378 vp_p.t1331 vdd.t168 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1605 vdd.t167 vp_p.t1332 out_p.t1009 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1606 vdd.t166 vp_p.t1333 out_p.t1008 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1607 vdd.t165 vp_p.t1334 out_p.t1435 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1608 vdd.t164 vp_p.t1335 out_p.t1434 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1609 out_p.t487 vp_p.t1336 vdd.t163 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1610 out_p.t486 vp_p.t1337 vdd.t162 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1611 vdd.t161 vp_p.t1338 out_p.t855 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1612 out_p.t854 vp_p.t1339 vdd.t160 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1613 out_p.t1499 vp_p.t1340 vdd.t159 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1614 out_p.t1498 vp_p.t1341 vdd.t158 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1615 out_p.t279 vp_p.t1342 vdd.t157 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1616 out_p.t1697 vp_n.t273 vss.t26 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1617 out_p.t1664 vp_n.t274 vss.t25 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1618 out_p.t278 vp_p.t1343 vdd.t156 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1619 vdd.t155 vp_p.t1344 out_p.t897 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1620 vss.t24 vp_n.t275 out_p.t1665 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1621 vdd.t154 vp_p.t1345 out_p.t896 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1622 vdd.t153 vp_p.t1346 out_p.t739 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1623 vdd.t152 vp_p.t1347 out_p.t738 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1624 vdd.t151 vp_p.t1348 out_p.t1141 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1625 out_p.t1140 vp_p.t1349 vdd.t150 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1626 out_p.t1179 vp_p.t1350 vdd.t149 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1627 out_p.t1178 vp_p.t1351 vdd.t148 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1628 vdd.t147 vp_p.t1352 out_p.t1117 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1629 vdd.t146 vp_p.t1353 out_p.t1116 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1630 out_p.t191 vp_p.t1354 vdd.t145 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1631 vdd.t144 vp_p.t1355 out_p.t190 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1632 out_p.t1676 vp_n.t276 vss.t23 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1633 out_p.t403 vp_p.t1356 vdd.t143 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1634 vdd.t142 vp_p.t1357 out_p.t402 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1635 vdd.t141 vp_p.t1358 out_p.t177 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1636 out_p.t176 vp_p.t1359 vdd.t140 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1637 out_p.t861 vp_p.t1360 vdd.t139 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1638 out_p.t860 vp_p.t1361 vdd.t138 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1639 out_p.t1399 vp_p.t1362 vdd.t137 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1640 vdd.t136 vp_p.t1363 out_p.t1398 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1641 out_p.t1013 vp_p.t1364 vdd.t135 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1642 vdd.t134 vp_p.t1365 out_p.t1012 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1643 vdd.t133 vp_p.t1366 out_p.t1479 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1644 out_p.t1478 vp_p.t1367 vdd.t132 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1645 vss.t22 vp_n.t277 out_p.t1677 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1646 vss.t21 vp_n.t278 out_p.t66 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1647 out_p.t973 vp_p.t1368 vdd.t131 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1648 vdd.t130 vp_p.t1369 out_p.t972 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1649 out_p.t1443 vp_p.t1370 vdd.t129 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1650 vdd.t128 vp_p.t1371 out_p.t1442 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1651 out_p.t67 vp_n.t279 vss.t20 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1652 vdd.t127 vp_p.t1372 out_p.t1161 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1653 out_p.t1160 vp_p.t1373 vdd.t126 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1654 out_p.t1421 vp_p.t1374 vdd.t125 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1655 out_p.t1420 vp_p.t1375 vdd.t124 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1656 out_p.t1641 vp_p.t1376 vdd.t123 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1657 out_p.t1640 vp_p.t1377 vdd.t122 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1658 out_p.t883 vp_p.t1378 vdd.t121 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1659 vdd.t120 vp_p.t1379 out_p.t882 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1660 vdd.t119 vp_p.t1380 out_p.t1429 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1661 vss.t19 vp_n.t280 out_p.t1688 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1662 vdd.t118 vp_p.t1381 out_p.t1428 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1663 vdd.t117 vp_p.t1382 out_p.t1447 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1664 out_p.t1446 vp_p.t1383 vdd.t116 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1665 out_p.t1419 vp_p.t1384 vdd.t115 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1666 out_p.t1418 vp_p.t1385 vdd.t114 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1667 out_p.t723 vp_p.t1386 vdd.t113 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1668 vss.t18 vp_n.t281 out_p.t1689 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1669 out_p.t722 vp_p.t1387 vdd.t112 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1670 vdd.t111 vp_p.t1388 out_p.t479 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1671 vdd.t110 vp_p.t1389 out_p.t478 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1672 vdd.t109 vp_p.t1390 out_p.t1021 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1673 out_p.t1020 vp_p.t1391 vdd.t108 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1674 out_p.t617 vp_p.t1392 vdd.t107 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1675 vdd.t106 vp_p.t1393 out_p.t616 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1676 out_p.t321 vp_p.t1394 vdd.t105 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1677 vdd.t104 vp_p.t1395 out_p.t320 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1678 vdd.t103 vp_p.t1396 out_p.t585 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1679 out_p.t584 vp_p.t1397 vdd.t102 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1680 out_p.t333 vp_p.t1398 vdd.t101 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1681 out_p.t332 vp_p.t1399 vdd.t100 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1682 vdd.t99 vp_p.t1400 out_p.t647 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1683 out_p.t44 vp_n.t282 vss.t17 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1684 vdd.t98 vp_p.t1401 out_p.t646 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1685 out_p.t289 vp_p.t1402 vdd.t97 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1686 out_p.t45 vp_n.t283 vss.t16 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1687 vdd.t96 vp_p.t1403 out_p.t288 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1688 out_p.t1233 vp_p.t1404 vdd.t95 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1689 out_p.t1232 vp_p.t1405 vdd.t94 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1690 out_p.t1145 vp_p.t1406 vdd.t93 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1691 vss.t15 vp_n.t284 out_p.t60 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1692 out_p.t1144 vp_p.t1407 vdd.t92 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1693 out_p.t467 vp_p.t1408 vdd.t91 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1694 vdd.t90 vp_p.t1409 out_p.t466 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1695 vdd.t89 vp_p.t1410 out_p.t1423 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1696 vdd.t88 vp_p.t1411 out_p.t1422 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1697 vdd.t87 vp_p.t1412 out_p.t1631 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1698 out_p.t1630 vp_p.t1413 vdd.t86 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1699 out_p.t1273 vp_p.t1414 vdd.t85 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1700 vdd.t84 vp_p.t1415 out_p.t1272 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1701 out_p.t1261 vp_p.t1416 vdd.t83 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1702 out_p.t1260 vp_p.t1417 vdd.t82 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1703 vdd.t81 vp_p.t1418 out_p.t1611 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1704 out_p.t1610 vp_p.t1419 vdd.t80 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1705 out_p.t789 vp_p.t1420 vdd.t79 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1706 out_p.t788 vp_p.t1421 vdd.t78 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1707 vdd.t77 vp_p.t1422 out_p.t927 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1708 out_p.t926 vp_p.t1423 vdd.t76 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1709 out_p.t169 vp_p.t1424 vdd.t75 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1710 out_p.t61 vp_n.t285 vss.t14 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1711 out_p.t168 vp_p.t1425 vdd.t74 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1712 out_p.t1557 vp_p.t1426 vdd.t73 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1713 out_p.t1556 vp_p.t1427 vdd.t72 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1714 vdd.t71 vp_p.t1428 out_p.t1569 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1715 vss.t13 vp_n.t286 out_p.t1776 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1716 vdd.t70 vp_p.t1429 out_p.t1568 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1717 vdd.t69 vp_p.t1430 out_p.t987 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1718 vdd.t68 vp_p.t1431 out_p.t986 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1719 vdd.t67 vp_p.t1432 out_p.t563 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1720 out_p.t562 vp_p.t1433 vdd.t66 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1721 vdd.t65 vp_p.t1434 out_p.t1121 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1722 out_p.t1120 vp_p.t1435 vdd.t64 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1723 vdd.t63 vp_p.t1436 out_p.t555 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1724 vdd.t62 vp_p.t1437 out_p.t554 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1725 out_p.t635 vp_p.t1438 vdd.t61 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1726 out_p.t1777 vp_n.t287 vss.t12 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1727 vdd.t60 vp_p.t1439 out_p.t634 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1728 vdd.t59 vp_p.t1440 out_p.t1113 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1729 vdd.t58 vp_p.t1441 out_p.t1112 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1730 vss.t11 vp_n.t288 out_p.t154 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1731 out_p.t715 vp_p.t1442 vdd.t57 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1732 out_p.t714 vp_p.t1443 vdd.t56 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1733 out_p.t399 vp_p.t1444 vdd.t55 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1734 out_p.t398 vp_p.t1445 vdd.t54 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1735 vdd.t53 vp_p.t1446 out_p.t277 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1736 vdd.t52 vp_p.t1447 out_p.t276 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1737 vss.t10 vp_n.t289 out_p.t155 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1738 vdd.t51 vp_p.t1448 out_p.t659 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1739 vdd.t50 vp_p.t1449 out_p.t658 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1740 out_p.t727 vp_p.t1450 vdd.t49 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1741 out_p.t726 vp_p.t1451 vdd.t48 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1742 out_p.t1173 vp_p.t1452 vdd.t47 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1743 out_p.t1172 vp_p.t1453 vdd.t46 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1744 out_p.t70 vp_n.t290 vss.t9 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1745 vdd.t45 vp_p.t1454 out_p.t477 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1746 vdd.t44 vp_p.t1455 out_p.t476 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1747 vdd.t43 vp_p.t1456 out_p.t499 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1748 vss.t8 vp_n.t291 out_p.t71 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1749 vss.t7 vp_n.t292 out_p.t1704 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1750 out_p.t498 vp_p.t1457 vdd.t42 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1751 out_p.t1559 vp_p.t1458 vdd.t41 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1752 vdd.t40 vp_p.t1459 out_p.t1558 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1753 vdd.t39 vp_p.t1460 out_p.t1171 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1754 out_p.t1170 vp_p.t1461 vdd.t38 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1755 out_p.t1539 vp_p.t1462 vdd.t37 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1756 vdd.t36 vp_p.t1463 out_p.t1538 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1757 out_p.t1235 vp_p.t1464 vdd.t35 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1758 vdd.t34 vp_p.t1465 out_p.t1234 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1759 vdd.t33 vp_p.t1466 out_p.t1425 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1760 out_p.t1705 vp_n.t293 vss.t6 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1761 out_p.t1424 vp_p.t1467 vdd.t32 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1762 vdd.t31 vp_p.t1468 out_p.t733 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1763 out_p.t732 vp_p.t1469 vdd.t30 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1764 out_p.t1143 vp_p.t1470 vdd.t29 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1765 vss.t5 vp_n.t294 out_p.t1698 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1766 out_p.t1142 vp_p.t1471 vdd.t28 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1767 vdd.t27 vp_p.t1472 out_p.t325 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1768 vdd.t26 vp_p.t1473 out_p.t324 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1769 out_p.t811 vp_p.t1474 vdd.t25 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1770 out_p.t810 vp_p.t1475 vdd.t24 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1771 out_p.t1699 vp_n.t295 vss.t4 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1772 out_p.t787 vp_p.t1476 vdd.t23 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1773 out_p.t786 vp_p.t1477 vdd.t22 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1774 out_p.t6 vp_n.t296 vss.t3 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1775 out_p.t163 vp_p.t1478 vdd.t21 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1776 vdd.t20 vp_p.t1479 out_p.t162 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1777 vdd.t19 vp_p.t1480 out_p.t1063 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1778 out_p.t1062 vp_p.t1481 vdd.t18 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1779 vdd.t17 vp_p.t1482 out_p.t1543 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1780 vdd.t16 vp_p.t1483 out_p.t1542 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1781 out_p.t1139 vp_p.t1484 vdd.t15 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1782 vdd.t14 vp_p.t1485 out_p.t1138 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1783 out_p.t1345 vp_p.t1486 vdd.t13 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1784 out_p.t1344 vp_p.t1487 vdd.t12 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1785 vdd.t11 vp_p.t1488 out_p.t411 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1786 vdd.t10 vp_p.t1489 out_p.t410 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1787 out_p.t553 vp_p.t1490 vdd.t9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1788 out_p.t552 vp_p.t1491 vdd.t8 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1789 vdd.t7 vp_p.t1492 out_p.t925 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1790 out_p.t924 vp_p.t1493 vdd.t6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1791 out_p.t158 vp_p.t1494 vdd.t5 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1792 vdd.t4 vp_p.t1495 out_p.t161 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1793 out_p.t156 vp_p.t1496 vdd.t3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1794 vdd.t2 vp_p.t1497 out_p.t157 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1795 out_p.t7 vp_n.t297 vss.t2 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1796 vss.t1 vp_n.t298 out_p.t1712 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1797 out_p.t160 vp_p.t1498 vdd.t1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1798 vdd.t0 vp_p.t1499 out_p.t159 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1799 vss.t0 vp_n.t299 out_p.t1713 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
C0 vdd out_p 4414.79fF
C1 vp_n out_p 102.35fF
C2 vdd vp_p 620.90fF
C3 out_p vp_p 548.19fF
R0 vp_p.n668 vp_p.t1456 756.008
R1 vp_p.n668 vp_p.t1242 756.008
R2 vp_p.n666 vp_p.t370 756.008
R3 vp_p.n666 vp_p.t157 756.008
R4 vp_p.n664 vp_p.t127 756.008
R5 vp_p.n664 vp_p.t1418 756.008
R6 vp_p.n662 vp_p.t534 756.008
R7 vp_p.n662 vp_p.t331 756.008
R8 vp_p.n660 vp_p.t939 756.008
R9 vp_p.n660 vp_p.t731 756.008
R10 vp_p.n658 vp_p.t877 756.008
R11 vp_p.n658 vp_p.t657 756.008
R12 vp_p.n656 vp_p.t1291 756.008
R13 vp_p.n656 vp_p.t1077 756.008
R14 vp_p.n654 vp_p.t1078 756.008
R15 vp_p.n654 vp_p.t865 756.008
R16 vp_p.n652 vp_p.t1497 756.008
R17 vp_p.n652 vp_p.t1281 756.008
R18 vp_p.n650 vp_p.t668 756.008
R19 vp_p.n650 vp_p.t465 756.008
R20 vp_p.n648 vp_p.t935 756.008
R21 vp_p.n648 vp_p.t720 756.008
R22 vp_p.n646 vp_p.t528 756.008
R23 vp_p.n646 vp_p.t320 756.008
R24 vp_p.n644 vp_p.t414 756.008
R25 vp_p.n644 vp_p.t211 756.008
R26 vp_p.n642 vp_p.t20 756.008
R27 vp_p.n642 vp_p.t1304 756.008
R28 vp_p.n640 vp_p.t243 756.008
R29 vp_p.n640 vp_p.t39 756.008
R30 vp_p.n638 vp_p.t1165 756.008
R31 vp_p.n638 vp_p.t958 756.008
R32 vp_p.n636 vp_p.t758 756.008
R33 vp_p.n636 vp_p.t550 756.008
R34 vp_p.n634 vp_p.t987 756.008
R35 vp_p.n634 vp_p.t775 756.008
R36 vp_p.n632 vp_p.t586 756.008
R37 vp_p.n632 vp_p.t380 756.008
R38 vp_p.n630 vp_p.t808 756.008
R39 vp_p.n630 vp_p.t607 756.008
R40 vp_p.n628 vp_p.t242 756.008
R41 vp_p.n628 vp_p.t38 756.008
R42 vp_p.n626 vp_p.t468 756.008
R43 vp_p.n626 vp_p.t271 756.008
R44 vp_p.n624 vp_p.t67 756.008
R45 vp_p.n624 vp_p.t1355 756.008
R46 vp_p.n622 vp_p.t1162 756.008
R47 vp_p.n622 vp_p.t951 756.008
R48 vp_p.n620 vp_p.t1388 756.008
R49 vp_p.n620 vp_p.t1183 756.008
R50 vp_p.n618 vp_p.t807 756.008
R51 vp_p.n618 vp_p.t606 756.008
R52 vp_p.n616 vp_p.t1037 756.008
R53 vp_p.n616 vp_p.t838 756.008
R54 vp_p.n614 vp_p.t635 756.008
R55 vp_p.n614 vp_p.t428 756.008
R56 vp_p.n612 vp_p.t240 756.008
R57 vp_p.n612 vp_p.t34 756.008
R58 vp_p.n610 vp_p.t466 756.008
R59 vp_p.n610 vp_p.t267 756.008
R60 vp_p.n608 vp_p.t1389 756.008
R61 vp_p.n608 vp_p.t1184 756.008
R62 vp_p.n606 vp_p.t128 756.008
R63 vp_p.n606 vp_p.t1422 756.008
R64 vp_p.n604 vp_p.t1221 756.008
R65 vp_p.n604 vp_p.t1002 756.008
R66 vp_p.n602 vp_p.t1237 756.008
R67 vp_p.n602 vp_p.t1020 756.008
R68 vp_p.n600 vp_p.t826 756.008
R69 vp_p.n600 vp_p.t621 756.008
R70 vp_p.n598 vp_p.t260 756.008
R71 vp_p.n598 vp_p.t53 756.008
R72 vp_p.n596 vp_p.t488 756.008
R73 vp_p.n596 vp_p.t288 756.008
R74 vp_p.n594 vp_p.t81 756.008
R75 vp_p.n594 vp_p.t1371 756.008
R76 vp_p.n592 vp_p.t321 756.008
R77 vp_p.n592 vp_p.t104 756.008
R78 vp_p.n590 vp_p.t1411 756.008
R79 vp_p.n590 vp_p.t1202 756.008
R80 vp_p.n588 vp_p.t1488 756.008
R81 vp_p.n588 vp_p.t1269 756.008
R82 vp_p.n586 vp_p.t1067 756.008
R83 vp_p.n586 vp_p.t857 756.008
R84 vp_p.n584 vp_p.t651 756.008
R85 vp_p.n584 vp_p.t442 756.008
R86 vp_p.n582 vp_p.t898 756.008
R87 vp_p.n582 vp_p.t678 756.008
R88 vp_p.n580 vp_p.t485 756.008
R89 vp_p.n580 vp_p.t283 756.008
R90 vp_p.n578 vp_p.t560 756.008
R91 vp_p.n578 vp_p.t350 756.008
R92 vp_p.n576 vp_p.t151 756.008
R93 vp_p.n576 vp_p.t1437 756.008
R94 vp_p.n574 vp_p.t1235 756.008
R95 vp_p.n574 vp_p.t1014 756.008
R96 vp_p.n572 vp_p.t1482 756.008
R97 vp_p.n572 vp_p.t1260 756.008
R98 vp_p.n570 vp_p.t1059 756.008
R99 vp_p.n570 vp_p.t850 756.008
R100 vp_p.n568 vp_p.t1132 756.008
R101 vp_p.n568 vp_p.t914 756.008
R102 vp_p.n566 vp_p.t716 756.008
R103 vp_p.n566 vp_p.t508 756.008
R104 vp_p.n564 vp_p.t961 756.008
R105 vp_p.n564 vp_p.t746 756.008
R106 vp_p.n562 vp_p.t554 756.008
R107 vp_p.n562 vp_p.t344 756.008
R108 vp_p.n560 vp_p.t144 756.008
R109 vp_p.n560 vp_p.t1432 756.008
R110 vp_p.n558 vp_p.t214 756.008
R111 vp_p.n558 vp_p.t9 756.008
R112 vp_p.n556 vp_p.t1311 756.008
R113 vp_p.n556 vp_p.t1093 756.008
R114 vp_p.n554 vp_p.t926 756.008
R115 vp_p.n554 vp_p.t710 756.008
R116 vp_p.n552 vp_p.t516 756.008
R117 vp_p.n552 vp_p.t308 756.008
R118 vp_p.n550 vp_p.t107 756.008
R119 vp_p.n550 vp_p.t1400 756.008
R120 vp_p.n548 vp_p.t186 756.008
R121 vp_p.n548 vp_p.t1472 756.008
R122 vp_p.n546 vp_p.t1272 756.008
R123 vp_p.n546 vp_p.t1051 756.008
R124 vp_p.n544 vp_p.t17 756.008
R125 vp_p.n544 vp_p.t1301 756.008
R126 vp_p.n542 vp_p.t1104 756.008
R127 vp_p.n542 vp_p.t885 756.008
R128 vp_p.n540 vp_p.t1333 756.008
R129 vp_p.n540 vp_p.t1121 756.008
R130 vp_p.n538 vp_p.t756 756.008
R131 vp_p.n538 vp_p.t546 756.008
R132 vp_p.n536 vp_p.t355 756.008
R133 vp_p.n536 vp_p.t137 756.008
R134 vp_p.n534 vp_p.t584 756.008
R135 vp_p.n534 vp_p.t377 756.008
R136 vp_p.n532 vp_p.t179 756.008
R137 vp_p.n532 vp_p.t1465 756.008
R138 vp_p.n530 vp_p.t407 756.008
R139 vp_p.n530 vp_p.t201 756.008
R140 vp_p.n528 vp_p.t1332 756.008
R141 vp_p.n528 vp_p.t1120 756.008
R142 vp_p.n526 vp_p.t65 756.008
R143 vp_p.n526 vp_p.t1353 756.008
R144 vp_p.n524 vp_p.t1159 756.008
R145 vp_p.n524 vp_p.t948 756.008
R146 vp_p.n522 vp_p.t750 756.008
R147 vp_p.n522 vp_p.t541 756.008
R148 vp_p.n521 vp_p.t982 756.008
R149 vp_p.n521 vp_p.t768 756.008
R150 vp_p.n519 vp_p.t1026 756.008
R151 vp_p.n519 vp_p.t467 756.008
R152 vp_p.n517 vp_p.t1452 756.008
R153 vp_p.n517 vp_p.t878 756.008
R154 vp_p.n515 vp_p.t365 756.008
R155 vp_p.n515 vp_p.t1292 756.008
R156 vp_p.n513 vp_p.t121 756.008
R157 vp_p.n513 vp_p.t1038 756.008
R158 vp_p.n511 vp_p.t531 756.008
R159 vp_p.n511 vp_p.t1461 756.008
R160 vp_p.n509 vp_p.t456 756.008
R161 vp_p.n509 vp_p.t1392 756.008
R162 vp_p.n507 vp_p.t871 756.008
R163 vp_p.n507 vp_p.t302 756.008
R164 vp_p.n505 vp_p.t1286 756.008
R165 vp_p.n505 vp_p.t700 756.008
R166 vp_p.n503 vp_p.t1069 756.008
R167 vp_p.n503 vp_p.t498 756.008
R168 vp_p.n501 vp_p.t1491 756.008
R169 vp_p.n501 vp_p.t906 756.008
R170 vp_p.n499 vp_p.t927 756.008
R171 vp_p.n499 vp_p.t371 756.008
R172 vp_p.n497 vp_p.t520 756.008
R173 vp_p.n497 vp_p.t1458 756.008
R174 vp_p.n495 vp_p.t410 756.008
R175 vp_p.n495 vp_p.t1342 756.008
R176 vp_p.n493 vp_p.t13 756.008
R177 vp_p.n493 vp_p.t933 756.008
R178 vp_p.n491 vp_p.t1096 756.008
R179 vp_p.n491 vp_p.t524 756.008
R180 vp_p.n489 vp_p.t1161 756.008
R181 vp_p.n489 vp_p.t593 756.008
R182 vp_p.n487 vp_p.t752 756.008
R183 vp_p.n487 vp_p.t192 756.008
R184 vp_p.n485 vp_p.t983 756.008
R185 vp_p.n485 vp_p.t416 756.008
R186 vp_p.n483 vp_p.t581 756.008
R187 vp_p.n483 vp_p.t24 756.008
R188 vp_p.n481 vp_p.t174 756.008
R189 vp_p.n481 vp_p.t1110 756.008
R190 vp_p.n479 vp_p.t238 756.008
R191 vp_p.n479 vp_p.t1168 756.008
R192 vp_p.n477 vp_p.t1329 756.008
R193 vp_p.n477 vp_p.t761 756.008
R194 vp_p.n475 vp_p.t63 756.008
R195 vp_p.n475 vp_p.t989 756.008
R196 vp_p.n473 vp_p.t1154 756.008
R197 vp_p.n473 vp_p.t590 756.008
R198 vp_p.n471 vp_p.t1385 756.008
R199 vp_p.n471 vp_p.t809 756.008
R200 vp_p.n469 vp_p.t803 756.008
R201 vp_p.n469 vp_p.t247 756.008
R202 vp_p.n467 vp_p.t404 756.008
R203 vp_p.n467 vp_p.t1339 756.008
R204 vp_p.n465 vp_p.t631 756.008
R205 vp_p.n465 vp_p.t69 756.008
R206 vp_p.n463 vp_p.t233 756.008
R207 vp_p.n463 vp_p.t1164 756.008
R208 vp_p.n461 vp_p.t462 756.008
R209 vp_p.n461 vp_p.t1394 756.008
R210 vp_p.n459 vp_p.t1386 756.008
R211 vp_p.n459 vp_p.t810 756.008
R212 vp_p.n457 vp_p.t123 756.008
R213 vp_p.n457 vp_p.t1040 756.008
R214 vp_p.n455 vp_p.t1217 756.008
R215 vp_p.n455 vp_p.t637 756.008
R216 vp_p.n453 vp_p.t798 756.008
R217 vp_p.n453 vp_p.t245 756.008
R218 vp_p.n451 vp_p.t822 756.008
R219 vp_p.n451 vp_p.t266 756.008
R220 vp_p.n449 vp_p.t254 756.008
R221 vp_p.n449 vp_p.t1182 756.008
R222 vp_p.n447 vp_p.t484 756.008
R223 vp_p.n447 vp_p.t1421 756.008
R224 vp_p.n445 vp_p.t77 756.008
R225 vp_p.n445 vp_p.t1001 756.008
R226 vp_p.n443 vp_p.t1173 756.008
R227 vp_p.n443 vp_p.t601 756.008
R228 vp_p.n441 vp_p.t1405 756.008
R229 vp_p.n441 vp_p.t831 756.008
R230 vp_p.n439 vp_p.t821 756.008
R231 vp_p.n439 vp_p.t265 756.008
R232 vp_p.n437 vp_p.t1058 756.008
R233 vp_p.n437 vp_p.t494 756.008
R234 vp_p.n435 vp_p.t645 756.008
R235 vp_p.n435 vp_p.t84 756.008
R236 vp_p.n433 vp_p.t890 756.008
R237 vp_p.n433 vp_p.t329 756.008
R238 vp_p.n431 vp_p.t477 756.008
R239 vp_p.n431 vp_p.t1417 756.008
R240 vp_p.n429 vp_p.t1406 756.008
R241 vp_p.n429 vp_p.t833 756.008
R242 vp_p.n427 vp_p.t142 756.008
R243 vp_p.n427 vp_p.t1073 756.008
R244 vp_p.n425 vp_p.t1228 756.008
R245 vp_p.n425 vp_p.t655 756.008
R246 vp_p.n423 vp_p.t1470 756.008
R247 vp_p.n423 vp_p.t901 756.008
R248 vp_p.n421 vp_p.t1048 756.008
R249 vp_p.n421 vp_p.t489 756.008
R250 vp_p.n419 vp_p.t1125 756.008
R251 vp_p.n419 vp_p.t565 756.008
R252 vp_p.n417 vp_p.t707 756.008
R253 vp_p.n417 vp_p.t154 756.008
R254 vp_p.n415 vp_p.t309 756.008
R255 vp_p.n415 vp_p.t1240 756.008
R256 vp_p.n413 vp_p.t545 756.008
R257 vp_p.n413 vp_p.t1487 756.008
R258 vp_p.n411 vp_p.t136 756.008
R259 vp_p.n411 vp_p.t1066 756.008
R260 vp_p.n409 vp_p.t208 756.008
R261 vp_p.n409 vp_p.t1136 756.008
R262 vp_p.n407 vp_p.t1302 756.008
R263 vp_p.n407 vp_p.t722 756.008
R264 vp_p.n405 vp_p.t884 756.008
R265 vp_p.n405 vp_p.t322 756.008
R266 vp_p.n403 vp_p.t507 756.008
R267 vp_p.n403 vp_p.t1451 756.008
R268 vp_p.n401 vp_p.t98 756.008
R269 vp_p.n401 vp_p.t1025 756.008
R270 vp_p.n399 vp_p.t177 756.008
R271 vp_p.n399 vp_p.t1112 756.008
R272 vp_p.n397 vp_p.t1262 756.008
R273 vp_p.n397 vp_p.t692 756.008
R274 vp_p.n395 vp_p.t8 756.008
R275 vp_p.n395 vp_p.t928 756.008
R276 vp_p.n393 vp_p.t1094 756.008
R277 vp_p.n393 vp_p.t523 756.008
R278 vp_p.n391 vp_p.t673 756.008
R279 vp_p.n391 vp_p.t112 756.008
R280 vp_p.n389 vp_p.t749 756.008
R281 vp_p.n389 vp_p.t190 756.008
R282 vp_p.n387 vp_p.t345 756.008
R283 vp_p.n387 vp_p.t1279 756.008
R284 vp_p.n385 vp_p.t577 756.008
R285 vp_p.n385 vp_p.t21 756.008
R286 vp_p.n383 vp_p.t171 756.008
R287 vp_p.n383 vp_p.t1109 756.008
R288 vp_p.n381 vp_p.t1255 756.008
R289 vp_p.n381 vp_p.t688 756.008
R290 vp_p.n379 vp_p.t1326 756.008
R291 vp_p.n379 vp_p.t759 756.008
R292 vp_p.n377 vp_p.t910 756.008
R293 vp_p.n377 vp_p.t360 756.008
R294 vp_p.n375 vp_p.t1151 756.008
R295 vp_p.n375 vp_p.t588 756.008
R296 vp_p.n373 vp_p.t741 756.008
R297 vp_p.n373 vp_p.t185 756.008
R298 vp_p.n372 vp_p.t978 756.008
R299 vp_p.n372 vp_p.t413 756.008
R300 vp_p.n370 vp_p.t667 756.008
R301 vp_p.n370 vp_p.t908 756.008
R302 vp_p.n368 vp_p.t1084 756.008
R303 vp_p.n368 vp_p.t1322 756.008
R304 vp_p.n366 vp_p.t842 756.008
R305 vp_p.n366 vp_p.t1087 756.008
R306 vp_p.n364 vp_p.t1252 756.008
R307 vp_p.n364 vp_p.t2 756.008
R308 vp_p.n362 vp_p.t166 756.008
R309 vp_p.n362 vp_p.t400 756.008
R310 vp_p.n360 vp_p.t92 756.008
R311 vp_p.n360 vp_p.t339 756.008
R312 vp_p.n358 vp_p.t499 756.008
R313 vp_p.n358 vp_p.t739 756.008
R314 vp_p.n356 vp_p.t300 756.008
R315 vp_p.n356 vp_p.t536 756.008
R316 vp_p.n354 vp_p.t699 756.008
R317 vp_p.n354 vp_p.t943 756.008
R318 vp_p.n352 vp_p.t1396 756.008
R319 vp_p.n352 vp_p.t138 756.008
R320 vp_p.n350 vp_p.t163 756.008
R321 vp_p.n350 vp_p.t396 756.008
R322 vp_p.n348 vp_p.t1248 756.008
R323 vp_p.n348 vp_p.t1499 756.008
R324 vp_p.n346 vp_p.t1139 756.008
R325 vp_p.n346 vp_p.t1369 756.008
R326 vp_p.n344 vp_p.t724 756.008
R327 vp_p.n344 vp_p.t971 756.008
R328 vp_p.n342 vp_p.t968 756.008
R329 vp_p.n342 vp_p.t1199 756.008
R330 vp_p.n340 vp_p.t393 756.008
R331 vp_p.n340 vp_p.t619 756.008
R332 vp_p.n338 vp_p.t1492 756.008
R333 vp_p.n338 vp_p.t224 756.008
R334 vp_p.n336 vp_p.t221 756.008
R335 vp_p.n336 vp_p.t439 756.008
R336 vp_p.n334 vp_p.t1316 756.008
R337 vp_p.n334 vp_p.t51 756.008
R338 vp_p.n332 vp_p.t48 756.008
R339 vp_p.n332 vp_p.t279 756.008
R340 vp_p.n330 vp_p.t967 756.008
R341 vp_p.n330 vp_p.t1198 756.008
R342 vp_p.n328 vp_p.t1196 756.008
R343 vp_p.n328 vp_p.t1434 756.008
R344 vp_p.n326 vp_p.t784 756.008
R345 vp_p.n326 vp_p.t1011 756.008
R346 vp_p.n324 vp_p.t391 756.008
R347 vp_p.n324 vp_p.t618 756.008
R348 vp_p.n322 vp_p.t613 756.008
R349 vp_p.n322 vp_p.t848 756.008
R350 vp_p.n320 vp_p.t47 756.008
R351 vp_p.n320 vp_p.t280 756.008
R352 vp_p.n318 vp_p.t277 756.008
R353 vp_p.n318 vp_p.t503 756.008
R354 vp_p.n316 vp_p.t1363 756.008
R355 vp_p.n316 vp_p.t96 756.008
R356 vp_p.n314 vp_p.t964 756.008
R357 vp_p.n314 vp_p.t1197 756.008
R358 vp_p.n312 vp_p.t1194 756.008
R359 vp_p.n312 vp_p.t1430 756.008
R360 vp_p.n310 vp_p.t615 756.008
R361 vp_p.n310 vp_p.t847 756.008
R362 vp_p.n308 vp_p.t844 756.008
R363 vp_p.n308 vp_p.t1090 756.008
R364 vp_p.n306 vp_p.t434 756.008
R365 vp_p.n306 vp_p.t672 756.008
R366 vp_p.n304 vp_p.t461 756.008
R367 vp_p.n304 vp_p.t698 756.008
R368 vp_p.n302 vp_p.t60 756.008
R369 vp_p.n302 vp_p.t299 756.008
R370 vp_p.n300 vp_p.t980 756.008
R371 vp_p.n300 vp_p.t1220 756.008
R372 vp_p.n298 vp_p.t1216 756.008
R373 vp_p.n298 vp_p.t1459 756.008
R374 vp_p.n296 vp_p.t797 756.008
R375 vp_p.n296 vp_p.t1034 756.008
R376 vp_p.n294 vp_p.t1029 756.008
R377 vp_p.n294 vp_p.t1290 756.008
R378 vp_p.n292 vp_p.t628 756.008
R379 vp_p.n292 vp_p.t875 756.008
R380 vp_p.n290 vp_p.t695 756.008
R381 vp_p.n290 vp_p.t938 756.008
R382 vp_p.n288 vp_p.t297 756.008
R383 vp_p.n288 vp_p.t532 756.008
R384 vp_p.n286 vp_p.t1380 756.008
R385 vp_p.n286 vp_p.t125 756.008
R386 vp_p.n284 vp_p.t119 756.008
R387 vp_p.n284 vp_p.t369 756.008
R388 vp_p.n282 vp_p.t1212 756.008
R389 vp_p.n282 vp_p.t1454 756.008
R390 vp_p.n280 vp_p.t1283 756.008
R391 vp_p.n280 vp_p.t27 756.008
R392 vp_p.n278 vp_p.t869 756.008
R393 vp_p.n278 vp_p.t1114 756.008
R394 vp_p.n276 vp_p.t454 756.008
R395 vp_p.n276 vp_p.t696 756.008
R396 vp_p.n274 vp_p.t691 756.008
R397 vp_p.n274 vp_p.t936 756.008
R398 vp_p.n272 vp_p.t292 756.008
R399 vp_p.n272 vp_p.t529 756.008
R400 vp_p.n270 vp_p.t363 756.008
R401 vp_p.n270 vp_p.t594 756.008
R402 vp_p.n268 vp_p.t1449 756.008
R403 vp_p.n268 vp_p.t194 756.008
R404 vp_p.n266 vp_p.t189 756.008
R405 vp_p.n266 vp_p.t417 756.008
R406 vp_p.n264 vp_p.t1277 756.008
R407 vp_p.n264 vp_p.t25 756.008
R408 vp_p.n262 vp_p.t864 756.008
R409 vp_p.n262 vp_p.t1111 756.008
R410 vp_p.n260 vp_p.t929 756.008
R411 vp_p.n260 vp_p.t1169 756.008
R412 vp_p.n258 vp_p.t522 756.008
R413 vp_p.n258 vp_p.t762 756.008
R414 vp_p.n256 vp_p.t156 756.008
R415 vp_p.n256 vp_p.t394 756.008
R416 vp_p.n254 vp_p.t1239 756.008
R417 vp_p.n254 vp_p.t1495 756.008
R418 vp_p.n252 vp_p.t827 756.008
R419 vp_p.n252 vp_p.t1076 756.008
R420 vp_p.n250 vp_p.t902 756.008
R421 vp_p.n250 vp_p.t1142 756.008
R422 vp_p.n248 vp_p.t490 756.008
R423 vp_p.n248 vp_p.t730 756.008
R424 vp_p.n246 vp_p.t721 756.008
R425 vp_p.n246 vp_p.t970 756.008
R426 vp_p.n244 vp_p.t323 756.008
R427 vp_p.n244 vp_p.t568 756.008
R428 vp_p.n242 vp_p.t562 756.008
R429 vp_p.n242 vp_p.t786 756.008
R430 vp_p.n240 vp_p.t1489 756.008
R431 vp_p.n240 vp_p.t223 756.008
R432 vp_p.n238 vp_p.t1068 756.008
R433 vp_p.n238 vp_p.t1319 756.008
R434 vp_p.n236 vp_p.t1315 756.008
R435 vp_p.n236 vp_p.t49 756.008
R436 vp_p.n234 vp_p.t899 756.008
R437 vp_p.n234 vp_p.t1137 756.008
R438 vp_p.n232 vp_p.t1133 756.008
R439 vp_p.n232 vp_p.t1365 756.008
R440 vp_p.n230 vp_p.t561 756.008
R441 vp_p.n230 vp_p.t787 756.008
R442 vp_p.n228 vp_p.t782 756.008
R443 vp_p.n228 vp_p.t1009 756.008
R444 vp_p.n226 vp_p.t390 756.008
R445 vp_p.n226 vp_p.t616 756.008
R446 vp_p.n224 vp_p.t1483 756.008
R447 vp_p.n224 vp_p.t220 756.008
R448 vp_p.n223 vp_p.t215 756.008
R449 vp_p.n223 vp_p.t437 756.008
R450 vp_p.n221 vp_p.t701 756.008
R451 vp_p.n221 vp_p.t834 756.008
R452 vp_p.n219 vp_p.t1117 756.008
R453 vp_p.n219 vp_p.t1245 756.008
R454 vp_p.n217 vp_p.t31 756.008
R455 vp_p.n217 vp_p.t160 756.008
R456 vp_p.n215 vp_p.t1295 756.008
R457 vp_p.n215 vp_p.t1424 756.008
R458 vp_p.n213 vp_p.t200 756.008
R459 vp_p.n213 vp_p.t334 756.008
R460 vp_p.n211 vp_p.t131 756.008
R461 vp_p.n211 vp_p.t269 756.008
R462 vp_p.n209 vp_p.t539 756.008
R463 vp_p.n209 vp_p.t664 756.008
R464 vp_p.n207 vp_p.t945 756.008
R465 vp_p.n207 vp_p.t1082 756.008
R466 vp_p.n205 vp_p.t735 756.008
R467 vp_p.n205 vp_p.t873 756.008
R468 vp_p.n203 vp_p.t1146 756.008
R469 vp_p.n203 vp_p.t1287 756.008
R470 vp_p.n201 vp_p.t597 756.008
R471 vp_p.n201 vp_p.t726 756.008
R472 vp_p.n199 vp_p.t196 756.008
R473 vp_p.n199 vp_p.t327 756.008
R474 vp_p.n197 vp_p.t74 756.008
R475 vp_p.n197 vp_p.t216 756.008
R476 vp_p.n195 vp_p.t1171 756.008
R477 vp_p.n195 vp_p.t1312 756.008
R478 vp_p.n193 vp_p.t764 756.008
R479 vp_p.n193 vp_p.t897 756.008
R480 vp_p.n191 vp_p.t817 756.008
R481 vp_p.n191 vp_p.t963 756.008
R482 vp_p.n189 vp_p.t419 756.008
R483 vp_p.n189 vp_p.t559 756.008
R484 vp_p.n187 vp_p.t642 756.008
R485 vp_p.n187 vp_p.t779 756.008
R486 vp_p.n185 vp_p.t250 756.008
R487 vp_p.n185 vp_p.t386 756.008
R488 vp_p.n183 vp_p.t1341 756.008
R489 vp_p.n183 vp_p.t1477 756.008
R490 vp_p.n181 vp_p.t1402 756.008
R491 vp_p.n181 vp_p.t44 756.008
R492 vp_p.n179 vp_p.t991 756.008
R493 vp_p.n179 vp_p.t1130 756.008
R494 vp_p.n177 vp_p.t1224 756.008
R495 vp_p.n177 vp_p.t1360 756.008
R496 vp_p.n175 vp_p.t814 756.008
R497 vp_p.n175 vp_p.t957 756.008
R498 vp_p.n173 vp_p.t1046 756.008
R499 vp_p.n173 vp_p.t1189 756.008
R500 vp_p.n171 vp_p.t474 756.008
R501 vp_p.n171 vp_p.t611 756.008
R502 vp_p.n169 vp_p.t71 756.008
R503 vp_p.n169 vp_p.t210 756.008
R504 vp_p.n167 vp_p.t305 756.008
R505 vp_p.n167 vp_p.t431 756.008
R506 vp_p.n165 vp_p.t1399 756.008
R507 vp_p.n165 vp_p.t40 756.008
R508 vp_p.n163 vp_p.t134 756.008
R509 vp_p.n163 vp_p.t270 756.008
R510 vp_p.n161 vp_p.t1045 756.008
R511 vp_p.n161 vp_p.t1188 756.008
R512 vp_p.n159 vp_p.t1298 756.008
R513 vp_p.n159 vp_p.t1425 756.008
R514 vp_p.n157 vp_p.t883 756.008
R515 vp_p.n157 vp_p.t1005 756.008
R516 vp_p.n155 vp_p.t471 756.008
R517 vp_p.n155 vp_p.t605 756.008
R518 vp_p.n153 vp_p.t496 756.008
R519 vp_p.n153 vp_p.t624 756.008
R520 vp_p.n151 vp_p.t1426 756.008
R521 vp_p.n151 vp_p.t55 756.008
R522 vp_p.n149 vp_p.t164 756.008
R523 vp_p.n149 vp_p.t291 756.008
R524 vp_p.n147 vp_p.t1249 756.008
R525 vp_p.n147 vp_p.t1374 756.008
R526 vp_p.n145 vp_p.t837 756.008
R527 vp_p.n145 vp_p.t973 756.008
R528 vp_p.n143 vp_p.t1081 756.008
R529 vp_p.n143 vp_p.t1206 756.008
R530 vp_p.n141 vp_p.t497 756.008
R531 vp_p.n141 vp_p.t623 756.008
R532 vp_p.n139 vp_p.t732 756.008
R533 vp_p.n139 vp_p.t861 756.008
R534 vp_p.n137 vp_p.t333 756.008
R535 vp_p.n137 vp_p.t447 756.008
R536 vp_p.n135 vp_p.t569 756.008
R537 vp_p.n135 vp_p.t685 756.008
R538 vp_p.n133 vp_p.t159 756.008
R539 vp_p.n133 vp_p.t287 756.008
R540 vp_p.n131 vp_p.t1080 756.008
R541 vp_p.n131 vp_p.t1205 756.008
R542 vp_p.n129 vp_p.t1320 756.008
R543 vp_p.n129 vp_p.t1444 756.008
R544 vp_p.n127 vp_p.t905 756.008
R545 vp_p.n127 vp_p.t1021 756.008
R546 vp_p.n125 vp_p.t1141 756.008
R547 vp_p.n125 vp_p.t1268 756.008
R548 vp_p.n123 vp_p.t728 756.008
R549 vp_p.n123 vp_p.t856 756.008
R550 vp_p.n121 vp_p.t789 756.008
R551 vp_p.n121 vp_p.t923 756.008
R552 vp_p.n119 vp_p.t395 756.008
R553 vp_p.n119 vp_p.t513 756.008
R554 vp_p.n117 vp_p.t1494 756.008
R555 vp_p.n117 vp_p.t105 756.008
R556 vp_p.n115 vp_p.t222 756.008
R557 vp_p.n115 vp_p.t351 756.008
R558 vp_p.n113 vp_p.t1317 756.008
R559 vp_p.n113 vp_p.t1438 756.008
R560 vp_p.n111 vp_p.t1367 756.008
R561 vp_p.n111 vp_p.t15 756.008
R562 vp_p.n109 vp_p.t969 756.008
R563 vp_p.n109 vp_p.t1100 756.008
R564 vp_p.n107 vp_p.t566 756.008
R565 vp_p.n107 vp_p.t680 756.008
R566 vp_p.n105 vp_p.t193 756.008
R567 vp_p.n105 vp_p.t316 756.008
R568 vp_p.n103 vp_p.t1285 756.008
R569 vp_p.n103 vp_p.t1407 756.008
R570 vp_p.n101 vp_p.t1343 756.008
R571 vp_p.n101 vp_p.t1481 756.008
R572 vp_p.n99 vp_p.t937 756.008
R573 vp_p.n99 vp_p.t1060 756.008
R574 vp_p.n97 vp_p.t1170 756.008
R575 vp_p.n97 vp_p.t1309 756.008
R576 vp_p.n95 vp_p.t763 756.008
R577 vp_p.n95 vp_p.t893 756.008
R578 vp_p.n93 vp_p.t368 756.008
R579 vp_p.n93 vp_p.t478 756.008
R580 vp_p.n91 vp_p.t418 756.008
R581 vp_p.n91 vp_p.t555 756.008
R582 vp_p.n89 vp_p.t26 756.008
R583 vp_p.n89 vp_p.t146 756.008
R584 vp_p.n87 vp_p.t248 756.008
R585 vp_p.n87 vp_p.t383 756.008
R586 vp_p.n85 vp_p.t1340 756.008
R587 vp_p.n85 vp_p.t1471 756.008
R588 vp_p.n83 vp_p.t931 756.008
R589 vp_p.n83 vp_p.t1050 756.008
R590 vp_p.n81 vp_p.t990 756.008
R591 vp_p.n81 vp_p.t1127 756.008
R592 vp_p.n79 vp_p.t592 756.008
R593 vp_p.n79 vp_p.t709 756.008
R594 vp_p.n77 vp_p.t811 756.008
R595 vp_p.n77 vp_p.t954 756.008
R596 vp_p.n75 vp_p.t415 756.008
R597 vp_p.n75 vp_p.t548 756.008
R598 vp_p.n74 vp_p.t638 756.008
R599 vp_p.n74 vp_p.t774 756.008
R600 vp_p.n970 vp_p.t629 756.008
R601 vp_p.n970 vp_p.t68 756.008
R602 vp_p.n968 vp_p.t1030 756.008
R603 vp_p.n968 vp_p.t469 756.008
R604 vp_p.n966 vp_p.t796 756.008
R605 vp_p.n966 vp_p.t244 756.008
R606 vp_p.n964 vp_p.t1215 756.008
R607 vp_p.n964 vp_p.t636 756.008
R608 vp_p.n962 vp_p.t124 756.008
R609 vp_p.n962 vp_p.t1042 756.008
R610 vp_p.n960 vp_p.t59 756.008
R611 vp_p.n960 vp_p.t988 756.008
R612 vp_p.n958 vp_p.t460 756.008
R613 vp_p.n958 vp_p.t1393 756.008
R614 vp_p.n956 vp_p.t261 756.008
R615 vp_p.n956 vp_p.t1190 756.008
R616 vp_p.n954 vp_p.t656 756.008
R617 vp_p.n954 vp_p.t91 756.008
R618 vp_p.n952 vp_p.t1358 756.008
R619 vp_p.n952 vp_p.t785 756.008
R620 vp_p.n950 vp_p.t114 756.008
R621 vp_p.n950 vp_p.t1036 756.008
R622 vp_p.n948 vp_p.t1209 756.008
R623 vp_p.n948 vp_p.t633 756.008
R624 vp_p.n946 vp_p.t1102 756.008
R625 vp_p.n946 vp_p.t530 756.008
R626 vp_p.n944 vp_p.t681 756.008
R627 vp_p.n944 vp_p.t120 756.008
R628 vp_p.n942 vp_p.t918 756.008
R629 vp_p.n942 vp_p.t367 756.008
R630 vp_p.n940 vp_p.t353 756.008
R631 vp_p.n940 vp_p.t1284 756.008
R632 vp_p.n938 vp_p.t1439 756.008
R633 vp_p.n938 vp_p.t872 756.008
R634 vp_p.n936 vp_p.t178 756.008
R635 vp_p.n936 vp_p.t1113 756.008
R636 vp_p.n934 vp_p.t1264 756.008
R637 vp_p.n934 vp_p.t693 756.008
R638 vp_p.n932 vp_p.t10 756.008
R639 vp_p.n932 vp_p.t930 756.008
R640 vp_p.n930 vp_p.t917 756.008
R641 vp_p.n930 vp_p.t366 756.008
R642 vp_p.n928 vp_p.t1158 756.008
R643 vp_p.n928 vp_p.t591 756.008
R644 vp_p.n926 vp_p.t747 756.008
R645 vp_p.n926 vp_p.t191 756.008
R646 vp_p.n924 vp_p.t346 756.008
R647 vp_p.n924 vp_p.t1280 756.008
R648 vp_p.n922 vp_p.t580 756.008
R649 vp_p.n922 vp_p.t23 756.008
R650 vp_p.n920 vp_p.t12 756.008
R651 vp_p.n920 vp_p.t932 756.008
R652 vp_p.n918 vp_p.t237 756.008
R653 vp_p.n918 vp_p.t1166 756.008
R654 vp_p.n916 vp_p.t1327 756.008
R655 vp_p.n916 vp_p.t760 756.008
R656 vp_p.n914 vp_p.t912 756.008
R657 vp_p.n914 vp_p.t361 756.008
R658 vp_p.n912 vp_p.t1153 756.008
R659 vp_p.n912 vp_p.t589 756.008
R660 vp_p.n910 vp_p.t579 756.008
R661 vp_p.n910 vp_p.t22 756.008
R662 vp_p.n908 vp_p.t802 756.008
R663 vp_p.n908 vp_p.t246 756.008
R664 vp_p.n906 vp_p.t403 756.008
R665 vp_p.n906 vp_p.t1338 756.008
R666 vp_p.n904 vp_p.t421 756.008
R667 vp_p.n904 vp_p.t1352 756.008
R668 vp_p.n902 vp_p.t28 756.008
R669 vp_p.n902 vp_p.t947 756.008
R670 vp_p.n900 vp_p.t940 756.008
R671 vp_p.n900 vp_p.t378 756.008
R672 vp_p.n898 vp_p.t1174 756.008
R673 vp_p.n898 vp_p.t603 756.008
R674 vp_p.n896 vp_p.t765 756.008
R675 vp_p.n896 vp_p.t202 756.008
R676 vp_p.n894 vp_p.t993 756.008
R677 vp_p.n894 vp_p.t427 756.008
R678 vp_p.n892 vp_p.t595 756.008
R679 vp_p.n892 vp_p.t33 756.008
R680 vp_p.n890 vp_p.t648 756.008
R681 vp_p.n890 vp_p.t88 756.008
R682 vp_p.n888 vp_p.t253 756.008
R683 vp_p.n888 vp_p.t1181 756.008
R684 vp_p.n886 vp_p.t1344 756.008
R685 vp_p.n886 vp_p.t769 756.008
R686 vp_p.n884 vp_p.t75 756.008
R687 vp_p.n884 vp_p.t999 756.008
R688 vp_p.n882 vp_p.t1172 756.008
R689 vp_p.n882 vp_p.t600 756.008
R690 vp_p.n880 vp_p.t1233 756.008
R691 vp_p.n880 vp_p.t661 756.008
R692 vp_p.n878 vp_p.t819 756.008
R693 vp_p.n878 vp_p.t263 756.008
R694 vp_p.n876 vp_p.t420 756.008
R695 vp_p.n876 vp_p.t1348 756.008
R696 vp_p.n874 vp_p.t643 756.008
R697 vp_p.n874 vp_p.t82 756.008
R698 vp_p.n872 vp_p.t251 756.008
R699 vp_p.n872 vp_p.t1179 756.008
R700 vp_p.n870 vp_p.t314 756.008
R701 vp_p.n870 vp_p.t1243 756.008
R702 vp_p.n868 vp_p.t1403 756.008
R703 vp_p.n868 vp_p.t830 756.008
R704 vp_p.n866 vp_p.t140 756.008
R705 vp_p.n866 vp_p.t1071 756.008
R706 vp_p.n864 vp_p.t1225 756.008
R707 vp_p.n864 vp_p.t653 756.008
R708 vp_p.n862 vp_p.t815 756.008
R709 vp_p.n862 vp_p.t259 756.008
R710 vp_p.n860 vp_p.t888 756.008
R711 vp_p.n860 vp_p.t326 756.008
R712 vp_p.n858 vp_p.t475 756.008
R713 vp_p.n858 vp_p.t1415 756.008
R714 vp_p.n856 vp_p.t102 756.008
R715 vp_p.n856 vp_p.t1027 756.008
R716 vp_p.n854 vp_p.t1201 756.008
R717 vp_p.n854 vp_p.t627 756.008
R718 vp_p.n852 vp_p.t788 756.008
R719 vp_p.n852 vp_p.t228 756.008
R720 vp_p.n850 vp_p.t855 756.008
R721 vp_p.n850 vp_p.t296 756.008
R722 vp_p.n848 vp_p.t441 756.008
R723 vp_p.n848 vp_p.t1379 756.008
R724 vp_p.n846 vp_p.t677 756.008
R725 vp_p.n846 vp_p.t118 756.008
R726 vp_p.n844 vp_p.t282 756.008
R727 vp_p.n844 vp_p.t1211 756.008
R728 vp_p.n842 vp_p.t505 756.008
R729 vp_p.n842 vp_p.t1447 756.008
R730 vp_p.n840 vp_p.t1436 756.008
R731 vp_p.n840 vp_p.t868 756.008
R732 vp_p.n838 vp_p.t1013 756.008
R733 vp_p.n838 vp_p.t452 756.008
R734 vp_p.n836 vp_p.t1259 756.008
R735 vp_p.n836 vp_p.t690 756.008
R736 vp_p.n834 vp_p.t849 756.008
R737 vp_p.n834 vp_p.t290 756.008
R738 vp_p.n832 vp_p.t1092 756.008
R739 vp_p.n832 vp_p.t521 756.008
R740 vp_p.n830 vp_p.t506 756.008
R741 vp_p.n830 vp_p.t1448 756.008
R742 vp_p.n828 vp_p.t744 756.008
R743 vp_p.n828 vp_p.t188 756.008
R744 vp_p.n826 vp_p.t343 756.008
R745 vp_p.n826 vp_p.t1276 756.008
R746 vp_p.n824 vp_p.t1431 756.008
R747 vp_p.n824 vp_p.t863 756.008
R748 vp_p.n823 vp_p.t170 756.008
R749 vp_p.n823 vp_p.t1108 756.008
R750 vp_p.n1119 vp_p.t1362 756.008
R751 vp_p.n1119 vp_p.t1236 756.008
R752 vp_p.n1117 vp_p.t275 756.008
R753 vp_p.n1117 vp_p.t152 756.008
R754 vp_p.n1115 vp_p.t670 756.008
R755 vp_p.n1115 vp_p.t564 756.008
R756 vp_p.n1113 vp_p.t433 756.008
R757 vp_p.n1113 vp_p.t325 756.008
R758 vp_p.n1111 vp_p.t845 756.008
R759 vp_p.n1111 vp_p.t725 756.008
R760 vp_p.n1109 vp_p.t781 756.008
R761 vp_p.n1109 vp_p.t652 756.008
R762 vp_p.n1107 vp_p.t1193 756.008
R763 vp_p.n1107 vp_p.t1070 756.008
R764 vp_p.n1105 vp_p.t93 756.008
R765 vp_p.n1105 vp_p.t1493 756.008
R766 vp_p.n1103 vp_p.t1391 756.008
R767 vp_p.n1103 vp_p.t1275 756.008
R768 vp_p.n1101 vp_p.t301 756.008
R769 vp_p.n1101 vp_p.t187 756.008
R770 vp_p.n1099 vp_p.t1250 756.008
R771 vp_p.n1099 vp_p.t1134 756.008
R772 vp_p.n1097 vp_p.t840 756.008
R773 vp_p.n1097 vp_p.t717 756.008
R774 vp_p.n1095 vp_p.t729 756.008
R775 vp_p.n1095 vp_p.t608 756.008
R776 vp_p.n1093 vp_p.t330 756.008
R777 vp_p.n1093 vp_p.t207 756.008
R778 vp_p.n1091 vp_p.t1419 756.008
R779 vp_p.n1091 vp_p.t1300 756.008
R780 vp_p.n1089 vp_p.t1496 756.008
R781 vp_p.n1089 vp_p.t1356 756.008
R782 vp_p.n1087 vp_p.t1074 756.008
R783 vp_p.n1087 vp_p.t952 756.008
R784 vp_p.n1085 vp_p.t1318 756.008
R785 vp_p.n1085 vp_p.t1186 756.008
R786 vp_p.n1083 vp_p.t903 756.008
R787 vp_p.n1083 vp_p.t771 756.008
R788 vp_p.n1081 vp_p.t491 756.008
R789 vp_p.n1081 vp_p.t375 756.008
R790 vp_p.n1079 vp_p.t567 756.008
R791 vp_p.n1079 vp_p.t429 756.008
R792 vp_p.n1077 vp_p.t158 756.008
R793 vp_p.n1077 vp_p.t36 756.008
R794 vp_p.n1075 vp_p.t392 756.008
R795 vp_p.n1075 vp_p.t268 756.008
R796 vp_p.n1073 vp_p.t1490 756.008
R797 vp_p.n1073 vp_p.t1351 756.008
R798 vp_p.n1071 vp_p.t219 756.008
R799 vp_p.n1071 vp_p.t86 756.008
R800 vp_p.n1069 vp_p.t1138 756.008
R801 vp_p.n1069 vp_p.t1003 756.008
R802 vp_p.n1067 vp_p.t723 756.008
R803 vp_p.n1067 vp_p.t602 756.008
R804 vp_p.n1065 vp_p.t966 756.008
R805 vp_p.n1065 vp_p.t835 756.008
R806 vp_p.n1063 vp_p.t563 756.008
R807 vp_p.n1063 vp_p.t426 756.008
R808 vp_p.n1061 vp_p.t783 756.008
R809 vp_p.n1061 vp_p.t659 756.008
R810 vp_p.n1059 vp_p.t218 756.008
R811 vp_p.n1059 vp_p.t85 756.008
R812 vp_p.n1057 vp_p.t436 756.008
R813 vp_p.n1057 vp_p.t332 756.008
R814 vp_p.n1055 vp_p.t46 756.008
R815 vp_p.n1055 vp_p.t1420 756.008
R816 vp_p.n1053 vp_p.t1135 756.008
R817 vp_p.n1053 vp_p.t998 756.008
R818 vp_p.n1051 vp_p.t1150 756.008
R819 vp_p.n1051 vp_p.t1015 756.008
R820 vp_p.n1049 vp_p.t578 756.008
R821 vp_p.n1049 vp_p.t443 756.008
R822 vp_p.n1047 vp_p.t801 756.008
R823 vp_p.n1047 vp_p.t682 756.008
R824 vp_p.n1045 vp_p.t402 756.008
R825 vp_p.n1045 vp_p.t284 756.008
R826 vp_p.n1043 vp_p.t4 756.008
R827 vp_p.n1043 vp_p.t1368 756.008
R828 vp_p.n1041 vp_p.t232 756.008
R829 vp_p.n1041 vp_p.t99 756.008
R830 vp_p.n1039 vp_p.t1152 756.008
R831 vp_p.n1039 vp_p.t1016 756.008
R832 vp_p.n1037 vp_p.t1383 756.008
R833 vp_p.n1037 vp_p.t1263 756.008
R834 vp_p.n1035 vp_p.t979 756.008
R835 vp_p.n1035 vp_p.t851 756.008
R836 vp_p.n1033 vp_p.t1214 756.008
R837 vp_p.n1033 vp_p.t1095 756.008
R838 vp_p.n1031 vp_p.t795 756.008
R839 vp_p.n1031 vp_p.t674 756.008
R840 vp_p.n1029 vp_p.t231 756.008
R841 vp_p.n1029 vp_p.t100 756.008
R842 vp_p.n1027 vp_p.t459 756.008
R843 vp_p.n1027 vp_p.t348 756.008
R844 vp_p.n1025 vp_p.t57 756.008
R845 vp_p.n1025 vp_p.t1433 756.008
R846 vp_p.n1023 vp_p.t294 756.008
R847 vp_p.n1023 vp_p.t172 756.008
R848 vp_p.n1021 vp_p.t1378 756.008
R849 vp_p.n1021 vp_p.t1257 756.008
R850 vp_p.n1019 vp_p.t1453 756.008
R851 vp_p.n1019 vp_p.t1328 756.008
R852 vp_p.n1017 vp_p.t1028 756.008
R853 vp_p.n1017 vp_p.t911 756.008
R854 vp_p.n1015 vp_p.t626 756.008
R855 vp_p.n1015 vp_p.t502 756.008
R856 vp_p.n1013 vp_p.t867 756.008
R857 vp_p.n1013 vp_p.t742 756.008
R858 vp_p.n1011 vp_p.t450 756.008
R859 vp_p.n1011 vp_p.t341 756.008
R860 vp_p.n1009 vp_p.t527 756.008
R861 vp_p.n1009 vp_p.t401 756.008
R862 vp_p.n1007 vp_p.t116 756.008
R863 vp_p.n1007 vp_p.t5 756.008
R864 vp_p.n1005 vp_p.t1210 756.008
R865 vp_p.n1005 vp_p.t1089 756.008
R866 vp_p.n1003 vp_p.t829 756.008
R867 vp_p.n1003 vp_p.t705 756.008
R868 vp_p.n1001 vp_p.t424 756.008
R869 vp_p.n1001 vp_p.t306 756.008
R870 vp_p.n999 vp_p.t493 756.008
R871 vp_p.n999 vp_p.t379 756.008
R872 vp_p.n997 vp_p.t83 756.008
R873 vp_p.n997 vp_p.t1467 756.008
R874 vp_p.n995 vp_p.t328 756.008
R875 vp_p.n995 vp_p.t205 756.008
R876 vp_p.n993 vp_p.t1416 756.008
R877 vp_p.n993 vp_p.t1299 756.008
R878 vp_p.n991 vp_p.t997 756.008
R879 vp_p.n991 vp_p.t882 756.008
R880 vp_p.n989 vp_p.t1072 756.008
R881 vp_p.n989 vp_p.t950 756.008
R882 vp_p.n987 vp_p.t654 756.008
R883 vp_p.n987 vp_p.t543 756.008
R884 vp_p.n985 vp_p.t900 756.008
R885 vp_p.n985 vp_p.t770 756.008
R886 vp_p.n983 vp_p.t487 756.008
R887 vp_p.n983 vp_p.t374 756.008
R888 vp_p.n981 vp_p.t80 756.008
R889 vp_p.n981 vp_p.t1464 756.008
R890 vp_p.n979 vp_p.t153 756.008
R891 vp_p.n979 vp_p.t35 756.008
R892 vp_p.n977 vp_p.t1238 756.008
R893 vp_p.n977 vp_p.t1119 756.008
R894 vp_p.n975 vp_p.t1486 756.008
R895 vp_p.n975 vp_p.t1349 756.008
R896 vp_p.n973 vp_p.t1065 756.008
R897 vp_p.n973 vp_p.t944 756.008
R898 vp_p.n972 vp_p.t1314 756.008
R899 vp_p.n972 vp_p.t1180 756.008
R900 vp_p.n1268 vp_p.t1446 756.008
R901 vp_p.n1268 vp_p.t1231 756.008
R902 vp_p.n1266 vp_p.t362 756.008
R903 vp_p.n1266 vp_p.t149 756.008
R904 vp_p.n1264 vp_p.t115 756.008
R905 vp_p.n1264 vp_p.t1409 756.008
R906 vp_p.n1262 vp_p.t525 756.008
R907 vp_p.n1262 vp_p.t319 756.008
R908 vp_p.n1260 vp_p.t934 756.008
R909 vp_p.n1260 vp_p.t719 756.008
R910 vp_p.n1258 vp_p.t866 756.008
R911 vp_p.n1258 vp_p.t649 756.008
R912 vp_p.n1256 vp_p.t1282 756.008
R913 vp_p.n1256 vp_p.t1062 756.008
R914 vp_p.n1254 vp_p.t1063 756.008
R915 vp_p.n1254 vp_p.t854 756.008
R916 vp_p.n1252 vp_p.t1485 756.008
R917 vp_p.n1252 vp_p.t1266 756.008
R918 vp_p.n1250 vp_p.t663 756.008
R919 vp_p.n1250 vp_p.t455 756.008
R920 vp_p.n1248 vp_p.t925 756.008
R921 vp_p.n1248 vp_p.t708 756.008
R922 vp_p.n1246 vp_p.t518 756.008
R923 vp_p.n1246 vp_p.t310 756.008
R924 vp_p.n1244 vp_p.t406 756.008
R925 vp_p.n1244 vp_p.t199 756.008
R926 vp_p.n1242 vp_p.t7 756.008
R927 vp_p.n1242 vp_p.t1296 756.008
R928 vp_p.n1240 vp_p.t236 756.008
R929 vp_p.n1240 vp_p.t30 756.008
R930 vp_p.n1238 vp_p.t1155 756.008
R931 vp_p.n1238 vp_p.t946 756.008
R932 vp_p.n1236 vp_p.t745 756.008
R933 vp_p.n1236 vp_p.t540 756.008
R934 vp_p.n1234 vp_p.t981 756.008
R935 vp_p.n1234 vp_p.t767 756.008
R936 vp_p.n1232 vp_p.t575 756.008
R937 vp_p.n1232 vp_p.t373 756.008
R938 vp_p.n1230 vp_p.t800 756.008
R939 vp_p.n1230 vp_p.t598 756.008
R940 vp_p.n1228 vp_p.t235 756.008
R941 vp_p.n1228 vp_p.t32 756.008
R942 vp_p.n1226 vp_p.t464 756.008
R943 vp_p.n1226 vp_p.t262 756.008
R944 vp_p.n1224 vp_p.t61 756.008
R945 vp_p.n1224 vp_p.t1347 756.008
R946 vp_p.n1222 vp_p.t1149 756.008
R947 vp_p.n1222 vp_p.t942 756.008
R948 vp_p.n1220 vp_p.t1382 756.008
R949 vp_p.n1220 vp_p.t1176 756.008
R950 vp_p.n1218 vp_p.t799 756.008
R951 vp_p.n1218 vp_p.t599 756.008
R952 vp_p.n1216 vp_p.t1032 756.008
R953 vp_p.n1216 vp_p.t828 756.008
R954 vp_p.n1214 vp_p.t630 756.008
R955 vp_p.n1214 vp_p.t423 756.008
R956 vp_p.n1212 vp_p.t230 756.008
R957 vp_p.n1212 vp_p.t29 756.008
R958 vp_p.n1210 vp_p.t457 756.008
R959 vp_p.n1210 vp_p.t256 756.008
R960 vp_p.n1208 vp_p.t1381 756.008
R961 vp_p.n1208 vp_p.t1177 756.008
R962 vp_p.n1206 vp_p.t122 756.008
R963 vp_p.n1206 vp_p.t1412 756.008
R964 vp_p.n1204 vp_p.t1213 756.008
R965 vp_p.n1204 vp_p.t996 756.008
R966 vp_p.n1202 vp_p.t1229 756.008
R967 vp_p.n1202 vp_p.t1010 756.008
R968 vp_p.n1200 vp_p.t816 756.008
R969 vp_p.n1200 vp_p.t617 756.008
R970 vp_p.n1198 vp_p.t252 756.008
R971 vp_p.n1198 vp_p.t50 756.008
R972 vp_p.n1196 vp_p.t479 756.008
R973 vp_p.n1196 vp_p.t278 756.008
R974 vp_p.n1194 vp_p.t73 756.008
R975 vp_p.n1194 vp_p.t1366 756.008
R976 vp_p.n1192 vp_p.t311 756.008
R977 vp_p.n1192 vp_p.t95 756.008
R978 vp_p.n1190 vp_p.t1401 756.008
R979 vp_p.n1190 vp_p.t1195 756.008
R980 vp_p.n1188 vp_p.t1473 756.008
R981 vp_p.n1188 vp_p.t1256 756.008
R982 vp_p.n1186 vp_p.t1052 756.008
R983 vp_p.n1186 vp_p.t846 756.008
R984 vp_p.n1184 vp_p.t641 756.008
R985 vp_p.n1184 vp_p.t438 756.008
R986 vp_p.n1182 vp_p.t886 756.008
R987 vp_p.n1182 vp_p.t671 756.008
R988 vp_p.n1180 vp_p.t472 756.008
R989 vp_p.n1180 vp_p.t276 756.008
R990 vp_p.n1178 vp_p.t549 756.008
R991 vp_p.n1178 vp_p.t340 756.008
R992 vp_p.n1176 vp_p.t139 756.008
R993 vp_p.n1176 vp_p.t1429 756.008
R994 vp_p.n1174 vp_p.t1223 756.008
R995 vp_p.n1174 vp_p.t1008 756.008
R996 vp_p.n1172 vp_p.t1466 756.008
R997 vp_p.n1172 vp_p.t1253 756.008
R998 vp_p.n1170 vp_p.t1044 756.008
R999 vp_p.n1170 vp_p.t843 756.008
R1000 vp_p.n1168 vp_p.t1123 756.008
R1001 vp_p.n1168 vp_p.t909 756.008
R1002 vp_p.n1166 vp_p.t704 756.008
R1003 vp_p.n1166 vp_p.t500 756.008
R1004 vp_p.n1164 vp_p.t949 756.008
R1005 vp_p.n1164 vp_p.t736 756.008
R1006 vp_p.n1162 vp_p.t542 756.008
R1007 vp_p.n1162 vp_p.t337 756.008
R1008 vp_p.n1160 vp_p.t133 756.008
R1009 vp_p.n1160 vp_p.t1428 756.008
R1010 vp_p.n1158 vp_p.t203 756.008
R1011 vp_p.n1158 vp_p.t0 756.008
R1012 vp_p.n1156 vp_p.t1297 756.008
R1013 vp_p.n1156 vp_p.t1085 756.008
R1014 vp_p.n1154 vp_p.t913 756.008
R1015 vp_p.n1154 vp_p.t703 756.008
R1016 vp_p.n1152 vp_p.t504 756.008
R1017 vp_p.n1152 vp_p.t304 756.008
R1018 vp_p.n1150 vp_p.t97 756.008
R1019 vp_p.n1150 vp_p.t1395 756.008
R1020 vp_p.n1148 vp_p.t173 756.008
R1021 vp_p.n1148 vp_p.t1463 756.008
R1022 vp_p.n1146 vp_p.t1258 756.008
R1023 vp_p.n1146 vp_p.t1041 756.008
R1024 vp_p.n1144 vp_p.t6 756.008
R1025 vp_p.n1144 vp_p.t1294 756.008
R1026 vp_p.n1142 vp_p.t1091 756.008
R1027 vp_p.n1142 vp_p.t880 756.008
R1028 vp_p.n1140 vp_p.t1324 756.008
R1029 vp_p.n1140 vp_p.t1115 756.008
R1030 vp_p.n1138 vp_p.t743 756.008
R1031 vp_p.n1138 vp_p.t538 756.008
R1032 vp_p.n1136 vp_p.t342 756.008
R1033 vp_p.n1136 vp_p.t130 756.008
R1034 vp_p.n1134 vp_p.t574 756.008
R1035 vp_p.n1134 vp_p.t372 756.008
R1036 vp_p.n1132 vp_p.t169 756.008
R1037 vp_p.n1132 vp_p.t1460 756.008
R1038 vp_p.n1130 vp_p.t398 756.008
R1039 vp_p.n1130 vp_p.t197 756.008
R1040 vp_p.n1128 vp_p.t1325 756.008
R1041 vp_p.n1128 vp_p.t1116 756.008
R1042 vp_p.n1126 vp_p.t58 756.008
R1043 vp_p.n1126 vp_p.t1345 756.008
R1044 vp_p.n1124 vp_p.t1147 756.008
R1045 vp_p.n1124 vp_p.t941 756.008
R1046 vp_p.n1122 vp_p.t738 756.008
R1047 vp_p.n1122 vp_p.t535 756.008
R1048 vp_p.n1121 vp_p.t976 756.008
R1049 vp_p.n1121 vp_p.t766 756.008
R1050 vp_p.n1417 vp_p.t1017 756.008
R1051 vp_p.n1417 vp_p.t458 756.008
R1052 vp_p.n1415 vp_p.t1443 756.008
R1053 vp_p.n1415 vp_p.t874 756.008
R1054 vp_p.n1413 vp_p.t358 756.008
R1055 vp_p.n1413 vp_p.t1289 756.008
R1056 vp_p.n1411 vp_p.t109 756.008
R1057 vp_p.n1411 vp_p.t1033 756.008
R1058 vp_p.n1409 vp_p.t519 756.008
R1059 vp_p.n1409 vp_p.t1457 756.008
R1060 vp_p.n1407 vp_p.t446 756.008
R1061 vp_p.n1407 vp_p.t1384 756.008
R1062 vp_p.n1405 vp_p.t860 756.008
R1063 vp_p.n1405 vp_p.t298 756.008
R1064 vp_p.n1403 vp_p.t1274 756.008
R1065 vp_p.n1403 vp_p.t697 756.008
R1066 vp_p.n1401 vp_p.t1054 756.008
R1067 vp_p.n1401 vp_p.t492 756.008
R1068 vp_p.n1399 vp_p.t1478 756.008
R1069 vp_p.n1399 vp_p.t904 756.008
R1070 vp_p.n1397 vp_p.t915 756.008
R1071 vp_p.n1397 vp_p.t364 756.008
R1072 vp_p.n1395 vp_p.t509 756.008
R1073 vp_p.n1395 vp_p.t1450 756.008
R1074 vp_p.n1393 vp_p.t399 756.008
R1075 vp_p.n1393 vp_p.t1336 756.008
R1076 vp_p.n1391 vp_p.t3 756.008
R1077 vp_p.n1391 vp_p.t922 756.008
R1078 vp_p.n1389 vp_p.t1088 756.008
R1079 vp_p.n1389 vp_p.t514 756.008
R1080 vp_p.n1387 vp_p.t1148 756.008
R1081 vp_p.n1387 vp_p.t587 756.008
R1082 vp_p.n1385 vp_p.t740 756.008
R1083 vp_p.n1385 vp_p.t183 756.008
R1084 vp_p.n1383 vp_p.t977 756.008
R1085 vp_p.n1383 vp_p.t411 756.008
R1086 vp_p.n1381 vp_p.t573 756.008
R1087 vp_p.n1381 vp_p.t16 756.008
R1088 vp_p.n1379 vp_p.t167 756.008
R1089 vp_p.n1379 vp_p.t1099 756.008
R1090 vp_p.n1377 vp_p.t229 756.008
R1091 vp_p.n1377 vp_p.t1163 756.008
R1092 vp_p.n1375 vp_p.t1323 756.008
R1093 vp_p.n1375 vp_p.t755 756.008
R1094 vp_p.n1373 vp_p.t56 756.008
R1095 vp_p.n1373 vp_p.t986 756.008
R1096 vp_p.n1371 vp_p.t1145 756.008
R1097 vp_p.n1371 vp_p.t583 756.008
R1098 vp_p.n1369 vp_p.t1376 756.008
R1099 vp_p.n1369 vp_p.t805 756.008
R1100 vp_p.n1367 vp_p.t794 756.008
R1101 vp_p.n1367 vp_p.t241 756.008
R1102 vp_p.n1365 vp_p.t397 756.008
R1103 vp_p.n1365 vp_p.t1331 756.008
R1104 vp_p.n1363 vp_p.t625 756.008
R1105 vp_p.n1363 vp_p.t64 756.008
R1106 vp_p.n1361 vp_p.t227 756.008
R1107 vp_p.n1361 vp_p.t1156 756.008
R1108 vp_p.n1359 vp_p.t448 756.008
R1109 vp_p.n1359 vp_p.t1387 756.008
R1110 vp_p.n1357 vp_p.t1377 756.008
R1111 vp_p.n1357 vp_p.t806 756.008
R1112 vp_p.n1355 vp_p.t113 756.008
R1113 vp_p.n1355 vp_p.t1035 756.008
R1114 vp_p.n1353 vp_p.t1208 756.008
R1115 vp_p.n1353 vp_p.t632 756.008
R1116 vp_p.n1351 vp_p.t792 756.008
R1117 vp_p.n1351 vp_p.t234 756.008
R1118 vp_p.n1349 vp_p.t812 756.008
R1119 vp_p.n1349 vp_p.t258 756.008
R1120 vp_p.n1347 vp_p.t249 756.008
R1121 vp_p.n1347 vp_p.t1178 756.008
R1122 vp_p.n1345 vp_p.t473 756.008
R1123 vp_p.n1345 vp_p.t1413 756.008
R1124 vp_p.n1343 vp_p.t70 756.008
R1125 vp_p.n1343 vp_p.t995 756.008
R1126 vp_p.n1341 vp_p.t1167 756.008
R1127 vp_p.n1341 vp_p.t596 756.008
R1128 vp_p.n1339 vp_p.t1397 756.008
R1129 vp_p.n1339 vp_p.t824 756.008
R1130 vp_p.n1337 vp_p.t813 756.008
R1131 vp_p.n1337 vp_p.t257 756.008
R1132 vp_p.n1335 vp_p.t1043 756.008
R1133 vp_p.n1335 vp_p.t486 756.008
R1134 vp_p.n1333 vp_p.t639 756.008
R1135 vp_p.n1333 vp_p.t78 756.008
R1136 vp_p.n1331 vp_p.t881 756.008
R1137 vp_p.n1331 vp_p.t318 756.008
R1138 vp_p.n1329 vp_p.t470 756.008
R1139 vp_p.n1329 vp_p.t1408 756.008
R1140 vp_p.n1327 vp_p.t1398 756.008
R1141 vp_p.n1327 vp_p.t823 756.008
R1142 vp_p.n1325 vp_p.t132 756.008
R1143 vp_p.n1325 vp_p.t1061 756.008
R1144 vp_p.n1323 vp_p.t1222 756.008
R1145 vp_p.n1323 vp_p.t647 756.008
R1146 vp_p.n1321 vp_p.t1462 756.008
R1147 vp_p.n1321 vp_p.t895 756.008
R1148 vp_p.n1319 vp_p.t1039 756.008
R1149 vp_p.n1319 vp_p.t481 756.008
R1150 vp_p.n1317 vp_p.t1118 756.008
R1151 vp_p.n1317 vp_p.t558 756.008
R1152 vp_p.n1315 vp_p.t702 756.008
R1153 vp_p.n1315 vp_p.t147 756.008
R1154 vp_p.n1313 vp_p.t303 756.008
R1155 vp_p.n1313 vp_p.t1230 756.008
R1156 vp_p.n1311 vp_p.t537 756.008
R1157 vp_p.n1311 vp_p.t1476 756.008
R1158 vp_p.n1309 vp_p.t129 756.008
R1159 vp_p.n1309 vp_p.t1053 756.008
R1160 vp_p.n1307 vp_p.t198 756.008
R1161 vp_p.n1307 vp_p.t1129 756.008
R1162 vp_p.n1305 vp_p.t1293 756.008
R1163 vp_p.n1305 vp_p.t712 756.008
R1164 vp_p.n1303 vp_p.t879 756.008
R1165 vp_p.n1303 vp_p.t312 756.008
R1166 vp_p.n1301 vp_p.t501 756.008
R1167 vp_p.n1301 vp_p.t1442 756.008
R1168 vp_p.n1299 vp_p.t94 756.008
R1169 vp_p.n1299 vp_p.t1018 756.008
R1170 vp_p.n1297 vp_p.t168 756.008
R1171 vp_p.n1297 vp_p.t1105 756.008
R1172 vp_p.n1295 vp_p.t1254 756.008
R1173 vp_p.n1295 vp_p.t684 756.008
R1174 vp_p.n1293 vp_p.t1 756.008
R1175 vp_p.n1293 vp_p.t921 756.008
R1176 vp_p.n1291 vp_p.t1086 756.008
R1177 vp_p.n1291 vp_p.t511 756.008
R1178 vp_p.n1289 vp_p.t669 756.008
R1179 vp_p.n1289 vp_p.t101 756.008
R1180 vp_p.n1287 vp_p.t737 756.008
R1181 vp_p.n1287 vp_p.t182 756.008
R1182 vp_p.n1285 vp_p.t338 756.008
R1183 vp_p.n1285 vp_p.t1267 756.008
R1184 vp_p.n1283 vp_p.t572 756.008
R1185 vp_p.n1283 vp_p.t14 756.008
R1186 vp_p.n1281 vp_p.t165 756.008
R1187 vp_p.n1281 vp_p.t1097 756.008
R1188 vp_p.n1279 vp_p.t1251 756.008
R1189 vp_p.n1279 vp_p.t675 756.008
R1190 vp_p.n1277 vp_p.t1321 756.008
R1191 vp_p.n1277 vp_p.t753 756.008
R1192 vp_p.n1275 vp_p.t907 756.008
R1193 vp_p.n1275 vp_p.t349 756.008
R1194 vp_p.n1273 vp_p.t1144 756.008
R1195 vp_p.n1273 vp_p.t582 756.008
R1196 vp_p.n1271 vp_p.t734 756.008
R1197 vp_p.n1271 vp_p.t175 756.008
R1198 vp_p.n1270 vp_p.t974 756.008
R1199 vp_p.n1270 vp_p.t405 756.008
R1200 vp_p.n670 vp_p.t1187 706.013
R1201 vp_p.n0 vp_p.t576 706.013
R1202 vp_p.n1419 vp_p.t206 706.013
R1203 vp_p.n749 vp_p.t376 705.989
R1204 vp_p.n743 vp_p.t1246 704.872
R1205 vp_p.n742 vp_p.t161 704.872
R1206 vp_p.n741 vp_p.t570 704.872
R1207 vp_p.n740 vp_p.t335 704.872
R1208 vp_p.n739 vp_p.t733 704.872
R1209 vp_p.n738 vp_p.t665 704.872
R1210 vp_p.n737 vp_p.t1083 704.872
R1211 vp_p.n736 vp_p.t1498 704.872
R1212 vp_p.n735 vp_p.t1288 704.872
R1213 vp_p.n734 vp_p.t195 704.872
R1214 vp_p.n733 vp_p.t1140 704.872
R1215 vp_p.n732 vp_p.t727 704.872
R1216 vp_p.n731 vp_p.t614 704.872
R1217 vp_p.n730 vp_p.t217 704.872
R1218 vp_p.n729 vp_p.t1313 704.872
R1219 vp_p.n728 vp_p.t1364 704.872
R1220 vp_p.n727 vp_p.t965 704.872
R1221 vp_p.n726 vp_p.t1192 704.872
R1222 vp_p.n725 vp_p.t780 704.872
R1223 vp_p.n724 vp_p.t387 704.872
R1224 vp_p.n723 vp_p.t435 704.872
R1225 vp_p.n722 vp_p.t45 704.872
R1226 vp_p.n721 vp_p.t274 704.872
R1227 vp_p.n720 vp_p.t1361 704.872
R1228 vp_p.n719 vp_p.t89 704.872
R1229 vp_p.n718 vp_p.t1007 704.872
R1230 vp_p.n717 vp_p.t612 704.872
R1231 vp_p.n716 vp_p.t841 704.872
R1232 vp_p.n715 vp_p.t432 704.872
R1233 vp_p.n714 vp_p.t666 704.872
R1234 vp_p.n713 vp_p.t90 704.872
R1235 vp_p.n712 vp_p.t336 704.872
R1236 vp_p.n711 vp_p.t1427 704.872
R1237 vp_p.n710 vp_p.t1006 704.872
R1238 vp_p.n709 vp_p.t1024 704.872
R1239 vp_p.n708 vp_p.t451 704.872
R1240 vp_p.n707 vp_p.t689 704.872
R1241 vp_p.n706 vp_p.t293 704.872
R1242 vp_p.n705 vp_p.t1375 704.872
R1243 vp_p.n704 vp_p.t110 704.872
R1244 vp_p.n703 vp_p.t1023 704.872
R1245 vp_p.n702 vp_p.t1278 704.872
R1246 vp_p.n701 vp_p.t862 704.872
R1247 vp_p.n700 vp_p.t1107 704.872
R1248 vp_p.n699 vp_p.t686 704.872
R1249 vp_p.n698 vp_p.t111 704.872
R1250 vp_p.n697 vp_p.t359 704.872
R1251 vp_p.n696 vp_p.t1445 704.872
R1252 vp_p.n695 vp_p.t184 704.872
R1253 vp_p.n694 vp_p.t1271 704.872
R1254 vp_p.n693 vp_p.t1337 704.872
R1255 vp_p.n692 vp_p.t924 704.872
R1256 vp_p.n691 vp_p.t517 704.872
R1257 vp_p.n690 vp_p.t754 704.872
R1258 vp_p.n689 vp_p.t352 704.872
R1259 vp_p.n688 vp_p.t412 704.872
R1260 vp_p.n687 vp_p.t18 704.872
R1261 vp_p.n686 vp_p.t1101 704.872
R1262 vp_p.n685 vp_p.t718 704.872
R1263 vp_p.n684 vp_p.t317 704.872
R1264 vp_p.n683 vp_p.t389 704.872
R1265 vp_p.n682 vp_p.t1484 704.872
R1266 vp_p.n681 vp_p.t213 704.872
R1267 vp_p.n680 vp_p.t1310 704.872
R1268 vp_p.n679 vp_p.t894 704.872
R1269 vp_p.n678 vp_p.t962 704.872
R1270 vp_p.n677 vp_p.t556 704.872
R1271 vp_p.n676 vp_p.t778 704.872
R1272 vp_p.n675 vp_p.t385 704.872
R1273 vp_p.n674 vp_p.t1475 704.872
R1274 vp_p.n673 vp_p.t43 704.872
R1275 vp_p.n672 vp_p.t1128 704.872
R1276 vp_p.n671 vp_p.t1359 704.872
R1277 vp_p.n670 vp_p.t955 704.872
R1278 vp_p.n0 vp_p.t347 704.872
R1279 vp_p.n1 vp_p.t748 704.872
R1280 vp_p.n2 vp_p.t1157 704.872
R1281 vp_p.n3 vp_p.t919 704.872
R1282 vp_p.n4 vp_p.t11 704.872
R1283 vp_p.n5 vp_p.t1261 704.872
R1284 vp_p.n6 vp_p.t176 704.872
R1285 vp_p.n7 vp_p.t1440 704.872
R1286 vp_p.n8 vp_p.t354 704.872
R1287 vp_p.n9 vp_p.t916 704.872
R1288 vp_p.n10 vp_p.t679 704.872
R1289 vp_p.n11 vp_p.t1103 704.872
R1290 vp_p.n12 vp_p.t858 704.872
R1291 vp_p.n13 vp_p.t1270 704.872
R1292 vp_p.n14 vp_p.t1203 704.872
R1293 vp_p.n15 vp_p.t106 704.872
R1294 vp_p.n16 vp_p.t515 704.872
R1295 vp_p.n17 vp_p.t891 704.872
R1296 vp_p.n18 vp_p.t1307 704.872
R1297 vp_p.n19 vp_p.t1227 704.872
R1298 vp_p.n20 vp_p.t143 704.872
R1299 vp_p.n21 vp_p.t553 704.872
R1300 vp_p.n22 vp_p.t315 704.872
R1301 vp_p.n23 vp_p.t715 704.872
R1302 vp_p.n24 vp_p.t646 704.872
R1303 vp_p.n25 vp_p.t1057 704.872
R1304 vp_p.n26 vp_p.t820 704.872
R1305 vp_p.n27 vp_p.t1234 704.872
R1306 vp_p.n28 vp_p.t150 704.872
R1307 vp_p.n29 vp_p.t76 704.872
R1308 vp_p.n30 vp_p.t483 704.872
R1309 vp_p.n31 vp_p.t255 704.872
R1310 vp_p.n32 vp_p.t650 704.872
R1311 vp_p.n33 vp_p.t1064 704.872
R1312 vp_p.n34 vp_p.t994 704.872
R1313 vp_p.n35 vp_p.t1410 704.872
R1314 vp_p.n36 vp_p.t1175 704.872
R1315 vp_p.n37 vp_p.t79 704.872
R1316 vp_p.n38 vp_p.t1346 704.872
R1317 vp_p.n39 vp_p.t422 704.872
R1318 vp_p.n40 vp_p.t825 704.872
R1319 vp_p.n41 vp_p.t804 704.872
R1320 vp_p.n42 vp_p.t1219 704.872
R1321 vp_p.n43 vp_p.t984 704.872
R1322 vp_p.n44 vp_p.t62 704.872
R1323 vp_p.n45 vp_p.t1330 704.872
R1324 vp_p.n46 vp_p.t239 704.872
R1325 vp_p.n47 vp_p.t634 704.872
R1326 vp_p.n48 vp_p.t408 704.872
R1327 vp_p.n49 vp_p.t985 704.872
R1328 vp_p.n50 vp_p.t751 704.872
R1329 vp_p.n51 vp_p.t1160 704.872
R1330 vp_p.n52 vp_p.t66 704.872
R1331 vp_p.n53 vp_p.t1335 704.872
R1332 vp_p.n54 vp_p.t409 704.872
R1333 vp_p.n55 vp_p.t181 704.872
R1334 vp_p.n56 vp_p.t585 704.872
R1335 vp_p.n57 vp_p.t357 704.872
R1336 vp_p.n58 vp_p.t757 704.872
R1337 vp_p.n59 vp_p.t1334 704.872
R1338 vp_p.n60 vp_p.t1106 704.872
R1339 vp_p.n61 vp_p.t19 704.872
R1340 vp_p.n62 vp_p.t117 704.872
R1341 vp_p.n63 vp_p.t526 704.872
R1342 vp_p.n64 vp_p.t273 704.872
R1343 vp_p.n65 vp_p.t1075 704.872
R1344 vp_p.n66 vp_p.t658 704.872
R1345 vp_p.n67 vp_p.t876 704.872
R1346 vp_p.n68 vp_p.t463 704.872
R1347 vp_p.n69 vp_p.t533 704.872
R1348 vp_p.n70 vp_p.t126 704.872
R1349 vp_p.n71 vp_p.t1218 704.872
R1350 vp_p.n72 vp_p.t1455 704.872
R1351 vp_p.n73 vp_p.t1031 704.872
R1352 vp_p.n749 vp_p.t135 704.872
R1353 vp_p.n750 vp_p.t544 704.872
R1354 vp_p.n751 vp_p.t307 704.872
R1355 vp_p.n752 vp_p.t706 704.872
R1356 vp_p.n753 vp_p.t640 704.872
R1357 vp_p.n754 vp_p.t1047 704.872
R1358 vp_p.n755 vp_p.t1469 704.872
R1359 vp_p.n756 vp_p.t1226 704.872
R1360 vp_p.n757 vp_p.t141 704.872
R1361 vp_p.n758 vp_p.t72 704.872
R1362 vp_p.n759 vp_p.t476 704.872
R1363 vp_p.n760 vp_p.t889 704.872
R1364 vp_p.n761 vp_p.t644 704.872
R1365 vp_p.n762 vp_p.t1056 704.872
R1366 vp_p.n763 vp_p.t992 704.872
R1367 vp_p.n764 vp_p.t1404 704.872
R1368 vp_p.n765 vp_p.t281 704.872
R1369 vp_p.n766 vp_p.t676 704.872
R1370 vp_p.n767 vp_p.t1098 704.872
R1371 vp_p.n768 vp_p.t1012 704.872
R1372 vp_p.n769 vp_p.t1435 704.872
R1373 vp_p.n770 vp_p.t1200 704.872
R1374 vp_p.n771 vp_p.t103 704.872
R1375 vp_p.n772 vp_p.t512 704.872
R1376 vp_p.n773 vp_p.t440 704.872
R1377 vp_p.n774 vp_p.t853 704.872
R1378 vp_p.n775 vp_p.t620 704.872
R1379 vp_p.n776 vp_p.t1019 704.872
R1380 vp_p.n777 vp_p.t790 704.872
R1381 vp_p.n778 vp_p.t1370 704.872
R1382 vp_p.n779 vp_p.t286 704.872
R1383 vp_p.n780 vp_p.t52 704.872
R1384 vp_p.n781 vp_p.t445 704.872
R1385 vp_p.n782 vp_p.t226 704.872
R1386 vp_p.n783 vp_p.t791 704.872
R1387 vp_p.n784 vp_p.t571 704.872
R1388 vp_p.n785 vp_p.t972 704.872
R1389 vp_p.n786 vp_p.t1373 704.872
R1390 vp_p.n787 vp_p.t1143 704.872
R1391 vp_p.n788 vp_p.t225 704.872
R1392 vp_p.n789 vp_p.t204 704.872
R1393 vp_p.n790 vp_p.t604 704.872
R1394 vp_p.n791 vp_p.t1004 704.872
R1395 vp_p.n792 vp_p.t772 704.872
R1396 vp_p.n793 vp_p.t1354 704.872
R1397 vp_p.n794 vp_p.t1122 704.872
R1398 vp_p.n795 vp_p.t37 704.872
R1399 vp_p.n796 vp_p.t1303 704.872
R1400 vp_p.n797 vp_p.t209 704.872
R1401 vp_p.n798 vp_p.t773 704.872
R1402 vp_p.n799 vp_p.t547 704.872
R1403 vp_p.n800 vp_p.t956 704.872
R1404 vp_p.n801 vp_p.t711 704.872
R1405 vp_p.n802 vp_p.t1126 704.872
R1406 vp_p.n803 vp_p.t1049 704.872
R1407 vp_p.n804 vp_p.t1474 704.872
R1408 vp_p.n805 vp_p.t384 704.872
R1409 vp_p.n806 vp_p.t145 704.872
R1410 vp_p.n807 vp_p.t557 704.872
R1411 vp_p.n808 vp_p.t480 704.872
R1412 vp_p.n809 vp_p.t892 704.872
R1413 vp_p.n810 vp_p.t1308 704.872
R1414 vp_p.n811 vp_p.t1414 704.872
R1415 vp_p.n812 vp_p.t324 704.872
R1416 vp_p.n813 vp_p.t870 704.872
R1417 vp_p.n814 vp_p.t453 704.872
R1418 vp_p.n815 vp_p.t662 704.872
R1419 vp_p.n816 vp_p.t264 704.872
R1420 vp_p.n817 vp_p.t1350 704.872
R1421 vp_p.n818 vp_p.t1423 704.872
R1422 vp_p.n819 vp_p.t1000 704.872
R1423 vp_p.n820 vp_p.t1244 704.872
R1424 vp_p.n821 vp_p.t832 704.872
R1425 vp_p.n822 vp_p.t425 704.872
R1426 vp_p.n1419 vp_p.t1468 704.872
R1427 vp_p.n1420 vp_p.t381 704.872
R1428 vp_p.n1421 vp_p.t776 704.872
R1429 vp_p.n1422 vp_p.t552 704.872
R1430 vp_p.n1423 vp_p.t1124 704.872
R1431 vp_p.n1424 vp_p.t887 704.872
R1432 vp_p.n1425 vp_p.t1305 704.872
R1433 vp_p.n1426 vp_p.t1055 704.872
R1434 vp_p.n1427 vp_p.t1479 704.872
R1435 vp_p.n1428 vp_p.t551 704.872
R1436 vp_p.n1429 vp_p.t313 704.872
R1437 vp_p.n1430 vp_p.t713 704.872
R1438 vp_p.n1431 vp_p.t482 704.872
R1439 vp_p.n1432 vp_p.t896 704.872
R1440 vp_p.n1433 vp_p.t818 704.872
R1441 vp_p.n1434 vp_p.t1232 704.872
R1442 vp_p.n1435 vp_p.t148 704.872
R1443 vp_p.n1436 vp_p.t510 704.872
R1444 vp_p.n1437 vp_p.t920 704.872
R1445 vp_p.n1438 vp_p.t852 704.872
R1446 vp_p.n1439 vp_p.t1265 704.872
R1447 vp_p.n1440 vp_p.t180 704.872
R1448 vp_p.n1441 vp_p.t1441 704.872
R1449 vp_p.n1442 vp_p.t356 704.872
R1450 vp_p.n1443 vp_p.t285 704.872
R1451 vp_p.n1444 vp_p.t683 704.872
R1452 vp_p.n1445 vp_p.t444 704.872
R1453 vp_p.n1446 vp_p.t859 704.872
R1454 vp_p.n1447 vp_p.t1273 704.872
R1455 vp_p.n1448 vp_p.t1204 704.872
R1456 vp_p.n1449 vp_p.t108 704.872
R1457 vp_p.n1450 vp_p.t1372 704.872
R1458 vp_p.n1451 vp_p.t289 704.872
R1459 vp_p.n1452 vp_p.t687 704.872
R1460 vp_p.n1453 vp_p.t622 704.872
R1461 vp_p.n1454 vp_p.t1022 704.872
R1462 vp_p.n1455 vp_p.t793 704.872
R1463 vp_p.n1456 vp_p.t1207 704.872
R1464 vp_p.n1457 vp_p.t975 704.872
R1465 vp_p.n1458 vp_p.t54 704.872
R1466 vp_p.n1459 vp_p.t449 704.872
R1467 vp_p.n1460 vp_p.t430 704.872
R1468 vp_p.n1461 vp_p.t839 704.872
R1469 vp_p.n1462 vp_p.t610 704.872
R1470 vp_p.n1463 vp_p.t1185 704.872
R1471 vp_p.n1464 vp_p.t953 704.872
R1472 vp_p.n1465 vp_p.t1357 704.872
R1473 vp_p.n1466 vp_p.t272 704.872
R1474 vp_p.n1467 vp_p.t42 704.872
R1475 vp_p.n1468 vp_p.t609 704.872
R1476 vp_p.n1469 vp_p.t382 704.872
R1477 vp_p.n1470 vp_p.t777 704.872
R1478 vp_p.n1471 vp_p.t1191 704.872
R1479 vp_p.n1472 vp_p.t960 704.872
R1480 vp_p.n1473 vp_p.t41 704.872
R1481 vp_p.n1474 vp_p.t1306 704.872
R1482 vp_p.n1475 vp_p.t212 704.872
R1483 vp_p.n1476 vp_p.t1480 704.872
R1484 vp_p.n1477 vp_p.t388 704.872
R1485 vp_p.n1478 vp_p.t959 704.872
R1486 vp_p.n1479 vp_p.t714 704.872
R1487 vp_p.n1480 vp_p.t1131 704.872
R1488 vp_p.n1481 vp_p.t1241 704.872
R1489 vp_p.n1482 vp_p.t155 704.872
R1490 vp_p.n1483 vp_p.t1390 704.872
R1491 vp_p.n1484 vp_p.t694 704.872
R1492 vp_p.n1485 vp_p.t295 704.872
R1493 vp_p.n1486 vp_p.t495 704.872
R1494 vp_p.n1487 vp_p.t87 704.872
R1495 vp_p.n1488 vp_p.t162 704.872
R1496 vp_p.n1489 vp_p.t1247 704.872
R1497 vp_p.n1490 vp_p.t836 704.872
R1498 vp_p.n1491 vp_p.t1079 704.872
R1499 vp_p.n1492 vp_p.t660 704.872
R1500 vp_p.n1493 vp_p.n1492 1.225
R1501 vp_p.n671 vp_p.n670 1.141
R1502 vp_p.n672 vp_p.n671 1.141
R1503 vp_p.n673 vp_p.n672 1.141
R1504 vp_p.n674 vp_p.n673 1.141
R1505 vp_p.n675 vp_p.n674 1.141
R1506 vp_p.n676 vp_p.n675 1.141
R1507 vp_p.n677 vp_p.n676 1.141
R1508 vp_p.n678 vp_p.n677 1.141
R1509 vp_p.n679 vp_p.n678 1.141
R1510 vp_p.n680 vp_p.n679 1.141
R1511 vp_p.n681 vp_p.n680 1.141
R1512 vp_p.n682 vp_p.n681 1.141
R1513 vp_p.n683 vp_p.n682 1.141
R1514 vp_p.n684 vp_p.n683 1.141
R1515 vp_p.n685 vp_p.n684 1.141
R1516 vp_p.n686 vp_p.n685 1.141
R1517 vp_p.n687 vp_p.n686 1.141
R1518 vp_p.n688 vp_p.n687 1.141
R1519 vp_p.n689 vp_p.n688 1.141
R1520 vp_p.n690 vp_p.n689 1.141
R1521 vp_p.n691 vp_p.n690 1.141
R1522 vp_p.n692 vp_p.n691 1.141
R1523 vp_p.n693 vp_p.n692 1.141
R1524 vp_p.n694 vp_p.n693 1.141
R1525 vp_p.n695 vp_p.n694 1.141
R1526 vp_p.n696 vp_p.n695 1.141
R1527 vp_p.n697 vp_p.n696 1.141
R1528 vp_p.n698 vp_p.n697 1.141
R1529 vp_p.n699 vp_p.n698 1.141
R1530 vp_p.n700 vp_p.n699 1.141
R1531 vp_p.n701 vp_p.n700 1.141
R1532 vp_p.n702 vp_p.n701 1.141
R1533 vp_p.n703 vp_p.n702 1.141
R1534 vp_p.n704 vp_p.n703 1.141
R1535 vp_p.n705 vp_p.n704 1.141
R1536 vp_p.n706 vp_p.n705 1.141
R1537 vp_p.n707 vp_p.n706 1.141
R1538 vp_p.n708 vp_p.n707 1.141
R1539 vp_p.n709 vp_p.n708 1.141
R1540 vp_p.n710 vp_p.n709 1.141
R1541 vp_p.n711 vp_p.n710 1.141
R1542 vp_p.n712 vp_p.n711 1.141
R1543 vp_p.n713 vp_p.n712 1.141
R1544 vp_p.n714 vp_p.n713 1.141
R1545 vp_p.n715 vp_p.n714 1.141
R1546 vp_p.n716 vp_p.n715 1.141
R1547 vp_p.n717 vp_p.n716 1.141
R1548 vp_p.n718 vp_p.n717 1.141
R1549 vp_p.n719 vp_p.n718 1.141
R1550 vp_p.n720 vp_p.n719 1.141
R1551 vp_p.n721 vp_p.n720 1.141
R1552 vp_p.n722 vp_p.n721 1.141
R1553 vp_p.n723 vp_p.n722 1.141
R1554 vp_p.n724 vp_p.n723 1.141
R1555 vp_p.n725 vp_p.n724 1.141
R1556 vp_p.n726 vp_p.n725 1.141
R1557 vp_p.n727 vp_p.n726 1.141
R1558 vp_p.n728 vp_p.n727 1.141
R1559 vp_p.n729 vp_p.n728 1.141
R1560 vp_p.n730 vp_p.n729 1.141
R1561 vp_p.n731 vp_p.n730 1.141
R1562 vp_p.n732 vp_p.n731 1.141
R1563 vp_p.n733 vp_p.n732 1.141
R1564 vp_p.n734 vp_p.n733 1.141
R1565 vp_p.n735 vp_p.n734 1.141
R1566 vp_p.n736 vp_p.n735 1.141
R1567 vp_p.n737 vp_p.n736 1.141
R1568 vp_p.n738 vp_p.n737 1.141
R1569 vp_p.n739 vp_p.n738 1.141
R1570 vp_p.n740 vp_p.n739 1.141
R1571 vp_p.n741 vp_p.n740 1.141
R1572 vp_p.n742 vp_p.n741 1.141
R1573 vp_p.n743 vp_p.n742 1.141
R1574 vp_p.n1 vp_p.n0 1.141
R1575 vp_p.n2 vp_p.n1 1.141
R1576 vp_p.n3 vp_p.n2 1.141
R1577 vp_p.n4 vp_p.n3 1.141
R1578 vp_p.n5 vp_p.n4 1.141
R1579 vp_p.n6 vp_p.n5 1.141
R1580 vp_p.n7 vp_p.n6 1.141
R1581 vp_p.n8 vp_p.n7 1.141
R1582 vp_p.n9 vp_p.n8 1.141
R1583 vp_p.n10 vp_p.n9 1.141
R1584 vp_p.n11 vp_p.n10 1.141
R1585 vp_p.n12 vp_p.n11 1.141
R1586 vp_p.n13 vp_p.n12 1.141
R1587 vp_p.n14 vp_p.n13 1.141
R1588 vp_p.n15 vp_p.n14 1.141
R1589 vp_p.n16 vp_p.n15 1.141
R1590 vp_p.n17 vp_p.n16 1.141
R1591 vp_p.n18 vp_p.n17 1.141
R1592 vp_p.n19 vp_p.n18 1.141
R1593 vp_p.n20 vp_p.n19 1.141
R1594 vp_p.n21 vp_p.n20 1.141
R1595 vp_p.n22 vp_p.n21 1.141
R1596 vp_p.n23 vp_p.n22 1.141
R1597 vp_p.n24 vp_p.n23 1.141
R1598 vp_p.n25 vp_p.n24 1.141
R1599 vp_p.n26 vp_p.n25 1.141
R1600 vp_p.n27 vp_p.n26 1.141
R1601 vp_p.n28 vp_p.n27 1.141
R1602 vp_p.n29 vp_p.n28 1.141
R1603 vp_p.n30 vp_p.n29 1.141
R1604 vp_p.n31 vp_p.n30 1.141
R1605 vp_p.n32 vp_p.n31 1.141
R1606 vp_p.n33 vp_p.n32 1.141
R1607 vp_p.n34 vp_p.n33 1.141
R1608 vp_p.n35 vp_p.n34 1.141
R1609 vp_p.n36 vp_p.n35 1.141
R1610 vp_p.n37 vp_p.n36 1.141
R1611 vp_p.n38 vp_p.n37 1.141
R1612 vp_p.n39 vp_p.n38 1.141
R1613 vp_p.n40 vp_p.n39 1.141
R1614 vp_p.n41 vp_p.n40 1.141
R1615 vp_p.n42 vp_p.n41 1.141
R1616 vp_p.n43 vp_p.n42 1.141
R1617 vp_p.n44 vp_p.n43 1.141
R1618 vp_p.n45 vp_p.n44 1.141
R1619 vp_p.n46 vp_p.n45 1.141
R1620 vp_p.n47 vp_p.n46 1.141
R1621 vp_p.n48 vp_p.n47 1.141
R1622 vp_p.n49 vp_p.n48 1.141
R1623 vp_p.n50 vp_p.n49 1.141
R1624 vp_p.n51 vp_p.n50 1.141
R1625 vp_p.n52 vp_p.n51 1.141
R1626 vp_p.n53 vp_p.n52 1.141
R1627 vp_p.n54 vp_p.n53 1.141
R1628 vp_p.n55 vp_p.n54 1.141
R1629 vp_p.n56 vp_p.n55 1.141
R1630 vp_p.n57 vp_p.n56 1.141
R1631 vp_p.n58 vp_p.n57 1.141
R1632 vp_p.n59 vp_p.n58 1.141
R1633 vp_p.n60 vp_p.n59 1.141
R1634 vp_p.n61 vp_p.n60 1.141
R1635 vp_p.n62 vp_p.n61 1.141
R1636 vp_p.n63 vp_p.n62 1.141
R1637 vp_p.n64 vp_p.n63 1.141
R1638 vp_p.n65 vp_p.n64 1.141
R1639 vp_p.n66 vp_p.n65 1.141
R1640 vp_p.n67 vp_p.n66 1.141
R1641 vp_p.n68 vp_p.n67 1.141
R1642 vp_p.n69 vp_p.n68 1.141
R1643 vp_p.n70 vp_p.n69 1.141
R1644 vp_p.n71 vp_p.n70 1.141
R1645 vp_p.n72 vp_p.n71 1.141
R1646 vp_p.n73 vp_p.n72 1.141
R1647 vp_p.n1420 vp_p.n1419 1.141
R1648 vp_p.n1421 vp_p.n1420 1.141
R1649 vp_p.n1422 vp_p.n1421 1.141
R1650 vp_p.n1423 vp_p.n1422 1.141
R1651 vp_p.n1424 vp_p.n1423 1.141
R1652 vp_p.n1425 vp_p.n1424 1.141
R1653 vp_p.n1426 vp_p.n1425 1.141
R1654 vp_p.n1427 vp_p.n1426 1.141
R1655 vp_p.n1428 vp_p.n1427 1.141
R1656 vp_p.n1429 vp_p.n1428 1.141
R1657 vp_p.n1430 vp_p.n1429 1.141
R1658 vp_p.n1431 vp_p.n1430 1.141
R1659 vp_p.n1432 vp_p.n1431 1.141
R1660 vp_p.n1433 vp_p.n1432 1.141
R1661 vp_p.n1434 vp_p.n1433 1.141
R1662 vp_p.n1435 vp_p.n1434 1.141
R1663 vp_p.n1436 vp_p.n1435 1.141
R1664 vp_p.n1437 vp_p.n1436 1.141
R1665 vp_p.n1438 vp_p.n1437 1.141
R1666 vp_p.n1439 vp_p.n1438 1.141
R1667 vp_p.n1440 vp_p.n1439 1.141
R1668 vp_p.n1441 vp_p.n1440 1.141
R1669 vp_p.n1442 vp_p.n1441 1.141
R1670 vp_p.n1443 vp_p.n1442 1.141
R1671 vp_p.n1444 vp_p.n1443 1.141
R1672 vp_p.n1445 vp_p.n1444 1.141
R1673 vp_p.n1446 vp_p.n1445 1.141
R1674 vp_p.n1447 vp_p.n1446 1.141
R1675 vp_p.n1448 vp_p.n1447 1.141
R1676 vp_p.n1449 vp_p.n1448 1.141
R1677 vp_p.n1450 vp_p.n1449 1.141
R1678 vp_p.n1451 vp_p.n1450 1.141
R1679 vp_p.n1452 vp_p.n1451 1.141
R1680 vp_p.n1453 vp_p.n1452 1.141
R1681 vp_p.n1454 vp_p.n1453 1.141
R1682 vp_p.n1455 vp_p.n1454 1.141
R1683 vp_p.n1456 vp_p.n1455 1.141
R1684 vp_p.n1457 vp_p.n1456 1.141
R1685 vp_p.n1458 vp_p.n1457 1.141
R1686 vp_p.n1459 vp_p.n1458 1.141
R1687 vp_p.n1460 vp_p.n1459 1.141
R1688 vp_p.n1461 vp_p.n1460 1.141
R1689 vp_p.n1462 vp_p.n1461 1.141
R1690 vp_p.n1463 vp_p.n1462 1.141
R1691 vp_p.n1464 vp_p.n1463 1.141
R1692 vp_p.n1465 vp_p.n1464 1.141
R1693 vp_p.n1466 vp_p.n1465 1.141
R1694 vp_p.n1467 vp_p.n1466 1.141
R1695 vp_p.n1468 vp_p.n1467 1.141
R1696 vp_p.n1469 vp_p.n1468 1.141
R1697 vp_p.n1470 vp_p.n1469 1.141
R1698 vp_p.n1471 vp_p.n1470 1.141
R1699 vp_p.n1472 vp_p.n1471 1.141
R1700 vp_p.n1473 vp_p.n1472 1.141
R1701 vp_p.n1474 vp_p.n1473 1.141
R1702 vp_p.n1475 vp_p.n1474 1.141
R1703 vp_p.n1476 vp_p.n1475 1.141
R1704 vp_p.n1477 vp_p.n1476 1.141
R1705 vp_p.n1478 vp_p.n1477 1.141
R1706 vp_p.n1479 vp_p.n1478 1.141
R1707 vp_p.n1480 vp_p.n1479 1.141
R1708 vp_p.n1481 vp_p.n1480 1.141
R1709 vp_p.n1482 vp_p.n1481 1.141
R1710 vp_p.n1483 vp_p.n1482 1.141
R1711 vp_p.n1484 vp_p.n1483 1.141
R1712 vp_p.n1485 vp_p.n1484 1.141
R1713 vp_p.n1486 vp_p.n1485 1.141
R1714 vp_p.n1487 vp_p.n1486 1.141
R1715 vp_p.n1488 vp_p.n1487 1.141
R1716 vp_p.n1489 vp_p.n1488 1.141
R1717 vp_p.n1490 vp_p.n1489 1.141
R1718 vp_p.n1491 vp_p.n1490 1.141
R1719 vp_p.n1492 vp_p.n1491 1.141
R1720 vp_p.n750 vp_p.n749 1.117
R1721 vp_p.n751 vp_p.n750 1.117
R1722 vp_p.n752 vp_p.n751 1.117
R1723 vp_p.n753 vp_p.n752 1.117
R1724 vp_p.n754 vp_p.n753 1.117
R1725 vp_p.n755 vp_p.n754 1.117
R1726 vp_p.n756 vp_p.n755 1.117
R1727 vp_p.n757 vp_p.n756 1.117
R1728 vp_p.n758 vp_p.n757 1.117
R1729 vp_p.n759 vp_p.n758 1.117
R1730 vp_p.n760 vp_p.n759 1.117
R1731 vp_p.n761 vp_p.n760 1.117
R1732 vp_p.n762 vp_p.n761 1.117
R1733 vp_p.n763 vp_p.n762 1.117
R1734 vp_p.n764 vp_p.n763 1.117
R1735 vp_p.n765 vp_p.n764 1.117
R1736 vp_p.n766 vp_p.n765 1.117
R1737 vp_p.n767 vp_p.n766 1.117
R1738 vp_p.n768 vp_p.n767 1.117
R1739 vp_p.n769 vp_p.n768 1.117
R1740 vp_p.n770 vp_p.n769 1.117
R1741 vp_p.n771 vp_p.n770 1.117
R1742 vp_p.n772 vp_p.n771 1.117
R1743 vp_p.n773 vp_p.n772 1.117
R1744 vp_p.n774 vp_p.n773 1.117
R1745 vp_p.n775 vp_p.n774 1.117
R1746 vp_p.n776 vp_p.n775 1.117
R1747 vp_p.n777 vp_p.n776 1.117
R1748 vp_p.n778 vp_p.n777 1.117
R1749 vp_p.n779 vp_p.n778 1.117
R1750 vp_p.n780 vp_p.n779 1.117
R1751 vp_p.n781 vp_p.n780 1.117
R1752 vp_p.n782 vp_p.n781 1.117
R1753 vp_p.n783 vp_p.n782 1.117
R1754 vp_p.n784 vp_p.n783 1.117
R1755 vp_p.n785 vp_p.n784 1.117
R1756 vp_p.n786 vp_p.n785 1.117
R1757 vp_p.n787 vp_p.n786 1.117
R1758 vp_p.n788 vp_p.n787 1.117
R1759 vp_p.n789 vp_p.n788 1.117
R1760 vp_p.n790 vp_p.n789 1.117
R1761 vp_p.n791 vp_p.n790 1.117
R1762 vp_p.n792 vp_p.n791 1.117
R1763 vp_p.n793 vp_p.n792 1.117
R1764 vp_p.n794 vp_p.n793 1.117
R1765 vp_p.n795 vp_p.n794 1.117
R1766 vp_p.n796 vp_p.n795 1.117
R1767 vp_p.n797 vp_p.n796 1.117
R1768 vp_p.n798 vp_p.n797 1.117
R1769 vp_p.n799 vp_p.n798 1.117
R1770 vp_p.n800 vp_p.n799 1.117
R1771 vp_p.n801 vp_p.n800 1.117
R1772 vp_p.n802 vp_p.n801 1.117
R1773 vp_p.n803 vp_p.n802 1.117
R1774 vp_p.n804 vp_p.n803 1.117
R1775 vp_p.n805 vp_p.n804 1.117
R1776 vp_p.n806 vp_p.n805 1.117
R1777 vp_p.n807 vp_p.n806 1.117
R1778 vp_p.n808 vp_p.n807 1.117
R1779 vp_p.n809 vp_p.n808 1.117
R1780 vp_p.n810 vp_p.n809 1.117
R1781 vp_p.n811 vp_p.n810 1.117
R1782 vp_p.n812 vp_p.n811 1.117
R1783 vp_p.n813 vp_p.n812 1.117
R1784 vp_p.n814 vp_p.n813 1.117
R1785 vp_p.n815 vp_p.n814 1.117
R1786 vp_p.n816 vp_p.n815 1.117
R1787 vp_p.n817 vp_p.n816 1.117
R1788 vp_p.n818 vp_p.n817 1.117
R1789 vp_p.n819 vp_p.n818 1.117
R1790 vp_p.n820 vp_p.n819 1.117
R1791 vp_p.n821 vp_p.n820 1.117
R1792 vp_p.n822 vp_p.n821 1.117
R1793 vp_p.n748 vp_p.n73 1.084
R1794 vp_p.n744 vp_p.n743 0.654
R1795 vp_p.n1497 vp_p.n822 0.509
R1796 vp_p.n523 vp_p.n521 0.356
R1797 vp_p.n374 vp_p.n372 0.356
R1798 vp_p.n225 vp_p.n223 0.356
R1799 vp_p.n76 vp_p.n74 0.356
R1800 vp_p.n825 vp_p.n823 0.356
R1801 vp_p.n974 vp_p.n972 0.356
R1802 vp_p.n1123 vp_p.n1121 0.356
R1803 vp_p.n1272 vp_p.n1270 0.356
R1804 vp_p.n744 vp_p.n669 0.319
R1805 vp_p.n746 vp_p.n371 0.319
R1806 vp_p.n1496 vp_p.n971 0.319
R1807 vp_p.n1494 vp_p.n1269 0.319
R1808 vp_p.n525 vp_p.n523 0.316
R1809 vp_p.n527 vp_p.n525 0.316
R1810 vp_p.n529 vp_p.n527 0.316
R1811 vp_p.n531 vp_p.n529 0.316
R1812 vp_p.n533 vp_p.n531 0.316
R1813 vp_p.n535 vp_p.n533 0.316
R1814 vp_p.n537 vp_p.n535 0.316
R1815 vp_p.n539 vp_p.n537 0.316
R1816 vp_p.n541 vp_p.n539 0.316
R1817 vp_p.n543 vp_p.n541 0.316
R1818 vp_p.n545 vp_p.n543 0.316
R1819 vp_p.n547 vp_p.n545 0.316
R1820 vp_p.n549 vp_p.n547 0.316
R1821 vp_p.n551 vp_p.n549 0.316
R1822 vp_p.n553 vp_p.n551 0.316
R1823 vp_p.n555 vp_p.n553 0.316
R1824 vp_p.n557 vp_p.n555 0.316
R1825 vp_p.n559 vp_p.n557 0.316
R1826 vp_p.n561 vp_p.n559 0.316
R1827 vp_p.n563 vp_p.n561 0.316
R1828 vp_p.n565 vp_p.n563 0.316
R1829 vp_p.n567 vp_p.n565 0.316
R1830 vp_p.n569 vp_p.n567 0.316
R1831 vp_p.n571 vp_p.n569 0.316
R1832 vp_p.n573 vp_p.n571 0.316
R1833 vp_p.n575 vp_p.n573 0.316
R1834 vp_p.n577 vp_p.n575 0.316
R1835 vp_p.n579 vp_p.n577 0.316
R1836 vp_p.n581 vp_p.n579 0.316
R1837 vp_p.n583 vp_p.n581 0.316
R1838 vp_p.n585 vp_p.n583 0.316
R1839 vp_p.n587 vp_p.n585 0.316
R1840 vp_p.n589 vp_p.n587 0.316
R1841 vp_p.n591 vp_p.n589 0.316
R1842 vp_p.n593 vp_p.n591 0.316
R1843 vp_p.n595 vp_p.n593 0.316
R1844 vp_p.n597 vp_p.n595 0.316
R1845 vp_p.n599 vp_p.n597 0.316
R1846 vp_p.n601 vp_p.n599 0.316
R1847 vp_p.n603 vp_p.n601 0.316
R1848 vp_p.n605 vp_p.n603 0.316
R1849 vp_p.n607 vp_p.n605 0.316
R1850 vp_p.n609 vp_p.n607 0.316
R1851 vp_p.n611 vp_p.n609 0.316
R1852 vp_p.n613 vp_p.n611 0.316
R1853 vp_p.n615 vp_p.n613 0.316
R1854 vp_p.n617 vp_p.n615 0.316
R1855 vp_p.n619 vp_p.n617 0.316
R1856 vp_p.n621 vp_p.n619 0.316
R1857 vp_p.n623 vp_p.n621 0.316
R1858 vp_p.n625 vp_p.n623 0.316
R1859 vp_p.n627 vp_p.n625 0.316
R1860 vp_p.n629 vp_p.n627 0.316
R1861 vp_p.n631 vp_p.n629 0.316
R1862 vp_p.n633 vp_p.n631 0.316
R1863 vp_p.n635 vp_p.n633 0.316
R1864 vp_p.n637 vp_p.n635 0.316
R1865 vp_p.n639 vp_p.n637 0.316
R1866 vp_p.n641 vp_p.n639 0.316
R1867 vp_p.n643 vp_p.n641 0.316
R1868 vp_p.n645 vp_p.n643 0.316
R1869 vp_p.n647 vp_p.n645 0.316
R1870 vp_p.n649 vp_p.n647 0.316
R1871 vp_p.n651 vp_p.n649 0.316
R1872 vp_p.n653 vp_p.n651 0.316
R1873 vp_p.n655 vp_p.n653 0.316
R1874 vp_p.n657 vp_p.n655 0.316
R1875 vp_p.n659 vp_p.n657 0.316
R1876 vp_p.n661 vp_p.n659 0.316
R1877 vp_p.n663 vp_p.n661 0.316
R1878 vp_p.n665 vp_p.n663 0.316
R1879 vp_p.n667 vp_p.n665 0.316
R1880 vp_p.n669 vp_p.n667 0.316
R1881 vp_p.n376 vp_p.n374 0.316
R1882 vp_p.n378 vp_p.n376 0.316
R1883 vp_p.n380 vp_p.n378 0.316
R1884 vp_p.n382 vp_p.n380 0.316
R1885 vp_p.n384 vp_p.n382 0.316
R1886 vp_p.n386 vp_p.n384 0.316
R1887 vp_p.n388 vp_p.n386 0.316
R1888 vp_p.n390 vp_p.n388 0.316
R1889 vp_p.n392 vp_p.n390 0.316
R1890 vp_p.n394 vp_p.n392 0.316
R1891 vp_p.n396 vp_p.n394 0.316
R1892 vp_p.n398 vp_p.n396 0.316
R1893 vp_p.n400 vp_p.n398 0.316
R1894 vp_p.n402 vp_p.n400 0.316
R1895 vp_p.n404 vp_p.n402 0.316
R1896 vp_p.n406 vp_p.n404 0.316
R1897 vp_p.n408 vp_p.n406 0.316
R1898 vp_p.n410 vp_p.n408 0.316
R1899 vp_p.n412 vp_p.n410 0.316
R1900 vp_p.n414 vp_p.n412 0.316
R1901 vp_p.n416 vp_p.n414 0.316
R1902 vp_p.n418 vp_p.n416 0.316
R1903 vp_p.n420 vp_p.n418 0.316
R1904 vp_p.n422 vp_p.n420 0.316
R1905 vp_p.n424 vp_p.n422 0.316
R1906 vp_p.n426 vp_p.n424 0.316
R1907 vp_p.n428 vp_p.n426 0.316
R1908 vp_p.n430 vp_p.n428 0.316
R1909 vp_p.n432 vp_p.n430 0.316
R1910 vp_p.n434 vp_p.n432 0.316
R1911 vp_p.n436 vp_p.n434 0.316
R1912 vp_p.n438 vp_p.n436 0.316
R1913 vp_p.n440 vp_p.n438 0.316
R1914 vp_p.n442 vp_p.n440 0.316
R1915 vp_p.n444 vp_p.n442 0.316
R1916 vp_p.n446 vp_p.n444 0.316
R1917 vp_p.n448 vp_p.n446 0.316
R1918 vp_p.n450 vp_p.n448 0.316
R1919 vp_p.n452 vp_p.n450 0.316
R1920 vp_p.n454 vp_p.n452 0.316
R1921 vp_p.n456 vp_p.n454 0.316
R1922 vp_p.n458 vp_p.n456 0.316
R1923 vp_p.n460 vp_p.n458 0.316
R1924 vp_p.n462 vp_p.n460 0.316
R1925 vp_p.n464 vp_p.n462 0.316
R1926 vp_p.n466 vp_p.n464 0.316
R1927 vp_p.n468 vp_p.n466 0.316
R1928 vp_p.n470 vp_p.n468 0.316
R1929 vp_p.n472 vp_p.n470 0.316
R1930 vp_p.n474 vp_p.n472 0.316
R1931 vp_p.n476 vp_p.n474 0.316
R1932 vp_p.n478 vp_p.n476 0.316
R1933 vp_p.n480 vp_p.n478 0.316
R1934 vp_p.n482 vp_p.n480 0.316
R1935 vp_p.n484 vp_p.n482 0.316
R1936 vp_p.n486 vp_p.n484 0.316
R1937 vp_p.n488 vp_p.n486 0.316
R1938 vp_p.n490 vp_p.n488 0.316
R1939 vp_p.n492 vp_p.n490 0.316
R1940 vp_p.n494 vp_p.n492 0.316
R1941 vp_p.n496 vp_p.n494 0.316
R1942 vp_p.n498 vp_p.n496 0.316
R1943 vp_p.n500 vp_p.n498 0.316
R1944 vp_p.n502 vp_p.n500 0.316
R1945 vp_p.n504 vp_p.n502 0.316
R1946 vp_p.n506 vp_p.n504 0.316
R1947 vp_p.n508 vp_p.n506 0.316
R1948 vp_p.n510 vp_p.n508 0.316
R1949 vp_p.n512 vp_p.n510 0.316
R1950 vp_p.n514 vp_p.n512 0.316
R1951 vp_p.n516 vp_p.n514 0.316
R1952 vp_p.n518 vp_p.n516 0.316
R1953 vp_p.n520 vp_p.n518 0.316
R1954 vp_p.n227 vp_p.n225 0.316
R1955 vp_p.n229 vp_p.n227 0.316
R1956 vp_p.n231 vp_p.n229 0.316
R1957 vp_p.n233 vp_p.n231 0.316
R1958 vp_p.n235 vp_p.n233 0.316
R1959 vp_p.n237 vp_p.n235 0.316
R1960 vp_p.n239 vp_p.n237 0.316
R1961 vp_p.n241 vp_p.n239 0.316
R1962 vp_p.n243 vp_p.n241 0.316
R1963 vp_p.n245 vp_p.n243 0.316
R1964 vp_p.n247 vp_p.n245 0.316
R1965 vp_p.n249 vp_p.n247 0.316
R1966 vp_p.n251 vp_p.n249 0.316
R1967 vp_p.n253 vp_p.n251 0.316
R1968 vp_p.n255 vp_p.n253 0.316
R1969 vp_p.n257 vp_p.n255 0.316
R1970 vp_p.n259 vp_p.n257 0.316
R1971 vp_p.n261 vp_p.n259 0.316
R1972 vp_p.n263 vp_p.n261 0.316
R1973 vp_p.n265 vp_p.n263 0.316
R1974 vp_p.n267 vp_p.n265 0.316
R1975 vp_p.n269 vp_p.n267 0.316
R1976 vp_p.n271 vp_p.n269 0.316
R1977 vp_p.n273 vp_p.n271 0.316
R1978 vp_p.n275 vp_p.n273 0.316
R1979 vp_p.n277 vp_p.n275 0.316
R1980 vp_p.n279 vp_p.n277 0.316
R1981 vp_p.n281 vp_p.n279 0.316
R1982 vp_p.n283 vp_p.n281 0.316
R1983 vp_p.n285 vp_p.n283 0.316
R1984 vp_p.n287 vp_p.n285 0.316
R1985 vp_p.n289 vp_p.n287 0.316
R1986 vp_p.n291 vp_p.n289 0.316
R1987 vp_p.n293 vp_p.n291 0.316
R1988 vp_p.n295 vp_p.n293 0.316
R1989 vp_p.n297 vp_p.n295 0.316
R1990 vp_p.n299 vp_p.n297 0.316
R1991 vp_p.n301 vp_p.n299 0.316
R1992 vp_p.n303 vp_p.n301 0.316
R1993 vp_p.n305 vp_p.n303 0.316
R1994 vp_p.n307 vp_p.n305 0.316
R1995 vp_p.n309 vp_p.n307 0.316
R1996 vp_p.n311 vp_p.n309 0.316
R1997 vp_p.n313 vp_p.n311 0.316
R1998 vp_p.n315 vp_p.n313 0.316
R1999 vp_p.n317 vp_p.n315 0.316
R2000 vp_p.n319 vp_p.n317 0.316
R2001 vp_p.n321 vp_p.n319 0.316
R2002 vp_p.n323 vp_p.n321 0.316
R2003 vp_p.n325 vp_p.n323 0.316
R2004 vp_p.n327 vp_p.n325 0.316
R2005 vp_p.n329 vp_p.n327 0.316
R2006 vp_p.n331 vp_p.n329 0.316
R2007 vp_p.n333 vp_p.n331 0.316
R2008 vp_p.n335 vp_p.n333 0.316
R2009 vp_p.n337 vp_p.n335 0.316
R2010 vp_p.n339 vp_p.n337 0.316
R2011 vp_p.n341 vp_p.n339 0.316
R2012 vp_p.n343 vp_p.n341 0.316
R2013 vp_p.n345 vp_p.n343 0.316
R2014 vp_p.n347 vp_p.n345 0.316
R2015 vp_p.n349 vp_p.n347 0.316
R2016 vp_p.n351 vp_p.n349 0.316
R2017 vp_p.n353 vp_p.n351 0.316
R2018 vp_p.n355 vp_p.n353 0.316
R2019 vp_p.n357 vp_p.n355 0.316
R2020 vp_p.n359 vp_p.n357 0.316
R2021 vp_p.n361 vp_p.n359 0.316
R2022 vp_p.n363 vp_p.n361 0.316
R2023 vp_p.n365 vp_p.n363 0.316
R2024 vp_p.n367 vp_p.n365 0.316
R2025 vp_p.n369 vp_p.n367 0.316
R2026 vp_p.n371 vp_p.n369 0.316
R2027 vp_p.n78 vp_p.n76 0.316
R2028 vp_p.n80 vp_p.n78 0.316
R2029 vp_p.n82 vp_p.n80 0.316
R2030 vp_p.n84 vp_p.n82 0.316
R2031 vp_p.n86 vp_p.n84 0.316
R2032 vp_p.n88 vp_p.n86 0.316
R2033 vp_p.n90 vp_p.n88 0.316
R2034 vp_p.n92 vp_p.n90 0.316
R2035 vp_p.n94 vp_p.n92 0.316
R2036 vp_p.n96 vp_p.n94 0.316
R2037 vp_p.n98 vp_p.n96 0.316
R2038 vp_p.n100 vp_p.n98 0.316
R2039 vp_p.n102 vp_p.n100 0.316
R2040 vp_p.n104 vp_p.n102 0.316
R2041 vp_p.n106 vp_p.n104 0.316
R2042 vp_p.n108 vp_p.n106 0.316
R2043 vp_p.n110 vp_p.n108 0.316
R2044 vp_p.n112 vp_p.n110 0.316
R2045 vp_p.n114 vp_p.n112 0.316
R2046 vp_p.n116 vp_p.n114 0.316
R2047 vp_p.n118 vp_p.n116 0.316
R2048 vp_p.n120 vp_p.n118 0.316
R2049 vp_p.n122 vp_p.n120 0.316
R2050 vp_p.n124 vp_p.n122 0.316
R2051 vp_p.n126 vp_p.n124 0.316
R2052 vp_p.n128 vp_p.n126 0.316
R2053 vp_p.n130 vp_p.n128 0.316
R2054 vp_p.n132 vp_p.n130 0.316
R2055 vp_p.n134 vp_p.n132 0.316
R2056 vp_p.n136 vp_p.n134 0.316
R2057 vp_p.n138 vp_p.n136 0.316
R2058 vp_p.n140 vp_p.n138 0.316
R2059 vp_p.n142 vp_p.n140 0.316
R2060 vp_p.n144 vp_p.n142 0.316
R2061 vp_p.n146 vp_p.n144 0.316
R2062 vp_p.n148 vp_p.n146 0.316
R2063 vp_p.n150 vp_p.n148 0.316
R2064 vp_p.n152 vp_p.n150 0.316
R2065 vp_p.n154 vp_p.n152 0.316
R2066 vp_p.n156 vp_p.n154 0.316
R2067 vp_p.n158 vp_p.n156 0.316
R2068 vp_p.n160 vp_p.n158 0.316
R2069 vp_p.n162 vp_p.n160 0.316
R2070 vp_p.n164 vp_p.n162 0.316
R2071 vp_p.n166 vp_p.n164 0.316
R2072 vp_p.n168 vp_p.n166 0.316
R2073 vp_p.n170 vp_p.n168 0.316
R2074 vp_p.n172 vp_p.n170 0.316
R2075 vp_p.n174 vp_p.n172 0.316
R2076 vp_p.n176 vp_p.n174 0.316
R2077 vp_p.n178 vp_p.n176 0.316
R2078 vp_p.n180 vp_p.n178 0.316
R2079 vp_p.n182 vp_p.n180 0.316
R2080 vp_p.n184 vp_p.n182 0.316
R2081 vp_p.n186 vp_p.n184 0.316
R2082 vp_p.n188 vp_p.n186 0.316
R2083 vp_p.n190 vp_p.n188 0.316
R2084 vp_p.n192 vp_p.n190 0.316
R2085 vp_p.n194 vp_p.n192 0.316
R2086 vp_p.n196 vp_p.n194 0.316
R2087 vp_p.n198 vp_p.n196 0.316
R2088 vp_p.n200 vp_p.n198 0.316
R2089 vp_p.n202 vp_p.n200 0.316
R2090 vp_p.n204 vp_p.n202 0.316
R2091 vp_p.n206 vp_p.n204 0.316
R2092 vp_p.n208 vp_p.n206 0.316
R2093 vp_p.n210 vp_p.n208 0.316
R2094 vp_p.n212 vp_p.n210 0.316
R2095 vp_p.n214 vp_p.n212 0.316
R2096 vp_p.n216 vp_p.n214 0.316
R2097 vp_p.n218 vp_p.n216 0.316
R2098 vp_p.n220 vp_p.n218 0.316
R2099 vp_p.n222 vp_p.n220 0.316
R2100 vp_p.n827 vp_p.n825 0.316
R2101 vp_p.n829 vp_p.n827 0.316
R2102 vp_p.n831 vp_p.n829 0.316
R2103 vp_p.n833 vp_p.n831 0.316
R2104 vp_p.n835 vp_p.n833 0.316
R2105 vp_p.n837 vp_p.n835 0.316
R2106 vp_p.n839 vp_p.n837 0.316
R2107 vp_p.n841 vp_p.n839 0.316
R2108 vp_p.n843 vp_p.n841 0.316
R2109 vp_p.n845 vp_p.n843 0.316
R2110 vp_p.n847 vp_p.n845 0.316
R2111 vp_p.n849 vp_p.n847 0.316
R2112 vp_p.n851 vp_p.n849 0.316
R2113 vp_p.n853 vp_p.n851 0.316
R2114 vp_p.n855 vp_p.n853 0.316
R2115 vp_p.n857 vp_p.n855 0.316
R2116 vp_p.n859 vp_p.n857 0.316
R2117 vp_p.n861 vp_p.n859 0.316
R2118 vp_p.n863 vp_p.n861 0.316
R2119 vp_p.n865 vp_p.n863 0.316
R2120 vp_p.n867 vp_p.n865 0.316
R2121 vp_p.n869 vp_p.n867 0.316
R2122 vp_p.n871 vp_p.n869 0.316
R2123 vp_p.n873 vp_p.n871 0.316
R2124 vp_p.n875 vp_p.n873 0.316
R2125 vp_p.n877 vp_p.n875 0.316
R2126 vp_p.n879 vp_p.n877 0.316
R2127 vp_p.n881 vp_p.n879 0.316
R2128 vp_p.n883 vp_p.n881 0.316
R2129 vp_p.n885 vp_p.n883 0.316
R2130 vp_p.n887 vp_p.n885 0.316
R2131 vp_p.n889 vp_p.n887 0.316
R2132 vp_p.n891 vp_p.n889 0.316
R2133 vp_p.n893 vp_p.n891 0.316
R2134 vp_p.n895 vp_p.n893 0.316
R2135 vp_p.n897 vp_p.n895 0.316
R2136 vp_p.n899 vp_p.n897 0.316
R2137 vp_p.n901 vp_p.n899 0.316
R2138 vp_p.n903 vp_p.n901 0.316
R2139 vp_p.n905 vp_p.n903 0.316
R2140 vp_p.n907 vp_p.n905 0.316
R2141 vp_p.n909 vp_p.n907 0.316
R2142 vp_p.n911 vp_p.n909 0.316
R2143 vp_p.n913 vp_p.n911 0.316
R2144 vp_p.n915 vp_p.n913 0.316
R2145 vp_p.n917 vp_p.n915 0.316
R2146 vp_p.n919 vp_p.n917 0.316
R2147 vp_p.n921 vp_p.n919 0.316
R2148 vp_p.n923 vp_p.n921 0.316
R2149 vp_p.n925 vp_p.n923 0.316
R2150 vp_p.n927 vp_p.n925 0.316
R2151 vp_p.n929 vp_p.n927 0.316
R2152 vp_p.n931 vp_p.n929 0.316
R2153 vp_p.n933 vp_p.n931 0.316
R2154 vp_p.n935 vp_p.n933 0.316
R2155 vp_p.n937 vp_p.n935 0.316
R2156 vp_p.n939 vp_p.n937 0.316
R2157 vp_p.n941 vp_p.n939 0.316
R2158 vp_p.n943 vp_p.n941 0.316
R2159 vp_p.n945 vp_p.n943 0.316
R2160 vp_p.n947 vp_p.n945 0.316
R2161 vp_p.n949 vp_p.n947 0.316
R2162 vp_p.n951 vp_p.n949 0.316
R2163 vp_p.n953 vp_p.n951 0.316
R2164 vp_p.n955 vp_p.n953 0.316
R2165 vp_p.n957 vp_p.n955 0.316
R2166 vp_p.n959 vp_p.n957 0.316
R2167 vp_p.n961 vp_p.n959 0.316
R2168 vp_p.n963 vp_p.n961 0.316
R2169 vp_p.n965 vp_p.n963 0.316
R2170 vp_p.n967 vp_p.n965 0.316
R2171 vp_p.n969 vp_p.n967 0.316
R2172 vp_p.n971 vp_p.n969 0.316
R2173 vp_p.n976 vp_p.n974 0.316
R2174 vp_p.n978 vp_p.n976 0.316
R2175 vp_p.n980 vp_p.n978 0.316
R2176 vp_p.n982 vp_p.n980 0.316
R2177 vp_p.n984 vp_p.n982 0.316
R2178 vp_p.n986 vp_p.n984 0.316
R2179 vp_p.n988 vp_p.n986 0.316
R2180 vp_p.n990 vp_p.n988 0.316
R2181 vp_p.n992 vp_p.n990 0.316
R2182 vp_p.n994 vp_p.n992 0.316
R2183 vp_p.n996 vp_p.n994 0.316
R2184 vp_p.n998 vp_p.n996 0.316
R2185 vp_p.n1000 vp_p.n998 0.316
R2186 vp_p.n1002 vp_p.n1000 0.316
R2187 vp_p.n1004 vp_p.n1002 0.316
R2188 vp_p.n1006 vp_p.n1004 0.316
R2189 vp_p.n1008 vp_p.n1006 0.316
R2190 vp_p.n1010 vp_p.n1008 0.316
R2191 vp_p.n1012 vp_p.n1010 0.316
R2192 vp_p.n1014 vp_p.n1012 0.316
R2193 vp_p.n1016 vp_p.n1014 0.316
R2194 vp_p.n1018 vp_p.n1016 0.316
R2195 vp_p.n1020 vp_p.n1018 0.316
R2196 vp_p.n1022 vp_p.n1020 0.316
R2197 vp_p.n1024 vp_p.n1022 0.316
R2198 vp_p.n1026 vp_p.n1024 0.316
R2199 vp_p.n1028 vp_p.n1026 0.316
R2200 vp_p.n1030 vp_p.n1028 0.316
R2201 vp_p.n1032 vp_p.n1030 0.316
R2202 vp_p.n1034 vp_p.n1032 0.316
R2203 vp_p.n1036 vp_p.n1034 0.316
R2204 vp_p.n1038 vp_p.n1036 0.316
R2205 vp_p.n1040 vp_p.n1038 0.316
R2206 vp_p.n1042 vp_p.n1040 0.316
R2207 vp_p.n1044 vp_p.n1042 0.316
R2208 vp_p.n1046 vp_p.n1044 0.316
R2209 vp_p.n1048 vp_p.n1046 0.316
R2210 vp_p.n1050 vp_p.n1048 0.316
R2211 vp_p.n1052 vp_p.n1050 0.316
R2212 vp_p.n1054 vp_p.n1052 0.316
R2213 vp_p.n1056 vp_p.n1054 0.316
R2214 vp_p.n1058 vp_p.n1056 0.316
R2215 vp_p.n1060 vp_p.n1058 0.316
R2216 vp_p.n1062 vp_p.n1060 0.316
R2217 vp_p.n1064 vp_p.n1062 0.316
R2218 vp_p.n1066 vp_p.n1064 0.316
R2219 vp_p.n1068 vp_p.n1066 0.316
R2220 vp_p.n1070 vp_p.n1068 0.316
R2221 vp_p.n1072 vp_p.n1070 0.316
R2222 vp_p.n1074 vp_p.n1072 0.316
R2223 vp_p.n1076 vp_p.n1074 0.316
R2224 vp_p.n1078 vp_p.n1076 0.316
R2225 vp_p.n1080 vp_p.n1078 0.316
R2226 vp_p.n1082 vp_p.n1080 0.316
R2227 vp_p.n1084 vp_p.n1082 0.316
R2228 vp_p.n1086 vp_p.n1084 0.316
R2229 vp_p.n1088 vp_p.n1086 0.316
R2230 vp_p.n1090 vp_p.n1088 0.316
R2231 vp_p.n1092 vp_p.n1090 0.316
R2232 vp_p.n1094 vp_p.n1092 0.316
R2233 vp_p.n1096 vp_p.n1094 0.316
R2234 vp_p.n1098 vp_p.n1096 0.316
R2235 vp_p.n1100 vp_p.n1098 0.316
R2236 vp_p.n1102 vp_p.n1100 0.316
R2237 vp_p.n1104 vp_p.n1102 0.316
R2238 vp_p.n1106 vp_p.n1104 0.316
R2239 vp_p.n1108 vp_p.n1106 0.316
R2240 vp_p.n1110 vp_p.n1108 0.316
R2241 vp_p.n1112 vp_p.n1110 0.316
R2242 vp_p.n1114 vp_p.n1112 0.316
R2243 vp_p.n1116 vp_p.n1114 0.316
R2244 vp_p.n1118 vp_p.n1116 0.316
R2245 vp_p.n1120 vp_p.n1118 0.316
R2246 vp_p.n1125 vp_p.n1123 0.316
R2247 vp_p.n1127 vp_p.n1125 0.316
R2248 vp_p.n1129 vp_p.n1127 0.316
R2249 vp_p.n1131 vp_p.n1129 0.316
R2250 vp_p.n1133 vp_p.n1131 0.316
R2251 vp_p.n1135 vp_p.n1133 0.316
R2252 vp_p.n1137 vp_p.n1135 0.316
R2253 vp_p.n1139 vp_p.n1137 0.316
R2254 vp_p.n1141 vp_p.n1139 0.316
R2255 vp_p.n1143 vp_p.n1141 0.316
R2256 vp_p.n1145 vp_p.n1143 0.316
R2257 vp_p.n1147 vp_p.n1145 0.316
R2258 vp_p.n1149 vp_p.n1147 0.316
R2259 vp_p.n1151 vp_p.n1149 0.316
R2260 vp_p.n1153 vp_p.n1151 0.316
R2261 vp_p.n1155 vp_p.n1153 0.316
R2262 vp_p.n1157 vp_p.n1155 0.316
R2263 vp_p.n1159 vp_p.n1157 0.316
R2264 vp_p.n1161 vp_p.n1159 0.316
R2265 vp_p.n1163 vp_p.n1161 0.316
R2266 vp_p.n1165 vp_p.n1163 0.316
R2267 vp_p.n1167 vp_p.n1165 0.316
R2268 vp_p.n1169 vp_p.n1167 0.316
R2269 vp_p.n1171 vp_p.n1169 0.316
R2270 vp_p.n1173 vp_p.n1171 0.316
R2271 vp_p.n1175 vp_p.n1173 0.316
R2272 vp_p.n1177 vp_p.n1175 0.316
R2273 vp_p.n1179 vp_p.n1177 0.316
R2274 vp_p.n1181 vp_p.n1179 0.316
R2275 vp_p.n1183 vp_p.n1181 0.316
R2276 vp_p.n1185 vp_p.n1183 0.316
R2277 vp_p.n1187 vp_p.n1185 0.316
R2278 vp_p.n1189 vp_p.n1187 0.316
R2279 vp_p.n1191 vp_p.n1189 0.316
R2280 vp_p.n1193 vp_p.n1191 0.316
R2281 vp_p.n1195 vp_p.n1193 0.316
R2282 vp_p.n1197 vp_p.n1195 0.316
R2283 vp_p.n1199 vp_p.n1197 0.316
R2284 vp_p.n1201 vp_p.n1199 0.316
R2285 vp_p.n1203 vp_p.n1201 0.316
R2286 vp_p.n1205 vp_p.n1203 0.316
R2287 vp_p.n1207 vp_p.n1205 0.316
R2288 vp_p.n1209 vp_p.n1207 0.316
R2289 vp_p.n1211 vp_p.n1209 0.316
R2290 vp_p.n1213 vp_p.n1211 0.316
R2291 vp_p.n1215 vp_p.n1213 0.316
R2292 vp_p.n1217 vp_p.n1215 0.316
R2293 vp_p.n1219 vp_p.n1217 0.316
R2294 vp_p.n1221 vp_p.n1219 0.316
R2295 vp_p.n1223 vp_p.n1221 0.316
R2296 vp_p.n1225 vp_p.n1223 0.316
R2297 vp_p.n1227 vp_p.n1225 0.316
R2298 vp_p.n1229 vp_p.n1227 0.316
R2299 vp_p.n1231 vp_p.n1229 0.316
R2300 vp_p.n1233 vp_p.n1231 0.316
R2301 vp_p.n1235 vp_p.n1233 0.316
R2302 vp_p.n1237 vp_p.n1235 0.316
R2303 vp_p.n1239 vp_p.n1237 0.316
R2304 vp_p.n1241 vp_p.n1239 0.316
R2305 vp_p.n1243 vp_p.n1241 0.316
R2306 vp_p.n1245 vp_p.n1243 0.316
R2307 vp_p.n1247 vp_p.n1245 0.316
R2308 vp_p.n1249 vp_p.n1247 0.316
R2309 vp_p.n1251 vp_p.n1249 0.316
R2310 vp_p.n1253 vp_p.n1251 0.316
R2311 vp_p.n1255 vp_p.n1253 0.316
R2312 vp_p.n1257 vp_p.n1255 0.316
R2313 vp_p.n1259 vp_p.n1257 0.316
R2314 vp_p.n1261 vp_p.n1259 0.316
R2315 vp_p.n1263 vp_p.n1261 0.316
R2316 vp_p.n1265 vp_p.n1263 0.316
R2317 vp_p.n1267 vp_p.n1265 0.316
R2318 vp_p.n1269 vp_p.n1267 0.316
R2319 vp_p.n1274 vp_p.n1272 0.316
R2320 vp_p.n1276 vp_p.n1274 0.316
R2321 vp_p.n1278 vp_p.n1276 0.316
R2322 vp_p.n1280 vp_p.n1278 0.316
R2323 vp_p.n1282 vp_p.n1280 0.316
R2324 vp_p.n1284 vp_p.n1282 0.316
R2325 vp_p.n1286 vp_p.n1284 0.316
R2326 vp_p.n1288 vp_p.n1286 0.316
R2327 vp_p.n1290 vp_p.n1288 0.316
R2328 vp_p.n1292 vp_p.n1290 0.316
R2329 vp_p.n1294 vp_p.n1292 0.316
R2330 vp_p.n1296 vp_p.n1294 0.316
R2331 vp_p.n1298 vp_p.n1296 0.316
R2332 vp_p.n1300 vp_p.n1298 0.316
R2333 vp_p.n1302 vp_p.n1300 0.316
R2334 vp_p.n1304 vp_p.n1302 0.316
R2335 vp_p.n1306 vp_p.n1304 0.316
R2336 vp_p.n1308 vp_p.n1306 0.316
R2337 vp_p.n1310 vp_p.n1308 0.316
R2338 vp_p.n1312 vp_p.n1310 0.316
R2339 vp_p.n1314 vp_p.n1312 0.316
R2340 vp_p.n1316 vp_p.n1314 0.316
R2341 vp_p.n1318 vp_p.n1316 0.316
R2342 vp_p.n1320 vp_p.n1318 0.316
R2343 vp_p.n1322 vp_p.n1320 0.316
R2344 vp_p.n1324 vp_p.n1322 0.316
R2345 vp_p.n1326 vp_p.n1324 0.316
R2346 vp_p.n1328 vp_p.n1326 0.316
R2347 vp_p.n1330 vp_p.n1328 0.316
R2348 vp_p.n1332 vp_p.n1330 0.316
R2349 vp_p.n1334 vp_p.n1332 0.316
R2350 vp_p.n1336 vp_p.n1334 0.316
R2351 vp_p.n1338 vp_p.n1336 0.316
R2352 vp_p.n1340 vp_p.n1338 0.316
R2353 vp_p.n1342 vp_p.n1340 0.316
R2354 vp_p.n1344 vp_p.n1342 0.316
R2355 vp_p.n1346 vp_p.n1344 0.316
R2356 vp_p.n1348 vp_p.n1346 0.316
R2357 vp_p.n1350 vp_p.n1348 0.316
R2358 vp_p.n1352 vp_p.n1350 0.316
R2359 vp_p.n1354 vp_p.n1352 0.316
R2360 vp_p.n1356 vp_p.n1354 0.316
R2361 vp_p.n1358 vp_p.n1356 0.316
R2362 vp_p.n1360 vp_p.n1358 0.316
R2363 vp_p.n1362 vp_p.n1360 0.316
R2364 vp_p.n1364 vp_p.n1362 0.316
R2365 vp_p.n1366 vp_p.n1364 0.316
R2366 vp_p.n1368 vp_p.n1366 0.316
R2367 vp_p.n1370 vp_p.n1368 0.316
R2368 vp_p.n1372 vp_p.n1370 0.316
R2369 vp_p.n1374 vp_p.n1372 0.316
R2370 vp_p.n1376 vp_p.n1374 0.316
R2371 vp_p.n1378 vp_p.n1376 0.316
R2372 vp_p.n1380 vp_p.n1378 0.316
R2373 vp_p.n1382 vp_p.n1380 0.316
R2374 vp_p.n1384 vp_p.n1382 0.316
R2375 vp_p.n1386 vp_p.n1384 0.316
R2376 vp_p.n1388 vp_p.n1386 0.316
R2377 vp_p.n1390 vp_p.n1388 0.316
R2378 vp_p.n1392 vp_p.n1390 0.316
R2379 vp_p.n1394 vp_p.n1392 0.316
R2380 vp_p.n1396 vp_p.n1394 0.316
R2381 vp_p.n1398 vp_p.n1396 0.316
R2382 vp_p.n1400 vp_p.n1398 0.316
R2383 vp_p.n1402 vp_p.n1400 0.316
R2384 vp_p.n1404 vp_p.n1402 0.316
R2385 vp_p.n1406 vp_p.n1404 0.316
R2386 vp_p.n1408 vp_p.n1406 0.316
R2387 vp_p.n1410 vp_p.n1408 0.316
R2388 vp_p.n1412 vp_p.n1410 0.316
R2389 vp_p.n1414 vp_p.n1412 0.316
R2390 vp_p.n1416 vp_p.n1414 0.316
R2391 vp_p.n1418 vp_p.n1416 0.316
R2392 vp_p.n745 vp_p.n744 0.149
R2393 vp_p.n746 vp_p.n745 0.149
R2394 vp_p.n747 vp_p.n746 0.149
R2395 vp_p.n1496 vp_p.n1495 0.149
R2396 vp_p.n1495 vp_p.n1494 0.149
R2397 vp_p.n1494 vp_p.n1493 0.149
R2398 vp_p.n748 vp_p.n747 0.141
R2399 vp_p.n1497 vp_p.n1496 0.141
R2400 vp_p.n745 vp_p.n520 0.134
R2401 vp_p.n747 vp_p.n222 0.134
R2402 vp_p.n1495 vp_p.n1120 0.134
R2403 vp_p.n1493 vp_p.n1418 0.134
R2404 vp_p.n669 vp_p.n668 0.04
R2405 vp_p.n667 vp_p.n666 0.04
R2406 vp_p.n665 vp_p.n664 0.04
R2407 vp_p.n663 vp_p.n662 0.04
R2408 vp_p.n661 vp_p.n660 0.04
R2409 vp_p.n659 vp_p.n658 0.04
R2410 vp_p.n657 vp_p.n656 0.04
R2411 vp_p.n655 vp_p.n654 0.04
R2412 vp_p.n653 vp_p.n652 0.04
R2413 vp_p.n651 vp_p.n650 0.04
R2414 vp_p.n649 vp_p.n648 0.04
R2415 vp_p.n647 vp_p.n646 0.04
R2416 vp_p.n645 vp_p.n644 0.04
R2417 vp_p.n643 vp_p.n642 0.04
R2418 vp_p.n641 vp_p.n640 0.04
R2419 vp_p.n639 vp_p.n638 0.04
R2420 vp_p.n637 vp_p.n636 0.04
R2421 vp_p.n635 vp_p.n634 0.04
R2422 vp_p.n633 vp_p.n632 0.04
R2423 vp_p.n631 vp_p.n630 0.04
R2424 vp_p.n629 vp_p.n628 0.04
R2425 vp_p.n627 vp_p.n626 0.04
R2426 vp_p.n625 vp_p.n624 0.04
R2427 vp_p.n623 vp_p.n622 0.04
R2428 vp_p.n621 vp_p.n620 0.04
R2429 vp_p.n619 vp_p.n618 0.04
R2430 vp_p.n617 vp_p.n616 0.04
R2431 vp_p.n615 vp_p.n614 0.04
R2432 vp_p.n613 vp_p.n612 0.04
R2433 vp_p.n611 vp_p.n610 0.04
R2434 vp_p.n609 vp_p.n608 0.04
R2435 vp_p.n607 vp_p.n606 0.04
R2436 vp_p.n605 vp_p.n604 0.04
R2437 vp_p.n603 vp_p.n602 0.04
R2438 vp_p.n601 vp_p.n600 0.04
R2439 vp_p.n599 vp_p.n598 0.04
R2440 vp_p.n597 vp_p.n596 0.04
R2441 vp_p.n595 vp_p.n594 0.04
R2442 vp_p.n593 vp_p.n592 0.04
R2443 vp_p.n591 vp_p.n590 0.04
R2444 vp_p.n589 vp_p.n588 0.04
R2445 vp_p.n587 vp_p.n586 0.04
R2446 vp_p.n585 vp_p.n584 0.04
R2447 vp_p.n583 vp_p.n582 0.04
R2448 vp_p.n581 vp_p.n580 0.04
R2449 vp_p.n579 vp_p.n578 0.04
R2450 vp_p.n577 vp_p.n576 0.04
R2451 vp_p.n575 vp_p.n574 0.04
R2452 vp_p.n573 vp_p.n572 0.04
R2453 vp_p.n571 vp_p.n570 0.04
R2454 vp_p.n569 vp_p.n568 0.04
R2455 vp_p.n567 vp_p.n566 0.04
R2456 vp_p.n565 vp_p.n564 0.04
R2457 vp_p.n563 vp_p.n562 0.04
R2458 vp_p.n561 vp_p.n560 0.04
R2459 vp_p.n559 vp_p.n558 0.04
R2460 vp_p.n557 vp_p.n556 0.04
R2461 vp_p.n555 vp_p.n554 0.04
R2462 vp_p.n553 vp_p.n552 0.04
R2463 vp_p.n551 vp_p.n550 0.04
R2464 vp_p.n549 vp_p.n548 0.04
R2465 vp_p.n547 vp_p.n546 0.04
R2466 vp_p.n545 vp_p.n544 0.04
R2467 vp_p.n543 vp_p.n542 0.04
R2468 vp_p.n541 vp_p.n540 0.04
R2469 vp_p.n539 vp_p.n538 0.04
R2470 vp_p.n537 vp_p.n536 0.04
R2471 vp_p.n535 vp_p.n534 0.04
R2472 vp_p.n533 vp_p.n532 0.04
R2473 vp_p.n531 vp_p.n530 0.04
R2474 vp_p.n529 vp_p.n528 0.04
R2475 vp_p.n527 vp_p.n526 0.04
R2476 vp_p.n525 vp_p.n524 0.04
R2477 vp_p.n523 vp_p.n522 0.04
R2478 vp_p.n520 vp_p.n519 0.04
R2479 vp_p.n518 vp_p.n517 0.04
R2480 vp_p.n516 vp_p.n515 0.04
R2481 vp_p.n514 vp_p.n513 0.04
R2482 vp_p.n512 vp_p.n511 0.04
R2483 vp_p.n510 vp_p.n509 0.04
R2484 vp_p.n508 vp_p.n507 0.04
R2485 vp_p.n506 vp_p.n505 0.04
R2486 vp_p.n504 vp_p.n503 0.04
R2487 vp_p.n502 vp_p.n501 0.04
R2488 vp_p.n500 vp_p.n499 0.04
R2489 vp_p.n498 vp_p.n497 0.04
R2490 vp_p.n496 vp_p.n495 0.04
R2491 vp_p.n494 vp_p.n493 0.04
R2492 vp_p.n492 vp_p.n491 0.04
R2493 vp_p.n490 vp_p.n489 0.04
R2494 vp_p.n488 vp_p.n487 0.04
R2495 vp_p.n486 vp_p.n485 0.04
R2496 vp_p.n484 vp_p.n483 0.04
R2497 vp_p.n482 vp_p.n481 0.04
R2498 vp_p.n480 vp_p.n479 0.04
R2499 vp_p.n478 vp_p.n477 0.04
R2500 vp_p.n476 vp_p.n475 0.04
R2501 vp_p.n474 vp_p.n473 0.04
R2502 vp_p.n472 vp_p.n471 0.04
R2503 vp_p.n470 vp_p.n469 0.04
R2504 vp_p.n468 vp_p.n467 0.04
R2505 vp_p.n466 vp_p.n465 0.04
R2506 vp_p.n464 vp_p.n463 0.04
R2507 vp_p.n462 vp_p.n461 0.04
R2508 vp_p.n460 vp_p.n459 0.04
R2509 vp_p.n458 vp_p.n457 0.04
R2510 vp_p.n456 vp_p.n455 0.04
R2511 vp_p.n454 vp_p.n453 0.04
R2512 vp_p.n452 vp_p.n451 0.04
R2513 vp_p.n450 vp_p.n449 0.04
R2514 vp_p.n448 vp_p.n447 0.04
R2515 vp_p.n446 vp_p.n445 0.04
R2516 vp_p.n444 vp_p.n443 0.04
R2517 vp_p.n442 vp_p.n441 0.04
R2518 vp_p.n440 vp_p.n439 0.04
R2519 vp_p.n438 vp_p.n437 0.04
R2520 vp_p.n436 vp_p.n435 0.04
R2521 vp_p.n434 vp_p.n433 0.04
R2522 vp_p.n432 vp_p.n431 0.04
R2523 vp_p.n430 vp_p.n429 0.04
R2524 vp_p.n428 vp_p.n427 0.04
R2525 vp_p.n426 vp_p.n425 0.04
R2526 vp_p.n424 vp_p.n423 0.04
R2527 vp_p.n422 vp_p.n421 0.04
R2528 vp_p.n420 vp_p.n419 0.04
R2529 vp_p.n418 vp_p.n417 0.04
R2530 vp_p.n416 vp_p.n415 0.04
R2531 vp_p.n414 vp_p.n413 0.04
R2532 vp_p.n412 vp_p.n411 0.04
R2533 vp_p.n410 vp_p.n409 0.04
R2534 vp_p.n408 vp_p.n407 0.04
R2535 vp_p.n406 vp_p.n405 0.04
R2536 vp_p.n404 vp_p.n403 0.04
R2537 vp_p.n402 vp_p.n401 0.04
R2538 vp_p.n400 vp_p.n399 0.04
R2539 vp_p.n398 vp_p.n397 0.04
R2540 vp_p.n396 vp_p.n395 0.04
R2541 vp_p.n394 vp_p.n393 0.04
R2542 vp_p.n392 vp_p.n391 0.04
R2543 vp_p.n390 vp_p.n389 0.04
R2544 vp_p.n388 vp_p.n387 0.04
R2545 vp_p.n386 vp_p.n385 0.04
R2546 vp_p.n384 vp_p.n383 0.04
R2547 vp_p.n382 vp_p.n381 0.04
R2548 vp_p.n380 vp_p.n379 0.04
R2549 vp_p.n378 vp_p.n377 0.04
R2550 vp_p.n376 vp_p.n375 0.04
R2551 vp_p.n374 vp_p.n373 0.04
R2552 vp_p.n371 vp_p.n370 0.04
R2553 vp_p.n369 vp_p.n368 0.04
R2554 vp_p.n367 vp_p.n366 0.04
R2555 vp_p.n365 vp_p.n364 0.04
R2556 vp_p.n363 vp_p.n362 0.04
R2557 vp_p.n361 vp_p.n360 0.04
R2558 vp_p.n359 vp_p.n358 0.04
R2559 vp_p.n357 vp_p.n356 0.04
R2560 vp_p.n355 vp_p.n354 0.04
R2561 vp_p.n353 vp_p.n352 0.04
R2562 vp_p.n351 vp_p.n350 0.04
R2563 vp_p.n349 vp_p.n348 0.04
R2564 vp_p.n347 vp_p.n346 0.04
R2565 vp_p.n345 vp_p.n344 0.04
R2566 vp_p.n343 vp_p.n342 0.04
R2567 vp_p.n341 vp_p.n340 0.04
R2568 vp_p.n339 vp_p.n338 0.04
R2569 vp_p.n337 vp_p.n336 0.04
R2570 vp_p.n335 vp_p.n334 0.04
R2571 vp_p.n333 vp_p.n332 0.04
R2572 vp_p.n331 vp_p.n330 0.04
R2573 vp_p.n329 vp_p.n328 0.04
R2574 vp_p.n327 vp_p.n326 0.04
R2575 vp_p.n325 vp_p.n324 0.04
R2576 vp_p.n323 vp_p.n322 0.04
R2577 vp_p.n321 vp_p.n320 0.04
R2578 vp_p.n319 vp_p.n318 0.04
R2579 vp_p.n317 vp_p.n316 0.04
R2580 vp_p.n315 vp_p.n314 0.04
R2581 vp_p.n313 vp_p.n312 0.04
R2582 vp_p.n311 vp_p.n310 0.04
R2583 vp_p.n309 vp_p.n308 0.04
R2584 vp_p.n307 vp_p.n306 0.04
R2585 vp_p.n305 vp_p.n304 0.04
R2586 vp_p.n303 vp_p.n302 0.04
R2587 vp_p.n301 vp_p.n300 0.04
R2588 vp_p.n299 vp_p.n298 0.04
R2589 vp_p.n297 vp_p.n296 0.04
R2590 vp_p.n295 vp_p.n294 0.04
R2591 vp_p.n293 vp_p.n292 0.04
R2592 vp_p.n291 vp_p.n290 0.04
R2593 vp_p.n289 vp_p.n288 0.04
R2594 vp_p.n287 vp_p.n286 0.04
R2595 vp_p.n285 vp_p.n284 0.04
R2596 vp_p.n283 vp_p.n282 0.04
R2597 vp_p.n281 vp_p.n280 0.04
R2598 vp_p.n279 vp_p.n278 0.04
R2599 vp_p.n277 vp_p.n276 0.04
R2600 vp_p.n275 vp_p.n274 0.04
R2601 vp_p.n273 vp_p.n272 0.04
R2602 vp_p.n271 vp_p.n270 0.04
R2603 vp_p.n269 vp_p.n268 0.04
R2604 vp_p.n267 vp_p.n266 0.04
R2605 vp_p.n265 vp_p.n264 0.04
R2606 vp_p.n263 vp_p.n262 0.04
R2607 vp_p.n261 vp_p.n260 0.04
R2608 vp_p.n259 vp_p.n258 0.04
R2609 vp_p.n257 vp_p.n256 0.04
R2610 vp_p.n255 vp_p.n254 0.04
R2611 vp_p.n253 vp_p.n252 0.04
R2612 vp_p.n251 vp_p.n250 0.04
R2613 vp_p.n249 vp_p.n248 0.04
R2614 vp_p.n247 vp_p.n246 0.04
R2615 vp_p.n245 vp_p.n244 0.04
R2616 vp_p.n243 vp_p.n242 0.04
R2617 vp_p.n241 vp_p.n240 0.04
R2618 vp_p.n239 vp_p.n238 0.04
R2619 vp_p.n237 vp_p.n236 0.04
R2620 vp_p.n235 vp_p.n234 0.04
R2621 vp_p.n233 vp_p.n232 0.04
R2622 vp_p.n231 vp_p.n230 0.04
R2623 vp_p.n229 vp_p.n228 0.04
R2624 vp_p.n227 vp_p.n226 0.04
R2625 vp_p.n225 vp_p.n224 0.04
R2626 vp_p.n222 vp_p.n221 0.04
R2627 vp_p.n220 vp_p.n219 0.04
R2628 vp_p.n218 vp_p.n217 0.04
R2629 vp_p.n216 vp_p.n215 0.04
R2630 vp_p.n214 vp_p.n213 0.04
R2631 vp_p.n212 vp_p.n211 0.04
R2632 vp_p.n210 vp_p.n209 0.04
R2633 vp_p.n208 vp_p.n207 0.04
R2634 vp_p.n206 vp_p.n205 0.04
R2635 vp_p.n204 vp_p.n203 0.04
R2636 vp_p.n202 vp_p.n201 0.04
R2637 vp_p.n200 vp_p.n199 0.04
R2638 vp_p.n198 vp_p.n197 0.04
R2639 vp_p.n196 vp_p.n195 0.04
R2640 vp_p.n194 vp_p.n193 0.04
R2641 vp_p.n192 vp_p.n191 0.04
R2642 vp_p.n190 vp_p.n189 0.04
R2643 vp_p.n188 vp_p.n187 0.04
R2644 vp_p.n186 vp_p.n185 0.04
R2645 vp_p.n184 vp_p.n183 0.04
R2646 vp_p.n182 vp_p.n181 0.04
R2647 vp_p.n180 vp_p.n179 0.04
R2648 vp_p.n178 vp_p.n177 0.04
R2649 vp_p.n176 vp_p.n175 0.04
R2650 vp_p.n174 vp_p.n173 0.04
R2651 vp_p.n172 vp_p.n171 0.04
R2652 vp_p.n170 vp_p.n169 0.04
R2653 vp_p.n168 vp_p.n167 0.04
R2654 vp_p.n166 vp_p.n165 0.04
R2655 vp_p.n164 vp_p.n163 0.04
R2656 vp_p.n162 vp_p.n161 0.04
R2657 vp_p.n160 vp_p.n159 0.04
R2658 vp_p.n158 vp_p.n157 0.04
R2659 vp_p.n156 vp_p.n155 0.04
R2660 vp_p.n154 vp_p.n153 0.04
R2661 vp_p.n152 vp_p.n151 0.04
R2662 vp_p.n150 vp_p.n149 0.04
R2663 vp_p.n148 vp_p.n147 0.04
R2664 vp_p.n146 vp_p.n145 0.04
R2665 vp_p.n144 vp_p.n143 0.04
R2666 vp_p.n142 vp_p.n141 0.04
R2667 vp_p.n140 vp_p.n139 0.04
R2668 vp_p.n138 vp_p.n137 0.04
R2669 vp_p.n136 vp_p.n135 0.04
R2670 vp_p.n134 vp_p.n133 0.04
R2671 vp_p.n132 vp_p.n131 0.04
R2672 vp_p.n130 vp_p.n129 0.04
R2673 vp_p.n128 vp_p.n127 0.04
R2674 vp_p.n126 vp_p.n125 0.04
R2675 vp_p.n124 vp_p.n123 0.04
R2676 vp_p.n122 vp_p.n121 0.04
R2677 vp_p.n120 vp_p.n119 0.04
R2678 vp_p.n118 vp_p.n117 0.04
R2679 vp_p.n116 vp_p.n115 0.04
R2680 vp_p.n114 vp_p.n113 0.04
R2681 vp_p.n112 vp_p.n111 0.04
R2682 vp_p.n110 vp_p.n109 0.04
R2683 vp_p.n108 vp_p.n107 0.04
R2684 vp_p.n106 vp_p.n105 0.04
R2685 vp_p.n104 vp_p.n103 0.04
R2686 vp_p.n102 vp_p.n101 0.04
R2687 vp_p.n100 vp_p.n99 0.04
R2688 vp_p.n98 vp_p.n97 0.04
R2689 vp_p.n96 vp_p.n95 0.04
R2690 vp_p.n94 vp_p.n93 0.04
R2691 vp_p.n92 vp_p.n91 0.04
R2692 vp_p.n90 vp_p.n89 0.04
R2693 vp_p.n88 vp_p.n87 0.04
R2694 vp_p.n86 vp_p.n85 0.04
R2695 vp_p.n84 vp_p.n83 0.04
R2696 vp_p.n82 vp_p.n81 0.04
R2697 vp_p.n80 vp_p.n79 0.04
R2698 vp_p.n78 vp_p.n77 0.04
R2699 vp_p.n76 vp_p.n75 0.04
R2700 vp_p.n971 vp_p.n970 0.04
R2701 vp_p.n969 vp_p.n968 0.04
R2702 vp_p.n967 vp_p.n966 0.04
R2703 vp_p.n965 vp_p.n964 0.04
R2704 vp_p.n963 vp_p.n962 0.04
R2705 vp_p.n961 vp_p.n960 0.04
R2706 vp_p.n959 vp_p.n958 0.04
R2707 vp_p.n957 vp_p.n956 0.04
R2708 vp_p.n955 vp_p.n954 0.04
R2709 vp_p.n953 vp_p.n952 0.04
R2710 vp_p.n951 vp_p.n950 0.04
R2711 vp_p.n949 vp_p.n948 0.04
R2712 vp_p.n947 vp_p.n946 0.04
R2713 vp_p.n945 vp_p.n944 0.04
R2714 vp_p.n943 vp_p.n942 0.04
R2715 vp_p.n941 vp_p.n940 0.04
R2716 vp_p.n939 vp_p.n938 0.04
R2717 vp_p.n937 vp_p.n936 0.04
R2718 vp_p.n935 vp_p.n934 0.04
R2719 vp_p.n933 vp_p.n932 0.04
R2720 vp_p.n931 vp_p.n930 0.04
R2721 vp_p.n929 vp_p.n928 0.04
R2722 vp_p.n927 vp_p.n926 0.04
R2723 vp_p.n925 vp_p.n924 0.04
R2724 vp_p.n923 vp_p.n922 0.04
R2725 vp_p.n921 vp_p.n920 0.04
R2726 vp_p.n919 vp_p.n918 0.04
R2727 vp_p.n917 vp_p.n916 0.04
R2728 vp_p.n915 vp_p.n914 0.04
R2729 vp_p.n913 vp_p.n912 0.04
R2730 vp_p.n911 vp_p.n910 0.04
R2731 vp_p.n909 vp_p.n908 0.04
R2732 vp_p.n907 vp_p.n906 0.04
R2733 vp_p.n905 vp_p.n904 0.04
R2734 vp_p.n903 vp_p.n902 0.04
R2735 vp_p.n901 vp_p.n900 0.04
R2736 vp_p.n899 vp_p.n898 0.04
R2737 vp_p.n897 vp_p.n896 0.04
R2738 vp_p.n895 vp_p.n894 0.04
R2739 vp_p.n893 vp_p.n892 0.04
R2740 vp_p.n891 vp_p.n890 0.04
R2741 vp_p.n889 vp_p.n888 0.04
R2742 vp_p.n887 vp_p.n886 0.04
R2743 vp_p.n885 vp_p.n884 0.04
R2744 vp_p.n883 vp_p.n882 0.04
R2745 vp_p.n881 vp_p.n880 0.04
R2746 vp_p.n879 vp_p.n878 0.04
R2747 vp_p.n877 vp_p.n876 0.04
R2748 vp_p.n875 vp_p.n874 0.04
R2749 vp_p.n873 vp_p.n872 0.04
R2750 vp_p.n871 vp_p.n870 0.04
R2751 vp_p.n869 vp_p.n868 0.04
R2752 vp_p.n867 vp_p.n866 0.04
R2753 vp_p.n865 vp_p.n864 0.04
R2754 vp_p.n863 vp_p.n862 0.04
R2755 vp_p.n861 vp_p.n860 0.04
R2756 vp_p.n859 vp_p.n858 0.04
R2757 vp_p.n857 vp_p.n856 0.04
R2758 vp_p.n855 vp_p.n854 0.04
R2759 vp_p.n853 vp_p.n852 0.04
R2760 vp_p.n851 vp_p.n850 0.04
R2761 vp_p.n849 vp_p.n848 0.04
R2762 vp_p.n847 vp_p.n846 0.04
R2763 vp_p.n845 vp_p.n844 0.04
R2764 vp_p.n843 vp_p.n842 0.04
R2765 vp_p.n841 vp_p.n840 0.04
R2766 vp_p.n839 vp_p.n838 0.04
R2767 vp_p.n837 vp_p.n836 0.04
R2768 vp_p.n835 vp_p.n834 0.04
R2769 vp_p.n833 vp_p.n832 0.04
R2770 vp_p.n831 vp_p.n830 0.04
R2771 vp_p.n829 vp_p.n828 0.04
R2772 vp_p.n827 vp_p.n826 0.04
R2773 vp_p.n825 vp_p.n824 0.04
R2774 vp_p.n1120 vp_p.n1119 0.04
R2775 vp_p.n1118 vp_p.n1117 0.04
R2776 vp_p.n1116 vp_p.n1115 0.04
R2777 vp_p.n1114 vp_p.n1113 0.04
R2778 vp_p.n1112 vp_p.n1111 0.04
R2779 vp_p.n1110 vp_p.n1109 0.04
R2780 vp_p.n1108 vp_p.n1107 0.04
R2781 vp_p.n1106 vp_p.n1105 0.04
R2782 vp_p.n1104 vp_p.n1103 0.04
R2783 vp_p.n1102 vp_p.n1101 0.04
R2784 vp_p.n1100 vp_p.n1099 0.04
R2785 vp_p.n1098 vp_p.n1097 0.04
R2786 vp_p.n1096 vp_p.n1095 0.04
R2787 vp_p.n1094 vp_p.n1093 0.04
R2788 vp_p.n1092 vp_p.n1091 0.04
R2789 vp_p.n1090 vp_p.n1089 0.04
R2790 vp_p.n1088 vp_p.n1087 0.04
R2791 vp_p.n1086 vp_p.n1085 0.04
R2792 vp_p.n1084 vp_p.n1083 0.04
R2793 vp_p.n1082 vp_p.n1081 0.04
R2794 vp_p.n1080 vp_p.n1079 0.04
R2795 vp_p.n1078 vp_p.n1077 0.04
R2796 vp_p.n1076 vp_p.n1075 0.04
R2797 vp_p.n1074 vp_p.n1073 0.04
R2798 vp_p.n1072 vp_p.n1071 0.04
R2799 vp_p.n1070 vp_p.n1069 0.04
R2800 vp_p.n1068 vp_p.n1067 0.04
R2801 vp_p.n1066 vp_p.n1065 0.04
R2802 vp_p.n1064 vp_p.n1063 0.04
R2803 vp_p.n1062 vp_p.n1061 0.04
R2804 vp_p.n1060 vp_p.n1059 0.04
R2805 vp_p.n1058 vp_p.n1057 0.04
R2806 vp_p.n1056 vp_p.n1055 0.04
R2807 vp_p.n1054 vp_p.n1053 0.04
R2808 vp_p.n1052 vp_p.n1051 0.04
R2809 vp_p.n1050 vp_p.n1049 0.04
R2810 vp_p.n1048 vp_p.n1047 0.04
R2811 vp_p.n1046 vp_p.n1045 0.04
R2812 vp_p.n1044 vp_p.n1043 0.04
R2813 vp_p.n1042 vp_p.n1041 0.04
R2814 vp_p.n1040 vp_p.n1039 0.04
R2815 vp_p.n1038 vp_p.n1037 0.04
R2816 vp_p.n1036 vp_p.n1035 0.04
R2817 vp_p.n1034 vp_p.n1033 0.04
R2818 vp_p.n1032 vp_p.n1031 0.04
R2819 vp_p.n1030 vp_p.n1029 0.04
R2820 vp_p.n1028 vp_p.n1027 0.04
R2821 vp_p.n1026 vp_p.n1025 0.04
R2822 vp_p.n1024 vp_p.n1023 0.04
R2823 vp_p.n1022 vp_p.n1021 0.04
R2824 vp_p.n1020 vp_p.n1019 0.04
R2825 vp_p.n1018 vp_p.n1017 0.04
R2826 vp_p.n1016 vp_p.n1015 0.04
R2827 vp_p.n1014 vp_p.n1013 0.04
R2828 vp_p.n1012 vp_p.n1011 0.04
R2829 vp_p.n1010 vp_p.n1009 0.04
R2830 vp_p.n1008 vp_p.n1007 0.04
R2831 vp_p.n1006 vp_p.n1005 0.04
R2832 vp_p.n1004 vp_p.n1003 0.04
R2833 vp_p.n1002 vp_p.n1001 0.04
R2834 vp_p.n1000 vp_p.n999 0.04
R2835 vp_p.n998 vp_p.n997 0.04
R2836 vp_p.n996 vp_p.n995 0.04
R2837 vp_p.n994 vp_p.n993 0.04
R2838 vp_p.n992 vp_p.n991 0.04
R2839 vp_p.n990 vp_p.n989 0.04
R2840 vp_p.n988 vp_p.n987 0.04
R2841 vp_p.n986 vp_p.n985 0.04
R2842 vp_p.n984 vp_p.n983 0.04
R2843 vp_p.n982 vp_p.n981 0.04
R2844 vp_p.n980 vp_p.n979 0.04
R2845 vp_p.n978 vp_p.n977 0.04
R2846 vp_p.n976 vp_p.n975 0.04
R2847 vp_p.n974 vp_p.n973 0.04
R2848 vp_p.n1269 vp_p.n1268 0.04
R2849 vp_p.n1267 vp_p.n1266 0.04
R2850 vp_p.n1265 vp_p.n1264 0.04
R2851 vp_p.n1263 vp_p.n1262 0.04
R2852 vp_p.n1261 vp_p.n1260 0.04
R2853 vp_p.n1259 vp_p.n1258 0.04
R2854 vp_p.n1257 vp_p.n1256 0.04
R2855 vp_p.n1255 vp_p.n1254 0.04
R2856 vp_p.n1253 vp_p.n1252 0.04
R2857 vp_p.n1251 vp_p.n1250 0.04
R2858 vp_p.n1249 vp_p.n1248 0.04
R2859 vp_p.n1247 vp_p.n1246 0.04
R2860 vp_p.n1245 vp_p.n1244 0.04
R2861 vp_p.n1243 vp_p.n1242 0.04
R2862 vp_p.n1241 vp_p.n1240 0.04
R2863 vp_p.n1239 vp_p.n1238 0.04
R2864 vp_p.n1237 vp_p.n1236 0.04
R2865 vp_p.n1235 vp_p.n1234 0.04
R2866 vp_p.n1233 vp_p.n1232 0.04
R2867 vp_p.n1231 vp_p.n1230 0.04
R2868 vp_p.n1229 vp_p.n1228 0.04
R2869 vp_p.n1227 vp_p.n1226 0.04
R2870 vp_p.n1225 vp_p.n1224 0.04
R2871 vp_p.n1223 vp_p.n1222 0.04
R2872 vp_p.n1221 vp_p.n1220 0.04
R2873 vp_p.n1219 vp_p.n1218 0.04
R2874 vp_p.n1217 vp_p.n1216 0.04
R2875 vp_p.n1215 vp_p.n1214 0.04
R2876 vp_p.n1213 vp_p.n1212 0.04
R2877 vp_p.n1211 vp_p.n1210 0.04
R2878 vp_p.n1209 vp_p.n1208 0.04
R2879 vp_p.n1207 vp_p.n1206 0.04
R2880 vp_p.n1205 vp_p.n1204 0.04
R2881 vp_p.n1203 vp_p.n1202 0.04
R2882 vp_p.n1201 vp_p.n1200 0.04
R2883 vp_p.n1199 vp_p.n1198 0.04
R2884 vp_p.n1197 vp_p.n1196 0.04
R2885 vp_p.n1195 vp_p.n1194 0.04
R2886 vp_p.n1193 vp_p.n1192 0.04
R2887 vp_p.n1191 vp_p.n1190 0.04
R2888 vp_p.n1189 vp_p.n1188 0.04
R2889 vp_p.n1187 vp_p.n1186 0.04
R2890 vp_p.n1185 vp_p.n1184 0.04
R2891 vp_p.n1183 vp_p.n1182 0.04
R2892 vp_p.n1181 vp_p.n1180 0.04
R2893 vp_p.n1179 vp_p.n1178 0.04
R2894 vp_p.n1177 vp_p.n1176 0.04
R2895 vp_p.n1175 vp_p.n1174 0.04
R2896 vp_p.n1173 vp_p.n1172 0.04
R2897 vp_p.n1171 vp_p.n1170 0.04
R2898 vp_p.n1169 vp_p.n1168 0.04
R2899 vp_p.n1167 vp_p.n1166 0.04
R2900 vp_p.n1165 vp_p.n1164 0.04
R2901 vp_p.n1163 vp_p.n1162 0.04
R2902 vp_p.n1161 vp_p.n1160 0.04
R2903 vp_p.n1159 vp_p.n1158 0.04
R2904 vp_p.n1157 vp_p.n1156 0.04
R2905 vp_p.n1155 vp_p.n1154 0.04
R2906 vp_p.n1153 vp_p.n1152 0.04
R2907 vp_p.n1151 vp_p.n1150 0.04
R2908 vp_p.n1149 vp_p.n1148 0.04
R2909 vp_p.n1147 vp_p.n1146 0.04
R2910 vp_p.n1145 vp_p.n1144 0.04
R2911 vp_p.n1143 vp_p.n1142 0.04
R2912 vp_p.n1141 vp_p.n1140 0.04
R2913 vp_p.n1139 vp_p.n1138 0.04
R2914 vp_p.n1137 vp_p.n1136 0.04
R2915 vp_p.n1135 vp_p.n1134 0.04
R2916 vp_p.n1133 vp_p.n1132 0.04
R2917 vp_p.n1131 vp_p.n1130 0.04
R2918 vp_p.n1129 vp_p.n1128 0.04
R2919 vp_p.n1127 vp_p.n1126 0.04
R2920 vp_p.n1125 vp_p.n1124 0.04
R2921 vp_p.n1123 vp_p.n1122 0.04
R2922 vp_p.n1418 vp_p.n1417 0.04
R2923 vp_p.n1416 vp_p.n1415 0.04
R2924 vp_p.n1414 vp_p.n1413 0.04
R2925 vp_p.n1412 vp_p.n1411 0.04
R2926 vp_p.n1410 vp_p.n1409 0.04
R2927 vp_p.n1408 vp_p.n1407 0.04
R2928 vp_p.n1406 vp_p.n1405 0.04
R2929 vp_p.n1404 vp_p.n1403 0.04
R2930 vp_p.n1402 vp_p.n1401 0.04
R2931 vp_p.n1400 vp_p.n1399 0.04
R2932 vp_p.n1398 vp_p.n1397 0.04
R2933 vp_p.n1396 vp_p.n1395 0.04
R2934 vp_p.n1394 vp_p.n1393 0.04
R2935 vp_p.n1392 vp_p.n1391 0.04
R2936 vp_p.n1390 vp_p.n1389 0.04
R2937 vp_p.n1388 vp_p.n1387 0.04
R2938 vp_p.n1386 vp_p.n1385 0.04
R2939 vp_p.n1384 vp_p.n1383 0.04
R2940 vp_p.n1382 vp_p.n1381 0.04
R2941 vp_p.n1380 vp_p.n1379 0.04
R2942 vp_p.n1378 vp_p.n1377 0.04
R2943 vp_p.n1376 vp_p.n1375 0.04
R2944 vp_p.n1374 vp_p.n1373 0.04
R2945 vp_p.n1372 vp_p.n1371 0.04
R2946 vp_p.n1370 vp_p.n1369 0.04
R2947 vp_p.n1368 vp_p.n1367 0.04
R2948 vp_p.n1366 vp_p.n1365 0.04
R2949 vp_p.n1364 vp_p.n1363 0.04
R2950 vp_p.n1362 vp_p.n1361 0.04
R2951 vp_p.n1360 vp_p.n1359 0.04
R2952 vp_p.n1358 vp_p.n1357 0.04
R2953 vp_p.n1356 vp_p.n1355 0.04
R2954 vp_p.n1354 vp_p.n1353 0.04
R2955 vp_p.n1352 vp_p.n1351 0.04
R2956 vp_p.n1350 vp_p.n1349 0.04
R2957 vp_p.n1348 vp_p.n1347 0.04
R2958 vp_p.n1346 vp_p.n1345 0.04
R2959 vp_p.n1344 vp_p.n1343 0.04
R2960 vp_p.n1342 vp_p.n1341 0.04
R2961 vp_p.n1340 vp_p.n1339 0.04
R2962 vp_p.n1338 vp_p.n1337 0.04
R2963 vp_p.n1336 vp_p.n1335 0.04
R2964 vp_p.n1334 vp_p.n1333 0.04
R2965 vp_p.n1332 vp_p.n1331 0.04
R2966 vp_p.n1330 vp_p.n1329 0.04
R2967 vp_p.n1328 vp_p.n1327 0.04
R2968 vp_p.n1326 vp_p.n1325 0.04
R2969 vp_p.n1324 vp_p.n1323 0.04
R2970 vp_p.n1322 vp_p.n1321 0.04
R2971 vp_p.n1320 vp_p.n1319 0.04
R2972 vp_p.n1318 vp_p.n1317 0.04
R2973 vp_p.n1316 vp_p.n1315 0.04
R2974 vp_p.n1314 vp_p.n1313 0.04
R2975 vp_p.n1312 vp_p.n1311 0.04
R2976 vp_p.n1310 vp_p.n1309 0.04
R2977 vp_p.n1308 vp_p.n1307 0.04
R2978 vp_p.n1306 vp_p.n1305 0.04
R2979 vp_p.n1304 vp_p.n1303 0.04
R2980 vp_p.n1302 vp_p.n1301 0.04
R2981 vp_p.n1300 vp_p.n1299 0.04
R2982 vp_p.n1298 vp_p.n1297 0.04
R2983 vp_p.n1296 vp_p.n1295 0.04
R2984 vp_p.n1294 vp_p.n1293 0.04
R2985 vp_p.n1292 vp_p.n1291 0.04
R2986 vp_p.n1290 vp_p.n1289 0.04
R2987 vp_p.n1288 vp_p.n1287 0.04
R2988 vp_p.n1286 vp_p.n1285 0.04
R2989 vp_p.n1284 vp_p.n1283 0.04
R2990 vp_p.n1282 vp_p.n1281 0.04
R2991 vp_p.n1280 vp_p.n1279 0.04
R2992 vp_p.n1278 vp_p.n1277 0.04
R2993 vp_p.n1276 vp_p.n1275 0.04
R2994 vp_p.n1274 vp_p.n1273 0.04
R2995 vp_p.n1272 vp_p.n1271 0.04
R2996 vp_p vp_p.n748 0.028
R2997 vp_p vp_p.n1497 0.005
R2998 out_p.n36 out_p.t782 8.126
R2999 out_p.n36 out_p.t1149 8.126
R3000 out_p.n37 out_p.t1137 8.126
R3001 out_p.n37 out_p.t779 8.126
R3002 out_p.n38 out_p.t319 8.126
R3003 out_p.n38 out_p.t1199 8.126
R3004 out_p.n39 out_p.t605 8.126
R3005 out_p.n39 out_p.t533 8.126
R3006 out_p.n40 out_p.t701 8.126
R3007 out_p.n40 out_p.t389 8.126
R3008 out_p.n41 out_p.t1385 8.126
R3009 out_p.n41 out_p.t1165 8.126
R3010 out_p.n42 out_p.t629 8.126
R3011 out_p.n42 out_p.t1010 8.126
R3012 out_p.n43 out_p.t1100 8.126
R3013 out_p.n43 out_p.t942 8.126
R3014 out_p.n44 out_p.t1259 8.126
R3015 out_p.n44 out_p.t283 8.126
R3016 out_p.n45 out_p.t824 8.126
R3017 out_p.n45 out_p.t845 8.126
R3018 out_p.n47 out_p.t968 8.126
R3019 out_p.n47 out_p.t733 8.126
R3020 out_p.n48 out_p.t443 8.126
R3021 out_p.n48 out_p.t1416 8.126
R3022 out_p.n49 out_p.t465 8.126
R3023 out_p.n49 out_p.t1361 8.126
R3024 out_p.n50 out_p.t244 8.126
R3025 out_p.n50 out_p.t1460 8.126
R3026 out_p.n51 out_p.t522 8.126
R3027 out_p.n51 out_p.t986 8.126
R3028 out_p.n52 out_p.t991 8.126
R3029 out_p.n52 out_p.t1340 8.126
R3030 out_p.n53 out_p.t1318 8.126
R3031 out_p.n53 out_p.t1529 8.126
R3032 out_p.n54 out_p.t492 8.126
R3033 out_p.n54 out_p.t1542 8.126
R3034 out_p.n55 out_p.t520 8.126
R3035 out_p.n55 out_p.t868 8.126
R3036 out_p.n56 out_p.t704 8.126
R3037 out_p.n56 out_p.t761 8.126
R3038 out_p.n58 out_p.t1527 8.126
R3039 out_p.n58 out_p.t450 8.126
R3040 out_p.n59 out_p.t551 8.126
R3041 out_p.n59 out_p.t1218 8.126
R3042 out_p.n60 out_p.t1140 8.126
R3043 out_p.n60 out_p.t890 8.126
R3044 out_p.n61 out_p.t1345 8.126
R3045 out_p.n61 out_p.t327 8.126
R3046 out_p.n62 out_p.t651 8.126
R3047 out_p.n62 out_p.t1574 8.126
R3048 out_p.n63 out_p.t705 8.126
R3049 out_p.n63 out_p.t421 8.126
R3050 out_p.n64 out_p.t1244 8.126
R3051 out_p.n64 out_p.t1353 8.126
R3052 out_p.n65 out_p.t919 8.126
R3053 out_p.n65 out_p.t817 8.126
R3054 out_p.n66 out_p.t1150 8.126
R3055 out_p.n66 out_p.t1001 8.126
R3056 out_p.n67 out_p.t176 8.126
R3057 out_p.n67 out_p.t1500 8.126
R3058 out_p.n69 out_p.t1372 8.126
R3059 out_p.n69 out_p.t1003 8.126
R3060 out_p.n70 out_p.t1296 8.126
R3061 out_p.n70 out_p.t896 8.126
R3062 out_p.n71 out_p.t980 8.126
R3063 out_p.n71 out_p.t1091 8.126
R3064 out_p.n72 out_p.t935 8.126
R3065 out_p.n72 out_p.t653 8.126
R3066 out_p.n73 out_p.t1588 8.126
R3067 out_p.n73 out_p.t807 8.126
R3068 out_p.n74 out_p.t1334 8.126
R3069 out_p.n74 out_p.t308 8.126
R3070 out_p.n75 out_p.t599 8.126
R3071 out_p.n75 out_p.t1130 8.126
R3072 out_p.n76 out_p.t293 8.126
R3073 out_p.n76 out_p.t243 8.126
R3074 out_p.n77 out_p.t1123 8.126
R3075 out_p.n77 out_p.t1116 8.126
R3076 out_p.n78 out_p.t1587 8.126
R3077 out_p.n78 out_p.t1034 8.126
R3078 out_p.n80 out_p.t458 8.126
R3079 out_p.n80 out_p.t1337 8.126
R3080 out_p.n81 out_p.t330 8.126
R3081 out_p.n81 out_p.t1329 8.126
R3082 out_p.n82 out_p.t436 8.126
R3083 out_p.n82 out_p.t904 8.126
R3084 out_p.n83 out_p.t1154 8.126
R3085 out_p.n83 out_p.t659 8.126
R3086 out_p.n84 out_p.t1585 8.126
R3087 out_p.n84 out_p.t1545 8.126
R3088 out_p.n85 out_p.t1070 8.126
R3089 out_p.n85 out_p.t830 8.126
R3090 out_p.n86 out_p.t597 8.126
R3091 out_p.n86 out_p.t954 8.126
R3092 out_p.n87 out_p.t1546 8.126
R3093 out_p.n87 out_p.t1124 8.126
R3094 out_p.n88 out_p.t1613 8.126
R3095 out_p.n88 out_p.t1279 8.126
R3096 out_p.n89 out_p.t1592 8.126
R3097 out_p.n89 out_p.t1009 8.126
R3098 out_p.n91 out_p.t998 8.126
R3099 out_p.n91 out_p.t497 8.126
R3100 out_p.n92 out_p.t768 8.126
R3101 out_p.n92 out_p.t380 8.126
R3102 out_p.n93 out_p.t1235 8.126
R3103 out_p.n93 out_p.t1465 8.126
R3104 out_p.n94 out_p.t547 8.126
R3105 out_p.n94 out_p.t920 8.126
R3106 out_p.n95 out_p.t863 8.126
R3107 out_p.n95 out_p.t1507 8.126
R3108 out_p.n96 out_p.t1277 8.126
R3109 out_p.n96 out_p.t262 8.126
R3110 out_p.n97 out_p.t1430 8.126
R3111 out_p.n97 out_p.t1012 8.126
R3112 out_p.n98 out_p.t215 8.126
R3113 out_p.n98 out_p.t1048 8.126
R3114 out_p.n99 out_p.t592 8.126
R3115 out_p.n99 out_p.t1616 8.126
R3116 out_p.n100 out_p.t810 8.126
R3117 out_p.n100 out_p.t1126 8.126
R3118 out_p.n102 out_p.t1166 8.126
R3119 out_p.n102 out_p.t1348 8.126
R3120 out_p.n103 out_p.t212 8.126
R3121 out_p.n103 out_p.t1171 8.126
R3122 out_p.n104 out_p.t693 8.126
R3123 out_p.n104 out_p.t1560 8.126
R3124 out_p.n105 out_p.t1408 8.126
R3125 out_p.n105 out_p.t799 8.126
R3126 out_p.n106 out_p.t1608 8.126
R3127 out_p.n106 out_p.t1386 8.126
R3128 out_p.n107 out_p.t1142 8.126
R3129 out_p.n107 out_p.t364 8.126
R3130 out_p.n108 out_p.t1499 8.126
R3131 out_p.n108 out_p.t706 8.126
R3132 out_p.n109 out_p.t532 8.126
R3133 out_p.n109 out_p.t1194 8.126
R3134 out_p.n110 out_p.t388 8.126
R3135 out_p.n110 out_p.t1234 8.126
R3136 out_p.n111 out_p.t260 8.126
R3137 out_p.n111 out_p.t232 8.126
R3138 out_p.n113 out_p.t639 8.126
R3139 out_p.n113 out_p.t316 8.126
R3140 out_p.n114 out_p.t485 8.126
R3141 out_p.n114 out_p.t1251 8.126
R3142 out_p.n115 out_p.t717 8.126
R3143 out_p.n115 out_p.t1065 8.126
R3144 out_p.n116 out_p.t1027 8.126
R3145 out_p.n116 out_p.t747 8.126
R3146 out_p.n117 out_p.t732 8.126
R3147 out_p.n117 out_p.t758 8.126
R3148 out_p.n118 out_p.t1572 8.126
R3149 out_p.n118 out_p.t1413 8.126
R3150 out_p.n119 out_p.t413 8.126
R3151 out_p.n119 out_p.t1356 8.126
R3152 out_p.n120 out_p.t580 8.126
R3153 out_p.n120 out_p.t604 8.126
R3154 out_p.n121 out_p.t1164 8.126
R3155 out_p.n121 out_p.t700 8.126
R3156 out_p.n122 out_p.t1509 8.126
R3157 out_p.n122 out_p.t219 8.126
R3158 out_p.n124 out_p.t1482 8.126
R3159 out_p.n124 out_p.t416 8.126
R3160 out_p.n125 out_p.t1475 8.126
R3161 out_p.n125 out_p.t979 8.126
R3162 out_p.n126 out_p.t448 8.126
R3163 out_p.n126 out_p.t1575 8.126
R3164 out_p.n127 out_p.t1275 8.126
R3165 out_p.n127 out_p.t895 8.126
R3166 out_p.n128 out_p.t203 8.126
R3167 out_p.n128 out_p.t1290 8.126
R3168 out_p.n129 out_p.t469 8.126
R3169 out_p.n129 out_p.t1113 8.126
R3170 out_p.n130 out_p.t1307 8.126
R3171 out_p.n130 out_p.t494 8.126
R3172 out_p.n131 out_p.t1204 8.126
R3173 out_p.n131 out_p.t803 8.126
R3174 out_p.n132 out_p.t1472 8.126
R3175 out_p.n132 out_p.t1346 8.126
R3176 out_p.n133 out_p.t473 8.126
R3177 out_p.n133 out_p.t264 8.126
R3178 out_p.n135 out_p.t1053 8.126
R3179 out_p.n135 out_p.t162 8.126
R3180 out_p.n136 out_p.t1224 8.126
R3181 out_p.n136 out_p.t1223 8.126
R3182 out_p.n137 out_p.t903 8.126
R3183 out_p.n137 out_p.t1324 8.126
R3184 out_p.n138 out_p.t315 8.126
R3185 out_p.n138 out_p.t729 8.126
R3186 out_p.n139 out_p.t406 8.126
R3187 out_p.n139 out_p.t555 8.126
R3188 out_p.n140 out_p.t274 8.126
R3189 out_p.n140 out_p.t265 8.126
R3190 out_p.n141 out_p.t387 8.126
R3191 out_p.n141 out_p.t512 8.126
R3192 out_p.n142 out_p.t985 8.126
R3193 out_p.n142 out_p.t410 8.126
R3194 out_p.n143 out_p.t420 8.126
R3195 out_p.n143 out_p.t337 8.126
R3196 out_p.n144 out_p.t1549 8.126
R3197 out_p.n144 out_p.t767 8.126
R3198 out_p.n146 out_p.t240 8.126
R3199 out_p.n146 out_p.t570 8.126
R3200 out_p.n147 out_p.t1104 8.126
R3201 out_p.n147 out_p.t694 8.126
R3202 out_p.n148 out_p.t1519 8.126
R3203 out_p.n148 out_p.t905 8.126
R3204 out_p.n149 out_p.t850 8.126
R3205 out_p.n149 out_p.t276 8.126
R3206 out_p.n150 out_p.t1383 8.126
R3207 out_p.n150 out_p.t418 8.126
R3208 out_p.n151 out_p.t1525 8.126
R3209 out_p.n151 out_p.t1453 8.126
R3210 out_p.n152 out_p.t179 8.126
R3211 out_p.n152 out_p.t955 8.126
R3212 out_p.n153 out_p.t1481 8.126
R3213 out_p.n153 out_p.t587 8.126
R3214 out_p.n154 out_p.t1088 8.126
R3215 out_p.n154 out_p.t1278 8.126
R3216 out_p.n155 out_p.t247 8.126
R3217 out_p.n155 out_p.t1008 8.126
R3218 out_p.n157 out_p.t376 8.126
R3219 out_p.n157 out_p.t1562 8.126
R3220 out_p.n158 out_p.t959 8.126
R3221 out_p.n158 out_p.t765 8.126
R3222 out_p.n159 out_p.t886 8.126
R3223 out_p.n159 out_p.t300 8.126
R3224 out_p.n160 out_p.t1261 8.126
R3225 out_p.n160 out_p.t1114 8.126
R3226 out_p.n161 out_p.t675 8.126
R3227 out_p.n161 out_p.t363 8.126
R3228 out_p.n162 out_p.t1208 8.126
R3229 out_p.n162 out_p.t1228 8.126
R3230 out_p.n163 out_p.t440 8.126
R3231 out_p.n163 out_p.t1331 8.126
R3232 out_p.n164 out_p.t1492 8.126
R3233 out_p.n164 out_p.t852 8.126
R3234 out_p.n165 out_p.t225 8.126
R3235 out_p.n165 out_p.t618 8.126
R3236 out_p.n166 out_p.t197 8.126
R3237 out_p.n166 out_p.t735 8.126
R3238 out_p.n168 out_p.t1308 8.126
R3239 out_p.n168 out_p.t1622 8.126
R3240 out_p.n169 out_p.t460 8.126
R3241 out_p.n169 out_p.t1397 8.126
R3242 out_p.n170 out_p.t166 8.126
R3243 out_p.n170 out_p.t1045 8.126
R3244 out_p.n171 out_p.t1571 8.126
R3245 out_p.n171 out_p.t1459 8.126
R3246 out_p.n172 out_p.t718 8.126
R3247 out_p.n172 out_p.t922 8.126
R3248 out_p.n173 out_p.t698 8.126
R3249 out_p.n173 out_p.t384 8.126
R3250 out_p.n174 out_p.t1395 8.126
R3251 out_p.n174 out_p.t1619 8.126
R3252 out_p.n175 out_p.t1655 8.126
R3253 out_p.n175 out_p.t916 8.126
R3254 out_p.n176 out_p.t1489 8.126
R3255 out_p.n176 out_p.t352 8.126
R3256 out_p.n177 out_p.t1060 8.126
R3257 out_p.n177 out_p.t296 8.126
R3258 out_p.n0 out_p.t871 8.126
R3259 out_p.n0 out_p.t1295 8.126
R3260 out_p.n1 out_p.t593 8.126
R3261 out_p.n1 out_p.t360 8.126
R3262 out_p.n2 out_p.t1424 8.126
R3263 out_p.n2 out_p.t759 8.126
R3264 out_p.n3 out_p.t180 8.126
R3265 out_p.n3 out_p.t882 8.126
R3266 out_p.n4 out_p.t771 8.126
R3267 out_p.n4 out_p.t516 8.126
R3268 out_p.n5 out_p.t187 8.126
R3269 out_p.n5 out_p.t785 8.126
R3270 out_p.n6 out_p.t648 8.126
R3271 out_p.n6 out_p.t1183 8.126
R3272 out_p.n7 out_p.t1037 8.126
R3273 out_p.n7 out_p.t199 8.126
R3274 out_p.n8 out_p.t875 8.126
R3275 out_p.n8 out_p.t1276 8.126
R3276 out_p.n9 out_p.t1139 8.126
R3277 out_p.n9 out_p.t1393 8.126
R3278 out_p.n183 out_p.t734 8.126
R3279 out_p.n183 out_p.t885 8.126
R3280 out_p.n184 out_p.t1561 8.126
R3281 out_p.n184 out_p.t1538 8.126
R3282 out_p.n185 out_p.t1368 8.126
R3283 out_p.n185 out_p.t474 8.126
R3284 out_p.n186 out_p.t454 8.126
R3285 out_p.n186 out_p.t1069 8.126
R3286 out_p.n187 out_p.t841 8.126
R3287 out_p.n187 out_p.t1214 8.126
R3288 out_p.n188 out_p.t1062 8.126
R3289 out_p.n188 out_p.t1627 8.126
R3290 out_p.n189 out_p.t278 8.126
R3291 out_p.n189 out_p.t453 8.126
R3292 out_p.n190 out_p.t249 8.126
R3293 out_p.n190 out_p.t165 8.126
R3294 out_p.n191 out_p.t1412 8.126
R3295 out_p.n191 out_p.t325 8.126
R3296 out_p.n192 out_p.t800 8.126
R3297 out_p.n192 out_p.t1227 8.126
R3298 out_p.n195 out_p.t509 8.126
R3299 out_p.n195 out_p.t427 8.126
R3300 out_p.n196 out_p.t1455 8.126
R3301 out_p.n196 out_p.t320 8.126
R3302 out_p.n197 out_p.t1589 8.126
R3303 out_p.n197 out_p.t534 8.126
R3304 out_p.n198 out_p.t253 8.126
R3305 out_p.n198 out_p.t357 8.126
R3306 out_p.n199 out_p.t373 8.126
R3307 out_p.n199 out_p.t685 8.126
R3308 out_p.n200 out_p.t1144 8.126
R3309 out_p.n200 out_p.t1380 8.126
R3310 out_p.n201 out_p.t390 8.126
R3311 out_p.n201 out_p.t1629 8.126
R3312 out_p.n202 out_p.t204 8.126
R3313 out_p.n202 out_p.t432 8.126
R3314 out_p.n203 out_p.t631 8.126
R3315 out_p.n203 out_p.t647 8.126
R3316 out_p.n204 out_p.t338 8.126
R3317 out_p.n204 out_p.t624 8.126
R3318 out_p.n207 out_p.t715 8.126
R3319 out_p.n207 out_p.t889 8.126
R3320 out_p.n208 out_p.t1602 8.126
R3321 out_p.n208 out_p.t1555 8.126
R3322 out_p.n209 out_p.t220 8.126
R3323 out_p.n209 out_p.t419 8.126
R3324 out_p.n210 out_p.t1018 8.126
R3325 out_p.n210 out_p.t504 8.126
R3326 out_p.n211 out_p.t1233 8.126
R3327 out_p.n211 out_p.t286 8.126
R3328 out_p.n212 out_p.t339 8.126
R3329 out_p.n212 out_p.t625 8.126
R3330 out_p.n213 out_p.t1092 8.126
R3331 out_p.n213 out_p.t161 8.126
R3332 out_p.n214 out_p.t726 8.126
R3333 out_p.n214 out_p.t934 8.126
R3334 out_p.n215 out_p.t1544 8.126
R3335 out_p.n215 out_p.t231 8.126
R3336 out_p.n216 out_p.t857 8.126
R3337 out_p.n216 out_p.t573 8.126
R3338 out_p.n219 out_p.t1563 8.126
R3339 out_p.n219 out_p.t173 8.126
R3340 out_p.n220 out_p.t866 8.126
R3341 out_p.n220 out_p.t938 8.126
R3342 out_p.n221 out_p.t992 8.126
R3343 out_p.n221 out_p.t1502 8.126
R3344 out_p.n222 out_p.t1115 8.126
R3345 out_p.n222 out_p.t1364 8.126
R3346 out_p.n223 out_p.t1496 8.126
R3347 out_p.n223 out_p.t1107 8.126
R3348 out_p.n224 out_p.t833 8.126
R3349 out_p.n224 out_p.t514 8.126
R3350 out_p.n225 out_p.t1371 8.126
R3351 out_p.n225 out_p.t1057 8.126
R3352 out_p.n226 out_p.t853 8.126
R3353 out_p.n226 out_p.t793 8.126
R3354 out_p.n227 out_p.t619 8.126
R3355 out_p.n227 out_p.t355 8.126
R3356 out_p.n228 out_p.t606 8.126
R3357 out_p.n228 out_p.t1565 8.126
R3358 out_p.n231 out_p.t1623 8.126
R3359 out_p.n231 out_p.t377 8.126
R3360 out_p.n232 out_p.t1248 8.126
R3361 out_p.n232 out_p.t1312 8.126
R3362 out_p.n233 out_p.t1032 8.126
R3363 out_p.n233 out_p.t1652 8.126
R3364 out_p.n234 out_p.t753 8.126
R3365 out_p.n234 out_p.t1272 8.126
R3366 out_p.n235 out_p.t923 8.126
R3367 out_p.n235 out_p.t228 8.126
R3368 out_p.n236 out_p.t607 8.126
R3369 out_p.n236 out_p.t1134 8.126
R3370 out_p.n237 out_p.t1202 8.126
R3371 out_p.n237 out_p.t441 8.126
R3372 out_p.n238 out_p.t689 8.126
R3373 out_p.n238 out_p.t1493 8.126
R3374 out_p.n239 out_p.t829 8.126
R3375 out_p.n239 out_p.t1506 8.126
R3376 out_p.n240 out_p.t207 8.126
R3377 out_p.n240 out_p.t196 8.126
R3378 out_p.n243 out_p.t1586 8.126
R3379 out_p.n243 out_p.t1309 8.126
R3380 out_p.n244 out_p.t1401 8.126
R3381 out_p.n244 out_p.t461 8.126
R3382 out_p.n245 out_p.t642 8.126
R3383 out_p.n245 out_p.t876 8.126
R3384 out_p.n246 out_p.t654 8.126
R3385 out_p.n246 out_p.t797 8.126
R3386 out_p.n247 out_p.t227 8.126
R3387 out_p.n247 out_p.t719 8.126
R3388 out_p.n248 out_p.t638 8.126
R3389 out_p.n248 out_p.t640 8.126
R3390 out_p.n249 out_p.t1478 8.126
R3391 out_p.n249 out_p.t1648 8.126
R3392 out_p.n250 out_p.t707 8.126
R3393 out_p.n250 out_p.t1654 8.126
R3394 out_p.n251 out_p.t667 8.126
R3395 out_p.n251 out_p.t1488 8.126
R3396 out_p.n252 out_p.t1101 8.126
R3397 out_p.n252 out_p.t943 8.126
R3398 out_p.n255 out_p.t672 8.126
R3399 out_p.n255 out_p.t819 8.126
R3400 out_p.n256 out_p.t680 8.126
R3401 out_p.n256 out_p.t1569 8.126
R3402 out_p.n257 out_p.t1362 8.126
R3403 out_p.n257 out_p.t846 8.126
R3404 out_p.n258 out_p.t1339 8.126
R3405 out_p.n258 out_p.t566 8.126
R3406 out_p.n259 out_p.t1291 8.126
R3407 out_p.n259 out_p.t488 8.126
R3408 out_p.n260 out_p.t635 8.126
R3409 out_p.n260 out_p.t202 8.126
R3410 out_p.n261 out_p.t1466 8.126
R3411 out_p.n261 out_p.t872 8.126
R3412 out_p.n262 out_p.t1433 8.126
R3413 out_p.n262 out_p.t349 8.126
R3414 out_p.n263 out_p.t1347 8.126
R3415 out_p.n263 out_p.t563 8.126
R3416 out_p.n264 out_p.t1299 8.126
R3417 out_p.n264 out_p.t1201 8.126
R3418 out_p.n267 out_p.t787 8.126
R3419 out_p.n267 out_p.t908 8.126
R3420 out_p.n268 out_p.t1038 8.126
R3421 out_p.n268 out_p.t540 8.126
R3422 out_p.n269 out_p.t1325 8.126
R3423 out_p.n269 out_p.t449 8.126
R3424 out_p.n270 out_p.t914 8.126
R3425 out_p.n270 out_p.t1310 8.126
R3426 out_p.n271 out_p.t1120 8.126
R3427 out_p.n271 out_p.t1152 8.126
R3428 out_p.n272 out_p.t1242 8.126
R3429 out_p.n272 out_p.t776 8.126
R3430 out_p.n273 out_p.t513 8.126
R3431 out_p.n273 out_p.t656 8.126
R3432 out_p.n274 out_p.t1344 8.126
R3433 out_p.n274 out_p.t326 8.126
R3434 out_p.n275 out_p.t650 8.126
R3435 out_p.n275 out_p.t1473 8.126
R3436 out_p.n276 out_p.t1187 8.126
R3437 out_p.n276 out_p.t275 8.126
R3438 out_p.n279 out_p.t1289 8.126
R3439 out_p.n279 out_p.t545 8.126
R3440 out_p.n280 out_p.t542 8.126
R3441 out_p.n280 out_p.t1225 8.126
R3442 out_p.n281 out_p.t879 8.126
R3443 out_p.n281 out_p.t1000 8.126
R3444 out_p.n282 out_p.t505 8.126
R3445 out_p.n282 out_p.t842 8.126
R3446 out_p.n283 out_p.t287 8.126
R3447 out_p.n283 out_p.t407 8.126
R3448 out_p.n284 out_p.t188 8.126
R3449 out_p.n284 out_p.t1336 8.126
R3450 out_p.n285 out_p.t158 8.126
R3451 out_p.n285 out_p.t740 8.126
R3452 out_p.n286 out_p.t743 8.126
R3453 out_p.n286 out_p.t652 8.126
R3454 out_p.n287 out_p.t230 8.126
R3455 out_p.n287 out_p.t1207 8.126
R3456 out_p.n288 out_p.t572 8.126
R3457 out_p.n288 out_p.t1270 8.126
R3458 out_p.n291 out_p.t468 8.126
R3459 out_p.n291 out_p.t1112 8.126
R3460 out_p.n292 out_p.t939 8.126
R3461 out_p.n292 out_p.t1603 8.126
R3462 out_p.n293 out_p.t1122 8.126
R3463 out_p.n293 out_p.t221 8.126
R3464 out_p.n294 out_p.t837 8.126
R3465 out_p.n294 out_p.t663 8.126
R3466 out_p.n295 out_p.t1106 8.126
R3467 out_p.n295 out_p.t288 8.126
R3468 out_p.n296 out_p.t578 8.126
R3469 out_p.n296 out_p.t1494 8.126
R3470 out_p.n297 out_p.t1056 8.126
R3471 out_p.n297 out_p.t1159 8.126
R3472 out_p.n298 out_p.t1437 8.126
R3473 out_p.n298 out_p.t658 8.126
R3474 out_p.n299 out_p.t1584 8.126
R3475 out_p.n299 out_p.t1283 8.126
R3476 out_p.n300 out_p.t259 8.126
R3477 out_p.n300 out_p.t815 8.126
R3478 out_p.n303 out_p.t1439 8.126
R3479 out_p.n303 out_p.t1047 8.126
R3480 out_p.n304 out_p.t981 8.126
R3481 out_p.n304 out_p.t1414 8.126
R3482 out_p.n305 out_p.t335 8.126
R3483 out_p.n305 out_p.t1086 8.126
R3484 out_p.n306 out_p.t1172 8.126
R3485 out_p.n306 out_p.t794 8.126
R3486 out_p.n307 out_p.t579 8.126
R3487 out_p.n307 out_p.t1495 8.126
R3488 out_p.n308 out_p.t906 8.126
R3489 out_p.n308 out_p.t470 8.126
R3490 out_p.n309 out_p.t684 8.126
R3491 out_p.n309 out_p.t1257 8.126
R3492 out_p.n310 out_p.t736 8.126
R3493 out_p.n310 out_p.t1650 8.126
R3494 out_p.n311 out_p.t496 8.126
R3495 out_p.n311 out_p.t823 8.126
R3496 out_p.n312 out_p.t486 8.126
R3497 out_p.n312 out_p.t1049 8.126
R3498 out_p.n315 out_p.t1280 8.126
R3499 out_p.n315 out_p.t690 8.126
R3500 out_p.n316 out_p.t502 8.126
R3501 out_p.n316 out_p.t1644 8.126
R3502 out_p.n317 out_p.t1040 8.126
R3503 out_p.n317 out_p.t1177 8.126
R3504 out_p.n318 out_p.t883 8.126
R3505 out_p.n318 out_p.t1264 8.126
R3506 out_p.n319 out_p.t517 8.126
R3507 out_p.n319 out_p.t392 8.126
R3508 out_p.n320 out_p.t835 8.126
R3509 out_p.n320 out_p.t1269 8.126
R3510 out_p.n321 out_p.t1477 8.126
R3511 out_p.n321 out_p.t1332 8.126
R3512 out_p.n322 out_p.t748 8.126
R3513 out_p.n322 out_p.t805 8.126
R3514 out_p.n323 out_p.t589 8.126
R3515 out_p.n323 out_p.t1097 8.126
R3516 out_p.n324 out_p.t1626 8.126
R3517 out_p.n324 out_p.t1220 8.126
R3518 out_p.n327 out_p.t246 8.126
R3519 out_p.n327 out_p.t1596 8.126
R3520 out_p.n328 out_p.t1539 8.126
R3521 out_p.n328 out_p.t1470 8.126
R3522 out_p.n329 out_p.t475 8.126
R3523 out_p.n329 out_p.t1425 8.126
R3524 out_p.n330 out_p.t281 8.126
R3525 out_p.n330 out_p.t181 8.126
R3526 out_p.n331 out_p.t818 8.126
R3527 out_p.n331 out_p.t1192 8.126
R3528 out_p.n332 out_p.t313 8.126
R3529 out_p.n332 out_p.t840 8.126
R3530 out_p.n333 out_p.t1246 8.126
R3531 out_p.n333 out_p.t649 8.126
R3532 out_p.n334 out_p.t1026 8.126
R3533 out_p.n334 out_p.t746 8.126
R3534 out_p.n335 out_p.t1143 8.126
R3535 out_p.n335 out_p.t365 8.126
R3536 out_p.n336 out_p.t493 8.126
R3537 out_p.n336 out_p.t1543 8.126
R3538 out_p.n339 out_p.t1268 8.126
R3539 out_p.n339 out_p.t1391 8.126
R3540 out_p.n340 out_p.t849 8.126
R3541 out_p.n340 out_p.t1131 8.126
R3542 out_p.n341 out_p.t562 8.126
R3543 out_p.n341 out_p.t848 8.126
R3544 out_p.n342 out_p.t1230 8.126
R3545 out_p.n342 out_p.t1141 8.126
R3546 out_p.n343 out_p.t601 8.126
R3547 out_p.n343 out_p.t953 8.126
R3548 out_p.n344 out_p.t790 8.126
R3549 out_p.n344 out_p.t171 8.126
R3550 out_p.n345 out_p.t500 8.126
R3551 out_p.n345 out_p.t899 8.126
R3552 out_p.n346 out_p.t1274 8.126
R3553 out_p.n346 out_p.t195 8.126
R3554 out_p.n347 out_p.t1315 8.126
R3555 out_p.n347 out_p.t1103 8.126
R3556 out_p.n348 out_p.t398 8.126
R3557 out_p.n348 out_p.t560 8.126
R3558 out_p.n351 out_p.t186 8.126
R3559 out_p.n351 out_p.t784 8.126
R3560 out_p.n352 out_p.t847 8.126
R3561 out_p.n352 out_p.t1568 8.126
R3562 out_p.n353 out_p.t1373 8.126
R3563 out_p.n353 out_p.t208 8.126
R3564 out_p.n354 out_p.t256 8.126
R3565 out_p.n354 out_p.t1510 8.126
R3566 out_p.n355 out_p.t508 8.126
R3567 out_p.n355 out_p.t426 8.126
R3568 out_p.n356 out_p.t399 8.126
R3569 out_p.n356 out_p.t561 8.126
R3570 out_p.n357 out_p.t331 8.126
R3571 out_p.n357 out_p.t695 8.126
R3572 out_p.n358 out_p.t314 8.126
R3573 out_p.n358 out_p.t728 8.126
R3574 out_p.n359 out_p.t777 8.126
R3575 out_p.n359 out_p.t554 8.126
R3576 out_p.n360 out_p.t668 8.126
R3577 out_p.n360 out_p.t564 8.126
R3578 out_p.n363 out_p.t1004 8.126
R3579 out_p.n363 out_p.t1392 8.126
R3580 out_p.n364 out_p.t333 8.126
R3581 out_p.n364 out_p.t1363 8.126
R3582 out_p.n365 out_p.t241 8.126
R3583 out_p.n365 out_p.t990 8.126
R3584 out_p.n366 out_p.t1030 8.126
R3585 out_p.n366 out_p.t812 8.126
R3586 out_p.n367 out_p.t995 8.126
R3587 out_p.n367 out_p.t888 8.126
R3588 out_p.n368 out_p.t1410 8.126
R3589 out_p.n368 out_p.t565 8.126
R3590 out_p.n369 out_p.t677 8.126
R3591 out_p.n369 out_p.t1306 8.126
R3592 out_p.n370 out_p.t614 8.126
R3593 out_p.n370 out_p.t1266 8.126
R3594 out_p.n371 out_p.t1145 8.126
R3595 out_p.n371 out_p.t1243 8.126
R3596 out_p.n372 out_p.t310 8.126
R3597 out_p.n372 out_p.t1125 8.126
R3598 out_p.n375 out_p.t467 8.126
R3599 out_p.n375 out_p.t1411 8.126
R3600 out_p.n376 out_p.t1635 8.126
R3601 out_p.n376 out_p.t809 8.126
R3602 out_p.n377 out_p.t999 8.126
R3603 out_p.n377 out_p.t463 8.126
R3604 out_p.n378 out_p.t1552 8.126
R3605 out_p.n378 out_p.t1083 8.126
R3606 out_p.n379 out_p.t1443 8.126
R3607 out_p.n379 out_p.t347 8.126
R3608 out_p.n380 out_p.t438 8.126
R3609 out_p.n380 out_p.t1303 8.126
R3610 out_p.n381 out_p.t424 8.126
R3611 out_p.n381 out_p.t477 8.126
R3612 out_p.n382 out_p.t1260 8.126
R3613 out_p.n382 out_p.t1157 8.126
R3614 out_p.n383 out_p.t674 8.126
R3615 out_p.n383 out_p.t362 8.126
R3616 out_p.n384 out_p.t595 8.126
R3617 out_p.n384 out_p.t1566 8.126
R3618 out_p.n387 out_p.t1647 8.126
R3619 out_p.n387 out_p.t343 8.126
R3620 out_p.n388 out_p.t764 8.126
R3621 out_p.n388 out_p.t1132 8.126
R3622 out_p.n389 out_p.t224 8.126
R3623 out_p.n389 out_p.t1349 8.126
R3624 out_p.n390 out_p.t537 8.126
R3625 out_p.n390 out_p.t1440 8.126
R3626 out_p.n391 out_p.t439 8.126
R3627 out_p.n391 out_p.t482 8.126
R3628 out_p.n392 out_p.t870 8.126
R3629 out_p.n392 out_p.t1294 8.126
R3630 out_p.n393 out_p.t1330 8.126
R3631 out_p.n393 out_p.t178 8.126
R3632 out_p.n394 out_p.t1570 8.126
R3633 out_p.n394 out_p.t1458 8.126
R3634 out_p.n395 out_p.t1135 8.126
R3635 out_p.n395 out_p.t1229 8.126
R3636 out_p.n396 out_p.t350 8.126
R3637 out_p.n396 out_p.t1195 8.126
R3638 out_p.n399 out_p.t1505 8.126
R3639 out_p.n399 out_p.t1161 8.126
R3640 out_p.n400 out_p.t628 8.126
R3641 out_p.n400 out_p.t1535 8.126
R3642 out_p.n401 out_p.t1096 8.126
R3643 out_p.n401 out_p.t862 8.126
R3644 out_p.n402 out_p.t1258 8.126
R3645 out_p.n402 out_p.t282 8.126
R3646 out_p.n403 out_p.t367 8.126
R3647 out_p.n403 out_p.t897 8.126
R3648 out_p.n404 out_p.t664 8.126
R3649 out_p.n404 out_p.t284 8.126
R3650 out_p.n405 out_p.t910 8.126
R3651 out_p.n405 out_p.t298 8.126
R3652 out_p.n406 out_p.t185 8.126
R3653 out_p.n406 out_p.t1429 8.126
R3654 out_p.n407 out_p.t770 8.126
R3655 out_p.n407 out_p.t697 8.126
R3656 out_p.n408 out_p.t1461 8.126
R3657 out_p.n408 out_p.t236 8.126
R3658 out_p.n411 out_p.t1409 8.126
R3659 out_p.n411 out_p.t526 8.126
R3660 out_p.n412 out_p.t414 8.126
R3661 out_p.n412 out_p.t1427 8.126
R3662 out_p.n413 out_p.t874 8.126
R3663 out_p.n413 out_p.t673 8.126
R3664 out_p.n414 out_p.t1446 8.126
R3665 out_p.n414 out_p.t318 8.126
R3666 out_p.n415 out_p.t1390 8.126
R3667 out_p.n415 out_p.t1444 8.126
R3668 out_p.n416 out_p.t970 8.126
R3669 out_p.n416 out_p.t237 8.126
R3670 out_p.n417 out_p.t1163 8.126
R3671 out_p.n417 out_p.t609 8.126
R3672 out_p.n418 out_p.t211 8.126
R3673 out_p.n418 out_p.t1068 8.126
R3674 out_p.n419 out_p.t1221 8.126
R3675 out_p.n419 out_p.t834 8.126
R3676 out_p.n420 out_p.t1205 8.126
R3677 out_p.n420 out_p.t1432 8.126
R3678 out_p.n423 out_p.t1638 8.126
R3679 out_p.n423 out_p.t594 8.126
R3680 out_p.n424 out_p.t1024 8.126
R3681 out_p.n424 out_p.t1041 8.126
R3682 out_p.n425 out_p.t307 8.126
R3683 out_p.n425 out_p.t324 8.126
R3684 out_p.n426 out_p.t507 8.126
R3685 out_p.n426 out_p.t395 8.126
R3686 out_p.n427 out_p.t371 8.126
R3687 out_p.n427 out_p.t945 8.126
R3688 out_p.n428 out_p.t510 8.126
R3689 out_p.n428 out_p.t245 8.126
R3690 out_p.n429 out_p.t358 8.126
R3691 out_p.n429 out_p.t1537 8.126
R3692 out_p.n430 out_p.t1358 8.126
R3693 out_p.n430 out_p.t1188 8.126
R3694 out_p.n431 out_p.t170 8.126
R3695 out_p.n431 out_p.t312 8.126
R3696 out_p.n432 out_p.t428 8.126
R3697 out_p.n432 out_p.t411 8.126
R3698 out_p.n435 out_p.t679 8.126
R3699 out_p.n435 out_p.t511 8.126
R3700 out_p.n436 out_p.t584 8.126
R3701 out_p.n436 out_p.t1110 8.126
R3702 out_p.n437 out_p.t630 8.126
R3703 out_p.n437 out_p.t646 8.126
R3704 out_p.n438 out_p.t721 8.126
R3705 out_p.n438 out_p.t1450 8.126
R3706 out_p.n439 out_p.t994 8.126
R3707 out_p.n439 out_p.t1256 8.126
R3708 out_p.n440 out_p.t1147 8.126
R3709 out_p.n440 out_p.t1403 8.126
R3710 out_p.n441 out_p.t676 8.126
R3711 out_p.n441 out_p.t1094 8.126
R3712 out_p.n442 out_p.t662 8.126
R3713 out_p.n442 out_p.t1457 8.126
R3714 out_p.n443 out_p.t1232 8.126
R3715 out_p.n443 out_p.t1381 8.126
R3716 out_p.n444 out_p.t311 8.126
R3717 out_p.n444 out_p.t1422 8.126
R3718 out_p.n447 out_p.t1119 8.126
R3719 out_p.n447 out_p.t429 8.126
R3720 out_p.n448 out_p.t268 8.126
R3721 out_p.n448 out_p.t1454 8.126
R3722 out_p.n449 out_p.t973 8.126
R3723 out_p.n449 out_p.t622 8.126
R3724 out_p.n450 out_p.t1033 8.126
R3725 out_p.n450 out_p.t644 8.126
R3726 out_p.n451 out_p.t1292 8.126
R3727 out_p.n451 out_p.t372 8.126
R3728 out_p.n452 out_p.t1080 8.126
R3729 out_p.n452 out_p.t1423 8.126
R3730 out_p.n453 out_p.t928 8.126
R3731 out_p.n453 out_p.t901 8.126
R3732 out_p.n454 out_p.t1082 8.126
R3733 out_p.n454 out_p.t836 8.126
R3734 out_p.n455 out_p.t346 8.126
R3735 out_p.n455 out_p.t189 8.126
R3736 out_p.n456 out_p.t1420 8.126
R3737 out_p.n456 out_p.t174 8.126
R3738 out_p.n459 out_p.t1402 8.126
R3739 out_p.n459 out_p.t254 8.126
R3740 out_p.n460 out_p.t375 8.126
R3741 out_p.n460 out_p.t1479 8.126
R3742 out_p.n461 out_p.t691 8.126
R3743 out_p.n461 out_p.t1382 8.126
R3744 out_p.n462 out_p.t983 8.126
R3745 out_p.n462 out_p.t877 8.126
R3746 out_p.n463 out_p.t1081 8.126
R3747 out_p.n463 out_p.t912 8.126
R3748 out_p.n464 out_p.t1421 8.126
R3749 out_p.n464 out_p.t530 8.126
R3750 out_p.n465 out_p.t1624 8.126
R3751 out_p.n465 out_p.t183 8.126
R3752 out_p.n466 out_p.t1054 8.126
R3753 out_p.n466 out_p.t712 8.126
R3754 out_p.n467 out_p.t1302 8.126
R3755 out_p.n467 out_p.t1442 8.126
R3756 out_p.n468 out_p.t804 8.126
R3757 out_p.n468 out_p.t546 8.126
R3758 out_p.n471 out_p.t1630 8.126
R3759 out_p.n471 out_p.t1146 8.126
R3760 out_p.n472 out_p.t462 8.126
R3761 out_p.n472 out_p.t273 8.126
R3762 out_p.n473 out_p.t1597 8.126
R3763 out_p.n473 out_p.t1524 8.126
R3764 out_p.n474 out_p.t322 8.126
R3765 out_p.n474 out_p.t988 8.126
R3766 out_p.n475 out_p.t1160 8.126
R3767 out_p.n475 out_p.t531 8.126
R3768 out_p.n476 out_p.t798 8.126
R3769 out_p.n476 out_p.t1504 8.126
R3770 out_p.n477 out_p.t213 8.126
R3771 out_p.n477 out_p.t1558 8.126
R3772 out_p.n478 out_p.t788 8.126
R3773 out_p.n478 out_p.t947 8.126
R3774 out_p.n479 out_p.t1567 8.126
R3775 out_p.n479 out_p.t527 8.126
R3776 out_p.n480 out_p.t214 8.126
R3777 out_p.n480 out_p.t749 8.126
R3778 out_p.n483 out_p.t1265 8.126
R3779 out_p.n483 out_p.t1136 8.126
R3780 out_p.n484 out_p.t412 8.126
R3781 out_p.n484 out_p.t745 8.126
R3782 out_p.n485 out_p.t696 8.126
R3783 out_p.n485 out_p.t1445 8.126
R3784 out_p.n486 out_p.t1531 8.126
R3785 out_p.n486 out_p.t1369 8.126
R3786 out_p.n487 out_p.t452 8.126
R3787 out_p.n487 out_p.t1219 8.126
R3788 out_p.n488 out_p.t222 8.126
R3789 out_p.n488 out_p.t739 8.126
R3790 out_p.n489 out_p.t1557 8.126
R3791 out_p.n489 out_p.t949 8.126
R3792 out_p.n490 out_p.t775 8.126
R3793 out_p.n490 out_p.t1079 8.126
R3794 out_p.n491 out_p.t285 8.126
R3795 out_p.n491 out_p.t366 8.126
R3796 out_p.n492 out_p.t1338 8.126
R3797 out_p.n492 out_p.t569 8.126
R3798 out_p.n495 out_p.t567 8.126
R3799 out_p.n495 out_p.t223 8.126
R3800 out_p.n496 out_p.t1025 8.126
R3801 out_p.n496 out_p.t1352 8.126
R3802 out_p.n497 out_p.t1102 8.126
R3803 out_p.n497 out_p.t881 8.126
R3804 out_p.n498 out_p.t1151 8.126
R3805 out_p.n498 out_p.t1520 8.126
R3806 out_p.n499 out_p.t1642 8.126
R3807 out_p.n499 out_p.t931 8.126
R3808 out_p.n500 out_p.t1591 8.126
R3809 out_p.n500 out_p.t1321 8.126
R3810 out_p.n501 out_p.t359 8.126
R3811 out_p.n501 out_p.t490 8.126
R3812 out_p.n502 out_p.t1253 8.126
R3813 out_p.n502 out_p.t933 8.126
R3814 out_p.n503 out_p.t1005 8.126
R3815 out_p.n503 out_p.t600 8.126
R3816 out_p.n504 out_p.t205 8.126
R3817 out_p.n504 out_p.t433 8.126
R3818 out_p.n507 out_p.t1023 8.126
R3819 out_p.n507 out_p.t964 8.126
R3820 out_p.n508 out_p.t255 8.126
R3821 out_p.n508 out_p.t577 8.126
R3822 out_p.n509 out_p.t1441 8.126
R3823 out_p.n509 out_p.t1314 8.126
R3824 out_p.n510 out_p.t710 8.126
R3825 out_p.n510 out_p.t1117 8.126
R3826 out_p.n511 out_p.t167 8.126
R3827 out_p.n511 out_p.t952 8.126
R3828 out_p.n512 out_p.t408 8.126
R3829 out_p.n512 out_p.t678 8.126
R3830 out_p.n513 out_p.t1634 8.126
R3831 out_p.n513 out_p.t827 8.126
R3832 out_p.n514 out_p.t858 8.126
R3833 out_p.n514 out_p.t1532 8.126
R3834 out_p.n515 out_p.t519 8.126
R3835 out_p.n515 out_p.t791 8.126
R3836 out_p.n516 out_p.t1323 8.126
R3837 out_p.n516 out_p.t444 8.126
R3838 out_p.n519 out_p.t751 8.126
R3839 out_p.n519 out_p.t1605 8.126
R3840 out_p.n520 out_p.t1621 8.126
R3841 out_p.n520 out_p.t851 8.126
R3842 out_p.n521 out_p.t789 8.126
R3843 out_p.n521 out_p.t1156 8.126
R3844 out_p.n522 out_p.t239 8.126
R3845 out_p.n522 out_p.t855 8.126
R3846 out_p.n523 out_p.t409 8.126
R3847 out_p.n523 out_p.t982 8.126
R3848 out_p.n524 out_p.t1374 8.126
R3849 out_p.n524 out_p.t1367 8.126
R3850 out_p.n525 out_p.t1518 8.126
R3851 out_p.n525 out_p.t1089 8.126
R3852 out_p.n526 out_p.t660 8.126
R3853 out_p.n526 out_p.t1263 8.126
R3854 out_p.n527 out_p.t946 8.126
R3855 out_p.n527 out_p.t1191 8.126
R3856 out_p.n528 out_p.t1556 8.126
R3857 out_p.n528 out_p.t948 8.126
R3858 out_p.n531 out_p.t182 8.126
R3859 out_p.n531 out_p.t250 8.126
R3860 out_p.n532 out_p.t1480 8.126
R3861 out_p.n532 out_p.t1631 8.126
R3862 out_p.n533 out_p.t911 8.126
R3863 out_p.n533 out_p.t583 8.126
R3864 out_p.n534 out_p.t1011 8.126
R3865 out_p.n534 out_p.t559 8.126
R3866 out_p.n535 out_p.t1375 8.126
R3867 out_p.n535 out_p.t217 8.126
R3868 out_p.n536 out_p.t168 8.126
R3869 out_p.n536 out_p.t1254 8.126
R3870 out_p.n537 out_p.t887 8.126
R3871 out_p.n537 out_p.t301 8.126
R3872 out_p.n538 out_p.t361 8.126
R3873 out_p.n538 out_p.t709 8.126
R3874 out_p.n539 out_p.t582 8.126
R3875 out_p.n539 out_p.t927 8.126
R3876 out_p.n540 out_p.t541 8.126
R3877 out_p.n540 out_p.t681 8.126
R3878 out_p.n543 out_p.t1379 8.126
R3879 out_p.n543 out_p.t941 8.126
R3880 out_p.n544 out_p.t1640 8.126
R3881 out_p.n544 out_p.t772 8.126
R3882 out_p.n545 out_p.t184 8.126
R3883 out_p.n545 out_p.t1428 8.126
R3884 out_p.n546 out_p.t369 8.126
R3885 out_p.n546 out_p.t383 8.126
R3886 out_p.n547 out_p.t295 8.126
R3887 out_p.n547 out_p.t1530 8.126
R3888 out_p.n548 out_p.t529 8.126
R3889 out_p.n548 out_p.t603 8.126
R3890 out_p.n549 out_p.t1176 8.126
R3891 out_p.n549 out_p.t1426 8.126
R3892 out_p.n550 out_p.t1245 8.126
R3893 out_p.n550 out_p.t610 8.126
R3894 out_p.n551 out_p.t723 8.126
R3895 out_p.n551 out_p.t975 8.126
R3896 out_p.n552 out_p.t435 8.126
R3897 out_p.n552 out_p.t478 8.126
R3898 out_p.n555 out_p.t722 8.126
R3899 out_p.n555 out_p.t974 8.126
R3900 out_p.n556 out_p.t965 8.126
R3901 out_p.n556 out_p.t1639 8.126
R3902 out_p.n557 out_p.t1342 8.126
R3903 out_p.n557 out_p.t966 8.126
R3904 out_p.n558 out_p.t242 8.126
R3905 out_p.n558 out_p.t918 8.126
R3906 out_p.n559 out_p.t191 8.126
R3907 out_p.n559 out_p.t506 8.126
R3908 out_p.n560 out_p.t1067 8.126
R3909 out_p.n560 out_p.t1405 8.126
R3910 out_p.n561 out_p.t523 8.126
R3911 out_p.n561 out_p.t987 8.126
R3912 out_p.n562 out_p.t321 8.126
R3913 out_p.n562 out_p.t1111 8.126
R3914 out_p.n563 out_p.t1581 8.126
R3915 out_p.n563 out_p.t1252 8.126
R3916 out_p.n564 out_p.t1029 8.126
R3917 out_p.n564 out_p.t731 8.126
R3918 out_p.n567 out_p.t309 8.126
R3919 out_p.n567 out_p.t1168 8.126
R3920 out_p.n568 out_p.t370 8.126
R3921 out_p.n568 out_p.t930 8.126
R3922 out_p.n569 out_p.t645 8.126
R3923 out_p.n569 out_p.t1031 8.126
R3924 out_p.n570 out_p.t586 8.126
R3925 out_p.n570 out_p.t292 8.126
R3926 out_p.n571 out_p.t1087 8.126
R3927 out_p.n571 out_p.t1503 8.126
R3928 out_p.n572 out_p.t457 8.126
R3929 out_p.n572 out_p.t379 8.126
R3930 out_p.n573 out_p.t332 8.126
R3931 out_p.n573 out_p.t1042 8.126
R3932 out_p.n574 out_p.t1583 8.126
R3933 out_p.n574 out_p.t1355 8.126
R3934 out_p.n575 out_p.t720 8.126
R3935 out_p.n575 out_p.t437 8.126
R3936 out_p.n576 out_p.t839 8.126
R3937 out_p.n576 out_p.t621 8.126
R3938 out_p.n579 out_p.t1035 8.126
R3939 out_p.n579 out_p.t402 8.126
R3940 out_p.n580 out_p.t1590 8.126
R3941 out_p.n580 out_p.t1320 8.126
R3942 out_p.n581 out_p.t1606 8.126
R3943 out_p.n581 out_p.t305 8.126
R3944 out_p.n582 out_p.t447 8.126
R3945 out_p.n582 out_p.t997 8.126
R3946 out_p.n583 out_p.t1050 8.126
R3947 out_p.n583 out_p.t1612 8.126
R3948 out_p.n584 out_p.t1604 8.126
R3949 out_p.n584 out_p.t1406 8.126
R3950 out_p.n585 out_p.t1554 8.126
R3951 out_p.n585 out_p.t535 8.126
R3952 out_p.n586 out_p.t1184 8.126
R3953 out_p.n586 out_p.t1398 8.126
R3954 out_p.n587 out_p.t304 8.126
R3955 out_p.n587 out_p.t431 8.126
R3956 out_p.n588 out_p.t1238 8.126
R3957 out_p.n588 out_p.t574 8.126
R3958 out_p.n591 out_p.t378 8.126
R3959 out_p.n591 out_p.t865 8.126
R3960 out_p.n592 out_p.t1076 8.126
R3961 out_p.n592 out_p.t1019 8.126
R3962 out_p.n593 out_p.t989 8.126
R3963 out_p.n593 out_p.t1515 8.126
R3964 out_p.n594 out_p.t688 8.126
R3965 out_p.n594 out_p.t269 8.126
R3966 out_p.n595 out_p.t828 8.126
R3967 out_p.n595 out_p.t702 8.126
R3968 out_p.n596 out_p.t481 8.126
R3969 out_p.n596 out_p.t575 8.126
R3970 out_p.n597 out_p.t374 8.126
R3971 out_p.n597 out_p.t878 8.126
R3972 out_p.n598 out_p.t854 8.126
R3973 out_p.n598 out_p.t808 8.126
R3974 out_p.n599 out_p.t783 8.126
R3975 out_p.n599 out_p.t251 8.126
R3976 out_p.n600 out_p.t1181 8.126
R3977 out_p.n600 out_p.t1462 8.126
R3978 out_p.n603 out_p.t620 8.126
R3979 out_p.n603 out_p.t1593 8.126
R3980 out_p.n604 out_p.t1553 8.126
R3981 out_p.n604 out_p.t1098 8.126
R3982 out_p.n605 out_p.t1190 8.126
R3983 out_p.n605 out_p.t518 8.126
R3984 out_p.n606 out_p.t1513 8.126
R3985 out_p.n606 out_p.t1317 8.126
R3986 out_p.n607 out_p.t666 8.126
R3987 out_p.n607 out_p.t1241 8.126
R3988 out_p.n608 out_p.t940 8.126
R3989 out_p.n608 out_p.t1327 8.126
R3990 out_p.n609 out_p.t229 8.126
R3991 out_p.n609 out_p.t1497 8.126
R3992 out_p.n610 out_p.t558 8.126
R3993 out_p.n610 out_p.t238 8.126
R3994 out_p.n611 out_p.t216 8.126
R3995 out_p.n611 out_p.t557 8.126
R3996 out_p.n612 out_p.t1322 8.126
R3997 out_p.n612 out_p.t1378 8.126
R3998 out_p.n615 out_p.t1366 8.126
R3999 out_p.n615 out_p.t950 8.126
R4000 out_p.n616 out_p.t1641 8.126
R4001 out_p.n616 out_p.t773 8.126
R4002 out_p.n617 out_p.t963 8.126
R4003 out_p.n617 out_p.t1447 8.126
R4004 out_p.n618 out_p.t368 8.126
R4005 out_p.n618 out_p.t382 8.126
R4006 out_p.n619 out_p.t294 8.126
R4007 out_p.n619 out_p.t1487 8.126
R4008 out_p.n620 out_p.t528 8.126
R4009 out_p.n620 out_p.t602 8.126
R4010 out_p.n621 out_p.t1609 8.126
R4011 out_p.n621 out_p.t1387 8.126
R4012 out_p.n622 out_p.t1058 8.126
R4013 out_p.n622 out_p.t1180 8.126
R4014 out_p.n623 out_p.t1418 8.126
R4015 out_p.n623 out_p.t774 8.126
R4016 out_p.n624 out_p.t394 8.126
R4017 out_p.n624 out_p.t479 8.126
R4018 out_p.n627 out_p.t1526 8.126
R4019 out_p.n627 out_p.t1573 8.126
R4020 out_p.n628 out_p.t550 8.126
R4021 out_p.n628 out_p.t1007 8.126
R4022 out_p.n629 out_p.t1178 8.126
R4023 out_p.n629 out_p.t1350 8.126
R4024 out_p.n630 out_p.t553 8.126
R4025 out_p.n630 out_p.t1389 8.126
R4026 out_p.n631 out_p.t336 8.126
R4027 out_p.n631 out_p.t1341 8.126
R4028 out_p.n632 out_p.t1632 8.126
R4029 out_p.n632 out_p.t760 8.126
R4030 out_p.n633 out_p.t489 8.126
R4031 out_p.n633 out_p.t1517 8.126
R4032 out_p.n634 out_p.t781 8.126
R4033 out_p.n634 out_p.t816 8.126
R4034 out_p.n635 out_p.t201 8.126
R4035 out_p.n635 out_p.t902 8.126
R4036 out_p.n636 out_p.t860 8.126
R4037 out_p.n636 out_p.t193 8.126
R4038 out_p.n639 out_p.t329 8.126
R4039 out_p.n639 out_p.t1002 8.126
R4040 out_p.n640 out_p.t1231 8.126
R4041 out_p.n640 out_p.t738 8.126
R4042 out_p.n641 out_p.t1175 8.126
R4043 out_p.n641 out_p.t932 8.126
R4044 out_p.n642 out_p.t1449 8.126
R4045 out_p.n642 out_p.t984 8.126
R4046 out_p.n643 out_p.t1633 8.126
R4047 out_p.n643 out_p.t1206 8.126
R4048 out_p.n644 out_p.t861 8.126
R4049 out_p.n644 out_p.t397 8.126
R4050 out_p.n645 out_p.t1153 8.126
R4051 out_p.n645 out_p.t576 8.126
R4052 out_p.n646 out_p.t1376 8.126
R4053 out_p.n646 out_p.t1485 8.126
R4054 out_p.n647 out_p.t1404 8.126
R4055 out_p.n647 out_p.t190 8.126
R4056 out_p.n648 out_p.t291 8.126
R4057 out_p.n648 out_p.t1072 8.126
R4058 out_p.n651 out_p.t1186 8.126
R4059 out_p.n651 out_p.t960 8.126
R4060 out_p.n652 out_p.t1304 8.126
R4061 out_p.n652 out_p.t1511 8.126
R4062 out_p.n653 out_p.t1051 8.126
R4063 out_p.n653 out_p.t1615 8.126
R4064 out_p.n654 out_p.t425 8.126
R4065 out_p.n654 out_p.t780 8.126
R4066 out_p.n655 out_p.t354 8.126
R4067 out_p.n655 out_p.t1501 8.126
R4068 out_p.n656 out_p.t1197 8.126
R4069 out_p.n656 out_p.t1073 8.126
R4070 out_p.n657 out_p.t596 8.126
R4071 out_p.n657 out_p.t1121 8.126
R4072 out_p.n658 out_p.t996 8.126
R4073 out_p.n658 out_p.t1043 8.126
R4074 out_p.n659 out_p.t334 8.126
R4075 out_p.n659 out_p.t1066 8.126
R4076 out_p.n660 out_p.t1600 8.126
R4077 out_p.n660 out_p.t1491 8.126
R4078 out_p.n663 out_p.t192 8.126
R4079 out_p.n663 out_p.t1271 8.126
R4080 out_p.n664 out_p.t356 8.126
R4081 out_p.n664 out_p.t1451 8.126
R4082 out_p.n665 out_p.t430 8.126
R4083 out_p.n665 out_p.t1022 8.126
R4084 out_p.n666 out_p.t1370 8.126
R4085 out_p.n666 out_p.t683 8.126
R4086 out_p.n667 out_p.t1071 8.126
R4087 out_p.n667 out_p.t1452 8.126
R4088 out_p.n668 out_p.t1601 8.126
R4089 out_p.n668 out_p.t1434 8.126
R4090 out_p.n669 out_p.t289 8.126
R4091 out_p.n669 out_p.t405 8.126
R4092 out_p.n670 out_p.t1649 8.126
R4093 out_p.n670 out_p.t446 8.126
R4094 out_p.n671 out_p.t1407 8.126
R4095 out_p.n671 out_p.t1551 8.126
R4096 out_p.n672 out_p.t1262 8.126
R4097 out_p.n672 out_p.t1301 8.126
R4098 out_p.n675 out_p.t226 8.126
R4099 out_p.n675 out_p.t456 8.126
R4100 out_p.n676 out_p.t762 8.126
R4101 out_p.n676 out_p.t1099 8.126
R4102 out_p.n677 out_p.t692 8.126
R4103 out_p.n677 out_p.t323 8.126
R4104 out_p.n678 out_p.t198 8.126
R4105 out_p.n678 out_p.t1431 8.126
R4106 out_p.n679 out_p.t588 8.126
R4107 out_p.n679 out_p.t263 8.126
R4108 out_p.n680 out_p.t786 8.126
R4109 out_p.n680 out_p.t1326 8.126
R4110 out_p.n681 out_p.t1498 8.126
R4111 out_p.n681 out_p.t272 8.126
R4112 out_p.n682 out_p.t873 8.126
R4113 out_p.n682 out_p.t1357 8.126
R4114 out_p.n683 out_p.t969 8.126
R4115 out_p.n683 out_p.t556 8.126
R4116 out_p.n684 out_p.t626 8.126
R4117 out_p.n684 out_p.t1059 8.126
R4118 out_p.n687 out_p.t297 8.126
R4119 out_p.n687 out_p.t641 8.126
R4120 out_p.n688 out_p.t484 8.126
R4121 out_p.n688 out_p.t1250 8.126
R4122 out_p.n689 out_p.t716 8.126
R4123 out_p.n689 out_p.t1064 8.126
R4124 out_p.n690 out_p.t164 8.126
R4125 out_p.n690 out_p.t1036 8.126
R4126 out_p.n691 out_p.t811 8.126
R4127 out_p.n691 out_p.t909 8.126
R4128 out_p.n692 out_p.t627 8.126
R4129 out_p.n692 out_p.t544 8.126
R4130 out_p.n693 out_p.t393 8.126
R4131 out_p.n693 out_p.t744 8.126
R4132 out_p.n694 out_p.t657 8.126
R4133 out_p.n694 out_p.t1467 8.126
R4134 out_p.n695 out_p.t1486 8.126
R4135 out_p.n695 out_p.t451 8.126
R4136 out_p.n696 out_p.t1287 8.126
R4137 out_p.n696 out_p.t341 8.126
R4138 out_p.n699 out_p.t400 8.126
R4139 out_p.n699 out_p.t1061 8.126
R4140 out_p.n700 out_p.t1198 8.126
R4141 out_p.n700 out_p.t778 8.126
R4142 out_p.n701 out_p.t825 8.126
R4143 out_p.n701 out_p.t1078 8.126
R4144 out_p.n702 out_p.t495 8.126
R4145 out_p.n702 out_p.t248 8.126
R4146 out_p.n703 out_p.t261 8.126
R4147 out_p.n703 out_p.t233 8.126
R4148 out_p.n704 out_p.t1508 8.126
R4149 out_p.n704 out_p.t218 8.126
R4150 out_p.n705 out_p.t1193 8.126
R4151 out_p.n705 out_p.t1534 8.126
R4152 out_p.n706 out_p.t741 8.126
R4153 out_p.n706 out_p.t1528 8.126
R4154 out_p.n707 out_p.t844 8.126
R4155 out_p.n707 out_p.t1384 8.126
R4156 out_p.n708 out_p.t613 8.126
R4157 out_p.n708 out_p.t328 8.126
R4158 out_p.n711 out_p.t1052 8.126
R4159 out_p.n711 out_p.t1063 8.126
R4160 out_p.n712 out_p.t521 8.126
R4161 out_p.n712 out_p.t869 8.126
R4162 out_p.n713 out_p.t1169 8.126
R4163 out_p.n713 out_p.t806 8.126
R4164 out_p.n714 out_p.t303 8.126
R4165 out_p.n714 out_p.t633 8.126
R4166 out_p.n715 out_p.t1200 8.126
R4167 out_p.n715 out_p.t634 8.126
R4168 out_p.n716 out_p.t1438 8.126
R4169 out_p.n716 out_p.t1046 8.126
R4170 out_p.n717 out_p.t386 8.126
R4171 out_p.n717 out_p.t1643 8.126
R4172 out_p.n718 out_p.t1093 8.126
R4173 out_p.n718 out_p.t925 8.126
R4174 out_p.n719 out_p.t459 8.126
R4175 out_p.n719 out_p.t571 8.126
R4176 out_p.n720 out_p.t1354 8.126
R4177 out_p.n720 out_p.t1547 8.126
R4178 out_p.n723 out_p.t340 8.126
R4179 out_p.n723 out_p.t801 8.126
R4180 out_p.n724 out_p.t1351 8.126
R4181 out_p.n724 out_p.t1521 8.126
R4182 out_p.n725 out_p.t403 8.126
R4183 out_p.n725 out_p.t200 8.126
R4184 out_p.n726 out_p.t156 8.126
R4185 out_p.n726 out_p.t391 8.126
R4186 out_p.n727 out_p.t472 8.126
R4187 out_p.n727 out_p.t1298 8.126
R4188 out_p.n728 out_p.t1548 8.126
R4189 out_p.n728 out_p.t766 8.126
R4190 out_p.n729 out_p.t880 8.126
R4191 out_p.n729 out_p.t1516 8.126
R4192 out_p.n730 out_p.t598 8.126
R4193 out_p.n730 out_p.t1448 8.126
R4194 out_p.n731 out_p.t396 8.126
R4195 out_p.n731 out_p.t977 8.126
R4196 out_p.n732 out_p.t1013 8.126
R4197 out_p.n732 out_p.t1582 8.126
R4198 out_p.n735 out_p.t515 8.126
R4199 out_p.n735 out_p.t976 8.126
R4200 out_p.n736 out_p.t993 8.126
R4201 out_p.n736 out_p.t1075 8.126
R4202 out_p.n737 out_p.t353 8.126
R4203 out_p.n737 out_p.t703 8.126
R4204 out_p.n738 out_p.t1610 8.126
R4205 out_p.n738 out_p.t682 8.126
R4206 out_p.n739 out_p.t1281 8.126
R4207 out_p.n739 out_p.t831 8.126
R4208 out_p.n740 out_p.t884 8.126
R4209 out_p.n740 out_p.t1435 8.126
R4210 out_p.n741 out_p.t913 8.126
R4211 out_p.n741 out_p.t404 8.126
R4212 out_p.n742 out_p.t1523 8.126
R4213 out_p.n742 out_p.t1203 8.126
R4214 out_p.n743 out_p.t1167 8.126
R4215 out_p.n743 out_p.t1550 8.126
R4216 out_p.n744 out_p.t1284 8.126
R4217 out_p.n744 out_p.t1300 8.126
R4218 out_p.n747 out_p.t907 8.126
R4219 out_p.n747 out_p.t471 8.126
R4220 out_p.n748 out_p.t1212 8.126
R4221 out_p.n748 out_p.t1653 8.126
R4222 out_p.n749 out_p.t1148 8.126
R4223 out_p.n749 out_p.t1044 8.126
R4224 out_p.n750 out_p.t821 8.126
R4225 out_p.n750 out_p.t725 8.126
R4226 out_p.n751 out_p.t1209 8.126
R4227 out_p.n751 out_p.t832 8.126
R4228 out_p.n752 out_p.t1285 8.126
R4229 out_p.n752 out_p.t351 8.126
R4230 out_p.n753 out_p.t1394 8.126
R4231 out_p.n753 out_p.t1618 8.126
R4232 out_p.n754 out_p.t1316 8.126
R4233 out_p.n754 out_p.t1015 8.126
R4234 out_p.n755 out_p.t1240 8.126
R4235 out_p.n755 out_p.t317 8.126
R4236 out_p.n756 out_p.t538 8.126
R4237 out_p.n756 out_p.t581 8.126
R4238 out_p.n759 out_p.t487 8.126
R4239 out_p.n759 out_p.t1196 8.126
R4240 out_p.n760 out_p.t1464 8.126
R4241 out_p.n760 out_p.t1400 8.126
R4242 out_p.n761 out_p.t951 8.126
R4243 out_p.n761 out_p.t1127 8.126
R4244 out_p.n762 out_p.t1476 8.126
R4245 out_p.n762 out_p.t637 8.126
R4246 out_p.n763 out_p.t699 8.126
R4247 out_p.n763 out_p.t385 8.126
R4248 out_p.n764 out_p.t539 8.126
R4249 out_p.n764 out_p.t206 8.126
R4250 out_p.n765 out_p.t483 8.126
R4251 out_p.n765 out_p.t972 8.126
R4252 out_p.n766 out_p.t279 8.126
R4253 out_p.n766 out_p.t1512 8.126
R4254 out_p.n767 out_p.t401 8.126
R4255 out_p.n767 out_p.t480 8.126
R4256 out_p.n768 out_p.t611 8.126
R4257 out_p.n768 out_p.t1319 8.126
R4258 out_p.n771 out_p.t727 8.126
R4259 out_p.n771 out_p.t742 8.126
R4260 out_p.n772 out_p.t1282 8.126
R4261 out_p.n772 out_p.t623 8.126
R4262 out_p.n773 out_p.t814 8.126
R4263 out_p.n773 out_p.t1109 8.126
R4264 out_p.n774 out_p.t1239 8.126
R4265 out_p.n774 out_p.t750 8.126
R4266 out_p.n775 out_p.t1273 8.126
R4267 out_p.n775 out_p.t1620 8.126
R4268 out_p.n776 out_p.t796 8.126
R4269 out_p.n776 out_p.t752 8.126
R4270 out_p.n777 out_p.t381 8.126
R4271 out_p.n777 out_p.t159 8.126
R4272 out_p.n778 out_p.t1559 8.126
R4273 out_p.n778 out_p.t1625 8.126
R4274 out_p.n779 out_p.t921 8.126
R4275 out_p.n779 out_p.t175 8.126
R4276 out_p.n780 out_p.t590 8.126
R4277 out_p.n780 out_p.t1333 8.126
R4278 out_p.n783 out_p.t1599 8.126
R4279 out_p.n783 out_p.t1436 8.126
R4280 out_p.n784 out_p.t822 8.126
R4281 out_p.n784 out_p.t1335 8.126
R4282 out_p.n785 out_p.t711 8.126
R4283 out_p.n785 out_p.t258 8.126
R4284 out_p.n786 out_p.t769 8.126
R4285 out_p.n786 out_p.t1463 8.126
R4286 out_p.n787 out_p.t1017 8.126
R4287 out_p.n787 out_p.t1577 8.126
R4288 out_p.n788 out_p.t591 8.126
R4289 out_p.n788 out_p.t655 8.126
R4290 out_p.n789 out_p.t1118 8.126
R4291 out_p.n789 out_p.t1077 8.126
R4292 out_p.n790 out_p.t1084 8.126
R4293 out_p.n790 out_p.t956 8.126
R4294 out_p.n791 out_p.t1564 8.126
R4295 out_p.n791 out_p.t917 8.126
R4296 out_p.n792 out_p.t1247 8.126
R4297 out_p.n792 out_p.t524 8.126
R4298 out_p.n795 out_p.t501 8.126
R4299 out_p.n795 out_p.t1021 8.126
R4300 out_p.n796 out_p.t163 8.126
R4301 out_p.n796 out_p.t194 8.126
R4302 out_p.n797 out_p.t1226 8.126
R4303 out_p.n797 out_p.t422 8.126
R4304 out_p.n798 out_p.t1210 8.126
R4305 out_p.n798 out_p.t1484 8.126
R4306 out_p.n799 out_p.t1469 8.126
R4307 out_p.n799 out_p.t177 8.126
R4308 out_p.n800 out_p.t1594 8.126
R4309 out_p.n800 out_p.t864 8.126
R4310 out_p.n801 out_p.t891 8.126
R4311 out_p.n801 out_p.t209 8.126
R4312 out_p.n802 out_p.t1297 8.126
R4313 out_p.n802 out_p.t585 8.126
R4314 out_p.n803 out_p.t552 8.126
R4315 out_p.n803 out_p.t1614 8.126
R4316 out_p.n804 out_p.t1158 8.126
R4317 out_p.n804 out_p.t1105 8.126
R4318 out_p.n807 out_p.t455 8.126
R4319 out_p.n807 out_p.t1189 8.126
R4320 out_p.n808 out_p.t417 8.126
R4321 out_p.n808 out_p.t1483 8.126
R4322 out_p.n809 out_p.t1236 8.126
R4323 out_p.n809 out_p.t1138 8.126
R4324 out_p.n810 out_p.t1020 8.126
R4325 out_p.n810 out_p.t434 8.126
R4326 out_p.n811 out_p.t894 8.126
R4327 out_p.n811 out_p.t267 8.126
R4328 out_p.n812 out_p.t632 8.126
R4329 out_p.n812 out_p.t302 8.126
R4330 out_p.n813 out_p.t442 8.126
R4331 out_p.n813 out_p.t1006 8.126
R4332 out_p.n814 out_p.t687 8.126
R4333 out_p.n814 out_p.t826 8.126
R4334 out_p.n815 out_p.t802 8.126
R4335 out_p.n815 out_p.t1388 8.126
R4336 out_p.n816 out_p.t893 8.126
R4337 out_p.n816 out_p.t157 8.126
R4338 out_p.n819 out_p.t898 8.126
R4339 out_p.n819 out_p.t280 8.126
R4340 out_p.n820 out_p.t1237 8.126
R4341 out_p.n820 out_p.t1215 8.126
R4342 out_p.n821 out_p.t924 8.126
R4343 out_p.n821 out_p.t1128 8.126
R4344 out_p.n822 out_p.t936 8.126
R4345 out_p.n822 out_p.t961 8.126
R4346 out_p.n823 out_p.t423 8.126
R4347 out_p.n823 out_p.t568 8.126
R4348 out_p.n824 out_p.t235 8.126
R4349 out_p.n824 out_p.t1343 8.126
R4350 out_p.n825 out_p.t464 8.126
R4351 out_p.n825 out_p.t1039 8.126
R4352 out_p.n826 out_p.t1637 8.126
R4353 out_p.n826 out_p.t1211 8.126
R4354 out_p.n827 out_p.t1595 8.126
R4355 out_p.n827 out_p.t348 8.126
R4356 out_p.n828 out_p.t160 8.126
R4357 out_p.n828 out_p.t755 8.126
R4358 out_p.n831 out_p.t491 8.126
R4359 out_p.n831 out_p.t210 8.126
R4360 out_p.n832 out_p.t971 8.126
R4361 out_p.n832 out_p.t1129 8.126
R4362 out_p.n833 out_p.t843 8.126
R4363 out_p.n833 out_p.t1267 8.126
R4364 out_p.n834 out_p.t612 8.126
R4365 out_p.n834 out_p.t616 8.126
R4366 out_p.n835 out_p.t1359 8.126
R4367 out_p.n835 out_p.t1533 8.126
R4368 out_p.n836 out_p.t1217 8.126
R4369 out_p.n836 out_p.t271 8.126
R4370 out_p.n837 out_p.t1222 8.126
R4371 out_p.n837 out_p.t1360 8.126
R4372 out_p.n838 out_p.t543 8.126
R4373 out_p.n838 out_p.t686 8.126
R4374 out_p.n839 out_p.t1468 8.126
R4375 out_p.n839 out_p.t1628 8.126
R4376 out_p.n840 out_p.t234 8.126
R4377 out_p.n840 out_p.t900 8.126
R4378 out_p.n843 out_p.t1419 8.126
R4379 out_p.n843 out_p.t962 8.126
R4380 out_p.n844 out_p.t665 8.126
R4381 out_p.n844 out_p.t944 8.126
R4382 out_p.n845 out_p.t1311 8.126
R4383 out_p.n845 out_p.t915 8.126
R4384 out_p.n846 out_p.t1286 8.126
R4385 out_p.n846 out_p.t1377 8.126
R4386 out_p.n847 out_p.t1179 8.126
R4387 out_p.n847 out_p.t1090 8.126
R4388 out_p.n848 out_p.t1174 8.126
R4389 out_p.n848 out_p.t1580 8.126
R4390 out_p.n849 out_p.t978 8.126
R4391 out_p.n849 out_p.t1474 8.126
R4392 out_p.n850 out_p.t617 8.126
R4393 out_p.n850 out_p.t937 8.126
R4394 out_p.n851 out_p.t967 8.126
R4395 out_p.n851 out_p.t266 8.126
R4396 out_p.n852 out_p.t1216 8.126
R4397 out_p.n852 out_p.t270 8.126
R4398 out_p.n855 out_p.t498 8.126
R4399 out_p.n855 out_p.t957 8.126
R4400 out_p.n856 out_p.t1108 8.126
R4401 out_p.n856 out_p.t856 8.126
R4402 out_p.n857 out_p.t1014 8.126
R4403 out_p.n857 out_p.t525 8.126
R4404 out_p.n858 out_p.t708 8.126
R4405 out_p.n858 out_p.t415 8.126
R4406 out_p.n859 out_p.t926 8.126
R4407 out_p.n859 out_p.t299 8.126
R4408 out_p.n860 out_p.t345 8.126
R4409 out_p.n860 out_p.t608 8.126
R4410 out_p.n861 out_p.t1617 8.126
R4411 out_p.n861 out_p.t643 8.126
R4412 out_p.n862 out_p.t1170 8.126
R4413 out_p.n862 out_p.t763 8.126
R4414 out_p.n863 out_p.t636 8.126
R4415 out_p.n863 out_p.t1182 8.126
R4416 out_p.n864 out_p.t1162 8.126
R4417 out_p.n864 out_p.t1536 8.126
R4418 out_p.n867 out_p.t1514 8.126
R4419 out_p.n867 out_p.t670 8.126
R4420 out_p.n868 out_p.t342 8.126
R4421 out_p.n868 out_p.t1646 8.126
R4422 out_p.n869 out_p.t1016 8.126
R4423 out_p.n869 out_p.t1522 8.126
R4424 out_p.n870 out_p.t838 8.126
R4425 out_p.n870 out_p.t661 8.126
R4426 out_p.n871 out_p.t1055 8.126
R4427 out_p.n871 out_p.t536 8.126
R4428 out_p.n872 out_p.t169 8.126
R4429 out_p.n872 out_p.t1579 8.126
R4430 out_p.n873 out_p.t1396 8.126
R4431 out_p.n873 out_p.t1213 8.126
R4432 out_p.n874 out_p.t503 8.126
R4433 out_p.n874 out_p.t1471 8.126
R4434 out_p.n875 out_p.t724 8.126
R4435 out_p.n875 out_p.t820 8.126
R4436 out_p.n876 out_p.t344 8.126
R4437 out_p.n876 out_p.t1417 8.126
R4438 out_p.n879 out_p.t892 8.126
R4439 out_p.n879 out_p.t929 8.126
R4440 out_p.n880 out_p.t669 8.126
R4441 out_p.n880 out_p.t466 8.126
R4442 out_p.n881 out_p.t737 8.126
R4443 out_p.n881 out_p.t1576 8.126
R4444 out_p.n882 out_p.t1133 8.126
R4445 out_p.n882 out_p.t859 8.126
R4446 out_p.n883 out_p.t757 8.126
R4447 out_p.n883 out_p.t713 8.126
R4448 out_p.n884 out_p.t1541 8.126
R4449 out_p.n884 out_p.t1255 8.126
R4450 out_p.n885 out_p.t1074 8.126
R4451 out_p.n885 out_p.t958 8.126
R4452 out_p.n886 out_p.t1249 8.126
R4453 out_p.n886 out_p.t1645 8.126
R4454 out_p.n887 out_p.t1598 8.126
R4455 out_p.n887 out_p.t1611 8.126
R4456 out_p.n888 out_p.t1293 8.126
R4457 out_p.n888 out_p.t1578 8.126
R4458 out_p.n891 out_p.t1095 8.126
R4459 out_p.n891 out_p.t754 8.126
R4460 out_p.n892 out_p.t714 8.126
R4461 out_p.n892 out_p.t172 8.126
R4462 out_p.n893 out_p.t1155 8.126
R4463 out_p.n893 out_p.t1651 8.126
R4464 out_p.n894 out_p.t290 8.126
R4465 out_p.n894 out_p.t1490 8.126
R4466 out_p.n895 out_p.t615 8.126
R4467 out_p.n895 out_p.t549 8.126
R4468 out_p.n896 out_p.t756 8.126
R4469 out_p.n896 out_p.t476 8.126
R4470 out_p.n897 out_p.t1328 8.126
R4471 out_p.n897 out_p.t1305 8.126
R4472 out_p.n898 out_p.t867 8.126
R4473 out_p.n898 out_p.t1313 8.126
R4474 out_p.n899 out_p.t1173 8.126
R4475 out_p.n899 out_p.t792 8.126
R4476 out_p.n900 out_p.t1540 8.126
R4477 out_p.n900 out_p.t1085 8.126
R4478 out_p.n903 out_p.t257 8.126
R4479 out_p.n903 out_p.t813 8.126
R4480 out_p.n904 out_p.t306 8.126
R4481 out_p.n904 out_p.t1288 8.126
R4482 out_p.n905 out_p.t445 8.126
R4483 out_p.n905 out_p.t277 8.126
R4484 out_p.n906 out_p.t1399 8.126
R4485 out_p.n906 out_p.t1185 8.126
R4486 out_p.n907 out_p.t252 8.126
R4487 out_p.n907 out_p.t1456 8.126
R4488 out_p.n908 out_p.t1607 8.126
R4489 out_p.n908 out_p.t548 8.126
R4490 out_p.n909 out_p.t1636 8.126
R4491 out_p.n909 out_p.t1415 8.126
R4492 out_p.n910 out_p.t730 8.126
R4493 out_p.n910 out_p.t1028 8.126
R4494 out_p.n911 out_p.t1365 8.126
R4495 out_p.n911 out_p.t795 8.126
R4496 out_p.n912 out_p.t671 8.126
R4497 out_p.n912 out_p.t499 8.126
R4498 out_p.n902 out_p.t1736 4.95
R4499 out_p.n902 out_p.t1702 4.95
R4500 out_p.n901 out_p.t79 4.95
R4501 out_p.n901 out_p.t18 4.95
R4502 out_p.n889 out_p.t1700 4.95
R4503 out_p.n889 out_p.t51 4.95
R4504 out_p.n890 out_p.t26 4.95
R4505 out_p.n890 out_p.t120 4.95
R4506 out_p.n877 out_p.t1746 4.95
R4507 out_p.n877 out_p.t30 4.95
R4508 out_p.n878 out_p.t140 4.95
R4509 out_p.n878 out_p.t1693 4.95
R4510 out_p.n865 out_p.t9 4.95
R4511 out_p.n865 out_p.t14 4.95
R4512 out_p.n866 out_p.t152 4.95
R4513 out_p.n866 out_p.t124 4.95
R4514 out_p.n853 out_p.t1790 4.95
R4515 out_p.n853 out_p.t112 4.95
R4516 out_p.n854 out_p.t1742 4.95
R4517 out_p.n854 out_p.t71 4.95
R4518 out_p.n841 out_p.t1738 4.95
R4519 out_p.n841 out_p.t1776 4.95
R4520 out_p.n842 out_p.t1661 4.95
R4521 out_p.n842 out_p.t1688 4.95
R4522 out_p.n829 out_p.t109 4.95
R4523 out_p.n829 out_p.t1767 4.95
R4524 out_p.n830 out_p.t123 4.95
R4525 out_p.n830 out_p.t48 4.95
R4526 out_p.n817 out_p.t1683 4.95
R4527 out_p.n817 out_p.t108 4.95
R4528 out_p.n818 out_p.t1706 4.95
R4529 out_p.n818 out_p.t122 4.95
R4530 out_p.n805 out_p.t1766 4.95
R4531 out_p.n805 out_p.t1682 4.95
R4532 out_p.n806 out_p.t1745 4.95
R4533 out_p.n806 out_p.t1711 4.95
R4534 out_p.n793 out_p.t1721 4.95
R4535 out_p.n793 out_p.t1734 4.95
R4536 out_p.n794 out_p.t83 4.95
R4537 out_p.n794 out_p.t1733 4.95
R4538 out_p.n781 out_p.t69 4.95
R4539 out_p.n781 out_p.t1713 4.95
R4540 out_p.n782 out_p.t1722 4.95
R4541 out_p.n782 out_p.t155 4.95
R4542 out_p.n769 out_p.t1759 4.95
R4543 out_p.n769 out_p.t77 4.95
R4544 out_p.n770 out_p.t89 4.95
R4545 out_p.n770 out_p.t1781 4.95
R4546 out_p.n757 out_p.t53 4.95
R4547 out_p.n757 out_p.t114 4.95
R4548 out_p.n758 out_p.t1762 4.95
R4549 out_p.n758 out_p.t1770 4.95
R4550 out_p.n745 out_p.t1671 4.95
R4551 out_p.n745 out_p.t1658 4.95
R4552 out_p.n746 out_p.t1775 4.95
R4553 out_p.n746 out_p.t1719 4.95
R4554 out_p.n733 out_p.t1783 4.95
R4555 out_p.n733 out_p.t1679 4.95
R4556 out_p.n734 out_p.t102 4.95
R4557 out_p.n734 out_p.t1669 4.95
R4558 out_p.n721 out_p.t1797 4.95
R4559 out_p.n721 out_p.t116 4.95
R4560 out_p.n722 out_p.t1788 4.95
R4561 out_p.n722 out_p.t46 4.95
R4562 out_p.n709 out_p.t42 4.95
R4563 out_p.n709 out_p.t98 4.95
R4564 out_p.n710 out_p.t6 4.95
R4565 out_p.n710 out_p.t96 4.95
R4566 out_p.n697 out_p.t95 4.95
R4567 out_p.n697 out_p.t22 4.95
R4568 out_p.n698 out_p.t33 4.95
R4569 out_p.n698 out_p.t106 4.95
R4570 out_p.n685 out_p.t1664 4.95
R4571 out_p.n685 out_p.t58 4.95
R4572 out_p.n686 out_p.t1754 4.95
R4573 out_p.n686 out_p.t80 4.95
R4574 out_p.n673 out_p.t1716 4.95
R4575 out_p.n673 out_p.t1677 4.95
R4576 out_p.n674 out_p.t40 4.95
R4577 out_p.n674 out_p.t99 4.95
R4578 out_p.n661 out_p.t57 4.95
R4579 out_p.n661 out_p.t118 4.95
R4580 out_p.n662 out_p.t111 4.95
R4581 out_p.n662 out_p.t1672 4.95
R4582 out_p.n649 out_p.t1726 4.95
R4583 out_p.n649 out_p.t1750 4.95
R4584 out_p.n650 out_p.t1779 4.95
R4585 out_p.n650 out_p.t73 4.95
R4586 out_p.n637 out_p.t1799 4.95
R4587 out_p.n637 out_p.t1769 4.95
R4588 out_p.n638 out_p.t1681 4.95
R4589 out_p.n638 out_p.t62 4.95
R4590 out_p.n625 out_p.t1796 4.95
R4591 out_p.n625 out_p.t1731 4.95
R4592 out_p.n626 out_p.t101 4.95
R4593 out_p.n626 out_p.t1725 4.95
R4594 out_p.n613 out_p.t0 4.95
R4595 out_p.n613 out_p.t75 4.95
R4596 out_p.n614 out_p.t1662 4.95
R4597 out_p.n614 out_p.t1709 4.95
R4598 out_p.n601 out_p.t1753 4.95
R4599 out_p.n601 out_p.t66 4.95
R4600 out_p.n602 out_p.t1748 4.95
R4601 out_p.n602 out_p.t1696 4.95
R4602 out_p.n589 out_p.t52 4.95
R4603 out_p.n589 out_p.t134 4.95
R4604 out_p.n590 out_p.t1747 4.95
R4605 out_p.n590 out_p.t1761 4.95
R4606 out_p.n577 out_p.t44 4.95
R4607 out_p.n577 out_p.t144 4.95
R4608 out_p.n578 out_p.t1676 4.95
R4609 out_p.n578 out_p.t59 4.95
R4610 out_p.n565 out_p.t56 4.95
R4611 out_p.n565 out_p.t1678 4.95
R4612 out_p.n566 out_p.t110 4.95
R4613 out_p.n566 out_p.t1668 4.95
R4614 out_p.n553 out_p.t1739 4.95
R4615 out_p.n553 out_p.t1757 4.95
R4616 out_p.n554 out_p.t1732 4.95
R4617 out_p.n554 out_p.t72 4.95
R4618 out_p.n541 out_p.t1 4.95
R4619 out_p.n541 out_p.t16 4.95
R4620 out_p.n542 out_p.t1663 4.95
R4621 out_p.n542 out_p.t1674 4.95
R4622 out_p.n529 out_p.t12 4.95
R4623 out_p.n529 out_p.t31 4.95
R4624 out_p.n530 out_p.t153 4.95
R4625 out_p.n530 out_p.t1694 4.95
R4626 out_p.n517 out_p.t126 4.95
R4627 out_p.n517 out_p.t1737 4.95
R4628 out_p.n518 out_p.t1657 4.95
R4629 out_p.n518 out_p.t117 4.95
R4630 out_p.n505 out_p.t1752 4.95
R4631 out_p.n505 out_p.t78 4.95
R4632 out_p.n506 out_p.t43 4.95
R4633 out_p.n506 out_p.t1741 4.95
R4634 out_p.n493 out_p.t130 4.95
R4635 out_p.n493 out_p.t1689 4.95
R4636 out_p.n494 out_p.t23 4.95
R4637 out_p.n494 out_p.t1665 4.95
R4638 out_p.n481 out_p.t1756 4.95
R4639 out_p.n481 out_p.t1798 4.95
R4640 out_p.n482 out_p.t115 4.95
R4641 out_p.n482 out_p.t1680 4.95
R4642 out_p.n469 out_p.t64 4.95
R4643 out_p.n469 out_p.t132 4.95
R4644 out_p.n470 out_p.t92 4.95
R4645 out_p.n470 out_p.t105 4.95
R4646 out_p.n457 out_p.t4 4.95
R4647 out_p.n457 out_p.t1695 4.95
R4648 out_p.n458 out_p.t119 4.95
R4649 out_p.n458 out_p.t1727 4.95
R4650 out_p.n445 out_p.t74 4.95
R4651 out_p.n445 out_p.t8 4.95
R4652 out_p.n446 out_p.t1708 4.95
R4653 out_p.n446 out_p.t1795 4.95
R4654 out_p.n433 out_p.t38 4.95
R4655 out_p.n433 out_p.t1703 4.95
R4656 out_p.n434 out_p.t1691 4.95
R4657 out_p.n434 out_p.t1656 4.95
R4658 out_p.n421 out_p.t131 4.95
R4659 out_p.n421 out_p.t147 4.95
R4660 out_p.n422 out_p.t1760 4.95
R4661 out_p.n422 out_p.t1710 4.95
R4662 out_p.n409 out_p.t1787 4.95
R4663 out_p.n409 out_p.t129 4.95
R4664 out_p.n410 out_p.t1744 4.95
R4665 out_p.n410 out_p.t37 4.95
R4666 out_p.n397 out_p.t61 4.95
R4667 out_p.n397 out_p.t93 4.95
R4668 out_p.n398 out_p.t67 4.95
R4669 out_p.n398 out_p.t1660 4.95
R4670 out_p.n385 out_p.t1685 4.95
R4671 out_p.n385 out_p.t1704 4.95
R4672 out_p.n386 out_p.t139 4.95
R4673 out_p.n386 out_p.t60 4.95
R4674 out_p.n373 out_p.t1743 4.95
R4675 out_p.n373 out_p.t125 4.95
R4676 out_p.n374 out_p.t145 4.95
R4677 out_p.n374 out_p.t104 4.95
R4678 out_p.n361 out_p.t39 4.95
R4679 out_p.n361 out_p.t1793 4.95
R4680 out_p.n362 out_p.t1692 4.95
R4681 out_p.n362 out_p.t137 4.95
R4682 out_p.n349 out_p.t50 4.95
R4683 out_p.n349 out_p.t87 4.95
R4684 out_p.n350 out_p.t11 4.95
R4685 out_p.n350 out_p.t3 4.95
R4686 out_p.n337 out_p.t1707 4.95
R4687 out_p.n337 out_p.t49 4.95
R4688 out_p.n338 out_p.t17 4.95
R4689 out_p.n338 out_p.t1740 4.95
R4690 out_p.n325 out_p.t1667 4.95
R4691 out_p.n325 out_p.t1715 4.95
R4692 out_p.n326 out_p.t25 4.95
R4693 out_p.n326 out_p.t142 4.95
R4694 out_p.n313 out_p.t103 4.95
R4695 out_p.n313 out_p.t128 4.95
R4696 out_p.n314 out_p.t150 4.95
R4697 out_p.n314 out_p.t36 4.95
R4698 out_p.n301 out_p.t35 4.95
R4699 out_p.n301 out_p.t68 4.95
R4700 out_p.n302 out_p.t1784 4.95
R4701 out_p.n302 out_p.t85 4.95
R4702 out_p.n289 out_p.t7 4.95
R4703 out_p.n289 out_p.t97 4.95
R4704 out_p.n290 out_p.t1777 4.95
R4705 out_p.n290 out_p.t1735 4.95
R4706 out_p.n277 out_p.t141 4.95
R4707 out_p.n277 out_p.t1772 4.95
R4708 out_p.n278 out_p.t1751 4.95
R4709 out_p.n278 out_p.t1698 4.95
R4710 out_p.n265 out_p.t20 4.95
R4711 out_p.n265 out_p.t81 4.95
R4712 out_p.n266 out_p.t90 4.95
R4713 out_p.n266 out_p.t133 4.95
R4714 out_p.n253 out_p.t148 4.95
R4715 out_p.n253 out_p.t86 4.95
R4716 out_p.n254 out_p.t5 4.95
R4717 out_p.n254 out_p.t2 4.95
R4718 out_p.n241 out_p.t1687 4.95
R4719 out_p.n241 out_p.t1673 4.95
R4720 out_p.n242 out_p.t55 4.95
R4721 out_p.n242 out_p.t1701 4.95
R4722 out_p.n229 out_p.t1764 4.95
R4723 out_p.n229 out_p.t1785 4.95
R4724 out_p.n230 out_p.t19 4.95
R4725 out_p.n230 out_p.t1728 4.95
R4726 out_p.n217 out_p.t1723 4.95
R4727 out_p.n217 out_p.t1712 4.95
R4728 out_p.n218 out_p.t135 4.95
R4729 out_p.n218 out_p.t154 4.95
R4730 out_p.n205 out_p.t1758 4.95
R4731 out_p.n205 out_p.t76 4.95
R4732 out_p.n206 out_p.t88 4.95
R4733 out_p.n206 out_p.t1780 4.95
R4734 out_p.n193 out_p.t121 4.95
R4735 out_p.n193 out_p.t27 4.95
R4736 out_p.n194 out_p.t1794 4.95
R4737 out_p.n194 out_p.t1690 4.95
R4738 out_p.n181 out_p.t1717 4.95
R4739 out_p.n181 out_p.t1720 4.95
R4740 out_p.n182 out_p.t41 4.95
R4741 out_p.n182 out_p.t82 4.95
R4742 out_p.n179 out_p.t146 4.95
R4743 out_p.n179 out_p.t1786 4.95
R4744 out_p.n180 out_p.t143 4.95
R4745 out_p.n180 out_p.t151 4.95
R4746 out_p.n10 out_p.t1670 4.95
R4747 out_p.n10 out_p.t1765 4.95
R4748 out_p.n11 out_p.t1774 4.95
R4749 out_p.n11 out_p.t1718 4.95
R4750 out_p.n12 out_p.t1782 4.95
R4751 out_p.n12 out_p.t1684 4.95
R4752 out_p.n13 out_p.t1729 4.95
R4753 out_p.n13 out_p.t138 4.95
R4754 out_p.n14 out_p.t70 4.95
R4755 out_p.n14 out_p.t1789 4.95
R4756 out_p.n15 out_p.t45 4.95
R4757 out_p.n15 out_p.t29 4.95
R4758 out_p.n16 out_p.t1773 4.95
R4759 out_p.n16 out_p.t21 4.95
R4760 out_p.n17 out_p.t1699 4.95
R4761 out_p.n17 out_p.t91 4.95
R4762 out_p.n18 out_p.t1792 4.95
R4763 out_p.n18 out_p.t149 4.95
R4764 out_p.n19 out_p.t136 4.95
R4765 out_p.n19 out_p.t10 4.95
R4766 out_p.n20 out_p.t1697 4.95
R4767 out_p.n20 out_p.t1763 4.95
R4768 out_p.n21 out_p.t1791 4.95
R4769 out_p.n21 out_p.t15 4.95
R4770 out_p.n22 out_p.t1771 4.95
R4771 out_p.n22 out_p.t1666 4.95
R4772 out_p.n23 out_p.t13 4.95
R4773 out_p.n23 out_p.t24 4.95
R4774 out_p.n24 out_p.t1714 4.95
R4775 out_p.n24 out_p.t1686 4.95
R4776 out_p.n25 out_p.t127 4.95
R4777 out_p.n25 out_p.t54 4.95
R4778 out_p.n26 out_p.t63 4.95
R4779 out_p.n26 out_p.t34 4.95
R4780 out_p.n27 out_p.t1778 4.95
R4781 out_p.n27 out_p.t28 4.95
R4782 out_p.n28 out_p.t47 4.95
R4783 out_p.n28 out_p.t1768 4.95
R4784 out_p.n29 out_p.t84 4.95
R4785 out_p.n29 out_p.t1659 4.95
R4786 out_p.n30 out_p.t1675 4.95
R4787 out_p.n30 out_p.t1730 4.95
R4788 out_p.n31 out_p.t100 4.95
R4789 out_p.n31 out_p.t1724 4.95
R4790 out_p.n32 out_p.t107 4.95
R4791 out_p.n32 out_p.t1755 4.95
R4792 out_p.n33 out_p.t1705 4.95
R4793 out_p.n33 out_p.t65 4.95
R4794 out_p.n34 out_p.t94 4.95
R4795 out_p.n34 out_p.t1749 4.95
R4796 out_p.n35 out_p.t32 4.95
R4797 out_p.n35 out_p.t113 4.95
R4798 out_p.n908 out_p.n907 0.866
R4799 out_p.n41 out_p.n40 0.85
R4800 out_p.n52 out_p.n51 0.85
R4801 out_p.n63 out_p.n62 0.85
R4802 out_p.n74 out_p.n73 0.85
R4803 out_p.n85 out_p.n84 0.85
R4804 out_p.n96 out_p.n95 0.85
R4805 out_p.n107 out_p.n106 0.85
R4806 out_p.n118 out_p.n117 0.85
R4807 out_p.n129 out_p.n128 0.85
R4808 out_p.n140 out_p.n139 0.85
R4809 out_p.n151 out_p.n150 0.85
R4810 out_p.n162 out_p.n161 0.85
R4811 out_p.n173 out_p.n172 0.85
R4812 out_p.n5 out_p.n4 0.85
R4813 out_p.n188 out_p.n187 0.85
R4814 out_p.n200 out_p.n199 0.85
R4815 out_p.n212 out_p.n211 0.85
R4816 out_p.n224 out_p.n223 0.85
R4817 out_p.n236 out_p.n235 0.85
R4818 out_p.n248 out_p.n247 0.85
R4819 out_p.n260 out_p.n259 0.85
R4820 out_p.n272 out_p.n271 0.85
R4821 out_p.n284 out_p.n283 0.85
R4822 out_p.n296 out_p.n295 0.85
R4823 out_p.n308 out_p.n307 0.85
R4824 out_p.n320 out_p.n319 0.85
R4825 out_p.n332 out_p.n331 0.85
R4826 out_p.n344 out_p.n343 0.85
R4827 out_p.n356 out_p.n355 0.85
R4828 out_p.n368 out_p.n367 0.85
R4829 out_p.n380 out_p.n379 0.85
R4830 out_p.n392 out_p.n391 0.85
R4831 out_p.n404 out_p.n403 0.85
R4832 out_p.n416 out_p.n415 0.85
R4833 out_p.n428 out_p.n427 0.85
R4834 out_p.n440 out_p.n439 0.85
R4835 out_p.n452 out_p.n451 0.85
R4836 out_p.n464 out_p.n463 0.85
R4837 out_p.n476 out_p.n475 0.85
R4838 out_p.n488 out_p.n487 0.85
R4839 out_p.n500 out_p.n499 0.85
R4840 out_p.n512 out_p.n511 0.85
R4841 out_p.n524 out_p.n523 0.85
R4842 out_p.n536 out_p.n535 0.85
R4843 out_p.n548 out_p.n547 0.85
R4844 out_p.n560 out_p.n559 0.85
R4845 out_p.n572 out_p.n571 0.85
R4846 out_p.n584 out_p.n583 0.85
R4847 out_p.n596 out_p.n595 0.85
R4848 out_p.n608 out_p.n607 0.85
R4849 out_p.n620 out_p.n619 0.85
R4850 out_p.n632 out_p.n631 0.85
R4851 out_p.n644 out_p.n643 0.85
R4852 out_p.n656 out_p.n655 0.85
R4853 out_p.n668 out_p.n667 0.85
R4854 out_p.n680 out_p.n679 0.85
R4855 out_p.n692 out_p.n691 0.85
R4856 out_p.n704 out_p.n703 0.85
R4857 out_p.n716 out_p.n715 0.85
R4858 out_p.n728 out_p.n727 0.85
R4859 out_p.n740 out_p.n739 0.85
R4860 out_p.n752 out_p.n751 0.85
R4861 out_p.n764 out_p.n763 0.85
R4862 out_p.n776 out_p.n775 0.85
R4863 out_p.n788 out_p.n787 0.85
R4864 out_p.n800 out_p.n799 0.85
R4865 out_p.n812 out_p.n811 0.85
R4866 out_p.n824 out_p.n823 0.85
R4867 out_p.n836 out_p.n835 0.85
R4868 out_p.n848 out_p.n847 0.85
R4869 out_p.n860 out_p.n859 0.85
R4870 out_p.n872 out_p.n871 0.85
R4871 out_p.n884 out_p.n883 0.85
R4872 out_p.n896 out_p.n895 0.85
R4873 out_p.n912 out_p.n911 0.77
R4874 out_p.n911 out_p.n910 0.77
R4875 out_p.n910 out_p.n909 0.77
R4876 out_p.n909 out_p.n908 0.77
R4877 out_p.n907 out_p.n906 0.77
R4878 out_p.n906 out_p.n905 0.77
R4879 out_p.n905 out_p.n904 0.77
R4880 out_p.n904 out_p.n903 0.77
R4881 out_p.n902 out_p.n901 0.76
R4882 out_p.n890 out_p.n889 0.76
R4883 out_p.n878 out_p.n877 0.76
R4884 out_p.n866 out_p.n865 0.76
R4885 out_p.n854 out_p.n853 0.76
R4886 out_p.n842 out_p.n841 0.76
R4887 out_p.n830 out_p.n829 0.76
R4888 out_p.n818 out_p.n817 0.76
R4889 out_p.n806 out_p.n805 0.76
R4890 out_p.n794 out_p.n793 0.76
R4891 out_p.n782 out_p.n781 0.76
R4892 out_p.n770 out_p.n769 0.76
R4893 out_p.n758 out_p.n757 0.76
R4894 out_p.n746 out_p.n745 0.76
R4895 out_p.n734 out_p.n733 0.76
R4896 out_p.n722 out_p.n721 0.76
R4897 out_p.n710 out_p.n709 0.76
R4898 out_p.n698 out_p.n697 0.76
R4899 out_p.n686 out_p.n685 0.76
R4900 out_p.n674 out_p.n673 0.76
R4901 out_p.n662 out_p.n661 0.76
R4902 out_p.n650 out_p.n649 0.76
R4903 out_p.n638 out_p.n637 0.76
R4904 out_p.n626 out_p.n625 0.76
R4905 out_p.n614 out_p.n613 0.76
R4906 out_p.n602 out_p.n601 0.76
R4907 out_p.n590 out_p.n589 0.76
R4908 out_p.n578 out_p.n577 0.76
R4909 out_p.n566 out_p.n565 0.76
R4910 out_p.n554 out_p.n553 0.76
R4911 out_p.n542 out_p.n541 0.76
R4912 out_p.n530 out_p.n529 0.76
R4913 out_p.n518 out_p.n517 0.76
R4914 out_p.n506 out_p.n505 0.76
R4915 out_p.n494 out_p.n493 0.76
R4916 out_p.n482 out_p.n481 0.76
R4917 out_p.n470 out_p.n469 0.76
R4918 out_p.n458 out_p.n457 0.76
R4919 out_p.n446 out_p.n445 0.76
R4920 out_p.n434 out_p.n433 0.76
R4921 out_p.n422 out_p.n421 0.76
R4922 out_p.n410 out_p.n409 0.76
R4923 out_p.n398 out_p.n397 0.76
R4924 out_p.n386 out_p.n385 0.76
R4925 out_p.n374 out_p.n373 0.76
R4926 out_p.n362 out_p.n361 0.76
R4927 out_p.n350 out_p.n349 0.76
R4928 out_p.n338 out_p.n337 0.76
R4929 out_p.n326 out_p.n325 0.76
R4930 out_p.n314 out_p.n313 0.76
R4931 out_p.n302 out_p.n301 0.76
R4932 out_p.n290 out_p.n289 0.76
R4933 out_p.n278 out_p.n277 0.76
R4934 out_p.n266 out_p.n265 0.76
R4935 out_p.n254 out_p.n253 0.76
R4936 out_p.n242 out_p.n241 0.76
R4937 out_p.n230 out_p.n229 0.76
R4938 out_p.n218 out_p.n217 0.76
R4939 out_p.n206 out_p.n205 0.76
R4940 out_p.n194 out_p.n193 0.76
R4941 out_p.n182 out_p.n181 0.76
R4942 out_p.n180 out_p.n179 0.76
R4943 out_p.n11 out_p.n10 0.76
R4944 out_p.n13 out_p.n12 0.76
R4945 out_p.n15 out_p.n14 0.76
R4946 out_p.n17 out_p.n16 0.76
R4947 out_p.n19 out_p.n18 0.76
R4948 out_p.n21 out_p.n20 0.76
R4949 out_p.n23 out_p.n22 0.76
R4950 out_p.n25 out_p.n24 0.76
R4951 out_p.n27 out_p.n26 0.76
R4952 out_p.n29 out_p.n28 0.76
R4953 out_p.n31 out_p.n30 0.76
R4954 out_p.n33 out_p.n32 0.76
R4955 out_p.n35 out_p.n34 0.76
R4956 out_p.n45 out_p.n44 0.754
R4957 out_p.n44 out_p.n43 0.754
R4958 out_p.n43 out_p.n42 0.754
R4959 out_p.n42 out_p.n41 0.754
R4960 out_p.n40 out_p.n39 0.754
R4961 out_p.n39 out_p.n38 0.754
R4962 out_p.n38 out_p.n37 0.754
R4963 out_p.n37 out_p.n36 0.754
R4964 out_p.n56 out_p.n55 0.754
R4965 out_p.n55 out_p.n54 0.754
R4966 out_p.n54 out_p.n53 0.754
R4967 out_p.n53 out_p.n52 0.754
R4968 out_p.n51 out_p.n50 0.754
R4969 out_p.n50 out_p.n49 0.754
R4970 out_p.n49 out_p.n48 0.754
R4971 out_p.n48 out_p.n47 0.754
R4972 out_p.n67 out_p.n66 0.754
R4973 out_p.n66 out_p.n65 0.754
R4974 out_p.n65 out_p.n64 0.754
R4975 out_p.n64 out_p.n63 0.754
R4976 out_p.n62 out_p.n61 0.754
R4977 out_p.n61 out_p.n60 0.754
R4978 out_p.n60 out_p.n59 0.754
R4979 out_p.n59 out_p.n58 0.754
R4980 out_p.n78 out_p.n77 0.754
R4981 out_p.n77 out_p.n76 0.754
R4982 out_p.n76 out_p.n75 0.754
R4983 out_p.n75 out_p.n74 0.754
R4984 out_p.n73 out_p.n72 0.754
R4985 out_p.n72 out_p.n71 0.754
R4986 out_p.n71 out_p.n70 0.754
R4987 out_p.n70 out_p.n69 0.754
R4988 out_p.n89 out_p.n88 0.754
R4989 out_p.n88 out_p.n87 0.754
R4990 out_p.n87 out_p.n86 0.754
R4991 out_p.n86 out_p.n85 0.754
R4992 out_p.n84 out_p.n83 0.754
R4993 out_p.n83 out_p.n82 0.754
R4994 out_p.n82 out_p.n81 0.754
R4995 out_p.n81 out_p.n80 0.754
R4996 out_p.n100 out_p.n99 0.754
R4997 out_p.n99 out_p.n98 0.754
R4998 out_p.n98 out_p.n97 0.754
R4999 out_p.n97 out_p.n96 0.754
R5000 out_p.n95 out_p.n94 0.754
R5001 out_p.n94 out_p.n93 0.754
R5002 out_p.n93 out_p.n92 0.754
R5003 out_p.n92 out_p.n91 0.754
R5004 out_p.n111 out_p.n110 0.754
R5005 out_p.n110 out_p.n109 0.754
R5006 out_p.n109 out_p.n108 0.754
R5007 out_p.n108 out_p.n107 0.754
R5008 out_p.n106 out_p.n105 0.754
R5009 out_p.n105 out_p.n104 0.754
R5010 out_p.n104 out_p.n103 0.754
R5011 out_p.n103 out_p.n102 0.754
R5012 out_p.n122 out_p.n121 0.754
R5013 out_p.n121 out_p.n120 0.754
R5014 out_p.n120 out_p.n119 0.754
R5015 out_p.n119 out_p.n118 0.754
R5016 out_p.n117 out_p.n116 0.754
R5017 out_p.n116 out_p.n115 0.754
R5018 out_p.n115 out_p.n114 0.754
R5019 out_p.n114 out_p.n113 0.754
R5020 out_p.n133 out_p.n132 0.754
R5021 out_p.n132 out_p.n131 0.754
R5022 out_p.n131 out_p.n130 0.754
R5023 out_p.n130 out_p.n129 0.754
R5024 out_p.n128 out_p.n127 0.754
R5025 out_p.n127 out_p.n126 0.754
R5026 out_p.n126 out_p.n125 0.754
R5027 out_p.n125 out_p.n124 0.754
R5028 out_p.n144 out_p.n143 0.754
R5029 out_p.n143 out_p.n142 0.754
R5030 out_p.n142 out_p.n141 0.754
R5031 out_p.n141 out_p.n140 0.754
R5032 out_p.n139 out_p.n138 0.754
R5033 out_p.n138 out_p.n137 0.754
R5034 out_p.n137 out_p.n136 0.754
R5035 out_p.n136 out_p.n135 0.754
R5036 out_p.n155 out_p.n154 0.754
R5037 out_p.n154 out_p.n153 0.754
R5038 out_p.n153 out_p.n152 0.754
R5039 out_p.n152 out_p.n151 0.754
R5040 out_p.n150 out_p.n149 0.754
R5041 out_p.n149 out_p.n148 0.754
R5042 out_p.n148 out_p.n147 0.754
R5043 out_p.n147 out_p.n146 0.754
R5044 out_p.n166 out_p.n165 0.754
R5045 out_p.n165 out_p.n164 0.754
R5046 out_p.n164 out_p.n163 0.754
R5047 out_p.n163 out_p.n162 0.754
R5048 out_p.n161 out_p.n160 0.754
R5049 out_p.n160 out_p.n159 0.754
R5050 out_p.n159 out_p.n158 0.754
R5051 out_p.n158 out_p.n157 0.754
R5052 out_p.n177 out_p.n176 0.754
R5053 out_p.n176 out_p.n175 0.754
R5054 out_p.n175 out_p.n174 0.754
R5055 out_p.n174 out_p.n173 0.754
R5056 out_p.n172 out_p.n171 0.754
R5057 out_p.n171 out_p.n170 0.754
R5058 out_p.n170 out_p.n169 0.754
R5059 out_p.n169 out_p.n168 0.754
R5060 out_p.n9 out_p.n8 0.754
R5061 out_p.n8 out_p.n7 0.754
R5062 out_p.n7 out_p.n6 0.754
R5063 out_p.n6 out_p.n5 0.754
R5064 out_p.n4 out_p.n3 0.754
R5065 out_p.n3 out_p.n2 0.754
R5066 out_p.n2 out_p.n1 0.754
R5067 out_p.n1 out_p.n0 0.754
R5068 out_p.n192 out_p.n191 0.754
R5069 out_p.n191 out_p.n190 0.754
R5070 out_p.n190 out_p.n189 0.754
R5071 out_p.n189 out_p.n188 0.754
R5072 out_p.n187 out_p.n186 0.754
R5073 out_p.n186 out_p.n185 0.754
R5074 out_p.n185 out_p.n184 0.754
R5075 out_p.n184 out_p.n183 0.754
R5076 out_p.n204 out_p.n203 0.754
R5077 out_p.n203 out_p.n202 0.754
R5078 out_p.n202 out_p.n201 0.754
R5079 out_p.n201 out_p.n200 0.754
R5080 out_p.n199 out_p.n198 0.754
R5081 out_p.n198 out_p.n197 0.754
R5082 out_p.n197 out_p.n196 0.754
R5083 out_p.n196 out_p.n195 0.754
R5084 out_p.n216 out_p.n215 0.754
R5085 out_p.n215 out_p.n214 0.754
R5086 out_p.n214 out_p.n213 0.754
R5087 out_p.n213 out_p.n212 0.754
R5088 out_p.n211 out_p.n210 0.754
R5089 out_p.n210 out_p.n209 0.754
R5090 out_p.n209 out_p.n208 0.754
R5091 out_p.n208 out_p.n207 0.754
R5092 out_p.n228 out_p.n227 0.754
R5093 out_p.n227 out_p.n226 0.754
R5094 out_p.n226 out_p.n225 0.754
R5095 out_p.n225 out_p.n224 0.754
R5096 out_p.n223 out_p.n222 0.754
R5097 out_p.n222 out_p.n221 0.754
R5098 out_p.n221 out_p.n220 0.754
R5099 out_p.n220 out_p.n219 0.754
R5100 out_p.n240 out_p.n239 0.754
R5101 out_p.n239 out_p.n238 0.754
R5102 out_p.n238 out_p.n237 0.754
R5103 out_p.n237 out_p.n236 0.754
R5104 out_p.n235 out_p.n234 0.754
R5105 out_p.n234 out_p.n233 0.754
R5106 out_p.n233 out_p.n232 0.754
R5107 out_p.n232 out_p.n231 0.754
R5108 out_p.n252 out_p.n251 0.754
R5109 out_p.n251 out_p.n250 0.754
R5110 out_p.n250 out_p.n249 0.754
R5111 out_p.n249 out_p.n248 0.754
R5112 out_p.n247 out_p.n246 0.754
R5113 out_p.n246 out_p.n245 0.754
R5114 out_p.n245 out_p.n244 0.754
R5115 out_p.n244 out_p.n243 0.754
R5116 out_p.n264 out_p.n263 0.754
R5117 out_p.n263 out_p.n262 0.754
R5118 out_p.n262 out_p.n261 0.754
R5119 out_p.n261 out_p.n260 0.754
R5120 out_p.n259 out_p.n258 0.754
R5121 out_p.n258 out_p.n257 0.754
R5122 out_p.n257 out_p.n256 0.754
R5123 out_p.n256 out_p.n255 0.754
R5124 out_p.n276 out_p.n275 0.754
R5125 out_p.n275 out_p.n274 0.754
R5126 out_p.n274 out_p.n273 0.754
R5127 out_p.n273 out_p.n272 0.754
R5128 out_p.n271 out_p.n270 0.754
R5129 out_p.n270 out_p.n269 0.754
R5130 out_p.n269 out_p.n268 0.754
R5131 out_p.n268 out_p.n267 0.754
R5132 out_p.n288 out_p.n287 0.754
R5133 out_p.n287 out_p.n286 0.754
R5134 out_p.n286 out_p.n285 0.754
R5135 out_p.n285 out_p.n284 0.754
R5136 out_p.n283 out_p.n282 0.754
R5137 out_p.n282 out_p.n281 0.754
R5138 out_p.n281 out_p.n280 0.754
R5139 out_p.n280 out_p.n279 0.754
R5140 out_p.n300 out_p.n299 0.754
R5141 out_p.n299 out_p.n298 0.754
R5142 out_p.n298 out_p.n297 0.754
R5143 out_p.n297 out_p.n296 0.754
R5144 out_p.n295 out_p.n294 0.754
R5145 out_p.n294 out_p.n293 0.754
R5146 out_p.n293 out_p.n292 0.754
R5147 out_p.n292 out_p.n291 0.754
R5148 out_p.n312 out_p.n311 0.754
R5149 out_p.n311 out_p.n310 0.754
R5150 out_p.n310 out_p.n309 0.754
R5151 out_p.n309 out_p.n308 0.754
R5152 out_p.n307 out_p.n306 0.754
R5153 out_p.n306 out_p.n305 0.754
R5154 out_p.n305 out_p.n304 0.754
R5155 out_p.n304 out_p.n303 0.754
R5156 out_p.n324 out_p.n323 0.754
R5157 out_p.n323 out_p.n322 0.754
R5158 out_p.n322 out_p.n321 0.754
R5159 out_p.n321 out_p.n320 0.754
R5160 out_p.n319 out_p.n318 0.754
R5161 out_p.n318 out_p.n317 0.754
R5162 out_p.n317 out_p.n316 0.754
R5163 out_p.n316 out_p.n315 0.754
R5164 out_p.n336 out_p.n335 0.754
R5165 out_p.n335 out_p.n334 0.754
R5166 out_p.n334 out_p.n333 0.754
R5167 out_p.n333 out_p.n332 0.754
R5168 out_p.n331 out_p.n330 0.754
R5169 out_p.n330 out_p.n329 0.754
R5170 out_p.n329 out_p.n328 0.754
R5171 out_p.n328 out_p.n327 0.754
R5172 out_p.n348 out_p.n347 0.754
R5173 out_p.n347 out_p.n346 0.754
R5174 out_p.n346 out_p.n345 0.754
R5175 out_p.n345 out_p.n344 0.754
R5176 out_p.n343 out_p.n342 0.754
R5177 out_p.n342 out_p.n341 0.754
R5178 out_p.n341 out_p.n340 0.754
R5179 out_p.n340 out_p.n339 0.754
R5180 out_p.n360 out_p.n359 0.754
R5181 out_p.n359 out_p.n358 0.754
R5182 out_p.n358 out_p.n357 0.754
R5183 out_p.n357 out_p.n356 0.754
R5184 out_p.n355 out_p.n354 0.754
R5185 out_p.n354 out_p.n353 0.754
R5186 out_p.n353 out_p.n352 0.754
R5187 out_p.n352 out_p.n351 0.754
R5188 out_p.n372 out_p.n371 0.754
R5189 out_p.n371 out_p.n370 0.754
R5190 out_p.n370 out_p.n369 0.754
R5191 out_p.n369 out_p.n368 0.754
R5192 out_p.n367 out_p.n366 0.754
R5193 out_p.n366 out_p.n365 0.754
R5194 out_p.n365 out_p.n364 0.754
R5195 out_p.n364 out_p.n363 0.754
R5196 out_p.n384 out_p.n383 0.754
R5197 out_p.n383 out_p.n382 0.754
R5198 out_p.n382 out_p.n381 0.754
R5199 out_p.n381 out_p.n380 0.754
R5200 out_p.n379 out_p.n378 0.754
R5201 out_p.n378 out_p.n377 0.754
R5202 out_p.n377 out_p.n376 0.754
R5203 out_p.n376 out_p.n375 0.754
R5204 out_p.n396 out_p.n395 0.754
R5205 out_p.n395 out_p.n394 0.754
R5206 out_p.n394 out_p.n393 0.754
R5207 out_p.n393 out_p.n392 0.754
R5208 out_p.n391 out_p.n390 0.754
R5209 out_p.n390 out_p.n389 0.754
R5210 out_p.n389 out_p.n388 0.754
R5211 out_p.n388 out_p.n387 0.754
R5212 out_p.n408 out_p.n407 0.754
R5213 out_p.n407 out_p.n406 0.754
R5214 out_p.n406 out_p.n405 0.754
R5215 out_p.n405 out_p.n404 0.754
R5216 out_p.n403 out_p.n402 0.754
R5217 out_p.n402 out_p.n401 0.754
R5218 out_p.n401 out_p.n400 0.754
R5219 out_p.n400 out_p.n399 0.754
R5220 out_p.n420 out_p.n419 0.754
R5221 out_p.n419 out_p.n418 0.754
R5222 out_p.n418 out_p.n417 0.754
R5223 out_p.n417 out_p.n416 0.754
R5224 out_p.n415 out_p.n414 0.754
R5225 out_p.n414 out_p.n413 0.754
R5226 out_p.n413 out_p.n412 0.754
R5227 out_p.n412 out_p.n411 0.754
R5228 out_p.n432 out_p.n431 0.754
R5229 out_p.n431 out_p.n430 0.754
R5230 out_p.n430 out_p.n429 0.754
R5231 out_p.n429 out_p.n428 0.754
R5232 out_p.n427 out_p.n426 0.754
R5233 out_p.n426 out_p.n425 0.754
R5234 out_p.n425 out_p.n424 0.754
R5235 out_p.n424 out_p.n423 0.754
R5236 out_p.n444 out_p.n443 0.754
R5237 out_p.n443 out_p.n442 0.754
R5238 out_p.n442 out_p.n441 0.754
R5239 out_p.n441 out_p.n440 0.754
R5240 out_p.n439 out_p.n438 0.754
R5241 out_p.n438 out_p.n437 0.754
R5242 out_p.n437 out_p.n436 0.754
R5243 out_p.n436 out_p.n435 0.754
R5244 out_p.n456 out_p.n455 0.754
R5245 out_p.n455 out_p.n454 0.754
R5246 out_p.n454 out_p.n453 0.754
R5247 out_p.n453 out_p.n452 0.754
R5248 out_p.n451 out_p.n450 0.754
R5249 out_p.n450 out_p.n449 0.754
R5250 out_p.n449 out_p.n448 0.754
R5251 out_p.n448 out_p.n447 0.754
R5252 out_p.n468 out_p.n467 0.754
R5253 out_p.n467 out_p.n466 0.754
R5254 out_p.n466 out_p.n465 0.754
R5255 out_p.n465 out_p.n464 0.754
R5256 out_p.n463 out_p.n462 0.754
R5257 out_p.n462 out_p.n461 0.754
R5258 out_p.n461 out_p.n460 0.754
R5259 out_p.n460 out_p.n459 0.754
R5260 out_p.n480 out_p.n479 0.754
R5261 out_p.n479 out_p.n478 0.754
R5262 out_p.n478 out_p.n477 0.754
R5263 out_p.n477 out_p.n476 0.754
R5264 out_p.n475 out_p.n474 0.754
R5265 out_p.n474 out_p.n473 0.754
R5266 out_p.n473 out_p.n472 0.754
R5267 out_p.n472 out_p.n471 0.754
R5268 out_p.n492 out_p.n491 0.754
R5269 out_p.n491 out_p.n490 0.754
R5270 out_p.n490 out_p.n489 0.754
R5271 out_p.n489 out_p.n488 0.754
R5272 out_p.n487 out_p.n486 0.754
R5273 out_p.n486 out_p.n485 0.754
R5274 out_p.n485 out_p.n484 0.754
R5275 out_p.n484 out_p.n483 0.754
R5276 out_p.n504 out_p.n503 0.754
R5277 out_p.n503 out_p.n502 0.754
R5278 out_p.n502 out_p.n501 0.754
R5279 out_p.n501 out_p.n500 0.754
R5280 out_p.n499 out_p.n498 0.754
R5281 out_p.n498 out_p.n497 0.754
R5282 out_p.n497 out_p.n496 0.754
R5283 out_p.n496 out_p.n495 0.754
R5284 out_p.n516 out_p.n515 0.754
R5285 out_p.n515 out_p.n514 0.754
R5286 out_p.n514 out_p.n513 0.754
R5287 out_p.n513 out_p.n512 0.754
R5288 out_p.n511 out_p.n510 0.754
R5289 out_p.n510 out_p.n509 0.754
R5290 out_p.n509 out_p.n508 0.754
R5291 out_p.n508 out_p.n507 0.754
R5292 out_p.n528 out_p.n527 0.754
R5293 out_p.n527 out_p.n526 0.754
R5294 out_p.n526 out_p.n525 0.754
R5295 out_p.n525 out_p.n524 0.754
R5296 out_p.n523 out_p.n522 0.754
R5297 out_p.n522 out_p.n521 0.754
R5298 out_p.n521 out_p.n520 0.754
R5299 out_p.n520 out_p.n519 0.754
R5300 out_p.n540 out_p.n539 0.754
R5301 out_p.n539 out_p.n538 0.754
R5302 out_p.n538 out_p.n537 0.754
R5303 out_p.n537 out_p.n536 0.754
R5304 out_p.n535 out_p.n534 0.754
R5305 out_p.n534 out_p.n533 0.754
R5306 out_p.n533 out_p.n532 0.754
R5307 out_p.n532 out_p.n531 0.754
R5308 out_p.n552 out_p.n551 0.754
R5309 out_p.n551 out_p.n550 0.754
R5310 out_p.n550 out_p.n549 0.754
R5311 out_p.n549 out_p.n548 0.754
R5312 out_p.n547 out_p.n546 0.754
R5313 out_p.n546 out_p.n545 0.754
R5314 out_p.n545 out_p.n544 0.754
R5315 out_p.n544 out_p.n543 0.754
R5316 out_p.n564 out_p.n563 0.754
R5317 out_p.n563 out_p.n562 0.754
R5318 out_p.n562 out_p.n561 0.754
R5319 out_p.n561 out_p.n560 0.754
R5320 out_p.n559 out_p.n558 0.754
R5321 out_p.n558 out_p.n557 0.754
R5322 out_p.n557 out_p.n556 0.754
R5323 out_p.n556 out_p.n555 0.754
R5324 out_p.n576 out_p.n575 0.754
R5325 out_p.n575 out_p.n574 0.754
R5326 out_p.n574 out_p.n573 0.754
R5327 out_p.n573 out_p.n572 0.754
R5328 out_p.n571 out_p.n570 0.754
R5329 out_p.n570 out_p.n569 0.754
R5330 out_p.n569 out_p.n568 0.754
R5331 out_p.n568 out_p.n567 0.754
R5332 out_p.n588 out_p.n587 0.754
R5333 out_p.n587 out_p.n586 0.754
R5334 out_p.n586 out_p.n585 0.754
R5335 out_p.n585 out_p.n584 0.754
R5336 out_p.n583 out_p.n582 0.754
R5337 out_p.n582 out_p.n581 0.754
R5338 out_p.n581 out_p.n580 0.754
R5339 out_p.n580 out_p.n579 0.754
R5340 out_p.n600 out_p.n599 0.754
R5341 out_p.n599 out_p.n598 0.754
R5342 out_p.n598 out_p.n597 0.754
R5343 out_p.n597 out_p.n596 0.754
R5344 out_p.n595 out_p.n594 0.754
R5345 out_p.n594 out_p.n593 0.754
R5346 out_p.n593 out_p.n592 0.754
R5347 out_p.n592 out_p.n591 0.754
R5348 out_p.n612 out_p.n611 0.754
R5349 out_p.n611 out_p.n610 0.754
R5350 out_p.n610 out_p.n609 0.754
R5351 out_p.n609 out_p.n608 0.754
R5352 out_p.n607 out_p.n606 0.754
R5353 out_p.n606 out_p.n605 0.754
R5354 out_p.n605 out_p.n604 0.754
R5355 out_p.n604 out_p.n603 0.754
R5356 out_p.n624 out_p.n623 0.754
R5357 out_p.n623 out_p.n622 0.754
R5358 out_p.n622 out_p.n621 0.754
R5359 out_p.n621 out_p.n620 0.754
R5360 out_p.n619 out_p.n618 0.754
R5361 out_p.n618 out_p.n617 0.754
R5362 out_p.n617 out_p.n616 0.754
R5363 out_p.n616 out_p.n615 0.754
R5364 out_p.n636 out_p.n635 0.754
R5365 out_p.n635 out_p.n634 0.754
R5366 out_p.n634 out_p.n633 0.754
R5367 out_p.n633 out_p.n632 0.754
R5368 out_p.n631 out_p.n630 0.754
R5369 out_p.n630 out_p.n629 0.754
R5370 out_p.n629 out_p.n628 0.754
R5371 out_p.n628 out_p.n627 0.754
R5372 out_p.n648 out_p.n647 0.754
R5373 out_p.n647 out_p.n646 0.754
R5374 out_p.n646 out_p.n645 0.754
R5375 out_p.n645 out_p.n644 0.754
R5376 out_p.n643 out_p.n642 0.754
R5377 out_p.n642 out_p.n641 0.754
R5378 out_p.n641 out_p.n640 0.754
R5379 out_p.n640 out_p.n639 0.754
R5380 out_p.n660 out_p.n659 0.754
R5381 out_p.n659 out_p.n658 0.754
R5382 out_p.n658 out_p.n657 0.754
R5383 out_p.n657 out_p.n656 0.754
R5384 out_p.n655 out_p.n654 0.754
R5385 out_p.n654 out_p.n653 0.754
R5386 out_p.n653 out_p.n652 0.754
R5387 out_p.n652 out_p.n651 0.754
R5388 out_p.n672 out_p.n671 0.754
R5389 out_p.n671 out_p.n670 0.754
R5390 out_p.n670 out_p.n669 0.754
R5391 out_p.n669 out_p.n668 0.754
R5392 out_p.n667 out_p.n666 0.754
R5393 out_p.n666 out_p.n665 0.754
R5394 out_p.n665 out_p.n664 0.754
R5395 out_p.n664 out_p.n663 0.754
R5396 out_p.n684 out_p.n683 0.754
R5397 out_p.n683 out_p.n682 0.754
R5398 out_p.n682 out_p.n681 0.754
R5399 out_p.n681 out_p.n680 0.754
R5400 out_p.n679 out_p.n678 0.754
R5401 out_p.n678 out_p.n677 0.754
R5402 out_p.n677 out_p.n676 0.754
R5403 out_p.n676 out_p.n675 0.754
R5404 out_p.n696 out_p.n695 0.754
R5405 out_p.n695 out_p.n694 0.754
R5406 out_p.n694 out_p.n693 0.754
R5407 out_p.n693 out_p.n692 0.754
R5408 out_p.n691 out_p.n690 0.754
R5409 out_p.n690 out_p.n689 0.754
R5410 out_p.n689 out_p.n688 0.754
R5411 out_p.n688 out_p.n687 0.754
R5412 out_p.n708 out_p.n707 0.754
R5413 out_p.n707 out_p.n706 0.754
R5414 out_p.n706 out_p.n705 0.754
R5415 out_p.n705 out_p.n704 0.754
R5416 out_p.n703 out_p.n702 0.754
R5417 out_p.n702 out_p.n701 0.754
R5418 out_p.n701 out_p.n700 0.754
R5419 out_p.n700 out_p.n699 0.754
R5420 out_p.n720 out_p.n719 0.754
R5421 out_p.n719 out_p.n718 0.754
R5422 out_p.n718 out_p.n717 0.754
R5423 out_p.n717 out_p.n716 0.754
R5424 out_p.n715 out_p.n714 0.754
R5425 out_p.n714 out_p.n713 0.754
R5426 out_p.n713 out_p.n712 0.754
R5427 out_p.n712 out_p.n711 0.754
R5428 out_p.n732 out_p.n731 0.754
R5429 out_p.n731 out_p.n730 0.754
R5430 out_p.n730 out_p.n729 0.754
R5431 out_p.n729 out_p.n728 0.754
R5432 out_p.n727 out_p.n726 0.754
R5433 out_p.n726 out_p.n725 0.754
R5434 out_p.n725 out_p.n724 0.754
R5435 out_p.n724 out_p.n723 0.754
R5436 out_p.n744 out_p.n743 0.754
R5437 out_p.n743 out_p.n742 0.754
R5438 out_p.n742 out_p.n741 0.754
R5439 out_p.n741 out_p.n740 0.754
R5440 out_p.n739 out_p.n738 0.754
R5441 out_p.n738 out_p.n737 0.754
R5442 out_p.n737 out_p.n736 0.754
R5443 out_p.n736 out_p.n735 0.754
R5444 out_p.n756 out_p.n755 0.754
R5445 out_p.n755 out_p.n754 0.754
R5446 out_p.n754 out_p.n753 0.754
R5447 out_p.n753 out_p.n752 0.754
R5448 out_p.n751 out_p.n750 0.754
R5449 out_p.n750 out_p.n749 0.754
R5450 out_p.n749 out_p.n748 0.754
R5451 out_p.n748 out_p.n747 0.754
R5452 out_p.n768 out_p.n767 0.754
R5453 out_p.n767 out_p.n766 0.754
R5454 out_p.n766 out_p.n765 0.754
R5455 out_p.n765 out_p.n764 0.754
R5456 out_p.n763 out_p.n762 0.754
R5457 out_p.n762 out_p.n761 0.754
R5458 out_p.n761 out_p.n760 0.754
R5459 out_p.n760 out_p.n759 0.754
R5460 out_p.n780 out_p.n779 0.754
R5461 out_p.n779 out_p.n778 0.754
R5462 out_p.n778 out_p.n777 0.754
R5463 out_p.n777 out_p.n776 0.754
R5464 out_p.n775 out_p.n774 0.754
R5465 out_p.n774 out_p.n773 0.754
R5466 out_p.n773 out_p.n772 0.754
R5467 out_p.n772 out_p.n771 0.754
R5468 out_p.n792 out_p.n791 0.754
R5469 out_p.n791 out_p.n790 0.754
R5470 out_p.n790 out_p.n789 0.754
R5471 out_p.n789 out_p.n788 0.754
R5472 out_p.n787 out_p.n786 0.754
R5473 out_p.n786 out_p.n785 0.754
R5474 out_p.n785 out_p.n784 0.754
R5475 out_p.n784 out_p.n783 0.754
R5476 out_p.n804 out_p.n803 0.754
R5477 out_p.n803 out_p.n802 0.754
R5478 out_p.n802 out_p.n801 0.754
R5479 out_p.n801 out_p.n800 0.754
R5480 out_p.n799 out_p.n798 0.754
R5481 out_p.n798 out_p.n797 0.754
R5482 out_p.n797 out_p.n796 0.754
R5483 out_p.n796 out_p.n795 0.754
R5484 out_p.n816 out_p.n815 0.754
R5485 out_p.n815 out_p.n814 0.754
R5486 out_p.n814 out_p.n813 0.754
R5487 out_p.n813 out_p.n812 0.754
R5488 out_p.n811 out_p.n810 0.754
R5489 out_p.n810 out_p.n809 0.754
R5490 out_p.n809 out_p.n808 0.754
R5491 out_p.n808 out_p.n807 0.754
R5492 out_p.n828 out_p.n827 0.754
R5493 out_p.n827 out_p.n826 0.754
R5494 out_p.n826 out_p.n825 0.754
R5495 out_p.n825 out_p.n824 0.754
R5496 out_p.n823 out_p.n822 0.754
R5497 out_p.n822 out_p.n821 0.754
R5498 out_p.n821 out_p.n820 0.754
R5499 out_p.n820 out_p.n819 0.754
R5500 out_p.n840 out_p.n839 0.754
R5501 out_p.n839 out_p.n838 0.754
R5502 out_p.n838 out_p.n837 0.754
R5503 out_p.n837 out_p.n836 0.754
R5504 out_p.n835 out_p.n834 0.754
R5505 out_p.n834 out_p.n833 0.754
R5506 out_p.n833 out_p.n832 0.754
R5507 out_p.n832 out_p.n831 0.754
R5508 out_p.n852 out_p.n851 0.754
R5509 out_p.n851 out_p.n850 0.754
R5510 out_p.n850 out_p.n849 0.754
R5511 out_p.n849 out_p.n848 0.754
R5512 out_p.n847 out_p.n846 0.754
R5513 out_p.n846 out_p.n845 0.754
R5514 out_p.n845 out_p.n844 0.754
R5515 out_p.n844 out_p.n843 0.754
R5516 out_p.n864 out_p.n863 0.754
R5517 out_p.n863 out_p.n862 0.754
R5518 out_p.n862 out_p.n861 0.754
R5519 out_p.n861 out_p.n860 0.754
R5520 out_p.n859 out_p.n858 0.754
R5521 out_p.n858 out_p.n857 0.754
R5522 out_p.n857 out_p.n856 0.754
R5523 out_p.n856 out_p.n855 0.754
R5524 out_p.n876 out_p.n875 0.754
R5525 out_p.n875 out_p.n874 0.754
R5526 out_p.n874 out_p.n873 0.754
R5527 out_p.n873 out_p.n872 0.754
R5528 out_p.n871 out_p.n870 0.754
R5529 out_p.n870 out_p.n869 0.754
R5530 out_p.n869 out_p.n868 0.754
R5531 out_p.n868 out_p.n867 0.754
R5532 out_p.n888 out_p.n887 0.754
R5533 out_p.n887 out_p.n886 0.754
R5534 out_p.n886 out_p.n885 0.754
R5535 out_p.n885 out_p.n884 0.754
R5536 out_p.n883 out_p.n882 0.754
R5537 out_p.n882 out_p.n881 0.754
R5538 out_p.n881 out_p.n880 0.754
R5539 out_p.n880 out_p.n879 0.754
R5540 out_p.n900 out_p.n899 0.754
R5541 out_p.n899 out_p.n898 0.754
R5542 out_p.n898 out_p.n897 0.754
R5543 out_p.n897 out_p.n896 0.754
R5544 out_p.n895 out_p.n894 0.754
R5545 out_p.n894 out_p.n893 0.754
R5546 out_p.n893 out_p.n892 0.754
R5547 out_p.n892 out_p.n891 0.754
R5548 out_p.n913 out_p.n902 0.554
R5549 out_p.n914 out_p.n890 0.554
R5550 out_p.n915 out_p.n878 0.554
R5551 out_p.n916 out_p.n866 0.554
R5552 out_p.n917 out_p.n854 0.554
R5553 out_p.n918 out_p.n842 0.554
R5554 out_p.n919 out_p.n830 0.554
R5555 out_p.n920 out_p.n818 0.554
R5556 out_p.n921 out_p.n806 0.554
R5557 out_p.n922 out_p.n794 0.554
R5558 out_p.n923 out_p.n782 0.554
R5559 out_p.n924 out_p.n770 0.554
R5560 out_p.n925 out_p.n758 0.554
R5561 out_p.n926 out_p.n746 0.554
R5562 out_p.n927 out_p.n734 0.554
R5563 out_p.n928 out_p.n722 0.554
R5564 out_p.n929 out_p.n710 0.554
R5565 out_p.n930 out_p.n698 0.554
R5566 out_p.n931 out_p.n686 0.554
R5567 out_p.n932 out_p.n674 0.554
R5568 out_p.n933 out_p.n662 0.554
R5569 out_p.n934 out_p.n650 0.554
R5570 out_p.n935 out_p.n638 0.554
R5571 out_p.n936 out_p.n626 0.554
R5572 out_p.n937 out_p.n614 0.554
R5573 out_p.n938 out_p.n602 0.554
R5574 out_p.n939 out_p.n590 0.554
R5575 out_p.n940 out_p.n578 0.554
R5576 out_p.n941 out_p.n566 0.554
R5577 out_p.n942 out_p.n554 0.554
R5578 out_p.n943 out_p.n542 0.554
R5579 out_p.n944 out_p.n530 0.554
R5580 out_p.n945 out_p.n518 0.554
R5581 out_p.n946 out_p.n506 0.554
R5582 out_p.n947 out_p.n494 0.554
R5583 out_p.n948 out_p.n482 0.554
R5584 out_p.n949 out_p.n470 0.554
R5585 out_p.n950 out_p.n458 0.554
R5586 out_p.n951 out_p.n446 0.554
R5587 out_p.n952 out_p.n434 0.554
R5588 out_p.n953 out_p.n422 0.554
R5589 out_p.n954 out_p.n410 0.554
R5590 out_p.n955 out_p.n398 0.554
R5591 out_p.n956 out_p.n386 0.554
R5592 out_p.n957 out_p.n374 0.554
R5593 out_p.n958 out_p.n362 0.554
R5594 out_p.n959 out_p.n350 0.554
R5595 out_p.n960 out_p.n338 0.554
R5596 out_p.n961 out_p.n326 0.554
R5597 out_p.n962 out_p.n314 0.554
R5598 out_p.n963 out_p.n302 0.554
R5599 out_p.n964 out_p.n290 0.554
R5600 out_p.n965 out_p.n278 0.554
R5601 out_p.n966 out_p.n266 0.554
R5602 out_p.n967 out_p.n254 0.554
R5603 out_p.n968 out_p.n242 0.554
R5604 out_p.n969 out_p.n230 0.554
R5605 out_p.n970 out_p.n218 0.554
R5606 out_p.n971 out_p.n206 0.554
R5607 out_p.n972 out_p.n194 0.554
R5608 out_p.n973 out_p.n182 0.554
R5609 out_p out_p.n180 0.554
R5610 out_p.n178 out_p.n11 0.554
R5611 out_p.n167 out_p.n13 0.554
R5612 out_p.n156 out_p.n15 0.554
R5613 out_p.n145 out_p.n17 0.554
R5614 out_p.n134 out_p.n19 0.554
R5615 out_p.n123 out_p.n21 0.554
R5616 out_p.n112 out_p.n23 0.554
R5617 out_p.n101 out_p.n25 0.554
R5618 out_p.n90 out_p.n27 0.554
R5619 out_p.n79 out_p.n29 0.554
R5620 out_p.n68 out_p.n31 0.554
R5621 out_p.n57 out_p.n33 0.554
R5622 out_p.n46 out_p.n35 0.554
R5623 out_p.n913 out_p.n912 0.541
R5624 out_p.n46 out_p.n45 0.524
R5625 out_p.n57 out_p.n56 0.524
R5626 out_p.n68 out_p.n67 0.524
R5627 out_p.n79 out_p.n78 0.524
R5628 out_p.n90 out_p.n89 0.524
R5629 out_p.n101 out_p.n100 0.524
R5630 out_p.n112 out_p.n111 0.524
R5631 out_p.n123 out_p.n122 0.524
R5632 out_p.n134 out_p.n133 0.524
R5633 out_p.n145 out_p.n144 0.524
R5634 out_p.n156 out_p.n155 0.524
R5635 out_p.n167 out_p.n166 0.524
R5636 out_p.n178 out_p.n177 0.524
R5637 out_p out_p.n9 0.524
R5638 out_p.n973 out_p.n192 0.524
R5639 out_p.n972 out_p.n204 0.524
R5640 out_p.n971 out_p.n216 0.524
R5641 out_p.n970 out_p.n228 0.524
R5642 out_p.n969 out_p.n240 0.524
R5643 out_p.n968 out_p.n252 0.524
R5644 out_p.n967 out_p.n264 0.524
R5645 out_p.n966 out_p.n276 0.524
R5646 out_p.n965 out_p.n288 0.524
R5647 out_p.n964 out_p.n300 0.524
R5648 out_p.n963 out_p.n312 0.524
R5649 out_p.n962 out_p.n324 0.524
R5650 out_p.n961 out_p.n336 0.524
R5651 out_p.n960 out_p.n348 0.524
R5652 out_p.n959 out_p.n360 0.524
R5653 out_p.n958 out_p.n372 0.524
R5654 out_p.n957 out_p.n384 0.524
R5655 out_p.n956 out_p.n396 0.524
R5656 out_p.n955 out_p.n408 0.524
R5657 out_p.n954 out_p.n420 0.524
R5658 out_p.n953 out_p.n432 0.524
R5659 out_p.n952 out_p.n444 0.524
R5660 out_p.n951 out_p.n456 0.524
R5661 out_p.n950 out_p.n468 0.524
R5662 out_p.n949 out_p.n480 0.524
R5663 out_p.n948 out_p.n492 0.524
R5664 out_p.n947 out_p.n504 0.524
R5665 out_p.n946 out_p.n516 0.524
R5666 out_p.n945 out_p.n528 0.524
R5667 out_p.n944 out_p.n540 0.524
R5668 out_p.n943 out_p.n552 0.524
R5669 out_p.n942 out_p.n564 0.524
R5670 out_p.n941 out_p.n576 0.524
R5671 out_p.n940 out_p.n588 0.524
R5672 out_p.n939 out_p.n600 0.524
R5673 out_p.n938 out_p.n612 0.524
R5674 out_p.n937 out_p.n624 0.524
R5675 out_p.n936 out_p.n636 0.524
R5676 out_p.n935 out_p.n648 0.524
R5677 out_p.n934 out_p.n660 0.524
R5678 out_p.n933 out_p.n672 0.524
R5679 out_p.n932 out_p.n684 0.524
R5680 out_p.n931 out_p.n696 0.524
R5681 out_p.n930 out_p.n708 0.524
R5682 out_p.n929 out_p.n720 0.524
R5683 out_p.n928 out_p.n732 0.524
R5684 out_p.n927 out_p.n744 0.524
R5685 out_p.n926 out_p.n756 0.524
R5686 out_p.n925 out_p.n768 0.524
R5687 out_p.n924 out_p.n780 0.524
R5688 out_p.n923 out_p.n792 0.524
R5689 out_p.n922 out_p.n804 0.524
R5690 out_p.n921 out_p.n816 0.524
R5691 out_p.n920 out_p.n828 0.524
R5692 out_p.n919 out_p.n840 0.524
R5693 out_p.n918 out_p.n852 0.524
R5694 out_p.n917 out_p.n864 0.524
R5695 out_p.n916 out_p.n876 0.524
R5696 out_p.n915 out_p.n888 0.524
R5697 out_p.n914 out_p.n900 0.524
R5698 out_p.n57 out_p.n46 0.002
R5699 out_p.n68 out_p.n57 0.002
R5700 out_p.n79 out_p.n68 0.002
R5701 out_p.n90 out_p.n79 0.002
R5702 out_p.n101 out_p.n90 0.002
R5703 out_p.n112 out_p.n101 0.002
R5704 out_p.n123 out_p.n112 0.002
R5705 out_p.n134 out_p.n123 0.002
R5706 out_p.n145 out_p.n134 0.002
R5707 out_p.n156 out_p.n145 0.002
R5708 out_p.n167 out_p.n156 0.002
R5709 out_p.n178 out_p.n167 0.002
R5710 out_p out_p.n178 0.002
R5711 out_p out_p.n973 0.002
R5712 out_p.n973 out_p.n972 0.002
R5713 out_p.n972 out_p.n971 0.002
R5714 out_p.n971 out_p.n970 0.002
R5715 out_p.n970 out_p.n969 0.002
R5716 out_p.n969 out_p.n968 0.002
R5717 out_p.n968 out_p.n967 0.002
R5718 out_p.n967 out_p.n966 0.002
R5719 out_p.n966 out_p.n965 0.002
R5720 out_p.n965 out_p.n964 0.002
R5721 out_p.n964 out_p.n963 0.002
R5722 out_p.n963 out_p.n962 0.002
R5723 out_p.n962 out_p.n961 0.002
R5724 out_p.n961 out_p.n960 0.002
R5725 out_p.n960 out_p.n959 0.002
R5726 out_p.n959 out_p.n958 0.002
R5727 out_p.n958 out_p.n957 0.002
R5728 out_p.n957 out_p.n956 0.002
R5729 out_p.n956 out_p.n955 0.002
R5730 out_p.n955 out_p.n954 0.002
R5731 out_p.n954 out_p.n953 0.002
R5732 out_p.n953 out_p.n952 0.002
R5733 out_p.n952 out_p.n951 0.002
R5734 out_p.n951 out_p.n950 0.002
R5735 out_p.n950 out_p.n949 0.002
R5736 out_p.n949 out_p.n948 0.002
R5737 out_p.n948 out_p.n947 0.002
R5738 out_p.n947 out_p.n946 0.002
R5739 out_p.n946 out_p.n945 0.002
R5740 out_p.n945 out_p.n944 0.002
R5741 out_p.n944 out_p.n943 0.002
R5742 out_p.n943 out_p.n942 0.002
R5743 out_p.n942 out_p.n941 0.002
R5744 out_p.n941 out_p.n940 0.002
R5745 out_p.n940 out_p.n939 0.002
R5746 out_p.n939 out_p.n938 0.002
R5747 out_p.n938 out_p.n937 0.002
R5748 out_p.n937 out_p.n936 0.002
R5749 out_p.n936 out_p.n935 0.002
R5750 out_p.n935 out_p.n934 0.002
R5751 out_p.n934 out_p.n933 0.002
R5752 out_p.n933 out_p.n932 0.002
R5753 out_p.n932 out_p.n931 0.002
R5754 out_p.n931 out_p.n930 0.002
R5755 out_p.n930 out_p.n929 0.002
R5756 out_p.n929 out_p.n928 0.002
R5757 out_p.n928 out_p.n927 0.002
R5758 out_p.n927 out_p.n926 0.002
R5759 out_p.n926 out_p.n925 0.002
R5760 out_p.n925 out_p.n924 0.002
R5761 out_p.n924 out_p.n923 0.002
R5762 out_p.n923 out_p.n922 0.002
R5763 out_p.n922 out_p.n921 0.002
R5764 out_p.n921 out_p.n920 0.002
R5765 out_p.n920 out_p.n919 0.002
R5766 out_p.n919 out_p.n918 0.002
R5767 out_p.n918 out_p.n917 0.002
R5768 out_p.n917 out_p.n916 0.002
R5769 out_p.n916 out_p.n915 0.002
R5770 out_p.n915 out_p.n914 0.002
R5771 out_p.n914 out_p.n913 0.002
R5772 vdd.n530 vdd.n529 9250.59
R5773 vdd.n536 vdd.n535 9250.59
R5774 vdd.n528 vdd.n527 2878.29
R5775 vdd.n534 vdd.n533 2869.55
R5776 vdd.n537 vdd.n530 2247.42
R5777 vdd.n537 vdd.n536 2247.42
R5778 vdd.n534 vdd.n531 940.477
R5779 vdd.n528 vdd.n525 940.476
R5780 vdd.n536 vdd.n534 940.476
R5781 vdd.n530 vdd.n528 940.476
R5782 vdd.n608 vdd.t253 10.284
R5783 vdd.n12 vdd.t517 8.711
R5784 vdd.n20 vdd.t1293 8.131
R5785 vdd.n19 vdd.t733 8.131
R5786 vdd.n18 vdd.t523 8.131
R5787 vdd.n17 vdd.t391 8.131
R5788 vdd.n16 vdd.t1329 8.131
R5789 vdd.n15 vdd.t923 8.131
R5790 vdd.n14 vdd.t1062 8.131
R5791 vdd.n13 vdd.t1284 8.131
R5792 vdd.n12 vdd.t731 8.131
R5793 vdd.n616 vdd.t1041 8.126
R5794 vdd.n615 vdd.t482 8.126
R5795 vdd.n614 vdd.t263 8.126
R5796 vdd.n613 vdd.t137 8.126
R5797 vdd.n612 vdd.t1074 8.126
R5798 vdd.n608 vdd.t473 8.126
R5799 vdd.n609 vdd.t1032 8.126
R5800 vdd.n610 vdd.t798 8.126
R5801 vdd.n611 vdd.t665 8.126
R5802 vdd.n618 vdd.t43 8.126
R5803 vdd.n618 vdd.t1338 8.126
R5804 vdd.n619 vdd.t257 8.126
R5805 vdd.n619 vdd.t47 8.126
R5806 vdd.n620 vdd.t832 8.126
R5807 vdd.n620 vdd.t621 8.126
R5808 vdd.n621 vdd.t591 8.126
R5809 vdd.n621 vdd.t382 8.126
R5810 vdd.n622 vdd.t468 8.126
R5811 vdd.n622 vdd.t254 8.126
R5812 vdd.n623 vdd.t870 8.126
R5813 vdd.n623 vdd.t667 8.126
R5814 vdd.n624 vdd.t1431 8.126
R5815 vdd.n624 vdd.t1224 8.126
R5816 vdd.n625 vdd.t53 8.126
R5817 vdd.n625 vdd.t1347 8.126
R5818 vdd.n626 vdd.t268 8.126
R5819 vdd.n626 vdd.t56 8.126
R5820 vdd.n627 vdd.t839 8.126
R5821 vdd.n627 vdd.t625 8.126
R5822 vdd.n630 vdd.t1129 8.126
R5823 vdd.n630 vdd.t929 8.126
R5824 vdd.n631 vdd.t1342 8.126
R5825 vdd.n631 vdd.t1134 8.126
R5826 vdd.n632 vdd.t415 8.126
R5827 vdd.n632 vdd.t207 8.126
R5828 vdd.n633 vdd.t177 8.126
R5829 vdd.n633 vdd.t1468 8.126
R5830 vdd.n634 vdd.t44 8.126
R5831 vdd.n634 vdd.t1339 8.126
R5832 vdd.n635 vdd.t469 8.126
R5833 vdd.n635 vdd.t255 8.126
R5834 vdd.n636 vdd.t1030 8.126
R5835 vdd.n636 vdd.t829 8.126
R5836 vdd.n637 vdd.t1137 8.126
R5837 vdd.n637 vdd.t935 8.126
R5838 vdd.n638 vdd.t1350 8.126
R5839 vdd.n638 vdd.t1141 8.126
R5840 vdd.n639 vdd.t420 8.126
R5841 vdd.n639 vdd.t210 8.126
R5842 vdd.n646 vdd.t1372 8.126
R5843 vdd.n646 vdd.t1164 8.126
R5844 vdd.n647 vdd.t81 8.126
R5845 vdd.n647 vdd.t1378 8.126
R5846 vdd.n648 vdd.t657 8.126
R5847 vdd.n648 vdd.t461 8.126
R5848 vdd.n649 vdd.t412 8.126
R5849 vdd.n649 vdd.t204 8.126
R5850 vdd.n650 vdd.t281 8.126
R5851 vdd.n650 vdd.t75 8.126
R5852 vdd.n651 vdd.t703 8.126
R5853 vdd.n651 vdd.t499 8.126
R5854 vdd.n652 vdd.t1255 8.126
R5855 vdd.n652 vdd.t1066 8.126
R5856 vdd.n653 vdd.t1384 8.126
R5857 vdd.n653 vdd.t1174 8.126
R5858 vdd.n654 vdd.t90 8.126
R5859 vdd.n654 vdd.t1390 8.126
R5860 vdd.n655 vdd.t663 8.126
R5861 vdd.n655 vdd.t466 8.126
R5862 vdd.n658 vdd.t965 8.126
R5863 vdd.n658 vdd.t766 8.126
R5864 vdd.n659 vdd.t1168 8.126
R5865 vdd.n659 vdd.t968 8.126
R5866 vdd.n660 vdd.t247 8.126
R5867 vdd.n660 vdd.t38 8.126
R5868 vdd.n661 vdd.t1497 8.126
R5869 vdd.n661 vdd.t1299 8.126
R5870 vdd.n662 vdd.t1373 8.126
R5871 vdd.n662 vdd.t1165 8.126
R5872 vdd.n663 vdd.t284 8.126
R5873 vdd.n663 vdd.t76 8.126
R5874 vdd.n664 vdd.t863 8.126
R5875 vdd.n664 vdd.t654 8.126
R5876 vdd.n665 vdd.t974 8.126
R5877 vdd.n665 vdd.t774 8.126
R5878 vdd.n666 vdd.t1180 8.126
R5879 vdd.n666 vdd.t980 8.126
R5880 vdd.n667 vdd.t252 8.126
R5881 vdd.n667 vdd.t42 8.126
R5882 vdd.n674 vdd.t560 8.126
R5883 vdd.n674 vdd.t834 8.126
R5884 vdd.n675 vdd.t768 8.126
R5885 vdd.n675 vdd.t1043 8.126
R5886 vdd.n676 vdd.t1333 8.126
R5887 vdd.n676 vdd.t107 8.126
R5888 vdd.n677 vdd.t1099 8.126
R5889 vdd.n677 vdd.t1368 8.126
R5890 vdd.n678 vdd.t966 8.126
R5891 vdd.n678 vdd.t1230 8.126
R5892 vdd.n679 vdd.t1375 8.126
R5893 vdd.n679 vdd.t149 8.126
R5894 vdd.n680 vdd.t457 8.126
R5895 vdd.n680 vdd.t718 8.126
R5896 vdd.n681 vdd.t565 8.126
R5897 vdd.n681 vdd.t847 8.126
R5898 vdd.n682 vdd.t780 8.126
R5899 vdd.n682 vdd.t1053 8.126
R5900 vdd.n683 vdd.t1337 8.126
R5901 vdd.n683 vdd.t115 8.126
R5902 vdd.n686 vdd.t622 8.126
R5903 vdd.n686 vdd.t416 8.126
R5904 vdd.n687 vdd.t842 8.126
R5905 vdd.n687 vdd.t628 8.126
R5906 vdd.n688 vdd.t1407 8.126
R5907 vdd.n688 vdd.t1197 8.126
R5908 vdd.n689 vdd.t1160 8.126
R5909 vdd.n689 vdd.t960 8.126
R5910 vdd.n690 vdd.t1036 8.126
R5911 vdd.n690 vdd.t835 8.126
R5912 vdd.n691 vdd.t1440 8.126
R5913 vdd.n691 vdd.t1235 8.126
R5914 vdd.n692 vdd.t511 8.126
R5915 vdd.n692 vdd.t306 8.126
R5916 vdd.n693 vdd.t633 8.126
R5917 vdd.n693 vdd.t429 8.126
R5918 vdd.n694 vdd.t850 8.126
R5919 vdd.n694 vdd.t639 8.126
R5920 vdd.n695 vdd.t1412 8.126
R5921 vdd.n695 vdd.t1201 8.126
R5922 vdd.n702 vdd.t208 8.126
R5923 vdd.n702 vdd.t1 8.126
R5924 vdd.n703 vdd.t422 8.126
R5925 vdd.n703 vdd.t213 8.126
R5926 vdd.n704 vdd.t1000 8.126
R5927 vdd.n704 vdd.t799 8.126
R5928 vdd.n705 vdd.t760 8.126
R5929 vdd.n705 vdd.t554 8.126
R5930 vdd.n706 vdd.t623 8.126
R5931 vdd.n706 vdd.t417 8.126
R5932 vdd.n707 vdd.t1039 8.126
R5933 vdd.n707 vdd.t837 8.126
R5934 vdd.n708 vdd.t106 8.126
R5935 vdd.n708 vdd.t1406 8.126
R5936 vdd.n709 vdd.t217 8.126
R5937 vdd.n709 vdd.t6 8.126
R5938 vdd.n710 vdd.t437 8.126
R5939 vdd.n710 vdd.t225 8.126
R5940 vdd.n711 vdd.t1004 8.126
R5941 vdd.n711 vdd.t802 8.126
R5942 vdd.n714 vdd.t421 8.126
R5943 vdd.n714 vdd.t211 8.126
R5944 vdd.n715 vdd.t634 8.126
R5945 vdd.n715 vdd.t430 8.126
R5946 vdd.n716 vdd.t1199 8.126
R5947 vdd.n716 vdd.t1001 8.126
R5948 vdd.n717 vdd.t963 8.126
R5949 vdd.n717 vdd.t764 8.126
R5950 vdd.n718 vdd.t841 8.126
R5951 vdd.n718 vdd.t626 8.126
R5952 vdd.n719 vdd.t1238 8.126
R5953 vdd.n719 vdd.t1046 8.126
R5954 vdd.n720 vdd.t309 8.126
R5955 vdd.n720 vdd.t108 8.126
R5956 vdd.n721 vdd.t436 8.126
R5957 vdd.n721 vdd.t224 8.126
R5958 vdd.n722 vdd.t645 8.126
R5959 vdd.n722 vdd.t445 8.126
R5960 vdd.n723 vdd.t1204 8.126
R5961 vdd.n723 vdd.t1007 8.126
R5962 vdd.n730 vdd.t2 8.126
R5963 vdd.n730 vdd.t1304 8.126
R5964 vdd.n731 vdd.t218 8.126
R5965 vdd.n731 vdd.t8 8.126
R5966 vdd.n732 vdd.t800 8.126
R5967 vdd.n732 vdd.t593 8.126
R5968 vdd.n733 vdd.t556 8.126
R5969 vdd.n733 vdd.t353 8.126
R5970 vdd.n734 vdd.t424 8.126
R5971 vdd.n734 vdd.t212 8.126
R5972 vdd.n735 vdd.t843 8.126
R5973 vdd.n735 vdd.t629 8.126
R5974 vdd.n736 vdd.t1408 8.126
R5975 vdd.n736 vdd.t1198 8.126
R5976 vdd.n737 vdd.t14 8.126
R5977 vdd.n737 vdd.t1312 8.126
R5978 vdd.n738 vdd.t233 8.126
R5979 vdd.n738 vdd.t21 8.126
R5980 vdd.n739 vdd.t805 8.126
R5981 vdd.n739 vdd.t595 8.126
R5982 vdd.n742 vdd.t831 8.126
R5983 vdd.n742 vdd.t359 8.126
R5984 vdd.n743 vdd.t1034 8.126
R5985 vdd.n743 vdd.t572 8.126
R5986 vdd.n744 vdd.t103 8.126
R5987 vdd.n744 vdd.t1128 8.126
R5988 vdd.n745 vdd.t1361 8.126
R5989 vdd.n745 vdd.t902 8.126
R5990 vdd.n746 vdd.t1226 8.126
R5991 vdd.n746 vdd.t773 8.126
R5992 vdd.n747 vdd.t141 8.126
R5993 vdd.n747 vdd.t1175 8.126
R5994 vdd.n748 vdd.t714 8.126
R5995 vdd.n748 vdd.t249 8.126
R5996 vdd.n749 vdd.t836 8.126
R5997 vdd.n749 vdd.t365 8.126
R5998 vdd.n750 vdd.t1044 8.126
R5999 vdd.n750 vdd.t584 8.126
R6000 vdd.n751 vdd.t109 8.126
R6001 vdd.n751 vdd.t1135 8.126
R6002 vdd.n758 vdd.t564 8.126
R6003 vdd.n758 vdd.t772 8.126
R6004 vdd.n759 vdd.t779 8.126
R6005 vdd.n759 vdd.t979 8.126
R6006 vdd.n760 vdd.t1336 8.126
R6007 vdd.n760 vdd.t41 8.126
R6008 vdd.n761 vdd.t1103 8.126
R6009 vdd.n761 vdd.t1303 8.126
R6010 vdd.n762 vdd.t973 8.126
R6011 vdd.n762 vdd.t1172 8.126
R6012 vdd.n763 vdd.t1385 8.126
R6013 vdd.n763 vdd.t85 8.126
R6014 vdd.n764 vdd.t463 8.126
R6015 vdd.n764 vdd.t659 8.126
R6016 vdd.n765 vdd.t574 8.126
R6017 vdd.n765 vdd.t782 8.126
R6018 vdd.n766 vdd.t791 8.126
R6019 vdd.n766 vdd.t990 8.126
R6020 vdd.n767 vdd.t1344 8.126
R6021 vdd.n767 vdd.t49 8.126
R6022 vdd.n770 vdd.t971 8.126
R6023 vdd.n770 vdd.t885 8.126
R6024 vdd.n771 vdd.t1179 8.126
R6025 vdd.n771 vdd.t1089 8.126
R6026 vdd.n772 vdd.t251 8.126
R6027 vdd.n772 vdd.t157 8.126
R6028 vdd.n773 vdd.t0 8.126
R6029 vdd.n773 vdd.t1425 8.126
R6030 vdd.n774 vdd.t1382 8.126
R6031 vdd.n774 vdd.t1283 8.126
R6032 vdd.n775 vdd.t290 8.126
R6033 vdd.n775 vdd.t191 8.126
R6034 vdd.n776 vdd.t866 8.126
R6035 vdd.n776 vdd.t770 8.126
R6036 vdd.n777 vdd.t981 8.126
R6037 vdd.n777 vdd.t891 8.126
R6038 vdd.n778 vdd.t1189 8.126
R6039 vdd.n778 vdd.t1100 8.126
R6040 vdd.n779 vdd.t258 8.126
R6041 vdd.n779 vdd.t163 8.126
R6042 vdd.n786 vdd.t1085 8.126
R6043 vdd.n786 vdd.t1282 8.126
R6044 vdd.n787 vdd.t1288 8.126
R6045 vdd.n787 vdd.t1486 8.126
R6046 vdd.n788 vdd.t360 8.126
R6047 vdd.n788 vdd.t566 8.126
R6048 vdd.n789 vdd.t130 8.126
R6049 vdd.n789 vdd.t328 8.126
R6050 vdd.n790 vdd.t1480 8.126
R6051 vdd.n790 vdd.t187 8.126
R6052 vdd.n791 vdd.t397 8.126
R6053 vdd.n791 vdd.t607 8.126
R6054 vdd.n792 vdd.t969 8.126
R6055 vdd.n792 vdd.t1169 8.126
R6056 vdd.n793 vdd.t1093 8.126
R6057 vdd.n793 vdd.t1292 8.126
R6058 vdd.n794 vdd.t1300 8.126
R6059 vdd.n794 vdd.t1496 8.126
R6060 vdd.n795 vdd.t368 8.126
R6061 vdd.n795 vdd.t577 8.126
R6062 vdd.n798 vdd.t1479 8.126
R6063 vdd.n798 vdd.t186 8.126
R6064 vdd.n799 vdd.t195 8.126
R6065 vdd.n799 vdd.t403 8.126
R6066 vdd.n800 vdd.t775 8.126
R6067 vdd.n800 vdd.t975 8.126
R6068 vdd.n801 vdd.t528 8.126
R6069 vdd.n801 vdd.t735 8.126
R6070 vdd.n802 vdd.t393 8.126
R6071 vdd.n802 vdd.t602 8.126
R6072 vdd.n803 vdd.t818 8.126
R6073 vdd.n803 vdd.t1019 8.126
R6074 vdd.n804 vdd.t1379 8.126
R6075 vdd.n804 vdd.t80 8.126
R6076 vdd.n805 vdd.t1492 8.126
R6077 vdd.n805 vdd.t199 8.126
R6078 vdd.n806 vdd.t203 8.126
R6079 vdd.n806 vdd.t411 8.126
R6080 vdd.n807 vdd.t785 8.126
R6081 vdd.n807 vdd.t985 8.126
R6082 vdd.n814 vdd.t1256 8.126
R6083 vdd.n814 vdd.t135 8.126
R6084 vdd.n815 vdd.t1460 8.126
R6085 vdd.n815 vdd.t338 8.126
R6086 vdd.n816 vdd.t531 8.126
R6087 vdd.n816 vdd.t906 8.126
R6088 vdd.n817 vdd.t300 8.126
R6089 vdd.n817 vdd.t682 8.126
R6090 vdd.n818 vdd.t165 8.126
R6091 vdd.n818 vdd.t536 8.126
R6092 vdd.n819 vdd.t581 8.126
R6093 vdd.n819 vdd.t942 8.126
R6094 vdd.n820 vdd.t1132 8.126
R6095 vdd.n820 vdd.t3 8.126
R6096 vdd.n821 vdd.t1263 8.126
R6097 vdd.n821 vdd.t143 8.126
R6098 vdd.n822 vdd.t1469 8.126
R6099 vdd.n822 vdd.t351 8.126
R6100 vdd.n823 vdd.t540 8.126
R6101 vdd.n823 vdd.t912 8.126
R6102 vdd.n826 vdd.t334 8.126
R6103 vdd.n826 vdd.t534 8.126
R6104 vdd.n827 vdd.t541 8.126
R6105 vdd.n827 vdd.t747 8.126
R6106 vdd.n828 vdd.t1106 8.126
R6107 vdd.n828 vdd.t1307 8.126
R6108 vdd.n829 vdd.t880 8.126
R6109 vdd.n829 vdd.t1080 8.126
R6110 vdd.n830 vdd.t742 8.126
R6111 vdd.n830 vdd.t940 8.126
R6112 vdd.n831 vdd.t1146 8.126
R6113 vdd.n831 vdd.t1354 8.126
R6114 vdd.n832 vdd.t215 8.126
R6115 vdd.n832 vdd.t425 8.126
R6116 vdd.n833 vdd.t344 8.126
R6117 vdd.n833 vdd.t547 8.126
R6118 vdd.n834 vdd.t553 8.126
R6119 vdd.n834 vdd.t759 8.126
R6120 vdd.n835 vdd.t1111 8.126
R6121 vdd.n835 vdd.t1316 8.126
R6122 vdd.n842 vdd.t741 8.126
R6123 vdd.n842 vdd.t307 8.126
R6124 vdd.n843 vdd.t949 8.126
R6125 vdd.n843 vdd.t516 8.126
R6126 vdd.n844 vdd.t7 8.126
R6127 vdd.n844 vdd.t1083 8.126
R6128 vdd.n845 vdd.t1275 8.126
R6129 vdd.n845 vdd.t857 8.126
R6130 vdd.n846 vdd.t1142 8.126
R6131 vdd.n846 vdd.t720 8.126
R6132 vdd.n847 vdd.t60 8.126
R6133 vdd.n847 vdd.t1115 8.126
R6134 vdd.n848 vdd.t627 8.126
R6135 vdd.n848 vdd.t181 8.126
R6136 vdd.n849 vdd.t754 8.126
R6137 vdd.n849 vdd.t313 8.126
R6138 vdd.n850 vdd.t959 8.126
R6139 vdd.n850 vdd.t522 8.126
R6140 vdd.n851 vdd.t19 8.126
R6141 vdd.n851 vdd.t1088 8.126
R6142 vdd.n854 vdd.t512 8.126
R6143 vdd.n854 vdd.t719 8.126
R6144 vdd.n855 vdd.t724 8.126
R6145 vdd.n855 vdd.t918 8.126
R6146 vdd.n856 vdd.t1278 8.126
R6147 vdd.n856 vdd.t1475 8.126
R6148 vdd.n857 vdd.t1060 8.126
R6149 vdd.n857 vdd.t1249 8.126
R6150 vdd.n858 vdd.t914 8.126
R6151 vdd.n858 vdd.t1113 8.126
R6152 vdd.n859 vdd.t1321 8.126
R6153 vdd.n859 vdd.t25 8.126
R6154 vdd.n860 vdd.t386 8.126
R6155 vdd.n860 vdd.t596 8.126
R6156 vdd.n861 vdd.t518 8.126
R6157 vdd.n861 vdd.t728 8.126
R6158 vdd.n862 vdd.t732 8.126
R6159 vdd.n862 vdd.t926 8.126
R6160 vdd.n863 vdd.t1287 8.126
R6161 vdd.n863 vdd.t1483 8.126
R6162 vdd.n870 vdd.t913 8.126
R6163 vdd.n870 vdd.t1112 8.126
R6164 vdd.n871 vdd.t1119 8.126
R6165 vdd.n871 vdd.t1325 8.126
R6166 vdd.n872 vdd.t183 8.126
R6167 vdd.n872 vdd.t389 8.126
R6168 vdd.n873 vdd.t1448 8.126
R6169 vdd.n873 vdd.t158 8.126
R6170 vdd.n874 vdd.t1318 8.126
R6171 vdd.n874 vdd.t22 8.126
R6172 vdd.n875 vdd.t235 8.126
R6173 vdd.n875 vdd.t450 8.126
R6174 vdd.n876 vdd.t806 8.126
R6175 vdd.n876 vdd.t1008 8.126
R6176 vdd.n877 vdd.t924 8.126
R6177 vdd.n877 vdd.t1124 8.126
R6178 vdd.n878 vdd.t1126 8.126
R6179 vdd.n878 vdd.t1332 8.126
R6180 vdd.n879 vdd.t193 8.126
R6181 vdd.n879 vdd.t400 8.126
R6182 vdd.n882 vdd.t691 8.126
R6183 vdd.n882 vdd.t1064 8.126
R6184 vdd.n883 vdd.t892 8.126
R6185 vdd.n883 vdd.t1261 8.126
R6186 vdd.n884 vdd.t1451 8.126
R6187 vdd.n884 vdd.t331 8.126
R6188 vdd.n885 vdd.t1220 8.126
R6189 vdd.n885 vdd.t97 8.126
R6190 vdd.n886 vdd.t1090 8.126
R6191 vdd.n886 vdd.t1455 8.126
R6192 vdd.n887 vdd.t1489 8.126
R6193 vdd.n887 vdd.t373 8.126
R6194 vdd.n888 vdd.t569 8.126
R6195 vdd.n888 vdd.t932 8.126
R6196 vdd.n889 vdd.t699 8.126
R6197 vdd.n889 vdd.t1070 8.126
R6198 vdd.n890 vdd.t901 8.126
R6199 vdd.n890 vdd.t1270 8.126
R6200 vdd.n891 vdd.t1458 8.126
R6201 vdd.n891 vdd.t336 8.126
R6202 vdd.n898 vdd.t1257 8.126
R6203 vdd.n898 vdd.t1454 8.126
R6204 vdd.n899 vdd.t1461 8.126
R6205 vdd.n899 vdd.t170 8.126
R6206 vdd.n900 vdd.t532 8.126
R6207 vdd.n900 vdd.t738 8.126
R6208 vdd.n901 vdd.t301 8.126
R6209 vdd.n901 vdd.t508 8.126
R6210 vdd.n902 vdd.t164 8.126
R6211 vdd.n902 vdd.t369 8.126
R6212 vdd.n903 vdd.t582 8.126
R6213 vdd.n903 vdd.t788 8.126
R6214 vdd.n904 vdd.t1133 8.126
R6215 vdd.n904 vdd.t1341 8.126
R6216 vdd.n905 vdd.t1264 8.126
R6217 vdd.n905 vdd.t1463 8.126
R6218 vdd.n906 vdd.t1467 8.126
R6219 vdd.n906 vdd.t176 8.126
R6220 vdd.n907 vdd.t539 8.126
R6221 vdd.n907 vdd.t744 8.126
R6222 vdd.n910 vdd.t1031 8.126
R6223 vdd.n910 vdd.t1225 8.126
R6224 vdd.n911 vdd.t1228 8.126
R6225 vdd.n911 vdd.t1436 8.126
R6226 vdd.n912 vdd.t303 8.126
R6227 vdd.n912 vdd.t510 8.126
R6228 vdd.n913 vdd.t65 8.126
R6229 vdd.n913 vdd.t275 8.126
R6230 vdd.n914 vdd.t1433 8.126
R6231 vdd.n914 vdd.t139 8.126
R6232 vdd.n915 vdd.t341 8.126
R6233 vdd.n915 vdd.t543 8.126
R6234 vdd.n916 vdd.t908 8.126
R6235 vdd.n916 vdd.t1107 8.126
R6236 vdd.n917 vdd.t1035 8.126
R6237 vdd.n917 vdd.t1231 8.126
R6238 vdd.n918 vdd.t1237 8.126
R6239 vdd.n918 vdd.t1443 8.126
R6240 vdd.n919 vdd.t308 8.126
R6241 vdd.n919 vdd.t513 8.126
R6242 vdd.n926 vdd.t1432 8.126
R6243 vdd.n926 vdd.t138 8.126
R6244 vdd.n927 vdd.t144 8.126
R6245 vdd.n927 vdd.t345 8.126
R6246 vdd.n928 vdd.t715 8.126
R6247 vdd.n928 vdd.t909 8.126
R6248 vdd.n929 vdd.t488 8.126
R6249 vdd.n929 vdd.t685 8.126
R6250 vdd.n930 vdd.t339 8.126
R6251 vdd.n930 vdd.t542 8.126
R6252 vdd.n931 vdd.t752 8.126
R6253 vdd.n931 vdd.t952 8.126
R6254 vdd.n932 vdd.t1308 8.126
R6255 vdd.n932 vdd.t9 8.126
R6256 vdd.n933 vdd.t1438 8.126
R6257 vdd.n933 vdd.t148 8.126
R6258 vdd.n934 vdd.t152 8.126
R6259 vdd.n934 vdd.t354 8.126
R6260 vdd.n935 vdd.t722 8.126
R6261 vdd.n935 vdd.t916 8.126
R6262 vdd.n938 vdd.t337 8.126
R6263 vdd.n938 vdd.t1410 8.126
R6264 vdd.n939 vdd.t548 8.126
R6265 vdd.n939 vdd.t114 8.126
R6266 vdd.n940 vdd.t1108 8.126
R6267 vdd.n940 vdd.t690 8.126
R6268 vdd.n941 vdd.t881 8.126
R6269 vdd.n941 vdd.t453 8.126
R6270 vdd.n942 vdd.t748 8.126
R6271 vdd.n942 vdd.t310 8.126
R6272 vdd.n943 vdd.t1153 8.126
R6273 vdd.n943 vdd.t726 8.126
R6274 vdd.n944 vdd.t219 8.126
R6275 vdd.n944 vdd.t1280 8.126
R6276 vdd.n945 vdd.t350 8.126
R6277 vdd.n945 vdd.t1413 8.126
R6278 vdd.n946 vdd.t557 8.126
R6279 vdd.n946 vdd.t123 8.126
R6280 vdd.n947 vdd.t1117 8.126
R6281 vdd.n947 vdd.t694 8.126
R6282 vdd.n954 vdd.t111 8.126
R6283 vdd.n954 vdd.t492 8.126
R6284 vdd.n955 vdd.t316 8.126
R6285 vdd.n955 vdd.t696 8.126
R6286 vdd.n956 vdd.t886 8.126
R6287 vdd.n956 vdd.t1252 8.126
R6288 vdd.n957 vdd.t651 8.126
R6289 vdd.n957 vdd.t1025 8.126
R6290 vdd.n958 vdd.t514 8.126
R6291 vdd.n958 vdd.t888 8.126
R6292 vdd.n959 vdd.t919 8.126
R6293 vdd.n959 vdd.t1290 8.126
R6294 vdd.n960 vdd.t1476 8.126
R6295 vdd.n960 vdd.t361 8.126
R6296 vdd.n961 vdd.t117 8.126
R6297 vdd.n961 vdd.t496 8.126
R6298 vdd.n962 vdd.t323 8.126
R6299 vdd.n962 vdd.t705 8.126
R6300 vdd.n963 vdd.t890 8.126
R6301 vdd.n963 vdd.t1258 8.126
R6302 vdd.n966 vdd.t692 8.126
R6303 vdd.n966 vdd.t887 8.126
R6304 vdd.n967 vdd.t893 8.126
R6305 vdd.n967 vdd.t1095 8.126
R6306 vdd.n968 vdd.t1452 8.126
R6307 vdd.n968 vdd.t160 8.126
R6308 vdd.n969 vdd.t1219 8.126
R6309 vdd.n969 vdd.t1428 8.126
R6310 vdd.n970 vdd.t1091 8.126
R6311 vdd.n970 vdd.t1289 8.126
R6312 vdd.n971 vdd.t1487 8.126
R6313 vdd.n971 vdd.t196 8.126
R6314 vdd.n972 vdd.t567 8.126
R6315 vdd.n972 vdd.t776 8.126
R6316 vdd.n973 vdd.t700 8.126
R6317 vdd.n973 vdd.t897 8.126
R6318 vdd.n974 vdd.t900 8.126
R6319 vdd.n974 vdd.t1102 8.126
R6320 vdd.n975 vdd.t1457 8.126
R6321 vdd.n975 vdd.t168 8.126
R6322 vdd.n982 vdd.t462 8.126
R6323 vdd.n982 vdd.t658 8.126
R6324 vdd.n983 vdd.t661 8.126
R6325 vdd.n983 vdd.t868 8.126
R6326 vdd.n984 vdd.t1222 8.126
R6327 vdd.n984 vdd.t1430 8.126
R6328 vdd.n985 vdd.t996 8.126
R6329 vdd.n985 vdd.t1194 8.126
R6330 vdd.n986 vdd.t865 8.126
R6331 vdd.n986 vdd.t1068 8.126
R6332 vdd.n987 vdd.t1262 8.126
R6333 vdd.n987 vdd.t1462 8.126
R6334 vdd.n988 vdd.t333 8.126
R6335 vdd.n988 vdd.t533 8.126
R6336 vdd.n989 vdd.t467 8.126
R6337 vdd.n989 vdd.t664 8.126
R6338 vdd.n990 vdd.t671 8.126
R6339 vdd.n990 vdd.t874 8.126
R6340 vdd.n991 vdd.t1227 8.126
R6341 vdd.n991 vdd.t1435 8.126
R6342 vdd.n994 vdd.t864 8.126
R6343 vdd.n994 vdd.t1067 8.126
R6344 vdd.n995 vdd.t1071 8.126
R6345 vdd.n995 vdd.t1266 8.126
R6346 vdd.n996 vdd.t136 8.126
R6347 vdd.n996 vdd.t335 8.126
R6348 vdd.n997 vdd.t1403 8.126
R6349 vdd.n997 vdd.t100 8.126
R6350 vdd.n998 vdd.t1260 8.126
R6351 vdd.n998 vdd.t1459 8.126
R6352 vdd.n999 vdd.t172 8.126
R6353 vdd.n999 vdd.t377 8.126
R6354 vdd.n1000 vdd.t739 8.126
R6355 vdd.n1000 vdd.t936 8.126
R6356 vdd.n1001 vdd.t869 8.126
R6357 vdd.n1001 vdd.t1073 8.126
R6358 vdd.n1002 vdd.t1076 8.126
R6359 vdd.n1002 vdd.t1272 8.126
R6360 vdd.n1003 vdd.t142 8.126
R6361 vdd.n1003 vdd.t343 8.126
R6362 vdd.n1010 vdd.t1259 8.126
R6363 vdd.n1010 vdd.t833 8.126
R6364 vdd.n1011 vdd.t1465 8.126
R6365 vdd.n1011 vdd.t1037 8.126
R6366 vdd.n1012 vdd.t535 8.126
R6367 vdd.n1012 vdd.t105 8.126
R6368 vdd.n1013 vdd.t302 8.126
R6369 vdd.n1013 vdd.t1365 8.126
R6370 vdd.n1014 vdd.t169 8.126
R6371 vdd.n1014 vdd.t1229 8.126
R6372 vdd.n1015 vdd.t587 8.126
R6373 vdd.n1015 vdd.t145 8.126
R6374 vdd.n1016 vdd.t1138 8.126
R6375 vdd.n1016 vdd.t716 8.126
R6376 vdd.n1017 vdd.t1269 8.126
R6377 vdd.n1017 vdd.t840 8.126
R6378 vdd.n1018 vdd.t1470 8.126
R6379 vdd.n1018 vdd.t1051 8.126
R6380 vdd.n1019 vdd.t546 8.126
R6381 vdd.n1019 vdd.t112 8.126
R6382 vdd.n1022 vdd.t1033 8.126
R6383 vdd.n1022 vdd.t1409 8.126
R6384 vdd.n1023 vdd.t1232 8.126
R6385 vdd.n1023 vdd.t113 8.126
R6386 vdd.n1024 vdd.t305 8.126
R6387 vdd.n1024 vdd.t689 8.126
R6388 vdd.n1025 vdd.t69 8.126
R6389 vdd.n1025 vdd.t454 8.126
R6390 vdd.n1026 vdd.t1437 8.126
R6391 vdd.n1026 vdd.t311 8.126
R6392 vdd.n1027 vdd.t346 8.126
R6393 vdd.n1027 vdd.t727 8.126
R6394 vdd.n1028 vdd.t910 8.126
R6395 vdd.n1028 vdd.t1281 8.126
R6396 vdd.n1029 vdd.t1042 8.126
R6397 vdd.n1029 vdd.t1414 8.126
R6398 vdd.n1030 vdd.t1243 8.126
R6399 vdd.n1030 vdd.t122 8.126
R6400 vdd.n1031 vdd.t314 8.126
R6401 vdd.n1031 vdd.t693 8.126
R6402 vdd.n1038 vdd.t110 8.126
R6403 vdd.n1038 vdd.t1163 8.126
R6404 vdd.n1039 vdd.t315 8.126
R6405 vdd.n1039 vdd.t1376 8.126
R6406 vdd.n1040 vdd.t884 8.126
R6407 vdd.n1040 vdd.t459 8.126
R6408 vdd.n1041 vdd.t652 8.126
R6409 vdd.n1041 vdd.t201 8.126
R6410 vdd.n1042 vdd.t515 8.126
R6411 vdd.n1042 vdd.t74 8.126
R6412 vdd.n1043 vdd.t920 8.126
R6413 vdd.n1043 vdd.t495 8.126
R6414 vdd.n1044 vdd.t1477 8.126
R6415 vdd.n1044 vdd.t1063 8.126
R6416 vdd.n1045 vdd.t118 8.126
R6417 vdd.n1045 vdd.t1167 8.126
R6418 vdd.n1046 vdd.t322 8.126
R6419 vdd.n1046 vdd.t1386 8.126
R6420 vdd.n1047 vdd.t889 8.126
R6421 vdd.n1047 vdd.t464 8.126
R6422 vdd.n1050 vdd.t1371 8.126
R6423 vdd.n1050 vdd.t72 8.126
R6424 vdd.n1051 vdd.t77 8.126
R6425 vdd.n1051 vdd.t282 8.126
R6426 vdd.n1052 vdd.t655 8.126
R6427 vdd.n1052 vdd.t862 8.126
R6428 vdd.n1053 vdd.t409 8.126
R6429 vdd.n1053 vdd.t616 8.126
R6430 vdd.n1054 vdd.t280 8.126
R6431 vdd.n1054 vdd.t494 8.126
R6432 vdd.n1055 vdd.t697 8.126
R6433 vdd.n1055 vdd.t895 8.126
R6434 vdd.n1056 vdd.t1253 8.126
R6435 vdd.n1056 vdd.t1453 8.126
R6436 vdd.n1057 vdd.t1377 8.126
R6437 vdd.n1057 vdd.t79 8.126
R6438 vdd.n1058 vdd.t87 8.126
R6439 vdd.n1058 vdd.t291 8.126
R6440 vdd.n1059 vdd.t660 8.126
R6441 vdd.n1059 vdd.t867 8.126
R6442 vdd.n0 vdd.t278 8.126
R6443 vdd.n0 vdd.t493 8.126
R6444 vdd.n1 vdd.t497 8.126
R6445 vdd.n1 vdd.t701 8.126
R6446 vdd.n2 vdd.t1065 8.126
R6447 vdd.n2 vdd.t1254 8.126
R6448 vdd.n3 vdd.t827 8.126
R6449 vdd.n3 vdd.t1028 8.126
R6450 vdd.n4 vdd.t695 8.126
R6451 vdd.n4 vdd.t894 8.126
R6452 vdd.n5 vdd.t1096 8.126
R6453 vdd.n5 vdd.t1295 8.126
R6454 vdd.n6 vdd.t161 8.126
R6455 vdd.n6 vdd.t364 8.126
R6456 vdd.n7 vdd.t286 8.126
R6457 vdd.n7 vdd.t501 8.126
R6458 vdd.n8 vdd.t503 8.126
R6459 vdd.n8 vdd.t707 8.126
R6460 vdd.n9 vdd.t1069 8.126
R6461 vdd.n9 vdd.t1265 8.126
R6462 vdd.n594 vdd.t262 8.126
R6463 vdd.n594 vdd.t475 8.126
R6464 vdd.n595 vdd.t479 8.126
R6465 vdd.n595 vdd.t677 8.126
R6466 vdd.n596 vdd.t1038 8.126
R6467 vdd.n596 vdd.t1233 8.126
R6468 vdd.n597 vdd.t801 8.126
R6469 vdd.n597 vdd.t1003 8.126
R6470 vdd.n598 vdd.t674 8.126
R6471 vdd.n598 vdd.t875 8.126
R6472 vdd.n599 vdd.t1078 8.126
R6473 vdd.n599 vdd.t1274 8.126
R6474 vdd.n600 vdd.t147 8.126
R6475 vdd.n600 vdd.t349 8.126
R6476 vdd.n601 vdd.t270 8.126
R6477 vdd.n601 vdd.t484 8.126
R6478 vdd.n602 vdd.t489 8.126
R6479 vdd.n602 vdd.t687 8.126
R6480 vdd.n603 vdd.t1050 8.126
R6481 vdd.n603 vdd.t1241 8.126
R6482 vdd.n582 vdd.t673 8.126
R6483 vdd.n582 vdd.t1048 8.126
R6484 vdd.n583 vdd.t878 8.126
R6485 vdd.n583 vdd.t1245 8.126
R6486 vdd.n584 vdd.t1439 8.126
R6487 vdd.n584 vdd.t317 8.126
R6488 vdd.n585 vdd.t1200 8.126
R6489 vdd.n585 vdd.t73 8.126
R6490 vdd.n586 vdd.t1077 8.126
R6491 vdd.n586 vdd.t1444 8.126
R6492 vdd.n587 vdd.t1471 8.126
R6493 vdd.n587 vdd.t356 8.126
R6494 vdd.n588 vdd.t552 8.126
R6495 vdd.n588 vdd.t921 8.126
R6496 vdd.n589 vdd.t683 8.126
R6497 vdd.n589 vdd.t1056 8.126
R6498 vdd.n590 vdd.t882 8.126
R6499 vdd.n590 vdd.t1250 8.126
R6500 vdd.n591 vdd.t1445 8.126
R6501 vdd.n591 vdd.t321 8.126
R6502 vdd.n566 vdd.t1239 8.126
R6503 vdd.n566 vdd.t810 8.126
R6504 vdd.n567 vdd.t1446 8.126
R6505 vdd.n567 vdd.t1015 8.126
R6506 vdd.n568 vdd.t519 8.126
R6507 vdd.n568 vdd.t78 8.126
R6508 vdd.n569 vdd.t279 8.126
R6509 vdd.n569 vdd.t1335 8.126
R6510 vdd.n570 vdd.t153 8.126
R6511 vdd.n570 vdd.t1208 8.126
R6512 vdd.n571 vdd.t559 8.126
R6513 vdd.n571 vdd.t126 8.126
R6514 vdd.n572 vdd.t1121 8.126
R6515 vdd.n572 vdd.t698 8.126
R6516 vdd.n573 vdd.t1247 8.126
R6517 vdd.n573 vdd.t817 8.126
R6518 vdd.n574 vdd.t1449 8.126
R6519 vdd.n574 vdd.t1026 8.126
R6520 vdd.n575 vdd.t524 8.126
R6521 vdd.n575 vdd.t86 8.126
R6522 vdd.n554 vdd.t1011 8.126
R6523 vdd.n554 vdd.t1206 8.126
R6524 vdd.n555 vdd.t1211 8.126
R6525 vdd.n555 vdd.t1422 8.126
R6526 vdd.n556 vdd.t283 8.126
R6527 vdd.n556 vdd.t498 8.126
R6528 vdd.n557 vdd.t40 8.126
R6529 vdd.n557 vdd.t250 8.126
R6530 vdd.n558 vdd.t1420 8.126
R6531 vdd.n558 vdd.t125 8.126
R6532 vdd.n559 vdd.t325 8.126
R6533 vdd.n559 vdd.t527 8.126
R6534 vdd.n560 vdd.t896 8.126
R6535 vdd.n560 vdd.t1097 8.126
R6536 vdd.n561 vdd.t1020 8.126
R6537 vdd.n561 vdd.t1215 8.126
R6538 vdd.n562 vdd.t1221 8.126
R6539 vdd.n562 vdd.t1429 8.126
R6540 vdd.n563 vdd.t292 8.126
R6541 vdd.n563 vdd.t504 8.126
R6542 vdd.n22 vdd.t749 8.126
R6543 vdd.n22 vdd.t312 8.126
R6544 vdd.n23 vdd.t958 8.126
R6545 vdd.n23 vdd.t521 8.126
R6546 vdd.n24 vdd.t16 8.126
R6547 vdd.n24 vdd.t1086 8.126
R6548 vdd.n25 vdd.t1279 8.126
R6549 vdd.n25 vdd.t861 8.126
R6550 vdd.n26 vdd.t1152 8.126
R6551 vdd.n26 vdd.t725 8.126
R6552 vdd.n27 vdd.t68 8.126
R6553 vdd.n27 vdd.t1123 8.126
R6554 vdd.n28 vdd.t636 8.126
R6555 vdd.n28 vdd.t185 8.126
R6556 vdd.n29 vdd.t761 8.126
R6557 vdd.n29 vdd.t319 8.126
R6558 vdd.n30 vdd.t964 8.126
R6559 vdd.n30 vdd.t525 8.126
R6560 vdd.n31 vdd.t31 8.126
R6561 vdd.n31 vdd.t1094 8.126
R6562 vdd.n38 vdd.t340 8.126
R6563 vdd.n38 vdd.t544 8.126
R6564 vdd.n39 vdd.t551 8.126
R6565 vdd.n39 vdd.t758 8.126
R6566 vdd.n40 vdd.t1109 8.126
R6567 vdd.n40 vdd.t1314 8.126
R6568 vdd.n41 vdd.t883 8.126
R6569 vdd.n41 vdd.t1084 8.126
R6570 vdd.n42 vdd.t751 8.126
R6571 vdd.n42 vdd.t951 8.126
R6572 vdd.n43 vdd.t1156 8.126
R6573 vdd.n43 vdd.t1364 8.126
R6574 vdd.n44 vdd.t223 8.126
R6575 vdd.n44 vdd.t434 8.126
R6576 vdd.n45 vdd.t352 8.126
R6577 vdd.n45 vdd.t555 8.126
R6578 vdd.n46 vdd.t558 8.126
R6579 vdd.n46 vdd.t765 8.126
R6580 vdd.n47 vdd.t1118 8.126
R6581 vdd.n47 vdd.t1324 8.126
R6582 vdd.n50 vdd.t1434 8.126
R6583 vdd.n50 vdd.t140 8.126
R6584 vdd.n51 vdd.t146 8.126
R6585 vdd.n51 vdd.t348 8.126
R6586 vdd.n52 vdd.t717 8.126
R6587 vdd.n52 vdd.t911 8.126
R6588 vdd.n53 vdd.t490 8.126
R6589 vdd.n53 vdd.t688 8.126
R6590 vdd.n54 vdd.t342 8.126
R6591 vdd.n54 vdd.t545 8.126
R6592 vdd.n55 vdd.t755 8.126
R6593 vdd.n55 vdd.t955 8.126
R6594 vdd.n56 vdd.t1311 8.126
R6595 vdd.n56 vdd.t13 8.126
R6596 vdd.n57 vdd.t1441 8.126
R6597 vdd.n57 vdd.t150 8.126
R6598 vdd.n58 vdd.t154 8.126
R6599 vdd.n58 vdd.t355 8.126
R6600 vdd.n59 vdd.t723 8.126
R6601 vdd.n59 vdd.t917 8.126
R6602 vdd.n66 vdd.t167 8.126
R6603 vdd.n66 vdd.t371 8.126
R6604 vdd.n67 vdd.t379 8.126
R6605 vdd.n67 vdd.t589 8.126
R6606 vdd.n68 vdd.t938 8.126
R6607 vdd.n68 vdd.t1139 8.126
R6608 vdd.n69 vdd.t712 8.126
R6609 vdd.n69 vdd.t907 8.126
R6610 vdd.n70 vdd.t580 8.126
R6611 vdd.n70 vdd.t790 8.126
R6612 vdd.n71 vdd.t993 8.126
R6613 vdd.n71 vdd.t1192 8.126
R6614 vdd.n72 vdd.t51 8.126
R6615 vdd.n72 vdd.t261 8.126
R6616 vdd.n73 vdd.t174 8.126
R6617 vdd.n73 vdd.t380 8.126
R6618 vdd.n74 vdd.t383 8.126
R6619 vdd.n74 vdd.t592 8.126
R6620 vdd.n75 vdd.t947 8.126
R6621 vdd.n75 vdd.t1150 8.126
R6622 vdd.n78 vdd.t1092 8.126
R6623 vdd.n78 vdd.t1456 8.126
R6624 vdd.n79 vdd.t1298 8.126
R6625 vdd.n79 vdd.t173 8.126
R6626 vdd.n80 vdd.t366 8.126
R6627 vdd.n80 vdd.t740 8.126
R6628 vdd.n81 vdd.t134 8.126
R6629 vdd.n81 vdd.t509 8.126
R6630 vdd.n82 vdd.t1488 8.126
R6631 vdd.n82 vdd.t372 8.126
R6632 vdd.n83 vdd.t407 8.126
R6633 vdd.n83 vdd.t793 8.126
R6634 vdd.n84 vdd.t978 8.126
R6635 vdd.n84 vdd.t1346 8.126
R6636 vdd.n85 vdd.t1101 8.126
R6637 vdd.n85 vdd.t1464 8.126
R6638 vdd.n86 vdd.t1302 8.126
R6639 vdd.n86 vdd.t178 8.126
R6640 vdd.n87 vdd.t375 8.126
R6641 vdd.n87 vdd.t746 8.126
R6642 vdd.n94 vdd.t1320 8.126
R6643 vdd.n94 vdd.t24 8.126
R6644 vdd.n95 vdd.t34 8.126
R6645 vdd.n95 vdd.t244 8.126
R6646 vdd.n96 vdd.t600 8.126
R6647 vdd.n96 vdd.t811 8.126
R6648 vdd.n97 vdd.t362 8.126
R6649 vdd.n97 vdd.t568 8.126
R6650 vdd.n98 vdd.t238 8.126
R6651 vdd.n98 vdd.t449 8.126
R6652 vdd.n99 vdd.t650 8.126
R6653 vdd.n99 vdd.t859 8.126
R6654 vdd.n100 vdd.t1209 8.126
R6655 vdd.n100 vdd.t1419 8.126
R6656 vdd.n101 vdd.t1330 8.126
R6657 vdd.n101 vdd.t35 8.126
R6658 vdd.n102 vdd.t39 8.126
R6659 vdd.n102 vdd.t248 8.126
R6660 vdd.n103 vdd.t612 8.126
R6661 vdd.n103 vdd.t824 8.126
R6662 vdd.n106 vdd.t915 8.126
R6663 vdd.n106 vdd.t1114 8.126
R6664 vdd.n107 vdd.t1122 8.126
R6665 vdd.n107 vdd.t1328 8.126
R6666 vdd.n108 vdd.t184 8.126
R6667 vdd.n108 vdd.t390 8.126
R6668 vdd.n109 vdd.t1450 8.126
R6669 vdd.n109 vdd.t159 8.126
R6670 vdd.n110 vdd.t1323 8.126
R6671 vdd.n110 vdd.t28 8.126
R6672 vdd.n111 vdd.t240 8.126
R6673 vdd.n111 vdd.t452 8.126
R6674 vdd.n112 vdd.t809 8.126
R6675 vdd.n112 vdd.t1012 8.126
R6676 vdd.n113 vdd.t925 8.126
R6677 vdd.n113 vdd.t1125 8.126
R6678 vdd.n114 vdd.t1127 8.126
R6679 vdd.n114 vdd.t1334 8.126
R6680 vdd.n115 vdd.t194 8.126
R6681 vdd.n115 vdd.t402 8.126
R6682 vdd.n122 vdd.t1144 8.126
R6683 vdd.n122 vdd.t721 8.126
R6684 vdd.n123 vdd.t1362 8.126
R6685 vdd.n123 vdd.t922 8.126
R6686 vdd.n124 vdd.t431 8.126
R6687 vdd.n124 vdd.t1478 8.126
R6688 vdd.n125 vdd.t180 8.126
R6689 vdd.n125 vdd.t1251 8.126
R6690 vdd.n126 vdd.t59 8.126
R6691 vdd.n126 vdd.t1116 8.126
R6692 vdd.n127 vdd.t486 8.126
R6693 vdd.n127 vdd.t30 8.126
R6694 vdd.n128 vdd.t1047 8.126
R6695 vdd.n128 vdd.t599 8.126
R6696 vdd.n129 vdd.t1157 8.126
R6697 vdd.n129 vdd.t729 8.126
R6698 vdd.n130 vdd.t1369 8.126
R6699 vdd.n130 vdd.t927 8.126
R6700 vdd.n131 vdd.t444 8.126
R6701 vdd.n131 vdd.t1485 8.126
R6702 vdd.n134 vdd.t743 8.126
R6703 vdd.n134 vdd.t943 8.126
R6704 vdd.n135 vdd.t953 8.126
R6705 vdd.n135 vdd.t1154 8.126
R6706 vdd.n136 vdd.t10 8.126
R6707 vdd.n136 vdd.t220 8.126
R6708 vdd.n137 vdd.t1276 8.126
R6709 vdd.n137 vdd.t1473 8.126
R6710 vdd.n138 vdd.t1145 8.126
R6711 vdd.n138 vdd.t1353 8.126
R6712 vdd.n139 vdd.t63 8.126
R6713 vdd.n139 vdd.t273 8.126
R6714 vdd.n140 vdd.t631 8.126
R6715 vdd.n140 vdd.t845 8.126
R6716 vdd.n141 vdd.t756 8.126
R6717 vdd.n141 vdd.t956 8.126
R6718 vdd.n142 vdd.t961 8.126
R6719 vdd.n142 vdd.t1161 8.126
R6720 vdd.n143 vdd.t20 8.126
R6721 vdd.n143 vdd.t232 8.126
R6722 vdd.n150 vdd.t166 8.126
R6723 vdd.n150 vdd.t537 8.126
R6724 vdd.n151 vdd.t378 8.126
R6725 vdd.n151 vdd.t750 8.126
R6726 vdd.n152 vdd.t937 8.126
R6727 vdd.n152 vdd.t1309 8.126
R6728 vdd.n153 vdd.t713 8.126
R6729 vdd.n153 vdd.t1081 8.126
R6730 vdd.n154 vdd.t583 8.126
R6731 vdd.n154 vdd.t944 8.126
R6732 vdd.n155 vdd.t994 8.126
R6733 vdd.n155 vdd.t1358 8.126
R6734 vdd.n156 vdd.t52 8.126
R6735 vdd.n156 vdd.t427 8.126
R6736 vdd.n157 vdd.t175 8.126
R6737 vdd.n157 vdd.t549 8.126
R6738 vdd.n158 vdd.t384 8.126
R6739 vdd.n158 vdd.t762 8.126
R6740 vdd.n159 vdd.t948 8.126
R6741 vdd.n159 vdd.t1317 8.126
R6742 vdd.n162 vdd.t395 8.126
R6743 vdd.n162 vdd.t605 8.126
R6744 vdd.n163 vdd.t614 8.126
R6745 vdd.n163 vdd.t826 8.126
R6746 vdd.n164 vdd.t1176 8.126
R6747 vdd.n164 vdd.t1387 8.126
R6748 vdd.n165 vdd.t931 8.126
R6749 vdd.n165 vdd.t1131 8.126
R6750 vdd.n166 vdd.t820 8.126
R6751 vdd.n166 vdd.t1021 8.126
R6752 vdd.n167 vdd.t1217 8.126
R6753 vdd.n167 vdd.t1427 8.126
R6754 vdd.n168 vdd.t288 8.126
R6755 vdd.n168 vdd.t502 8.126
R6756 vdd.n169 vdd.t408 8.126
R6757 vdd.n169 vdd.t617 8.126
R6758 vdd.n170 vdd.t619 8.126
R6759 vdd.n170 vdd.t830 8.126
R6760 vdd.n171 vdd.t1186 8.126
R6761 vdd.n171 vdd.t1398 8.126
R6762 vdd.n178 vdd.t1482 8.126
R6763 vdd.n178 vdd.t189 8.126
R6764 vdd.n179 vdd.t198 8.126
R6765 vdd.n179 vdd.t405 8.126
R6766 vdd.n180 vdd.t778 8.126
R6767 vdd.n180 vdd.t976 8.126
R6768 vdd.n181 vdd.t529 8.126
R6769 vdd.n181 vdd.t736 8.126
R6770 vdd.n182 vdd.t396 8.126
R6771 vdd.n182 vdd.t606 8.126
R6772 vdd.n183 vdd.t822 8.126
R6773 vdd.n183 vdd.t1023 8.126
R6774 vdd.n184 vdd.t1381 8.126
R6775 vdd.n184 vdd.t83 8.126
R6776 vdd.n185 vdd.t1493 8.126
R6777 vdd.n185 vdd.t200 8.126
R6778 vdd.n186 vdd.t205 8.126
R6779 vdd.n186 vdd.t413 8.126
R6780 vdd.n187 vdd.t786 8.126
R6781 vdd.n187 vdd.t988 8.126
R6782 vdd.n190 vdd.t227 8.126
R6783 vdd.n190 vdd.t1286 8.126
R6784 vdd.n191 vdd.t448 8.126
R6785 vdd.n191 vdd.t1491 8.126
R6786 vdd.n192 vdd.t1009 8.126
R6787 vdd.n192 vdd.t571 8.126
R6788 vdd.n193 vdd.t769 8.126
R6789 vdd.n193 vdd.t329 8.126
R6790 vdd.n194 vdd.t641 8.126
R6791 vdd.n194 vdd.t190 8.126
R6792 vdd.n195 vdd.t1058 8.126
R6793 vdd.n195 vdd.t610 8.126
R6794 vdd.n196 vdd.t120 8.126
R6795 vdd.n196 vdd.t1171 8.126
R6796 vdd.n197 vdd.t241 8.126
R6797 vdd.n197 vdd.t1294 8.126
R6798 vdd.n198 vdd.t458 8.126
R6799 vdd.n198 vdd.t1498 8.126
R6800 vdd.n199 vdd.t1017 8.126
R6801 vdd.n199 vdd.t578 8.126
R6802 vdd.n206 vdd.t1313 8.126
R6803 vdd.n206 vdd.t15 8.126
R6804 vdd.n207 vdd.t27 8.126
R6805 vdd.n207 vdd.t237 8.126
R6806 vdd.n208 vdd.t597 8.126
R6807 vdd.n208 vdd.t807 8.126
R6808 vdd.n209 vdd.t357 8.126
R6809 vdd.n209 vdd.t562 8.126
R6810 vdd.n210 vdd.t229 8.126
R6811 vdd.n210 vdd.t439 8.126
R6812 vdd.n211 vdd.t644 8.126
R6813 vdd.n211 vdd.t855 8.126
R6814 vdd.n212 vdd.t1203 8.126
R6815 vdd.n212 vdd.t1416 8.126
R6816 vdd.n213 vdd.t1326 8.126
R6817 vdd.n213 vdd.t32 8.126
R6818 vdd.n214 vdd.t36 8.126
R6819 vdd.n214 vdd.t245 8.126
R6820 vdd.n215 vdd.t603 8.126
R6821 vdd.n215 vdd.t815 8.126
R6822 vdd.n218 vdd.t1392 8.126
R6823 vdd.n218 vdd.t1110 8.126
R6824 vdd.n219 vdd.t99 8.126
R6825 vdd.n219 vdd.t1322 8.126
R6826 vdd.n220 vdd.t672 8.126
R6827 vdd.n220 vdd.t387 8.126
R6828 vdd.n221 vdd.t423 8.126
R6829 vdd.n221 vdd.t156 8.126
R6830 vdd.n222 vdd.t296 8.126
R6831 vdd.n222 vdd.t18 8.126
R6832 vdd.n223 vdd.t711 8.126
R6833 vdd.n223 vdd.t443 8.126
R6834 vdd.n224 vdd.t1271 8.126
R6835 vdd.n224 vdd.t1006 8.126
R6836 vdd.n225 vdd.t1402 8.126
R6837 vdd.n225 vdd.t1120 8.126
R6838 vdd.n226 vdd.t104 8.126
R6839 vdd.n226 vdd.t1331 8.126
R6840 vdd.n227 vdd.t681 8.126
R6841 vdd.n227 vdd.t394 8.126
R6842 vdd.n234 vdd.t983 8.126
R6843 vdd.n234 vdd.t1182 8.126
R6844 vdd.n235 vdd.t1191 8.126
R6845 vdd.n235 vdd.t1401 8.126
R6846 vdd.n236 vdd.t260 8.126
R6847 vdd.n236 vdd.t474 8.126
R6848 vdd.n237 vdd.t4 8.126
R6849 vdd.n237 vdd.t214 8.126
R6850 vdd.n238 vdd.t1393 8.126
R6851 vdd.n238 vdd.t92 8.126
R6852 vdd.n239 vdd.t298 8.126
R6853 vdd.n239 vdd.t507 8.126
R6854 vdd.n240 vdd.t872 8.126
R6855 vdd.n240 vdd.t1075 8.126
R6856 vdd.n241 vdd.t995 8.126
R6857 vdd.n241 vdd.t1193 8.126
R6858 vdd.n242 vdd.t1195 8.126
R6859 vdd.n242 vdd.t1405 8.126
R6860 vdd.n243 vdd.t267 8.126
R6861 vdd.n243 vdd.t481 8.126
R6862 vdd.n246 vdd.t573 8.126
R6863 vdd.n246 vdd.t781 8.126
R6864 vdd.n247 vdd.t789 8.126
R6865 vdd.n247 vdd.t992 8.126
R6866 vdd.n248 vdd.t1343 8.126
R6867 vdd.n248 vdd.t48 8.126
R6868 vdd.n249 vdd.t1105 8.126
R6869 vdd.n249 vdd.t1306 8.126
R6870 vdd.n250 vdd.t984 8.126
R6871 vdd.n250 vdd.t1183 8.126
R6872 vdd.n251 vdd.t1397 8.126
R6873 vdd.n251 vdd.t95 8.126
R6874 vdd.n252 vdd.t472 8.126
R6875 vdd.n252 vdd.t670 8.126
R6876 vdd.n253 vdd.t586 8.126
R6877 vdd.n253 vdd.t794 8.126
R6878 vdd.n254 vdd.t796 8.126
R6879 vdd.n254 vdd.t998 8.126
R6880 vdd.n255 vdd.t1351 8.126
R6881 vdd.n255 vdd.t57 8.126
R6882 vdd.n262 vdd.t188 8.126
R6883 vdd.n262 vdd.t398 8.126
R6884 vdd.n263 vdd.t406 8.126
R6885 vdd.n263 vdd.t615 8.126
R6886 vdd.n264 vdd.t977 8.126
R6887 vdd.n264 vdd.t1177 8.126
R6888 vdd.n265 vdd.t737 8.126
R6889 vdd.n265 vdd.t933 8.126
R6890 vdd.n266 vdd.t608 8.126
R6891 vdd.n266 vdd.t819 8.126
R6892 vdd.n267 vdd.t1024 8.126
R6893 vdd.n267 vdd.t1218 8.126
R6894 vdd.n268 vdd.t84 8.126
R6895 vdd.n268 vdd.t289 8.126
R6896 vdd.n269 vdd.t202 8.126
R6897 vdd.n269 vdd.t410 8.126
R6898 vdd.n270 vdd.t414 8.126
R6899 vdd.n270 vdd.t620 8.126
R6900 vdd.n271 vdd.t989 8.126
R6901 vdd.n271 vdd.t1187 8.126
R6902 vdd.n274 vdd.t1285 8.126
R6903 vdd.n274 vdd.t1481 8.126
R6904 vdd.n275 vdd.t1490 8.126
R6905 vdd.n275 vdd.t197 8.126
R6906 vdd.n276 vdd.t570 8.126
R6907 vdd.n276 vdd.t777 8.126
R6908 vdd.n277 vdd.t330 8.126
R6909 vdd.n277 vdd.t530 8.126
R6910 vdd.n278 vdd.t192 8.126
R6911 vdd.n278 vdd.t399 8.126
R6912 vdd.n279 vdd.t611 8.126
R6913 vdd.n279 vdd.t823 8.126
R6914 vdd.n280 vdd.t1173 8.126
R6915 vdd.n280 vdd.t1383 8.126
R6916 vdd.n281 vdd.t1296 8.126
R6917 vdd.n281 vdd.t1494 8.126
R6918 vdd.n282 vdd.t1499 8.126
R6919 vdd.n282 vdd.t206 8.126
R6920 vdd.n283 vdd.t579 8.126
R6921 vdd.n283 vdd.t787 8.126
R6922 vdd.n290 vdd.t1355 8.126
R6923 vdd.n290 vdd.t1087 8.126
R6924 vdd.n291 vdd.t67 8.126
R6925 vdd.n291 vdd.t1291 8.126
R6926 vdd.n292 vdd.t635 8.126
R6927 vdd.n292 vdd.t363 8.126
R6928 vdd.n293 vdd.t388 8.126
R6929 vdd.n293 vdd.t132 8.126
R6930 vdd.n294 vdd.t272 8.126
R6931 vdd.n294 vdd.t1484 8.126
R6932 vdd.n295 vdd.t684 8.126
R6933 vdd.n295 vdd.t401 8.126
R6934 vdd.n296 vdd.t1240 8.126
R6935 vdd.n296 vdd.t972 8.126
R6936 vdd.n297 vdd.t1366 8.126
R6937 vdd.n297 vdd.t1098 8.126
R6938 vdd.n298 vdd.t71 8.126
R6939 vdd.n298 vdd.t1301 8.126
R6940 vdd.n299 vdd.t647 8.126
R6941 vdd.n299 vdd.t370 8.126
R6942 vdd.n302 vdd.t945 8.126
R6943 vdd.n302 vdd.t1147 8.126
R6944 vdd.n303 vdd.t1155 8.126
R6945 vdd.n303 vdd.t1363 8.126
R6946 vdd.n304 vdd.t222 8.126
R6947 vdd.n304 vdd.t433 8.126
R6948 vdd.n305 vdd.t1474 8.126
R6949 vdd.n305 vdd.t182 8.126
R6950 vdd.n306 vdd.t1356 8.126
R6951 vdd.n306 vdd.t61 8.126
R6952 vdd.n307 vdd.t274 8.126
R6953 vdd.n307 vdd.t487 8.126
R6954 vdd.n308 vdd.t846 8.126
R6955 vdd.n308 vdd.t1049 8.126
R6956 vdd.n309 vdd.t957 8.126
R6957 vdd.n309 vdd.t1158 8.126
R6958 vdd.n310 vdd.t1162 8.126
R6959 vdd.n310 vdd.t1370 8.126
R6960 vdd.n311 vdd.t234 8.126
R6961 vdd.n311 vdd.t446 8.126
R6962 vdd.n318 vdd.t538 8.126
R6963 vdd.n318 vdd.t745 8.126
R6964 vdd.n319 vdd.t753 8.126
R6965 vdd.n319 vdd.t954 8.126
R6966 vdd.n320 vdd.t1310 8.126
R6967 vdd.n320 vdd.t12 8.126
R6968 vdd.n321 vdd.t1082 8.126
R6969 vdd.n321 vdd.t1277 8.126
R6970 vdd.n322 vdd.t946 8.126
R6971 vdd.n322 vdd.t1148 8.126
R6972 vdd.n323 vdd.t1359 8.126
R6973 vdd.n323 vdd.t64 8.126
R6974 vdd.n324 vdd.t428 8.126
R6975 vdd.n324 vdd.t632 8.126
R6976 vdd.n325 vdd.t550 8.126
R6977 vdd.n325 vdd.t757 8.126
R6978 vdd.n326 vdd.t763 8.126
R6979 vdd.n326 vdd.t962 8.126
R6980 vdd.n327 vdd.t1319 8.126
R6981 vdd.n327 vdd.t23 8.126
R6982 vdd.n330 vdd.t783 8.126
R6983 vdd.n330 vdd.t982 8.126
R6984 vdd.n331 vdd.t991 8.126
R6985 vdd.n331 vdd.t1190 8.126
R6986 vdd.n332 vdd.t50 8.126
R6987 vdd.n332 vdd.t259 8.126
R6988 vdd.n333 vdd.t1305 8.126
R6989 vdd.n333 vdd.t5 8.126
R6990 vdd.n334 vdd.t1184 8.126
R6991 vdd.n334 vdd.t1394 8.126
R6992 vdd.n335 vdd.t96 8.126
R6993 vdd.n335 vdd.t299 8.126
R6994 vdd.n336 vdd.t669 8.126
R6995 vdd.n336 vdd.t873 8.126
R6996 vdd.n337 vdd.t795 8.126
R6997 vdd.n337 vdd.t997 8.126
R6998 vdd.n338 vdd.t999 8.126
R6999 vdd.n338 vdd.t1196 8.126
R7000 vdd.n339 vdd.t58 8.126
R7001 vdd.n339 vdd.t269 8.126
R7002 vdd.n346 vdd.t367 8.126
R7003 vdd.n346 vdd.t575 8.126
R7004 vdd.n347 vdd.t585 8.126
R7005 vdd.n347 vdd.t792 8.126
R7006 vdd.n348 vdd.t1136 8.126
R7007 vdd.n348 vdd.t1345 8.126
R7008 vdd.n349 vdd.t905 8.126
R7009 vdd.n349 vdd.t1104 8.126
R7010 vdd.n350 vdd.t784 8.126
R7011 vdd.n350 vdd.t986 8.126
R7012 vdd.n351 vdd.t1185 8.126
R7013 vdd.n351 vdd.t1396 8.126
R7014 vdd.n352 vdd.t256 8.126
R7015 vdd.n352 vdd.t471 8.126
R7016 vdd.n353 vdd.t376 8.126
R7017 vdd.n353 vdd.t588 8.126
R7018 vdd.n354 vdd.t590 8.126
R7019 vdd.n354 vdd.t797 8.126
R7020 vdd.n355 vdd.t1143 8.126
R7021 vdd.n355 vdd.t1352 8.126
R7022 vdd.n358 vdd.t440 8.126
R7023 vdd.n358 vdd.t162 8.126
R7024 vdd.n359 vdd.t649 8.126
R7025 vdd.n359 vdd.t374 8.126
R7026 vdd.n360 vdd.t1207 8.126
R7027 vdd.n360 vdd.t934 8.126
R7028 vdd.n361 vdd.t970 8.126
R7029 vdd.n361 vdd.t710 8.126
R7030 vdd.n362 vdd.t853 8.126
R7031 vdd.n362 vdd.t576 8.126
R7032 vdd.n363 vdd.t1248 8.126
R7033 vdd.n363 vdd.t987 8.126
R7034 vdd.n364 vdd.t320 8.126
R7035 vdd.n364 vdd.t46 8.126
R7036 vdd.n365 vdd.t455 8.126
R7037 vdd.n365 vdd.t171 8.126
R7038 vdd.n366 vdd.t656 8.126
R7039 vdd.n366 vdd.t381 8.126
R7040 vdd.n367 vdd.t1214 8.126
R7041 vdd.n367 vdd.t941 8.126
R7042 vdd.n374 vdd.t17 8.126
R7043 vdd.n374 vdd.t228 8.126
R7044 vdd.n375 vdd.t239 8.126
R7045 vdd.n375 vdd.t451 8.126
R7046 vdd.n376 vdd.t808 8.126
R7047 vdd.n376 vdd.t1010 8.126
R7048 vdd.n377 vdd.t563 8.126
R7049 vdd.n377 vdd.t771 8.126
R7050 vdd.n378 vdd.t442 8.126
R7051 vdd.n378 vdd.t643 8.126
R7052 vdd.n379 vdd.t856 8.126
R7053 vdd.n379 vdd.t1059 8.126
R7054 vdd.n380 vdd.t1417 8.126
R7055 vdd.n380 vdd.t121 8.126
R7056 vdd.n381 vdd.t33 8.126
R7057 vdd.n381 vdd.t242 8.126
R7058 vdd.n382 vdd.t246 8.126
R7059 vdd.n382 vdd.t460 8.126
R7060 vdd.n383 vdd.t816 8.126
R7061 vdd.n383 vdd.t1018 8.126
R7062 vdd.n386 vdd.t264 8.126
R7063 vdd.n386 vdd.t1315 8.126
R7064 vdd.n387 vdd.t485 8.126
R7065 vdd.n387 vdd.t29 8.126
R7066 vdd.n388 vdd.t1045 8.126
R7067 vdd.n388 vdd.t598 8.126
R7068 vdd.n389 vdd.t803 8.126
R7069 vdd.n389 vdd.t358 8.126
R7070 vdd.n390 vdd.t679 8.126
R7071 vdd.n390 vdd.t231 8.126
R7072 vdd.n391 vdd.t1079 8.126
R7073 vdd.n391 vdd.t646 8.126
R7074 vdd.n392 vdd.t151 8.126
R7075 vdd.n392 vdd.t1205 8.126
R7076 vdd.n393 vdd.t276 8.126
R7077 vdd.n393 vdd.t1327 8.126
R7078 vdd.n394 vdd.t491 8.126
R7079 vdd.n394 vdd.t37 8.126
R7080 vdd.n395 vdd.t1055 8.126
R7081 vdd.n395 vdd.t604 8.126
R7082 vdd.n402 vdd.t1348 8.126
R7083 vdd.n402 vdd.t54 8.126
R7084 vdd.n403 vdd.t62 8.126
R7085 vdd.n403 vdd.t271 8.126
R7086 vdd.n404 vdd.t630 8.126
R7087 vdd.n404 vdd.t844 8.126
R7088 vdd.n405 vdd.t385 8.126
R7089 vdd.n405 vdd.t594 8.126
R7090 vdd.n406 vdd.t265 8.126
R7091 vdd.n406 vdd.t478 8.126
R7092 vdd.n407 vdd.t680 8.126
R7093 vdd.n407 vdd.t879 8.126
R7094 vdd.n408 vdd.t1236 8.126
R7095 vdd.n408 vdd.t1442 8.126
R7096 vdd.n409 vdd.t1360 8.126
R7097 vdd.n409 vdd.t66 8.126
R7098 vdd.n410 vdd.t70 8.126
R7099 vdd.n410 vdd.t277 8.126
R7100 vdd.n411 vdd.t640 8.126
R7101 vdd.n411 vdd.t852 8.126
R7102 vdd.n414 vdd.t939 8.126
R7103 vdd.n414 vdd.t1140 8.126
R7104 vdd.n415 vdd.t1149 8.126
R7105 vdd.n415 vdd.t1357 8.126
R7106 vdd.n416 vdd.t216 8.126
R7107 vdd.n416 vdd.t426 8.126
R7108 vdd.n417 vdd.t1472 8.126
R7109 vdd.n417 vdd.t179 8.126
R7110 vdd.n418 vdd.t1349 8.126
R7111 vdd.n418 vdd.t55 8.126
R7112 vdd.n419 vdd.t266 8.126
R7113 vdd.n419 vdd.t480 8.126
R7114 vdd.n420 vdd.t838 8.126
R7115 vdd.n420 vdd.t1040 8.126
R7116 vdd.n421 vdd.t950 8.126
R7117 vdd.n421 vdd.t1151 8.126
R7118 vdd.n422 vdd.t1159 8.126
R7119 vdd.n422 vdd.t1367 8.126
R7120 vdd.n423 vdd.t226 8.126
R7121 vdd.n423 vdd.t438 8.126
R7122 vdd.n430 vdd.t1014 8.126
R7123 vdd.n430 vdd.t1388 8.126
R7124 vdd.n431 vdd.t1216 8.126
R7125 vdd.n431 vdd.t93 8.126
R7126 vdd.n432 vdd.t287 8.126
R7127 vdd.n432 vdd.t666 8.126
R7128 vdd.n433 vdd.t45 8.126
R7129 vdd.n433 vdd.t419 8.126
R7130 vdd.n434 vdd.t1423 8.126
R7131 vdd.n434 vdd.t294 8.126
R7132 vdd.n435 vdd.t327 8.126
R7133 vdd.n435 vdd.t709 8.126
R7134 vdd.n436 vdd.t899 8.126
R7135 vdd.n436 vdd.t1268 8.126
R7136 vdd.n437 vdd.t1027 8.126
R7137 vdd.n437 vdd.t1399 8.126
R7138 vdd.n438 vdd.t1223 8.126
R7139 vdd.n438 vdd.t101 8.126
R7140 vdd.n439 vdd.t295 8.126
R7141 vdd.n439 vdd.t676 8.126
R7142 vdd.n442 vdd.t601 8.126
R7143 vdd.n442 vdd.t813 8.126
R7144 vdd.n443 vdd.t821 8.126
R7145 vdd.n443 vdd.t1022 8.126
R7146 vdd.n444 vdd.t1380 8.126
R7147 vdd.n444 vdd.t82 8.126
R7148 vdd.n445 vdd.t1130 8.126
R7149 vdd.n445 vdd.t1340 8.126
R7150 vdd.n446 vdd.t1016 8.126
R7151 vdd.n446 vdd.t1212 8.126
R7152 vdd.n447 vdd.t1424 8.126
R7153 vdd.n447 vdd.t129 8.126
R7154 vdd.n448 vdd.t500 8.126
R7155 vdd.n448 vdd.t704 8.126
R7156 vdd.n449 vdd.t613 8.126
R7157 vdd.n449 vdd.t825 8.126
R7158 vdd.n450 vdd.t828 8.126
R7159 vdd.n450 vdd.t1029 8.126
R7160 vdd.n451 vdd.t1391 8.126
R7161 vdd.n451 vdd.t91 8.126
R7162 vdd.n458 vdd.t848 8.126
R7163 vdd.n458 vdd.t392 8.126
R7164 vdd.n459 vdd.t1057 8.126
R7165 vdd.n459 vdd.t609 8.126
R7166 vdd.n460 vdd.t119 8.126
R7167 vdd.n460 vdd.t1170 8.126
R7168 vdd.n461 vdd.t1374 8.126
R7169 vdd.n461 vdd.t930 8.126
R7170 vdd.n462 vdd.t1244 8.126
R7171 vdd.n462 vdd.t814 8.126
R7172 vdd.n463 vdd.t155 8.126
R7173 vdd.n463 vdd.t1213 8.126
R7174 vdd.n464 vdd.t730 8.126
R7175 vdd.n464 vdd.t285 8.126
R7176 vdd.n465 vdd.t858 8.126
R7177 vdd.n465 vdd.t404 8.126
R7178 vdd.n466 vdd.t1061 8.126
R7179 vdd.n466 vdd.t618 8.126
R7180 vdd.n467 vdd.t127 8.126
R7181 vdd.n467 vdd.t1181 8.126
R7182 vdd.n470 vdd.t432 8.126
R7183 vdd.n470 vdd.t637 8.126
R7184 vdd.n471 vdd.t642 8.126
R7185 vdd.n471 vdd.t854 8.126
R7186 vdd.n472 vdd.t1202 8.126
R7187 vdd.n472 vdd.t1415 8.126
R7188 vdd.n473 vdd.t967 8.126
R7189 vdd.n473 vdd.t1166 8.126
R7190 vdd.n474 vdd.t849 8.126
R7191 vdd.n474 vdd.t1052 8.126
R7192 vdd.n475 vdd.t1246 8.126
R7193 vdd.n475 vdd.t1447 8.126
R7194 vdd.n476 vdd.t318 8.126
R7195 vdd.n476 vdd.t520 8.126
R7196 vdd.n477 vdd.t447 8.126
R7197 vdd.n477 vdd.t648 8.126
R7198 vdd.n478 vdd.t653 8.126
R7199 vdd.n478 vdd.t860 8.126
R7200 vdd.n479 vdd.t1210 8.126
R7201 vdd.n479 vdd.t1421 8.126
R7202 vdd.n486 vdd.t11 8.126
R7203 vdd.n486 vdd.t221 8.126
R7204 vdd.n487 vdd.t230 8.126
R7205 vdd.n487 vdd.t441 8.126
R7206 vdd.n488 vdd.t804 8.126
R7207 vdd.n488 vdd.t1005 8.126
R7208 vdd.n489 vdd.t561 8.126
R7209 vdd.n489 vdd.t767 8.126
R7210 vdd.n490 vdd.t435 8.126
R7211 vdd.n490 vdd.t638 8.126
R7212 vdd.n491 vdd.t851 8.126
R7213 vdd.n491 vdd.t1054 8.126
R7214 vdd.n492 vdd.t1411 8.126
R7215 vdd.n492 vdd.t116 8.126
R7216 vdd.n493 vdd.t26 8.126
R7217 vdd.n493 vdd.t236 8.126
R7218 vdd.n494 vdd.t243 8.126
R7219 vdd.n494 vdd.t456 8.126
R7220 vdd.n495 vdd.t812 8.126
R7221 vdd.n495 vdd.t1013 8.126
R7222 vdd.n498 vdd.t88 8.126
R7223 vdd.n498 vdd.t476 8.126
R7224 vdd.n499 vdd.t297 8.126
R7225 vdd.n499 vdd.t678 8.126
R7226 vdd.n500 vdd.t871 8.126
R7227 vdd.n500 vdd.t1234 8.126
R7228 vdd.n501 vdd.t624 8.126
R7229 vdd.n501 vdd.t1002 8.126
R7230 vdd.n502 vdd.t505 8.126
R7231 vdd.n502 vdd.t876 8.126
R7232 vdd.n503 vdd.t904 8.126
R7233 vdd.n503 vdd.t1273 8.126
R7234 vdd.n504 vdd.t1466 8.126
R7235 vdd.n504 vdd.t347 8.126
R7236 vdd.n505 vdd.t98 8.126
R7237 vdd.n505 vdd.t483 8.126
R7238 vdd.n506 vdd.t304 8.126
R7239 vdd.n506 vdd.t686 8.126
R7240 vdd.n507 vdd.t877 8.126
R7241 vdd.n507 vdd.t1242 8.126
R7242 vdd.n513 vdd.t1178 8.126
R7243 vdd.n513 vdd.t1389 8.126
R7244 vdd.n514 vdd.t1395 8.126
R7245 vdd.n514 vdd.t94 8.126
R7246 vdd.n515 vdd.t470 8.126
R7247 vdd.n515 vdd.t668 8.126
R7248 vdd.n516 vdd.t209 8.126
R7249 vdd.n516 vdd.t418 8.126
R7250 vdd.n517 vdd.t89 8.126
R7251 vdd.n517 vdd.t293 8.126
R7252 vdd.n518 vdd.t506 8.126
R7253 vdd.n518 vdd.t708 8.126
R7254 vdd.n519 vdd.t1072 8.126
R7255 vdd.n519 vdd.t1267 8.126
R7256 vdd.n520 vdd.t1188 8.126
R7257 vdd.n520 vdd.t1400 8.126
R7258 vdd.n521 vdd.t1404 8.126
R7259 vdd.n521 vdd.t102 8.126
R7260 vdd.n522 vdd.t477 8.126
R7261 vdd.n522 vdd.t675 8.126
R7262 vdd.n540 vdd.t1418 8.126
R7263 vdd.n540 vdd.t124 8.126
R7264 vdd.n541 vdd.t128 8.126
R7265 vdd.n541 vdd.t326 8.126
R7266 vdd.n542 vdd.t702 8.126
R7267 vdd.n542 vdd.t898 8.126
R7268 vdd.n543 vdd.t465 8.126
R7269 vdd.n543 vdd.t662 8.126
R7270 vdd.n544 vdd.t324 8.126
R7271 vdd.n544 vdd.t526 8.126
R7272 vdd.n545 vdd.t734 8.126
R7273 vdd.n545 vdd.t928 8.126
R7274 vdd.n546 vdd.t1297 8.126
R7275 vdd.n546 vdd.t1495 8.126
R7276 vdd.n547 vdd.t1426 8.126
R7277 vdd.n547 vdd.t131 8.126
R7278 vdd.n548 vdd.t133 8.126
R7279 vdd.n548 vdd.t332 8.126
R7280 vdd.n549 vdd.t706 8.126
R7281 vdd.n549 vdd.t903 8.126
R7282 vdd.n533 vdd.n532 7.5
R7283 vdd.n527 vdd.n526 3.75
R7284 vdd.n612 vdd.n611 2.427
R7285 vdd.n609 vdd.n608 2.158
R7286 vdd.n610 vdd.n609 2.158
R7287 vdd.n611 vdd.n610 2.158
R7288 vdd.n613 vdd.n612 2.158
R7289 vdd.n614 vdd.n613 2.158
R7290 vdd.n615 vdd.n614 2.158
R7291 vdd.n616 vdd.n615 2.158
R7292 vdd.n617 vdd.n616 1.211
R7293 vdd.n623 vdd.n622 0.866
R7294 vdd.n635 vdd.n634 0.85
R7295 vdd.n651 vdd.n650 0.85
R7296 vdd.n663 vdd.n662 0.85
R7297 vdd.n679 vdd.n678 0.85
R7298 vdd.n691 vdd.n690 0.85
R7299 vdd.n707 vdd.n706 0.85
R7300 vdd.n719 vdd.n718 0.85
R7301 vdd.n735 vdd.n734 0.85
R7302 vdd.n747 vdd.n746 0.85
R7303 vdd.n763 vdd.n762 0.85
R7304 vdd.n775 vdd.n774 0.85
R7305 vdd.n791 vdd.n790 0.85
R7306 vdd.n803 vdd.n802 0.85
R7307 vdd.n819 vdd.n818 0.85
R7308 vdd.n831 vdd.n830 0.85
R7309 vdd.n847 vdd.n846 0.85
R7310 vdd.n859 vdd.n858 0.85
R7311 vdd.n875 vdd.n874 0.85
R7312 vdd.n887 vdd.n886 0.85
R7313 vdd.n903 vdd.n902 0.85
R7314 vdd.n915 vdd.n914 0.85
R7315 vdd.n931 vdd.n930 0.85
R7316 vdd.n943 vdd.n942 0.85
R7317 vdd.n959 vdd.n958 0.85
R7318 vdd.n971 vdd.n970 0.85
R7319 vdd.n987 vdd.n986 0.85
R7320 vdd.n999 vdd.n998 0.85
R7321 vdd.n1015 vdd.n1014 0.85
R7322 vdd.n1027 vdd.n1026 0.85
R7323 vdd.n1043 vdd.n1042 0.85
R7324 vdd.n1055 vdd.n1054 0.85
R7325 vdd.n5 vdd.n4 0.85
R7326 vdd.n599 vdd.n598 0.85
R7327 vdd.n587 vdd.n586 0.85
R7328 vdd.n571 vdd.n570 0.85
R7329 vdd.n559 vdd.n558 0.85
R7330 vdd.n27 vdd.n26 0.85
R7331 vdd.n43 vdd.n42 0.85
R7332 vdd.n55 vdd.n54 0.85
R7333 vdd.n71 vdd.n70 0.85
R7334 vdd.n83 vdd.n82 0.85
R7335 vdd.n99 vdd.n98 0.85
R7336 vdd.n111 vdd.n110 0.85
R7337 vdd.n127 vdd.n126 0.85
R7338 vdd.n139 vdd.n138 0.85
R7339 vdd.n155 vdd.n154 0.85
R7340 vdd.n167 vdd.n166 0.85
R7341 vdd.n183 vdd.n182 0.85
R7342 vdd.n195 vdd.n194 0.85
R7343 vdd.n211 vdd.n210 0.85
R7344 vdd.n223 vdd.n222 0.85
R7345 vdd.n239 vdd.n238 0.85
R7346 vdd.n251 vdd.n250 0.85
R7347 vdd.n267 vdd.n266 0.85
R7348 vdd.n279 vdd.n278 0.85
R7349 vdd.n295 vdd.n294 0.85
R7350 vdd.n307 vdd.n306 0.85
R7351 vdd.n323 vdd.n322 0.85
R7352 vdd.n335 vdd.n334 0.85
R7353 vdd.n351 vdd.n350 0.85
R7354 vdd.n363 vdd.n362 0.85
R7355 vdd.n379 vdd.n378 0.85
R7356 vdd.n391 vdd.n390 0.85
R7357 vdd.n407 vdd.n406 0.85
R7358 vdd.n419 vdd.n418 0.85
R7359 vdd.n435 vdd.n434 0.85
R7360 vdd.n447 vdd.n446 0.85
R7361 vdd.n463 vdd.n462 0.85
R7362 vdd.n475 vdd.n474 0.85
R7363 vdd.n491 vdd.n490 0.85
R7364 vdd.n503 vdd.n502 0.85
R7365 vdd.n518 vdd.n517 0.85
R7366 vdd.n545 vdd.n544 0.85
R7367 vdd.n619 vdd.n618 0.77
R7368 vdd.n620 vdd.n619 0.77
R7369 vdd.n621 vdd.n620 0.77
R7370 vdd.n622 vdd.n621 0.77
R7371 vdd.n624 vdd.n623 0.77
R7372 vdd.n625 vdd.n624 0.77
R7373 vdd.n626 vdd.n625 0.77
R7374 vdd.n627 vdd.n626 0.77
R7375 vdd.n639 vdd.n638 0.754
R7376 vdd.n638 vdd.n637 0.754
R7377 vdd.n637 vdd.n636 0.754
R7378 vdd.n636 vdd.n635 0.754
R7379 vdd.n634 vdd.n633 0.754
R7380 vdd.n633 vdd.n632 0.754
R7381 vdd.n632 vdd.n631 0.754
R7382 vdd.n631 vdd.n630 0.754
R7383 vdd.n655 vdd.n654 0.754
R7384 vdd.n654 vdd.n653 0.754
R7385 vdd.n653 vdd.n652 0.754
R7386 vdd.n652 vdd.n651 0.754
R7387 vdd.n650 vdd.n649 0.754
R7388 vdd.n649 vdd.n648 0.754
R7389 vdd.n648 vdd.n647 0.754
R7390 vdd.n647 vdd.n646 0.754
R7391 vdd.n667 vdd.n666 0.754
R7392 vdd.n666 vdd.n665 0.754
R7393 vdd.n665 vdd.n664 0.754
R7394 vdd.n664 vdd.n663 0.754
R7395 vdd.n662 vdd.n661 0.754
R7396 vdd.n661 vdd.n660 0.754
R7397 vdd.n660 vdd.n659 0.754
R7398 vdd.n659 vdd.n658 0.754
R7399 vdd.n683 vdd.n682 0.754
R7400 vdd.n682 vdd.n681 0.754
R7401 vdd.n681 vdd.n680 0.754
R7402 vdd.n680 vdd.n679 0.754
R7403 vdd.n678 vdd.n677 0.754
R7404 vdd.n677 vdd.n676 0.754
R7405 vdd.n676 vdd.n675 0.754
R7406 vdd.n675 vdd.n674 0.754
R7407 vdd.n695 vdd.n694 0.754
R7408 vdd.n694 vdd.n693 0.754
R7409 vdd.n693 vdd.n692 0.754
R7410 vdd.n692 vdd.n691 0.754
R7411 vdd.n690 vdd.n689 0.754
R7412 vdd.n689 vdd.n688 0.754
R7413 vdd.n688 vdd.n687 0.754
R7414 vdd.n687 vdd.n686 0.754
R7415 vdd.n711 vdd.n710 0.754
R7416 vdd.n710 vdd.n709 0.754
R7417 vdd.n709 vdd.n708 0.754
R7418 vdd.n708 vdd.n707 0.754
R7419 vdd.n706 vdd.n705 0.754
R7420 vdd.n705 vdd.n704 0.754
R7421 vdd.n704 vdd.n703 0.754
R7422 vdd.n703 vdd.n702 0.754
R7423 vdd.n723 vdd.n722 0.754
R7424 vdd.n722 vdd.n721 0.754
R7425 vdd.n721 vdd.n720 0.754
R7426 vdd.n720 vdd.n719 0.754
R7427 vdd.n718 vdd.n717 0.754
R7428 vdd.n717 vdd.n716 0.754
R7429 vdd.n716 vdd.n715 0.754
R7430 vdd.n715 vdd.n714 0.754
R7431 vdd.n739 vdd.n738 0.754
R7432 vdd.n738 vdd.n737 0.754
R7433 vdd.n737 vdd.n736 0.754
R7434 vdd.n736 vdd.n735 0.754
R7435 vdd.n734 vdd.n733 0.754
R7436 vdd.n733 vdd.n732 0.754
R7437 vdd.n732 vdd.n731 0.754
R7438 vdd.n731 vdd.n730 0.754
R7439 vdd.n751 vdd.n750 0.754
R7440 vdd.n750 vdd.n749 0.754
R7441 vdd.n749 vdd.n748 0.754
R7442 vdd.n748 vdd.n747 0.754
R7443 vdd.n746 vdd.n745 0.754
R7444 vdd.n745 vdd.n744 0.754
R7445 vdd.n744 vdd.n743 0.754
R7446 vdd.n743 vdd.n742 0.754
R7447 vdd.n767 vdd.n766 0.754
R7448 vdd.n766 vdd.n765 0.754
R7449 vdd.n765 vdd.n764 0.754
R7450 vdd.n764 vdd.n763 0.754
R7451 vdd.n762 vdd.n761 0.754
R7452 vdd.n761 vdd.n760 0.754
R7453 vdd.n760 vdd.n759 0.754
R7454 vdd.n759 vdd.n758 0.754
R7455 vdd.n779 vdd.n778 0.754
R7456 vdd.n778 vdd.n777 0.754
R7457 vdd.n777 vdd.n776 0.754
R7458 vdd.n776 vdd.n775 0.754
R7459 vdd.n774 vdd.n773 0.754
R7460 vdd.n773 vdd.n772 0.754
R7461 vdd.n772 vdd.n771 0.754
R7462 vdd.n771 vdd.n770 0.754
R7463 vdd.n795 vdd.n794 0.754
R7464 vdd.n794 vdd.n793 0.754
R7465 vdd.n793 vdd.n792 0.754
R7466 vdd.n792 vdd.n791 0.754
R7467 vdd.n790 vdd.n789 0.754
R7468 vdd.n789 vdd.n788 0.754
R7469 vdd.n788 vdd.n787 0.754
R7470 vdd.n787 vdd.n786 0.754
R7471 vdd.n807 vdd.n806 0.754
R7472 vdd.n806 vdd.n805 0.754
R7473 vdd.n805 vdd.n804 0.754
R7474 vdd.n804 vdd.n803 0.754
R7475 vdd.n802 vdd.n801 0.754
R7476 vdd.n801 vdd.n800 0.754
R7477 vdd.n800 vdd.n799 0.754
R7478 vdd.n799 vdd.n798 0.754
R7479 vdd.n823 vdd.n822 0.754
R7480 vdd.n822 vdd.n821 0.754
R7481 vdd.n821 vdd.n820 0.754
R7482 vdd.n820 vdd.n819 0.754
R7483 vdd.n818 vdd.n817 0.754
R7484 vdd.n817 vdd.n816 0.754
R7485 vdd.n816 vdd.n815 0.754
R7486 vdd.n815 vdd.n814 0.754
R7487 vdd.n835 vdd.n834 0.754
R7488 vdd.n834 vdd.n833 0.754
R7489 vdd.n833 vdd.n832 0.754
R7490 vdd.n832 vdd.n831 0.754
R7491 vdd.n830 vdd.n829 0.754
R7492 vdd.n829 vdd.n828 0.754
R7493 vdd.n828 vdd.n827 0.754
R7494 vdd.n827 vdd.n826 0.754
R7495 vdd.n851 vdd.n850 0.754
R7496 vdd.n850 vdd.n849 0.754
R7497 vdd.n849 vdd.n848 0.754
R7498 vdd.n848 vdd.n847 0.754
R7499 vdd.n846 vdd.n845 0.754
R7500 vdd.n845 vdd.n844 0.754
R7501 vdd.n844 vdd.n843 0.754
R7502 vdd.n843 vdd.n842 0.754
R7503 vdd.n863 vdd.n862 0.754
R7504 vdd.n862 vdd.n861 0.754
R7505 vdd.n861 vdd.n860 0.754
R7506 vdd.n860 vdd.n859 0.754
R7507 vdd.n858 vdd.n857 0.754
R7508 vdd.n857 vdd.n856 0.754
R7509 vdd.n856 vdd.n855 0.754
R7510 vdd.n855 vdd.n854 0.754
R7511 vdd.n879 vdd.n878 0.754
R7512 vdd.n878 vdd.n877 0.754
R7513 vdd.n877 vdd.n876 0.754
R7514 vdd.n876 vdd.n875 0.754
R7515 vdd.n874 vdd.n873 0.754
R7516 vdd.n873 vdd.n872 0.754
R7517 vdd.n872 vdd.n871 0.754
R7518 vdd.n871 vdd.n870 0.754
R7519 vdd.n891 vdd.n890 0.754
R7520 vdd.n890 vdd.n889 0.754
R7521 vdd.n889 vdd.n888 0.754
R7522 vdd.n888 vdd.n887 0.754
R7523 vdd.n886 vdd.n885 0.754
R7524 vdd.n885 vdd.n884 0.754
R7525 vdd.n884 vdd.n883 0.754
R7526 vdd.n883 vdd.n882 0.754
R7527 vdd.n907 vdd.n906 0.754
R7528 vdd.n906 vdd.n905 0.754
R7529 vdd.n905 vdd.n904 0.754
R7530 vdd.n904 vdd.n903 0.754
R7531 vdd.n902 vdd.n901 0.754
R7532 vdd.n901 vdd.n900 0.754
R7533 vdd.n900 vdd.n899 0.754
R7534 vdd.n899 vdd.n898 0.754
R7535 vdd.n919 vdd.n918 0.754
R7536 vdd.n918 vdd.n917 0.754
R7537 vdd.n917 vdd.n916 0.754
R7538 vdd.n916 vdd.n915 0.754
R7539 vdd.n914 vdd.n913 0.754
R7540 vdd.n913 vdd.n912 0.754
R7541 vdd.n912 vdd.n911 0.754
R7542 vdd.n911 vdd.n910 0.754
R7543 vdd.n935 vdd.n934 0.754
R7544 vdd.n934 vdd.n933 0.754
R7545 vdd.n933 vdd.n932 0.754
R7546 vdd.n932 vdd.n931 0.754
R7547 vdd.n930 vdd.n929 0.754
R7548 vdd.n929 vdd.n928 0.754
R7549 vdd.n928 vdd.n927 0.754
R7550 vdd.n927 vdd.n926 0.754
R7551 vdd.n947 vdd.n946 0.754
R7552 vdd.n946 vdd.n945 0.754
R7553 vdd.n945 vdd.n944 0.754
R7554 vdd.n944 vdd.n943 0.754
R7555 vdd.n942 vdd.n941 0.754
R7556 vdd.n941 vdd.n940 0.754
R7557 vdd.n940 vdd.n939 0.754
R7558 vdd.n939 vdd.n938 0.754
R7559 vdd.n963 vdd.n962 0.754
R7560 vdd.n962 vdd.n961 0.754
R7561 vdd.n961 vdd.n960 0.754
R7562 vdd.n960 vdd.n959 0.754
R7563 vdd.n958 vdd.n957 0.754
R7564 vdd.n957 vdd.n956 0.754
R7565 vdd.n956 vdd.n955 0.754
R7566 vdd.n955 vdd.n954 0.754
R7567 vdd.n975 vdd.n974 0.754
R7568 vdd.n974 vdd.n973 0.754
R7569 vdd.n973 vdd.n972 0.754
R7570 vdd.n972 vdd.n971 0.754
R7571 vdd.n970 vdd.n969 0.754
R7572 vdd.n969 vdd.n968 0.754
R7573 vdd.n968 vdd.n967 0.754
R7574 vdd.n967 vdd.n966 0.754
R7575 vdd.n991 vdd.n990 0.754
R7576 vdd.n990 vdd.n989 0.754
R7577 vdd.n989 vdd.n988 0.754
R7578 vdd.n988 vdd.n987 0.754
R7579 vdd.n986 vdd.n985 0.754
R7580 vdd.n985 vdd.n984 0.754
R7581 vdd.n984 vdd.n983 0.754
R7582 vdd.n983 vdd.n982 0.754
R7583 vdd.n1003 vdd.n1002 0.754
R7584 vdd.n1002 vdd.n1001 0.754
R7585 vdd.n1001 vdd.n1000 0.754
R7586 vdd.n1000 vdd.n999 0.754
R7587 vdd.n998 vdd.n997 0.754
R7588 vdd.n997 vdd.n996 0.754
R7589 vdd.n996 vdd.n995 0.754
R7590 vdd.n995 vdd.n994 0.754
R7591 vdd.n1019 vdd.n1018 0.754
R7592 vdd.n1018 vdd.n1017 0.754
R7593 vdd.n1017 vdd.n1016 0.754
R7594 vdd.n1016 vdd.n1015 0.754
R7595 vdd.n1014 vdd.n1013 0.754
R7596 vdd.n1013 vdd.n1012 0.754
R7597 vdd.n1012 vdd.n1011 0.754
R7598 vdd.n1011 vdd.n1010 0.754
R7599 vdd.n1031 vdd.n1030 0.754
R7600 vdd.n1030 vdd.n1029 0.754
R7601 vdd.n1029 vdd.n1028 0.754
R7602 vdd.n1028 vdd.n1027 0.754
R7603 vdd.n1026 vdd.n1025 0.754
R7604 vdd.n1025 vdd.n1024 0.754
R7605 vdd.n1024 vdd.n1023 0.754
R7606 vdd.n1023 vdd.n1022 0.754
R7607 vdd.n1047 vdd.n1046 0.754
R7608 vdd.n1046 vdd.n1045 0.754
R7609 vdd.n1045 vdd.n1044 0.754
R7610 vdd.n1044 vdd.n1043 0.754
R7611 vdd.n1042 vdd.n1041 0.754
R7612 vdd.n1041 vdd.n1040 0.754
R7613 vdd.n1040 vdd.n1039 0.754
R7614 vdd.n1039 vdd.n1038 0.754
R7615 vdd.n1059 vdd.n1058 0.754
R7616 vdd.n1058 vdd.n1057 0.754
R7617 vdd.n1057 vdd.n1056 0.754
R7618 vdd.n1056 vdd.n1055 0.754
R7619 vdd.n1054 vdd.n1053 0.754
R7620 vdd.n1053 vdd.n1052 0.754
R7621 vdd.n1052 vdd.n1051 0.754
R7622 vdd.n1051 vdd.n1050 0.754
R7623 vdd.n9 vdd.n8 0.754
R7624 vdd.n8 vdd.n7 0.754
R7625 vdd.n7 vdd.n6 0.754
R7626 vdd.n6 vdd.n5 0.754
R7627 vdd.n4 vdd.n3 0.754
R7628 vdd.n3 vdd.n2 0.754
R7629 vdd.n2 vdd.n1 0.754
R7630 vdd.n1 vdd.n0 0.754
R7631 vdd.n603 vdd.n602 0.754
R7632 vdd.n602 vdd.n601 0.754
R7633 vdd.n601 vdd.n600 0.754
R7634 vdd.n600 vdd.n599 0.754
R7635 vdd.n598 vdd.n597 0.754
R7636 vdd.n597 vdd.n596 0.754
R7637 vdd.n596 vdd.n595 0.754
R7638 vdd.n595 vdd.n594 0.754
R7639 vdd.n591 vdd.n590 0.754
R7640 vdd.n590 vdd.n589 0.754
R7641 vdd.n589 vdd.n588 0.754
R7642 vdd.n588 vdd.n587 0.754
R7643 vdd.n586 vdd.n585 0.754
R7644 vdd.n585 vdd.n584 0.754
R7645 vdd.n584 vdd.n583 0.754
R7646 vdd.n583 vdd.n582 0.754
R7647 vdd.n575 vdd.n574 0.754
R7648 vdd.n574 vdd.n573 0.754
R7649 vdd.n573 vdd.n572 0.754
R7650 vdd.n572 vdd.n571 0.754
R7651 vdd.n570 vdd.n569 0.754
R7652 vdd.n569 vdd.n568 0.754
R7653 vdd.n568 vdd.n567 0.754
R7654 vdd.n567 vdd.n566 0.754
R7655 vdd.n563 vdd.n562 0.754
R7656 vdd.n562 vdd.n561 0.754
R7657 vdd.n561 vdd.n560 0.754
R7658 vdd.n560 vdd.n559 0.754
R7659 vdd.n558 vdd.n557 0.754
R7660 vdd.n557 vdd.n556 0.754
R7661 vdd.n556 vdd.n555 0.754
R7662 vdd.n555 vdd.n554 0.754
R7663 vdd.n31 vdd.n30 0.754
R7664 vdd.n30 vdd.n29 0.754
R7665 vdd.n29 vdd.n28 0.754
R7666 vdd.n28 vdd.n27 0.754
R7667 vdd.n26 vdd.n25 0.754
R7668 vdd.n25 vdd.n24 0.754
R7669 vdd.n24 vdd.n23 0.754
R7670 vdd.n23 vdd.n22 0.754
R7671 vdd.n47 vdd.n46 0.754
R7672 vdd.n46 vdd.n45 0.754
R7673 vdd.n45 vdd.n44 0.754
R7674 vdd.n44 vdd.n43 0.754
R7675 vdd.n42 vdd.n41 0.754
R7676 vdd.n41 vdd.n40 0.754
R7677 vdd.n40 vdd.n39 0.754
R7678 vdd.n39 vdd.n38 0.754
R7679 vdd.n59 vdd.n58 0.754
R7680 vdd.n58 vdd.n57 0.754
R7681 vdd.n57 vdd.n56 0.754
R7682 vdd.n56 vdd.n55 0.754
R7683 vdd.n54 vdd.n53 0.754
R7684 vdd.n53 vdd.n52 0.754
R7685 vdd.n52 vdd.n51 0.754
R7686 vdd.n51 vdd.n50 0.754
R7687 vdd.n75 vdd.n74 0.754
R7688 vdd.n74 vdd.n73 0.754
R7689 vdd.n73 vdd.n72 0.754
R7690 vdd.n72 vdd.n71 0.754
R7691 vdd.n70 vdd.n69 0.754
R7692 vdd.n69 vdd.n68 0.754
R7693 vdd.n68 vdd.n67 0.754
R7694 vdd.n67 vdd.n66 0.754
R7695 vdd.n87 vdd.n86 0.754
R7696 vdd.n86 vdd.n85 0.754
R7697 vdd.n85 vdd.n84 0.754
R7698 vdd.n84 vdd.n83 0.754
R7699 vdd.n82 vdd.n81 0.754
R7700 vdd.n81 vdd.n80 0.754
R7701 vdd.n80 vdd.n79 0.754
R7702 vdd.n79 vdd.n78 0.754
R7703 vdd.n103 vdd.n102 0.754
R7704 vdd.n102 vdd.n101 0.754
R7705 vdd.n101 vdd.n100 0.754
R7706 vdd.n100 vdd.n99 0.754
R7707 vdd.n98 vdd.n97 0.754
R7708 vdd.n97 vdd.n96 0.754
R7709 vdd.n96 vdd.n95 0.754
R7710 vdd.n95 vdd.n94 0.754
R7711 vdd.n115 vdd.n114 0.754
R7712 vdd.n114 vdd.n113 0.754
R7713 vdd.n113 vdd.n112 0.754
R7714 vdd.n112 vdd.n111 0.754
R7715 vdd.n110 vdd.n109 0.754
R7716 vdd.n109 vdd.n108 0.754
R7717 vdd.n108 vdd.n107 0.754
R7718 vdd.n107 vdd.n106 0.754
R7719 vdd.n131 vdd.n130 0.754
R7720 vdd.n130 vdd.n129 0.754
R7721 vdd.n129 vdd.n128 0.754
R7722 vdd.n128 vdd.n127 0.754
R7723 vdd.n126 vdd.n125 0.754
R7724 vdd.n125 vdd.n124 0.754
R7725 vdd.n124 vdd.n123 0.754
R7726 vdd.n123 vdd.n122 0.754
R7727 vdd.n143 vdd.n142 0.754
R7728 vdd.n142 vdd.n141 0.754
R7729 vdd.n141 vdd.n140 0.754
R7730 vdd.n140 vdd.n139 0.754
R7731 vdd.n138 vdd.n137 0.754
R7732 vdd.n137 vdd.n136 0.754
R7733 vdd.n136 vdd.n135 0.754
R7734 vdd.n135 vdd.n134 0.754
R7735 vdd.n159 vdd.n158 0.754
R7736 vdd.n158 vdd.n157 0.754
R7737 vdd.n157 vdd.n156 0.754
R7738 vdd.n156 vdd.n155 0.754
R7739 vdd.n154 vdd.n153 0.754
R7740 vdd.n153 vdd.n152 0.754
R7741 vdd.n152 vdd.n151 0.754
R7742 vdd.n151 vdd.n150 0.754
R7743 vdd.n171 vdd.n170 0.754
R7744 vdd.n170 vdd.n169 0.754
R7745 vdd.n169 vdd.n168 0.754
R7746 vdd.n168 vdd.n167 0.754
R7747 vdd.n166 vdd.n165 0.754
R7748 vdd.n165 vdd.n164 0.754
R7749 vdd.n164 vdd.n163 0.754
R7750 vdd.n163 vdd.n162 0.754
R7751 vdd.n187 vdd.n186 0.754
R7752 vdd.n186 vdd.n185 0.754
R7753 vdd.n185 vdd.n184 0.754
R7754 vdd.n184 vdd.n183 0.754
R7755 vdd.n182 vdd.n181 0.754
R7756 vdd.n181 vdd.n180 0.754
R7757 vdd.n180 vdd.n179 0.754
R7758 vdd.n179 vdd.n178 0.754
R7759 vdd.n199 vdd.n198 0.754
R7760 vdd.n198 vdd.n197 0.754
R7761 vdd.n197 vdd.n196 0.754
R7762 vdd.n196 vdd.n195 0.754
R7763 vdd.n194 vdd.n193 0.754
R7764 vdd.n193 vdd.n192 0.754
R7765 vdd.n192 vdd.n191 0.754
R7766 vdd.n191 vdd.n190 0.754
R7767 vdd.n215 vdd.n214 0.754
R7768 vdd.n214 vdd.n213 0.754
R7769 vdd.n213 vdd.n212 0.754
R7770 vdd.n212 vdd.n211 0.754
R7771 vdd.n210 vdd.n209 0.754
R7772 vdd.n209 vdd.n208 0.754
R7773 vdd.n208 vdd.n207 0.754
R7774 vdd.n207 vdd.n206 0.754
R7775 vdd.n227 vdd.n226 0.754
R7776 vdd.n226 vdd.n225 0.754
R7777 vdd.n225 vdd.n224 0.754
R7778 vdd.n224 vdd.n223 0.754
R7779 vdd.n222 vdd.n221 0.754
R7780 vdd.n221 vdd.n220 0.754
R7781 vdd.n220 vdd.n219 0.754
R7782 vdd.n219 vdd.n218 0.754
R7783 vdd.n243 vdd.n242 0.754
R7784 vdd.n242 vdd.n241 0.754
R7785 vdd.n241 vdd.n240 0.754
R7786 vdd.n240 vdd.n239 0.754
R7787 vdd.n238 vdd.n237 0.754
R7788 vdd.n237 vdd.n236 0.754
R7789 vdd.n236 vdd.n235 0.754
R7790 vdd.n235 vdd.n234 0.754
R7791 vdd.n255 vdd.n254 0.754
R7792 vdd.n254 vdd.n253 0.754
R7793 vdd.n253 vdd.n252 0.754
R7794 vdd.n252 vdd.n251 0.754
R7795 vdd.n250 vdd.n249 0.754
R7796 vdd.n249 vdd.n248 0.754
R7797 vdd.n248 vdd.n247 0.754
R7798 vdd.n247 vdd.n246 0.754
R7799 vdd.n271 vdd.n270 0.754
R7800 vdd.n270 vdd.n269 0.754
R7801 vdd.n269 vdd.n268 0.754
R7802 vdd.n268 vdd.n267 0.754
R7803 vdd.n266 vdd.n265 0.754
R7804 vdd.n265 vdd.n264 0.754
R7805 vdd.n264 vdd.n263 0.754
R7806 vdd.n263 vdd.n262 0.754
R7807 vdd.n283 vdd.n282 0.754
R7808 vdd.n282 vdd.n281 0.754
R7809 vdd.n281 vdd.n280 0.754
R7810 vdd.n280 vdd.n279 0.754
R7811 vdd.n278 vdd.n277 0.754
R7812 vdd.n277 vdd.n276 0.754
R7813 vdd.n276 vdd.n275 0.754
R7814 vdd.n275 vdd.n274 0.754
R7815 vdd.n299 vdd.n298 0.754
R7816 vdd.n298 vdd.n297 0.754
R7817 vdd.n297 vdd.n296 0.754
R7818 vdd.n296 vdd.n295 0.754
R7819 vdd.n294 vdd.n293 0.754
R7820 vdd.n293 vdd.n292 0.754
R7821 vdd.n292 vdd.n291 0.754
R7822 vdd.n291 vdd.n290 0.754
R7823 vdd.n311 vdd.n310 0.754
R7824 vdd.n310 vdd.n309 0.754
R7825 vdd.n309 vdd.n308 0.754
R7826 vdd.n308 vdd.n307 0.754
R7827 vdd.n306 vdd.n305 0.754
R7828 vdd.n305 vdd.n304 0.754
R7829 vdd.n304 vdd.n303 0.754
R7830 vdd.n303 vdd.n302 0.754
R7831 vdd.n327 vdd.n326 0.754
R7832 vdd.n326 vdd.n325 0.754
R7833 vdd.n325 vdd.n324 0.754
R7834 vdd.n324 vdd.n323 0.754
R7835 vdd.n322 vdd.n321 0.754
R7836 vdd.n321 vdd.n320 0.754
R7837 vdd.n320 vdd.n319 0.754
R7838 vdd.n319 vdd.n318 0.754
R7839 vdd.n339 vdd.n338 0.754
R7840 vdd.n338 vdd.n337 0.754
R7841 vdd.n337 vdd.n336 0.754
R7842 vdd.n336 vdd.n335 0.754
R7843 vdd.n334 vdd.n333 0.754
R7844 vdd.n333 vdd.n332 0.754
R7845 vdd.n332 vdd.n331 0.754
R7846 vdd.n331 vdd.n330 0.754
R7847 vdd.n355 vdd.n354 0.754
R7848 vdd.n354 vdd.n353 0.754
R7849 vdd.n353 vdd.n352 0.754
R7850 vdd.n352 vdd.n351 0.754
R7851 vdd.n350 vdd.n349 0.754
R7852 vdd.n349 vdd.n348 0.754
R7853 vdd.n348 vdd.n347 0.754
R7854 vdd.n347 vdd.n346 0.754
R7855 vdd.n367 vdd.n366 0.754
R7856 vdd.n366 vdd.n365 0.754
R7857 vdd.n365 vdd.n364 0.754
R7858 vdd.n364 vdd.n363 0.754
R7859 vdd.n362 vdd.n361 0.754
R7860 vdd.n361 vdd.n360 0.754
R7861 vdd.n360 vdd.n359 0.754
R7862 vdd.n359 vdd.n358 0.754
R7863 vdd.n383 vdd.n382 0.754
R7864 vdd.n382 vdd.n381 0.754
R7865 vdd.n381 vdd.n380 0.754
R7866 vdd.n380 vdd.n379 0.754
R7867 vdd.n378 vdd.n377 0.754
R7868 vdd.n377 vdd.n376 0.754
R7869 vdd.n376 vdd.n375 0.754
R7870 vdd.n375 vdd.n374 0.754
R7871 vdd.n395 vdd.n394 0.754
R7872 vdd.n394 vdd.n393 0.754
R7873 vdd.n393 vdd.n392 0.754
R7874 vdd.n392 vdd.n391 0.754
R7875 vdd.n390 vdd.n389 0.754
R7876 vdd.n389 vdd.n388 0.754
R7877 vdd.n388 vdd.n387 0.754
R7878 vdd.n387 vdd.n386 0.754
R7879 vdd.n411 vdd.n410 0.754
R7880 vdd.n410 vdd.n409 0.754
R7881 vdd.n409 vdd.n408 0.754
R7882 vdd.n408 vdd.n407 0.754
R7883 vdd.n406 vdd.n405 0.754
R7884 vdd.n405 vdd.n404 0.754
R7885 vdd.n404 vdd.n403 0.754
R7886 vdd.n403 vdd.n402 0.754
R7887 vdd.n423 vdd.n422 0.754
R7888 vdd.n422 vdd.n421 0.754
R7889 vdd.n421 vdd.n420 0.754
R7890 vdd.n420 vdd.n419 0.754
R7891 vdd.n418 vdd.n417 0.754
R7892 vdd.n417 vdd.n416 0.754
R7893 vdd.n416 vdd.n415 0.754
R7894 vdd.n415 vdd.n414 0.754
R7895 vdd.n439 vdd.n438 0.754
R7896 vdd.n438 vdd.n437 0.754
R7897 vdd.n437 vdd.n436 0.754
R7898 vdd.n436 vdd.n435 0.754
R7899 vdd.n434 vdd.n433 0.754
R7900 vdd.n433 vdd.n432 0.754
R7901 vdd.n432 vdd.n431 0.754
R7902 vdd.n431 vdd.n430 0.754
R7903 vdd.n451 vdd.n450 0.754
R7904 vdd.n450 vdd.n449 0.754
R7905 vdd.n449 vdd.n448 0.754
R7906 vdd.n448 vdd.n447 0.754
R7907 vdd.n446 vdd.n445 0.754
R7908 vdd.n445 vdd.n444 0.754
R7909 vdd.n444 vdd.n443 0.754
R7910 vdd.n443 vdd.n442 0.754
R7911 vdd.n467 vdd.n466 0.754
R7912 vdd.n466 vdd.n465 0.754
R7913 vdd.n465 vdd.n464 0.754
R7914 vdd.n464 vdd.n463 0.754
R7915 vdd.n462 vdd.n461 0.754
R7916 vdd.n461 vdd.n460 0.754
R7917 vdd.n460 vdd.n459 0.754
R7918 vdd.n459 vdd.n458 0.754
R7919 vdd.n479 vdd.n478 0.754
R7920 vdd.n478 vdd.n477 0.754
R7921 vdd.n477 vdd.n476 0.754
R7922 vdd.n476 vdd.n475 0.754
R7923 vdd.n474 vdd.n473 0.754
R7924 vdd.n473 vdd.n472 0.754
R7925 vdd.n472 vdd.n471 0.754
R7926 vdd.n471 vdd.n470 0.754
R7927 vdd.n495 vdd.n494 0.754
R7928 vdd.n494 vdd.n493 0.754
R7929 vdd.n493 vdd.n492 0.754
R7930 vdd.n492 vdd.n491 0.754
R7931 vdd.n490 vdd.n489 0.754
R7932 vdd.n489 vdd.n488 0.754
R7933 vdd.n488 vdd.n487 0.754
R7934 vdd.n487 vdd.n486 0.754
R7935 vdd.n507 vdd.n506 0.754
R7936 vdd.n506 vdd.n505 0.754
R7937 vdd.n505 vdd.n504 0.754
R7938 vdd.n504 vdd.n503 0.754
R7939 vdd.n502 vdd.n501 0.754
R7940 vdd.n501 vdd.n500 0.754
R7941 vdd.n500 vdd.n499 0.754
R7942 vdd.n499 vdd.n498 0.754
R7943 vdd.n522 vdd.n521 0.754
R7944 vdd.n521 vdd.n520 0.754
R7945 vdd.n520 vdd.n519 0.754
R7946 vdd.n519 vdd.n518 0.754
R7947 vdd.n517 vdd.n516 0.754
R7948 vdd.n516 vdd.n515 0.754
R7949 vdd.n515 vdd.n514 0.754
R7950 vdd.n514 vdd.n513 0.754
R7951 vdd.n549 vdd.n548 0.754
R7952 vdd.n548 vdd.n547 0.754
R7953 vdd.n547 vdd.n546 0.754
R7954 vdd.n546 vdd.n545 0.754
R7955 vdd.n544 vdd.n543 0.754
R7956 vdd.n543 vdd.n542 0.754
R7957 vdd.n542 vdd.n541 0.754
R7958 vdd.n541 vdd.n540 0.754
R7959 vdd.n16 vdd.n15 0.726
R7960 vdd.n13 vdd.n12 0.58
R7961 vdd.n14 vdd.n13 0.58
R7962 vdd.n15 vdd.n14 0.58
R7963 vdd.n17 vdd.n16 0.58
R7964 vdd.n18 vdd.n17 0.58
R7965 vdd.n19 vdd.n18 0.58
R7966 vdd.n20 vdd.n19 0.58
R7967 vdd.n21 vdd.n20 0.495
R7968 vdd.n550 vdd.n549 0.427
R7969 vdd.n628 vdd.n627 0.426
R7970 vdd.n640 vdd.n639 0.426
R7971 vdd.n656 vdd.n655 0.426
R7972 vdd.n668 vdd.n667 0.426
R7973 vdd.n684 vdd.n683 0.426
R7974 vdd.n696 vdd.n695 0.426
R7975 vdd.n712 vdd.n711 0.426
R7976 vdd.n724 vdd.n723 0.426
R7977 vdd.n740 vdd.n739 0.426
R7978 vdd.n752 vdd.n751 0.426
R7979 vdd.n768 vdd.n767 0.426
R7980 vdd.n780 vdd.n779 0.426
R7981 vdd.n796 vdd.n795 0.426
R7982 vdd.n808 vdd.n807 0.426
R7983 vdd.n824 vdd.n823 0.426
R7984 vdd.n836 vdd.n835 0.426
R7985 vdd.n852 vdd.n851 0.426
R7986 vdd.n864 vdd.n863 0.426
R7987 vdd.n880 vdd.n879 0.426
R7988 vdd.n892 vdd.n891 0.426
R7989 vdd.n908 vdd.n907 0.426
R7990 vdd.n920 vdd.n919 0.426
R7991 vdd.n936 vdd.n935 0.426
R7992 vdd.n948 vdd.n947 0.426
R7993 vdd.n964 vdd.n963 0.426
R7994 vdd.n976 vdd.n975 0.426
R7995 vdd.n992 vdd.n991 0.426
R7996 vdd.n1004 vdd.n1003 0.426
R7997 vdd.n1020 vdd.n1019 0.426
R7998 vdd.n1032 vdd.n1031 0.426
R7999 vdd.n1048 vdd.n1047 0.426
R8000 vdd.n1060 vdd.n1059 0.426
R8001 vdd.n10 vdd.n9 0.426
R8002 vdd.n604 vdd.n603 0.426
R8003 vdd.n592 vdd.n591 0.426
R8004 vdd.n576 vdd.n575 0.426
R8005 vdd.n564 vdd.n563 0.426
R8006 vdd.n32 vdd.n31 0.426
R8007 vdd.n48 vdd.n47 0.426
R8008 vdd.n60 vdd.n59 0.426
R8009 vdd.n76 vdd.n75 0.426
R8010 vdd.n88 vdd.n87 0.426
R8011 vdd.n104 vdd.n103 0.426
R8012 vdd.n116 vdd.n115 0.426
R8013 vdd.n132 vdd.n131 0.426
R8014 vdd.n144 vdd.n143 0.426
R8015 vdd.n160 vdd.n159 0.426
R8016 vdd.n172 vdd.n171 0.426
R8017 vdd.n188 vdd.n187 0.426
R8018 vdd.n200 vdd.n199 0.426
R8019 vdd.n216 vdd.n215 0.426
R8020 vdd.n228 vdd.n227 0.426
R8021 vdd.n244 vdd.n243 0.426
R8022 vdd.n256 vdd.n255 0.426
R8023 vdd.n272 vdd.n271 0.426
R8024 vdd.n284 vdd.n283 0.426
R8025 vdd.n300 vdd.n299 0.426
R8026 vdd.n312 vdd.n311 0.426
R8027 vdd.n328 vdd.n327 0.426
R8028 vdd.n340 vdd.n339 0.426
R8029 vdd.n356 vdd.n355 0.426
R8030 vdd.n368 vdd.n367 0.426
R8031 vdd.n384 vdd.n383 0.426
R8032 vdd.n396 vdd.n395 0.426
R8033 vdd.n412 vdd.n411 0.426
R8034 vdd.n424 vdd.n423 0.426
R8035 vdd.n440 vdd.n439 0.426
R8036 vdd.n452 vdd.n451 0.426
R8037 vdd.n468 vdd.n467 0.426
R8038 vdd.n480 vdd.n479 0.426
R8039 vdd.n496 vdd.n495 0.426
R8040 vdd.n508 vdd.n507 0.426
R8041 vdd.n523 vdd.n522 0.426
R8042 vdd.n642 vdd.n641 0.094
R8043 vdd.n645 vdd.n644 0.094
R8044 vdd.n670 vdd.n669 0.094
R8045 vdd.n673 vdd.n672 0.094
R8046 vdd.n698 vdd.n697 0.094
R8047 vdd.n701 vdd.n700 0.094
R8048 vdd.n726 vdd.n725 0.094
R8049 vdd.n729 vdd.n728 0.094
R8050 vdd.n754 vdd.n753 0.094
R8051 vdd.n757 vdd.n756 0.094
R8052 vdd.n782 vdd.n781 0.094
R8053 vdd.n785 vdd.n784 0.094
R8054 vdd.n810 vdd.n809 0.094
R8055 vdd.n813 vdd.n812 0.094
R8056 vdd.n838 vdd.n837 0.094
R8057 vdd.n841 vdd.n840 0.094
R8058 vdd.n866 vdd.n865 0.094
R8059 vdd.n869 vdd.n868 0.094
R8060 vdd.n894 vdd.n893 0.094
R8061 vdd.n897 vdd.n896 0.094
R8062 vdd.n922 vdd.n921 0.094
R8063 vdd.n925 vdd.n924 0.094
R8064 vdd.n950 vdd.n949 0.094
R8065 vdd.n953 vdd.n952 0.094
R8066 vdd.n978 vdd.n977 0.094
R8067 vdd.n981 vdd.n980 0.094
R8068 vdd.n1006 vdd.n1005 0.094
R8069 vdd.n1009 vdd.n1008 0.094
R8070 vdd.n1034 vdd.n1033 0.094
R8071 vdd.n1037 vdd.n1036 0.094
R8072 vdd.n1062 vdd.n1061 0.094
R8073 vdd.n1065 vdd.n1064 0.094
R8074 vdd.n606 vdd.n605 0.094
R8075 vdd.n581 vdd.n580 0.094
R8076 vdd.n578 vdd.n577 0.094
R8077 vdd.n553 vdd.n552 0.094
R8078 vdd.n34 vdd.n33 0.094
R8079 vdd.n37 vdd.n36 0.094
R8080 vdd.n62 vdd.n61 0.094
R8081 vdd.n65 vdd.n64 0.094
R8082 vdd.n90 vdd.n89 0.094
R8083 vdd.n93 vdd.n92 0.094
R8084 vdd.n118 vdd.n117 0.094
R8085 vdd.n121 vdd.n120 0.094
R8086 vdd.n146 vdd.n145 0.094
R8087 vdd.n149 vdd.n148 0.094
R8088 vdd.n174 vdd.n173 0.094
R8089 vdd.n177 vdd.n176 0.094
R8090 vdd.n202 vdd.n201 0.094
R8091 vdd.n205 vdd.n204 0.094
R8092 vdd.n230 vdd.n229 0.094
R8093 vdd.n233 vdd.n232 0.094
R8094 vdd.n258 vdd.n257 0.094
R8095 vdd.n261 vdd.n260 0.094
R8096 vdd.n286 vdd.n285 0.094
R8097 vdd.n289 vdd.n288 0.094
R8098 vdd.n314 vdd.n313 0.094
R8099 vdd.n317 vdd.n316 0.094
R8100 vdd.n342 vdd.n341 0.094
R8101 vdd.n345 vdd.n344 0.094
R8102 vdd.n370 vdd.n369 0.094
R8103 vdd.n373 vdd.n372 0.094
R8104 vdd.n398 vdd.n397 0.094
R8105 vdd.n401 vdd.n400 0.094
R8106 vdd.n426 vdd.n425 0.094
R8107 vdd.n429 vdd.n428 0.094
R8108 vdd.n454 vdd.n453 0.094
R8109 vdd.n457 vdd.n456 0.094
R8110 vdd.n482 vdd.n481 0.094
R8111 vdd.n485 vdd.n484 0.094
R8112 vdd.n510 vdd.n509 0.094
R8113 vdd.n551 vdd.n539 0.093
R8114 vdd.n21 vdd.n11 0.082
R8115 vdd.n35 vdd.n21 0.021
R8116 vdd.n49 vdd.n35 0.002
R8117 vdd.n63 vdd.n49 0.002
R8118 vdd.n77 vdd.n63 0.002
R8119 vdd.n91 vdd.n77 0.002
R8120 vdd.n105 vdd.n91 0.002
R8121 vdd.n119 vdd.n105 0.002
R8122 vdd.n133 vdd.n119 0.002
R8123 vdd.n147 vdd.n133 0.002
R8124 vdd.n161 vdd.n147 0.002
R8125 vdd.n175 vdd.n161 0.002
R8126 vdd.n189 vdd.n175 0.002
R8127 vdd.n203 vdd.n189 0.002
R8128 vdd.n217 vdd.n203 0.002
R8129 vdd.n231 vdd.n217 0.002
R8130 vdd.n245 vdd.n231 0.002
R8131 vdd.n259 vdd.n245 0.002
R8132 vdd.n273 vdd.n259 0.002
R8133 vdd.n287 vdd.n273 0.002
R8134 vdd.n301 vdd.n287 0.002
R8135 vdd.n315 vdd.n301 0.002
R8136 vdd.n329 vdd.n315 0.002
R8137 vdd.n343 vdd.n329 0.002
R8138 vdd.n357 vdd.n343 0.002
R8139 vdd.n371 vdd.n357 0.002
R8140 vdd.n385 vdd.n371 0.002
R8141 vdd.n399 vdd.n385 0.002
R8142 vdd.n413 vdd.n399 0.002
R8143 vdd.n427 vdd.n413 0.002
R8144 vdd.n441 vdd.n427 0.002
R8145 vdd.n455 vdd.n441 0.002
R8146 vdd.n469 vdd.n455 0.002
R8147 vdd.n483 vdd.n469 0.002
R8148 vdd.n497 vdd.n483 0.002
R8149 vdd.n511 vdd.n497 0.002
R8150 vdd.n524 vdd.n511 0.002
R8151 vdd.n551 vdd.n524 0.002
R8152 vdd.n565 vdd.n551 0.002
R8153 vdd.n579 vdd.n565 0.002
R8154 vdd.n593 vdd.n579 0.002
R8155 vdd.n607 vdd.n593 0.002
R8156 vdd vdd.n607 0.002
R8157 vdd vdd.n1063 0.002
R8158 vdd.n1063 vdd.n1049 0.002
R8159 vdd.n1049 vdd.n1035 0.002
R8160 vdd.n1035 vdd.n1021 0.002
R8161 vdd.n1021 vdd.n1007 0.002
R8162 vdd.n1007 vdd.n993 0.002
R8163 vdd.n993 vdd.n979 0.002
R8164 vdd.n979 vdd.n965 0.002
R8165 vdd.n965 vdd.n951 0.002
R8166 vdd.n951 vdd.n937 0.002
R8167 vdd.n937 vdd.n923 0.002
R8168 vdd.n923 vdd.n909 0.002
R8169 vdd.n909 vdd.n895 0.002
R8170 vdd.n895 vdd.n881 0.002
R8171 vdd.n881 vdd.n867 0.002
R8172 vdd.n867 vdd.n853 0.002
R8173 vdd.n853 vdd.n839 0.002
R8174 vdd.n839 vdd.n825 0.002
R8175 vdd.n825 vdd.n811 0.002
R8176 vdd.n811 vdd.n797 0.002
R8177 vdd.n797 vdd.n783 0.002
R8178 vdd.n783 vdd.n769 0.002
R8179 vdd.n769 vdd.n755 0.002
R8180 vdd.n755 vdd.n741 0.002
R8181 vdd.n741 vdd.n727 0.002
R8182 vdd.n727 vdd.n713 0.002
R8183 vdd.n713 vdd.n699 0.002
R8184 vdd.n699 vdd.n685 0.002
R8185 vdd.n685 vdd.n671 0.002
R8186 vdd.n671 vdd.n657 0.002
R8187 vdd.n657 vdd.n643 0.002
R8188 vdd.n643 vdd.n629 0.002
R8189 vdd.n551 vdd.n550 0.001
R8190 vdd.n629 vdd.n628 0.001
R8191 vdd.n643 vdd.n640 0.001
R8192 vdd.n657 vdd.n656 0.001
R8193 vdd.n671 vdd.n668 0.001
R8194 vdd.n685 vdd.n684 0.001
R8195 vdd.n699 vdd.n696 0.001
R8196 vdd.n713 vdd.n712 0.001
R8197 vdd.n727 vdd.n724 0.001
R8198 vdd.n741 vdd.n740 0.001
R8199 vdd.n755 vdd.n752 0.001
R8200 vdd.n769 vdd.n768 0.001
R8201 vdd.n783 vdd.n780 0.001
R8202 vdd.n797 vdd.n796 0.001
R8203 vdd.n811 vdd.n808 0.001
R8204 vdd.n825 vdd.n824 0.001
R8205 vdd.n839 vdd.n836 0.001
R8206 vdd.n853 vdd.n852 0.001
R8207 vdd.n867 vdd.n864 0.001
R8208 vdd.n881 vdd.n880 0.001
R8209 vdd.n895 vdd.n892 0.001
R8210 vdd.n909 vdd.n908 0.001
R8211 vdd.n923 vdd.n920 0.001
R8212 vdd.n937 vdd.n936 0.001
R8213 vdd.n951 vdd.n948 0.001
R8214 vdd.n965 vdd.n964 0.001
R8215 vdd.n979 vdd.n976 0.001
R8216 vdd.n993 vdd.n992 0.001
R8217 vdd.n1007 vdd.n1004 0.001
R8218 vdd.n1021 vdd.n1020 0.001
R8219 vdd.n1035 vdd.n1032 0.001
R8220 vdd.n1049 vdd.n1048 0.001
R8221 vdd.n1063 vdd.n1060 0.001
R8222 vdd vdd.n10 0.001
R8223 vdd.n607 vdd.n604 0.001
R8224 vdd.n593 vdd.n592 0.001
R8225 vdd.n579 vdd.n576 0.001
R8226 vdd.n565 vdd.n564 0.001
R8227 vdd.n35 vdd.n32 0.001
R8228 vdd.n49 vdd.n48 0.001
R8229 vdd.n63 vdd.n60 0.001
R8230 vdd.n77 vdd.n76 0.001
R8231 vdd.n91 vdd.n88 0.001
R8232 vdd.n105 vdd.n104 0.001
R8233 vdd.n119 vdd.n116 0.001
R8234 vdd.n133 vdd.n132 0.001
R8235 vdd.n147 vdd.n144 0.001
R8236 vdd.n161 vdd.n160 0.001
R8237 vdd.n175 vdd.n172 0.001
R8238 vdd.n189 vdd.n188 0.001
R8239 vdd.n203 vdd.n200 0.001
R8240 vdd.n217 vdd.n216 0.001
R8241 vdd.n231 vdd.n228 0.001
R8242 vdd.n245 vdd.n244 0.001
R8243 vdd.n259 vdd.n256 0.001
R8244 vdd.n273 vdd.n272 0.001
R8245 vdd.n287 vdd.n284 0.001
R8246 vdd.n301 vdd.n300 0.001
R8247 vdd.n315 vdd.n312 0.001
R8248 vdd.n329 vdd.n328 0.001
R8249 vdd.n343 vdd.n340 0.001
R8250 vdd.n357 vdd.n356 0.001
R8251 vdd.n371 vdd.n368 0.001
R8252 vdd.n385 vdd.n384 0.001
R8253 vdd.n399 vdd.n396 0.001
R8254 vdd.n413 vdd.n412 0.001
R8255 vdd.n427 vdd.n424 0.001
R8256 vdd.n441 vdd.n440 0.001
R8257 vdd.n455 vdd.n452 0.001
R8258 vdd.n469 vdd.n468 0.001
R8259 vdd.n483 vdd.n480 0.001
R8260 vdd.n497 vdd.n496 0.001
R8261 vdd.n511 vdd.n508 0.001
R8262 vdd.n524 vdd.n523 0.001
R8263 vdd.n539 vdd.n538 0.001
R8264 vdd.n539 vdd.n537 0.001
R8265 vdd.n629 vdd.n617 0.001
R8266 vdd.n643 vdd.n642 0.001
R8267 vdd.n657 vdd.n645 0.001
R8268 vdd.n671 vdd.n670 0.001
R8269 vdd.n685 vdd.n673 0.001
R8270 vdd.n699 vdd.n698 0.001
R8271 vdd.n713 vdd.n701 0.001
R8272 vdd.n727 vdd.n726 0.001
R8273 vdd.n741 vdd.n729 0.001
R8274 vdd.n755 vdd.n754 0.001
R8275 vdd.n769 vdd.n757 0.001
R8276 vdd.n783 vdd.n782 0.001
R8277 vdd.n797 vdd.n785 0.001
R8278 vdd.n811 vdd.n810 0.001
R8279 vdd.n825 vdd.n813 0.001
R8280 vdd.n839 vdd.n838 0.001
R8281 vdd.n853 vdd.n841 0.001
R8282 vdd.n867 vdd.n866 0.001
R8283 vdd.n881 vdd.n869 0.001
R8284 vdd.n895 vdd.n894 0.001
R8285 vdd.n909 vdd.n897 0.001
R8286 vdd.n923 vdd.n922 0.001
R8287 vdd.n937 vdd.n925 0.001
R8288 vdd.n951 vdd.n950 0.001
R8289 vdd.n965 vdd.n953 0.001
R8290 vdd.n979 vdd.n978 0.001
R8291 vdd.n993 vdd.n981 0.001
R8292 vdd.n1007 vdd.n1006 0.001
R8293 vdd.n1021 vdd.n1009 0.001
R8294 vdd.n1035 vdd.n1034 0.001
R8295 vdd.n1049 vdd.n1037 0.001
R8296 vdd.n1063 vdd.n1062 0.001
R8297 vdd.n1065 vdd 0.001
R8298 vdd.n607 vdd.n606 0.001
R8299 vdd.n593 vdd.n581 0.001
R8300 vdd.n579 vdd.n578 0.001
R8301 vdd.n565 vdd.n553 0.001
R8302 vdd.n524 vdd.n512 0.001
R8303 vdd.n511 vdd.n510 0.001
R8304 vdd.n497 vdd.n485 0.001
R8305 vdd.n483 vdd.n482 0.001
R8306 vdd.n469 vdd.n457 0.001
R8307 vdd.n455 vdd.n454 0.001
R8308 vdd.n441 vdd.n429 0.001
R8309 vdd.n427 vdd.n426 0.001
R8310 vdd.n413 vdd.n401 0.001
R8311 vdd.n399 vdd.n398 0.001
R8312 vdd.n385 vdd.n373 0.001
R8313 vdd.n371 vdd.n370 0.001
R8314 vdd.n357 vdd.n345 0.001
R8315 vdd.n343 vdd.n342 0.001
R8316 vdd.n329 vdd.n317 0.001
R8317 vdd.n315 vdd.n314 0.001
R8318 vdd.n301 vdd.n289 0.001
R8319 vdd.n287 vdd.n286 0.001
R8320 vdd.n273 vdd.n261 0.001
R8321 vdd.n259 vdd.n258 0.001
R8322 vdd.n245 vdd.n233 0.001
R8323 vdd.n231 vdd.n230 0.001
R8324 vdd.n217 vdd.n205 0.001
R8325 vdd.n203 vdd.n202 0.001
R8326 vdd.n189 vdd.n177 0.001
R8327 vdd.n175 vdd.n174 0.001
R8328 vdd.n161 vdd.n149 0.001
R8329 vdd.n147 vdd.n146 0.001
R8330 vdd.n133 vdd.n121 0.001
R8331 vdd.n119 vdd.n118 0.001
R8332 vdd.n105 vdd.n93 0.001
R8333 vdd.n91 vdd.n90 0.001
R8334 vdd.n77 vdd.n65 0.001
R8335 vdd.n63 vdd.n62 0.001
R8336 vdd.n49 vdd.n37 0.001
R8337 vdd.n35 vdd.n34 0.001
R8338 vp_n.n221 vp_n.t104 721.861
R8339 vp_n.n219 vp_n.t191 721.861
R8340 vp_n.n217 vp_n.t142 721.861
R8341 vp_n.n215 vp_n.t226 721.861
R8342 vp_n.n213 vp_n.t0 721.861
R8343 vp_n.n211 vp_n.t286 721.861
R8344 vp_n.n209 vp_n.t69 721.861
R8345 vp_n.n207 vp_n.t28 721.861
R8346 vp_n.n205 vp_n.t112 721.861
R8347 vp_n.n203 vp_n.t250 721.861
R8348 vp_n.n201 vp_n.t299 721.861
R8349 vp_n.n199 vp_n.t225 721.861
R8350 vp_n.n197 vp_n.t202 721.861
R8351 vp_n.n195 vp_n.t118 721.861
R8352 vp_n.n193 vp_n.t167 721.861
R8353 vp_n.n191 vp_n.t46 721.861
R8354 vp_n.n189 vp_n.t270 721.861
R8355 vp_n.n187 vp_n.t10 721.861
R8356 vp_n.n185 vp_n.t236 721.861
R8357 vp_n.n183 vp_n.t277 721.861
R8358 vp_n.n181 vp_n.t168 721.861
R8359 vp_n.n179 vp_n.t212 721.861
R8360 vp_n.n177 vp_n.t127 721.861
R8361 vp_n.n175 vp_n.t45 721.861
R8362 vp_n.n173 vp_n.t91 721.861
R8363 vp_n.n171 vp_n.t278 721.861
R8364 vp_n.n169 vp_n.t22 721.861
R8365 vp_n.n167 vp_n.t244 721.861
R8366 vp_n.n165 vp_n.t166 721.861
R8367 vp_n.n163 vp_n.t211 721.861
R8368 vp_n.n161 vp_n.t92 721.861
R8369 vp_n.n159 vp_n.t143 721.861
R8370 vp_n.n157 vp_n.t53 721.861
R8371 vp_n.n155 vp_n.t60 721.861
R8372 vp_n.n153 vp_n.t281 721.861
R8373 vp_n.n151 vp_n.t170 721.861
R8374 vp_n.n149 vp_n.t218 721.861
R8375 vp_n.n147 vp_n.t133 721.861
R8376 vp_n.n145 vp_n.t182 721.861
R8377 vp_n.n143 vp_n.t95 721.861
R8378 vp_n.n141 vp_n.t111 721.861
R8379 vp_n.n139 vp_n.t27 721.861
R8380 vp_n.n137 vp_n.t247 721.861
R8381 vp_n.n135 vp_n.t292 721.861
R8382 vp_n.n133 vp_n.t217 721.861
R8383 vp_n.n131 vp_n.t231 721.861
R8384 vp_n.n129 vp_n.t149 721.861
R8385 vp_n.n127 vp_n.t59 721.861
R8386 vp_n.n125 vp_n.t109 721.861
R8387 vp_n.n123 vp_n.t26 721.861
R8388 vp_n.n121 vp_n.t40 721.861
R8389 vp_n.n119 vp_n.t261 721.861
R8390 vp_n.n117 vp_n.t4 721.861
R8391 vp_n.n115 vp_n.t229 721.861
R8392 vp_n.n113 vp_n.t148 721.861
R8393 vp_n.n111 vp_n.t161 721.861
R8394 vp_n.n109 vp_n.t73 721.861
R8395 vp_n.n107 vp_n.t298 721.861
R8396 vp_n.n105 vp_n.t224 721.861
R8397 vp_n.n103 vp_n.t139 721.861
R8398 vp_n.n101 vp_n.t156 721.861
R8399 vp_n.n99 vp_n.t66 721.861
R8400 vp_n.n97 vp_n.t117 721.861
R8401 vp_n.n95 vp_n.t34 721.861
R8402 vp_n.n93 vp_n.t79 721.861
R8403 vp_n.n91 vp_n.t269 721.861
R8404 vp_n.n89 vp_n.t189 721.861
R8405 vp_n.n87 vp_n.t235 721.861
R8406 vp_n.n85 vp_n.t154 721.861
R8407 vp_n.n83 vp_n.t200 721.861
R8408 vp_n.n81 vp_n.t80 721.861
R8409 vp_n.n79 vp_n.t126 721.861
R8410 vp_n.n77 vp_n.t44 721.861
R8411 vp_n.n75 vp_n.t267 721.861
R8412 vp_n.n74 vp_n.t9 721.861
R8413 vp_n.n221 vp_n.t94 721.861
R8414 vp_n.n219 vp_n.t180 721.861
R8415 vp_n.n217 vp_n.t131 721.861
R8416 vp_n.n215 vp_n.t216 721.861
R8417 vp_n.n213 vp_n.t291 721.861
R8418 vp_n.n211 vp_n.t280 721.861
R8419 vp_n.n209 vp_n.t58 721.861
R8420 vp_n.n207 vp_n.t18 721.861
R8421 vp_n.n205 vp_n.t101 721.861
R8422 vp_n.n203 vp_n.t243 721.861
R8423 vp_n.n201 vp_n.t289 721.861
R8424 vp_n.n199 vp_n.t215 721.861
R8425 vp_n.n197 vp_n.t194 721.861
R8426 vp_n.n195 vp_n.t107 721.861
R8427 vp_n.n193 vp_n.t159 721.861
R8428 vp_n.n191 vp_n.t38 721.861
R8429 vp_n.n189 vp_n.t260 721.861
R8430 vp_n.n187 vp_n.t2 721.861
R8431 vp_n.n185 vp_n.t228 721.861
R8432 vp_n.n183 vp_n.t271 721.861
R8433 vp_n.n181 vp_n.t160 721.861
R8434 vp_n.n179 vp_n.t205 721.861
R8435 vp_n.n177 vp_n.t120 721.861
R8436 vp_n.n175 vp_n.t37 721.861
R8437 vp_n.n173 vp_n.t83 721.861
R8438 vp_n.n171 vp_n.t272 721.861
R8439 vp_n.n169 vp_n.t13 721.861
R8440 vp_n.n167 vp_n.t237 721.861
R8441 vp_n.n165 vp_n.t158 721.861
R8442 vp_n.n163 vp_n.t204 721.861
R8443 vp_n.n161 vp_n.t84 721.861
R8444 vp_n.n159 vp_n.t132 721.861
R8445 vp_n.n157 vp_n.t47 721.861
R8446 vp_n.n155 vp_n.t51 721.861
R8447 vp_n.n153 vp_n.t275 721.861
R8448 vp_n.n151 vp_n.t164 721.861
R8449 vp_n.n149 vp_n.t209 721.861
R8450 vp_n.n147 vp_n.t123 721.861
R8451 vp_n.n145 vp_n.t173 721.861
R8452 vp_n.n143 vp_n.t88 721.861
R8453 vp_n.n141 vp_n.t100 721.861
R8454 vp_n.n139 vp_n.t17 721.861
R8455 vp_n.n137 vp_n.t240 721.861
R8456 vp_n.n135 vp_n.t284 721.861
R8457 vp_n.n133 vp_n.t208 721.861
R8458 vp_n.n131 vp_n.t221 721.861
R8459 vp_n.n129 vp_n.t137 721.861
R8460 vp_n.n127 vp_n.t50 721.861
R8461 vp_n.n125 vp_n.t98 721.861
R8462 vp_n.n123 vp_n.t16 721.861
R8463 vp_n.n121 vp_n.t31 721.861
R8464 vp_n.n119 vp_n.t251 721.861
R8465 vp_n.n117 vp_n.t294 721.861
R8466 vp_n.n115 vp_n.t219 721.861
R8467 vp_n.n113 vp_n.t136 721.861
R8468 vp_n.n111 vp_n.t151 721.861
R8469 vp_n.n109 vp_n.t62 721.861
R8470 vp_n.n107 vp_n.t288 721.861
R8471 vp_n.n105 vp_n.t214 721.861
R8472 vp_n.n103 vp_n.t128 721.861
R8473 vp_n.n101 vp_n.t146 721.861
R8474 vp_n.n99 vp_n.t55 721.861
R8475 vp_n.n97 vp_n.t106 721.861
R8476 vp_n.n95 vp_n.t24 721.861
R8477 vp_n.n93 vp_n.t71 721.861
R8478 vp_n.n91 vp_n.t259 721.861
R8479 vp_n.n89 vp_n.t178 721.861
R8480 vp_n.n87 vp_n.t227 721.861
R8481 vp_n.n85 vp_n.t144 721.861
R8482 vp_n.n83 vp_n.t192 721.861
R8483 vp_n.n81 vp_n.t70 721.861
R8484 vp_n.n79 vp_n.t119 721.861
R8485 vp_n.n77 vp_n.t36 721.861
R8486 vp_n.n75 vp_n.t257 721.861
R8487 vp_n.n74 vp_n.t1 721.861
R8488 vp_n.n0 vp_n.t48 691.553
R8489 vp_n.n223 vp_n.t42 691.553
R8490 vp_n.n73 vp_n.t61 690.412
R8491 vp_n.n72 vp_n.t150 690.412
R8492 vp_n.n71 vp_n.t232 690.412
R8493 vp_n.n70 vp_n.t183 690.412
R8494 vp_n.n69 vp_n.t264 690.412
R8495 vp_n.n68 vp_n.t248 690.412
R8496 vp_n.n67 vp_n.t29 690.412
R8497 vp_n.n66 vp_n.t113 690.412
R8498 vp_n.n65 vp_n.t68 690.412
R8499 vp_n.n64 vp_n.t157 690.412
R8500 vp_n.n63 vp_n.t41 690.412
R8501 vp_n.n62 vp_n.t263 690.412
R8502 vp_n.n61 vp_n.t239 690.412
R8503 vp_n.n60 vp_n.t163 690.412
R8504 vp_n.n59 vp_n.t75 690.412
R8505 vp_n.n58 vp_n.t87 690.412
R8506 vp_n.n57 vp_n.t6 690.412
R8507 vp_n.n56 vp_n.t49 690.412
R8508 vp_n.n55 vp_n.t274 690.412
R8509 vp_n.n54 vp_n.t196 690.412
R8510 vp_n.n53 vp_n.t207 690.412
R8511 vp_n.n52 vp_n.t122 690.412
R8512 vp_n.n51 vp_n.t171 690.412
R8513 vp_n.n50 vp_n.t86 690.412
R8514 vp_n.n49 vp_n.t134 690.412
R8515 vp_n.n48 vp_n.t15 690.412
R8516 vp_n.n47 vp_n.t238 690.412
R8517 vp_n.n46 vp_n.t282 690.412
R8518 vp_n.n45 vp_n.t206 690.412
R8519 vp_n.n44 vp_n.t249 690.412
R8520 vp_n.n43 vp_n.t135 690.412
R8521 vp_n.n42 vp_n.t184 690.412
R8522 vp_n.n41 vp_n.t96 690.412
R8523 vp_n.n40 vp_n.t14 690.412
R8524 vp_n.n39 vp_n.t20 690.412
R8525 vp_n.n38 vp_n.t210 690.412
R8526 vp_n.n37 vp_n.t256 690.412
R8527 vp_n.n36 vp_n.t176 690.412
R8528 vp_n.n35 vp_n.t90 690.412
R8529 vp_n.n34 vp_n.t140 690.412
R8530 vp_n.n33 vp_n.t21 690.412
R8531 vp_n.n32 vp_n.t67 690.412
R8532 vp_n.n31 vp_n.t285 690.412
R8533 vp_n.n30 vp_n.t35 690.412
R8534 vp_n.n29 vp_n.t255 690.412
R8535 vp_n.n28 vp_n.t141 690.412
R8536 vp_n.n27 vp_n.t190 690.412
R8537 vp_n.n26 vp_n.t103 690.412
R8538 vp_n.n25 vp_n.t155 690.412
R8539 vp_n.n24 vp_n.t65 690.412
R8540 vp_n.n23 vp_n.t81 690.412
R8541 vp_n.n22 vp_n.t297 690.412
R8542 vp_n.n21 vp_n.t223 690.412
R8543 vp_n.n20 vp_n.t268 690.412
R8544 vp_n.n19 vp_n.t188 690.412
R8545 vp_n.n18 vp_n.t201 690.412
R8546 vp_n.n17 vp_n.t116 690.412
R8547 vp_n.n16 vp_n.t33 690.412
R8548 vp_n.n15 vp_n.t262 690.412
R8549 vp_n.n14 vp_n.t181 690.412
R8550 vp_n.n13 vp_n.t197 690.412
R8551 vp_n.n12 vp_n.t110 690.412
R8552 vp_n.n11 vp_n.t162 690.412
R8553 vp_n.n10 vp_n.t74 690.412
R8554 vp_n.n9 vp_n.t290 690.412
R8555 vp_n.n8 vp_n.t5 690.412
R8556 vp_n.n7 vp_n.t230 690.412
R8557 vp_n.n6 vp_n.t273 690.412
R8558 vp_n.n5 vp_n.t195 690.412
R8559 vp_n.n4 vp_n.t108 690.412
R8560 vp_n.n3 vp_n.t121 690.412
R8561 vp_n.n2 vp_n.t39 690.412
R8562 vp_n.n1 vp_n.t85 690.412
R8563 vp_n.n0 vp_n.t3 690.412
R8564 vp_n.n223 vp_n.t293 690.412
R8565 vp_n.n224 vp_n.t76 690.412
R8566 vp_n.n225 vp_n.t30 690.412
R8567 vp_n.n226 vp_n.t114 690.412
R8568 vp_n.n227 vp_n.t97 690.412
R8569 vp_n.n228 vp_n.t185 690.412
R8570 vp_n.n229 vp_n.t265 690.412
R8571 vp_n.n230 vp_n.t220 690.412
R8572 vp_n.n231 vp_n.t295 690.412
R8573 vp_n.n232 vp_n.t283 690.412
R8574 vp_n.n233 vp_n.t63 690.412
R8575 vp_n.n234 vp_n.t152 690.412
R8576 vp_n.n235 vp_n.t99 690.412
R8577 vp_n.n236 vp_n.t187 690.412
R8578 vp_n.n237 vp_n.t172 690.412
R8579 vp_n.n238 vp_n.t252 690.412
R8580 vp_n.n239 vp_n.t23 690.412
R8581 vp_n.n240 vp_n.t105 690.412
R8582 vp_n.n241 vp_n.t193 690.412
R8583 vp_n.n242 vp_n.t177 690.412
R8584 vp_n.n243 vp_n.t258 690.412
R8585 vp_n.n244 vp_n.t213 690.412
R8586 vp_n.n245 vp_n.t287 690.412
R8587 vp_n.n246 vp_n.t72 690.412
R8588 vp_n.n247 vp_n.t54 690.412
R8589 vp_n.n248 vp_n.t145 690.412
R8590 vp_n.n249 vp_n.t93 690.412
R8591 vp_n.n250 vp_n.t179 690.412
R8592 vp_n.n251 vp_n.t130 690.412
R8593 vp_n.n252 vp_n.t245 690.412
R8594 vp_n.n253 vp_n.t25 690.412
R8595 vp_n.n254 vp_n.t279 690.412
R8596 vp_n.n255 vp_n.t56 690.412
R8597 vp_n.n256 vp_n.t12 690.412
R8598 vp_n.n257 vp_n.t129 690.412
R8599 vp_n.n258 vp_n.t82 690.412
R8600 vp_n.n259 vp_n.t169 690.412
R8601 vp_n.n260 vp_n.t246 690.412
R8602 vp_n.n261 vp_n.t203 690.412
R8603 vp_n.n262 vp_n.t11 690.412
R8604 vp_n.n263 vp_n.t7 690.412
R8605 vp_n.n264 vp_n.t89 690.412
R8606 vp_n.n265 vp_n.t175 690.412
R8607 vp_n.n266 vp_n.t125 690.412
R8608 vp_n.n267 vp_n.t242 690.412
R8609 vp_n.n268 vp_n.t198 690.412
R8610 vp_n.n269 vp_n.t276 690.412
R8611 vp_n.n270 vp_n.t233 690.412
R8612 vp_n.n271 vp_n.t8 690.412
R8613 vp_n.n272 vp_n.t124 690.412
R8614 vp_n.n273 vp_n.t77 690.412
R8615 vp_n.n274 vp_n.t165 690.412
R8616 vp_n.n275 vp_n.t115 690.412
R8617 vp_n.n276 vp_n.t199 690.412
R8618 vp_n.n277 vp_n.t186 690.412
R8619 vp_n.n278 vp_n.t266 690.412
R8620 vp_n.n279 vp_n.t43 690.412
R8621 vp_n.n280 vp_n.t296 690.412
R8622 vp_n.n281 vp_n.t78 690.412
R8623 vp_n.n282 vp_n.t64 690.412
R8624 vp_n.n283 vp_n.t153 690.412
R8625 vp_n.n284 vp_n.t234 690.412
R8626 vp_n.n285 vp_n.t253 690.412
R8627 vp_n.n286 vp_n.t32 690.412
R8628 vp_n.n287 vp_n.t147 690.412
R8629 vp_n.n288 vp_n.t57 690.412
R8630 vp_n.n289 vp_n.t102 690.412
R8631 vp_n.n290 vp_n.t19 690.412
R8632 vp_n.n291 vp_n.t241 690.412
R8633 vp_n.n292 vp_n.t254 690.412
R8634 vp_n.n293 vp_n.t174 690.412
R8635 vp_n.n294 vp_n.t222 690.412
R8636 vp_n.n295 vp_n.t138 690.412
R8637 vp_n.n296 vp_n.t52 690.412
R8638 vp_n.n76 vp_n.n74 6.382
R8639 vp_n.n76 vp_n.n75 6.013
R8640 vp_n.n78 vp_n.n77 6.013
R8641 vp_n.n80 vp_n.n79 6.013
R8642 vp_n.n82 vp_n.n81 6.013
R8643 vp_n.n84 vp_n.n83 6.013
R8644 vp_n.n86 vp_n.n85 6.013
R8645 vp_n.n88 vp_n.n87 6.013
R8646 vp_n.n90 vp_n.n89 6.013
R8647 vp_n.n92 vp_n.n91 6.013
R8648 vp_n.n94 vp_n.n93 6.013
R8649 vp_n.n96 vp_n.n95 6.013
R8650 vp_n.n98 vp_n.n97 6.013
R8651 vp_n.n100 vp_n.n99 6.013
R8652 vp_n.n102 vp_n.n101 6.013
R8653 vp_n.n104 vp_n.n103 6.013
R8654 vp_n.n106 vp_n.n105 6.013
R8655 vp_n.n108 vp_n.n107 6.013
R8656 vp_n.n110 vp_n.n109 6.013
R8657 vp_n.n112 vp_n.n111 6.013
R8658 vp_n.n114 vp_n.n113 6.013
R8659 vp_n.n116 vp_n.n115 6.013
R8660 vp_n.n118 vp_n.n117 6.013
R8661 vp_n.n120 vp_n.n119 6.013
R8662 vp_n.n122 vp_n.n121 6.013
R8663 vp_n.n124 vp_n.n123 6.013
R8664 vp_n.n126 vp_n.n125 6.013
R8665 vp_n.n128 vp_n.n127 6.013
R8666 vp_n.n130 vp_n.n129 6.013
R8667 vp_n.n132 vp_n.n131 6.013
R8668 vp_n.n134 vp_n.n133 6.013
R8669 vp_n.n136 vp_n.n135 6.013
R8670 vp_n.n138 vp_n.n137 6.013
R8671 vp_n.n140 vp_n.n139 6.013
R8672 vp_n.n142 vp_n.n141 6.013
R8673 vp_n.n144 vp_n.n143 6.013
R8674 vp_n.n146 vp_n.n145 6.013
R8675 vp_n.n148 vp_n.n147 6.013
R8676 vp_n.n150 vp_n.n149 6.013
R8677 vp_n.n152 vp_n.n151 6.013
R8678 vp_n.n154 vp_n.n153 6.013
R8679 vp_n.n156 vp_n.n155 6.013
R8680 vp_n.n158 vp_n.n157 6.013
R8681 vp_n.n160 vp_n.n159 6.013
R8682 vp_n.n162 vp_n.n161 6.013
R8683 vp_n.n164 vp_n.n163 6.013
R8684 vp_n.n166 vp_n.n165 6.013
R8685 vp_n.n168 vp_n.n167 6.013
R8686 vp_n.n170 vp_n.n169 6.013
R8687 vp_n.n172 vp_n.n171 6.013
R8688 vp_n.n174 vp_n.n173 6.013
R8689 vp_n.n176 vp_n.n175 6.013
R8690 vp_n.n178 vp_n.n177 6.013
R8691 vp_n.n180 vp_n.n179 6.013
R8692 vp_n.n182 vp_n.n181 6.013
R8693 vp_n.n184 vp_n.n183 6.013
R8694 vp_n.n186 vp_n.n185 6.013
R8695 vp_n.n188 vp_n.n187 6.013
R8696 vp_n.n190 vp_n.n189 6.013
R8697 vp_n.n192 vp_n.n191 6.013
R8698 vp_n.n194 vp_n.n193 6.013
R8699 vp_n.n196 vp_n.n195 6.013
R8700 vp_n.n198 vp_n.n197 6.013
R8701 vp_n.n200 vp_n.n199 6.013
R8702 vp_n.n202 vp_n.n201 6.013
R8703 vp_n.n204 vp_n.n203 6.013
R8704 vp_n.n206 vp_n.n205 6.013
R8705 vp_n.n208 vp_n.n207 6.013
R8706 vp_n.n210 vp_n.n209 6.013
R8707 vp_n.n212 vp_n.n211 6.013
R8708 vp_n.n214 vp_n.n213 6.013
R8709 vp_n.n216 vp_n.n215 6.013
R8710 vp_n.n218 vp_n.n217 6.013
R8711 vp_n.n220 vp_n.n219 6.013
R8712 vp_n.n222 vp_n.n221 6.013
R8713 vp_n.n1 vp_n.n0 1.141
R8714 vp_n.n2 vp_n.n1 1.141
R8715 vp_n.n3 vp_n.n2 1.141
R8716 vp_n.n4 vp_n.n3 1.141
R8717 vp_n.n5 vp_n.n4 1.141
R8718 vp_n.n6 vp_n.n5 1.141
R8719 vp_n.n7 vp_n.n6 1.141
R8720 vp_n.n8 vp_n.n7 1.141
R8721 vp_n.n9 vp_n.n8 1.141
R8722 vp_n.n10 vp_n.n9 1.141
R8723 vp_n.n11 vp_n.n10 1.141
R8724 vp_n.n12 vp_n.n11 1.141
R8725 vp_n.n13 vp_n.n12 1.141
R8726 vp_n.n14 vp_n.n13 1.141
R8727 vp_n.n15 vp_n.n14 1.141
R8728 vp_n.n16 vp_n.n15 1.141
R8729 vp_n.n17 vp_n.n16 1.141
R8730 vp_n.n18 vp_n.n17 1.141
R8731 vp_n.n19 vp_n.n18 1.141
R8732 vp_n.n20 vp_n.n19 1.141
R8733 vp_n.n21 vp_n.n20 1.141
R8734 vp_n.n22 vp_n.n21 1.141
R8735 vp_n.n23 vp_n.n22 1.141
R8736 vp_n.n24 vp_n.n23 1.141
R8737 vp_n.n25 vp_n.n24 1.141
R8738 vp_n.n26 vp_n.n25 1.141
R8739 vp_n.n27 vp_n.n26 1.141
R8740 vp_n.n28 vp_n.n27 1.141
R8741 vp_n.n29 vp_n.n28 1.141
R8742 vp_n.n30 vp_n.n29 1.141
R8743 vp_n.n31 vp_n.n30 1.141
R8744 vp_n.n32 vp_n.n31 1.141
R8745 vp_n.n33 vp_n.n32 1.141
R8746 vp_n.n34 vp_n.n33 1.141
R8747 vp_n.n35 vp_n.n34 1.141
R8748 vp_n.n36 vp_n.n35 1.141
R8749 vp_n.n37 vp_n.n36 1.141
R8750 vp_n.n38 vp_n.n37 1.141
R8751 vp_n.n39 vp_n.n38 1.141
R8752 vp_n.n40 vp_n.n39 1.141
R8753 vp_n.n41 vp_n.n40 1.141
R8754 vp_n.n42 vp_n.n41 1.141
R8755 vp_n.n43 vp_n.n42 1.141
R8756 vp_n.n44 vp_n.n43 1.141
R8757 vp_n.n45 vp_n.n44 1.141
R8758 vp_n.n46 vp_n.n45 1.141
R8759 vp_n.n47 vp_n.n46 1.141
R8760 vp_n.n48 vp_n.n47 1.141
R8761 vp_n.n49 vp_n.n48 1.141
R8762 vp_n.n50 vp_n.n49 1.141
R8763 vp_n.n51 vp_n.n50 1.141
R8764 vp_n.n52 vp_n.n51 1.141
R8765 vp_n.n53 vp_n.n52 1.141
R8766 vp_n.n54 vp_n.n53 1.141
R8767 vp_n.n55 vp_n.n54 1.141
R8768 vp_n.n56 vp_n.n55 1.141
R8769 vp_n.n57 vp_n.n56 1.141
R8770 vp_n.n58 vp_n.n57 1.141
R8771 vp_n.n59 vp_n.n58 1.141
R8772 vp_n.n60 vp_n.n59 1.141
R8773 vp_n.n61 vp_n.n60 1.141
R8774 vp_n.n62 vp_n.n61 1.141
R8775 vp_n.n63 vp_n.n62 1.141
R8776 vp_n.n64 vp_n.n63 1.141
R8777 vp_n.n65 vp_n.n64 1.141
R8778 vp_n.n66 vp_n.n65 1.141
R8779 vp_n.n67 vp_n.n66 1.141
R8780 vp_n.n68 vp_n.n67 1.141
R8781 vp_n.n69 vp_n.n68 1.141
R8782 vp_n.n70 vp_n.n69 1.141
R8783 vp_n.n71 vp_n.n70 1.141
R8784 vp_n.n72 vp_n.n71 1.141
R8785 vp_n.n73 vp_n.n72 1.141
R8786 vp_n.n224 vp_n.n223 1.141
R8787 vp_n.n225 vp_n.n224 1.141
R8788 vp_n.n226 vp_n.n225 1.141
R8789 vp_n.n227 vp_n.n226 1.141
R8790 vp_n.n228 vp_n.n227 1.141
R8791 vp_n.n229 vp_n.n228 1.141
R8792 vp_n.n230 vp_n.n229 1.141
R8793 vp_n.n231 vp_n.n230 1.141
R8794 vp_n.n232 vp_n.n231 1.141
R8795 vp_n.n233 vp_n.n232 1.141
R8796 vp_n.n234 vp_n.n233 1.141
R8797 vp_n.n235 vp_n.n234 1.141
R8798 vp_n.n236 vp_n.n235 1.141
R8799 vp_n.n237 vp_n.n236 1.141
R8800 vp_n.n238 vp_n.n237 1.141
R8801 vp_n.n239 vp_n.n238 1.141
R8802 vp_n.n240 vp_n.n239 1.141
R8803 vp_n.n241 vp_n.n240 1.141
R8804 vp_n.n242 vp_n.n241 1.141
R8805 vp_n.n243 vp_n.n242 1.141
R8806 vp_n.n244 vp_n.n243 1.141
R8807 vp_n.n245 vp_n.n244 1.141
R8808 vp_n.n246 vp_n.n245 1.141
R8809 vp_n.n247 vp_n.n246 1.141
R8810 vp_n.n248 vp_n.n247 1.141
R8811 vp_n.n249 vp_n.n248 1.141
R8812 vp_n.n250 vp_n.n249 1.141
R8813 vp_n.n251 vp_n.n250 1.141
R8814 vp_n.n252 vp_n.n251 1.141
R8815 vp_n.n253 vp_n.n252 1.141
R8816 vp_n.n254 vp_n.n253 1.141
R8817 vp_n.n255 vp_n.n254 1.141
R8818 vp_n.n256 vp_n.n255 1.141
R8819 vp_n.n257 vp_n.n256 1.141
R8820 vp_n.n258 vp_n.n257 1.141
R8821 vp_n.n259 vp_n.n258 1.141
R8822 vp_n.n260 vp_n.n259 1.141
R8823 vp_n.n261 vp_n.n260 1.141
R8824 vp_n.n262 vp_n.n261 1.141
R8825 vp_n.n263 vp_n.n262 1.141
R8826 vp_n.n264 vp_n.n263 1.141
R8827 vp_n.n265 vp_n.n264 1.141
R8828 vp_n.n266 vp_n.n265 1.141
R8829 vp_n.n267 vp_n.n266 1.141
R8830 vp_n.n268 vp_n.n267 1.141
R8831 vp_n.n269 vp_n.n268 1.141
R8832 vp_n.n270 vp_n.n269 1.141
R8833 vp_n.n271 vp_n.n270 1.141
R8834 vp_n.n272 vp_n.n271 1.141
R8835 vp_n.n273 vp_n.n272 1.141
R8836 vp_n.n274 vp_n.n273 1.141
R8837 vp_n.n275 vp_n.n274 1.141
R8838 vp_n.n276 vp_n.n275 1.141
R8839 vp_n.n277 vp_n.n276 1.141
R8840 vp_n.n278 vp_n.n277 1.141
R8841 vp_n.n279 vp_n.n278 1.141
R8842 vp_n.n280 vp_n.n279 1.141
R8843 vp_n.n281 vp_n.n280 1.141
R8844 vp_n.n282 vp_n.n281 1.141
R8845 vp_n.n283 vp_n.n282 1.141
R8846 vp_n.n284 vp_n.n283 1.141
R8847 vp_n.n285 vp_n.n284 1.141
R8848 vp_n.n286 vp_n.n285 1.141
R8849 vp_n.n287 vp_n.n286 1.141
R8850 vp_n.n288 vp_n.n287 1.141
R8851 vp_n.n289 vp_n.n288 1.141
R8852 vp_n.n290 vp_n.n289 1.141
R8853 vp_n.n291 vp_n.n290 1.141
R8854 vp_n.n292 vp_n.n291 1.141
R8855 vp_n.n293 vp_n.n292 1.141
R8856 vp_n.n294 vp_n.n293 1.141
R8857 vp_n.n295 vp_n.n294 1.141
R8858 vp_n.n296 vp_n.n295 1.141
R8859 vp_n.n297 vp_n.n296 0.948
R8860 vp_n vp_n.n73 0.917
R8861 vp_n.n297 vp_n.n222 0.413
R8862 vp_n.n78 vp_n.n76 0.369
R8863 vp_n.n80 vp_n.n78 0.369
R8864 vp_n.n82 vp_n.n80 0.369
R8865 vp_n.n84 vp_n.n82 0.369
R8866 vp_n.n86 vp_n.n84 0.369
R8867 vp_n.n88 vp_n.n86 0.369
R8868 vp_n.n90 vp_n.n88 0.369
R8869 vp_n.n92 vp_n.n90 0.369
R8870 vp_n.n94 vp_n.n92 0.369
R8871 vp_n.n96 vp_n.n94 0.369
R8872 vp_n.n98 vp_n.n96 0.369
R8873 vp_n.n100 vp_n.n98 0.369
R8874 vp_n.n102 vp_n.n100 0.369
R8875 vp_n.n104 vp_n.n102 0.369
R8876 vp_n.n106 vp_n.n104 0.369
R8877 vp_n.n108 vp_n.n106 0.369
R8878 vp_n.n110 vp_n.n108 0.369
R8879 vp_n.n112 vp_n.n110 0.369
R8880 vp_n.n114 vp_n.n112 0.369
R8881 vp_n.n116 vp_n.n114 0.369
R8882 vp_n.n118 vp_n.n116 0.369
R8883 vp_n.n120 vp_n.n118 0.369
R8884 vp_n.n122 vp_n.n120 0.369
R8885 vp_n.n124 vp_n.n122 0.369
R8886 vp_n.n126 vp_n.n124 0.369
R8887 vp_n.n128 vp_n.n126 0.369
R8888 vp_n.n130 vp_n.n128 0.369
R8889 vp_n.n132 vp_n.n130 0.369
R8890 vp_n.n134 vp_n.n132 0.369
R8891 vp_n.n136 vp_n.n134 0.369
R8892 vp_n.n138 vp_n.n136 0.369
R8893 vp_n.n140 vp_n.n138 0.369
R8894 vp_n.n142 vp_n.n140 0.369
R8895 vp_n.n144 vp_n.n142 0.369
R8896 vp_n.n146 vp_n.n144 0.369
R8897 vp_n.n148 vp_n.n146 0.369
R8898 vp_n.n150 vp_n.n148 0.369
R8899 vp_n.n152 vp_n.n150 0.369
R8900 vp_n.n154 vp_n.n152 0.369
R8901 vp_n.n156 vp_n.n154 0.369
R8902 vp_n.n158 vp_n.n156 0.369
R8903 vp_n.n160 vp_n.n158 0.369
R8904 vp_n.n162 vp_n.n160 0.369
R8905 vp_n.n164 vp_n.n162 0.369
R8906 vp_n.n166 vp_n.n164 0.369
R8907 vp_n.n168 vp_n.n166 0.369
R8908 vp_n.n170 vp_n.n168 0.369
R8909 vp_n.n172 vp_n.n170 0.369
R8910 vp_n.n174 vp_n.n172 0.369
R8911 vp_n.n176 vp_n.n174 0.369
R8912 vp_n.n178 vp_n.n176 0.369
R8913 vp_n.n180 vp_n.n178 0.369
R8914 vp_n.n182 vp_n.n180 0.369
R8915 vp_n.n184 vp_n.n182 0.369
R8916 vp_n.n186 vp_n.n184 0.369
R8917 vp_n.n188 vp_n.n186 0.369
R8918 vp_n.n190 vp_n.n188 0.369
R8919 vp_n.n192 vp_n.n190 0.369
R8920 vp_n.n194 vp_n.n192 0.369
R8921 vp_n.n196 vp_n.n194 0.369
R8922 vp_n.n198 vp_n.n196 0.369
R8923 vp_n.n200 vp_n.n198 0.369
R8924 vp_n.n202 vp_n.n200 0.369
R8925 vp_n.n204 vp_n.n202 0.369
R8926 vp_n.n206 vp_n.n204 0.369
R8927 vp_n.n208 vp_n.n206 0.369
R8928 vp_n.n210 vp_n.n208 0.369
R8929 vp_n.n212 vp_n.n210 0.369
R8930 vp_n.n214 vp_n.n212 0.369
R8931 vp_n.n216 vp_n.n214 0.369
R8932 vp_n.n218 vp_n.n216 0.369
R8933 vp_n.n220 vp_n.n218 0.369
R8934 vp_n.n222 vp_n.n220 0.369
R8935 vp_n vp_n.n297 0.03
R8936 vss.n191 vss.t247 7.272
R8937 vss.n2 vss.t298 6.619
R8938 vss.n2 vss.t290 4.955
R8939 vss.n191 vss.t238 4.95
R8940 vss.n193 vss.t205 4.95
R8941 vss.n193 vss.t161 4.95
R8942 vss.n194 vss.t195 4.95
R8943 vss.n194 vss.t149 4.95
R8944 vss.n197 vss.t119 4.95
R8945 vss.n197 vss.t77 4.95
R8946 vss.n198 vss.t108 4.95
R8947 vss.n198 vss.t67 4.95
R8948 vss.n201 vss.t168 4.95
R8949 vss.n201 vss.t125 4.95
R8950 vss.n202 vss.t157 4.95
R8951 vss.n202 vss.t116 4.95
R8952 vss.n205 vss.t83 4.95
R8953 vss.n205 vss.t45 4.95
R8954 vss.n206 vss.t73 4.95
R8955 vss.n206 vss.t35 4.95
R8956 vss.n209 vss.t8 4.95
R8957 vss.n209 vss.t58 4.95
R8958 vss.n210 vss.t299 4.95
R8959 vss.n210 vss.t51 4.95
R8960 vss.n213 vss.t19 4.95
R8961 vss.n213 vss.t280 4.95
R8962 vss.n214 vss.t13 4.95
R8963 vss.n214 vss.t270 4.95
R8964 vss.n217 vss.t241 4.95
R8965 vss.n217 vss.t197 4.95
R8966 vss.n218 vss.t230 4.95
R8967 vss.n218 vss.t186 4.95
R8968 vss.n221 vss.t281 4.95
R8969 vss.n221 vss.t242 4.95
R8970 vss.n222 vss.t271 4.95
R8971 vss.n222 vss.t231 4.95
R8972 vss.n225 vss.t198 4.95
R8973 vss.n225 vss.t152 4.95
R8974 vss.n226 vss.t187 4.95
R8975 vss.n226 vss.t142 4.95
R8976 vss.n229 vss.t56 4.95
R8977 vss.n229 vss.t267 4.95
R8978 vss.n230 vss.t49 4.95
R8979 vss.n230 vss.t258 4.95
R8980 vss.n233 vss.t10 4.95
R8981 vss.n233 vss.t46 4.95
R8982 vss.n234 vss.t0 4.95
R8983 vss.n234 vss.t36 4.95
R8984 vss.n237 vss.t84 4.95
R8985 vss.n237 vss.t65 4.95
R8986 vss.n238 vss.t74 4.95
R8987 vss.n238 vss.t60 4.95
R8988 vss.n241 vss.t105 4.95
R8989 vss.n241 vss.t146 4.95
R8990 vss.n242 vss.t97 4.95
R8991 vss.n242 vss.t136 4.95
R8992 vss.n245 vss.t192 4.95
R8993 vss.n245 vss.t235 4.95
R8994 vss.n246 vss.t181 4.95
R8995 vss.n246 vss.t224 4.95
R8996 vss.n249 vss.t140 4.95
R8997 vss.n249 vss.t221 4.95
R8998 vss.n250 vss.t132 4.95
R8999 vss.n250 vss.t212 4.95
R9000 vss.n253 vss.t261 4.95
R9001 vss.n253 vss.t3 4.95
R9002 vss.n254 vss.t253 4.95
R9003 vss.n254 vss.t293 4.95
R9004 vss.n257 vss.t39 4.95
R9005 vss.n257 vss.t256 4.95
R9006 vss.n258 vss.t29 4.95
R9007 vss.n258 vss.t250 4.95
R9008 vss.n261 vss.t297 4.95
R9009 vss.n261 vss.t33 4.95
R9010 vss.n262 vss.t289 4.95
R9011 vss.n262 vss.t25 4.95
R9012 vss.n265 vss.t71 4.95
R9013 vss.n265 vss.t113 4.95
R9014 vss.n266 vss.t63 4.95
R9015 vss.n266 vss.t103 4.95
R9016 vss.n269 vss.t28 4.95
R9017 vss.n269 vss.t100 4.95
R9018 vss.n270 vss.t22 4.95
R9019 vss.n270 vss.t92 4.95
R9020 vss.n273 vss.t139 4.95
R9021 vss.n273 vss.t184 4.95
R9022 vss.n274 vss.t131 4.95
R9023 vss.n274 vss.t177 4.95
R9024 vss.n277 vss.t94 4.95
R9025 vss.n277 vss.t134 4.95
R9026 vss.n278 vss.t87 4.95
R9027 vss.n278 vss.t128 4.95
R9028 vss.n281 vss.t179 4.95
R9029 vss.n281 vss.t222 4.95
R9030 vss.n282 vss.t172 4.95
R9031 vss.n282 vss.t213 4.95
R9032 vss.n285 vss.t262 4.95
R9033 vss.n285 vss.t175 4.95
R9034 vss.n286 vss.t254 4.95
R9035 vss.n286 vss.t165 4.95
R9036 vss.n289 vss.t216 4.95
R9037 vss.n289 vss.t291 4.95
R9038 vss.n290 vss.t208 4.95
R9039 vss.n290 vss.t284 4.95
R9040 vss.n293 vss.t27 4.95
R9041 vss.n293 vss.t66 4.95
R9042 vss.n294 vss.t21 4.95
R9043 vss.n294 vss.t61 4.95
R9044 vss.n0 vss.t286 4.95
R9045 vss.n0 vss.t23 4.95
R9046 vss.n1 vss.t277 4.95
R9047 vss.n1 vss.t17 4.95
R9048 vss.n188 vss.t62 4.95
R9049 vss.n188 vss.t101 4.95
R9050 vss.n189 vss.t55 4.95
R9051 vss.n189 vss.t93 4.95
R9052 vss.n184 vss.t141 4.95
R9053 vss.n184 vss.t57 4.95
R9054 vss.n185 vss.t133 4.95
R9055 vss.n185 vss.t50 4.95
R9056 vss.n180 vss.t95 4.95
R9057 vss.n180 vss.t174 4.95
R9058 vss.n181 vss.t88 4.95
R9059 vss.n181 vss.t164 4.95
R9060 vss.n176 vss.t215 4.95
R9061 vss.n176 vss.t124 4.95
R9062 vss.n177 vss.t207 4.95
R9063 vss.n177 vss.t115 4.95
R9064 vss.n172 vss.t167 4.95
R9065 vss.n172 vss.t210 4.95
R9066 vss.n173 vss.t156 4.95
R9067 vss.n173 vss.t203 4.95
R9068 vss.n168 vss.t252 4.95
R9069 vss.n168 vss.t292 4.95
R9070 vss.n169 vss.t246 4.95
R9071 vss.n169 vss.t285 4.95
R9072 vss.n164 vss.t248 4.95
R9073 vss.n164 vss.t288 4.95
R9074 vss.n165 vss.t239 4.95
R9075 vss.n165 vss.t279 4.95
R9076 vss.n160 vss.t24 4.95
R9077 vss.n160 vss.t96 4.95
R9078 vss.n161 vss.t18 4.95
R9079 vss.n161 vss.t89 4.95
R9080 vss.n156 vss.t135 4.95
R9081 vss.n156 vss.t53 4.95
R9082 vss.n157 vss.t129 4.95
R9083 vss.n157 vss.t43 4.95
R9084 vss.n152 vss.t90 4.95
R9085 vss.n152 vss.t130 4.95
R9086 vss.n153 vss.t81 4.95
R9087 vss.n153 vss.t123 4.95
R9088 vss.n148 vss.t176 4.95
R9089 vss.n148 vss.t217 4.95
R9090 vss.n149 vss.t166 4.95
R9091 vss.n149 vss.t209 4.95
R9092 vss.n144 vss.t126 4.95
R9093 vss.n144 vss.t170 4.95
R9094 vss.n145 vss.t117 4.95
R9095 vss.n145 vss.t159 4.95
R9096 vss.n140 vss.t211 4.95
R9097 vss.n140 vss.t287 4.95
R9098 vss.n141 vss.t204 4.95
R9099 vss.n141 vss.t278 4.95
R9100 vss.n136 vss.t199 4.95
R9101 vss.n136 vss.t243 4.95
R9102 vss.n137 vss.t188 4.95
R9103 vss.n137 vss.t232 4.95
R9104 vss.n132 vss.t282 4.95
R9105 vss.n132 vss.t20 4.95
R9106 vss.n133 vss.t272 4.95
R9107 vss.n133 vss.t14 4.95
R9108 vss.n128 vss.t59 4.95
R9109 vss.n128 vss.t274 4.95
R9110 vss.n129 vss.t52 4.95
R9111 vss.n129 vss.t264 4.95
R9112 vss.n124 vss.t15 4.95
R9113 vss.n124 vss.t54 4.95
R9114 vss.n125 vss.t7 4.95
R9115 vss.n125 vss.t44 4.95
R9116 vss.n120 vss.t91 4.95
R9117 vss.n120 vss.t169 4.95
R9118 vss.n121 vss.t82 4.95
R9119 vss.n121 vss.t158 4.95
R9120 vss.n116 vss.t78 4.95
R9121 vss.n116 vss.t120 4.95
R9122 vss.n117 vss.t68 4.95
R9123 vss.n117 vss.t109 4.95
R9124 vss.n112 vss.t162 4.95
R9125 vss.n112 vss.t206 4.95
R9126 vss.n113 vss.t150 4.95
R9127 vss.n113 vss.t196 4.95
R9128 vss.n108 vss.t249 4.95
R9129 vss.n108 vss.t154 4.95
R9130 vss.n109 vss.t240 4.95
R9131 vss.n109 vss.t144 4.95
R9132 vss.n104 vss.t201 4.95
R9133 vss.n104 vss.t245 4.95
R9134 vss.n105 vss.t190 4.95
R9135 vss.n105 vss.t234 4.95
R9136 vss.n100 vss.t283 4.95
R9137 vss.n100 vss.t227 4.95
R9138 vss.n101 vss.t273 4.95
R9139 vss.n101 vss.t218 4.95
R9140 vss.n96 vss.t268 4.95
R9141 vss.n96 vss.t12 4.95
R9142 vss.n97 vss.t259 4.95
R9143 vss.n97 vss.t2 4.95
R9144 vss.n92 vss.t48 4.95
R9145 vss.n92 vss.t86 4.95
R9146 vss.n93 vss.t38 4.95
R9147 vss.n93 vss.t76 4.95
R9148 vss.n88 vss.t5 4.95
R9149 vss.n88 vss.t41 4.95
R9150 vss.n89 vss.t295 4.95
R9151 vss.n89 vss.t31 4.95
R9152 vss.n84 vss.t80 4.95
R9153 vss.n84 vss.t122 4.95
R9154 vss.n85 vss.t70 4.95
R9155 vss.n85 vss.t111 4.95
R9156 vss.n80 vss.t163 4.95
R9157 vss.n80 vss.t106 4.95
R9158 vss.n81 vss.t151 4.95
R9159 vss.n81 vss.t98 4.95
R9160 vss.n76 vss.t148 4.95
R9161 vss.n76 vss.t194 4.95
R9162 vss.n77 vss.t138 4.95
R9163 vss.n77 vss.t183 4.95
R9164 vss.n72 vss.t237 4.95
R9165 vss.n72 vss.t276 4.95
R9166 vss.n73 vss.t226 4.95
R9167 vss.n73 vss.t266 4.95
R9168 vss.n68 vss.t11 4.95
R9169 vss.n68 vss.t47 4.95
R9170 vss.n69 vss.t1 4.95
R9171 vss.n69 vss.t37 4.95
R9172 vss.n64 vss.t85 4.95
R9173 vss.n64 vss.t127 4.95
R9174 vss.n65 vss.t75 4.95
R9175 vss.n65 vss.t118 4.95
R9176 vss.n60 vss.t171 4.95
R9177 vss.n60 vss.t112 4.95
R9178 vss.n61 vss.t160 4.95
R9179 vss.n61 vss.t102 4.95
R9180 vss.n56 vss.t153 4.95
R9181 vss.n56 vss.t200 4.95
R9182 vss.n57 vss.t143 4.95
R9183 vss.n57 vss.t189 4.95
R9184 vss.n52 vss.t244 4.95
R9185 vss.n52 vss.t147 4.95
R9186 vss.n53 vss.t233 4.95
R9187 vss.n53 vss.t137 4.95
R9188 vss.n48 vss.t193 4.95
R9189 vss.n48 vss.t236 4.95
R9190 vss.n49 vss.t182 4.95
R9191 vss.n49 vss.t225 4.95
R9192 vss.n44 vss.t275 4.95
R9193 vss.n44 vss.t16 4.95
R9194 vss.n45 vss.t265 4.95
R9195 vss.n45 vss.t9 4.95
R9196 vss.n40 vss.t228 4.95
R9197 vss.n40 vss.t4 4.95
R9198 vss.n41 vss.t220 4.95
R9199 vss.n41 vss.t294 4.95
R9200 vss.n36 vss.t40 4.95
R9201 vss.n36 vss.t79 4.95
R9202 vss.n37 vss.t30 4.95
R9203 vss.n37 vss.t69 4.95
R9204 vss.n32 vss.t121 4.95
R9205 vss.n32 vss.t34 4.95
R9206 vss.n33 vss.t110 4.95
R9207 vss.n33 vss.t26 4.95
R9208 vss.n28 vss.t72 4.95
R9209 vss.n28 vss.t114 4.95
R9210 vss.n29 vss.t64 4.95
R9211 vss.n29 vss.t104 4.95
R9212 vss.n24 vss.t155 4.95
R9213 vss.n24 vss.t202 4.95
R9214 vss.n25 vss.t145 4.95
R9215 vss.n25 vss.t191 4.95
R9216 vss.n20 vss.t107 4.95
R9217 vss.n20 vss.t185 4.95
R9218 vss.n21 vss.t99 4.95
R9219 vss.n21 vss.t178 4.95
R9220 vss.n16 vss.t229 4.95
R9221 vss.n16 vss.t269 4.95
R9222 vss.n17 vss.t219 4.95
R9223 vss.n17 vss.t260 4.95
R9224 vss.n12 vss.t180 4.95
R9225 vss.n12 vss.t223 4.95
R9226 vss.n13 vss.t173 4.95
R9227 vss.n13 vss.t214 4.95
R9228 vss.n8 vss.t263 4.95
R9229 vss.n8 vss.t6 4.95
R9230 vss.n9 vss.t255 4.95
R9231 vss.n9 vss.t296 4.95
R9232 vss.n4 vss.t42 4.95
R9233 vss.n4 vss.t257 4.95
R9234 vss.n5 vss.t32 4.95
R9235 vss.n5 vss.t251 4.95
R9236 vss.n192 vss.n191 1.3
R9237 vss.n3 vss.n2 0.989
R9238 vss.n194 vss.n193 0.76
R9239 vss.n198 vss.n197 0.76
R9240 vss.n202 vss.n201 0.76
R9241 vss.n206 vss.n205 0.76
R9242 vss.n210 vss.n209 0.76
R9243 vss.n214 vss.n213 0.76
R9244 vss.n218 vss.n217 0.76
R9245 vss.n222 vss.n221 0.76
R9246 vss.n226 vss.n225 0.76
R9247 vss.n230 vss.n229 0.76
R9248 vss.n234 vss.n233 0.76
R9249 vss.n238 vss.n237 0.76
R9250 vss.n242 vss.n241 0.76
R9251 vss.n246 vss.n245 0.76
R9252 vss.n250 vss.n249 0.76
R9253 vss.n254 vss.n253 0.76
R9254 vss.n258 vss.n257 0.76
R9255 vss.n262 vss.n261 0.76
R9256 vss.n266 vss.n265 0.76
R9257 vss.n270 vss.n269 0.76
R9258 vss.n274 vss.n273 0.76
R9259 vss.n278 vss.n277 0.76
R9260 vss.n282 vss.n281 0.76
R9261 vss.n286 vss.n285 0.76
R9262 vss.n290 vss.n289 0.76
R9263 vss.n294 vss.n293 0.76
R9264 vss.n1 vss.n0 0.76
R9265 vss.n189 vss.n188 0.76
R9266 vss.n185 vss.n184 0.76
R9267 vss.n181 vss.n180 0.76
R9268 vss.n177 vss.n176 0.76
R9269 vss.n173 vss.n172 0.76
R9270 vss.n169 vss.n168 0.76
R9271 vss.n165 vss.n164 0.76
R9272 vss.n161 vss.n160 0.76
R9273 vss.n157 vss.n156 0.76
R9274 vss.n153 vss.n152 0.76
R9275 vss.n149 vss.n148 0.76
R9276 vss.n145 vss.n144 0.76
R9277 vss.n141 vss.n140 0.76
R9278 vss.n137 vss.n136 0.76
R9279 vss.n133 vss.n132 0.76
R9280 vss.n129 vss.n128 0.76
R9281 vss.n125 vss.n124 0.76
R9282 vss.n121 vss.n120 0.76
R9283 vss.n117 vss.n116 0.76
R9284 vss.n113 vss.n112 0.76
R9285 vss.n109 vss.n108 0.76
R9286 vss.n105 vss.n104 0.76
R9287 vss.n101 vss.n100 0.76
R9288 vss.n97 vss.n96 0.76
R9289 vss.n93 vss.n92 0.76
R9290 vss.n89 vss.n88 0.76
R9291 vss.n85 vss.n84 0.76
R9292 vss.n81 vss.n80 0.76
R9293 vss.n77 vss.n76 0.76
R9294 vss.n73 vss.n72 0.76
R9295 vss.n69 vss.n68 0.76
R9296 vss.n65 vss.n64 0.76
R9297 vss.n61 vss.n60 0.76
R9298 vss.n57 vss.n56 0.76
R9299 vss.n53 vss.n52 0.76
R9300 vss.n49 vss.n48 0.76
R9301 vss.n45 vss.n44 0.76
R9302 vss.n41 vss.n40 0.76
R9303 vss.n37 vss.n36 0.76
R9304 vss.n33 vss.n32 0.76
R9305 vss.n29 vss.n28 0.76
R9306 vss.n25 vss.n24 0.76
R9307 vss.n21 vss.n20 0.76
R9308 vss.n17 vss.n16 0.76
R9309 vss.n13 vss.n12 0.76
R9310 vss.n9 vss.n8 0.76
R9311 vss.n5 vss.n4 0.76
R9312 vss.n195 vss.n194 0.419
R9313 vss.n199 vss.n198 0.419
R9314 vss.n203 vss.n202 0.419
R9315 vss.n207 vss.n206 0.419
R9316 vss.n211 vss.n210 0.419
R9317 vss.n215 vss.n214 0.419
R9318 vss.n219 vss.n218 0.419
R9319 vss.n223 vss.n222 0.419
R9320 vss.n227 vss.n226 0.419
R9321 vss.n231 vss.n230 0.419
R9322 vss.n235 vss.n234 0.419
R9323 vss.n239 vss.n238 0.419
R9324 vss.n243 vss.n242 0.419
R9325 vss.n247 vss.n246 0.419
R9326 vss.n251 vss.n250 0.419
R9327 vss.n255 vss.n254 0.419
R9328 vss.n259 vss.n258 0.419
R9329 vss.n263 vss.n262 0.419
R9330 vss.n267 vss.n266 0.419
R9331 vss.n271 vss.n270 0.419
R9332 vss.n275 vss.n274 0.419
R9333 vss.n279 vss.n278 0.419
R9334 vss.n283 vss.n282 0.419
R9335 vss.n287 vss.n286 0.419
R9336 vss.n291 vss.n290 0.419
R9337 vss.n295 vss.n294 0.419
R9338 vss vss.n1 0.419
R9339 vss.n190 vss.n189 0.419
R9340 vss.n186 vss.n185 0.419
R9341 vss.n182 vss.n181 0.419
R9342 vss.n178 vss.n177 0.419
R9343 vss.n174 vss.n173 0.419
R9344 vss.n170 vss.n169 0.419
R9345 vss.n166 vss.n165 0.419
R9346 vss.n162 vss.n161 0.419
R9347 vss.n158 vss.n157 0.419
R9348 vss.n154 vss.n153 0.419
R9349 vss.n150 vss.n149 0.419
R9350 vss.n146 vss.n145 0.419
R9351 vss.n142 vss.n141 0.419
R9352 vss.n138 vss.n137 0.419
R9353 vss.n134 vss.n133 0.419
R9354 vss.n130 vss.n129 0.419
R9355 vss.n126 vss.n125 0.419
R9356 vss.n122 vss.n121 0.419
R9357 vss.n118 vss.n117 0.419
R9358 vss.n114 vss.n113 0.419
R9359 vss.n110 vss.n109 0.419
R9360 vss.n106 vss.n105 0.419
R9361 vss.n102 vss.n101 0.419
R9362 vss.n98 vss.n97 0.419
R9363 vss.n94 vss.n93 0.419
R9364 vss.n90 vss.n89 0.419
R9365 vss.n86 vss.n85 0.419
R9366 vss.n82 vss.n81 0.419
R9367 vss.n78 vss.n77 0.419
R9368 vss.n74 vss.n73 0.419
R9369 vss.n70 vss.n69 0.419
R9370 vss.n66 vss.n65 0.419
R9371 vss.n62 vss.n61 0.419
R9372 vss.n58 vss.n57 0.419
R9373 vss.n54 vss.n53 0.419
R9374 vss.n50 vss.n49 0.419
R9375 vss.n46 vss.n45 0.419
R9376 vss.n42 vss.n41 0.419
R9377 vss.n38 vss.n37 0.419
R9378 vss.n34 vss.n33 0.419
R9379 vss.n30 vss.n29 0.419
R9380 vss.n26 vss.n25 0.419
R9381 vss.n22 vss.n21 0.419
R9382 vss.n18 vss.n17 0.419
R9383 vss.n14 vss.n13 0.419
R9384 vss.n10 vss.n9 0.419
R9385 vss.n6 vss.n5 0.419
R9386 vss.n10 vss.n6 0.002
R9387 vss.n14 vss.n10 0.002
R9388 vss.n18 vss.n14 0.002
R9389 vss.n22 vss.n18 0.002
R9390 vss.n26 vss.n22 0.002
R9391 vss.n30 vss.n26 0.002
R9392 vss.n34 vss.n30 0.002
R9393 vss.n38 vss.n34 0.002
R9394 vss.n42 vss.n38 0.002
R9395 vss.n46 vss.n42 0.002
R9396 vss.n50 vss.n46 0.002
R9397 vss.n54 vss.n50 0.002
R9398 vss.n58 vss.n54 0.002
R9399 vss.n62 vss.n58 0.002
R9400 vss.n66 vss.n62 0.002
R9401 vss.n70 vss.n66 0.002
R9402 vss.n74 vss.n70 0.002
R9403 vss.n78 vss.n74 0.002
R9404 vss.n82 vss.n78 0.002
R9405 vss.n86 vss.n82 0.002
R9406 vss.n90 vss.n86 0.002
R9407 vss.n94 vss.n90 0.002
R9408 vss.n98 vss.n94 0.002
R9409 vss.n102 vss.n98 0.002
R9410 vss.n106 vss.n102 0.002
R9411 vss.n110 vss.n106 0.002
R9412 vss.n114 vss.n110 0.002
R9413 vss.n118 vss.n114 0.002
R9414 vss.n122 vss.n118 0.002
R9415 vss.n126 vss.n122 0.002
R9416 vss.n130 vss.n126 0.002
R9417 vss.n134 vss.n130 0.002
R9418 vss.n138 vss.n134 0.002
R9419 vss.n142 vss.n138 0.002
R9420 vss.n146 vss.n142 0.002
R9421 vss.n150 vss.n146 0.002
R9422 vss.n154 vss.n150 0.002
R9423 vss.n158 vss.n154 0.002
R9424 vss.n162 vss.n158 0.002
R9425 vss.n166 vss.n162 0.002
R9426 vss.n170 vss.n166 0.002
R9427 vss.n174 vss.n170 0.002
R9428 vss.n178 vss.n174 0.002
R9429 vss.n182 vss.n178 0.002
R9430 vss.n186 vss.n182 0.002
R9431 vss.n190 vss.n186 0.002
R9432 vss vss.n190 0.002
R9433 vss vss.n295 0.002
R9434 vss.n295 vss.n291 0.002
R9435 vss.n291 vss.n287 0.002
R9436 vss.n287 vss.n283 0.002
R9437 vss.n283 vss.n279 0.002
R9438 vss.n279 vss.n275 0.002
R9439 vss.n275 vss.n271 0.002
R9440 vss.n271 vss.n267 0.002
R9441 vss.n267 vss.n263 0.002
R9442 vss.n263 vss.n259 0.002
R9443 vss.n259 vss.n255 0.002
R9444 vss.n255 vss.n251 0.002
R9445 vss.n251 vss.n247 0.002
R9446 vss.n247 vss.n243 0.002
R9447 vss.n243 vss.n239 0.002
R9448 vss.n239 vss.n235 0.002
R9449 vss.n235 vss.n231 0.002
R9450 vss.n231 vss.n227 0.002
R9451 vss.n227 vss.n223 0.002
R9452 vss.n223 vss.n219 0.002
R9453 vss.n219 vss.n215 0.002
R9454 vss.n215 vss.n211 0.002
R9455 vss.n211 vss.n207 0.002
R9456 vss.n207 vss.n203 0.002
R9457 vss.n203 vss.n199 0.002
R9458 vss.n199 vss.n195 0.002
R9459 vss.n10 vss.n7 0.001
R9460 vss.n14 vss.n11 0.001
R9461 vss.n18 vss.n15 0.001
R9462 vss.n22 vss.n19 0.001
R9463 vss.n26 vss.n23 0.001
R9464 vss.n30 vss.n27 0.001
R9465 vss.n34 vss.n31 0.001
R9466 vss.n38 vss.n35 0.001
R9467 vss.n42 vss.n39 0.001
R9468 vss.n46 vss.n43 0.001
R9469 vss.n50 vss.n47 0.001
R9470 vss.n54 vss.n51 0.001
R9471 vss.n58 vss.n55 0.001
R9472 vss.n62 vss.n59 0.001
R9473 vss.n66 vss.n63 0.001
R9474 vss.n70 vss.n67 0.001
R9475 vss.n74 vss.n71 0.001
R9476 vss.n78 vss.n75 0.001
R9477 vss.n82 vss.n79 0.001
R9478 vss.n86 vss.n83 0.001
R9479 vss.n90 vss.n87 0.001
R9480 vss.n94 vss.n91 0.001
R9481 vss.n98 vss.n95 0.001
R9482 vss.n102 vss.n99 0.001
R9483 vss.n106 vss.n103 0.001
R9484 vss.n110 vss.n107 0.001
R9485 vss.n114 vss.n111 0.001
R9486 vss.n118 vss.n115 0.001
R9487 vss.n122 vss.n119 0.001
R9488 vss.n126 vss.n123 0.001
R9489 vss.n130 vss.n127 0.001
R9490 vss.n134 vss.n131 0.001
R9491 vss.n138 vss.n135 0.001
R9492 vss.n142 vss.n139 0.001
R9493 vss.n146 vss.n143 0.001
R9494 vss.n154 vss.n151 0.001
R9495 vss.n158 vss.n155 0.001
R9496 vss.n162 vss.n159 0.001
R9497 vss.n166 vss.n163 0.001
R9498 vss.n170 vss.n167 0.001
R9499 vss.n174 vss.n171 0.001
R9500 vss.n178 vss.n175 0.001
R9501 vss.n182 vss.n179 0.001
R9502 vss.n186 vss.n183 0.001
R9503 vss.n190 vss.n187 0.001
R9504 vss.n296 vss 0.001
R9505 vss.n295 vss.n292 0.001
R9506 vss.n291 vss.n288 0.001
R9507 vss.n287 vss.n284 0.001
R9508 vss.n283 vss.n280 0.001
R9509 vss.n279 vss.n276 0.001
R9510 vss.n275 vss.n272 0.001
R9511 vss.n271 vss.n268 0.001
R9512 vss.n267 vss.n264 0.001
R9513 vss.n263 vss.n260 0.001
R9514 vss.n259 vss.n256 0.001
R9515 vss.n255 vss.n252 0.001
R9516 vss.n251 vss.n248 0.001
R9517 vss.n247 vss.n244 0.001
R9518 vss.n243 vss.n240 0.001
R9519 vss.n239 vss.n236 0.001
R9520 vss.n235 vss.n232 0.001
R9521 vss.n231 vss.n228 0.001
R9522 vss.n227 vss.n224 0.001
R9523 vss.n223 vss.n220 0.001
R9524 vss.n219 vss.n216 0.001
R9525 vss.n215 vss.n212 0.001
R9526 vss.n211 vss.n208 0.001
R9527 vss.n207 vss.n204 0.001
R9528 vss.n203 vss.n200 0.001
R9529 vss.n199 vss.n196 0.001
R9530 vss.n150 vss.n147 0.001
R9531 vss.n195 vss.n192 0.001
R9532 vss.n6 vss.n3 0.001
C4 vp_p vss 345.28fF
C5 out_p vss 1048.44fF
C6 vp_n vss 211.11fF
C7 vdd vss 1210.44fF
C8 vp_n.n0 vss 1.10fF $ **FLOATING
C9 vp_n.n73 vss 1.25fF $ **FLOATING
C10 vp_n.n76 vss 1.56fF $ **FLOATING
C11 vp_n.n78 vss 1.00fF $ **FLOATING
C12 vp_n.n80 vss 1.00fF $ **FLOATING
C13 vp_n.n82 vss 1.00fF $ **FLOATING
C14 vp_n.n84 vss 1.00fF $ **FLOATING
C15 vp_n.n86 vss 1.00fF $ **FLOATING
C16 vp_n.n88 vss 1.00fF $ **FLOATING
C17 vp_n.n90 vss 1.00fF $ **FLOATING
C18 vp_n.n92 vss 1.00fF $ **FLOATING
C19 vp_n.n94 vss 1.00fF $ **FLOATING
C20 vp_n.n96 vss 1.00fF $ **FLOATING
C21 vp_n.n98 vss 1.00fF $ **FLOATING
C22 vp_n.n100 vss 1.00fF $ **FLOATING
C23 vp_n.n102 vss 1.00fF $ **FLOATING
C24 vp_n.n104 vss 1.00fF $ **FLOATING
C25 vp_n.n106 vss 1.00fF $ **FLOATING
C26 vp_n.n108 vss 1.00fF $ **FLOATING
C27 vp_n.n110 vss 1.00fF $ **FLOATING
C28 vp_n.n112 vss 1.00fF $ **FLOATING
C29 vp_n.n114 vss 1.00fF $ **FLOATING
C30 vp_n.n116 vss 1.00fF $ **FLOATING
C31 vp_n.n118 vss 1.00fF $ **FLOATING
C32 vp_n.n120 vss 1.00fF $ **FLOATING
C33 vp_n.n122 vss 1.00fF $ **FLOATING
C34 vp_n.n124 vss 1.00fF $ **FLOATING
C35 vp_n.n126 vss 1.00fF $ **FLOATING
C36 vp_n.n128 vss 1.00fF $ **FLOATING
C37 vp_n.n130 vss 1.00fF $ **FLOATING
C38 vp_n.n132 vss 1.00fF $ **FLOATING
C39 vp_n.n134 vss 1.00fF $ **FLOATING
C40 vp_n.n136 vss 1.00fF $ **FLOATING
C41 vp_n.n138 vss 1.00fF $ **FLOATING
C42 vp_n.n140 vss 1.00fF $ **FLOATING
C43 vp_n.n142 vss 1.00fF $ **FLOATING
C44 vp_n.n144 vss 1.00fF $ **FLOATING
C45 vp_n.n146 vss 1.00fF $ **FLOATING
C46 vp_n.n148 vss 1.00fF $ **FLOATING
C47 vp_n.n150 vss 1.00fF $ **FLOATING
C48 vp_n.n152 vss 1.00fF $ **FLOATING
C49 vp_n.n154 vss 1.00fF $ **FLOATING
C50 vp_n.n156 vss 1.00fF $ **FLOATING
C51 vp_n.n158 vss 1.00fF $ **FLOATING
C52 vp_n.n160 vss 1.00fF $ **FLOATING
C53 vp_n.n162 vss 1.00fF $ **FLOATING
C54 vp_n.n164 vss 1.00fF $ **FLOATING
C55 vp_n.n166 vss 1.00fF $ **FLOATING
C56 vp_n.n168 vss 1.00fF $ **FLOATING
C57 vp_n.n170 vss 1.00fF $ **FLOATING
C58 vp_n.n172 vss 1.00fF $ **FLOATING
C59 vp_n.n174 vss 1.00fF $ **FLOATING
C60 vp_n.n176 vss 1.00fF $ **FLOATING
C61 vp_n.n178 vss 1.00fF $ **FLOATING
C62 vp_n.n180 vss 1.00fF $ **FLOATING
C63 vp_n.n182 vss 1.00fF $ **FLOATING
C64 vp_n.n184 vss 1.00fF $ **FLOATING
C65 vp_n.n186 vss 1.00fF $ **FLOATING
C66 vp_n.n188 vss 1.00fF $ **FLOATING
C67 vp_n.n190 vss 1.00fF $ **FLOATING
C68 vp_n.n192 vss 1.00fF $ **FLOATING
C69 vp_n.n194 vss 1.00fF $ **FLOATING
C70 vp_n.n196 vss 1.00fF $ **FLOATING
C71 vp_n.n198 vss 1.00fF $ **FLOATING
C72 vp_n.n200 vss 1.00fF $ **FLOATING
C73 vp_n.n202 vss 1.00fF $ **FLOATING
C74 vp_n.n204 vss 1.00fF $ **FLOATING
C75 vp_n.n206 vss 1.00fF $ **FLOATING
C76 vp_n.n208 vss 1.00fF $ **FLOATING
C77 vp_n.n210 vss 1.00fF $ **FLOATING
C78 vp_n.n212 vss 1.00fF $ **FLOATING
C79 vp_n.n214 vss 1.00fF $ **FLOATING
C80 vp_n.n216 vss 1.00fF $ **FLOATING
C81 vp_n.n218 vss 1.00fF $ **FLOATING
C82 vp_n.n220 vss 1.00fF $ **FLOATING
C83 vp_n.n222 vss 1.06fF $ **FLOATING
C84 vp_n.n223 vss 1.16fF $ **FLOATING
C85 vp_n.n296 vss 1.58fF $ **FLOATING
C86 vp_n.n297 vss 12.55fF $ **FLOATING
C87 vdd.n0 vss 4.21fF $ **FLOATING
C88 vdd.n1 vss 4.42fF $ **FLOATING
C89 vdd.n2 vss 4.42fF $ **FLOATING
C90 vdd.n3 vss 4.42fF $ **FLOATING
C91 vdd.n4 vss 4.53fF $ **FLOATING
C92 vdd.n5 vss 4.53fF $ **FLOATING
C93 vdd.n6 vss 4.42fF $ **FLOATING
C94 vdd.n7 vss 4.42fF $ **FLOATING
C95 vdd.n8 vss 4.42fF $ **FLOATING
C96 vdd.n9 vss 4.02fF $ **FLOATING
C97 vdd.n12 vss 5.67fF $ **FLOATING
C98 vdd.n13 vss 3.04fF $ **FLOATING
C99 vdd.n14 vss 3.04fF $ **FLOATING
C100 vdd.n15 vss 3.08fF $ **FLOATING
C101 vdd.n16 vss 3.14fF $ **FLOATING
C102 vdd.n17 vss 3.04fF $ **FLOATING
C103 vdd.n18 vss 3.04fF $ **FLOATING
C104 vdd.n19 vss 3.04fF $ **FLOATING
C105 vdd.n20 vss 2.69fF $ **FLOATING
C106 vdd.n21 vss 4.63fF $ **FLOATING
C107 vdd.n22 vss 4.21fF $ **FLOATING
C108 vdd.n23 vss 4.42fF $ **FLOATING
C109 vdd.n24 vss 4.42fF $ **FLOATING
C110 vdd.n25 vss 4.42fF $ **FLOATING
C111 vdd.n26 vss 4.53fF $ **FLOATING
C112 vdd.n27 vss 4.53fF $ **FLOATING
C113 vdd.n28 vss 4.42fF $ **FLOATING
C114 vdd.n29 vss 4.42fF $ **FLOATING
C115 vdd.n30 vss 4.42fF $ **FLOATING
C116 vdd.n31 vss 4.02fF $ **FLOATING
C117 vdd.n35 vss 61.16fF $ **FLOATING
C118 vdd.n38 vss 4.21fF $ **FLOATING
C119 vdd.n39 vss 4.42fF $ **FLOATING
C120 vdd.n40 vss 4.42fF $ **FLOATING
C121 vdd.n41 vss 4.42fF $ **FLOATING
C122 vdd.n42 vss 4.53fF $ **FLOATING
C123 vdd.n43 vss 4.53fF $ **FLOATING
C124 vdd.n44 vss 4.42fF $ **FLOATING
C125 vdd.n45 vss 4.42fF $ **FLOATING
C126 vdd.n46 vss 4.42fF $ **FLOATING
C127 vdd.n47 vss 4.02fF $ **FLOATING
C128 vdd.n49 vss 32.58fF $ **FLOATING
C129 vdd.n50 vss 4.21fF $ **FLOATING
C130 vdd.n51 vss 4.42fF $ **FLOATING
C131 vdd.n52 vss 4.42fF $ **FLOATING
C132 vdd.n53 vss 4.42fF $ **FLOATING
C133 vdd.n54 vss 4.53fF $ **FLOATING
C134 vdd.n55 vss 4.53fF $ **FLOATING
C135 vdd.n56 vss 4.42fF $ **FLOATING
C136 vdd.n57 vss 4.42fF $ **FLOATING
C137 vdd.n58 vss 4.42fF $ **FLOATING
C138 vdd.n59 vss 4.02fF $ **FLOATING
C139 vdd.n63 vss 32.58fF $ **FLOATING
C140 vdd.n66 vss 4.21fF $ **FLOATING
C141 vdd.n67 vss 4.42fF $ **FLOATING
C142 vdd.n68 vss 4.42fF $ **FLOATING
C143 vdd.n69 vss 4.42fF $ **FLOATING
C144 vdd.n70 vss 4.53fF $ **FLOATING
C145 vdd.n71 vss 4.53fF $ **FLOATING
C146 vdd.n72 vss 4.42fF $ **FLOATING
C147 vdd.n73 vss 4.42fF $ **FLOATING
C148 vdd.n74 vss 4.42fF $ **FLOATING
C149 vdd.n75 vss 4.02fF $ **FLOATING
C150 vdd.n77 vss 32.58fF $ **FLOATING
C151 vdd.n78 vss 4.21fF $ **FLOATING
C152 vdd.n79 vss 4.42fF $ **FLOATING
C153 vdd.n80 vss 4.42fF $ **FLOATING
C154 vdd.n81 vss 4.42fF $ **FLOATING
C155 vdd.n82 vss 4.53fF $ **FLOATING
C156 vdd.n83 vss 4.53fF $ **FLOATING
C157 vdd.n84 vss 4.42fF $ **FLOATING
C158 vdd.n85 vss 4.42fF $ **FLOATING
C159 vdd.n86 vss 4.42fF $ **FLOATING
C160 vdd.n87 vss 4.02fF $ **FLOATING
C161 vdd.n91 vss 32.58fF $ **FLOATING
C162 vdd.n94 vss 4.21fF $ **FLOATING
C163 vdd.n95 vss 4.42fF $ **FLOATING
C164 vdd.n96 vss 4.42fF $ **FLOATING
C165 vdd.n97 vss 4.42fF $ **FLOATING
C166 vdd.n98 vss 4.53fF $ **FLOATING
C167 vdd.n99 vss 4.53fF $ **FLOATING
C168 vdd.n100 vss 4.42fF $ **FLOATING
C169 vdd.n101 vss 4.42fF $ **FLOATING
C170 vdd.n102 vss 4.42fF $ **FLOATING
C171 vdd.n103 vss 4.02fF $ **FLOATING
C172 vdd.n105 vss 32.58fF $ **FLOATING
C173 vdd.n106 vss 4.21fF $ **FLOATING
C174 vdd.n107 vss 4.42fF $ **FLOATING
C175 vdd.n108 vss 4.42fF $ **FLOATING
C176 vdd.n109 vss 4.42fF $ **FLOATING
C177 vdd.n110 vss 4.53fF $ **FLOATING
C178 vdd.n111 vss 4.53fF $ **FLOATING
C179 vdd.n112 vss 4.42fF $ **FLOATING
C180 vdd.n113 vss 4.42fF $ **FLOATING
C181 vdd.n114 vss 4.42fF $ **FLOATING
C182 vdd.n115 vss 4.02fF $ **FLOATING
C183 vdd.n119 vss 32.58fF $ **FLOATING
C184 vdd.n122 vss 4.21fF $ **FLOATING
C185 vdd.n123 vss 4.42fF $ **FLOATING
C186 vdd.n124 vss 4.42fF $ **FLOATING
C187 vdd.n125 vss 4.42fF $ **FLOATING
C188 vdd.n126 vss 4.53fF $ **FLOATING
C189 vdd.n127 vss 4.53fF $ **FLOATING
C190 vdd.n128 vss 4.42fF $ **FLOATING
C191 vdd.n129 vss 4.42fF $ **FLOATING
C192 vdd.n130 vss 4.42fF $ **FLOATING
C193 vdd.n131 vss 4.02fF $ **FLOATING
C194 vdd.n133 vss 32.58fF $ **FLOATING
C195 vdd.n134 vss 4.21fF $ **FLOATING
C196 vdd.n135 vss 4.42fF $ **FLOATING
C197 vdd.n136 vss 4.42fF $ **FLOATING
C198 vdd.n137 vss 4.42fF $ **FLOATING
C199 vdd.n138 vss 4.53fF $ **FLOATING
C200 vdd.n139 vss 4.53fF $ **FLOATING
C201 vdd.n140 vss 4.42fF $ **FLOATING
C202 vdd.n141 vss 4.42fF $ **FLOATING
C203 vdd.n142 vss 4.42fF $ **FLOATING
C204 vdd.n143 vss 4.02fF $ **FLOATING
C205 vdd.n147 vss 32.58fF $ **FLOATING
C206 vdd.n150 vss 4.21fF $ **FLOATING
C207 vdd.n151 vss 4.42fF $ **FLOATING
C208 vdd.n152 vss 4.42fF $ **FLOATING
C209 vdd.n153 vss 4.42fF $ **FLOATING
C210 vdd.n154 vss 4.53fF $ **FLOATING
C211 vdd.n155 vss 4.53fF $ **FLOATING
C212 vdd.n156 vss 4.42fF $ **FLOATING
C213 vdd.n157 vss 4.42fF $ **FLOATING
C214 vdd.n158 vss 4.42fF $ **FLOATING
C215 vdd.n159 vss 4.02fF $ **FLOATING
C216 vdd.n161 vss 32.58fF $ **FLOATING
C217 vdd.n162 vss 4.21fF $ **FLOATING
C218 vdd.n163 vss 4.42fF $ **FLOATING
C219 vdd.n164 vss 4.42fF $ **FLOATING
C220 vdd.n165 vss 4.42fF $ **FLOATING
C221 vdd.n166 vss 4.53fF $ **FLOATING
C222 vdd.n167 vss 4.53fF $ **FLOATING
C223 vdd.n168 vss 4.42fF $ **FLOATING
C224 vdd.n169 vss 4.42fF $ **FLOATING
C225 vdd.n170 vss 4.42fF $ **FLOATING
C226 vdd.n171 vss 4.02fF $ **FLOATING
C227 vdd.n175 vss 32.58fF $ **FLOATING
C228 vdd.n178 vss 4.21fF $ **FLOATING
C229 vdd.n179 vss 4.42fF $ **FLOATING
C230 vdd.n180 vss 4.42fF $ **FLOATING
C231 vdd.n181 vss 4.42fF $ **FLOATING
C232 vdd.n182 vss 4.53fF $ **FLOATING
C233 vdd.n183 vss 4.53fF $ **FLOATING
C234 vdd.n184 vss 4.42fF $ **FLOATING
C235 vdd.n185 vss 4.42fF $ **FLOATING
C236 vdd.n186 vss 4.42fF $ **FLOATING
C237 vdd.n187 vss 4.02fF $ **FLOATING
C238 vdd.n189 vss 32.58fF $ **FLOATING
C239 vdd.n190 vss 4.21fF $ **FLOATING
C240 vdd.n191 vss 4.42fF $ **FLOATING
C241 vdd.n192 vss 4.42fF $ **FLOATING
C242 vdd.n193 vss 4.42fF $ **FLOATING
C243 vdd.n194 vss 4.53fF $ **FLOATING
C244 vdd.n195 vss 4.53fF $ **FLOATING
C245 vdd.n196 vss 4.42fF $ **FLOATING
C246 vdd.n197 vss 4.42fF $ **FLOATING
C247 vdd.n198 vss 4.42fF $ **FLOATING
C248 vdd.n199 vss 4.02fF $ **FLOATING
C249 vdd.n203 vss 32.58fF $ **FLOATING
C250 vdd.n206 vss 4.21fF $ **FLOATING
C251 vdd.n207 vss 4.42fF $ **FLOATING
C252 vdd.n208 vss 4.42fF $ **FLOATING
C253 vdd.n209 vss 4.42fF $ **FLOATING
C254 vdd.n210 vss 4.53fF $ **FLOATING
C255 vdd.n211 vss 4.53fF $ **FLOATING
C256 vdd.n212 vss 4.42fF $ **FLOATING
C257 vdd.n213 vss 4.42fF $ **FLOATING
C258 vdd.n214 vss 4.42fF $ **FLOATING
C259 vdd.n215 vss 4.02fF $ **FLOATING
C260 vdd.n217 vss 32.58fF $ **FLOATING
C261 vdd.n218 vss 4.21fF $ **FLOATING
C262 vdd.n219 vss 4.42fF $ **FLOATING
C263 vdd.n220 vss 4.42fF $ **FLOATING
C264 vdd.n221 vss 4.42fF $ **FLOATING
C265 vdd.n222 vss 4.53fF $ **FLOATING
C266 vdd.n223 vss 4.53fF $ **FLOATING
C267 vdd.n224 vss 4.42fF $ **FLOATING
C268 vdd.n225 vss 4.42fF $ **FLOATING
C269 vdd.n226 vss 4.42fF $ **FLOATING
C270 vdd.n227 vss 4.02fF $ **FLOATING
C271 vdd.n231 vss 32.58fF $ **FLOATING
C272 vdd.n234 vss 4.21fF $ **FLOATING
C273 vdd.n235 vss 4.42fF $ **FLOATING
C274 vdd.n236 vss 4.42fF $ **FLOATING
C275 vdd.n237 vss 4.42fF $ **FLOATING
C276 vdd.n238 vss 4.53fF $ **FLOATING
C277 vdd.n239 vss 4.53fF $ **FLOATING
C278 vdd.n240 vss 4.42fF $ **FLOATING
C279 vdd.n241 vss 4.42fF $ **FLOATING
C280 vdd.n242 vss 4.42fF $ **FLOATING
C281 vdd.n243 vss 4.02fF $ **FLOATING
C282 vdd.n245 vss 32.58fF $ **FLOATING
C283 vdd.n246 vss 4.21fF $ **FLOATING
C284 vdd.n247 vss 4.42fF $ **FLOATING
C285 vdd.n248 vss 4.42fF $ **FLOATING
C286 vdd.n249 vss 4.42fF $ **FLOATING
C287 vdd.n250 vss 4.53fF $ **FLOATING
C288 vdd.n251 vss 4.53fF $ **FLOATING
C289 vdd.n252 vss 4.42fF $ **FLOATING
C290 vdd.n253 vss 4.42fF $ **FLOATING
C291 vdd.n254 vss 4.42fF $ **FLOATING
C292 vdd.n255 vss 4.02fF $ **FLOATING
C293 vdd.n259 vss 32.58fF $ **FLOATING
C294 vdd.n262 vss 4.21fF $ **FLOATING
C295 vdd.n263 vss 4.42fF $ **FLOATING
C296 vdd.n264 vss 4.42fF $ **FLOATING
C297 vdd.n265 vss 4.42fF $ **FLOATING
C298 vdd.n266 vss 4.53fF $ **FLOATING
C299 vdd.n267 vss 4.53fF $ **FLOATING
C300 vdd.n268 vss 4.42fF $ **FLOATING
C301 vdd.n269 vss 4.42fF $ **FLOATING
C302 vdd.n270 vss 4.42fF $ **FLOATING
C303 vdd.n271 vss 4.02fF $ **FLOATING
C304 vdd.n273 vss 32.58fF $ **FLOATING
C305 vdd.n274 vss 4.21fF $ **FLOATING
C306 vdd.n275 vss 4.42fF $ **FLOATING
C307 vdd.n276 vss 4.42fF $ **FLOATING
C308 vdd.n277 vss 4.42fF $ **FLOATING
C309 vdd.n278 vss 4.53fF $ **FLOATING
C310 vdd.n279 vss 4.53fF $ **FLOATING
C311 vdd.n280 vss 4.42fF $ **FLOATING
C312 vdd.n281 vss 4.42fF $ **FLOATING
C313 vdd.n282 vss 4.42fF $ **FLOATING
C314 vdd.n283 vss 4.02fF $ **FLOATING
C315 vdd.n287 vss 32.58fF $ **FLOATING
C316 vdd.n290 vss 4.21fF $ **FLOATING
C317 vdd.n291 vss 4.42fF $ **FLOATING
C318 vdd.n292 vss 4.42fF $ **FLOATING
C319 vdd.n293 vss 4.42fF $ **FLOATING
C320 vdd.n294 vss 4.53fF $ **FLOATING
C321 vdd.n295 vss 4.53fF $ **FLOATING
C322 vdd.n296 vss 4.42fF $ **FLOATING
C323 vdd.n297 vss 4.42fF $ **FLOATING
C324 vdd.n298 vss 4.42fF $ **FLOATING
C325 vdd.n299 vss 4.02fF $ **FLOATING
C326 vdd.n301 vss 32.58fF $ **FLOATING
C327 vdd.n302 vss 4.21fF $ **FLOATING
C328 vdd.n303 vss 4.42fF $ **FLOATING
C329 vdd.n304 vss 4.42fF $ **FLOATING
C330 vdd.n305 vss 4.42fF $ **FLOATING
C331 vdd.n306 vss 4.53fF $ **FLOATING
C332 vdd.n307 vss 4.53fF $ **FLOATING
C333 vdd.n308 vss 4.42fF $ **FLOATING
C334 vdd.n309 vss 4.42fF $ **FLOATING
C335 vdd.n310 vss 4.42fF $ **FLOATING
C336 vdd.n311 vss 4.02fF $ **FLOATING
C337 vdd.n315 vss 32.58fF $ **FLOATING
C338 vdd.n318 vss 4.21fF $ **FLOATING
C339 vdd.n319 vss 4.42fF $ **FLOATING
C340 vdd.n320 vss 4.42fF $ **FLOATING
C341 vdd.n321 vss 4.42fF $ **FLOATING
C342 vdd.n322 vss 4.53fF $ **FLOATING
C343 vdd.n323 vss 4.53fF $ **FLOATING
C344 vdd.n324 vss 4.42fF $ **FLOATING
C345 vdd.n325 vss 4.42fF $ **FLOATING
C346 vdd.n326 vss 4.42fF $ **FLOATING
C347 vdd.n327 vss 4.02fF $ **FLOATING
C348 vdd.n329 vss 32.58fF $ **FLOATING
C349 vdd.n330 vss 4.21fF $ **FLOATING
C350 vdd.n331 vss 4.42fF $ **FLOATING
C351 vdd.n332 vss 4.42fF $ **FLOATING
C352 vdd.n333 vss 4.42fF $ **FLOATING
C353 vdd.n334 vss 4.53fF $ **FLOATING
C354 vdd.n335 vss 4.53fF $ **FLOATING
C355 vdd.n336 vss 4.42fF $ **FLOATING
C356 vdd.n337 vss 4.42fF $ **FLOATING
C357 vdd.n338 vss 4.42fF $ **FLOATING
C358 vdd.n339 vss 4.02fF $ **FLOATING
C359 vdd.n343 vss 32.58fF $ **FLOATING
C360 vdd.n346 vss 4.21fF $ **FLOATING
C361 vdd.n347 vss 4.42fF $ **FLOATING
C362 vdd.n348 vss 4.42fF $ **FLOATING
C363 vdd.n349 vss 4.42fF $ **FLOATING
C364 vdd.n350 vss 4.53fF $ **FLOATING
C365 vdd.n351 vss 4.53fF $ **FLOATING
C366 vdd.n352 vss 4.42fF $ **FLOATING
C367 vdd.n353 vss 4.42fF $ **FLOATING
C368 vdd.n354 vss 4.42fF $ **FLOATING
C369 vdd.n355 vss 4.02fF $ **FLOATING
C370 vdd.n357 vss 32.58fF $ **FLOATING
C371 vdd.n358 vss 4.21fF $ **FLOATING
C372 vdd.n359 vss 4.42fF $ **FLOATING
C373 vdd.n360 vss 4.42fF $ **FLOATING
C374 vdd.n361 vss 4.42fF $ **FLOATING
C375 vdd.n362 vss 4.53fF $ **FLOATING
C376 vdd.n363 vss 4.53fF $ **FLOATING
C377 vdd.n364 vss 4.42fF $ **FLOATING
C378 vdd.n365 vss 4.42fF $ **FLOATING
C379 vdd.n366 vss 4.42fF $ **FLOATING
C380 vdd.n367 vss 4.02fF $ **FLOATING
C381 vdd.n371 vss 32.58fF $ **FLOATING
C382 vdd.n374 vss 4.21fF $ **FLOATING
C383 vdd.n375 vss 4.42fF $ **FLOATING
C384 vdd.n376 vss 4.42fF $ **FLOATING
C385 vdd.n377 vss 4.42fF $ **FLOATING
C386 vdd.n378 vss 4.53fF $ **FLOATING
C387 vdd.n379 vss 4.53fF $ **FLOATING
C388 vdd.n380 vss 4.42fF $ **FLOATING
C389 vdd.n381 vss 4.42fF $ **FLOATING
C390 vdd.n382 vss 4.42fF $ **FLOATING
C391 vdd.n383 vss 4.02fF $ **FLOATING
C392 vdd.n385 vss 32.58fF $ **FLOATING
C393 vdd.n386 vss 4.21fF $ **FLOATING
C394 vdd.n387 vss 4.42fF $ **FLOATING
C395 vdd.n388 vss 4.42fF $ **FLOATING
C396 vdd.n389 vss 4.42fF $ **FLOATING
C397 vdd.n390 vss 4.53fF $ **FLOATING
C398 vdd.n391 vss 4.53fF $ **FLOATING
C399 vdd.n392 vss 4.42fF $ **FLOATING
C400 vdd.n393 vss 4.42fF $ **FLOATING
C401 vdd.n394 vss 4.42fF $ **FLOATING
C402 vdd.n395 vss 4.02fF $ **FLOATING
C403 vdd.n399 vss 32.58fF $ **FLOATING
C404 vdd.n402 vss 4.21fF $ **FLOATING
C405 vdd.n403 vss 4.42fF $ **FLOATING
C406 vdd.n404 vss 4.42fF $ **FLOATING
C407 vdd.n405 vss 4.42fF $ **FLOATING
C408 vdd.n406 vss 4.53fF $ **FLOATING
C409 vdd.n407 vss 4.53fF $ **FLOATING
C410 vdd.n408 vss 4.42fF $ **FLOATING
C411 vdd.n409 vss 4.42fF $ **FLOATING
C412 vdd.n410 vss 4.42fF $ **FLOATING
C413 vdd.n411 vss 4.02fF $ **FLOATING
C414 vdd.n413 vss 32.58fF $ **FLOATING
C415 vdd.n414 vss 4.21fF $ **FLOATING
C416 vdd.n415 vss 4.42fF $ **FLOATING
C417 vdd.n416 vss 4.42fF $ **FLOATING
C418 vdd.n417 vss 4.42fF $ **FLOATING
C419 vdd.n418 vss 4.53fF $ **FLOATING
C420 vdd.n419 vss 4.53fF $ **FLOATING
C421 vdd.n420 vss 4.42fF $ **FLOATING
C422 vdd.n421 vss 4.42fF $ **FLOATING
C423 vdd.n422 vss 4.42fF $ **FLOATING
C424 vdd.n423 vss 4.02fF $ **FLOATING
C425 vdd.n427 vss 32.58fF $ **FLOATING
C426 vdd.n430 vss 4.21fF $ **FLOATING
C427 vdd.n431 vss 4.42fF $ **FLOATING
C428 vdd.n432 vss 4.42fF $ **FLOATING
C429 vdd.n433 vss 4.42fF $ **FLOATING
C430 vdd.n434 vss 4.53fF $ **FLOATING
C431 vdd.n435 vss 4.53fF $ **FLOATING
C432 vdd.n436 vss 4.42fF $ **FLOATING
C433 vdd.n437 vss 4.42fF $ **FLOATING
C434 vdd.n438 vss 4.42fF $ **FLOATING
C435 vdd.n439 vss 4.02fF $ **FLOATING
C436 vdd.n441 vss 32.58fF $ **FLOATING
C437 vdd.n442 vss 4.21fF $ **FLOATING
C438 vdd.n443 vss 4.42fF $ **FLOATING
C439 vdd.n444 vss 4.42fF $ **FLOATING
C440 vdd.n445 vss 4.42fF $ **FLOATING
C441 vdd.n446 vss 4.53fF $ **FLOATING
C442 vdd.n447 vss 4.53fF $ **FLOATING
C443 vdd.n448 vss 4.42fF $ **FLOATING
C444 vdd.n449 vss 4.42fF $ **FLOATING
C445 vdd.n450 vss 4.42fF $ **FLOATING
C446 vdd.n451 vss 4.02fF $ **FLOATING
C447 vdd.n455 vss 32.58fF $ **FLOATING
C448 vdd.n458 vss 4.21fF $ **FLOATING
C449 vdd.n459 vss 4.42fF $ **FLOATING
C450 vdd.n460 vss 4.42fF $ **FLOATING
C451 vdd.n461 vss 4.42fF $ **FLOATING
C452 vdd.n462 vss 4.53fF $ **FLOATING
C453 vdd.n463 vss 4.53fF $ **FLOATING
C454 vdd.n464 vss 4.42fF $ **FLOATING
C455 vdd.n465 vss 4.42fF $ **FLOATING
C456 vdd.n466 vss 4.42fF $ **FLOATING
C457 vdd.n467 vss 4.02fF $ **FLOATING
C458 vdd.n469 vss 32.58fF $ **FLOATING
C459 vdd.n470 vss 4.21fF $ **FLOATING
C460 vdd.n471 vss 4.42fF $ **FLOATING
C461 vdd.n472 vss 4.42fF $ **FLOATING
C462 vdd.n473 vss 4.42fF $ **FLOATING
C463 vdd.n474 vss 4.53fF $ **FLOATING
C464 vdd.n475 vss 4.53fF $ **FLOATING
C465 vdd.n476 vss 4.42fF $ **FLOATING
C466 vdd.n477 vss 4.42fF $ **FLOATING
C467 vdd.n478 vss 4.42fF $ **FLOATING
C468 vdd.n479 vss 4.02fF $ **FLOATING
C469 vdd.n483 vss 32.58fF $ **FLOATING
C470 vdd.n486 vss 4.21fF $ **FLOATING
C471 vdd.n487 vss 4.42fF $ **FLOATING
C472 vdd.n488 vss 4.42fF $ **FLOATING
C473 vdd.n489 vss 4.42fF $ **FLOATING
C474 vdd.n490 vss 4.53fF $ **FLOATING
C475 vdd.n491 vss 4.53fF $ **FLOATING
C476 vdd.n492 vss 4.42fF $ **FLOATING
C477 vdd.n493 vss 4.42fF $ **FLOATING
C478 vdd.n494 vss 4.42fF $ **FLOATING
C479 vdd.n495 vss 4.02fF $ **FLOATING
C480 vdd.n497 vss 32.58fF $ **FLOATING
C481 vdd.n498 vss 4.21fF $ **FLOATING
C482 vdd.n499 vss 4.42fF $ **FLOATING
C483 vdd.n500 vss 4.42fF $ **FLOATING
C484 vdd.n501 vss 4.42fF $ **FLOATING
C485 vdd.n502 vss 4.53fF $ **FLOATING
C486 vdd.n503 vss 4.53fF $ **FLOATING
C487 vdd.n504 vss 4.42fF $ **FLOATING
C488 vdd.n505 vss 4.42fF $ **FLOATING
C489 vdd.n506 vss 4.42fF $ **FLOATING
C490 vdd.n507 vss 4.02fF $ **FLOATING
C491 vdd.n511 vss 32.58fF $ **FLOATING
C492 vdd.n513 vss 4.21fF $ **FLOATING
C493 vdd.n514 vss 4.42fF $ **FLOATING
C494 vdd.n515 vss 4.42fF $ **FLOATING
C495 vdd.n516 vss 4.42fF $ **FLOATING
C496 vdd.n517 vss 4.53fF $ **FLOATING
C497 vdd.n518 vss 4.53fF $ **FLOATING
C498 vdd.n519 vss 4.42fF $ **FLOATING
C499 vdd.n520 vss 4.42fF $ **FLOATING
C500 vdd.n521 vss 4.42fF $ **FLOATING
C501 vdd.n522 vss 4.02fF $ **FLOATING
C502 vdd.n524 vss 32.58fF $ **FLOATING
C503 vdd.n525 vss 13.80fF $ **FLOATING
C504 vdd.n526 vss 5.45fF $ **FLOATING
C505 vdd.n527 vss 5.45fF $ **FLOATING
C506 vdd.n528 vss 6.37fF $ **FLOATING
C507 vdd.n529 vss 6.37fF $ **FLOATING
C508 vdd.n530 vss 11.61fF $ **FLOATING
C509 vdd.n531 vss 13.80fF $ **FLOATING
C510 vdd.n532 vss 5.44fF $ **FLOATING
C511 vdd.n533 vss 5.44fF $ **FLOATING
C512 vdd.n534 vss 6.35fF $ **FLOATING
C513 vdd.n535 vss 6.35fF $ **FLOATING
C514 vdd.n536 vss 11.61fF $ **FLOATING
C515 vdd.n537 vss 6.44fF $ **FLOATING
C516 vdd.n539 vss 32.33fF $ **FLOATING
C517 vdd.n540 vss 4.21fF $ **FLOATING
C518 vdd.n541 vss 4.42fF $ **FLOATING
C519 vdd.n542 vss 4.42fF $ **FLOATING
C520 vdd.n543 vss 4.42fF $ **FLOATING
C521 vdd.n544 vss 4.53fF $ **FLOATING
C522 vdd.n545 vss 4.53fF $ **FLOATING
C523 vdd.n546 vss 4.42fF $ **FLOATING
C524 vdd.n547 vss 4.42fF $ **FLOATING
C525 vdd.n548 vss 4.42fF $ **FLOATING
C526 vdd.n549 vss 4.03fF $ **FLOATING
C527 vdd.n550 vss 1.01fF $ **FLOATING
C528 vdd.n551 vss 32.83fF $ **FLOATING
C529 vdd.n554 vss 4.21fF $ **FLOATING
C530 vdd.n555 vss 4.42fF $ **FLOATING
C531 vdd.n556 vss 4.42fF $ **FLOATING
C532 vdd.n557 vss 4.42fF $ **FLOATING
C533 vdd.n558 vss 4.53fF $ **FLOATING
C534 vdd.n559 vss 4.53fF $ **FLOATING
C535 vdd.n560 vss 4.42fF $ **FLOATING
C536 vdd.n561 vss 4.42fF $ **FLOATING
C537 vdd.n562 vss 4.42fF $ **FLOATING
C538 vdd.n563 vss 4.02fF $ **FLOATING
C539 vdd.n565 vss 32.58fF $ **FLOATING
C540 vdd.n566 vss 4.21fF $ **FLOATING
C541 vdd.n567 vss 4.42fF $ **FLOATING
C542 vdd.n568 vss 4.42fF $ **FLOATING
C543 vdd.n569 vss 4.42fF $ **FLOATING
C544 vdd.n570 vss 4.53fF $ **FLOATING
C545 vdd.n571 vss 4.53fF $ **FLOATING
C546 vdd.n572 vss 4.42fF $ **FLOATING
C547 vdd.n573 vss 4.42fF $ **FLOATING
C548 vdd.n574 vss 4.42fF $ **FLOATING
C549 vdd.n575 vss 4.02fF $ **FLOATING
C550 vdd.n579 vss 32.58fF $ **FLOATING
C551 vdd.n582 vss 4.21fF $ **FLOATING
C552 vdd.n583 vss 4.42fF $ **FLOATING
C553 vdd.n584 vss 4.42fF $ **FLOATING
C554 vdd.n585 vss 4.42fF $ **FLOATING
C555 vdd.n586 vss 4.53fF $ **FLOATING
C556 vdd.n587 vss 4.53fF $ **FLOATING
C557 vdd.n588 vss 4.42fF $ **FLOATING
C558 vdd.n589 vss 4.42fF $ **FLOATING
C559 vdd.n590 vss 4.42fF $ **FLOATING
C560 vdd.n591 vss 4.02fF $ **FLOATING
C561 vdd.n593 vss 32.58fF $ **FLOATING
C562 vdd.n594 vss 4.21fF $ **FLOATING
C563 vdd.n595 vss 4.42fF $ **FLOATING
C564 vdd.n596 vss 4.42fF $ **FLOATING
C565 vdd.n597 vss 4.42fF $ **FLOATING
C566 vdd.n598 vss 4.53fF $ **FLOATING
C567 vdd.n599 vss 4.53fF $ **FLOATING
C568 vdd.n600 vss 4.42fF $ **FLOATING
C569 vdd.n601 vss 4.42fF $ **FLOATING
C570 vdd.n602 vss 4.42fF $ **FLOATING
C571 vdd.n603 vss 4.02fF $ **FLOATING
C572 vdd.n607 vss 32.58fF $ **FLOATING
C573 vdd.n608 vss 3.29fF $ **FLOATING
C574 vdd.n609 vss 1.87fF $ **FLOATING
C575 vdd.n610 vss 1.87fF $ **FLOATING
C576 vdd.n611 vss 1.91fF $ **FLOATING
C577 vdd.n612 vss 1.96fF $ **FLOATING
C578 vdd.n613 vss 1.92fF $ **FLOATING
C579 vdd.n614 vss 1.92fF $ **FLOATING
C580 vdd.n615 vss 1.92fF $ **FLOATING
C581 vdd.n616 vss 1.83fF $ **FLOATING
C582 vdd.n617 vss 4.83fF $ **FLOATING
C583 vdd.n618 vss 4.21fF $ **FLOATING
C584 vdd.n619 vss 4.42fF $ **FLOATING
C585 vdd.n620 vss 4.42fF $ **FLOATING
C586 vdd.n621 vss 4.42fF $ **FLOATING
C587 vdd.n622 vss 4.53fF $ **FLOATING
C588 vdd.n623 vss 4.53fF $ **FLOATING
C589 vdd.n624 vss 4.42fF $ **FLOATING
C590 vdd.n625 vss 4.42fF $ **FLOATING
C591 vdd.n626 vss 4.42fF $ **FLOATING
C592 vdd.n627 vss 4.02fF $ **FLOATING
C593 vdd.n629 vss 52.58fF $ **FLOATING
C594 vdd.n630 vss 4.21fF $ **FLOATING
C595 vdd.n631 vss 4.42fF $ **FLOATING
C596 vdd.n632 vss 4.42fF $ **FLOATING
C597 vdd.n633 vss 4.42fF $ **FLOATING
C598 vdd.n634 vss 4.53fF $ **FLOATING
C599 vdd.n635 vss 4.53fF $ **FLOATING
C600 vdd.n636 vss 4.42fF $ **FLOATING
C601 vdd.n637 vss 4.42fF $ **FLOATING
C602 vdd.n638 vss 4.42fF $ **FLOATING
C603 vdd.n639 vss 4.02fF $ **FLOATING
C604 vdd.n643 vss 32.58fF $ **FLOATING
C605 vdd.n646 vss 4.21fF $ **FLOATING
C606 vdd.n647 vss 4.42fF $ **FLOATING
C607 vdd.n648 vss 4.42fF $ **FLOATING
C608 vdd.n649 vss 4.42fF $ **FLOATING
C609 vdd.n650 vss 4.53fF $ **FLOATING
C610 vdd.n651 vss 4.53fF $ **FLOATING
C611 vdd.n652 vss 4.42fF $ **FLOATING
C612 vdd.n653 vss 4.42fF $ **FLOATING
C613 vdd.n654 vss 4.42fF $ **FLOATING
C614 vdd.n655 vss 4.02fF $ **FLOATING
C615 vdd.n657 vss 32.58fF $ **FLOATING
C616 vdd.n658 vss 4.21fF $ **FLOATING
C617 vdd.n659 vss 4.42fF $ **FLOATING
C618 vdd.n660 vss 4.42fF $ **FLOATING
C619 vdd.n661 vss 4.42fF $ **FLOATING
C620 vdd.n662 vss 4.53fF $ **FLOATING
C621 vdd.n663 vss 4.53fF $ **FLOATING
C622 vdd.n664 vss 4.42fF $ **FLOATING
C623 vdd.n665 vss 4.42fF $ **FLOATING
C624 vdd.n666 vss 4.42fF $ **FLOATING
C625 vdd.n667 vss 4.02fF $ **FLOATING
C626 vdd.n671 vss 32.58fF $ **FLOATING
C627 vdd.n674 vss 4.21fF $ **FLOATING
C628 vdd.n675 vss 4.42fF $ **FLOATING
C629 vdd.n676 vss 4.42fF $ **FLOATING
C630 vdd.n677 vss 4.42fF $ **FLOATING
C631 vdd.n678 vss 4.53fF $ **FLOATING
C632 vdd.n679 vss 4.53fF $ **FLOATING
C633 vdd.n680 vss 4.42fF $ **FLOATING
C634 vdd.n681 vss 4.42fF $ **FLOATING
C635 vdd.n682 vss 4.42fF $ **FLOATING
C636 vdd.n683 vss 4.02fF $ **FLOATING
C637 vdd.n685 vss 32.58fF $ **FLOATING
C638 vdd.n686 vss 4.21fF $ **FLOATING
C639 vdd.n687 vss 4.42fF $ **FLOATING
C640 vdd.n688 vss 4.42fF $ **FLOATING
C641 vdd.n689 vss 4.42fF $ **FLOATING
C642 vdd.n690 vss 4.53fF $ **FLOATING
C643 vdd.n691 vss 4.53fF $ **FLOATING
C644 vdd.n692 vss 4.42fF $ **FLOATING
C645 vdd.n693 vss 4.42fF $ **FLOATING
C646 vdd.n694 vss 4.42fF $ **FLOATING
C647 vdd.n695 vss 4.02fF $ **FLOATING
C648 vdd.n699 vss 32.58fF $ **FLOATING
C649 vdd.n702 vss 4.21fF $ **FLOATING
C650 vdd.n703 vss 4.42fF $ **FLOATING
C651 vdd.n704 vss 4.42fF $ **FLOATING
C652 vdd.n705 vss 4.42fF $ **FLOATING
C653 vdd.n706 vss 4.53fF $ **FLOATING
C654 vdd.n707 vss 4.53fF $ **FLOATING
C655 vdd.n708 vss 4.42fF $ **FLOATING
C656 vdd.n709 vss 4.42fF $ **FLOATING
C657 vdd.n710 vss 4.42fF $ **FLOATING
C658 vdd.n711 vss 4.02fF $ **FLOATING
C659 vdd.n713 vss 32.58fF $ **FLOATING
C660 vdd.n714 vss 4.21fF $ **FLOATING
C661 vdd.n715 vss 4.42fF $ **FLOATING
C662 vdd.n716 vss 4.42fF $ **FLOATING
C663 vdd.n717 vss 4.42fF $ **FLOATING
C664 vdd.n718 vss 4.53fF $ **FLOATING
C665 vdd.n719 vss 4.53fF $ **FLOATING
C666 vdd.n720 vss 4.42fF $ **FLOATING
C667 vdd.n721 vss 4.42fF $ **FLOATING
C668 vdd.n722 vss 4.42fF $ **FLOATING
C669 vdd.n723 vss 4.02fF $ **FLOATING
C670 vdd.n727 vss 32.58fF $ **FLOATING
C671 vdd.n730 vss 4.21fF $ **FLOATING
C672 vdd.n731 vss 4.42fF $ **FLOATING
C673 vdd.n732 vss 4.42fF $ **FLOATING
C674 vdd.n733 vss 4.42fF $ **FLOATING
C675 vdd.n734 vss 4.53fF $ **FLOATING
C676 vdd.n735 vss 4.53fF $ **FLOATING
C677 vdd.n736 vss 4.42fF $ **FLOATING
C678 vdd.n737 vss 4.42fF $ **FLOATING
C679 vdd.n738 vss 4.42fF $ **FLOATING
C680 vdd.n739 vss 4.02fF $ **FLOATING
C681 vdd.n741 vss 32.58fF $ **FLOATING
C682 vdd.n742 vss 4.21fF $ **FLOATING
C683 vdd.n743 vss 4.42fF $ **FLOATING
C684 vdd.n744 vss 4.42fF $ **FLOATING
C685 vdd.n745 vss 4.42fF $ **FLOATING
C686 vdd.n746 vss 4.53fF $ **FLOATING
C687 vdd.n747 vss 4.53fF $ **FLOATING
C688 vdd.n748 vss 4.42fF $ **FLOATING
C689 vdd.n749 vss 4.42fF $ **FLOATING
C690 vdd.n750 vss 4.42fF $ **FLOATING
C691 vdd.n751 vss 4.02fF $ **FLOATING
C692 vdd.n755 vss 32.58fF $ **FLOATING
C693 vdd.n758 vss 4.21fF $ **FLOATING
C694 vdd.n759 vss 4.42fF $ **FLOATING
C695 vdd.n760 vss 4.42fF $ **FLOATING
C696 vdd.n761 vss 4.42fF $ **FLOATING
C697 vdd.n762 vss 4.53fF $ **FLOATING
C698 vdd.n763 vss 4.53fF $ **FLOATING
C699 vdd.n764 vss 4.42fF $ **FLOATING
C700 vdd.n765 vss 4.42fF $ **FLOATING
C701 vdd.n766 vss 4.42fF $ **FLOATING
C702 vdd.n767 vss 4.02fF $ **FLOATING
C703 vdd.n769 vss 32.58fF $ **FLOATING
C704 vdd.n770 vss 4.21fF $ **FLOATING
C705 vdd.n771 vss 4.42fF $ **FLOATING
C706 vdd.n772 vss 4.42fF $ **FLOATING
C707 vdd.n773 vss 4.42fF $ **FLOATING
C708 vdd.n774 vss 4.53fF $ **FLOATING
C709 vdd.n775 vss 4.53fF $ **FLOATING
C710 vdd.n776 vss 4.42fF $ **FLOATING
C711 vdd.n777 vss 4.42fF $ **FLOATING
C712 vdd.n778 vss 4.42fF $ **FLOATING
C713 vdd.n779 vss 4.02fF $ **FLOATING
C714 vdd.n783 vss 32.58fF $ **FLOATING
C715 vdd.n786 vss 4.21fF $ **FLOATING
C716 vdd.n787 vss 4.42fF $ **FLOATING
C717 vdd.n788 vss 4.42fF $ **FLOATING
C718 vdd.n789 vss 4.42fF $ **FLOATING
C719 vdd.n790 vss 4.53fF $ **FLOATING
C720 vdd.n791 vss 4.53fF $ **FLOATING
C721 vdd.n792 vss 4.42fF $ **FLOATING
C722 vdd.n793 vss 4.42fF $ **FLOATING
C723 vdd.n794 vss 4.42fF $ **FLOATING
C724 vdd.n795 vss 4.02fF $ **FLOATING
C725 vdd.n797 vss 32.58fF $ **FLOATING
C726 vdd.n798 vss 4.21fF $ **FLOATING
C727 vdd.n799 vss 4.42fF $ **FLOATING
C728 vdd.n800 vss 4.42fF $ **FLOATING
C729 vdd.n801 vss 4.42fF $ **FLOATING
C730 vdd.n802 vss 4.53fF $ **FLOATING
C731 vdd.n803 vss 4.53fF $ **FLOATING
C732 vdd.n804 vss 4.42fF $ **FLOATING
C733 vdd.n805 vss 4.42fF $ **FLOATING
C734 vdd.n806 vss 4.42fF $ **FLOATING
C735 vdd.n807 vss 4.02fF $ **FLOATING
C736 vdd.n811 vss 32.58fF $ **FLOATING
C737 vdd.n814 vss 4.21fF $ **FLOATING
C738 vdd.n815 vss 4.42fF $ **FLOATING
C739 vdd.n816 vss 4.42fF $ **FLOATING
C740 vdd.n817 vss 4.42fF $ **FLOATING
C741 vdd.n818 vss 4.53fF $ **FLOATING
C742 vdd.n819 vss 4.53fF $ **FLOATING
C743 vdd.n820 vss 4.42fF $ **FLOATING
C744 vdd.n821 vss 4.42fF $ **FLOATING
C745 vdd.n822 vss 4.42fF $ **FLOATING
C746 vdd.n823 vss 4.02fF $ **FLOATING
C747 vdd.n825 vss 32.58fF $ **FLOATING
C748 vdd.n826 vss 4.21fF $ **FLOATING
C749 vdd.n827 vss 4.42fF $ **FLOATING
C750 vdd.n828 vss 4.42fF $ **FLOATING
C751 vdd.n829 vss 4.42fF $ **FLOATING
C752 vdd.n830 vss 4.53fF $ **FLOATING
C753 vdd.n831 vss 4.53fF $ **FLOATING
C754 vdd.n832 vss 4.42fF $ **FLOATING
C755 vdd.n833 vss 4.42fF $ **FLOATING
C756 vdd.n834 vss 4.42fF $ **FLOATING
C757 vdd.n835 vss 4.02fF $ **FLOATING
C758 vdd.n839 vss 32.58fF $ **FLOATING
C759 vdd.n842 vss 4.21fF $ **FLOATING
C760 vdd.n843 vss 4.42fF $ **FLOATING
C761 vdd.n844 vss 4.42fF $ **FLOATING
C762 vdd.n845 vss 4.42fF $ **FLOATING
C763 vdd.n846 vss 4.53fF $ **FLOATING
C764 vdd.n847 vss 4.53fF $ **FLOATING
C765 vdd.n848 vss 4.42fF $ **FLOATING
C766 vdd.n849 vss 4.42fF $ **FLOATING
C767 vdd.n850 vss 4.42fF $ **FLOATING
C768 vdd.n851 vss 4.02fF $ **FLOATING
C769 vdd.n853 vss 32.58fF $ **FLOATING
C770 vdd.n854 vss 4.21fF $ **FLOATING
C771 vdd.n855 vss 4.42fF $ **FLOATING
C772 vdd.n856 vss 4.42fF $ **FLOATING
C773 vdd.n857 vss 4.42fF $ **FLOATING
C774 vdd.n858 vss 4.53fF $ **FLOATING
C775 vdd.n859 vss 4.53fF $ **FLOATING
C776 vdd.n860 vss 4.42fF $ **FLOATING
C777 vdd.n861 vss 4.42fF $ **FLOATING
C778 vdd.n862 vss 4.42fF $ **FLOATING
C779 vdd.n863 vss 4.02fF $ **FLOATING
C780 vdd.n867 vss 32.58fF $ **FLOATING
C781 vdd.n870 vss 4.21fF $ **FLOATING
C782 vdd.n871 vss 4.42fF $ **FLOATING
C783 vdd.n872 vss 4.42fF $ **FLOATING
C784 vdd.n873 vss 4.42fF $ **FLOATING
C785 vdd.n874 vss 4.53fF $ **FLOATING
C786 vdd.n875 vss 4.53fF $ **FLOATING
C787 vdd.n876 vss 4.42fF $ **FLOATING
C788 vdd.n877 vss 4.42fF $ **FLOATING
C789 vdd.n878 vss 4.42fF $ **FLOATING
C790 vdd.n879 vss 4.02fF $ **FLOATING
C791 vdd.n881 vss 32.58fF $ **FLOATING
C792 vdd.n882 vss 4.21fF $ **FLOATING
C793 vdd.n883 vss 4.42fF $ **FLOATING
C794 vdd.n884 vss 4.42fF $ **FLOATING
C795 vdd.n885 vss 4.42fF $ **FLOATING
C796 vdd.n886 vss 4.53fF $ **FLOATING
C797 vdd.n887 vss 4.53fF $ **FLOATING
C798 vdd.n888 vss 4.42fF $ **FLOATING
C799 vdd.n889 vss 4.42fF $ **FLOATING
C800 vdd.n890 vss 4.42fF $ **FLOATING
C801 vdd.n891 vss 4.02fF $ **FLOATING
C802 vdd.n895 vss 32.58fF $ **FLOATING
C803 vdd.n898 vss 4.21fF $ **FLOATING
C804 vdd.n899 vss 4.42fF $ **FLOATING
C805 vdd.n900 vss 4.42fF $ **FLOATING
C806 vdd.n901 vss 4.42fF $ **FLOATING
C807 vdd.n902 vss 4.53fF $ **FLOATING
C808 vdd.n903 vss 4.53fF $ **FLOATING
C809 vdd.n904 vss 4.42fF $ **FLOATING
C810 vdd.n905 vss 4.42fF $ **FLOATING
C811 vdd.n906 vss 4.42fF $ **FLOATING
C812 vdd.n907 vss 4.02fF $ **FLOATING
C813 vdd.n909 vss 32.58fF $ **FLOATING
C814 vdd.n910 vss 4.21fF $ **FLOATING
C815 vdd.n911 vss 4.42fF $ **FLOATING
C816 vdd.n912 vss 4.42fF $ **FLOATING
C817 vdd.n913 vss 4.42fF $ **FLOATING
C818 vdd.n914 vss 4.53fF $ **FLOATING
C819 vdd.n915 vss 4.53fF $ **FLOATING
C820 vdd.n916 vss 4.42fF $ **FLOATING
C821 vdd.n917 vss 4.42fF $ **FLOATING
C822 vdd.n918 vss 4.42fF $ **FLOATING
C823 vdd.n919 vss 4.02fF $ **FLOATING
C824 vdd.n923 vss 32.58fF $ **FLOATING
C825 vdd.n926 vss 4.21fF $ **FLOATING
C826 vdd.n927 vss 4.42fF $ **FLOATING
C827 vdd.n928 vss 4.42fF $ **FLOATING
C828 vdd.n929 vss 4.42fF $ **FLOATING
C829 vdd.n930 vss 4.53fF $ **FLOATING
C830 vdd.n931 vss 4.53fF $ **FLOATING
C831 vdd.n932 vss 4.42fF $ **FLOATING
C832 vdd.n933 vss 4.42fF $ **FLOATING
C833 vdd.n934 vss 4.42fF $ **FLOATING
C834 vdd.n935 vss 4.02fF $ **FLOATING
C835 vdd.n937 vss 32.58fF $ **FLOATING
C836 vdd.n938 vss 4.21fF $ **FLOATING
C837 vdd.n939 vss 4.42fF $ **FLOATING
C838 vdd.n940 vss 4.42fF $ **FLOATING
C839 vdd.n941 vss 4.42fF $ **FLOATING
C840 vdd.n942 vss 4.53fF $ **FLOATING
C841 vdd.n943 vss 4.53fF $ **FLOATING
C842 vdd.n944 vss 4.42fF $ **FLOATING
C843 vdd.n945 vss 4.42fF $ **FLOATING
C844 vdd.n946 vss 4.42fF $ **FLOATING
C845 vdd.n947 vss 4.02fF $ **FLOATING
C846 vdd.n951 vss 32.58fF $ **FLOATING
C847 vdd.n954 vss 4.21fF $ **FLOATING
C848 vdd.n955 vss 4.42fF $ **FLOATING
C849 vdd.n956 vss 4.42fF $ **FLOATING
C850 vdd.n957 vss 4.42fF $ **FLOATING
C851 vdd.n958 vss 4.53fF $ **FLOATING
C852 vdd.n959 vss 4.53fF $ **FLOATING
C853 vdd.n960 vss 4.42fF $ **FLOATING
C854 vdd.n961 vss 4.42fF $ **FLOATING
C855 vdd.n962 vss 4.42fF $ **FLOATING
C856 vdd.n963 vss 4.02fF $ **FLOATING
C857 vdd.n965 vss 32.58fF $ **FLOATING
C858 vdd.n966 vss 4.21fF $ **FLOATING
C859 vdd.n967 vss 4.42fF $ **FLOATING
C860 vdd.n968 vss 4.42fF $ **FLOATING
C861 vdd.n969 vss 4.42fF $ **FLOATING
C862 vdd.n970 vss 4.53fF $ **FLOATING
C863 vdd.n971 vss 4.53fF $ **FLOATING
C864 vdd.n972 vss 4.42fF $ **FLOATING
C865 vdd.n973 vss 4.42fF $ **FLOATING
C866 vdd.n974 vss 4.42fF $ **FLOATING
C867 vdd.n975 vss 4.02fF $ **FLOATING
C868 vdd.n979 vss 32.58fF $ **FLOATING
C869 vdd.n982 vss 4.21fF $ **FLOATING
C870 vdd.n983 vss 4.42fF $ **FLOATING
C871 vdd.n984 vss 4.42fF $ **FLOATING
C872 vdd.n985 vss 4.42fF $ **FLOATING
C873 vdd.n986 vss 4.53fF $ **FLOATING
C874 vdd.n987 vss 4.53fF $ **FLOATING
C875 vdd.n988 vss 4.42fF $ **FLOATING
C876 vdd.n989 vss 4.42fF $ **FLOATING
C877 vdd.n990 vss 4.42fF $ **FLOATING
C878 vdd.n991 vss 4.02fF $ **FLOATING
C879 vdd.n993 vss 32.58fF $ **FLOATING
C880 vdd.n994 vss 4.21fF $ **FLOATING
C881 vdd.n995 vss 4.42fF $ **FLOATING
C882 vdd.n996 vss 4.42fF $ **FLOATING
C883 vdd.n997 vss 4.42fF $ **FLOATING
C884 vdd.n998 vss 4.53fF $ **FLOATING
C885 vdd.n999 vss 4.53fF $ **FLOATING
C886 vdd.n1000 vss 4.42fF $ **FLOATING
C887 vdd.n1001 vss 4.42fF $ **FLOATING
C888 vdd.n1002 vss 4.42fF $ **FLOATING
C889 vdd.n1003 vss 4.02fF $ **FLOATING
C890 vdd.n1007 vss 32.58fF $ **FLOATING
C891 vdd.n1010 vss 4.21fF $ **FLOATING
C892 vdd.n1011 vss 4.42fF $ **FLOATING
C893 vdd.n1012 vss 4.42fF $ **FLOATING
C894 vdd.n1013 vss 4.42fF $ **FLOATING
C895 vdd.n1014 vss 4.53fF $ **FLOATING
C896 vdd.n1015 vss 4.53fF $ **FLOATING
C897 vdd.n1016 vss 4.42fF $ **FLOATING
C898 vdd.n1017 vss 4.42fF $ **FLOATING
C899 vdd.n1018 vss 4.42fF $ **FLOATING
C900 vdd.n1019 vss 4.02fF $ **FLOATING
C901 vdd.n1021 vss 32.58fF $ **FLOATING
C902 vdd.n1022 vss 4.21fF $ **FLOATING
C903 vdd.n1023 vss 4.42fF $ **FLOATING
C904 vdd.n1024 vss 4.42fF $ **FLOATING
C905 vdd.n1025 vss 4.42fF $ **FLOATING
C906 vdd.n1026 vss 4.53fF $ **FLOATING
C907 vdd.n1027 vss 4.53fF $ **FLOATING
C908 vdd.n1028 vss 4.42fF $ **FLOATING
C909 vdd.n1029 vss 4.42fF $ **FLOATING
C910 vdd.n1030 vss 4.42fF $ **FLOATING
C911 vdd.n1031 vss 4.02fF $ **FLOATING
C912 vdd.n1035 vss 32.58fF $ **FLOATING
C913 vdd.n1038 vss 4.21fF $ **FLOATING
C914 vdd.n1039 vss 4.42fF $ **FLOATING
C915 vdd.n1040 vss 4.42fF $ **FLOATING
C916 vdd.n1041 vss 4.42fF $ **FLOATING
C917 vdd.n1042 vss 4.53fF $ **FLOATING
C918 vdd.n1043 vss 4.53fF $ **FLOATING
C919 vdd.n1044 vss 4.42fF $ **FLOATING
C920 vdd.n1045 vss 4.42fF $ **FLOATING
C921 vdd.n1046 vss 4.42fF $ **FLOATING
C922 vdd.n1047 vss 4.02fF $ **FLOATING
C923 vdd.n1049 vss 32.58fF $ **FLOATING
C924 vdd.n1050 vss 4.21fF $ **FLOATING
C925 vdd.n1051 vss 4.42fF $ **FLOATING
C926 vdd.n1052 vss 4.42fF $ **FLOATING
C927 vdd.n1053 vss 4.42fF $ **FLOATING
C928 vdd.n1054 vss 4.53fF $ **FLOATING
C929 vdd.n1055 vss 4.53fF $ **FLOATING
C930 vdd.n1056 vss 4.42fF $ **FLOATING
C931 vdd.n1057 vss 4.42fF $ **FLOATING
C932 vdd.n1058 vss 4.42fF $ **FLOATING
C933 vdd.n1059 vss 4.02fF $ **FLOATING
C934 vdd.n1063 vss 29.96fF $ **FLOATING
C935 out_p.n0 vss 3.87fF $ **FLOATING
C936 out_p.n1 vss 4.05fF $ **FLOATING
C937 out_p.n2 vss 4.05fF $ **FLOATING
C938 out_p.n3 vss 4.05fF $ **FLOATING
C939 out_p.n4 vss 4.15fF $ **FLOATING
C940 out_p.n5 vss 4.15fF $ **FLOATING
C941 out_p.n6 vss 4.05fF $ **FLOATING
C942 out_p.n7 vss 4.05fF $ **FLOATING
C943 out_p.n8 vss 4.05fF $ **FLOATING
C944 out_p.n9 vss 3.80fF $ **FLOATING
C945 out_p.n10 vss 3.85fF $ **FLOATING
C946 out_p.n11 vss 3.81fF $ **FLOATING
C947 out_p.n12 vss 3.85fF $ **FLOATING
C948 out_p.n13 vss 3.81fF $ **FLOATING
C949 out_p.n14 vss 3.85fF $ **FLOATING
C950 out_p.n15 vss 3.81fF $ **FLOATING
C951 out_p.n16 vss 3.85fF $ **FLOATING
C952 out_p.n17 vss 3.81fF $ **FLOATING
C953 out_p.n18 vss 3.85fF $ **FLOATING
C954 out_p.n19 vss 3.81fF $ **FLOATING
C955 out_p.n20 vss 3.85fF $ **FLOATING
C956 out_p.n21 vss 3.81fF $ **FLOATING
C957 out_p.n22 vss 3.85fF $ **FLOATING
C958 out_p.n23 vss 3.81fF $ **FLOATING
C959 out_p.n24 vss 3.85fF $ **FLOATING
C960 out_p.n25 vss 3.81fF $ **FLOATING
C961 out_p.n26 vss 3.85fF $ **FLOATING
C962 out_p.n27 vss 3.81fF $ **FLOATING
C963 out_p.n28 vss 3.85fF $ **FLOATING
C964 out_p.n29 vss 3.81fF $ **FLOATING
C965 out_p.n30 vss 3.85fF $ **FLOATING
C966 out_p.n31 vss 3.81fF $ **FLOATING
C967 out_p.n32 vss 3.85fF $ **FLOATING
C968 out_p.n33 vss 3.81fF $ **FLOATING
C969 out_p.n34 vss 3.85fF $ **FLOATING
C970 out_p.n35 vss 3.81fF $ **FLOATING
C971 out_p.n36 vss 3.87fF $ **FLOATING
C972 out_p.n37 vss 4.05fF $ **FLOATING
C973 out_p.n38 vss 4.05fF $ **FLOATING
C974 out_p.n39 vss 4.05fF $ **FLOATING
C975 out_p.n40 vss 4.15fF $ **FLOATING
C976 out_p.n41 vss 4.15fF $ **FLOATING
C977 out_p.n42 vss 4.05fF $ **FLOATING
C978 out_p.n43 vss 4.05fF $ **FLOATING
C979 out_p.n44 vss 4.05fF $ **FLOATING
C980 out_p.n45 vss 3.80fF $ **FLOATING
C981 out_p.n46 vss 33.39fF $ **FLOATING
C982 out_p.n47 vss 3.87fF $ **FLOATING
C983 out_p.n48 vss 4.05fF $ **FLOATING
C984 out_p.n49 vss 4.05fF $ **FLOATING
C985 out_p.n50 vss 4.05fF $ **FLOATING
C986 out_p.n51 vss 4.15fF $ **FLOATING
C987 out_p.n52 vss 4.15fF $ **FLOATING
C988 out_p.n53 vss 4.05fF $ **FLOATING
C989 out_p.n54 vss 4.05fF $ **FLOATING
C990 out_p.n55 vss 4.05fF $ **FLOATING
C991 out_p.n56 vss 3.80fF $ **FLOATING
C992 out_p.n57 vss 30.23fF $ **FLOATING
C993 out_p.n58 vss 3.87fF $ **FLOATING
C994 out_p.n59 vss 4.05fF $ **FLOATING
C995 out_p.n60 vss 4.05fF $ **FLOATING
C996 out_p.n61 vss 4.05fF $ **FLOATING
C997 out_p.n62 vss 4.15fF $ **FLOATING
C998 out_p.n63 vss 4.15fF $ **FLOATING
C999 out_p.n64 vss 4.05fF $ **FLOATING
C1000 out_p.n65 vss 4.05fF $ **FLOATING
C1001 out_p.n66 vss 4.05fF $ **FLOATING
C1002 out_p.n67 vss 3.80fF $ **FLOATING
C1003 out_p.n68 vss 30.23fF $ **FLOATING
C1004 out_p.n69 vss 3.87fF $ **FLOATING
C1005 out_p.n70 vss 4.05fF $ **FLOATING
C1006 out_p.n71 vss 4.05fF $ **FLOATING
C1007 out_p.n72 vss 4.05fF $ **FLOATING
C1008 out_p.n73 vss 4.15fF $ **FLOATING
C1009 out_p.n74 vss 4.15fF $ **FLOATING
C1010 out_p.n75 vss 4.05fF $ **FLOATING
C1011 out_p.n76 vss 4.05fF $ **FLOATING
C1012 out_p.n77 vss 4.05fF $ **FLOATING
C1013 out_p.n78 vss 3.80fF $ **FLOATING
C1014 out_p.n79 vss 30.23fF $ **FLOATING
C1015 out_p.n80 vss 3.87fF $ **FLOATING
C1016 out_p.n81 vss 4.05fF $ **FLOATING
C1017 out_p.n82 vss 4.05fF $ **FLOATING
C1018 out_p.n83 vss 4.05fF $ **FLOATING
C1019 out_p.n84 vss 4.15fF $ **FLOATING
C1020 out_p.n85 vss 4.15fF $ **FLOATING
C1021 out_p.n86 vss 4.05fF $ **FLOATING
C1022 out_p.n87 vss 4.05fF $ **FLOATING
C1023 out_p.n88 vss 4.05fF $ **FLOATING
C1024 out_p.n89 vss 3.80fF $ **FLOATING
C1025 out_p.n90 vss 30.23fF $ **FLOATING
C1026 out_p.n91 vss 3.87fF $ **FLOATING
C1027 out_p.n92 vss 4.05fF $ **FLOATING
C1028 out_p.n93 vss 4.05fF $ **FLOATING
C1029 out_p.n94 vss 4.05fF $ **FLOATING
C1030 out_p.n95 vss 4.15fF $ **FLOATING
C1031 out_p.n96 vss 4.15fF $ **FLOATING
C1032 out_p.n97 vss 4.05fF $ **FLOATING
C1033 out_p.n98 vss 4.05fF $ **FLOATING
C1034 out_p.n99 vss 4.05fF $ **FLOATING
C1035 out_p.n100 vss 3.80fF $ **FLOATING
C1036 out_p.n101 vss 30.23fF $ **FLOATING
C1037 out_p.n102 vss 3.87fF $ **FLOATING
C1038 out_p.n103 vss 4.05fF $ **FLOATING
C1039 out_p.n104 vss 4.05fF $ **FLOATING
C1040 out_p.n105 vss 4.05fF $ **FLOATING
C1041 out_p.n106 vss 4.15fF $ **FLOATING
C1042 out_p.n107 vss 4.15fF $ **FLOATING
C1043 out_p.n108 vss 4.05fF $ **FLOATING
C1044 out_p.n109 vss 4.05fF $ **FLOATING
C1045 out_p.n110 vss 4.05fF $ **FLOATING
C1046 out_p.n111 vss 3.80fF $ **FLOATING
C1047 out_p.n112 vss 30.23fF $ **FLOATING
C1048 out_p.n113 vss 3.87fF $ **FLOATING
C1049 out_p.n114 vss 4.05fF $ **FLOATING
C1050 out_p.n115 vss 4.05fF $ **FLOATING
C1051 out_p.n116 vss 4.05fF $ **FLOATING
C1052 out_p.n117 vss 4.15fF $ **FLOATING
C1053 out_p.n118 vss 4.15fF $ **FLOATING
C1054 out_p.n119 vss 4.05fF $ **FLOATING
C1055 out_p.n120 vss 4.05fF $ **FLOATING
C1056 out_p.n121 vss 4.05fF $ **FLOATING
C1057 out_p.n122 vss 3.80fF $ **FLOATING
C1058 out_p.n123 vss 30.23fF $ **FLOATING
C1059 out_p.n124 vss 3.87fF $ **FLOATING
C1060 out_p.n125 vss 4.05fF $ **FLOATING
C1061 out_p.n126 vss 4.05fF $ **FLOATING
C1062 out_p.n127 vss 4.05fF $ **FLOATING
C1063 out_p.n128 vss 4.15fF $ **FLOATING
C1064 out_p.n129 vss 4.15fF $ **FLOATING
C1065 out_p.n130 vss 4.05fF $ **FLOATING
C1066 out_p.n131 vss 4.05fF $ **FLOATING
C1067 out_p.n132 vss 4.05fF $ **FLOATING
C1068 out_p.n133 vss 3.80fF $ **FLOATING
C1069 out_p.n134 vss 30.23fF $ **FLOATING
C1070 out_p.n135 vss 3.87fF $ **FLOATING
C1071 out_p.n136 vss 4.05fF $ **FLOATING
C1072 out_p.n137 vss 4.05fF $ **FLOATING
C1073 out_p.n138 vss 4.05fF $ **FLOATING
C1074 out_p.n139 vss 4.15fF $ **FLOATING
C1075 out_p.n140 vss 4.15fF $ **FLOATING
C1076 out_p.n141 vss 4.05fF $ **FLOATING
C1077 out_p.n142 vss 4.05fF $ **FLOATING
C1078 out_p.n143 vss 4.05fF $ **FLOATING
C1079 out_p.n144 vss 3.80fF $ **FLOATING
C1080 out_p.n145 vss 30.23fF $ **FLOATING
C1081 out_p.n146 vss 3.87fF $ **FLOATING
C1082 out_p.n147 vss 4.05fF $ **FLOATING
C1083 out_p.n148 vss 4.05fF $ **FLOATING
C1084 out_p.n149 vss 4.05fF $ **FLOATING
C1085 out_p.n150 vss 4.15fF $ **FLOATING
C1086 out_p.n151 vss 4.15fF $ **FLOATING
C1087 out_p.n152 vss 4.05fF $ **FLOATING
C1088 out_p.n153 vss 4.05fF $ **FLOATING
C1089 out_p.n154 vss 4.05fF $ **FLOATING
C1090 out_p.n155 vss 3.80fF $ **FLOATING
C1091 out_p.n156 vss 30.23fF $ **FLOATING
C1092 out_p.n157 vss 3.87fF $ **FLOATING
C1093 out_p.n158 vss 4.05fF $ **FLOATING
C1094 out_p.n159 vss 4.05fF $ **FLOATING
C1095 out_p.n160 vss 4.05fF $ **FLOATING
C1096 out_p.n161 vss 4.15fF $ **FLOATING
C1097 out_p.n162 vss 4.15fF $ **FLOATING
C1098 out_p.n163 vss 4.05fF $ **FLOATING
C1099 out_p.n164 vss 4.05fF $ **FLOATING
C1100 out_p.n165 vss 4.05fF $ **FLOATING
C1101 out_p.n166 vss 3.80fF $ **FLOATING
C1102 out_p.n167 vss 30.23fF $ **FLOATING
C1103 out_p.n168 vss 3.87fF $ **FLOATING
C1104 out_p.n169 vss 4.05fF $ **FLOATING
C1105 out_p.n170 vss 4.05fF $ **FLOATING
C1106 out_p.n171 vss 4.05fF $ **FLOATING
C1107 out_p.n172 vss 4.15fF $ **FLOATING
C1108 out_p.n173 vss 4.15fF $ **FLOATING
C1109 out_p.n174 vss 4.05fF $ **FLOATING
C1110 out_p.n175 vss 4.05fF $ **FLOATING
C1111 out_p.n176 vss 4.05fF $ **FLOATING
C1112 out_p.n177 vss 3.80fF $ **FLOATING
C1113 out_p.n178 vss 30.23fF $ **FLOATING
C1114 out_p.n179 vss 3.85fF $ **FLOATING
C1115 out_p.n180 vss 3.81fF $ **FLOATING
C1116 out_p.n181 vss 3.85fF $ **FLOATING
C1117 out_p.n182 vss 3.81fF $ **FLOATING
C1118 out_p.n183 vss 3.87fF $ **FLOATING
C1119 out_p.n184 vss 4.05fF $ **FLOATING
C1120 out_p.n185 vss 4.05fF $ **FLOATING
C1121 out_p.n186 vss 4.05fF $ **FLOATING
C1122 out_p.n187 vss 4.15fF $ **FLOATING
C1123 out_p.n188 vss 4.15fF $ **FLOATING
C1124 out_p.n189 vss 4.05fF $ **FLOATING
C1125 out_p.n190 vss 4.05fF $ **FLOATING
C1126 out_p.n191 vss 4.05fF $ **FLOATING
C1127 out_p.n192 vss 3.80fF $ **FLOATING
C1128 out_p.n193 vss 3.85fF $ **FLOATING
C1129 out_p.n194 vss 3.81fF $ **FLOATING
C1130 out_p.n195 vss 3.87fF $ **FLOATING
C1131 out_p.n196 vss 4.05fF $ **FLOATING
C1132 out_p.n197 vss 4.05fF $ **FLOATING
C1133 out_p.n198 vss 4.05fF $ **FLOATING
C1134 out_p.n199 vss 4.15fF $ **FLOATING
C1135 out_p.n200 vss 4.15fF $ **FLOATING
C1136 out_p.n201 vss 4.05fF $ **FLOATING
C1137 out_p.n202 vss 4.05fF $ **FLOATING
C1138 out_p.n203 vss 4.05fF $ **FLOATING
C1139 out_p.n204 vss 3.80fF $ **FLOATING
C1140 out_p.n205 vss 3.85fF $ **FLOATING
C1141 out_p.n206 vss 3.81fF $ **FLOATING
C1142 out_p.n207 vss 3.87fF $ **FLOATING
C1143 out_p.n208 vss 4.05fF $ **FLOATING
C1144 out_p.n209 vss 4.05fF $ **FLOATING
C1145 out_p.n210 vss 4.05fF $ **FLOATING
C1146 out_p.n211 vss 4.15fF $ **FLOATING
C1147 out_p.n212 vss 4.15fF $ **FLOATING
C1148 out_p.n213 vss 4.05fF $ **FLOATING
C1149 out_p.n214 vss 4.05fF $ **FLOATING
C1150 out_p.n215 vss 4.05fF $ **FLOATING
C1151 out_p.n216 vss 3.80fF $ **FLOATING
C1152 out_p.n217 vss 3.85fF $ **FLOATING
C1153 out_p.n218 vss 3.81fF $ **FLOATING
C1154 out_p.n219 vss 3.87fF $ **FLOATING
C1155 out_p.n220 vss 4.05fF $ **FLOATING
C1156 out_p.n221 vss 4.05fF $ **FLOATING
C1157 out_p.n222 vss 4.05fF $ **FLOATING
C1158 out_p.n223 vss 4.15fF $ **FLOATING
C1159 out_p.n224 vss 4.15fF $ **FLOATING
C1160 out_p.n225 vss 4.05fF $ **FLOATING
C1161 out_p.n226 vss 4.05fF $ **FLOATING
C1162 out_p.n227 vss 4.05fF $ **FLOATING
C1163 out_p.n228 vss 3.80fF $ **FLOATING
C1164 out_p.n229 vss 3.85fF $ **FLOATING
C1165 out_p.n230 vss 3.81fF $ **FLOATING
C1166 out_p.n231 vss 3.87fF $ **FLOATING
C1167 out_p.n232 vss 4.05fF $ **FLOATING
C1168 out_p.n233 vss 4.05fF $ **FLOATING
C1169 out_p.n234 vss 4.05fF $ **FLOATING
C1170 out_p.n235 vss 4.15fF $ **FLOATING
C1171 out_p.n236 vss 4.15fF $ **FLOATING
C1172 out_p.n237 vss 4.05fF $ **FLOATING
C1173 out_p.n238 vss 4.05fF $ **FLOATING
C1174 out_p.n239 vss 4.05fF $ **FLOATING
C1175 out_p.n240 vss 3.80fF $ **FLOATING
C1176 out_p.n241 vss 3.85fF $ **FLOATING
C1177 out_p.n242 vss 3.81fF $ **FLOATING
C1178 out_p.n243 vss 3.87fF $ **FLOATING
C1179 out_p.n244 vss 4.05fF $ **FLOATING
C1180 out_p.n245 vss 4.05fF $ **FLOATING
C1181 out_p.n246 vss 4.05fF $ **FLOATING
C1182 out_p.n247 vss 4.15fF $ **FLOATING
C1183 out_p.n248 vss 4.15fF $ **FLOATING
C1184 out_p.n249 vss 4.05fF $ **FLOATING
C1185 out_p.n250 vss 4.05fF $ **FLOATING
C1186 out_p.n251 vss 4.05fF $ **FLOATING
C1187 out_p.n252 vss 3.80fF $ **FLOATING
C1188 out_p.n253 vss 3.85fF $ **FLOATING
C1189 out_p.n254 vss 3.81fF $ **FLOATING
C1190 out_p.n255 vss 3.87fF $ **FLOATING
C1191 out_p.n256 vss 4.05fF $ **FLOATING
C1192 out_p.n257 vss 4.05fF $ **FLOATING
C1193 out_p.n258 vss 4.05fF $ **FLOATING
C1194 out_p.n259 vss 4.15fF $ **FLOATING
C1195 out_p.n260 vss 4.15fF $ **FLOATING
C1196 out_p.n261 vss 4.05fF $ **FLOATING
C1197 out_p.n262 vss 4.05fF $ **FLOATING
C1198 out_p.n263 vss 4.05fF $ **FLOATING
C1199 out_p.n264 vss 3.80fF $ **FLOATING
C1200 out_p.n265 vss 3.85fF $ **FLOATING
C1201 out_p.n266 vss 3.81fF $ **FLOATING
C1202 out_p.n267 vss 3.87fF $ **FLOATING
C1203 out_p.n268 vss 4.05fF $ **FLOATING
C1204 out_p.n269 vss 4.05fF $ **FLOATING
C1205 out_p.n270 vss 4.05fF $ **FLOATING
C1206 out_p.n271 vss 4.15fF $ **FLOATING
C1207 out_p.n272 vss 4.15fF $ **FLOATING
C1208 out_p.n273 vss 4.05fF $ **FLOATING
C1209 out_p.n274 vss 4.05fF $ **FLOATING
C1210 out_p.n275 vss 4.05fF $ **FLOATING
C1211 out_p.n276 vss 3.80fF $ **FLOATING
C1212 out_p.n277 vss 3.85fF $ **FLOATING
C1213 out_p.n278 vss 3.81fF $ **FLOATING
C1214 out_p.n279 vss 3.87fF $ **FLOATING
C1215 out_p.n280 vss 4.05fF $ **FLOATING
C1216 out_p.n281 vss 4.05fF $ **FLOATING
C1217 out_p.n282 vss 4.05fF $ **FLOATING
C1218 out_p.n283 vss 4.15fF $ **FLOATING
C1219 out_p.n284 vss 4.15fF $ **FLOATING
C1220 out_p.n285 vss 4.05fF $ **FLOATING
C1221 out_p.n286 vss 4.05fF $ **FLOATING
C1222 out_p.n287 vss 4.05fF $ **FLOATING
C1223 out_p.n288 vss 3.80fF $ **FLOATING
C1224 out_p.n289 vss 3.85fF $ **FLOATING
C1225 out_p.n290 vss 3.81fF $ **FLOATING
C1226 out_p.n291 vss 3.87fF $ **FLOATING
C1227 out_p.n292 vss 4.05fF $ **FLOATING
C1228 out_p.n293 vss 4.05fF $ **FLOATING
C1229 out_p.n294 vss 4.05fF $ **FLOATING
C1230 out_p.n295 vss 4.15fF $ **FLOATING
C1231 out_p.n296 vss 4.15fF $ **FLOATING
C1232 out_p.n297 vss 4.05fF $ **FLOATING
C1233 out_p.n298 vss 4.05fF $ **FLOATING
C1234 out_p.n299 vss 4.05fF $ **FLOATING
C1235 out_p.n300 vss 3.80fF $ **FLOATING
C1236 out_p.n301 vss 3.85fF $ **FLOATING
C1237 out_p.n302 vss 3.81fF $ **FLOATING
C1238 out_p.n303 vss 3.87fF $ **FLOATING
C1239 out_p.n304 vss 4.05fF $ **FLOATING
C1240 out_p.n305 vss 4.05fF $ **FLOATING
C1241 out_p.n306 vss 4.05fF $ **FLOATING
C1242 out_p.n307 vss 4.15fF $ **FLOATING
C1243 out_p.n308 vss 4.15fF $ **FLOATING
C1244 out_p.n309 vss 4.05fF $ **FLOATING
C1245 out_p.n310 vss 4.05fF $ **FLOATING
C1246 out_p.n311 vss 4.05fF $ **FLOATING
C1247 out_p.n312 vss 3.80fF $ **FLOATING
C1248 out_p.n313 vss 3.85fF $ **FLOATING
C1249 out_p.n314 vss 3.81fF $ **FLOATING
C1250 out_p.n315 vss 3.87fF $ **FLOATING
C1251 out_p.n316 vss 4.05fF $ **FLOATING
C1252 out_p.n317 vss 4.05fF $ **FLOATING
C1253 out_p.n318 vss 4.05fF $ **FLOATING
C1254 out_p.n319 vss 4.15fF $ **FLOATING
C1255 out_p.n320 vss 4.15fF $ **FLOATING
C1256 out_p.n321 vss 4.05fF $ **FLOATING
C1257 out_p.n322 vss 4.05fF $ **FLOATING
C1258 out_p.n323 vss 4.05fF $ **FLOATING
C1259 out_p.n324 vss 3.80fF $ **FLOATING
C1260 out_p.n325 vss 3.85fF $ **FLOATING
C1261 out_p.n326 vss 3.81fF $ **FLOATING
C1262 out_p.n327 vss 3.87fF $ **FLOATING
C1263 out_p.n328 vss 4.05fF $ **FLOATING
C1264 out_p.n329 vss 4.05fF $ **FLOATING
C1265 out_p.n330 vss 4.05fF $ **FLOATING
C1266 out_p.n331 vss 4.15fF $ **FLOATING
C1267 out_p.n332 vss 4.15fF $ **FLOATING
C1268 out_p.n333 vss 4.05fF $ **FLOATING
C1269 out_p.n334 vss 4.05fF $ **FLOATING
C1270 out_p.n335 vss 4.05fF $ **FLOATING
C1271 out_p.n336 vss 3.80fF $ **FLOATING
C1272 out_p.n337 vss 3.85fF $ **FLOATING
C1273 out_p.n338 vss 3.81fF $ **FLOATING
C1274 out_p.n339 vss 3.87fF $ **FLOATING
C1275 out_p.n340 vss 4.05fF $ **FLOATING
C1276 out_p.n341 vss 4.05fF $ **FLOATING
C1277 out_p.n342 vss 4.05fF $ **FLOATING
C1278 out_p.n343 vss 4.15fF $ **FLOATING
C1279 out_p.n344 vss 4.15fF $ **FLOATING
C1280 out_p.n345 vss 4.05fF $ **FLOATING
C1281 out_p.n346 vss 4.05fF $ **FLOATING
C1282 out_p.n347 vss 4.05fF $ **FLOATING
C1283 out_p.n348 vss 3.80fF $ **FLOATING
C1284 out_p.n349 vss 3.85fF $ **FLOATING
C1285 out_p.n350 vss 3.81fF $ **FLOATING
C1286 out_p.n351 vss 3.87fF $ **FLOATING
C1287 out_p.n352 vss 4.05fF $ **FLOATING
C1288 out_p.n353 vss 4.05fF $ **FLOATING
C1289 out_p.n354 vss 4.05fF $ **FLOATING
C1290 out_p.n355 vss 4.15fF $ **FLOATING
C1291 out_p.n356 vss 4.15fF $ **FLOATING
C1292 out_p.n357 vss 4.05fF $ **FLOATING
C1293 out_p.n358 vss 4.05fF $ **FLOATING
C1294 out_p.n359 vss 4.05fF $ **FLOATING
C1295 out_p.n360 vss 3.80fF $ **FLOATING
C1296 out_p.n361 vss 3.85fF $ **FLOATING
C1297 out_p.n362 vss 3.81fF $ **FLOATING
C1298 out_p.n363 vss 3.87fF $ **FLOATING
C1299 out_p.n364 vss 4.05fF $ **FLOATING
C1300 out_p.n365 vss 4.05fF $ **FLOATING
C1301 out_p.n366 vss 4.05fF $ **FLOATING
C1302 out_p.n367 vss 4.15fF $ **FLOATING
C1303 out_p.n368 vss 4.15fF $ **FLOATING
C1304 out_p.n369 vss 4.05fF $ **FLOATING
C1305 out_p.n370 vss 4.05fF $ **FLOATING
C1306 out_p.n371 vss 4.05fF $ **FLOATING
C1307 out_p.n372 vss 3.80fF $ **FLOATING
C1308 out_p.n373 vss 3.85fF $ **FLOATING
C1309 out_p.n374 vss 3.81fF $ **FLOATING
C1310 out_p.n375 vss 3.87fF $ **FLOATING
C1311 out_p.n376 vss 4.05fF $ **FLOATING
C1312 out_p.n377 vss 4.05fF $ **FLOATING
C1313 out_p.n378 vss 4.05fF $ **FLOATING
C1314 out_p.n379 vss 4.15fF $ **FLOATING
C1315 out_p.n380 vss 4.15fF $ **FLOATING
C1316 out_p.n381 vss 4.05fF $ **FLOATING
C1317 out_p.n382 vss 4.05fF $ **FLOATING
C1318 out_p.n383 vss 4.05fF $ **FLOATING
C1319 out_p.n384 vss 3.80fF $ **FLOATING
C1320 out_p.n385 vss 3.85fF $ **FLOATING
C1321 out_p.n386 vss 3.81fF $ **FLOATING
C1322 out_p.n387 vss 3.87fF $ **FLOATING
C1323 out_p.n388 vss 4.05fF $ **FLOATING
C1324 out_p.n389 vss 4.05fF $ **FLOATING
C1325 out_p.n390 vss 4.05fF $ **FLOATING
C1326 out_p.n391 vss 4.15fF $ **FLOATING
C1327 out_p.n392 vss 4.15fF $ **FLOATING
C1328 out_p.n393 vss 4.05fF $ **FLOATING
C1329 out_p.n394 vss 4.05fF $ **FLOATING
C1330 out_p.n395 vss 4.05fF $ **FLOATING
C1331 out_p.n396 vss 3.80fF $ **FLOATING
C1332 out_p.n397 vss 3.85fF $ **FLOATING
C1333 out_p.n398 vss 3.81fF $ **FLOATING
C1334 out_p.n399 vss 3.87fF $ **FLOATING
C1335 out_p.n400 vss 4.05fF $ **FLOATING
C1336 out_p.n401 vss 4.05fF $ **FLOATING
C1337 out_p.n402 vss 4.05fF $ **FLOATING
C1338 out_p.n403 vss 4.15fF $ **FLOATING
C1339 out_p.n404 vss 4.15fF $ **FLOATING
C1340 out_p.n405 vss 4.05fF $ **FLOATING
C1341 out_p.n406 vss 4.05fF $ **FLOATING
C1342 out_p.n407 vss 4.05fF $ **FLOATING
C1343 out_p.n408 vss 3.80fF $ **FLOATING
C1344 out_p.n409 vss 3.85fF $ **FLOATING
C1345 out_p.n410 vss 3.81fF $ **FLOATING
C1346 out_p.n411 vss 3.87fF $ **FLOATING
C1347 out_p.n412 vss 4.05fF $ **FLOATING
C1348 out_p.n413 vss 4.05fF $ **FLOATING
C1349 out_p.n414 vss 4.05fF $ **FLOATING
C1350 out_p.n415 vss 4.15fF $ **FLOATING
C1351 out_p.n416 vss 4.15fF $ **FLOATING
C1352 out_p.n417 vss 4.05fF $ **FLOATING
C1353 out_p.n418 vss 4.05fF $ **FLOATING
C1354 out_p.n419 vss 4.05fF $ **FLOATING
C1355 out_p.n420 vss 3.80fF $ **FLOATING
C1356 out_p.n421 vss 3.85fF $ **FLOATING
C1357 out_p.n422 vss 3.81fF $ **FLOATING
C1358 out_p.n423 vss 3.87fF $ **FLOATING
C1359 out_p.n424 vss 4.05fF $ **FLOATING
C1360 out_p.n425 vss 4.05fF $ **FLOATING
C1361 out_p.n426 vss 4.05fF $ **FLOATING
C1362 out_p.n427 vss 4.15fF $ **FLOATING
C1363 out_p.n428 vss 4.15fF $ **FLOATING
C1364 out_p.n429 vss 4.05fF $ **FLOATING
C1365 out_p.n430 vss 4.05fF $ **FLOATING
C1366 out_p.n431 vss 4.05fF $ **FLOATING
C1367 out_p.n432 vss 3.80fF $ **FLOATING
C1368 out_p.n433 vss 3.85fF $ **FLOATING
C1369 out_p.n434 vss 3.81fF $ **FLOATING
C1370 out_p.n435 vss 3.87fF $ **FLOATING
C1371 out_p.n436 vss 4.05fF $ **FLOATING
C1372 out_p.n437 vss 4.05fF $ **FLOATING
C1373 out_p.n438 vss 4.05fF $ **FLOATING
C1374 out_p.n439 vss 4.15fF $ **FLOATING
C1375 out_p.n440 vss 4.15fF $ **FLOATING
C1376 out_p.n441 vss 4.05fF $ **FLOATING
C1377 out_p.n442 vss 4.05fF $ **FLOATING
C1378 out_p.n443 vss 4.05fF $ **FLOATING
C1379 out_p.n444 vss 3.80fF $ **FLOATING
C1380 out_p.n445 vss 3.85fF $ **FLOATING
C1381 out_p.n446 vss 3.81fF $ **FLOATING
C1382 out_p.n447 vss 3.87fF $ **FLOATING
C1383 out_p.n448 vss 4.05fF $ **FLOATING
C1384 out_p.n449 vss 4.05fF $ **FLOATING
C1385 out_p.n450 vss 4.05fF $ **FLOATING
C1386 out_p.n451 vss 4.15fF $ **FLOATING
C1387 out_p.n452 vss 4.15fF $ **FLOATING
C1388 out_p.n453 vss 4.05fF $ **FLOATING
C1389 out_p.n454 vss 4.05fF $ **FLOATING
C1390 out_p.n455 vss 4.05fF $ **FLOATING
C1391 out_p.n456 vss 3.80fF $ **FLOATING
C1392 out_p.n457 vss 3.85fF $ **FLOATING
C1393 out_p.n458 vss 3.81fF $ **FLOATING
C1394 out_p.n459 vss 3.87fF $ **FLOATING
C1395 out_p.n460 vss 4.05fF $ **FLOATING
C1396 out_p.n461 vss 4.05fF $ **FLOATING
C1397 out_p.n462 vss 4.05fF $ **FLOATING
C1398 out_p.n463 vss 4.15fF $ **FLOATING
C1399 out_p.n464 vss 4.15fF $ **FLOATING
C1400 out_p.n465 vss 4.05fF $ **FLOATING
C1401 out_p.n466 vss 4.05fF $ **FLOATING
C1402 out_p.n467 vss 4.05fF $ **FLOATING
C1403 out_p.n468 vss 3.80fF $ **FLOATING
C1404 out_p.n469 vss 3.85fF $ **FLOATING
C1405 out_p.n470 vss 3.81fF $ **FLOATING
C1406 out_p.n471 vss 3.87fF $ **FLOATING
C1407 out_p.n472 vss 4.05fF $ **FLOATING
C1408 out_p.n473 vss 4.05fF $ **FLOATING
C1409 out_p.n474 vss 4.05fF $ **FLOATING
C1410 out_p.n475 vss 4.15fF $ **FLOATING
C1411 out_p.n476 vss 4.15fF $ **FLOATING
C1412 out_p.n477 vss 4.05fF $ **FLOATING
C1413 out_p.n478 vss 4.05fF $ **FLOATING
C1414 out_p.n479 vss 4.05fF $ **FLOATING
C1415 out_p.n480 vss 3.80fF $ **FLOATING
C1416 out_p.n481 vss 3.85fF $ **FLOATING
C1417 out_p.n482 vss 3.81fF $ **FLOATING
C1418 out_p.n483 vss 3.87fF $ **FLOATING
C1419 out_p.n484 vss 4.05fF $ **FLOATING
C1420 out_p.n485 vss 4.05fF $ **FLOATING
C1421 out_p.n486 vss 4.05fF $ **FLOATING
C1422 out_p.n487 vss 4.15fF $ **FLOATING
C1423 out_p.n488 vss 4.15fF $ **FLOATING
C1424 out_p.n489 vss 4.05fF $ **FLOATING
C1425 out_p.n490 vss 4.05fF $ **FLOATING
C1426 out_p.n491 vss 4.05fF $ **FLOATING
C1427 out_p.n492 vss 3.80fF $ **FLOATING
C1428 out_p.n493 vss 3.85fF $ **FLOATING
C1429 out_p.n494 vss 3.81fF $ **FLOATING
C1430 out_p.n495 vss 3.87fF $ **FLOATING
C1431 out_p.n496 vss 4.05fF $ **FLOATING
C1432 out_p.n497 vss 4.05fF $ **FLOATING
C1433 out_p.n498 vss 4.05fF $ **FLOATING
C1434 out_p.n499 vss 4.15fF $ **FLOATING
C1435 out_p.n500 vss 4.15fF $ **FLOATING
C1436 out_p.n501 vss 4.05fF $ **FLOATING
C1437 out_p.n502 vss 4.05fF $ **FLOATING
C1438 out_p.n503 vss 4.05fF $ **FLOATING
C1439 out_p.n504 vss 3.80fF $ **FLOATING
C1440 out_p.n505 vss 3.85fF $ **FLOATING
C1441 out_p.n506 vss 3.81fF $ **FLOATING
C1442 out_p.n507 vss 3.87fF $ **FLOATING
C1443 out_p.n508 vss 4.05fF $ **FLOATING
C1444 out_p.n509 vss 4.05fF $ **FLOATING
C1445 out_p.n510 vss 4.05fF $ **FLOATING
C1446 out_p.n511 vss 4.15fF $ **FLOATING
C1447 out_p.n512 vss 4.15fF $ **FLOATING
C1448 out_p.n513 vss 4.05fF $ **FLOATING
C1449 out_p.n514 vss 4.05fF $ **FLOATING
C1450 out_p.n515 vss 4.05fF $ **FLOATING
C1451 out_p.n516 vss 3.80fF $ **FLOATING
C1452 out_p.n517 vss 3.85fF $ **FLOATING
C1453 out_p.n518 vss 3.81fF $ **FLOATING
C1454 out_p.n519 vss 3.87fF $ **FLOATING
C1455 out_p.n520 vss 4.05fF $ **FLOATING
C1456 out_p.n521 vss 4.05fF $ **FLOATING
C1457 out_p.n522 vss 4.05fF $ **FLOATING
C1458 out_p.n523 vss 4.15fF $ **FLOATING
C1459 out_p.n524 vss 4.15fF $ **FLOATING
C1460 out_p.n525 vss 4.05fF $ **FLOATING
C1461 out_p.n526 vss 4.05fF $ **FLOATING
C1462 out_p.n527 vss 4.05fF $ **FLOATING
C1463 out_p.n528 vss 3.80fF $ **FLOATING
C1464 out_p.n529 vss 3.85fF $ **FLOATING
C1465 out_p.n530 vss 3.81fF $ **FLOATING
C1466 out_p.n531 vss 3.87fF $ **FLOATING
C1467 out_p.n532 vss 4.05fF $ **FLOATING
C1468 out_p.n533 vss 4.05fF $ **FLOATING
C1469 out_p.n534 vss 4.05fF $ **FLOATING
C1470 out_p.n535 vss 4.15fF $ **FLOATING
C1471 out_p.n536 vss 4.15fF $ **FLOATING
C1472 out_p.n537 vss 4.05fF $ **FLOATING
C1473 out_p.n538 vss 4.05fF $ **FLOATING
C1474 out_p.n539 vss 4.05fF $ **FLOATING
C1475 out_p.n540 vss 3.80fF $ **FLOATING
C1476 out_p.n541 vss 3.85fF $ **FLOATING
C1477 out_p.n542 vss 3.81fF $ **FLOATING
C1478 out_p.n543 vss 3.87fF $ **FLOATING
C1479 out_p.n544 vss 4.05fF $ **FLOATING
C1480 out_p.n545 vss 4.05fF $ **FLOATING
C1481 out_p.n546 vss 4.05fF $ **FLOATING
C1482 out_p.n547 vss 4.15fF $ **FLOATING
C1483 out_p.n548 vss 4.15fF $ **FLOATING
C1484 out_p.n549 vss 4.05fF $ **FLOATING
C1485 out_p.n550 vss 4.05fF $ **FLOATING
C1486 out_p.n551 vss 4.05fF $ **FLOATING
C1487 out_p.n552 vss 3.80fF $ **FLOATING
C1488 out_p.n553 vss 3.85fF $ **FLOATING
C1489 out_p.n554 vss 3.81fF $ **FLOATING
C1490 out_p.n555 vss 3.87fF $ **FLOATING
C1491 out_p.n556 vss 4.05fF $ **FLOATING
C1492 out_p.n557 vss 4.05fF $ **FLOATING
C1493 out_p.n558 vss 4.05fF $ **FLOATING
C1494 out_p.n559 vss 4.15fF $ **FLOATING
C1495 out_p.n560 vss 4.15fF $ **FLOATING
C1496 out_p.n561 vss 4.05fF $ **FLOATING
C1497 out_p.n562 vss 4.05fF $ **FLOATING
C1498 out_p.n563 vss 4.05fF $ **FLOATING
C1499 out_p.n564 vss 3.80fF $ **FLOATING
C1500 out_p.n565 vss 3.85fF $ **FLOATING
C1501 out_p.n566 vss 3.81fF $ **FLOATING
C1502 out_p.n567 vss 3.87fF $ **FLOATING
C1503 out_p.n568 vss 4.05fF $ **FLOATING
C1504 out_p.n569 vss 4.05fF $ **FLOATING
C1505 out_p.n570 vss 4.05fF $ **FLOATING
C1506 out_p.n571 vss 4.15fF $ **FLOATING
C1507 out_p.n572 vss 4.15fF $ **FLOATING
C1508 out_p.n573 vss 4.05fF $ **FLOATING
C1509 out_p.n574 vss 4.05fF $ **FLOATING
C1510 out_p.n575 vss 4.05fF $ **FLOATING
C1511 out_p.n576 vss 3.80fF $ **FLOATING
C1512 out_p.n577 vss 3.85fF $ **FLOATING
C1513 out_p.n578 vss 3.81fF $ **FLOATING
C1514 out_p.n579 vss 3.87fF $ **FLOATING
C1515 out_p.n580 vss 4.05fF $ **FLOATING
C1516 out_p.n581 vss 4.05fF $ **FLOATING
C1517 out_p.n582 vss 4.05fF $ **FLOATING
C1518 out_p.n583 vss 4.15fF $ **FLOATING
C1519 out_p.n584 vss 4.15fF $ **FLOATING
C1520 out_p.n585 vss 4.05fF $ **FLOATING
C1521 out_p.n586 vss 4.05fF $ **FLOATING
C1522 out_p.n587 vss 4.05fF $ **FLOATING
C1523 out_p.n588 vss 3.80fF $ **FLOATING
C1524 out_p.n589 vss 3.85fF $ **FLOATING
C1525 out_p.n590 vss 3.81fF $ **FLOATING
C1526 out_p.n591 vss 3.87fF $ **FLOATING
C1527 out_p.n592 vss 4.05fF $ **FLOATING
C1528 out_p.n593 vss 4.05fF $ **FLOATING
C1529 out_p.n594 vss 4.05fF $ **FLOATING
C1530 out_p.n595 vss 4.15fF $ **FLOATING
C1531 out_p.n596 vss 4.15fF $ **FLOATING
C1532 out_p.n597 vss 4.05fF $ **FLOATING
C1533 out_p.n598 vss 4.05fF $ **FLOATING
C1534 out_p.n599 vss 4.05fF $ **FLOATING
C1535 out_p.n600 vss 3.80fF $ **FLOATING
C1536 out_p.n601 vss 3.85fF $ **FLOATING
C1537 out_p.n602 vss 3.81fF $ **FLOATING
C1538 out_p.n603 vss 3.87fF $ **FLOATING
C1539 out_p.n604 vss 4.05fF $ **FLOATING
C1540 out_p.n605 vss 4.05fF $ **FLOATING
C1541 out_p.n606 vss 4.05fF $ **FLOATING
C1542 out_p.n607 vss 4.15fF $ **FLOATING
C1543 out_p.n608 vss 4.15fF $ **FLOATING
C1544 out_p.n609 vss 4.05fF $ **FLOATING
C1545 out_p.n610 vss 4.05fF $ **FLOATING
C1546 out_p.n611 vss 4.05fF $ **FLOATING
C1547 out_p.n612 vss 3.80fF $ **FLOATING
C1548 out_p.n613 vss 3.85fF $ **FLOATING
C1549 out_p.n614 vss 3.81fF $ **FLOATING
C1550 out_p.n615 vss 3.87fF $ **FLOATING
C1551 out_p.n616 vss 4.05fF $ **FLOATING
C1552 out_p.n617 vss 4.05fF $ **FLOATING
C1553 out_p.n618 vss 4.05fF $ **FLOATING
C1554 out_p.n619 vss 4.15fF $ **FLOATING
C1555 out_p.n620 vss 4.15fF $ **FLOATING
C1556 out_p.n621 vss 4.05fF $ **FLOATING
C1557 out_p.n622 vss 4.05fF $ **FLOATING
C1558 out_p.n623 vss 4.05fF $ **FLOATING
C1559 out_p.n624 vss 3.80fF $ **FLOATING
C1560 out_p.n625 vss 3.85fF $ **FLOATING
C1561 out_p.n626 vss 3.81fF $ **FLOATING
C1562 out_p.n627 vss 3.87fF $ **FLOATING
C1563 out_p.n628 vss 4.05fF $ **FLOATING
C1564 out_p.n629 vss 4.05fF $ **FLOATING
C1565 out_p.n630 vss 4.05fF $ **FLOATING
C1566 out_p.n631 vss 4.15fF $ **FLOATING
C1567 out_p.n632 vss 4.15fF $ **FLOATING
C1568 out_p.n633 vss 4.05fF $ **FLOATING
C1569 out_p.n634 vss 4.05fF $ **FLOATING
C1570 out_p.n635 vss 4.05fF $ **FLOATING
C1571 out_p.n636 vss 3.80fF $ **FLOATING
C1572 out_p.n637 vss 3.85fF $ **FLOATING
C1573 out_p.n638 vss 3.81fF $ **FLOATING
C1574 out_p.n639 vss 3.87fF $ **FLOATING
C1575 out_p.n640 vss 4.05fF $ **FLOATING
C1576 out_p.n641 vss 4.05fF $ **FLOATING
C1577 out_p.n642 vss 4.05fF $ **FLOATING
C1578 out_p.n643 vss 4.15fF $ **FLOATING
C1579 out_p.n644 vss 4.15fF $ **FLOATING
C1580 out_p.n645 vss 4.05fF $ **FLOATING
C1581 out_p.n646 vss 4.05fF $ **FLOATING
C1582 out_p.n647 vss 4.05fF $ **FLOATING
C1583 out_p.n648 vss 3.80fF $ **FLOATING
C1584 out_p.n649 vss 3.85fF $ **FLOATING
C1585 out_p.n650 vss 3.81fF $ **FLOATING
C1586 out_p.n651 vss 3.87fF $ **FLOATING
C1587 out_p.n652 vss 4.05fF $ **FLOATING
C1588 out_p.n653 vss 4.05fF $ **FLOATING
C1589 out_p.n654 vss 4.05fF $ **FLOATING
C1590 out_p.n655 vss 4.15fF $ **FLOATING
C1591 out_p.n656 vss 4.15fF $ **FLOATING
C1592 out_p.n657 vss 4.05fF $ **FLOATING
C1593 out_p.n658 vss 4.05fF $ **FLOATING
C1594 out_p.n659 vss 4.05fF $ **FLOATING
C1595 out_p.n660 vss 3.80fF $ **FLOATING
C1596 out_p.n661 vss 3.85fF $ **FLOATING
C1597 out_p.n662 vss 3.81fF $ **FLOATING
C1598 out_p.n663 vss 3.87fF $ **FLOATING
C1599 out_p.n664 vss 4.05fF $ **FLOATING
C1600 out_p.n665 vss 4.05fF $ **FLOATING
C1601 out_p.n666 vss 4.05fF $ **FLOATING
C1602 out_p.n667 vss 4.15fF $ **FLOATING
C1603 out_p.n668 vss 4.15fF $ **FLOATING
C1604 out_p.n669 vss 4.05fF $ **FLOATING
C1605 out_p.n670 vss 4.05fF $ **FLOATING
C1606 out_p.n671 vss 4.05fF $ **FLOATING
C1607 out_p.n672 vss 3.80fF $ **FLOATING
C1608 out_p.n673 vss 3.85fF $ **FLOATING
C1609 out_p.n674 vss 3.81fF $ **FLOATING
C1610 out_p.n675 vss 3.87fF $ **FLOATING
C1611 out_p.n676 vss 4.05fF $ **FLOATING
C1612 out_p.n677 vss 4.05fF $ **FLOATING
C1613 out_p.n678 vss 4.05fF $ **FLOATING
C1614 out_p.n679 vss 4.15fF $ **FLOATING
C1615 out_p.n680 vss 4.15fF $ **FLOATING
C1616 out_p.n681 vss 4.05fF $ **FLOATING
C1617 out_p.n682 vss 4.05fF $ **FLOATING
C1618 out_p.n683 vss 4.05fF $ **FLOATING
C1619 out_p.n684 vss 3.80fF $ **FLOATING
C1620 out_p.n685 vss 3.85fF $ **FLOATING
C1621 out_p.n686 vss 3.81fF $ **FLOATING
C1622 out_p.n687 vss 3.87fF $ **FLOATING
C1623 out_p.n688 vss 4.05fF $ **FLOATING
C1624 out_p.n689 vss 4.05fF $ **FLOATING
C1625 out_p.n690 vss 4.05fF $ **FLOATING
C1626 out_p.n691 vss 4.15fF $ **FLOATING
C1627 out_p.n692 vss 4.15fF $ **FLOATING
C1628 out_p.n693 vss 4.05fF $ **FLOATING
C1629 out_p.n694 vss 4.05fF $ **FLOATING
C1630 out_p.n695 vss 4.05fF $ **FLOATING
C1631 out_p.n696 vss 3.80fF $ **FLOATING
C1632 out_p.n697 vss 3.85fF $ **FLOATING
C1633 out_p.n698 vss 3.81fF $ **FLOATING
C1634 out_p.n699 vss 3.87fF $ **FLOATING
C1635 out_p.n700 vss 4.05fF $ **FLOATING
C1636 out_p.n701 vss 4.05fF $ **FLOATING
C1637 out_p.n702 vss 4.05fF $ **FLOATING
C1638 out_p.n703 vss 4.15fF $ **FLOATING
C1639 out_p.n704 vss 4.15fF $ **FLOATING
C1640 out_p.n705 vss 4.05fF $ **FLOATING
C1641 out_p.n706 vss 4.05fF $ **FLOATING
C1642 out_p.n707 vss 4.05fF $ **FLOATING
C1643 out_p.n708 vss 3.80fF $ **FLOATING
C1644 out_p.n709 vss 3.85fF $ **FLOATING
C1645 out_p.n710 vss 3.81fF $ **FLOATING
C1646 out_p.n711 vss 3.87fF $ **FLOATING
C1647 out_p.n712 vss 4.05fF $ **FLOATING
C1648 out_p.n713 vss 4.05fF $ **FLOATING
C1649 out_p.n714 vss 4.05fF $ **FLOATING
C1650 out_p.n715 vss 4.15fF $ **FLOATING
C1651 out_p.n716 vss 4.15fF $ **FLOATING
C1652 out_p.n717 vss 4.05fF $ **FLOATING
C1653 out_p.n718 vss 4.05fF $ **FLOATING
C1654 out_p.n719 vss 4.05fF $ **FLOATING
C1655 out_p.n720 vss 3.80fF $ **FLOATING
C1656 out_p.n721 vss 3.85fF $ **FLOATING
C1657 out_p.n722 vss 3.81fF $ **FLOATING
C1658 out_p.n723 vss 3.87fF $ **FLOATING
C1659 out_p.n724 vss 4.05fF $ **FLOATING
C1660 out_p.n725 vss 4.05fF $ **FLOATING
C1661 out_p.n726 vss 4.05fF $ **FLOATING
C1662 out_p.n727 vss 4.15fF $ **FLOATING
C1663 out_p.n728 vss 4.15fF $ **FLOATING
C1664 out_p.n729 vss 4.05fF $ **FLOATING
C1665 out_p.n730 vss 4.05fF $ **FLOATING
C1666 out_p.n731 vss 4.05fF $ **FLOATING
C1667 out_p.n732 vss 3.80fF $ **FLOATING
C1668 out_p.n733 vss 3.85fF $ **FLOATING
C1669 out_p.n734 vss 3.81fF $ **FLOATING
C1670 out_p.n735 vss 3.87fF $ **FLOATING
C1671 out_p.n736 vss 4.05fF $ **FLOATING
C1672 out_p.n737 vss 4.05fF $ **FLOATING
C1673 out_p.n738 vss 4.05fF $ **FLOATING
C1674 out_p.n739 vss 4.15fF $ **FLOATING
C1675 out_p.n740 vss 4.15fF $ **FLOATING
C1676 out_p.n741 vss 4.05fF $ **FLOATING
C1677 out_p.n742 vss 4.05fF $ **FLOATING
C1678 out_p.n743 vss 4.05fF $ **FLOATING
C1679 out_p.n744 vss 3.80fF $ **FLOATING
C1680 out_p.n745 vss 3.85fF $ **FLOATING
C1681 out_p.n746 vss 3.81fF $ **FLOATING
C1682 out_p.n747 vss 3.87fF $ **FLOATING
C1683 out_p.n748 vss 4.05fF $ **FLOATING
C1684 out_p.n749 vss 4.05fF $ **FLOATING
C1685 out_p.n750 vss 4.05fF $ **FLOATING
C1686 out_p.n751 vss 4.15fF $ **FLOATING
C1687 out_p.n752 vss 4.15fF $ **FLOATING
C1688 out_p.n753 vss 4.05fF $ **FLOATING
C1689 out_p.n754 vss 4.05fF $ **FLOATING
C1690 out_p.n755 vss 4.05fF $ **FLOATING
C1691 out_p.n756 vss 3.80fF $ **FLOATING
C1692 out_p.n757 vss 3.85fF $ **FLOATING
C1693 out_p.n758 vss 3.81fF $ **FLOATING
C1694 out_p.n759 vss 3.87fF $ **FLOATING
C1695 out_p.n760 vss 4.05fF $ **FLOATING
C1696 out_p.n761 vss 4.05fF $ **FLOATING
C1697 out_p.n762 vss 4.05fF $ **FLOATING
C1698 out_p.n763 vss 4.15fF $ **FLOATING
C1699 out_p.n764 vss 4.15fF $ **FLOATING
C1700 out_p.n765 vss 4.05fF $ **FLOATING
C1701 out_p.n766 vss 4.05fF $ **FLOATING
C1702 out_p.n767 vss 4.05fF $ **FLOATING
C1703 out_p.n768 vss 3.80fF $ **FLOATING
C1704 out_p.n769 vss 3.85fF $ **FLOATING
C1705 out_p.n770 vss 3.81fF $ **FLOATING
C1706 out_p.n771 vss 3.87fF $ **FLOATING
C1707 out_p.n772 vss 4.05fF $ **FLOATING
C1708 out_p.n773 vss 4.05fF $ **FLOATING
C1709 out_p.n774 vss 4.05fF $ **FLOATING
C1710 out_p.n775 vss 4.15fF $ **FLOATING
C1711 out_p.n776 vss 4.15fF $ **FLOATING
C1712 out_p.n777 vss 4.05fF $ **FLOATING
C1713 out_p.n778 vss 4.05fF $ **FLOATING
C1714 out_p.n779 vss 4.05fF $ **FLOATING
C1715 out_p.n780 vss 3.80fF $ **FLOATING
C1716 out_p.n781 vss 3.85fF $ **FLOATING
C1717 out_p.n782 vss 3.81fF $ **FLOATING
C1718 out_p.n783 vss 3.87fF $ **FLOATING
C1719 out_p.n784 vss 4.05fF $ **FLOATING
C1720 out_p.n785 vss 4.05fF $ **FLOATING
C1721 out_p.n786 vss 4.05fF $ **FLOATING
C1722 out_p.n787 vss 4.15fF $ **FLOATING
C1723 out_p.n788 vss 4.15fF $ **FLOATING
C1724 out_p.n789 vss 4.05fF $ **FLOATING
C1725 out_p.n790 vss 4.05fF $ **FLOATING
C1726 out_p.n791 vss 4.05fF $ **FLOATING
C1727 out_p.n792 vss 3.80fF $ **FLOATING
C1728 out_p.n793 vss 3.85fF $ **FLOATING
C1729 out_p.n794 vss 3.81fF $ **FLOATING
C1730 out_p.n795 vss 3.87fF $ **FLOATING
C1731 out_p.n796 vss 4.05fF $ **FLOATING
C1732 out_p.n797 vss 4.05fF $ **FLOATING
C1733 out_p.n798 vss 4.05fF $ **FLOATING
C1734 out_p.n799 vss 4.15fF $ **FLOATING
C1735 out_p.n800 vss 4.15fF $ **FLOATING
C1736 out_p.n801 vss 4.05fF $ **FLOATING
C1737 out_p.n802 vss 4.05fF $ **FLOATING
C1738 out_p.n803 vss 4.05fF $ **FLOATING
C1739 out_p.n804 vss 3.80fF $ **FLOATING
C1740 out_p.n805 vss 3.85fF $ **FLOATING
C1741 out_p.n806 vss 3.81fF $ **FLOATING
C1742 out_p.n807 vss 3.87fF $ **FLOATING
C1743 out_p.n808 vss 4.05fF $ **FLOATING
C1744 out_p.n809 vss 4.05fF $ **FLOATING
C1745 out_p.n810 vss 4.05fF $ **FLOATING
C1746 out_p.n811 vss 4.15fF $ **FLOATING
C1747 out_p.n812 vss 4.15fF $ **FLOATING
C1748 out_p.n813 vss 4.05fF $ **FLOATING
C1749 out_p.n814 vss 4.05fF $ **FLOATING
C1750 out_p.n815 vss 4.05fF $ **FLOATING
C1751 out_p.n816 vss 3.80fF $ **FLOATING
C1752 out_p.n817 vss 3.85fF $ **FLOATING
C1753 out_p.n818 vss 3.81fF $ **FLOATING
C1754 out_p.n819 vss 3.87fF $ **FLOATING
C1755 out_p.n820 vss 4.05fF $ **FLOATING
C1756 out_p.n821 vss 4.05fF $ **FLOATING
C1757 out_p.n822 vss 4.05fF $ **FLOATING
C1758 out_p.n823 vss 4.15fF $ **FLOATING
C1759 out_p.n824 vss 4.15fF $ **FLOATING
C1760 out_p.n825 vss 4.05fF $ **FLOATING
C1761 out_p.n826 vss 4.05fF $ **FLOATING
C1762 out_p.n827 vss 4.05fF $ **FLOATING
C1763 out_p.n828 vss 3.80fF $ **FLOATING
C1764 out_p.n829 vss 3.85fF $ **FLOATING
C1765 out_p.n830 vss 3.81fF $ **FLOATING
C1766 out_p.n831 vss 3.87fF $ **FLOATING
C1767 out_p.n832 vss 4.05fF $ **FLOATING
C1768 out_p.n833 vss 4.05fF $ **FLOATING
C1769 out_p.n834 vss 4.05fF $ **FLOATING
C1770 out_p.n835 vss 4.15fF $ **FLOATING
C1771 out_p.n836 vss 4.15fF $ **FLOATING
C1772 out_p.n837 vss 4.05fF $ **FLOATING
C1773 out_p.n838 vss 4.05fF $ **FLOATING
C1774 out_p.n839 vss 4.05fF $ **FLOATING
C1775 out_p.n840 vss 3.80fF $ **FLOATING
C1776 out_p.n841 vss 3.85fF $ **FLOATING
C1777 out_p.n842 vss 3.81fF $ **FLOATING
C1778 out_p.n843 vss 3.87fF $ **FLOATING
C1779 out_p.n844 vss 4.05fF $ **FLOATING
C1780 out_p.n845 vss 4.05fF $ **FLOATING
C1781 out_p.n846 vss 4.05fF $ **FLOATING
C1782 out_p.n847 vss 4.15fF $ **FLOATING
C1783 out_p.n848 vss 4.15fF $ **FLOATING
C1784 out_p.n849 vss 4.05fF $ **FLOATING
C1785 out_p.n850 vss 4.05fF $ **FLOATING
C1786 out_p.n851 vss 4.05fF $ **FLOATING
C1787 out_p.n852 vss 3.80fF $ **FLOATING
C1788 out_p.n853 vss 3.85fF $ **FLOATING
C1789 out_p.n854 vss 3.81fF $ **FLOATING
C1790 out_p.n855 vss 3.87fF $ **FLOATING
C1791 out_p.n856 vss 4.05fF $ **FLOATING
C1792 out_p.n857 vss 4.05fF $ **FLOATING
C1793 out_p.n858 vss 4.05fF $ **FLOATING
C1794 out_p.n859 vss 4.15fF $ **FLOATING
C1795 out_p.n860 vss 4.15fF $ **FLOATING
C1796 out_p.n861 vss 4.05fF $ **FLOATING
C1797 out_p.n862 vss 4.05fF $ **FLOATING
C1798 out_p.n863 vss 4.05fF $ **FLOATING
C1799 out_p.n864 vss 3.80fF $ **FLOATING
C1800 out_p.n865 vss 3.85fF $ **FLOATING
C1801 out_p.n866 vss 3.81fF $ **FLOATING
C1802 out_p.n867 vss 3.87fF $ **FLOATING
C1803 out_p.n868 vss 4.05fF $ **FLOATING
C1804 out_p.n869 vss 4.05fF $ **FLOATING
C1805 out_p.n870 vss 4.05fF $ **FLOATING
C1806 out_p.n871 vss 4.15fF $ **FLOATING
C1807 out_p.n872 vss 4.15fF $ **FLOATING
C1808 out_p.n873 vss 4.05fF $ **FLOATING
C1809 out_p.n874 vss 4.05fF $ **FLOATING
C1810 out_p.n875 vss 4.05fF $ **FLOATING
C1811 out_p.n876 vss 3.80fF $ **FLOATING
C1812 out_p.n877 vss 3.85fF $ **FLOATING
C1813 out_p.n878 vss 3.81fF $ **FLOATING
C1814 out_p.n879 vss 3.87fF $ **FLOATING
C1815 out_p.n880 vss 4.05fF $ **FLOATING
C1816 out_p.n881 vss 4.05fF $ **FLOATING
C1817 out_p.n882 vss 4.05fF $ **FLOATING
C1818 out_p.n883 vss 4.15fF $ **FLOATING
C1819 out_p.n884 vss 4.15fF $ **FLOATING
C1820 out_p.n885 vss 4.05fF $ **FLOATING
C1821 out_p.n886 vss 4.05fF $ **FLOATING
C1822 out_p.n887 vss 4.05fF $ **FLOATING
C1823 out_p.n888 vss 3.80fF $ **FLOATING
C1824 out_p.n889 vss 3.85fF $ **FLOATING
C1825 out_p.n890 vss 3.81fF $ **FLOATING
C1826 out_p.n891 vss 3.87fF $ **FLOATING
C1827 out_p.n892 vss 4.05fF $ **FLOATING
C1828 out_p.n893 vss 4.05fF $ **FLOATING
C1829 out_p.n894 vss 4.05fF $ **FLOATING
C1830 out_p.n895 vss 4.15fF $ **FLOATING
C1831 out_p.n896 vss 4.15fF $ **FLOATING
C1832 out_p.n897 vss 4.05fF $ **FLOATING
C1833 out_p.n898 vss 4.05fF $ **FLOATING
C1834 out_p.n899 vss 4.05fF $ **FLOATING
C1835 out_p.n900 vss 3.80fF $ **FLOATING
C1836 out_p.n901 vss 3.85fF $ **FLOATING
C1837 out_p.n902 vss 3.81fF $ **FLOATING
C1838 out_p.n903 vss 3.86fF $ **FLOATING
C1839 out_p.n904 vss 4.05fF $ **FLOATING
C1840 out_p.n905 vss 4.05fF $ **FLOATING
C1841 out_p.n906 vss 4.05fF $ **FLOATING
C1842 out_p.n907 vss 4.15fF $ **FLOATING
C1843 out_p.n908 vss 4.15fF $ **FLOATING
C1844 out_p.n909 vss 4.05fF $ **FLOATING
C1845 out_p.n910 vss 4.05fF $ **FLOATING
C1846 out_p.n911 vss 4.05fF $ **FLOATING
C1847 out_p.n912 vss 3.81fF $ **FLOATING
C1848 out_p.n913 vss 23.47fF $ **FLOATING
C1849 out_p.n914 vss 30.23fF $ **FLOATING
C1850 out_p.n915 vss 30.23fF $ **FLOATING
C1851 out_p.n916 vss 30.23fF $ **FLOATING
C1852 out_p.n917 vss 30.23fF $ **FLOATING
C1853 out_p.n918 vss 30.23fF $ **FLOATING
C1854 out_p.n919 vss 30.23fF $ **FLOATING
C1855 out_p.n920 vss 30.23fF $ **FLOATING
C1856 out_p.n921 vss 30.23fF $ **FLOATING
C1857 out_p.n922 vss 30.23fF $ **FLOATING
C1858 out_p.n923 vss 30.23fF $ **FLOATING
C1859 out_p.n924 vss 30.23fF $ **FLOATING
C1860 out_p.n925 vss 30.23fF $ **FLOATING
C1861 out_p.n926 vss 30.23fF $ **FLOATING
C1862 out_p.n927 vss 30.23fF $ **FLOATING
C1863 out_p.n928 vss 30.23fF $ **FLOATING
C1864 out_p.n929 vss 30.23fF $ **FLOATING
C1865 out_p.n930 vss 30.23fF $ **FLOATING
C1866 out_p.n931 vss 30.23fF $ **FLOATING
C1867 out_p.n932 vss 30.23fF $ **FLOATING
C1868 out_p.n933 vss 30.23fF $ **FLOATING
C1869 out_p.n934 vss 30.23fF $ **FLOATING
C1870 out_p.n935 vss 30.23fF $ **FLOATING
C1871 out_p.n936 vss 30.23fF $ **FLOATING
C1872 out_p.n937 vss 30.23fF $ **FLOATING
C1873 out_p.n938 vss 30.23fF $ **FLOATING
C1874 out_p.n939 vss 30.23fF $ **FLOATING
C1875 out_p.n940 vss 30.23fF $ **FLOATING
C1876 out_p.n941 vss 30.23fF $ **FLOATING
C1877 out_p.n942 vss 30.23fF $ **FLOATING
C1878 out_p.n943 vss 30.23fF $ **FLOATING
C1879 out_p.n944 vss 30.23fF $ **FLOATING
C1880 out_p.n945 vss 30.23fF $ **FLOATING
C1881 out_p.n946 vss 30.23fF $ **FLOATING
C1882 out_p.n947 vss 30.23fF $ **FLOATING
C1883 out_p.n948 vss 30.23fF $ **FLOATING
C1884 out_p.n949 vss 30.23fF $ **FLOATING
C1885 out_p.n950 vss 30.23fF $ **FLOATING
C1886 out_p.n951 vss 30.23fF $ **FLOATING
C1887 out_p.n952 vss 30.23fF $ **FLOATING
C1888 out_p.n953 vss 30.23fF $ **FLOATING
C1889 out_p.n954 vss 30.23fF $ **FLOATING
C1890 out_p.n955 vss 30.23fF $ **FLOATING
C1891 out_p.n956 vss 30.23fF $ **FLOATING
C1892 out_p.n957 vss 30.23fF $ **FLOATING
C1893 out_p.n958 vss 30.23fF $ **FLOATING
C1894 out_p.n959 vss 30.23fF $ **FLOATING
C1895 out_p.n960 vss 30.23fF $ **FLOATING
C1896 out_p.n961 vss 30.23fF $ **FLOATING
C1897 out_p.n962 vss 30.23fF $ **FLOATING
C1898 out_p.n963 vss 30.23fF $ **FLOATING
C1899 out_p.n964 vss 30.23fF $ **FLOATING
C1900 out_p.n965 vss 30.23fF $ **FLOATING
C1901 out_p.n966 vss 30.23fF $ **FLOATING
C1902 out_p.n967 vss 30.23fF $ **FLOATING
C1903 out_p.n968 vss 30.23fF $ **FLOATING
C1904 out_p.n969 vss 30.23fF $ **FLOATING
C1905 out_p.n970 vss 30.23fF $ **FLOATING
C1906 out_p.n971 vss 30.23fF $ **FLOATING
C1907 out_p.n972 vss 30.23fF $ **FLOATING
C1908 out_p.n973 vss 29.52fF $ **FLOATING
C1909 vp_p.n0 vss 1.04fF $ **FLOATING
C1910 vp_p.n76 vss 1.09fF $ **FLOATING
C1911 vp_p.n78 vss 1.03fF $ **FLOATING
C1912 vp_p.n80 vss 1.03fF $ **FLOATING
C1913 vp_p.n82 vss 1.03fF $ **FLOATING
C1914 vp_p.n84 vss 1.03fF $ **FLOATING
C1915 vp_p.n86 vss 1.03fF $ **FLOATING
C1916 vp_p.n88 vss 1.03fF $ **FLOATING
C1917 vp_p.n90 vss 1.03fF $ **FLOATING
C1918 vp_p.n92 vss 1.03fF $ **FLOATING
C1919 vp_p.n94 vss 1.03fF $ **FLOATING
C1920 vp_p.n96 vss 1.03fF $ **FLOATING
C1921 vp_p.n98 vss 1.03fF $ **FLOATING
C1922 vp_p.n100 vss 1.03fF $ **FLOATING
C1923 vp_p.n102 vss 1.03fF $ **FLOATING
C1924 vp_p.n104 vss 1.03fF $ **FLOATING
C1925 vp_p.n106 vss 1.03fF $ **FLOATING
C1926 vp_p.n108 vss 1.03fF $ **FLOATING
C1927 vp_p.n110 vss 1.03fF $ **FLOATING
C1928 vp_p.n112 vss 1.03fF $ **FLOATING
C1929 vp_p.n114 vss 1.03fF $ **FLOATING
C1930 vp_p.n116 vss 1.03fF $ **FLOATING
C1931 vp_p.n118 vss 1.03fF $ **FLOATING
C1932 vp_p.n120 vss 1.03fF $ **FLOATING
C1933 vp_p.n122 vss 1.03fF $ **FLOATING
C1934 vp_p.n124 vss 1.03fF $ **FLOATING
C1935 vp_p.n126 vss 1.03fF $ **FLOATING
C1936 vp_p.n128 vss 1.03fF $ **FLOATING
C1937 vp_p.n130 vss 1.03fF $ **FLOATING
C1938 vp_p.n132 vss 1.03fF $ **FLOATING
C1939 vp_p.n134 vss 1.03fF $ **FLOATING
C1940 vp_p.n136 vss 1.03fF $ **FLOATING
C1941 vp_p.n138 vss 1.03fF $ **FLOATING
C1942 vp_p.n140 vss 1.03fF $ **FLOATING
C1943 vp_p.n142 vss 1.03fF $ **FLOATING
C1944 vp_p.n144 vss 1.03fF $ **FLOATING
C1945 vp_p.n146 vss 1.03fF $ **FLOATING
C1946 vp_p.n148 vss 1.03fF $ **FLOATING
C1947 vp_p.n150 vss 1.03fF $ **FLOATING
C1948 vp_p.n152 vss 1.03fF $ **FLOATING
C1949 vp_p.n154 vss 1.03fF $ **FLOATING
C1950 vp_p.n156 vss 1.03fF $ **FLOATING
C1951 vp_p.n158 vss 1.03fF $ **FLOATING
C1952 vp_p.n160 vss 1.03fF $ **FLOATING
C1953 vp_p.n162 vss 1.03fF $ **FLOATING
C1954 vp_p.n164 vss 1.03fF $ **FLOATING
C1955 vp_p.n166 vss 1.03fF $ **FLOATING
C1956 vp_p.n168 vss 1.03fF $ **FLOATING
C1957 vp_p.n170 vss 1.03fF $ **FLOATING
C1958 vp_p.n172 vss 1.03fF $ **FLOATING
C1959 vp_p.n174 vss 1.03fF $ **FLOATING
C1960 vp_p.n176 vss 1.03fF $ **FLOATING
C1961 vp_p.n178 vss 1.03fF $ **FLOATING
C1962 vp_p.n180 vss 1.03fF $ **FLOATING
C1963 vp_p.n182 vss 1.03fF $ **FLOATING
C1964 vp_p.n184 vss 1.03fF $ **FLOATING
C1965 vp_p.n186 vss 1.03fF $ **FLOATING
C1966 vp_p.n188 vss 1.03fF $ **FLOATING
C1967 vp_p.n190 vss 1.03fF $ **FLOATING
C1968 vp_p.n192 vss 1.03fF $ **FLOATING
C1969 vp_p.n194 vss 1.03fF $ **FLOATING
C1970 vp_p.n196 vss 1.03fF $ **FLOATING
C1971 vp_p.n198 vss 1.03fF $ **FLOATING
C1972 vp_p.n200 vss 1.03fF $ **FLOATING
C1973 vp_p.n202 vss 1.03fF $ **FLOATING
C1974 vp_p.n204 vss 1.03fF $ **FLOATING
C1975 vp_p.n206 vss 1.03fF $ **FLOATING
C1976 vp_p.n208 vss 1.03fF $ **FLOATING
C1977 vp_p.n210 vss 1.03fF $ **FLOATING
C1978 vp_p.n212 vss 1.03fF $ **FLOATING
C1979 vp_p.n214 vss 1.03fF $ **FLOATING
C1980 vp_p.n216 vss 1.03fF $ **FLOATING
C1981 vp_p.n218 vss 1.03fF $ **FLOATING
C1982 vp_p.n220 vss 1.03fF $ **FLOATING
C1983 vp_p.n225 vss 1.09fF $ **FLOATING
C1984 vp_p.n227 vss 1.03fF $ **FLOATING
C1985 vp_p.n229 vss 1.03fF $ **FLOATING
C1986 vp_p.n231 vss 1.03fF $ **FLOATING
C1987 vp_p.n233 vss 1.03fF $ **FLOATING
C1988 vp_p.n235 vss 1.03fF $ **FLOATING
C1989 vp_p.n237 vss 1.03fF $ **FLOATING
C1990 vp_p.n239 vss 1.03fF $ **FLOATING
C1991 vp_p.n241 vss 1.03fF $ **FLOATING
C1992 vp_p.n243 vss 1.03fF $ **FLOATING
C1993 vp_p.n245 vss 1.03fF $ **FLOATING
C1994 vp_p.n247 vss 1.03fF $ **FLOATING
C1995 vp_p.n249 vss 1.03fF $ **FLOATING
C1996 vp_p.n251 vss 1.03fF $ **FLOATING
C1997 vp_p.n253 vss 1.03fF $ **FLOATING
C1998 vp_p.n255 vss 1.03fF $ **FLOATING
C1999 vp_p.n257 vss 1.03fF $ **FLOATING
C2000 vp_p.n259 vss 1.03fF $ **FLOATING
C2001 vp_p.n261 vss 1.03fF $ **FLOATING
C2002 vp_p.n263 vss 1.03fF $ **FLOATING
C2003 vp_p.n265 vss 1.03fF $ **FLOATING
C2004 vp_p.n267 vss 1.03fF $ **FLOATING
C2005 vp_p.n269 vss 1.03fF $ **FLOATING
C2006 vp_p.n271 vss 1.03fF $ **FLOATING
C2007 vp_p.n273 vss 1.03fF $ **FLOATING
C2008 vp_p.n275 vss 1.03fF $ **FLOATING
C2009 vp_p.n277 vss 1.03fF $ **FLOATING
C2010 vp_p.n279 vss 1.03fF $ **FLOATING
C2011 vp_p.n281 vss 1.03fF $ **FLOATING
C2012 vp_p.n283 vss 1.03fF $ **FLOATING
C2013 vp_p.n285 vss 1.03fF $ **FLOATING
C2014 vp_p.n287 vss 1.03fF $ **FLOATING
C2015 vp_p.n289 vss 1.03fF $ **FLOATING
C2016 vp_p.n291 vss 1.03fF $ **FLOATING
C2017 vp_p.n293 vss 1.03fF $ **FLOATING
C2018 vp_p.n295 vss 1.03fF $ **FLOATING
C2019 vp_p.n297 vss 1.03fF $ **FLOATING
C2020 vp_p.n299 vss 1.03fF $ **FLOATING
C2021 vp_p.n301 vss 1.03fF $ **FLOATING
C2022 vp_p.n303 vss 1.03fF $ **FLOATING
C2023 vp_p.n305 vss 1.03fF $ **FLOATING
C2024 vp_p.n307 vss 1.03fF $ **FLOATING
C2025 vp_p.n309 vss 1.03fF $ **FLOATING
C2026 vp_p.n311 vss 1.03fF $ **FLOATING
C2027 vp_p.n313 vss 1.03fF $ **FLOATING
C2028 vp_p.n315 vss 1.03fF $ **FLOATING
C2029 vp_p.n317 vss 1.03fF $ **FLOATING
C2030 vp_p.n319 vss 1.03fF $ **FLOATING
C2031 vp_p.n321 vss 1.03fF $ **FLOATING
C2032 vp_p.n323 vss 1.03fF $ **FLOATING
C2033 vp_p.n325 vss 1.03fF $ **FLOATING
C2034 vp_p.n327 vss 1.03fF $ **FLOATING
C2035 vp_p.n329 vss 1.03fF $ **FLOATING
C2036 vp_p.n331 vss 1.03fF $ **FLOATING
C2037 vp_p.n333 vss 1.03fF $ **FLOATING
C2038 vp_p.n335 vss 1.03fF $ **FLOATING
C2039 vp_p.n337 vss 1.03fF $ **FLOATING
C2040 vp_p.n339 vss 1.03fF $ **FLOATING
C2041 vp_p.n341 vss 1.03fF $ **FLOATING
C2042 vp_p.n343 vss 1.03fF $ **FLOATING
C2043 vp_p.n345 vss 1.03fF $ **FLOATING
C2044 vp_p.n347 vss 1.03fF $ **FLOATING
C2045 vp_p.n349 vss 1.03fF $ **FLOATING
C2046 vp_p.n351 vss 1.03fF $ **FLOATING
C2047 vp_p.n353 vss 1.03fF $ **FLOATING
C2048 vp_p.n355 vss 1.03fF $ **FLOATING
C2049 vp_p.n357 vss 1.03fF $ **FLOATING
C2050 vp_p.n359 vss 1.03fF $ **FLOATING
C2051 vp_p.n361 vss 1.03fF $ **FLOATING
C2052 vp_p.n363 vss 1.03fF $ **FLOATING
C2053 vp_p.n365 vss 1.03fF $ **FLOATING
C2054 vp_p.n367 vss 1.03fF $ **FLOATING
C2055 vp_p.n369 vss 1.03fF $ **FLOATING
C2056 vp_p.n374 vss 1.09fF $ **FLOATING
C2057 vp_p.n376 vss 1.03fF $ **FLOATING
C2058 vp_p.n378 vss 1.03fF $ **FLOATING
C2059 vp_p.n380 vss 1.03fF $ **FLOATING
C2060 vp_p.n382 vss 1.03fF $ **FLOATING
C2061 vp_p.n384 vss 1.03fF $ **FLOATING
C2062 vp_p.n386 vss 1.03fF $ **FLOATING
C2063 vp_p.n388 vss 1.03fF $ **FLOATING
C2064 vp_p.n390 vss 1.03fF $ **FLOATING
C2065 vp_p.n392 vss 1.03fF $ **FLOATING
C2066 vp_p.n394 vss 1.03fF $ **FLOATING
C2067 vp_p.n396 vss 1.03fF $ **FLOATING
C2068 vp_p.n398 vss 1.03fF $ **FLOATING
C2069 vp_p.n400 vss 1.03fF $ **FLOATING
C2070 vp_p.n402 vss 1.03fF $ **FLOATING
C2071 vp_p.n404 vss 1.03fF $ **FLOATING
C2072 vp_p.n406 vss 1.03fF $ **FLOATING
C2073 vp_p.n408 vss 1.03fF $ **FLOATING
C2074 vp_p.n410 vss 1.03fF $ **FLOATING
C2075 vp_p.n412 vss 1.03fF $ **FLOATING
C2076 vp_p.n414 vss 1.03fF $ **FLOATING
C2077 vp_p.n416 vss 1.03fF $ **FLOATING
C2078 vp_p.n418 vss 1.03fF $ **FLOATING
C2079 vp_p.n420 vss 1.03fF $ **FLOATING
C2080 vp_p.n422 vss 1.03fF $ **FLOATING
C2081 vp_p.n424 vss 1.03fF $ **FLOATING
C2082 vp_p.n426 vss 1.03fF $ **FLOATING
C2083 vp_p.n428 vss 1.03fF $ **FLOATING
C2084 vp_p.n430 vss 1.03fF $ **FLOATING
C2085 vp_p.n432 vss 1.03fF $ **FLOATING
C2086 vp_p.n434 vss 1.03fF $ **FLOATING
C2087 vp_p.n436 vss 1.03fF $ **FLOATING
C2088 vp_p.n438 vss 1.03fF $ **FLOATING
C2089 vp_p.n440 vss 1.03fF $ **FLOATING
C2090 vp_p.n442 vss 1.03fF $ **FLOATING
C2091 vp_p.n444 vss 1.03fF $ **FLOATING
C2092 vp_p.n446 vss 1.03fF $ **FLOATING
C2093 vp_p.n448 vss 1.03fF $ **FLOATING
C2094 vp_p.n450 vss 1.03fF $ **FLOATING
C2095 vp_p.n452 vss 1.03fF $ **FLOATING
C2096 vp_p.n454 vss 1.03fF $ **FLOATING
C2097 vp_p.n456 vss 1.03fF $ **FLOATING
C2098 vp_p.n458 vss 1.03fF $ **FLOATING
C2099 vp_p.n460 vss 1.03fF $ **FLOATING
C2100 vp_p.n462 vss 1.03fF $ **FLOATING
C2101 vp_p.n464 vss 1.03fF $ **FLOATING
C2102 vp_p.n466 vss 1.03fF $ **FLOATING
C2103 vp_p.n468 vss 1.03fF $ **FLOATING
C2104 vp_p.n470 vss 1.03fF $ **FLOATING
C2105 vp_p.n472 vss 1.03fF $ **FLOATING
C2106 vp_p.n474 vss 1.03fF $ **FLOATING
C2107 vp_p.n476 vss 1.03fF $ **FLOATING
C2108 vp_p.n478 vss 1.03fF $ **FLOATING
C2109 vp_p.n480 vss 1.03fF $ **FLOATING
C2110 vp_p.n482 vss 1.03fF $ **FLOATING
C2111 vp_p.n484 vss 1.03fF $ **FLOATING
C2112 vp_p.n486 vss 1.03fF $ **FLOATING
C2113 vp_p.n488 vss 1.03fF $ **FLOATING
C2114 vp_p.n490 vss 1.03fF $ **FLOATING
C2115 vp_p.n492 vss 1.03fF $ **FLOATING
C2116 vp_p.n494 vss 1.03fF $ **FLOATING
C2117 vp_p.n496 vss 1.03fF $ **FLOATING
C2118 vp_p.n498 vss 1.03fF $ **FLOATING
C2119 vp_p.n500 vss 1.03fF $ **FLOATING
C2120 vp_p.n502 vss 1.03fF $ **FLOATING
C2121 vp_p.n504 vss 1.03fF $ **FLOATING
C2122 vp_p.n506 vss 1.03fF $ **FLOATING
C2123 vp_p.n508 vss 1.03fF $ **FLOATING
C2124 vp_p.n510 vss 1.03fF $ **FLOATING
C2125 vp_p.n512 vss 1.03fF $ **FLOATING
C2126 vp_p.n514 vss 1.03fF $ **FLOATING
C2127 vp_p.n516 vss 1.03fF $ **FLOATING
C2128 vp_p.n518 vss 1.03fF $ **FLOATING
C2129 vp_p.n523 vss 1.09fF $ **FLOATING
C2130 vp_p.n525 vss 1.03fF $ **FLOATING
C2131 vp_p.n527 vss 1.03fF $ **FLOATING
C2132 vp_p.n529 vss 1.03fF $ **FLOATING
C2133 vp_p.n531 vss 1.03fF $ **FLOATING
C2134 vp_p.n533 vss 1.03fF $ **FLOATING
C2135 vp_p.n535 vss 1.03fF $ **FLOATING
C2136 vp_p.n537 vss 1.03fF $ **FLOATING
C2137 vp_p.n539 vss 1.03fF $ **FLOATING
C2138 vp_p.n541 vss 1.03fF $ **FLOATING
C2139 vp_p.n543 vss 1.03fF $ **FLOATING
C2140 vp_p.n545 vss 1.03fF $ **FLOATING
C2141 vp_p.n547 vss 1.03fF $ **FLOATING
C2142 vp_p.n549 vss 1.03fF $ **FLOATING
C2143 vp_p.n551 vss 1.03fF $ **FLOATING
C2144 vp_p.n553 vss 1.03fF $ **FLOATING
C2145 vp_p.n555 vss 1.03fF $ **FLOATING
C2146 vp_p.n557 vss 1.03fF $ **FLOATING
C2147 vp_p.n559 vss 1.03fF $ **FLOATING
C2148 vp_p.n561 vss 1.03fF $ **FLOATING
C2149 vp_p.n563 vss 1.03fF $ **FLOATING
C2150 vp_p.n565 vss 1.03fF $ **FLOATING
C2151 vp_p.n567 vss 1.03fF $ **FLOATING
C2152 vp_p.n569 vss 1.03fF $ **FLOATING
C2153 vp_p.n571 vss 1.03fF $ **FLOATING
C2154 vp_p.n573 vss 1.03fF $ **FLOATING
C2155 vp_p.n575 vss 1.03fF $ **FLOATING
C2156 vp_p.n577 vss 1.03fF $ **FLOATING
C2157 vp_p.n579 vss 1.03fF $ **FLOATING
C2158 vp_p.n581 vss 1.03fF $ **FLOATING
C2159 vp_p.n583 vss 1.03fF $ **FLOATING
C2160 vp_p.n585 vss 1.03fF $ **FLOATING
C2161 vp_p.n587 vss 1.03fF $ **FLOATING
C2162 vp_p.n589 vss 1.03fF $ **FLOATING
C2163 vp_p.n591 vss 1.03fF $ **FLOATING
C2164 vp_p.n593 vss 1.03fF $ **FLOATING
C2165 vp_p.n595 vss 1.03fF $ **FLOATING
C2166 vp_p.n597 vss 1.03fF $ **FLOATING
C2167 vp_p.n599 vss 1.03fF $ **FLOATING
C2168 vp_p.n601 vss 1.03fF $ **FLOATING
C2169 vp_p.n603 vss 1.03fF $ **FLOATING
C2170 vp_p.n605 vss 1.03fF $ **FLOATING
C2171 vp_p.n607 vss 1.03fF $ **FLOATING
C2172 vp_p.n609 vss 1.03fF $ **FLOATING
C2173 vp_p.n611 vss 1.03fF $ **FLOATING
C2174 vp_p.n613 vss 1.03fF $ **FLOATING
C2175 vp_p.n615 vss 1.03fF $ **FLOATING
C2176 vp_p.n617 vss 1.03fF $ **FLOATING
C2177 vp_p.n619 vss 1.03fF $ **FLOATING
C2178 vp_p.n621 vss 1.03fF $ **FLOATING
C2179 vp_p.n623 vss 1.03fF $ **FLOATING
C2180 vp_p.n625 vss 1.03fF $ **FLOATING
C2181 vp_p.n627 vss 1.03fF $ **FLOATING
C2182 vp_p.n629 vss 1.03fF $ **FLOATING
C2183 vp_p.n631 vss 1.03fF $ **FLOATING
C2184 vp_p.n633 vss 1.03fF $ **FLOATING
C2185 vp_p.n635 vss 1.03fF $ **FLOATING
C2186 vp_p.n637 vss 1.03fF $ **FLOATING
C2187 vp_p.n639 vss 1.03fF $ **FLOATING
C2188 vp_p.n641 vss 1.03fF $ **FLOATING
C2189 vp_p.n643 vss 1.03fF $ **FLOATING
C2190 vp_p.n645 vss 1.03fF $ **FLOATING
C2191 vp_p.n647 vss 1.03fF $ **FLOATING
C2192 vp_p.n649 vss 1.03fF $ **FLOATING
C2193 vp_p.n651 vss 1.03fF $ **FLOATING
C2194 vp_p.n653 vss 1.03fF $ **FLOATING
C2195 vp_p.n655 vss 1.03fF $ **FLOATING
C2196 vp_p.n657 vss 1.03fF $ **FLOATING
C2197 vp_p.n659 vss 1.03fF $ **FLOATING
C2198 vp_p.n661 vss 1.03fF $ **FLOATING
C2199 vp_p.n663 vss 1.03fF $ **FLOATING
C2200 vp_p.n665 vss 1.03fF $ **FLOATING
C2201 vp_p.n667 vss 1.03fF $ **FLOATING
C2202 vp_p.n670 vss 1.10fF $ **FLOATING
C2203 vp_p.n743 vss 1.92fF $ **FLOATING
C2204 vp_p.n744 vss 18.53fF $ **FLOATING
C2205 vp_p.n745 vss 13.44fF $ **FLOATING
C2206 vp_p.n746 vss 13.65fF $ **FLOATING
C2207 vp_p.n747 vss 13.09fF $ **FLOATING
C2208 vp_p.n748 vss 7.69fF $ **FLOATING
C2209 vp_p.n749 vss 1.05fF $ **FLOATING
C2210 vp_p.n825 vss 1.09fF $ **FLOATING
C2211 vp_p.n827 vss 1.03fF $ **FLOATING
C2212 vp_p.n829 vss 1.03fF $ **FLOATING
C2213 vp_p.n831 vss 1.03fF $ **FLOATING
C2214 vp_p.n833 vss 1.03fF $ **FLOATING
C2215 vp_p.n835 vss 1.03fF $ **FLOATING
C2216 vp_p.n837 vss 1.03fF $ **FLOATING
C2217 vp_p.n839 vss 1.03fF $ **FLOATING
C2218 vp_p.n841 vss 1.03fF $ **FLOATING
C2219 vp_p.n843 vss 1.03fF $ **FLOATING
C2220 vp_p.n845 vss 1.03fF $ **FLOATING
C2221 vp_p.n847 vss 1.03fF $ **FLOATING
C2222 vp_p.n849 vss 1.03fF $ **FLOATING
C2223 vp_p.n851 vss 1.03fF $ **FLOATING
C2224 vp_p.n853 vss 1.03fF $ **FLOATING
C2225 vp_p.n855 vss 1.03fF $ **FLOATING
C2226 vp_p.n857 vss 1.03fF $ **FLOATING
C2227 vp_p.n859 vss 1.03fF $ **FLOATING
C2228 vp_p.n861 vss 1.03fF $ **FLOATING
C2229 vp_p.n863 vss 1.03fF $ **FLOATING
C2230 vp_p.n865 vss 1.03fF $ **FLOATING
C2231 vp_p.n867 vss 1.03fF $ **FLOATING
C2232 vp_p.n869 vss 1.03fF $ **FLOATING
C2233 vp_p.n871 vss 1.03fF $ **FLOATING
C2234 vp_p.n873 vss 1.03fF $ **FLOATING
C2235 vp_p.n875 vss 1.03fF $ **FLOATING
C2236 vp_p.n877 vss 1.03fF $ **FLOATING
C2237 vp_p.n879 vss 1.03fF $ **FLOATING
C2238 vp_p.n881 vss 1.03fF $ **FLOATING
C2239 vp_p.n883 vss 1.03fF $ **FLOATING
C2240 vp_p.n885 vss 1.03fF $ **FLOATING
C2241 vp_p.n887 vss 1.03fF $ **FLOATING
C2242 vp_p.n889 vss 1.03fF $ **FLOATING
C2243 vp_p.n891 vss 1.03fF $ **FLOATING
C2244 vp_p.n893 vss 1.03fF $ **FLOATING
C2245 vp_p.n895 vss 1.03fF $ **FLOATING
C2246 vp_p.n897 vss 1.03fF $ **FLOATING
C2247 vp_p.n899 vss 1.03fF $ **FLOATING
C2248 vp_p.n901 vss 1.03fF $ **FLOATING
C2249 vp_p.n903 vss 1.03fF $ **FLOATING
C2250 vp_p.n905 vss 1.03fF $ **FLOATING
C2251 vp_p.n907 vss 1.03fF $ **FLOATING
C2252 vp_p.n909 vss 1.03fF $ **FLOATING
C2253 vp_p.n911 vss 1.03fF $ **FLOATING
C2254 vp_p.n913 vss 1.03fF $ **FLOATING
C2255 vp_p.n915 vss 1.03fF $ **FLOATING
C2256 vp_p.n917 vss 1.03fF $ **FLOATING
C2257 vp_p.n919 vss 1.03fF $ **FLOATING
C2258 vp_p.n921 vss 1.03fF $ **FLOATING
C2259 vp_p.n923 vss 1.03fF $ **FLOATING
C2260 vp_p.n925 vss 1.03fF $ **FLOATING
C2261 vp_p.n927 vss 1.03fF $ **FLOATING
C2262 vp_p.n929 vss 1.03fF $ **FLOATING
C2263 vp_p.n931 vss 1.03fF $ **FLOATING
C2264 vp_p.n933 vss 1.03fF $ **FLOATING
C2265 vp_p.n935 vss 1.03fF $ **FLOATING
C2266 vp_p.n937 vss 1.03fF $ **FLOATING
C2267 vp_p.n939 vss 1.03fF $ **FLOATING
C2268 vp_p.n941 vss 1.03fF $ **FLOATING
C2269 vp_p.n943 vss 1.03fF $ **FLOATING
C2270 vp_p.n945 vss 1.03fF $ **FLOATING
C2271 vp_p.n947 vss 1.03fF $ **FLOATING
C2272 vp_p.n949 vss 1.03fF $ **FLOATING
C2273 vp_p.n951 vss 1.03fF $ **FLOATING
C2274 vp_p.n953 vss 1.03fF $ **FLOATING
C2275 vp_p.n955 vss 1.03fF $ **FLOATING
C2276 vp_p.n957 vss 1.03fF $ **FLOATING
C2277 vp_p.n959 vss 1.03fF $ **FLOATING
C2278 vp_p.n961 vss 1.03fF $ **FLOATING
C2279 vp_p.n963 vss 1.03fF $ **FLOATING
C2280 vp_p.n965 vss 1.03fF $ **FLOATING
C2281 vp_p.n967 vss 1.03fF $ **FLOATING
C2282 vp_p.n969 vss 1.03fF $ **FLOATING
C2283 vp_p.n974 vss 1.09fF $ **FLOATING
C2284 vp_p.n976 vss 1.03fF $ **FLOATING
C2285 vp_p.n978 vss 1.03fF $ **FLOATING
C2286 vp_p.n980 vss 1.03fF $ **FLOATING
C2287 vp_p.n982 vss 1.03fF $ **FLOATING
C2288 vp_p.n984 vss 1.03fF $ **FLOATING
C2289 vp_p.n986 vss 1.03fF $ **FLOATING
C2290 vp_p.n988 vss 1.03fF $ **FLOATING
C2291 vp_p.n990 vss 1.03fF $ **FLOATING
C2292 vp_p.n992 vss 1.03fF $ **FLOATING
C2293 vp_p.n994 vss 1.03fF $ **FLOATING
C2294 vp_p.n996 vss 1.03fF $ **FLOATING
C2295 vp_p.n998 vss 1.03fF $ **FLOATING
C2296 vp_p.n1000 vss 1.03fF $ **FLOATING
C2297 vp_p.n1002 vss 1.03fF $ **FLOATING
C2298 vp_p.n1004 vss 1.03fF $ **FLOATING
C2299 vp_p.n1006 vss 1.03fF $ **FLOATING
C2300 vp_p.n1008 vss 1.03fF $ **FLOATING
C2301 vp_p.n1010 vss 1.03fF $ **FLOATING
C2302 vp_p.n1012 vss 1.03fF $ **FLOATING
C2303 vp_p.n1014 vss 1.03fF $ **FLOATING
C2304 vp_p.n1016 vss 1.03fF $ **FLOATING
C2305 vp_p.n1018 vss 1.03fF $ **FLOATING
C2306 vp_p.n1020 vss 1.03fF $ **FLOATING
C2307 vp_p.n1022 vss 1.03fF $ **FLOATING
C2308 vp_p.n1024 vss 1.03fF $ **FLOATING
C2309 vp_p.n1026 vss 1.03fF $ **FLOATING
C2310 vp_p.n1028 vss 1.03fF $ **FLOATING
C2311 vp_p.n1030 vss 1.03fF $ **FLOATING
C2312 vp_p.n1032 vss 1.03fF $ **FLOATING
C2313 vp_p.n1034 vss 1.03fF $ **FLOATING
C2314 vp_p.n1036 vss 1.03fF $ **FLOATING
C2315 vp_p.n1038 vss 1.03fF $ **FLOATING
C2316 vp_p.n1040 vss 1.03fF $ **FLOATING
C2317 vp_p.n1042 vss 1.03fF $ **FLOATING
C2318 vp_p.n1044 vss 1.03fF $ **FLOATING
C2319 vp_p.n1046 vss 1.03fF $ **FLOATING
C2320 vp_p.n1048 vss 1.03fF $ **FLOATING
C2321 vp_p.n1050 vss 1.03fF $ **FLOATING
C2322 vp_p.n1052 vss 1.03fF $ **FLOATING
C2323 vp_p.n1054 vss 1.03fF $ **FLOATING
C2324 vp_p.n1056 vss 1.03fF $ **FLOATING
C2325 vp_p.n1058 vss 1.03fF $ **FLOATING
C2326 vp_p.n1060 vss 1.03fF $ **FLOATING
C2327 vp_p.n1062 vss 1.03fF $ **FLOATING
C2328 vp_p.n1064 vss 1.03fF $ **FLOATING
C2329 vp_p.n1066 vss 1.03fF $ **FLOATING
C2330 vp_p.n1068 vss 1.03fF $ **FLOATING
C2331 vp_p.n1070 vss 1.03fF $ **FLOATING
C2332 vp_p.n1072 vss 1.03fF $ **FLOATING
C2333 vp_p.n1074 vss 1.03fF $ **FLOATING
C2334 vp_p.n1076 vss 1.03fF $ **FLOATING
C2335 vp_p.n1078 vss 1.03fF $ **FLOATING
C2336 vp_p.n1080 vss 1.03fF $ **FLOATING
C2337 vp_p.n1082 vss 1.03fF $ **FLOATING
C2338 vp_p.n1084 vss 1.03fF $ **FLOATING
C2339 vp_p.n1086 vss 1.03fF $ **FLOATING
C2340 vp_p.n1088 vss 1.03fF $ **FLOATING
C2341 vp_p.n1090 vss 1.03fF $ **FLOATING
C2342 vp_p.n1092 vss 1.03fF $ **FLOATING
C2343 vp_p.n1094 vss 1.03fF $ **FLOATING
C2344 vp_p.n1096 vss 1.03fF $ **FLOATING
C2345 vp_p.n1098 vss 1.03fF $ **FLOATING
C2346 vp_p.n1100 vss 1.03fF $ **FLOATING
C2347 vp_p.n1102 vss 1.03fF $ **FLOATING
C2348 vp_p.n1104 vss 1.03fF $ **FLOATING
C2349 vp_p.n1106 vss 1.03fF $ **FLOATING
C2350 vp_p.n1108 vss 1.03fF $ **FLOATING
C2351 vp_p.n1110 vss 1.03fF $ **FLOATING
C2352 vp_p.n1112 vss 1.03fF $ **FLOATING
C2353 vp_p.n1114 vss 1.03fF $ **FLOATING
C2354 vp_p.n1116 vss 1.03fF $ **FLOATING
C2355 vp_p.n1118 vss 1.03fF $ **FLOATING
C2356 vp_p.n1123 vss 1.09fF $ **FLOATING
C2357 vp_p.n1125 vss 1.03fF $ **FLOATING
C2358 vp_p.n1127 vss 1.03fF $ **FLOATING
C2359 vp_p.n1129 vss 1.03fF $ **FLOATING
C2360 vp_p.n1131 vss 1.03fF $ **FLOATING
C2361 vp_p.n1133 vss 1.03fF $ **FLOATING
C2362 vp_p.n1135 vss 1.03fF $ **FLOATING
C2363 vp_p.n1137 vss 1.03fF $ **FLOATING
C2364 vp_p.n1139 vss 1.03fF $ **FLOATING
C2365 vp_p.n1141 vss 1.03fF $ **FLOATING
C2366 vp_p.n1143 vss 1.03fF $ **FLOATING
C2367 vp_p.n1145 vss 1.03fF $ **FLOATING
C2368 vp_p.n1147 vss 1.03fF $ **FLOATING
C2369 vp_p.n1149 vss 1.03fF $ **FLOATING
C2370 vp_p.n1151 vss 1.03fF $ **FLOATING
C2371 vp_p.n1153 vss 1.03fF $ **FLOATING
C2372 vp_p.n1155 vss 1.03fF $ **FLOATING
C2373 vp_p.n1157 vss 1.03fF $ **FLOATING
C2374 vp_p.n1159 vss 1.03fF $ **FLOATING
C2375 vp_p.n1161 vss 1.03fF $ **FLOATING
C2376 vp_p.n1163 vss 1.03fF $ **FLOATING
C2377 vp_p.n1165 vss 1.03fF $ **FLOATING
C2378 vp_p.n1167 vss 1.03fF $ **FLOATING
C2379 vp_p.n1169 vss 1.03fF $ **FLOATING
C2380 vp_p.n1171 vss 1.03fF $ **FLOATING
C2381 vp_p.n1173 vss 1.03fF $ **FLOATING
C2382 vp_p.n1175 vss 1.03fF $ **FLOATING
C2383 vp_p.n1177 vss 1.03fF $ **FLOATING
C2384 vp_p.n1179 vss 1.03fF $ **FLOATING
C2385 vp_p.n1181 vss 1.03fF $ **FLOATING
C2386 vp_p.n1183 vss 1.03fF $ **FLOATING
C2387 vp_p.n1185 vss 1.03fF $ **FLOATING
C2388 vp_p.n1187 vss 1.03fF $ **FLOATING
C2389 vp_p.n1189 vss 1.03fF $ **FLOATING
C2390 vp_p.n1191 vss 1.03fF $ **FLOATING
C2391 vp_p.n1193 vss 1.03fF $ **FLOATING
C2392 vp_p.n1195 vss 1.03fF $ **FLOATING
C2393 vp_p.n1197 vss 1.03fF $ **FLOATING
C2394 vp_p.n1199 vss 1.03fF $ **FLOATING
C2395 vp_p.n1201 vss 1.03fF $ **FLOATING
C2396 vp_p.n1203 vss 1.03fF $ **FLOATING
C2397 vp_p.n1205 vss 1.03fF $ **FLOATING
C2398 vp_p.n1207 vss 1.03fF $ **FLOATING
C2399 vp_p.n1209 vss 1.03fF $ **FLOATING
C2400 vp_p.n1211 vss 1.03fF $ **FLOATING
C2401 vp_p.n1213 vss 1.03fF $ **FLOATING
C2402 vp_p.n1215 vss 1.03fF $ **FLOATING
C2403 vp_p.n1217 vss 1.03fF $ **FLOATING
C2404 vp_p.n1219 vss 1.03fF $ **FLOATING
C2405 vp_p.n1221 vss 1.03fF $ **FLOATING
C2406 vp_p.n1223 vss 1.03fF $ **FLOATING
C2407 vp_p.n1225 vss 1.03fF $ **FLOATING
C2408 vp_p.n1227 vss 1.03fF $ **FLOATING
C2409 vp_p.n1229 vss 1.03fF $ **FLOATING
C2410 vp_p.n1231 vss 1.03fF $ **FLOATING
C2411 vp_p.n1233 vss 1.03fF $ **FLOATING
C2412 vp_p.n1235 vss 1.03fF $ **FLOATING
C2413 vp_p.n1237 vss 1.03fF $ **FLOATING
C2414 vp_p.n1239 vss 1.03fF $ **FLOATING
C2415 vp_p.n1241 vss 1.03fF $ **FLOATING
C2416 vp_p.n1243 vss 1.03fF $ **FLOATING
C2417 vp_p.n1245 vss 1.03fF $ **FLOATING
C2418 vp_p.n1247 vss 1.03fF $ **FLOATING
C2419 vp_p.n1249 vss 1.03fF $ **FLOATING
C2420 vp_p.n1251 vss 1.03fF $ **FLOATING
C2421 vp_p.n1253 vss 1.03fF $ **FLOATING
C2422 vp_p.n1255 vss 1.03fF $ **FLOATING
C2423 vp_p.n1257 vss 1.03fF $ **FLOATING
C2424 vp_p.n1259 vss 1.03fF $ **FLOATING
C2425 vp_p.n1261 vss 1.03fF $ **FLOATING
C2426 vp_p.n1263 vss 1.03fF $ **FLOATING
C2427 vp_p.n1265 vss 1.03fF $ **FLOATING
C2428 vp_p.n1267 vss 1.03fF $ **FLOATING
C2429 vp_p.n1272 vss 1.09fF $ **FLOATING
C2430 vp_p.n1274 vss 1.03fF $ **FLOATING
C2431 vp_p.n1276 vss 1.03fF $ **FLOATING
C2432 vp_p.n1278 vss 1.03fF $ **FLOATING
C2433 vp_p.n1280 vss 1.03fF $ **FLOATING
C2434 vp_p.n1282 vss 1.03fF $ **FLOATING
C2435 vp_p.n1284 vss 1.03fF $ **FLOATING
C2436 vp_p.n1286 vss 1.03fF $ **FLOATING
C2437 vp_p.n1288 vss 1.03fF $ **FLOATING
C2438 vp_p.n1290 vss 1.03fF $ **FLOATING
C2439 vp_p.n1292 vss 1.03fF $ **FLOATING
C2440 vp_p.n1294 vss 1.03fF $ **FLOATING
C2441 vp_p.n1296 vss 1.03fF $ **FLOATING
C2442 vp_p.n1298 vss 1.03fF $ **FLOATING
C2443 vp_p.n1300 vss 1.03fF $ **FLOATING
C2444 vp_p.n1302 vss 1.03fF $ **FLOATING
C2445 vp_p.n1304 vss 1.03fF $ **FLOATING
C2446 vp_p.n1306 vss 1.03fF $ **FLOATING
C2447 vp_p.n1308 vss 1.03fF $ **FLOATING
C2448 vp_p.n1310 vss 1.03fF $ **FLOATING
C2449 vp_p.n1312 vss 1.03fF $ **FLOATING
C2450 vp_p.n1314 vss 1.03fF $ **FLOATING
C2451 vp_p.n1316 vss 1.03fF $ **FLOATING
C2452 vp_p.n1318 vss 1.03fF $ **FLOATING
C2453 vp_p.n1320 vss 1.03fF $ **FLOATING
C2454 vp_p.n1322 vss 1.03fF $ **FLOATING
C2455 vp_p.n1324 vss 1.03fF $ **FLOATING
C2456 vp_p.n1326 vss 1.03fF $ **FLOATING
C2457 vp_p.n1328 vss 1.03fF $ **FLOATING
C2458 vp_p.n1330 vss 1.03fF $ **FLOATING
C2459 vp_p.n1332 vss 1.03fF $ **FLOATING
C2460 vp_p.n1334 vss 1.03fF $ **FLOATING
C2461 vp_p.n1336 vss 1.03fF $ **FLOATING
C2462 vp_p.n1338 vss 1.03fF $ **FLOATING
C2463 vp_p.n1340 vss 1.03fF $ **FLOATING
C2464 vp_p.n1342 vss 1.03fF $ **FLOATING
C2465 vp_p.n1344 vss 1.03fF $ **FLOATING
C2466 vp_p.n1346 vss 1.03fF $ **FLOATING
C2467 vp_p.n1348 vss 1.03fF $ **FLOATING
C2468 vp_p.n1350 vss 1.03fF $ **FLOATING
C2469 vp_p.n1352 vss 1.03fF $ **FLOATING
C2470 vp_p.n1354 vss 1.03fF $ **FLOATING
C2471 vp_p.n1356 vss 1.03fF $ **FLOATING
C2472 vp_p.n1358 vss 1.03fF $ **FLOATING
C2473 vp_p.n1360 vss 1.03fF $ **FLOATING
C2474 vp_p.n1362 vss 1.03fF $ **FLOATING
C2475 vp_p.n1364 vss 1.03fF $ **FLOATING
C2476 vp_p.n1366 vss 1.03fF $ **FLOATING
C2477 vp_p.n1368 vss 1.03fF $ **FLOATING
C2478 vp_p.n1370 vss 1.03fF $ **FLOATING
C2479 vp_p.n1372 vss 1.03fF $ **FLOATING
C2480 vp_p.n1374 vss 1.03fF $ **FLOATING
C2481 vp_p.n1376 vss 1.03fF $ **FLOATING
C2482 vp_p.n1378 vss 1.03fF $ **FLOATING
C2483 vp_p.n1380 vss 1.03fF $ **FLOATING
C2484 vp_p.n1382 vss 1.03fF $ **FLOATING
C2485 vp_p.n1384 vss 1.03fF $ **FLOATING
C2486 vp_p.n1386 vss 1.03fF $ **FLOATING
C2487 vp_p.n1388 vss 1.03fF $ **FLOATING
C2488 vp_p.n1390 vss 1.03fF $ **FLOATING
C2489 vp_p.n1392 vss 1.03fF $ **FLOATING
C2490 vp_p.n1394 vss 1.03fF $ **FLOATING
C2491 vp_p.n1396 vss 1.03fF $ **FLOATING
C2492 vp_p.n1398 vss 1.03fF $ **FLOATING
C2493 vp_p.n1400 vss 1.03fF $ **FLOATING
C2494 vp_p.n1402 vss 1.03fF $ **FLOATING
C2495 vp_p.n1404 vss 1.03fF $ **FLOATING
C2496 vp_p.n1406 vss 1.03fF $ **FLOATING
C2497 vp_p.n1408 vss 1.03fF $ **FLOATING
C2498 vp_p.n1410 vss 1.03fF $ **FLOATING
C2499 vp_p.n1412 vss 1.03fF $ **FLOATING
C2500 vp_p.n1414 vss 1.03fF $ **FLOATING
C2501 vp_p.n1416 vss 1.03fF $ **FLOATING
C2502 vp_p.n1419 vss 1.04fF $ **FLOATING
C2503 vp_p.n1492 vss 1.34fF $ **FLOATING
C2504 vp_p.n1493 vss 19.04fF $ **FLOATING
C2505 vp_p.n1494 vss 13.65fF $ **FLOATING
C2506 vp_p.n1495 vss 13.44fF $ **FLOATING
C2507 vp_p.n1496 vss 13.30fF $ **FLOATING
C2508 vp_p.n1497 vss 6.61fF $ **FLOATING
.ends
