magic
tech sky130A
magscale 1 2
timestamp 1628437795
<< nwell >>
rect -596 2790 -482 2850
rect -596 2590 -474 2790
rect -596 2288 -482 2590
<< pwell >>
rect -622 1922 -278 2152
<< psubdiffcont >>
rect -574 1966 -510 2108
<< nsubdiffcont >>
rect -550 2620 -510 2736
<< poly >>
rect -416 2220 -350 2296
<< locali >>
rect -570 2736 -492 2756
rect -570 2620 -550 2736
rect -510 2620 -492 2736
rect -570 2600 -492 2620
rect -592 2108 -494 2124
rect -592 1966 -574 2108
rect -510 1966 -494 2108
rect -592 1950 -494 1966
<< viali >>
rect -550 2620 -510 2736
rect -400 2170 -366 2342
rect -574 1966 -510 2108
<< metal1 >>
rect -466 2892 -456 2918
rect -556 2854 -456 2892
rect -556 2736 -494 2854
rect -466 2852 -456 2854
rect -392 2852 -382 2918
rect -450 2788 -404 2852
rect -556 2620 -550 2736
rect -510 2620 -494 2736
rect -556 2608 -494 2620
rect -316 2388 -280 2416
rect -406 2342 -360 2354
rect -406 2302 -400 2342
rect -412 2278 -400 2302
rect -492 2232 -400 2278
rect -412 2210 -400 2232
rect -406 2170 -400 2210
rect -366 2170 -360 2342
rect -406 2164 -360 2170
rect -310 2132 -280 2388
rect -580 2108 -504 2120
rect -580 1966 -574 2108
rect -510 1966 -504 2108
rect -316 2092 -280 2132
rect -580 1954 -504 1966
rect -556 1898 -512 1954
rect -450 1898 -404 1932
rect -556 1884 -404 1898
rect -556 1840 -458 1884
rect -468 1820 -458 1840
rect -394 1820 -384 1884
<< via1 >>
rect -456 2852 -392 2918
rect -458 1820 -394 1884
<< metal2 >>
rect -462 2924 -380 2934
rect -462 2830 -380 2840
rect -462 1892 -386 1902
rect -462 1806 -386 1816
<< via2 >>
rect -462 2918 -380 2924
rect -462 2852 -456 2918
rect -456 2852 -392 2918
rect -392 2852 -380 2918
rect -462 2840 -380 2852
rect -462 1884 -386 1892
rect -462 1820 -458 1884
rect -458 1820 -394 1884
rect -394 1820 -386 1884
rect -462 1816 -386 1820
<< metal3 >>
rect -472 2926 -370 2930
rect -472 2834 -462 2926
rect -380 2834 -370 2926
rect -474 1898 -372 1904
rect -476 1810 -466 1898
rect -378 1810 -368 1898
rect -474 1804 -372 1810
<< via3 >>
rect -462 2924 -380 2926
rect -462 2840 -380 2924
rect -462 2834 -380 2840
rect -466 1892 -378 1898
rect -466 1816 -462 1892
rect -462 1816 -386 1892
rect -386 1816 -378 1892
rect -466 1810 -378 1816
<< metal4 >>
rect -466 2926 -296 2930
rect -466 2834 -462 2926
rect -380 2834 -296 2926
rect -466 2830 -296 2834
rect -470 1898 -300 1904
rect -470 1810 -466 1898
rect -378 1810 -300 1898
rect -470 1804 -300 1810
use sky130_fd_pr__pfet_01v8_L4T9AL  sky130_fd_pr__pfet_01v8_L4T9AL_0
timestamp 1627366162
transform 1 0 -383 0 1 2552
box -109 -264 109 298
use sky130_fd_pr__nfet_01v8_UPT43B  sky130_fd_pr__nfet_01v8_UPT43B_0
timestamp 1627366162
transform 1 0 -383 0 1 2063
box -73 -157 73 157
<< labels >>
flabel metal4 -328 2880 -328 2880 0 FreeSans 1600 0 0 0 vdd
port 0 nsew
flabel metal1 -472 2252 -472 2252 0 FreeSans 1600 0 0 0 A
port 1 nsew
flabel metal1 -296 2230 -296 2230 0 FreeSans 1600 0 0 0 B
port 2 nsew
flabel metal4 -330 1812 -330 1812 0 FreeSans 1600 0 0 0 vss
port 3 nsew
<< end >>
