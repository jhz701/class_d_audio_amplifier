magic
tech sky130A
magscale 1 2
timestamp 1627297958
<< pwell >>
rect 1990 9144 2062 9308
<< locali >>
rect 1288 6670 1862 6896
rect 1336 2830 1862 3050
<< viali >>
rect 820 6560 1288 6976
rect 868 2744 1336 3160
<< metal1 >>
rect 2100 28464 3236 29310
rect 2100 22838 2398 28464
rect 28940 28458 30158 28980
rect 3986 25552 4258 25668
rect 2006 21990 2016 22838
rect 2838 21990 2848 22838
rect 32286 22252 32296 23036
rect 33112 22252 33122 23036
rect 1990 12038 3234 12908
rect 29302 12124 29882 12646
rect 1990 9144 2062 12038
rect 4006 9148 4252 9264
rect 808 6976 1300 6982
rect 808 6560 820 6976
rect 1288 6560 1300 6976
rect 808 6554 1300 6560
rect 1990 5980 2062 6536
rect 1970 5454 1980 5980
rect 2496 5454 2506 5980
rect 1990 4980 2062 5454
rect 856 3160 1348 3166
rect 856 2744 868 3160
rect 1336 2744 1348 3160
rect 856 2738 1348 2744
rect 32302 2486 32762 22252
rect 1990 2122 2062 2314
rect 1980 1572 1990 2122
rect 2534 1572 2544 2122
rect 32190 1618 32200 2486
rect 33018 1618 33028 2486
<< via1 >>
rect 2016 21990 2838 22838
rect 32296 22252 33112 23036
rect 820 6560 1288 6976
rect 1980 5454 2496 5980
rect 868 2744 1336 3160
rect 1990 1572 2534 2122
rect 32200 1618 33018 2486
<< metal2 >>
rect 32296 23036 33112 23046
rect 2016 22838 2838 22848
rect 2838 22068 15808 22600
rect 18912 22258 32296 22700
rect 32296 22242 33112 22252
rect 2016 21980 2838 21990
rect 820 6976 1288 6986
rect 820 6550 1288 6560
rect 1980 5980 2496 5990
rect 2496 5524 15814 5912
rect 1980 5444 2496 5454
rect 18908 4870 19408 5364
rect 868 3160 1336 3170
rect 868 2734 1336 2744
rect 32200 2486 33018 2496
rect 1990 2122 2534 2132
rect 2534 1620 32200 2062
rect 32200 1608 33018 1618
rect 1990 1562 2534 1572
<< via2 >>
rect 820 6560 1288 6976
rect 868 2744 1336 3160
<< metal3 >>
rect 810 6976 1298 6981
rect 810 6560 820 6976
rect 1288 6560 1298 6976
rect 810 6555 1298 6560
rect 858 3160 1346 3165
rect 858 2744 868 3160
rect 1336 2744 1346 3160
rect 858 2739 1346 2744
<< via3 >>
rect 820 6560 1288 6976
rect 868 2744 1336 3160
<< metal4 >>
rect 32064 23692 35064 25224
rect -2 16322 28546 16504
rect 33850 8822 35064 23692
rect 32064 7290 35064 8822
rect 819 6976 1289 6977
rect 819 6560 820 6976
rect 1288 6560 1289 6976
rect 819 6559 1289 6560
rect 867 3160 1337 3161
rect 867 2744 868 3160
rect 1336 2744 1337 3160
rect 867 2743 1337 2744
use OTA  OTA_0 ~/magic/class_d_audio_amplifier/OTA
timestamp 1627028181
transform 1 0 19206 0 1 19408
box -19208 -19408 12858 -3006
use OTA  OTA_1
timestamp 1627028181
transform 1 0 19206 0 1 35810
box -19208 -19408 12858 -3006
use sky130_fd_pr__res_xhigh_po_0p35_X24WYH  sky130_fd_pr__res_xhigh_po_0p35_X24WYH_0
timestamp 1627296012
transform 1 0 2026 0 1 3709
box -201 -1598 201 1598
use sky130_fd_pr__res_xhigh_po_0p35_X24WYH  sky130_fd_pr__res_xhigh_po_0p35_X24WYH_1
timestamp 1627296012
transform 1 0 2026 0 1 7743
box -201 -1598 201 1598
<< labels >>
flabel metal2 19304 5158 19304 5158 0 FreeSans 3200 0 0 0 vref
port 4 nsew
flabel metal1 32464 14304 32464 14304 0 FreeSans 3200 0 0 0 vi
port 3 nsew
flabel metal1 4088 25610 4088 25610 0 FreeSans 3200 0 0 0 vbias1
port 1 nsew
flabel metal1 4066 9202 4066 9202 0 FreeSans 3200 0 0 0 vbias2
port 2 nsew
flabel metal4 2570 16386 2570 16386 0 FreeSans 3200 0 0 0 vss
port 5 nsew
flabel metal4 34766 13506 34766 13506 0 FreeSans 3200 0 0 0 vdd
port 0 nsew
flabel metal1 29396 28690 29396 28690 0 FreeSans 3200 0 0 0 vp
port 7 nsew
flabel metal1 29618 12410 29618 12410 0 FreeSans 3200 0 0 0 vn
port 6 nsew
<< end >>
