magic
tech sky130A
magscale 1 2
timestamp 1632368578
<< nwell >>
rect 61629 13567 91905 43843
<< pwell >>
rect 61491 43843 92043 43981
rect 61491 13567 61629 43843
rect 91905 13567 92043 43843
rect 61491 13429 92043 13567
rect 61637 -30343 91913 -67
<< psubdiff >>
rect 61527 43911 61623 43945
rect 91911 43911 92007 43945
rect 61527 43849 61561 43911
rect 91973 43849 92007 43911
rect 61527 13499 61561 13561
rect 91973 13499 92007 13561
rect 61527 13465 61623 13499
rect 91911 13465 92007 13499
rect 61673 -137 61769 -103
rect 91781 -137 91877 -103
rect 61673 -199 61707 -137
rect 91843 -199 91877 -137
rect 61673 -30273 61707 -30211
rect 91843 -30273 91877 -30211
rect 61673 -30307 61769 -30273
rect 91781 -30307 91877 -30273
<< nsubdiff >>
rect 61665 43773 61761 43807
rect 91773 43773 91869 43807
rect 61665 43711 61699 43773
rect 91835 43711 91869 43773
rect 61665 13637 61699 13699
rect 91835 13637 91869 13699
rect 61665 13603 61761 13637
rect 91773 13603 91869 13637
<< psubdiffcont >>
rect 61623 43911 91911 43945
rect 61527 13561 61561 43849
rect 91973 13561 92007 43849
rect 61623 13465 91911 13499
rect 61769 -137 91781 -103
rect 61673 -30211 61707 -199
rect 91843 -30211 91877 -199
rect 61769 -30307 91781 -30273
<< nsubdiffcont >>
rect 61761 43773 91773 43807
rect 61665 13699 61699 43711
rect 91835 13699 91869 43711
rect 61761 13603 91773 13637
<< pdiode >>
rect 61767 43693 91767 43705
rect 61767 13717 61779 43693
rect 91755 13717 91767 43693
rect 61767 13705 91767 13717
<< ndiode >>
rect 61775 -217 91775 -205
rect 61775 -30193 61787 -217
rect 91763 -30193 91775 -217
rect 61775 -30205 91775 -30193
<< pdiodec >>
rect 61779 13717 91755 43693
<< ndiodec >>
rect 61787 -30193 91763 -217
<< locali >>
rect 61527 43911 61623 43945
rect 91911 43911 92007 43945
rect 61527 43849 61561 43911
rect 91973 43849 92007 43911
rect 61665 43773 61761 43807
rect 91773 43773 91869 43807
rect 61665 43711 61699 43773
rect 91835 43711 91869 43773
rect 61763 13717 61779 43693
rect 91755 13717 91771 43693
rect 61665 13637 61699 13699
rect 91835 13637 91869 13699
rect 61665 13603 61761 13637
rect 91773 13603 91869 13637
rect 61527 13499 61561 13561
rect 91973 13499 92007 13561
rect 61527 13465 61623 13499
rect 91911 13465 92007 13499
rect 61673 -137 61769 -103
rect 91781 -137 91877 -103
rect 61673 -199 61707 -137
rect 91843 -199 91877 -137
rect 61771 -30193 61787 -217
rect 91763 -30193 91779 -217
rect 61673 -30273 61707 -30211
rect 91843 -30273 91877 -30211
rect 61673 -30307 61769 -30273
rect 91781 -30307 91877 -30273
<< viali >>
rect 61779 13717 91755 43693
rect 61787 -30193 91763 -217
<< metal1 >>
rect 61767 43693 91767 43699
rect 61767 13717 61779 43693
rect 91755 13850 91767 43693
rect 91755 13717 91770 13850
rect 61767 13711 91770 13717
rect 61780 -211 91770 13711
rect 61775 -217 91775 -211
rect 61775 -30193 61787 -217
rect 91763 -30193 91775 -217
rect 61775 -30199 91775 -30193
<< labels >>
flabel metal1 66220 9000 66220 9000 0 FreeSans 32000 0 0 0 vin
flabel locali 61550 13490 61550 13490 0 FreeSans 8000 0 0 0 vss
flabel nsubdiffcont 61680 14660 61680 14660 0 FreeSans 8000 0 0 0 vdd
<< end >>
