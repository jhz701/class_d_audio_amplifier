magic
tech sky130A
magscale 1 2
timestamp 1629189135
<< nwell >>
rect 18539 9687 30663 11797
rect 20027 5063 23223 9409
<< pwell >>
rect 23653 5739 24055 7495
rect 20027 2841 29175 4715
<< pmoslvt >>
rect 18735 11178 18935 11578
rect 19107 11178 19307 11578
rect 19479 11178 19679 11578
rect 19851 11178 20051 11578
rect 20223 11178 20423 11578
rect 20595 11178 20795 11578
rect 20967 11178 21167 11578
rect 21339 11178 21539 11578
rect 21711 11178 21911 11578
rect 22083 11178 22283 11578
rect 22455 11178 22655 11578
rect 22827 11178 23027 11578
rect 23199 11178 23399 11578
rect 23571 11178 23771 11578
rect 23943 11178 24143 11578
rect 24315 11178 24515 11578
rect 24687 11178 24887 11578
rect 25059 11178 25259 11578
rect 25431 11178 25631 11578
rect 25803 11178 26003 11578
rect 26175 11178 26375 11578
rect 26547 11178 26747 11578
rect 26919 11178 27119 11578
rect 27291 11178 27491 11578
rect 27663 11178 27863 11578
rect 28035 11178 28235 11578
rect 28407 11178 28607 11578
rect 28779 11178 28979 11578
rect 29151 11178 29351 11578
rect 29523 11178 29723 11578
rect 29895 11178 30095 11578
rect 30267 11178 30467 11578
rect 18735 10542 18935 10942
rect 19107 10542 19307 10942
rect 19479 10542 19679 10942
rect 19851 10542 20051 10942
rect 20223 10542 20423 10942
rect 20595 10542 20795 10942
rect 20967 10542 21167 10942
rect 21339 10542 21539 10942
rect 21711 10542 21911 10942
rect 22083 10542 22283 10942
rect 22455 10542 22655 10942
rect 22827 10542 23027 10942
rect 23199 10542 23399 10942
rect 23571 10542 23771 10942
rect 23943 10542 24143 10942
rect 24315 10542 24515 10942
rect 24687 10542 24887 10942
rect 25059 10542 25259 10942
rect 25431 10542 25631 10942
rect 25803 10542 26003 10942
rect 26175 10542 26375 10942
rect 26547 10542 26747 10942
rect 26919 10542 27119 10942
rect 27291 10542 27491 10942
rect 27663 10542 27863 10942
rect 28035 10542 28235 10942
rect 28407 10542 28607 10942
rect 28779 10542 28979 10942
rect 29151 10542 29351 10942
rect 29523 10542 29723 10942
rect 29895 10542 30095 10942
rect 30267 10542 30467 10942
rect 18735 9906 18935 10306
rect 19107 9906 19307 10306
rect 19479 9906 19679 10306
rect 19851 9906 20051 10306
rect 20223 9906 20423 10306
rect 20595 9906 20795 10306
rect 20967 9906 21167 10306
rect 21339 9906 21539 10306
rect 21711 9906 21911 10306
rect 22083 9906 22283 10306
rect 22455 9906 22655 10306
rect 22827 9906 23027 10306
rect 23199 9906 23399 10306
rect 23571 9906 23771 10306
rect 23943 9906 24143 10306
rect 24315 9906 24515 10306
rect 24687 9906 24887 10306
rect 25059 9906 25259 10306
rect 25431 9906 25631 10306
rect 25803 9906 26003 10306
rect 26175 9906 26375 10306
rect 26547 9906 26747 10306
rect 26919 9906 27119 10306
rect 27291 9906 27491 10306
rect 27663 9906 27863 10306
rect 28035 9906 28235 10306
rect 28407 9906 28607 10306
rect 28779 9906 28979 10306
rect 29151 9906 29351 10306
rect 29523 9906 29723 10306
rect 29895 9906 30095 10306
rect 30267 9906 30467 10306
rect 20223 8390 20423 9190
rect 20595 8390 20795 9190
rect 20967 8390 21167 9190
rect 21339 8390 21539 9190
rect 21711 8390 21911 9190
rect 22083 8390 22283 9190
rect 22455 8390 22655 9190
rect 22827 8390 23027 9190
rect 20223 7354 20423 8154
rect 20595 7354 20795 8154
rect 20967 7354 21167 8154
rect 21339 7354 21539 8154
rect 21711 7354 21911 8154
rect 22083 7354 22283 8154
rect 22455 7354 22655 8154
rect 22827 7354 23027 8154
rect 20223 6318 20423 7118
rect 20595 6318 20795 7118
rect 20967 6318 21167 7118
rect 21339 6318 21539 7118
rect 21711 6318 21911 7118
rect 22083 6318 22283 7118
rect 22455 6318 22655 7118
rect 22827 6318 23027 7118
rect 20223 5282 20423 6082
rect 20595 5282 20795 6082
rect 20967 5282 21167 6082
rect 21339 5282 21539 6082
rect 21711 5282 21911 6082
rect 22083 5282 22283 6082
rect 22455 5282 22655 6082
rect 22827 5282 23027 6082
<< nmoslvt >>
rect 20223 4305 20423 4505
rect 20595 4305 20795 4505
rect 20967 4305 21167 4505
rect 21339 4305 21539 4505
rect 21711 4305 21911 4505
rect 22083 4305 22283 4505
rect 22455 4305 22655 4505
rect 22827 4305 23027 4505
rect 23199 4305 23399 4505
rect 23571 4305 23771 4505
rect 23943 4305 24143 4505
rect 24315 4305 24515 4505
rect 24687 4305 24887 4505
rect 25059 4305 25259 4505
rect 25431 4305 25631 4505
rect 25803 4305 26003 4505
rect 26175 4305 26375 4505
rect 26547 4305 26747 4505
rect 26919 4305 27119 4505
rect 27291 4305 27491 4505
rect 27663 4305 27863 4505
rect 28035 4305 28235 4505
rect 28407 4305 28607 4505
rect 28779 4305 28979 4505
rect 20223 3887 20423 4087
rect 20595 3887 20795 4087
rect 20967 3887 21167 4087
rect 21339 3887 21539 4087
rect 21711 3887 21911 4087
rect 22083 3887 22283 4087
rect 22455 3887 22655 4087
rect 22827 3887 23027 4087
rect 23199 3887 23399 4087
rect 23571 3887 23771 4087
rect 23943 3887 24143 4087
rect 24315 3887 24515 4087
rect 24687 3887 24887 4087
rect 25059 3887 25259 4087
rect 25431 3887 25631 4087
rect 25803 3887 26003 4087
rect 26175 3887 26375 4087
rect 26547 3887 26747 4087
rect 26919 3887 27119 4087
rect 27291 3887 27491 4087
rect 27663 3887 27863 4087
rect 28035 3887 28235 4087
rect 28407 3887 28607 4087
rect 28779 3887 28979 4087
rect 20223 3469 20423 3669
rect 20595 3469 20795 3669
rect 20967 3469 21167 3669
rect 21339 3469 21539 3669
rect 21711 3469 21911 3669
rect 22083 3469 22283 3669
rect 22455 3469 22655 3669
rect 22827 3469 23027 3669
rect 23199 3469 23399 3669
rect 23571 3469 23771 3669
rect 23943 3469 24143 3669
rect 24315 3469 24515 3669
rect 24687 3469 24887 3669
rect 25059 3469 25259 3669
rect 25431 3469 25631 3669
rect 25803 3469 26003 3669
rect 26175 3469 26375 3669
rect 26547 3469 26747 3669
rect 26919 3469 27119 3669
rect 27291 3469 27491 3669
rect 27663 3469 27863 3669
rect 28035 3469 28235 3669
rect 28407 3469 28607 3669
rect 28779 3469 28979 3669
rect 20223 3051 20423 3251
rect 20595 3051 20795 3251
rect 20967 3051 21167 3251
rect 21339 3051 21539 3251
rect 21711 3051 21911 3251
rect 22083 3051 22283 3251
rect 22455 3051 22655 3251
rect 22827 3051 23027 3251
rect 23199 3051 23399 3251
rect 23571 3051 23771 3251
rect 23943 3051 24143 3251
rect 24315 3051 24515 3251
rect 24687 3051 24887 3251
rect 25059 3051 25259 3251
rect 25431 3051 25631 3251
rect 25803 3051 26003 3251
rect 26175 3051 26375 3251
rect 26547 3051 26747 3251
rect 26919 3051 27119 3251
rect 27291 3051 27491 3251
rect 27663 3051 27863 3251
rect 28035 3051 28235 3251
rect 28407 3051 28607 3251
rect 28779 3051 28979 3251
<< ndiff >>
rect 20165 4493 20223 4505
rect 20165 4317 20177 4493
rect 20211 4317 20223 4493
rect 20165 4305 20223 4317
rect 20423 4493 20481 4505
rect 20423 4317 20435 4493
rect 20469 4317 20481 4493
rect 20423 4305 20481 4317
rect 20537 4493 20595 4505
rect 20537 4317 20549 4493
rect 20583 4317 20595 4493
rect 20537 4305 20595 4317
rect 20795 4493 20853 4505
rect 20795 4317 20807 4493
rect 20841 4317 20853 4493
rect 20795 4305 20853 4317
rect 20909 4493 20967 4505
rect 20909 4317 20921 4493
rect 20955 4317 20967 4493
rect 20909 4305 20967 4317
rect 21167 4493 21225 4505
rect 21167 4317 21179 4493
rect 21213 4317 21225 4493
rect 21167 4305 21225 4317
rect 21281 4493 21339 4505
rect 21281 4317 21293 4493
rect 21327 4317 21339 4493
rect 21281 4305 21339 4317
rect 21539 4493 21597 4505
rect 21539 4317 21551 4493
rect 21585 4317 21597 4493
rect 21539 4305 21597 4317
rect 21653 4493 21711 4505
rect 21653 4317 21665 4493
rect 21699 4317 21711 4493
rect 21653 4305 21711 4317
rect 21911 4493 21969 4505
rect 21911 4317 21923 4493
rect 21957 4317 21969 4493
rect 21911 4305 21969 4317
rect 22025 4493 22083 4505
rect 22025 4317 22037 4493
rect 22071 4317 22083 4493
rect 22025 4305 22083 4317
rect 22283 4493 22341 4505
rect 22283 4317 22295 4493
rect 22329 4317 22341 4493
rect 22283 4305 22341 4317
rect 22397 4493 22455 4505
rect 22397 4317 22409 4493
rect 22443 4317 22455 4493
rect 22397 4305 22455 4317
rect 22655 4493 22713 4505
rect 22655 4317 22667 4493
rect 22701 4317 22713 4493
rect 22655 4305 22713 4317
rect 22769 4493 22827 4505
rect 22769 4317 22781 4493
rect 22815 4317 22827 4493
rect 22769 4305 22827 4317
rect 23027 4493 23085 4505
rect 23027 4317 23039 4493
rect 23073 4317 23085 4493
rect 23027 4305 23085 4317
rect 23141 4493 23199 4505
rect 23141 4317 23153 4493
rect 23187 4317 23199 4493
rect 23141 4305 23199 4317
rect 23399 4493 23457 4505
rect 23399 4317 23411 4493
rect 23445 4317 23457 4493
rect 23399 4305 23457 4317
rect 23513 4493 23571 4505
rect 23513 4317 23525 4493
rect 23559 4317 23571 4493
rect 23513 4305 23571 4317
rect 23771 4493 23829 4505
rect 23771 4317 23783 4493
rect 23817 4317 23829 4493
rect 23771 4305 23829 4317
rect 23885 4493 23943 4505
rect 23885 4317 23897 4493
rect 23931 4317 23943 4493
rect 23885 4305 23943 4317
rect 24143 4493 24201 4505
rect 24143 4317 24155 4493
rect 24189 4317 24201 4493
rect 24143 4305 24201 4317
rect 24257 4493 24315 4505
rect 24257 4317 24269 4493
rect 24303 4317 24315 4493
rect 24257 4305 24315 4317
rect 24515 4493 24573 4505
rect 24515 4317 24527 4493
rect 24561 4317 24573 4493
rect 24515 4305 24573 4317
rect 24629 4493 24687 4505
rect 24629 4317 24641 4493
rect 24675 4317 24687 4493
rect 24629 4305 24687 4317
rect 24887 4493 24945 4505
rect 24887 4317 24899 4493
rect 24933 4317 24945 4493
rect 24887 4305 24945 4317
rect 25001 4493 25059 4505
rect 25001 4317 25013 4493
rect 25047 4317 25059 4493
rect 25001 4305 25059 4317
rect 25259 4493 25317 4505
rect 25259 4317 25271 4493
rect 25305 4317 25317 4493
rect 25259 4305 25317 4317
rect 25373 4493 25431 4505
rect 25373 4317 25385 4493
rect 25419 4317 25431 4493
rect 25373 4305 25431 4317
rect 25631 4493 25689 4505
rect 25631 4317 25643 4493
rect 25677 4317 25689 4493
rect 25631 4305 25689 4317
rect 25745 4493 25803 4505
rect 25745 4317 25757 4493
rect 25791 4317 25803 4493
rect 25745 4305 25803 4317
rect 26003 4493 26061 4505
rect 26003 4317 26015 4493
rect 26049 4317 26061 4493
rect 26003 4305 26061 4317
rect 26117 4493 26175 4505
rect 26117 4317 26129 4493
rect 26163 4317 26175 4493
rect 26117 4305 26175 4317
rect 26375 4493 26433 4505
rect 26375 4317 26387 4493
rect 26421 4317 26433 4493
rect 26375 4305 26433 4317
rect 26489 4493 26547 4505
rect 26489 4317 26501 4493
rect 26535 4317 26547 4493
rect 26489 4305 26547 4317
rect 26747 4493 26805 4505
rect 26747 4317 26759 4493
rect 26793 4317 26805 4493
rect 26747 4305 26805 4317
rect 26861 4493 26919 4505
rect 26861 4317 26873 4493
rect 26907 4317 26919 4493
rect 26861 4305 26919 4317
rect 27119 4493 27177 4505
rect 27119 4317 27131 4493
rect 27165 4317 27177 4493
rect 27119 4305 27177 4317
rect 27233 4493 27291 4505
rect 27233 4317 27245 4493
rect 27279 4317 27291 4493
rect 27233 4305 27291 4317
rect 27491 4493 27549 4505
rect 27491 4317 27503 4493
rect 27537 4317 27549 4493
rect 27491 4305 27549 4317
rect 27605 4493 27663 4505
rect 27605 4317 27617 4493
rect 27651 4317 27663 4493
rect 27605 4305 27663 4317
rect 27863 4493 27921 4505
rect 27863 4317 27875 4493
rect 27909 4317 27921 4493
rect 27863 4305 27921 4317
rect 27977 4493 28035 4505
rect 27977 4317 27989 4493
rect 28023 4317 28035 4493
rect 27977 4305 28035 4317
rect 28235 4493 28293 4505
rect 28235 4317 28247 4493
rect 28281 4317 28293 4493
rect 28235 4305 28293 4317
rect 28349 4493 28407 4505
rect 28349 4317 28361 4493
rect 28395 4317 28407 4493
rect 28349 4305 28407 4317
rect 28607 4493 28665 4505
rect 28607 4317 28619 4493
rect 28653 4317 28665 4493
rect 28607 4305 28665 4317
rect 28721 4493 28779 4505
rect 28721 4317 28733 4493
rect 28767 4317 28779 4493
rect 28721 4305 28779 4317
rect 28979 4493 29037 4505
rect 28979 4317 28991 4493
rect 29025 4317 29037 4493
rect 28979 4305 29037 4317
rect 20165 4075 20223 4087
rect 20165 3899 20177 4075
rect 20211 3899 20223 4075
rect 20165 3887 20223 3899
rect 20423 4075 20481 4087
rect 20423 3899 20435 4075
rect 20469 3899 20481 4075
rect 20423 3887 20481 3899
rect 20537 4075 20595 4087
rect 20537 3899 20549 4075
rect 20583 3899 20595 4075
rect 20537 3887 20595 3899
rect 20795 4075 20853 4087
rect 20795 3899 20807 4075
rect 20841 3899 20853 4075
rect 20795 3887 20853 3899
rect 20909 4075 20967 4087
rect 20909 3899 20921 4075
rect 20955 3899 20967 4075
rect 20909 3887 20967 3899
rect 21167 4075 21225 4087
rect 21167 3899 21179 4075
rect 21213 3899 21225 4075
rect 21167 3887 21225 3899
rect 21281 4075 21339 4087
rect 21281 3899 21293 4075
rect 21327 3899 21339 4075
rect 21281 3887 21339 3899
rect 21539 4075 21597 4087
rect 21539 3899 21551 4075
rect 21585 3899 21597 4075
rect 21539 3887 21597 3899
rect 21653 4075 21711 4087
rect 21653 3899 21665 4075
rect 21699 3899 21711 4075
rect 21653 3887 21711 3899
rect 21911 4075 21969 4087
rect 21911 3899 21923 4075
rect 21957 3899 21969 4075
rect 21911 3887 21969 3899
rect 22025 4075 22083 4087
rect 22025 3899 22037 4075
rect 22071 3899 22083 4075
rect 22025 3887 22083 3899
rect 22283 4075 22341 4087
rect 22283 3899 22295 4075
rect 22329 3899 22341 4075
rect 22283 3887 22341 3899
rect 22397 4075 22455 4087
rect 22397 3899 22409 4075
rect 22443 3899 22455 4075
rect 22397 3887 22455 3899
rect 22655 4075 22713 4087
rect 22655 3899 22667 4075
rect 22701 3899 22713 4075
rect 22655 3887 22713 3899
rect 22769 4075 22827 4087
rect 22769 3899 22781 4075
rect 22815 3899 22827 4075
rect 22769 3887 22827 3899
rect 23027 4075 23085 4087
rect 23027 3899 23039 4075
rect 23073 3899 23085 4075
rect 23027 3887 23085 3899
rect 23141 4075 23199 4087
rect 23141 3899 23153 4075
rect 23187 3899 23199 4075
rect 23141 3887 23199 3899
rect 23399 4075 23457 4087
rect 23399 3899 23411 4075
rect 23445 3899 23457 4075
rect 23399 3887 23457 3899
rect 23513 4075 23571 4087
rect 23513 3899 23525 4075
rect 23559 3899 23571 4075
rect 23513 3887 23571 3899
rect 23771 4075 23829 4087
rect 23771 3899 23783 4075
rect 23817 3899 23829 4075
rect 23771 3887 23829 3899
rect 23885 4075 23943 4087
rect 23885 3899 23897 4075
rect 23931 3899 23943 4075
rect 23885 3887 23943 3899
rect 24143 4075 24201 4087
rect 24143 3899 24155 4075
rect 24189 3899 24201 4075
rect 24143 3887 24201 3899
rect 24257 4075 24315 4087
rect 24257 3899 24269 4075
rect 24303 3899 24315 4075
rect 24257 3887 24315 3899
rect 24515 4075 24573 4087
rect 24515 3899 24527 4075
rect 24561 3899 24573 4075
rect 24515 3887 24573 3899
rect 24629 4075 24687 4087
rect 24629 3899 24641 4075
rect 24675 3899 24687 4075
rect 24629 3887 24687 3899
rect 24887 4075 24945 4087
rect 24887 3899 24899 4075
rect 24933 3899 24945 4075
rect 24887 3887 24945 3899
rect 25001 4075 25059 4087
rect 25001 3899 25013 4075
rect 25047 3899 25059 4075
rect 25001 3887 25059 3899
rect 25259 4075 25317 4087
rect 25259 3899 25271 4075
rect 25305 3899 25317 4075
rect 25259 3887 25317 3899
rect 25373 4075 25431 4087
rect 25373 3899 25385 4075
rect 25419 3899 25431 4075
rect 25373 3887 25431 3899
rect 25631 4075 25689 4087
rect 25631 3899 25643 4075
rect 25677 3899 25689 4075
rect 25631 3887 25689 3899
rect 25745 4075 25803 4087
rect 25745 3899 25757 4075
rect 25791 3899 25803 4075
rect 25745 3887 25803 3899
rect 26003 4075 26061 4087
rect 26003 3899 26015 4075
rect 26049 3899 26061 4075
rect 26003 3887 26061 3899
rect 26117 4075 26175 4087
rect 26117 3899 26129 4075
rect 26163 3899 26175 4075
rect 26117 3887 26175 3899
rect 26375 4075 26433 4087
rect 26375 3899 26387 4075
rect 26421 3899 26433 4075
rect 26375 3887 26433 3899
rect 26489 4075 26547 4087
rect 26489 3899 26501 4075
rect 26535 3899 26547 4075
rect 26489 3887 26547 3899
rect 26747 4075 26805 4087
rect 26747 3899 26759 4075
rect 26793 3899 26805 4075
rect 26747 3887 26805 3899
rect 26861 4075 26919 4087
rect 26861 3899 26873 4075
rect 26907 3899 26919 4075
rect 26861 3887 26919 3899
rect 27119 4075 27177 4087
rect 27119 3899 27131 4075
rect 27165 3899 27177 4075
rect 27119 3887 27177 3899
rect 27233 4075 27291 4087
rect 27233 3899 27245 4075
rect 27279 3899 27291 4075
rect 27233 3887 27291 3899
rect 27491 4075 27549 4087
rect 27491 3899 27503 4075
rect 27537 3899 27549 4075
rect 27491 3887 27549 3899
rect 27605 4075 27663 4087
rect 27605 3899 27617 4075
rect 27651 3899 27663 4075
rect 27605 3887 27663 3899
rect 27863 4075 27921 4087
rect 27863 3899 27875 4075
rect 27909 3899 27921 4075
rect 27863 3887 27921 3899
rect 27977 4075 28035 4087
rect 27977 3899 27989 4075
rect 28023 3899 28035 4075
rect 27977 3887 28035 3899
rect 28235 4075 28293 4087
rect 28235 3899 28247 4075
rect 28281 3899 28293 4075
rect 28235 3887 28293 3899
rect 28349 4075 28407 4087
rect 28349 3899 28361 4075
rect 28395 3899 28407 4075
rect 28349 3887 28407 3899
rect 28607 4075 28665 4087
rect 28607 3899 28619 4075
rect 28653 3899 28665 4075
rect 28607 3887 28665 3899
rect 28721 4075 28779 4087
rect 28721 3899 28733 4075
rect 28767 3899 28779 4075
rect 28721 3887 28779 3899
rect 28979 4075 29037 4087
rect 28979 3899 28991 4075
rect 29025 3899 29037 4075
rect 28979 3887 29037 3899
rect 20165 3657 20223 3669
rect 20165 3481 20177 3657
rect 20211 3481 20223 3657
rect 20165 3469 20223 3481
rect 20423 3657 20481 3669
rect 20423 3481 20435 3657
rect 20469 3481 20481 3657
rect 20423 3469 20481 3481
rect 20537 3657 20595 3669
rect 20537 3481 20549 3657
rect 20583 3481 20595 3657
rect 20537 3469 20595 3481
rect 20795 3657 20853 3669
rect 20795 3481 20807 3657
rect 20841 3481 20853 3657
rect 20795 3469 20853 3481
rect 20909 3657 20967 3669
rect 20909 3481 20921 3657
rect 20955 3481 20967 3657
rect 20909 3469 20967 3481
rect 21167 3657 21225 3669
rect 21167 3481 21179 3657
rect 21213 3481 21225 3657
rect 21167 3469 21225 3481
rect 21281 3657 21339 3669
rect 21281 3481 21293 3657
rect 21327 3481 21339 3657
rect 21281 3469 21339 3481
rect 21539 3657 21597 3669
rect 21539 3481 21551 3657
rect 21585 3481 21597 3657
rect 21539 3469 21597 3481
rect 21653 3657 21711 3669
rect 21653 3481 21665 3657
rect 21699 3481 21711 3657
rect 21653 3469 21711 3481
rect 21911 3657 21969 3669
rect 21911 3481 21923 3657
rect 21957 3481 21969 3657
rect 21911 3469 21969 3481
rect 22025 3657 22083 3669
rect 22025 3481 22037 3657
rect 22071 3481 22083 3657
rect 22025 3469 22083 3481
rect 22283 3657 22341 3669
rect 22283 3481 22295 3657
rect 22329 3481 22341 3657
rect 22283 3469 22341 3481
rect 22397 3657 22455 3669
rect 22397 3481 22409 3657
rect 22443 3481 22455 3657
rect 22397 3469 22455 3481
rect 22655 3657 22713 3669
rect 22655 3481 22667 3657
rect 22701 3481 22713 3657
rect 22655 3469 22713 3481
rect 22769 3657 22827 3669
rect 22769 3481 22781 3657
rect 22815 3481 22827 3657
rect 22769 3469 22827 3481
rect 23027 3657 23085 3669
rect 23027 3481 23039 3657
rect 23073 3481 23085 3657
rect 23027 3469 23085 3481
rect 23141 3657 23199 3669
rect 23141 3481 23153 3657
rect 23187 3481 23199 3657
rect 23141 3469 23199 3481
rect 23399 3657 23457 3669
rect 23399 3481 23411 3657
rect 23445 3481 23457 3657
rect 23399 3469 23457 3481
rect 23513 3657 23571 3669
rect 23513 3481 23525 3657
rect 23559 3481 23571 3657
rect 23513 3469 23571 3481
rect 23771 3657 23829 3669
rect 23771 3481 23783 3657
rect 23817 3481 23829 3657
rect 23771 3469 23829 3481
rect 23885 3657 23943 3669
rect 23885 3481 23897 3657
rect 23931 3481 23943 3657
rect 23885 3469 23943 3481
rect 24143 3657 24201 3669
rect 24143 3481 24155 3657
rect 24189 3481 24201 3657
rect 24143 3469 24201 3481
rect 24257 3657 24315 3669
rect 24257 3481 24269 3657
rect 24303 3481 24315 3657
rect 24257 3469 24315 3481
rect 24515 3657 24573 3669
rect 24515 3481 24527 3657
rect 24561 3481 24573 3657
rect 24515 3469 24573 3481
rect 24629 3657 24687 3669
rect 24629 3481 24641 3657
rect 24675 3481 24687 3657
rect 24629 3469 24687 3481
rect 24887 3657 24945 3669
rect 24887 3481 24899 3657
rect 24933 3481 24945 3657
rect 24887 3469 24945 3481
rect 25001 3657 25059 3669
rect 25001 3481 25013 3657
rect 25047 3481 25059 3657
rect 25001 3469 25059 3481
rect 25259 3657 25317 3669
rect 25259 3481 25271 3657
rect 25305 3481 25317 3657
rect 25259 3469 25317 3481
rect 25373 3657 25431 3669
rect 25373 3481 25385 3657
rect 25419 3481 25431 3657
rect 25373 3469 25431 3481
rect 25631 3657 25689 3669
rect 25631 3481 25643 3657
rect 25677 3481 25689 3657
rect 25631 3469 25689 3481
rect 25745 3657 25803 3669
rect 25745 3481 25757 3657
rect 25791 3481 25803 3657
rect 25745 3469 25803 3481
rect 26003 3657 26061 3669
rect 26003 3481 26015 3657
rect 26049 3481 26061 3657
rect 26003 3469 26061 3481
rect 26117 3657 26175 3669
rect 26117 3481 26129 3657
rect 26163 3481 26175 3657
rect 26117 3469 26175 3481
rect 26375 3657 26433 3669
rect 26375 3481 26387 3657
rect 26421 3481 26433 3657
rect 26375 3469 26433 3481
rect 26489 3657 26547 3669
rect 26489 3481 26501 3657
rect 26535 3481 26547 3657
rect 26489 3469 26547 3481
rect 26747 3657 26805 3669
rect 26747 3481 26759 3657
rect 26793 3481 26805 3657
rect 26747 3469 26805 3481
rect 26861 3657 26919 3669
rect 26861 3481 26873 3657
rect 26907 3481 26919 3657
rect 26861 3469 26919 3481
rect 27119 3657 27177 3669
rect 27119 3481 27131 3657
rect 27165 3481 27177 3657
rect 27119 3469 27177 3481
rect 27233 3657 27291 3669
rect 27233 3481 27245 3657
rect 27279 3481 27291 3657
rect 27233 3469 27291 3481
rect 27491 3657 27549 3669
rect 27491 3481 27503 3657
rect 27537 3481 27549 3657
rect 27491 3469 27549 3481
rect 27605 3657 27663 3669
rect 27605 3481 27617 3657
rect 27651 3481 27663 3657
rect 27605 3469 27663 3481
rect 27863 3657 27921 3669
rect 27863 3481 27875 3657
rect 27909 3481 27921 3657
rect 27863 3469 27921 3481
rect 27977 3657 28035 3669
rect 27977 3481 27989 3657
rect 28023 3481 28035 3657
rect 27977 3469 28035 3481
rect 28235 3657 28293 3669
rect 28235 3481 28247 3657
rect 28281 3481 28293 3657
rect 28235 3469 28293 3481
rect 28349 3657 28407 3669
rect 28349 3481 28361 3657
rect 28395 3481 28407 3657
rect 28349 3469 28407 3481
rect 28607 3657 28665 3669
rect 28607 3481 28619 3657
rect 28653 3481 28665 3657
rect 28607 3469 28665 3481
rect 28721 3657 28779 3669
rect 28721 3481 28733 3657
rect 28767 3481 28779 3657
rect 28721 3469 28779 3481
rect 28979 3657 29037 3669
rect 28979 3481 28991 3657
rect 29025 3481 29037 3657
rect 28979 3469 29037 3481
rect 20165 3239 20223 3251
rect 20165 3063 20177 3239
rect 20211 3063 20223 3239
rect 20165 3051 20223 3063
rect 20423 3239 20481 3251
rect 20423 3063 20435 3239
rect 20469 3063 20481 3239
rect 20423 3051 20481 3063
rect 20537 3239 20595 3251
rect 20537 3063 20549 3239
rect 20583 3063 20595 3239
rect 20537 3051 20595 3063
rect 20795 3239 20853 3251
rect 20795 3063 20807 3239
rect 20841 3063 20853 3239
rect 20795 3051 20853 3063
rect 20909 3239 20967 3251
rect 20909 3063 20921 3239
rect 20955 3063 20967 3239
rect 20909 3051 20967 3063
rect 21167 3239 21225 3251
rect 21167 3063 21179 3239
rect 21213 3063 21225 3239
rect 21167 3051 21225 3063
rect 21281 3239 21339 3251
rect 21281 3063 21293 3239
rect 21327 3063 21339 3239
rect 21281 3051 21339 3063
rect 21539 3239 21597 3251
rect 21539 3063 21551 3239
rect 21585 3063 21597 3239
rect 21539 3051 21597 3063
rect 21653 3239 21711 3251
rect 21653 3063 21665 3239
rect 21699 3063 21711 3239
rect 21653 3051 21711 3063
rect 21911 3239 21969 3251
rect 21911 3063 21923 3239
rect 21957 3063 21969 3239
rect 21911 3051 21969 3063
rect 22025 3239 22083 3251
rect 22025 3063 22037 3239
rect 22071 3063 22083 3239
rect 22025 3051 22083 3063
rect 22283 3239 22341 3251
rect 22283 3063 22295 3239
rect 22329 3063 22341 3239
rect 22283 3051 22341 3063
rect 22397 3239 22455 3251
rect 22397 3063 22409 3239
rect 22443 3063 22455 3239
rect 22397 3051 22455 3063
rect 22655 3239 22713 3251
rect 22655 3063 22667 3239
rect 22701 3063 22713 3239
rect 22655 3051 22713 3063
rect 22769 3239 22827 3251
rect 22769 3063 22781 3239
rect 22815 3063 22827 3239
rect 22769 3051 22827 3063
rect 23027 3239 23085 3251
rect 23027 3063 23039 3239
rect 23073 3063 23085 3239
rect 23027 3051 23085 3063
rect 23141 3239 23199 3251
rect 23141 3063 23153 3239
rect 23187 3063 23199 3239
rect 23141 3051 23199 3063
rect 23399 3239 23457 3251
rect 23399 3063 23411 3239
rect 23445 3063 23457 3239
rect 23399 3051 23457 3063
rect 23513 3239 23571 3251
rect 23513 3063 23525 3239
rect 23559 3063 23571 3239
rect 23513 3051 23571 3063
rect 23771 3239 23829 3251
rect 23771 3063 23783 3239
rect 23817 3063 23829 3239
rect 23771 3051 23829 3063
rect 23885 3239 23943 3251
rect 23885 3063 23897 3239
rect 23931 3063 23943 3239
rect 23885 3051 23943 3063
rect 24143 3239 24201 3251
rect 24143 3063 24155 3239
rect 24189 3063 24201 3239
rect 24143 3051 24201 3063
rect 24257 3239 24315 3251
rect 24257 3063 24269 3239
rect 24303 3063 24315 3239
rect 24257 3051 24315 3063
rect 24515 3239 24573 3251
rect 24515 3063 24527 3239
rect 24561 3063 24573 3239
rect 24515 3051 24573 3063
rect 24629 3239 24687 3251
rect 24629 3063 24641 3239
rect 24675 3063 24687 3239
rect 24629 3051 24687 3063
rect 24887 3239 24945 3251
rect 24887 3063 24899 3239
rect 24933 3063 24945 3239
rect 24887 3051 24945 3063
rect 25001 3239 25059 3251
rect 25001 3063 25013 3239
rect 25047 3063 25059 3239
rect 25001 3051 25059 3063
rect 25259 3239 25317 3251
rect 25259 3063 25271 3239
rect 25305 3063 25317 3239
rect 25259 3051 25317 3063
rect 25373 3239 25431 3251
rect 25373 3063 25385 3239
rect 25419 3063 25431 3239
rect 25373 3051 25431 3063
rect 25631 3239 25689 3251
rect 25631 3063 25643 3239
rect 25677 3063 25689 3239
rect 25631 3051 25689 3063
rect 25745 3239 25803 3251
rect 25745 3063 25757 3239
rect 25791 3063 25803 3239
rect 25745 3051 25803 3063
rect 26003 3239 26061 3251
rect 26003 3063 26015 3239
rect 26049 3063 26061 3239
rect 26003 3051 26061 3063
rect 26117 3239 26175 3251
rect 26117 3063 26129 3239
rect 26163 3063 26175 3239
rect 26117 3051 26175 3063
rect 26375 3239 26433 3251
rect 26375 3063 26387 3239
rect 26421 3063 26433 3239
rect 26375 3051 26433 3063
rect 26489 3239 26547 3251
rect 26489 3063 26501 3239
rect 26535 3063 26547 3239
rect 26489 3051 26547 3063
rect 26747 3239 26805 3251
rect 26747 3063 26759 3239
rect 26793 3063 26805 3239
rect 26747 3051 26805 3063
rect 26861 3239 26919 3251
rect 26861 3063 26873 3239
rect 26907 3063 26919 3239
rect 26861 3051 26919 3063
rect 27119 3239 27177 3251
rect 27119 3063 27131 3239
rect 27165 3063 27177 3239
rect 27119 3051 27177 3063
rect 27233 3239 27291 3251
rect 27233 3063 27245 3239
rect 27279 3063 27291 3239
rect 27233 3051 27291 3063
rect 27491 3239 27549 3251
rect 27491 3063 27503 3239
rect 27537 3063 27549 3239
rect 27491 3051 27549 3063
rect 27605 3239 27663 3251
rect 27605 3063 27617 3239
rect 27651 3063 27663 3239
rect 27605 3051 27663 3063
rect 27863 3239 27921 3251
rect 27863 3063 27875 3239
rect 27909 3063 27921 3239
rect 27863 3051 27921 3063
rect 27977 3239 28035 3251
rect 27977 3063 27989 3239
rect 28023 3063 28035 3239
rect 27977 3051 28035 3063
rect 28235 3239 28293 3251
rect 28235 3063 28247 3239
rect 28281 3063 28293 3239
rect 28235 3051 28293 3063
rect 28349 3239 28407 3251
rect 28349 3063 28361 3239
rect 28395 3063 28407 3239
rect 28349 3051 28407 3063
rect 28607 3239 28665 3251
rect 28607 3063 28619 3239
rect 28653 3063 28665 3239
rect 28607 3051 28665 3063
rect 28721 3239 28779 3251
rect 28721 3063 28733 3239
rect 28767 3063 28779 3239
rect 28721 3051 28779 3063
rect 28979 3239 29037 3251
rect 28979 3063 28991 3239
rect 29025 3063 29037 3239
rect 28979 3051 29037 3063
<< pdiff >>
rect 18677 11566 18735 11578
rect 18677 11190 18689 11566
rect 18723 11190 18735 11566
rect 18677 11178 18735 11190
rect 18935 11566 18993 11578
rect 18935 11190 18947 11566
rect 18981 11190 18993 11566
rect 18935 11178 18993 11190
rect 19049 11566 19107 11578
rect 19049 11190 19061 11566
rect 19095 11190 19107 11566
rect 19049 11178 19107 11190
rect 19307 11566 19365 11578
rect 19307 11190 19319 11566
rect 19353 11190 19365 11566
rect 19307 11178 19365 11190
rect 19421 11566 19479 11578
rect 19421 11190 19433 11566
rect 19467 11190 19479 11566
rect 19421 11178 19479 11190
rect 19679 11566 19737 11578
rect 19679 11190 19691 11566
rect 19725 11190 19737 11566
rect 19679 11178 19737 11190
rect 19793 11566 19851 11578
rect 19793 11190 19805 11566
rect 19839 11190 19851 11566
rect 19793 11178 19851 11190
rect 20051 11566 20109 11578
rect 20051 11190 20063 11566
rect 20097 11190 20109 11566
rect 20051 11178 20109 11190
rect 20165 11566 20223 11578
rect 20165 11190 20177 11566
rect 20211 11190 20223 11566
rect 20165 11178 20223 11190
rect 20423 11566 20481 11578
rect 20423 11190 20435 11566
rect 20469 11190 20481 11566
rect 20423 11178 20481 11190
rect 20537 11566 20595 11578
rect 20537 11190 20549 11566
rect 20583 11190 20595 11566
rect 20537 11178 20595 11190
rect 20795 11566 20853 11578
rect 20795 11190 20807 11566
rect 20841 11190 20853 11566
rect 20795 11178 20853 11190
rect 20909 11566 20967 11578
rect 20909 11190 20921 11566
rect 20955 11190 20967 11566
rect 20909 11178 20967 11190
rect 21167 11566 21225 11578
rect 21167 11190 21179 11566
rect 21213 11190 21225 11566
rect 21167 11178 21225 11190
rect 21281 11566 21339 11578
rect 21281 11190 21293 11566
rect 21327 11190 21339 11566
rect 21281 11178 21339 11190
rect 21539 11566 21597 11578
rect 21539 11190 21551 11566
rect 21585 11190 21597 11566
rect 21539 11178 21597 11190
rect 21653 11566 21711 11578
rect 21653 11190 21665 11566
rect 21699 11190 21711 11566
rect 21653 11178 21711 11190
rect 21911 11566 21969 11578
rect 21911 11190 21923 11566
rect 21957 11190 21969 11566
rect 21911 11178 21969 11190
rect 22025 11566 22083 11578
rect 22025 11190 22037 11566
rect 22071 11190 22083 11566
rect 22025 11178 22083 11190
rect 22283 11566 22341 11578
rect 22283 11190 22295 11566
rect 22329 11190 22341 11566
rect 22283 11178 22341 11190
rect 22397 11566 22455 11578
rect 22397 11190 22409 11566
rect 22443 11190 22455 11566
rect 22397 11178 22455 11190
rect 22655 11566 22713 11578
rect 22655 11190 22667 11566
rect 22701 11190 22713 11566
rect 22655 11178 22713 11190
rect 22769 11566 22827 11578
rect 22769 11190 22781 11566
rect 22815 11190 22827 11566
rect 22769 11178 22827 11190
rect 23027 11566 23085 11578
rect 23027 11190 23039 11566
rect 23073 11190 23085 11566
rect 23027 11178 23085 11190
rect 23141 11566 23199 11578
rect 23141 11190 23153 11566
rect 23187 11190 23199 11566
rect 23141 11178 23199 11190
rect 23399 11566 23457 11578
rect 23399 11190 23411 11566
rect 23445 11190 23457 11566
rect 23399 11178 23457 11190
rect 23513 11566 23571 11578
rect 23513 11190 23525 11566
rect 23559 11190 23571 11566
rect 23513 11178 23571 11190
rect 23771 11566 23829 11578
rect 23771 11190 23783 11566
rect 23817 11190 23829 11566
rect 23771 11178 23829 11190
rect 23885 11566 23943 11578
rect 23885 11190 23897 11566
rect 23931 11190 23943 11566
rect 23885 11178 23943 11190
rect 24143 11566 24201 11578
rect 24143 11190 24155 11566
rect 24189 11190 24201 11566
rect 24143 11178 24201 11190
rect 24257 11566 24315 11578
rect 24257 11190 24269 11566
rect 24303 11190 24315 11566
rect 24257 11178 24315 11190
rect 24515 11566 24573 11578
rect 24515 11190 24527 11566
rect 24561 11190 24573 11566
rect 24515 11178 24573 11190
rect 24629 11566 24687 11578
rect 24629 11190 24641 11566
rect 24675 11190 24687 11566
rect 24629 11178 24687 11190
rect 24887 11566 24945 11578
rect 24887 11190 24899 11566
rect 24933 11190 24945 11566
rect 24887 11178 24945 11190
rect 25001 11566 25059 11578
rect 25001 11190 25013 11566
rect 25047 11190 25059 11566
rect 25001 11178 25059 11190
rect 25259 11566 25317 11578
rect 25259 11190 25271 11566
rect 25305 11190 25317 11566
rect 25259 11178 25317 11190
rect 25373 11566 25431 11578
rect 25373 11190 25385 11566
rect 25419 11190 25431 11566
rect 25373 11178 25431 11190
rect 25631 11566 25689 11578
rect 25631 11190 25643 11566
rect 25677 11190 25689 11566
rect 25631 11178 25689 11190
rect 25745 11566 25803 11578
rect 25745 11190 25757 11566
rect 25791 11190 25803 11566
rect 25745 11178 25803 11190
rect 26003 11566 26061 11578
rect 26003 11190 26015 11566
rect 26049 11190 26061 11566
rect 26003 11178 26061 11190
rect 26117 11566 26175 11578
rect 26117 11190 26129 11566
rect 26163 11190 26175 11566
rect 26117 11178 26175 11190
rect 26375 11566 26433 11578
rect 26375 11190 26387 11566
rect 26421 11190 26433 11566
rect 26375 11178 26433 11190
rect 26489 11566 26547 11578
rect 26489 11190 26501 11566
rect 26535 11190 26547 11566
rect 26489 11178 26547 11190
rect 26747 11566 26805 11578
rect 26747 11190 26759 11566
rect 26793 11190 26805 11566
rect 26747 11178 26805 11190
rect 26861 11566 26919 11578
rect 26861 11190 26873 11566
rect 26907 11190 26919 11566
rect 26861 11178 26919 11190
rect 27119 11566 27177 11578
rect 27119 11190 27131 11566
rect 27165 11190 27177 11566
rect 27119 11178 27177 11190
rect 27233 11566 27291 11578
rect 27233 11190 27245 11566
rect 27279 11190 27291 11566
rect 27233 11178 27291 11190
rect 27491 11566 27549 11578
rect 27491 11190 27503 11566
rect 27537 11190 27549 11566
rect 27491 11178 27549 11190
rect 27605 11566 27663 11578
rect 27605 11190 27617 11566
rect 27651 11190 27663 11566
rect 27605 11178 27663 11190
rect 27863 11566 27921 11578
rect 27863 11190 27875 11566
rect 27909 11190 27921 11566
rect 27863 11178 27921 11190
rect 27977 11566 28035 11578
rect 27977 11190 27989 11566
rect 28023 11190 28035 11566
rect 27977 11178 28035 11190
rect 28235 11566 28293 11578
rect 28235 11190 28247 11566
rect 28281 11190 28293 11566
rect 28235 11178 28293 11190
rect 28349 11566 28407 11578
rect 28349 11190 28361 11566
rect 28395 11190 28407 11566
rect 28349 11178 28407 11190
rect 28607 11566 28665 11578
rect 28607 11190 28619 11566
rect 28653 11190 28665 11566
rect 28607 11178 28665 11190
rect 28721 11566 28779 11578
rect 28721 11190 28733 11566
rect 28767 11190 28779 11566
rect 28721 11178 28779 11190
rect 28979 11566 29037 11578
rect 28979 11190 28991 11566
rect 29025 11190 29037 11566
rect 28979 11178 29037 11190
rect 29093 11566 29151 11578
rect 29093 11190 29105 11566
rect 29139 11190 29151 11566
rect 29093 11178 29151 11190
rect 29351 11566 29409 11578
rect 29351 11190 29363 11566
rect 29397 11190 29409 11566
rect 29351 11178 29409 11190
rect 29465 11566 29523 11578
rect 29465 11190 29477 11566
rect 29511 11190 29523 11566
rect 29465 11178 29523 11190
rect 29723 11566 29781 11578
rect 29723 11190 29735 11566
rect 29769 11190 29781 11566
rect 29723 11178 29781 11190
rect 29837 11566 29895 11578
rect 29837 11190 29849 11566
rect 29883 11190 29895 11566
rect 29837 11178 29895 11190
rect 30095 11566 30153 11578
rect 30095 11190 30107 11566
rect 30141 11190 30153 11566
rect 30095 11178 30153 11190
rect 30209 11566 30267 11578
rect 30209 11190 30221 11566
rect 30255 11190 30267 11566
rect 30209 11178 30267 11190
rect 30467 11566 30525 11578
rect 30467 11190 30479 11566
rect 30513 11190 30525 11566
rect 30467 11178 30525 11190
rect 18677 10930 18735 10942
rect 18677 10554 18689 10930
rect 18723 10554 18735 10930
rect 18677 10542 18735 10554
rect 18935 10930 18993 10942
rect 18935 10554 18947 10930
rect 18981 10554 18993 10930
rect 18935 10542 18993 10554
rect 19049 10930 19107 10942
rect 19049 10554 19061 10930
rect 19095 10554 19107 10930
rect 19049 10542 19107 10554
rect 19307 10930 19365 10942
rect 19307 10554 19319 10930
rect 19353 10554 19365 10930
rect 19307 10542 19365 10554
rect 19421 10930 19479 10942
rect 19421 10554 19433 10930
rect 19467 10554 19479 10930
rect 19421 10542 19479 10554
rect 19679 10930 19737 10942
rect 19679 10554 19691 10930
rect 19725 10554 19737 10930
rect 19679 10542 19737 10554
rect 19793 10930 19851 10942
rect 19793 10554 19805 10930
rect 19839 10554 19851 10930
rect 19793 10542 19851 10554
rect 20051 10930 20109 10942
rect 20051 10554 20063 10930
rect 20097 10554 20109 10930
rect 20051 10542 20109 10554
rect 20165 10930 20223 10942
rect 20165 10554 20177 10930
rect 20211 10554 20223 10930
rect 20165 10542 20223 10554
rect 20423 10930 20481 10942
rect 20423 10554 20435 10930
rect 20469 10554 20481 10930
rect 20423 10542 20481 10554
rect 20537 10930 20595 10942
rect 20537 10554 20549 10930
rect 20583 10554 20595 10930
rect 20537 10542 20595 10554
rect 20795 10930 20853 10942
rect 20795 10554 20807 10930
rect 20841 10554 20853 10930
rect 20795 10542 20853 10554
rect 20909 10930 20967 10942
rect 20909 10554 20921 10930
rect 20955 10554 20967 10930
rect 20909 10542 20967 10554
rect 21167 10930 21225 10942
rect 21167 10554 21179 10930
rect 21213 10554 21225 10930
rect 21167 10542 21225 10554
rect 21281 10930 21339 10942
rect 21281 10554 21293 10930
rect 21327 10554 21339 10930
rect 21281 10542 21339 10554
rect 21539 10930 21597 10942
rect 21539 10554 21551 10930
rect 21585 10554 21597 10930
rect 21539 10542 21597 10554
rect 21653 10930 21711 10942
rect 21653 10554 21665 10930
rect 21699 10554 21711 10930
rect 21653 10542 21711 10554
rect 21911 10930 21969 10942
rect 21911 10554 21923 10930
rect 21957 10554 21969 10930
rect 21911 10542 21969 10554
rect 22025 10930 22083 10942
rect 22025 10554 22037 10930
rect 22071 10554 22083 10930
rect 22025 10542 22083 10554
rect 22283 10930 22341 10942
rect 22283 10554 22295 10930
rect 22329 10554 22341 10930
rect 22283 10542 22341 10554
rect 22397 10930 22455 10942
rect 22397 10554 22409 10930
rect 22443 10554 22455 10930
rect 22397 10542 22455 10554
rect 22655 10930 22713 10942
rect 22655 10554 22667 10930
rect 22701 10554 22713 10930
rect 22655 10542 22713 10554
rect 22769 10930 22827 10942
rect 22769 10554 22781 10930
rect 22815 10554 22827 10930
rect 22769 10542 22827 10554
rect 23027 10930 23085 10942
rect 23027 10554 23039 10930
rect 23073 10554 23085 10930
rect 23027 10542 23085 10554
rect 23141 10930 23199 10942
rect 23141 10554 23153 10930
rect 23187 10554 23199 10930
rect 23141 10542 23199 10554
rect 23399 10930 23457 10942
rect 23399 10554 23411 10930
rect 23445 10554 23457 10930
rect 23399 10542 23457 10554
rect 23513 10930 23571 10942
rect 23513 10554 23525 10930
rect 23559 10554 23571 10930
rect 23513 10542 23571 10554
rect 23771 10930 23829 10942
rect 23771 10554 23783 10930
rect 23817 10554 23829 10930
rect 23771 10542 23829 10554
rect 23885 10930 23943 10942
rect 23885 10554 23897 10930
rect 23931 10554 23943 10930
rect 23885 10542 23943 10554
rect 24143 10930 24201 10942
rect 24143 10554 24155 10930
rect 24189 10554 24201 10930
rect 24143 10542 24201 10554
rect 24257 10930 24315 10942
rect 24257 10554 24269 10930
rect 24303 10554 24315 10930
rect 24257 10542 24315 10554
rect 24515 10930 24573 10942
rect 24515 10554 24527 10930
rect 24561 10554 24573 10930
rect 24515 10542 24573 10554
rect 24629 10930 24687 10942
rect 24629 10554 24641 10930
rect 24675 10554 24687 10930
rect 24629 10542 24687 10554
rect 24887 10930 24945 10942
rect 24887 10554 24899 10930
rect 24933 10554 24945 10930
rect 24887 10542 24945 10554
rect 25001 10930 25059 10942
rect 25001 10554 25013 10930
rect 25047 10554 25059 10930
rect 25001 10542 25059 10554
rect 25259 10930 25317 10942
rect 25259 10554 25271 10930
rect 25305 10554 25317 10930
rect 25259 10542 25317 10554
rect 25373 10930 25431 10942
rect 25373 10554 25385 10930
rect 25419 10554 25431 10930
rect 25373 10542 25431 10554
rect 25631 10930 25689 10942
rect 25631 10554 25643 10930
rect 25677 10554 25689 10930
rect 25631 10542 25689 10554
rect 25745 10930 25803 10942
rect 25745 10554 25757 10930
rect 25791 10554 25803 10930
rect 25745 10542 25803 10554
rect 26003 10930 26061 10942
rect 26003 10554 26015 10930
rect 26049 10554 26061 10930
rect 26003 10542 26061 10554
rect 26117 10930 26175 10942
rect 26117 10554 26129 10930
rect 26163 10554 26175 10930
rect 26117 10542 26175 10554
rect 26375 10930 26433 10942
rect 26375 10554 26387 10930
rect 26421 10554 26433 10930
rect 26375 10542 26433 10554
rect 26489 10930 26547 10942
rect 26489 10554 26501 10930
rect 26535 10554 26547 10930
rect 26489 10542 26547 10554
rect 26747 10930 26805 10942
rect 26747 10554 26759 10930
rect 26793 10554 26805 10930
rect 26747 10542 26805 10554
rect 26861 10930 26919 10942
rect 26861 10554 26873 10930
rect 26907 10554 26919 10930
rect 26861 10542 26919 10554
rect 27119 10930 27177 10942
rect 27119 10554 27131 10930
rect 27165 10554 27177 10930
rect 27119 10542 27177 10554
rect 27233 10930 27291 10942
rect 27233 10554 27245 10930
rect 27279 10554 27291 10930
rect 27233 10542 27291 10554
rect 27491 10930 27549 10942
rect 27491 10554 27503 10930
rect 27537 10554 27549 10930
rect 27491 10542 27549 10554
rect 27605 10930 27663 10942
rect 27605 10554 27617 10930
rect 27651 10554 27663 10930
rect 27605 10542 27663 10554
rect 27863 10930 27921 10942
rect 27863 10554 27875 10930
rect 27909 10554 27921 10930
rect 27863 10542 27921 10554
rect 27977 10930 28035 10942
rect 27977 10554 27989 10930
rect 28023 10554 28035 10930
rect 27977 10542 28035 10554
rect 28235 10930 28293 10942
rect 28235 10554 28247 10930
rect 28281 10554 28293 10930
rect 28235 10542 28293 10554
rect 28349 10930 28407 10942
rect 28349 10554 28361 10930
rect 28395 10554 28407 10930
rect 28349 10542 28407 10554
rect 28607 10930 28665 10942
rect 28607 10554 28619 10930
rect 28653 10554 28665 10930
rect 28607 10542 28665 10554
rect 28721 10930 28779 10942
rect 28721 10554 28733 10930
rect 28767 10554 28779 10930
rect 28721 10542 28779 10554
rect 28979 10930 29037 10942
rect 28979 10554 28991 10930
rect 29025 10554 29037 10930
rect 28979 10542 29037 10554
rect 29093 10930 29151 10942
rect 29093 10554 29105 10930
rect 29139 10554 29151 10930
rect 29093 10542 29151 10554
rect 29351 10930 29409 10942
rect 29351 10554 29363 10930
rect 29397 10554 29409 10930
rect 29351 10542 29409 10554
rect 29465 10930 29523 10942
rect 29465 10554 29477 10930
rect 29511 10554 29523 10930
rect 29465 10542 29523 10554
rect 29723 10930 29781 10942
rect 29723 10554 29735 10930
rect 29769 10554 29781 10930
rect 29723 10542 29781 10554
rect 29837 10930 29895 10942
rect 29837 10554 29849 10930
rect 29883 10554 29895 10930
rect 29837 10542 29895 10554
rect 30095 10930 30153 10942
rect 30095 10554 30107 10930
rect 30141 10554 30153 10930
rect 30095 10542 30153 10554
rect 30209 10930 30267 10942
rect 30209 10554 30221 10930
rect 30255 10554 30267 10930
rect 30209 10542 30267 10554
rect 30467 10930 30525 10942
rect 30467 10554 30479 10930
rect 30513 10554 30525 10930
rect 30467 10542 30525 10554
rect 18677 10294 18735 10306
rect 18677 9918 18689 10294
rect 18723 9918 18735 10294
rect 18677 9906 18735 9918
rect 18935 10294 18993 10306
rect 18935 9918 18947 10294
rect 18981 9918 18993 10294
rect 18935 9906 18993 9918
rect 19049 10294 19107 10306
rect 19049 9918 19061 10294
rect 19095 9918 19107 10294
rect 19049 9906 19107 9918
rect 19307 10294 19365 10306
rect 19307 9918 19319 10294
rect 19353 9918 19365 10294
rect 19307 9906 19365 9918
rect 19421 10294 19479 10306
rect 19421 9918 19433 10294
rect 19467 9918 19479 10294
rect 19421 9906 19479 9918
rect 19679 10294 19737 10306
rect 19679 9918 19691 10294
rect 19725 9918 19737 10294
rect 19679 9906 19737 9918
rect 19793 10294 19851 10306
rect 19793 9918 19805 10294
rect 19839 9918 19851 10294
rect 19793 9906 19851 9918
rect 20051 10294 20109 10306
rect 20051 9918 20063 10294
rect 20097 9918 20109 10294
rect 20051 9906 20109 9918
rect 20165 10294 20223 10306
rect 20165 9918 20177 10294
rect 20211 9918 20223 10294
rect 20165 9906 20223 9918
rect 20423 10294 20481 10306
rect 20423 9918 20435 10294
rect 20469 9918 20481 10294
rect 20423 9906 20481 9918
rect 20537 10294 20595 10306
rect 20537 9918 20549 10294
rect 20583 9918 20595 10294
rect 20537 9906 20595 9918
rect 20795 10294 20853 10306
rect 20795 9918 20807 10294
rect 20841 9918 20853 10294
rect 20795 9906 20853 9918
rect 20909 10294 20967 10306
rect 20909 9918 20921 10294
rect 20955 9918 20967 10294
rect 20909 9906 20967 9918
rect 21167 10294 21225 10306
rect 21167 9918 21179 10294
rect 21213 9918 21225 10294
rect 21167 9906 21225 9918
rect 21281 10294 21339 10306
rect 21281 9918 21293 10294
rect 21327 9918 21339 10294
rect 21281 9906 21339 9918
rect 21539 10294 21597 10306
rect 21539 9918 21551 10294
rect 21585 9918 21597 10294
rect 21539 9906 21597 9918
rect 21653 10294 21711 10306
rect 21653 9918 21665 10294
rect 21699 9918 21711 10294
rect 21653 9906 21711 9918
rect 21911 10294 21969 10306
rect 21911 9918 21923 10294
rect 21957 9918 21969 10294
rect 21911 9906 21969 9918
rect 22025 10294 22083 10306
rect 22025 9918 22037 10294
rect 22071 9918 22083 10294
rect 22025 9906 22083 9918
rect 22283 10294 22341 10306
rect 22283 9918 22295 10294
rect 22329 9918 22341 10294
rect 22283 9906 22341 9918
rect 22397 10294 22455 10306
rect 22397 9918 22409 10294
rect 22443 9918 22455 10294
rect 22397 9906 22455 9918
rect 22655 10294 22713 10306
rect 22655 9918 22667 10294
rect 22701 9918 22713 10294
rect 22655 9906 22713 9918
rect 22769 10294 22827 10306
rect 22769 9918 22781 10294
rect 22815 9918 22827 10294
rect 22769 9906 22827 9918
rect 23027 10294 23085 10306
rect 23027 9918 23039 10294
rect 23073 9918 23085 10294
rect 23027 9906 23085 9918
rect 23141 10294 23199 10306
rect 23141 9918 23153 10294
rect 23187 9918 23199 10294
rect 23141 9906 23199 9918
rect 23399 10294 23457 10306
rect 23399 9918 23411 10294
rect 23445 9918 23457 10294
rect 23399 9906 23457 9918
rect 23513 10294 23571 10306
rect 23513 9918 23525 10294
rect 23559 9918 23571 10294
rect 23513 9906 23571 9918
rect 23771 10294 23829 10306
rect 23771 9918 23783 10294
rect 23817 9918 23829 10294
rect 23771 9906 23829 9918
rect 23885 10294 23943 10306
rect 23885 9918 23897 10294
rect 23931 9918 23943 10294
rect 23885 9906 23943 9918
rect 24143 10294 24201 10306
rect 24143 9918 24155 10294
rect 24189 9918 24201 10294
rect 24143 9906 24201 9918
rect 24257 10294 24315 10306
rect 24257 9918 24269 10294
rect 24303 9918 24315 10294
rect 24257 9906 24315 9918
rect 24515 10294 24573 10306
rect 24515 9918 24527 10294
rect 24561 9918 24573 10294
rect 24515 9906 24573 9918
rect 24629 10294 24687 10306
rect 24629 9918 24641 10294
rect 24675 9918 24687 10294
rect 24629 9906 24687 9918
rect 24887 10294 24945 10306
rect 24887 9918 24899 10294
rect 24933 9918 24945 10294
rect 24887 9906 24945 9918
rect 25001 10294 25059 10306
rect 25001 9918 25013 10294
rect 25047 9918 25059 10294
rect 25001 9906 25059 9918
rect 25259 10294 25317 10306
rect 25259 9918 25271 10294
rect 25305 9918 25317 10294
rect 25259 9906 25317 9918
rect 25373 10294 25431 10306
rect 25373 9918 25385 10294
rect 25419 9918 25431 10294
rect 25373 9906 25431 9918
rect 25631 10294 25689 10306
rect 25631 9918 25643 10294
rect 25677 9918 25689 10294
rect 25631 9906 25689 9918
rect 25745 10294 25803 10306
rect 25745 9918 25757 10294
rect 25791 9918 25803 10294
rect 25745 9906 25803 9918
rect 26003 10294 26061 10306
rect 26003 9918 26015 10294
rect 26049 9918 26061 10294
rect 26003 9906 26061 9918
rect 26117 10294 26175 10306
rect 26117 9918 26129 10294
rect 26163 9918 26175 10294
rect 26117 9906 26175 9918
rect 26375 10294 26433 10306
rect 26375 9918 26387 10294
rect 26421 9918 26433 10294
rect 26375 9906 26433 9918
rect 26489 10294 26547 10306
rect 26489 9918 26501 10294
rect 26535 9918 26547 10294
rect 26489 9906 26547 9918
rect 26747 10294 26805 10306
rect 26747 9918 26759 10294
rect 26793 9918 26805 10294
rect 26747 9906 26805 9918
rect 26861 10294 26919 10306
rect 26861 9918 26873 10294
rect 26907 9918 26919 10294
rect 26861 9906 26919 9918
rect 27119 10294 27177 10306
rect 27119 9918 27131 10294
rect 27165 9918 27177 10294
rect 27119 9906 27177 9918
rect 27233 10294 27291 10306
rect 27233 9918 27245 10294
rect 27279 9918 27291 10294
rect 27233 9906 27291 9918
rect 27491 10294 27549 10306
rect 27491 9918 27503 10294
rect 27537 9918 27549 10294
rect 27491 9906 27549 9918
rect 27605 10294 27663 10306
rect 27605 9918 27617 10294
rect 27651 9918 27663 10294
rect 27605 9906 27663 9918
rect 27863 10294 27921 10306
rect 27863 9918 27875 10294
rect 27909 9918 27921 10294
rect 27863 9906 27921 9918
rect 27977 10294 28035 10306
rect 27977 9918 27989 10294
rect 28023 9918 28035 10294
rect 27977 9906 28035 9918
rect 28235 10294 28293 10306
rect 28235 9918 28247 10294
rect 28281 9918 28293 10294
rect 28235 9906 28293 9918
rect 28349 10294 28407 10306
rect 28349 9918 28361 10294
rect 28395 9918 28407 10294
rect 28349 9906 28407 9918
rect 28607 10294 28665 10306
rect 28607 9918 28619 10294
rect 28653 9918 28665 10294
rect 28607 9906 28665 9918
rect 28721 10294 28779 10306
rect 28721 9918 28733 10294
rect 28767 9918 28779 10294
rect 28721 9906 28779 9918
rect 28979 10294 29037 10306
rect 28979 9918 28991 10294
rect 29025 9918 29037 10294
rect 28979 9906 29037 9918
rect 29093 10294 29151 10306
rect 29093 9918 29105 10294
rect 29139 9918 29151 10294
rect 29093 9906 29151 9918
rect 29351 10294 29409 10306
rect 29351 9918 29363 10294
rect 29397 9918 29409 10294
rect 29351 9906 29409 9918
rect 29465 10294 29523 10306
rect 29465 9918 29477 10294
rect 29511 9918 29523 10294
rect 29465 9906 29523 9918
rect 29723 10294 29781 10306
rect 29723 9918 29735 10294
rect 29769 9918 29781 10294
rect 29723 9906 29781 9918
rect 29837 10294 29895 10306
rect 29837 9918 29849 10294
rect 29883 9918 29895 10294
rect 29837 9906 29895 9918
rect 30095 10294 30153 10306
rect 30095 9918 30107 10294
rect 30141 9918 30153 10294
rect 30095 9906 30153 9918
rect 30209 10294 30267 10306
rect 30209 9918 30221 10294
rect 30255 9918 30267 10294
rect 30209 9906 30267 9918
rect 30467 10294 30525 10306
rect 30467 9918 30479 10294
rect 30513 9918 30525 10294
rect 30467 9906 30525 9918
rect 20165 9178 20223 9190
rect 20165 8402 20177 9178
rect 20211 8402 20223 9178
rect 20165 8390 20223 8402
rect 20423 9178 20481 9190
rect 20423 8402 20435 9178
rect 20469 8402 20481 9178
rect 20423 8390 20481 8402
rect 20537 9178 20595 9190
rect 20537 8402 20549 9178
rect 20583 8402 20595 9178
rect 20537 8390 20595 8402
rect 20795 9178 20853 9190
rect 20795 8402 20807 9178
rect 20841 8402 20853 9178
rect 20795 8390 20853 8402
rect 20909 9178 20967 9190
rect 20909 8402 20921 9178
rect 20955 8402 20967 9178
rect 20909 8390 20967 8402
rect 21167 9178 21225 9190
rect 21167 8402 21179 9178
rect 21213 8402 21225 9178
rect 21167 8390 21225 8402
rect 21281 9178 21339 9190
rect 21281 8402 21293 9178
rect 21327 8402 21339 9178
rect 21281 8390 21339 8402
rect 21539 9178 21597 9190
rect 21539 8402 21551 9178
rect 21585 8402 21597 9178
rect 21539 8390 21597 8402
rect 21653 9178 21711 9190
rect 21653 8402 21665 9178
rect 21699 8402 21711 9178
rect 21653 8390 21711 8402
rect 21911 9178 21969 9190
rect 21911 8402 21923 9178
rect 21957 8402 21969 9178
rect 21911 8390 21969 8402
rect 22025 9178 22083 9190
rect 22025 8402 22037 9178
rect 22071 8402 22083 9178
rect 22025 8390 22083 8402
rect 22283 9178 22341 9190
rect 22283 8402 22295 9178
rect 22329 8402 22341 9178
rect 22283 8390 22341 8402
rect 22397 9178 22455 9190
rect 22397 8402 22409 9178
rect 22443 8402 22455 9178
rect 22397 8390 22455 8402
rect 22655 9178 22713 9190
rect 22655 8402 22667 9178
rect 22701 8402 22713 9178
rect 22655 8390 22713 8402
rect 22769 9178 22827 9190
rect 22769 8402 22781 9178
rect 22815 8402 22827 9178
rect 22769 8390 22827 8402
rect 23027 9178 23085 9190
rect 23027 8402 23039 9178
rect 23073 8402 23085 9178
rect 23027 8390 23085 8402
rect 20165 8142 20223 8154
rect 20165 7366 20177 8142
rect 20211 7366 20223 8142
rect 20165 7354 20223 7366
rect 20423 8142 20481 8154
rect 20423 7366 20435 8142
rect 20469 7366 20481 8142
rect 20423 7354 20481 7366
rect 20537 8142 20595 8154
rect 20537 7366 20549 8142
rect 20583 7366 20595 8142
rect 20537 7354 20595 7366
rect 20795 8142 20853 8154
rect 20795 7366 20807 8142
rect 20841 7366 20853 8142
rect 20795 7354 20853 7366
rect 20909 8142 20967 8154
rect 20909 7366 20921 8142
rect 20955 7366 20967 8142
rect 20909 7354 20967 7366
rect 21167 8142 21225 8154
rect 21167 7366 21179 8142
rect 21213 7366 21225 8142
rect 21167 7354 21225 7366
rect 21281 8142 21339 8154
rect 21281 7366 21293 8142
rect 21327 7366 21339 8142
rect 21281 7354 21339 7366
rect 21539 8142 21597 8154
rect 21539 7366 21551 8142
rect 21585 7366 21597 8142
rect 21539 7354 21597 7366
rect 21653 8142 21711 8154
rect 21653 7366 21665 8142
rect 21699 7366 21711 8142
rect 21653 7354 21711 7366
rect 21911 8142 21969 8154
rect 21911 7366 21923 8142
rect 21957 7366 21969 8142
rect 21911 7354 21969 7366
rect 22025 8142 22083 8154
rect 22025 7366 22037 8142
rect 22071 7366 22083 8142
rect 22025 7354 22083 7366
rect 22283 8142 22341 8154
rect 22283 7366 22295 8142
rect 22329 7366 22341 8142
rect 22283 7354 22341 7366
rect 22397 8142 22455 8154
rect 22397 7366 22409 8142
rect 22443 7366 22455 8142
rect 22397 7354 22455 7366
rect 22655 8142 22713 8154
rect 22655 7366 22667 8142
rect 22701 7366 22713 8142
rect 22655 7354 22713 7366
rect 22769 8142 22827 8154
rect 22769 7366 22781 8142
rect 22815 7366 22827 8142
rect 22769 7354 22827 7366
rect 23027 8142 23085 8154
rect 23027 7366 23039 8142
rect 23073 7366 23085 8142
rect 23027 7354 23085 7366
rect 20165 7106 20223 7118
rect 20165 6330 20177 7106
rect 20211 6330 20223 7106
rect 20165 6318 20223 6330
rect 20423 7106 20481 7118
rect 20423 6330 20435 7106
rect 20469 6330 20481 7106
rect 20423 6318 20481 6330
rect 20537 7106 20595 7118
rect 20537 6330 20549 7106
rect 20583 6330 20595 7106
rect 20537 6318 20595 6330
rect 20795 7106 20853 7118
rect 20795 6330 20807 7106
rect 20841 6330 20853 7106
rect 20795 6318 20853 6330
rect 20909 7106 20967 7118
rect 20909 6330 20921 7106
rect 20955 6330 20967 7106
rect 20909 6318 20967 6330
rect 21167 7106 21225 7118
rect 21167 6330 21179 7106
rect 21213 6330 21225 7106
rect 21167 6318 21225 6330
rect 21281 7106 21339 7118
rect 21281 6330 21293 7106
rect 21327 6330 21339 7106
rect 21281 6318 21339 6330
rect 21539 7106 21597 7118
rect 21539 6330 21551 7106
rect 21585 6330 21597 7106
rect 21539 6318 21597 6330
rect 21653 7106 21711 7118
rect 21653 6330 21665 7106
rect 21699 6330 21711 7106
rect 21653 6318 21711 6330
rect 21911 7106 21969 7118
rect 21911 6330 21923 7106
rect 21957 6330 21969 7106
rect 21911 6318 21969 6330
rect 22025 7106 22083 7118
rect 22025 6330 22037 7106
rect 22071 6330 22083 7106
rect 22025 6318 22083 6330
rect 22283 7106 22341 7118
rect 22283 6330 22295 7106
rect 22329 6330 22341 7106
rect 22283 6318 22341 6330
rect 22397 7106 22455 7118
rect 22397 6330 22409 7106
rect 22443 6330 22455 7106
rect 22397 6318 22455 6330
rect 22655 7106 22713 7118
rect 22655 6330 22667 7106
rect 22701 6330 22713 7106
rect 22655 6318 22713 6330
rect 22769 7106 22827 7118
rect 22769 6330 22781 7106
rect 22815 6330 22827 7106
rect 22769 6318 22827 6330
rect 23027 7106 23085 7118
rect 23027 6330 23039 7106
rect 23073 6330 23085 7106
rect 23027 6318 23085 6330
rect 20165 6070 20223 6082
rect 20165 5294 20177 6070
rect 20211 5294 20223 6070
rect 20165 5282 20223 5294
rect 20423 6070 20481 6082
rect 20423 5294 20435 6070
rect 20469 5294 20481 6070
rect 20423 5282 20481 5294
rect 20537 6070 20595 6082
rect 20537 5294 20549 6070
rect 20583 5294 20595 6070
rect 20537 5282 20595 5294
rect 20795 6070 20853 6082
rect 20795 5294 20807 6070
rect 20841 5294 20853 6070
rect 20795 5282 20853 5294
rect 20909 6070 20967 6082
rect 20909 5294 20921 6070
rect 20955 5294 20967 6070
rect 20909 5282 20967 5294
rect 21167 6070 21225 6082
rect 21167 5294 21179 6070
rect 21213 5294 21225 6070
rect 21167 5282 21225 5294
rect 21281 6070 21339 6082
rect 21281 5294 21293 6070
rect 21327 5294 21339 6070
rect 21281 5282 21339 5294
rect 21539 6070 21597 6082
rect 21539 5294 21551 6070
rect 21585 5294 21597 6070
rect 21539 5282 21597 5294
rect 21653 6070 21711 6082
rect 21653 5294 21665 6070
rect 21699 5294 21711 6070
rect 21653 5282 21711 5294
rect 21911 6070 21969 6082
rect 21911 5294 21923 6070
rect 21957 5294 21969 6070
rect 21911 5282 21969 5294
rect 22025 6070 22083 6082
rect 22025 5294 22037 6070
rect 22071 5294 22083 6070
rect 22025 5282 22083 5294
rect 22283 6070 22341 6082
rect 22283 5294 22295 6070
rect 22329 5294 22341 6070
rect 22283 5282 22341 5294
rect 22397 6070 22455 6082
rect 22397 5294 22409 6070
rect 22443 5294 22455 6070
rect 22397 5282 22455 5294
rect 22655 6070 22713 6082
rect 22655 5294 22667 6070
rect 22701 5294 22713 6070
rect 22655 5282 22713 5294
rect 22769 6070 22827 6082
rect 22769 5294 22781 6070
rect 22815 5294 22827 6070
rect 22769 5282 22827 5294
rect 23027 6070 23085 6082
rect 23027 5294 23039 6070
rect 23073 5294 23085 6070
rect 23027 5282 23085 5294
<< ndiffc >>
rect 20177 4317 20211 4493
rect 20435 4317 20469 4493
rect 20549 4317 20583 4493
rect 20807 4317 20841 4493
rect 20921 4317 20955 4493
rect 21179 4317 21213 4493
rect 21293 4317 21327 4493
rect 21551 4317 21585 4493
rect 21665 4317 21699 4493
rect 21923 4317 21957 4493
rect 22037 4317 22071 4493
rect 22295 4317 22329 4493
rect 22409 4317 22443 4493
rect 22667 4317 22701 4493
rect 22781 4317 22815 4493
rect 23039 4317 23073 4493
rect 23153 4317 23187 4493
rect 23411 4317 23445 4493
rect 23525 4317 23559 4493
rect 23783 4317 23817 4493
rect 23897 4317 23931 4493
rect 24155 4317 24189 4493
rect 24269 4317 24303 4493
rect 24527 4317 24561 4493
rect 24641 4317 24675 4493
rect 24899 4317 24933 4493
rect 25013 4317 25047 4493
rect 25271 4317 25305 4493
rect 25385 4317 25419 4493
rect 25643 4317 25677 4493
rect 25757 4317 25791 4493
rect 26015 4317 26049 4493
rect 26129 4317 26163 4493
rect 26387 4317 26421 4493
rect 26501 4317 26535 4493
rect 26759 4317 26793 4493
rect 26873 4317 26907 4493
rect 27131 4317 27165 4493
rect 27245 4317 27279 4493
rect 27503 4317 27537 4493
rect 27617 4317 27651 4493
rect 27875 4317 27909 4493
rect 27989 4317 28023 4493
rect 28247 4317 28281 4493
rect 28361 4317 28395 4493
rect 28619 4317 28653 4493
rect 28733 4317 28767 4493
rect 28991 4317 29025 4493
rect 20177 3899 20211 4075
rect 20435 3899 20469 4075
rect 20549 3899 20583 4075
rect 20807 3899 20841 4075
rect 20921 3899 20955 4075
rect 21179 3899 21213 4075
rect 21293 3899 21327 4075
rect 21551 3899 21585 4075
rect 21665 3899 21699 4075
rect 21923 3899 21957 4075
rect 22037 3899 22071 4075
rect 22295 3899 22329 4075
rect 22409 3899 22443 4075
rect 22667 3899 22701 4075
rect 22781 3899 22815 4075
rect 23039 3899 23073 4075
rect 23153 3899 23187 4075
rect 23411 3899 23445 4075
rect 23525 3899 23559 4075
rect 23783 3899 23817 4075
rect 23897 3899 23931 4075
rect 24155 3899 24189 4075
rect 24269 3899 24303 4075
rect 24527 3899 24561 4075
rect 24641 3899 24675 4075
rect 24899 3899 24933 4075
rect 25013 3899 25047 4075
rect 25271 3899 25305 4075
rect 25385 3899 25419 4075
rect 25643 3899 25677 4075
rect 25757 3899 25791 4075
rect 26015 3899 26049 4075
rect 26129 3899 26163 4075
rect 26387 3899 26421 4075
rect 26501 3899 26535 4075
rect 26759 3899 26793 4075
rect 26873 3899 26907 4075
rect 27131 3899 27165 4075
rect 27245 3899 27279 4075
rect 27503 3899 27537 4075
rect 27617 3899 27651 4075
rect 27875 3899 27909 4075
rect 27989 3899 28023 4075
rect 28247 3899 28281 4075
rect 28361 3899 28395 4075
rect 28619 3899 28653 4075
rect 28733 3899 28767 4075
rect 28991 3899 29025 4075
rect 20177 3481 20211 3657
rect 20435 3481 20469 3657
rect 20549 3481 20583 3657
rect 20807 3481 20841 3657
rect 20921 3481 20955 3657
rect 21179 3481 21213 3657
rect 21293 3481 21327 3657
rect 21551 3481 21585 3657
rect 21665 3481 21699 3657
rect 21923 3481 21957 3657
rect 22037 3481 22071 3657
rect 22295 3481 22329 3657
rect 22409 3481 22443 3657
rect 22667 3481 22701 3657
rect 22781 3481 22815 3657
rect 23039 3481 23073 3657
rect 23153 3481 23187 3657
rect 23411 3481 23445 3657
rect 23525 3481 23559 3657
rect 23783 3481 23817 3657
rect 23897 3481 23931 3657
rect 24155 3481 24189 3657
rect 24269 3481 24303 3657
rect 24527 3481 24561 3657
rect 24641 3481 24675 3657
rect 24899 3481 24933 3657
rect 25013 3481 25047 3657
rect 25271 3481 25305 3657
rect 25385 3481 25419 3657
rect 25643 3481 25677 3657
rect 25757 3481 25791 3657
rect 26015 3481 26049 3657
rect 26129 3481 26163 3657
rect 26387 3481 26421 3657
rect 26501 3481 26535 3657
rect 26759 3481 26793 3657
rect 26873 3481 26907 3657
rect 27131 3481 27165 3657
rect 27245 3481 27279 3657
rect 27503 3481 27537 3657
rect 27617 3481 27651 3657
rect 27875 3481 27909 3657
rect 27989 3481 28023 3657
rect 28247 3481 28281 3657
rect 28361 3481 28395 3657
rect 28619 3481 28653 3657
rect 28733 3481 28767 3657
rect 28991 3481 29025 3657
rect 20177 3063 20211 3239
rect 20435 3063 20469 3239
rect 20549 3063 20583 3239
rect 20807 3063 20841 3239
rect 20921 3063 20955 3239
rect 21179 3063 21213 3239
rect 21293 3063 21327 3239
rect 21551 3063 21585 3239
rect 21665 3063 21699 3239
rect 21923 3063 21957 3239
rect 22037 3063 22071 3239
rect 22295 3063 22329 3239
rect 22409 3063 22443 3239
rect 22667 3063 22701 3239
rect 22781 3063 22815 3239
rect 23039 3063 23073 3239
rect 23153 3063 23187 3239
rect 23411 3063 23445 3239
rect 23525 3063 23559 3239
rect 23783 3063 23817 3239
rect 23897 3063 23931 3239
rect 24155 3063 24189 3239
rect 24269 3063 24303 3239
rect 24527 3063 24561 3239
rect 24641 3063 24675 3239
rect 24899 3063 24933 3239
rect 25013 3063 25047 3239
rect 25271 3063 25305 3239
rect 25385 3063 25419 3239
rect 25643 3063 25677 3239
rect 25757 3063 25791 3239
rect 26015 3063 26049 3239
rect 26129 3063 26163 3239
rect 26387 3063 26421 3239
rect 26501 3063 26535 3239
rect 26759 3063 26793 3239
rect 26873 3063 26907 3239
rect 27131 3063 27165 3239
rect 27245 3063 27279 3239
rect 27503 3063 27537 3239
rect 27617 3063 27651 3239
rect 27875 3063 27909 3239
rect 27989 3063 28023 3239
rect 28247 3063 28281 3239
rect 28361 3063 28395 3239
rect 28619 3063 28653 3239
rect 28733 3063 28767 3239
rect 28991 3063 29025 3239
<< pdiffc >>
rect 18689 11190 18723 11566
rect 18947 11190 18981 11566
rect 19061 11190 19095 11566
rect 19319 11190 19353 11566
rect 19433 11190 19467 11566
rect 19691 11190 19725 11566
rect 19805 11190 19839 11566
rect 20063 11190 20097 11566
rect 20177 11190 20211 11566
rect 20435 11190 20469 11566
rect 20549 11190 20583 11566
rect 20807 11190 20841 11566
rect 20921 11190 20955 11566
rect 21179 11190 21213 11566
rect 21293 11190 21327 11566
rect 21551 11190 21585 11566
rect 21665 11190 21699 11566
rect 21923 11190 21957 11566
rect 22037 11190 22071 11566
rect 22295 11190 22329 11566
rect 22409 11190 22443 11566
rect 22667 11190 22701 11566
rect 22781 11190 22815 11566
rect 23039 11190 23073 11566
rect 23153 11190 23187 11566
rect 23411 11190 23445 11566
rect 23525 11190 23559 11566
rect 23783 11190 23817 11566
rect 23897 11190 23931 11566
rect 24155 11190 24189 11566
rect 24269 11190 24303 11566
rect 24527 11190 24561 11566
rect 24641 11190 24675 11566
rect 24899 11190 24933 11566
rect 25013 11190 25047 11566
rect 25271 11190 25305 11566
rect 25385 11190 25419 11566
rect 25643 11190 25677 11566
rect 25757 11190 25791 11566
rect 26015 11190 26049 11566
rect 26129 11190 26163 11566
rect 26387 11190 26421 11566
rect 26501 11190 26535 11566
rect 26759 11190 26793 11566
rect 26873 11190 26907 11566
rect 27131 11190 27165 11566
rect 27245 11190 27279 11566
rect 27503 11190 27537 11566
rect 27617 11190 27651 11566
rect 27875 11190 27909 11566
rect 27989 11190 28023 11566
rect 28247 11190 28281 11566
rect 28361 11190 28395 11566
rect 28619 11190 28653 11566
rect 28733 11190 28767 11566
rect 28991 11190 29025 11566
rect 29105 11190 29139 11566
rect 29363 11190 29397 11566
rect 29477 11190 29511 11566
rect 29735 11190 29769 11566
rect 29849 11190 29883 11566
rect 30107 11190 30141 11566
rect 30221 11190 30255 11566
rect 30479 11190 30513 11566
rect 18689 10554 18723 10930
rect 18947 10554 18981 10930
rect 19061 10554 19095 10930
rect 19319 10554 19353 10930
rect 19433 10554 19467 10930
rect 19691 10554 19725 10930
rect 19805 10554 19839 10930
rect 20063 10554 20097 10930
rect 20177 10554 20211 10930
rect 20435 10554 20469 10930
rect 20549 10554 20583 10930
rect 20807 10554 20841 10930
rect 20921 10554 20955 10930
rect 21179 10554 21213 10930
rect 21293 10554 21327 10930
rect 21551 10554 21585 10930
rect 21665 10554 21699 10930
rect 21923 10554 21957 10930
rect 22037 10554 22071 10930
rect 22295 10554 22329 10930
rect 22409 10554 22443 10930
rect 22667 10554 22701 10930
rect 22781 10554 22815 10930
rect 23039 10554 23073 10930
rect 23153 10554 23187 10930
rect 23411 10554 23445 10930
rect 23525 10554 23559 10930
rect 23783 10554 23817 10930
rect 23897 10554 23931 10930
rect 24155 10554 24189 10930
rect 24269 10554 24303 10930
rect 24527 10554 24561 10930
rect 24641 10554 24675 10930
rect 24899 10554 24933 10930
rect 25013 10554 25047 10930
rect 25271 10554 25305 10930
rect 25385 10554 25419 10930
rect 25643 10554 25677 10930
rect 25757 10554 25791 10930
rect 26015 10554 26049 10930
rect 26129 10554 26163 10930
rect 26387 10554 26421 10930
rect 26501 10554 26535 10930
rect 26759 10554 26793 10930
rect 26873 10554 26907 10930
rect 27131 10554 27165 10930
rect 27245 10554 27279 10930
rect 27503 10554 27537 10930
rect 27617 10554 27651 10930
rect 27875 10554 27909 10930
rect 27989 10554 28023 10930
rect 28247 10554 28281 10930
rect 28361 10554 28395 10930
rect 28619 10554 28653 10930
rect 28733 10554 28767 10930
rect 28991 10554 29025 10930
rect 29105 10554 29139 10930
rect 29363 10554 29397 10930
rect 29477 10554 29511 10930
rect 29735 10554 29769 10930
rect 29849 10554 29883 10930
rect 30107 10554 30141 10930
rect 30221 10554 30255 10930
rect 30479 10554 30513 10930
rect 18689 9918 18723 10294
rect 18947 9918 18981 10294
rect 19061 9918 19095 10294
rect 19319 9918 19353 10294
rect 19433 9918 19467 10294
rect 19691 9918 19725 10294
rect 19805 9918 19839 10294
rect 20063 9918 20097 10294
rect 20177 9918 20211 10294
rect 20435 9918 20469 10294
rect 20549 9918 20583 10294
rect 20807 9918 20841 10294
rect 20921 9918 20955 10294
rect 21179 9918 21213 10294
rect 21293 9918 21327 10294
rect 21551 9918 21585 10294
rect 21665 9918 21699 10294
rect 21923 9918 21957 10294
rect 22037 9918 22071 10294
rect 22295 9918 22329 10294
rect 22409 9918 22443 10294
rect 22667 9918 22701 10294
rect 22781 9918 22815 10294
rect 23039 9918 23073 10294
rect 23153 9918 23187 10294
rect 23411 9918 23445 10294
rect 23525 9918 23559 10294
rect 23783 9918 23817 10294
rect 23897 9918 23931 10294
rect 24155 9918 24189 10294
rect 24269 9918 24303 10294
rect 24527 9918 24561 10294
rect 24641 9918 24675 10294
rect 24899 9918 24933 10294
rect 25013 9918 25047 10294
rect 25271 9918 25305 10294
rect 25385 9918 25419 10294
rect 25643 9918 25677 10294
rect 25757 9918 25791 10294
rect 26015 9918 26049 10294
rect 26129 9918 26163 10294
rect 26387 9918 26421 10294
rect 26501 9918 26535 10294
rect 26759 9918 26793 10294
rect 26873 9918 26907 10294
rect 27131 9918 27165 10294
rect 27245 9918 27279 10294
rect 27503 9918 27537 10294
rect 27617 9918 27651 10294
rect 27875 9918 27909 10294
rect 27989 9918 28023 10294
rect 28247 9918 28281 10294
rect 28361 9918 28395 10294
rect 28619 9918 28653 10294
rect 28733 9918 28767 10294
rect 28991 9918 29025 10294
rect 29105 9918 29139 10294
rect 29363 9918 29397 10294
rect 29477 9918 29511 10294
rect 29735 9918 29769 10294
rect 29849 9918 29883 10294
rect 30107 9918 30141 10294
rect 30221 9918 30255 10294
rect 30479 9918 30513 10294
rect 20177 8402 20211 9178
rect 20435 8402 20469 9178
rect 20549 8402 20583 9178
rect 20807 8402 20841 9178
rect 20921 8402 20955 9178
rect 21179 8402 21213 9178
rect 21293 8402 21327 9178
rect 21551 8402 21585 9178
rect 21665 8402 21699 9178
rect 21923 8402 21957 9178
rect 22037 8402 22071 9178
rect 22295 8402 22329 9178
rect 22409 8402 22443 9178
rect 22667 8402 22701 9178
rect 22781 8402 22815 9178
rect 23039 8402 23073 9178
rect 20177 7366 20211 8142
rect 20435 7366 20469 8142
rect 20549 7366 20583 8142
rect 20807 7366 20841 8142
rect 20921 7366 20955 8142
rect 21179 7366 21213 8142
rect 21293 7366 21327 8142
rect 21551 7366 21585 8142
rect 21665 7366 21699 8142
rect 21923 7366 21957 8142
rect 22037 7366 22071 8142
rect 22295 7366 22329 8142
rect 22409 7366 22443 8142
rect 22667 7366 22701 8142
rect 22781 7366 22815 8142
rect 23039 7366 23073 8142
rect 20177 6330 20211 7106
rect 20435 6330 20469 7106
rect 20549 6330 20583 7106
rect 20807 6330 20841 7106
rect 20921 6330 20955 7106
rect 21179 6330 21213 7106
rect 21293 6330 21327 7106
rect 21551 6330 21585 7106
rect 21665 6330 21699 7106
rect 21923 6330 21957 7106
rect 22037 6330 22071 7106
rect 22295 6330 22329 7106
rect 22409 6330 22443 7106
rect 22667 6330 22701 7106
rect 22781 6330 22815 7106
rect 23039 6330 23073 7106
rect 20177 5294 20211 6070
rect 20435 5294 20469 6070
rect 20549 5294 20583 6070
rect 20807 5294 20841 6070
rect 20921 5294 20955 6070
rect 21179 5294 21213 6070
rect 21293 5294 21327 6070
rect 21551 5294 21585 6070
rect 21665 5294 21699 6070
rect 21923 5294 21957 6070
rect 22037 5294 22071 6070
rect 22295 5294 22329 6070
rect 22409 5294 22443 6070
rect 22667 5294 22701 6070
rect 22781 5294 22815 6070
rect 23039 5294 23073 6070
<< psubdiff >>
rect 23689 7425 23785 7459
rect 23923 7425 24019 7459
rect 23689 7363 23723 7425
rect 23985 7363 24019 7425
rect 23689 5809 23723 5871
rect 23985 5809 24019 5871
rect 23689 5775 23785 5809
rect 23923 5775 24019 5809
rect 20063 4645 20159 4679
rect 29043 4645 29139 4679
rect 20063 4583 20097 4645
rect 29105 4583 29139 4645
rect 20063 2911 20097 2973
rect 29105 2911 29139 2973
rect 20063 2877 20159 2911
rect 29043 2877 29139 2911
<< nsubdiff >>
rect 18575 11727 18671 11761
rect 30531 11727 30627 11761
rect 18575 11665 18609 11727
rect 30593 11665 30627 11727
rect 18575 9757 18609 9819
rect 30593 9757 30627 9819
rect 18575 9723 18671 9757
rect 30531 9723 30627 9757
rect 20063 9339 20159 9373
rect 23091 9339 23187 9373
rect 20063 9277 20097 9339
rect 23153 9277 23187 9339
rect 20063 5133 20097 5195
rect 23153 5133 23187 5195
rect 20063 5099 20159 5133
rect 23091 5099 23187 5133
<< psubdiffcont >>
rect 23785 7425 23923 7459
rect 23689 5871 23723 7363
rect 23985 5871 24019 7363
rect 23785 5775 23923 5809
rect 20159 4645 29043 4679
rect 20063 2973 20097 4583
rect 29105 2973 29139 4583
rect 20159 2877 29043 2911
<< nsubdiffcont >>
rect 18671 11727 30531 11761
rect 18575 9819 18609 11665
rect 30593 9819 30627 11665
rect 18671 9723 30531 9757
rect 20159 9339 23091 9373
rect 20063 5195 20097 9277
rect 23153 5195 23187 9277
rect 20159 5099 23091 5133
<< poly >>
rect 18735 11659 18935 11675
rect 18735 11625 18751 11659
rect 18919 11625 18935 11659
rect 18735 11578 18935 11625
rect 19107 11659 19307 11675
rect 19107 11625 19123 11659
rect 19291 11625 19307 11659
rect 19107 11578 19307 11625
rect 19479 11659 19679 11675
rect 19479 11625 19495 11659
rect 19663 11625 19679 11659
rect 19479 11578 19679 11625
rect 19851 11659 20051 11675
rect 19851 11625 19867 11659
rect 20035 11625 20051 11659
rect 19851 11578 20051 11625
rect 20223 11659 20423 11675
rect 20223 11625 20239 11659
rect 20407 11625 20423 11659
rect 20223 11578 20423 11625
rect 20595 11659 20795 11675
rect 20595 11625 20611 11659
rect 20779 11625 20795 11659
rect 20595 11578 20795 11625
rect 20967 11659 21167 11675
rect 20967 11625 20983 11659
rect 21151 11625 21167 11659
rect 20967 11578 21167 11625
rect 21339 11659 21539 11675
rect 21339 11625 21355 11659
rect 21523 11625 21539 11659
rect 21339 11578 21539 11625
rect 21711 11659 21911 11675
rect 21711 11625 21727 11659
rect 21895 11625 21911 11659
rect 21711 11578 21911 11625
rect 22083 11659 22283 11675
rect 22083 11625 22099 11659
rect 22267 11625 22283 11659
rect 22083 11578 22283 11625
rect 22455 11659 22655 11675
rect 22455 11625 22471 11659
rect 22639 11625 22655 11659
rect 22455 11578 22655 11625
rect 22827 11659 23027 11675
rect 22827 11625 22843 11659
rect 23011 11625 23027 11659
rect 22827 11578 23027 11625
rect 23199 11659 23399 11675
rect 23199 11625 23215 11659
rect 23383 11625 23399 11659
rect 23199 11578 23399 11625
rect 23571 11659 23771 11675
rect 23571 11625 23587 11659
rect 23755 11625 23771 11659
rect 23571 11578 23771 11625
rect 23943 11659 24143 11675
rect 23943 11625 23959 11659
rect 24127 11625 24143 11659
rect 23943 11578 24143 11625
rect 24315 11659 24515 11675
rect 24315 11625 24331 11659
rect 24499 11625 24515 11659
rect 24315 11578 24515 11625
rect 24687 11659 24887 11675
rect 24687 11625 24703 11659
rect 24871 11625 24887 11659
rect 24687 11578 24887 11625
rect 25059 11659 25259 11675
rect 25059 11625 25075 11659
rect 25243 11625 25259 11659
rect 25059 11578 25259 11625
rect 25431 11659 25631 11675
rect 25431 11625 25447 11659
rect 25615 11625 25631 11659
rect 25431 11578 25631 11625
rect 25803 11659 26003 11675
rect 25803 11625 25819 11659
rect 25987 11625 26003 11659
rect 25803 11578 26003 11625
rect 26175 11659 26375 11675
rect 26175 11625 26191 11659
rect 26359 11625 26375 11659
rect 26175 11578 26375 11625
rect 26547 11659 26747 11675
rect 26547 11625 26563 11659
rect 26731 11625 26747 11659
rect 26547 11578 26747 11625
rect 26919 11659 27119 11675
rect 26919 11625 26935 11659
rect 27103 11625 27119 11659
rect 26919 11578 27119 11625
rect 27291 11659 27491 11675
rect 27291 11625 27307 11659
rect 27475 11625 27491 11659
rect 27291 11578 27491 11625
rect 27663 11659 27863 11675
rect 27663 11625 27679 11659
rect 27847 11625 27863 11659
rect 27663 11578 27863 11625
rect 28035 11659 28235 11675
rect 28035 11625 28051 11659
rect 28219 11625 28235 11659
rect 28035 11578 28235 11625
rect 28407 11659 28607 11675
rect 28407 11625 28423 11659
rect 28591 11625 28607 11659
rect 28407 11578 28607 11625
rect 28779 11659 28979 11675
rect 28779 11625 28795 11659
rect 28963 11625 28979 11659
rect 28779 11578 28979 11625
rect 29151 11659 29351 11675
rect 29151 11625 29167 11659
rect 29335 11625 29351 11659
rect 29151 11578 29351 11625
rect 29523 11659 29723 11675
rect 29523 11625 29539 11659
rect 29707 11625 29723 11659
rect 29523 11578 29723 11625
rect 29895 11659 30095 11675
rect 29895 11625 29911 11659
rect 30079 11625 30095 11659
rect 29895 11578 30095 11625
rect 30267 11659 30467 11675
rect 30267 11625 30283 11659
rect 30451 11625 30467 11659
rect 30267 11578 30467 11625
rect 18735 11131 18935 11178
rect 18735 11097 18751 11131
rect 18919 11097 18935 11131
rect 18735 11081 18935 11097
rect 19107 11131 19307 11178
rect 19107 11097 19123 11131
rect 19291 11097 19307 11131
rect 19107 11081 19307 11097
rect 19479 11131 19679 11178
rect 19479 11097 19495 11131
rect 19663 11097 19679 11131
rect 19479 11081 19679 11097
rect 19851 11131 20051 11178
rect 19851 11097 19867 11131
rect 20035 11097 20051 11131
rect 19851 11081 20051 11097
rect 20223 11131 20423 11178
rect 20223 11097 20239 11131
rect 20407 11097 20423 11131
rect 20223 11081 20423 11097
rect 20595 11131 20795 11178
rect 20595 11097 20611 11131
rect 20779 11097 20795 11131
rect 20595 11081 20795 11097
rect 20967 11131 21167 11178
rect 20967 11097 20983 11131
rect 21151 11097 21167 11131
rect 20967 11081 21167 11097
rect 21339 11131 21539 11178
rect 21339 11097 21355 11131
rect 21523 11097 21539 11131
rect 21339 11081 21539 11097
rect 21711 11131 21911 11178
rect 21711 11097 21727 11131
rect 21895 11097 21911 11131
rect 21711 11081 21911 11097
rect 22083 11131 22283 11178
rect 22083 11097 22099 11131
rect 22267 11097 22283 11131
rect 22083 11081 22283 11097
rect 22455 11131 22655 11178
rect 22455 11097 22471 11131
rect 22639 11097 22655 11131
rect 22455 11081 22655 11097
rect 22827 11131 23027 11178
rect 22827 11097 22843 11131
rect 23011 11097 23027 11131
rect 22827 11081 23027 11097
rect 23199 11131 23399 11178
rect 23199 11097 23215 11131
rect 23383 11097 23399 11131
rect 23199 11081 23399 11097
rect 23571 11131 23771 11178
rect 23571 11097 23587 11131
rect 23755 11097 23771 11131
rect 23571 11081 23771 11097
rect 23943 11131 24143 11178
rect 23943 11097 23959 11131
rect 24127 11097 24143 11131
rect 23943 11081 24143 11097
rect 24315 11131 24515 11178
rect 24315 11097 24331 11131
rect 24499 11097 24515 11131
rect 24315 11081 24515 11097
rect 24687 11131 24887 11178
rect 24687 11097 24703 11131
rect 24871 11097 24887 11131
rect 24687 11081 24887 11097
rect 25059 11131 25259 11178
rect 25059 11097 25075 11131
rect 25243 11097 25259 11131
rect 25059 11081 25259 11097
rect 25431 11131 25631 11178
rect 25431 11097 25447 11131
rect 25615 11097 25631 11131
rect 25431 11081 25631 11097
rect 25803 11131 26003 11178
rect 25803 11097 25819 11131
rect 25987 11097 26003 11131
rect 25803 11081 26003 11097
rect 26175 11131 26375 11178
rect 26175 11097 26191 11131
rect 26359 11097 26375 11131
rect 26175 11081 26375 11097
rect 26547 11131 26747 11178
rect 26547 11097 26563 11131
rect 26731 11097 26747 11131
rect 26547 11081 26747 11097
rect 26919 11131 27119 11178
rect 26919 11097 26935 11131
rect 27103 11097 27119 11131
rect 26919 11081 27119 11097
rect 27291 11131 27491 11178
rect 27291 11097 27307 11131
rect 27475 11097 27491 11131
rect 27291 11081 27491 11097
rect 27663 11131 27863 11178
rect 27663 11097 27679 11131
rect 27847 11097 27863 11131
rect 27663 11081 27863 11097
rect 28035 11131 28235 11178
rect 28035 11097 28051 11131
rect 28219 11097 28235 11131
rect 28035 11081 28235 11097
rect 28407 11131 28607 11178
rect 28407 11097 28423 11131
rect 28591 11097 28607 11131
rect 28407 11081 28607 11097
rect 28779 11131 28979 11178
rect 28779 11097 28795 11131
rect 28963 11097 28979 11131
rect 28779 11081 28979 11097
rect 29151 11131 29351 11178
rect 29151 11097 29167 11131
rect 29335 11097 29351 11131
rect 29151 11081 29351 11097
rect 29523 11131 29723 11178
rect 29523 11097 29539 11131
rect 29707 11097 29723 11131
rect 29523 11081 29723 11097
rect 29895 11131 30095 11178
rect 29895 11097 29911 11131
rect 30079 11097 30095 11131
rect 29895 11081 30095 11097
rect 30267 11131 30467 11178
rect 30267 11097 30283 11131
rect 30451 11097 30467 11131
rect 30267 11081 30467 11097
rect 18735 11023 18935 11039
rect 18735 10989 18751 11023
rect 18919 10989 18935 11023
rect 18735 10942 18935 10989
rect 19107 11023 19307 11039
rect 19107 10989 19123 11023
rect 19291 10989 19307 11023
rect 19107 10942 19307 10989
rect 19479 11023 19679 11039
rect 19479 10989 19495 11023
rect 19663 10989 19679 11023
rect 19479 10942 19679 10989
rect 19851 11023 20051 11039
rect 19851 10989 19867 11023
rect 20035 10989 20051 11023
rect 19851 10942 20051 10989
rect 20223 11023 20423 11039
rect 20223 10989 20239 11023
rect 20407 10989 20423 11023
rect 20223 10942 20423 10989
rect 20595 11023 20795 11039
rect 20595 10989 20611 11023
rect 20779 10989 20795 11023
rect 20595 10942 20795 10989
rect 20967 11023 21167 11039
rect 20967 10989 20983 11023
rect 21151 10989 21167 11023
rect 20967 10942 21167 10989
rect 21339 11023 21539 11039
rect 21339 10989 21355 11023
rect 21523 10989 21539 11023
rect 21339 10942 21539 10989
rect 21711 11023 21911 11039
rect 21711 10989 21727 11023
rect 21895 10989 21911 11023
rect 21711 10942 21911 10989
rect 22083 11023 22283 11039
rect 22083 10989 22099 11023
rect 22267 10989 22283 11023
rect 22083 10942 22283 10989
rect 22455 11023 22655 11039
rect 22455 10989 22471 11023
rect 22639 10989 22655 11023
rect 22455 10942 22655 10989
rect 22827 11023 23027 11039
rect 22827 10989 22843 11023
rect 23011 10989 23027 11023
rect 22827 10942 23027 10989
rect 23199 11023 23399 11039
rect 23199 10989 23215 11023
rect 23383 10989 23399 11023
rect 23199 10942 23399 10989
rect 23571 11023 23771 11039
rect 23571 10989 23587 11023
rect 23755 10989 23771 11023
rect 23571 10942 23771 10989
rect 23943 11023 24143 11039
rect 23943 10989 23959 11023
rect 24127 10989 24143 11023
rect 23943 10942 24143 10989
rect 24315 11023 24515 11039
rect 24315 10989 24331 11023
rect 24499 10989 24515 11023
rect 24315 10942 24515 10989
rect 24687 11023 24887 11039
rect 24687 10989 24703 11023
rect 24871 10989 24887 11023
rect 24687 10942 24887 10989
rect 25059 11023 25259 11039
rect 25059 10989 25075 11023
rect 25243 10989 25259 11023
rect 25059 10942 25259 10989
rect 25431 11023 25631 11039
rect 25431 10989 25447 11023
rect 25615 10989 25631 11023
rect 25431 10942 25631 10989
rect 25803 11023 26003 11039
rect 25803 10989 25819 11023
rect 25987 10989 26003 11023
rect 25803 10942 26003 10989
rect 26175 11023 26375 11039
rect 26175 10989 26191 11023
rect 26359 10989 26375 11023
rect 26175 10942 26375 10989
rect 26547 11023 26747 11039
rect 26547 10989 26563 11023
rect 26731 10989 26747 11023
rect 26547 10942 26747 10989
rect 26919 11023 27119 11039
rect 26919 10989 26935 11023
rect 27103 10989 27119 11023
rect 26919 10942 27119 10989
rect 27291 11023 27491 11039
rect 27291 10989 27307 11023
rect 27475 10989 27491 11023
rect 27291 10942 27491 10989
rect 27663 11023 27863 11039
rect 27663 10989 27679 11023
rect 27847 10989 27863 11023
rect 27663 10942 27863 10989
rect 28035 11023 28235 11039
rect 28035 10989 28051 11023
rect 28219 10989 28235 11023
rect 28035 10942 28235 10989
rect 28407 11023 28607 11039
rect 28407 10989 28423 11023
rect 28591 10989 28607 11023
rect 28407 10942 28607 10989
rect 28779 11023 28979 11039
rect 28779 10989 28795 11023
rect 28963 10989 28979 11023
rect 28779 10942 28979 10989
rect 29151 11023 29351 11039
rect 29151 10989 29167 11023
rect 29335 10989 29351 11023
rect 29151 10942 29351 10989
rect 29523 11023 29723 11039
rect 29523 10989 29539 11023
rect 29707 10989 29723 11023
rect 29523 10942 29723 10989
rect 29895 11023 30095 11039
rect 29895 10989 29911 11023
rect 30079 10989 30095 11023
rect 29895 10942 30095 10989
rect 30267 11023 30467 11039
rect 30267 10989 30283 11023
rect 30451 10989 30467 11023
rect 30267 10942 30467 10989
rect 18735 10495 18935 10542
rect 18735 10461 18751 10495
rect 18919 10461 18935 10495
rect 18735 10445 18935 10461
rect 19107 10495 19307 10542
rect 19107 10461 19123 10495
rect 19291 10461 19307 10495
rect 19107 10445 19307 10461
rect 19479 10495 19679 10542
rect 19479 10461 19495 10495
rect 19663 10461 19679 10495
rect 19479 10445 19679 10461
rect 19851 10495 20051 10542
rect 19851 10461 19867 10495
rect 20035 10461 20051 10495
rect 19851 10445 20051 10461
rect 20223 10495 20423 10542
rect 20223 10461 20239 10495
rect 20407 10461 20423 10495
rect 20223 10445 20423 10461
rect 20595 10495 20795 10542
rect 20595 10461 20611 10495
rect 20779 10461 20795 10495
rect 20595 10445 20795 10461
rect 20967 10495 21167 10542
rect 20967 10461 20983 10495
rect 21151 10461 21167 10495
rect 20967 10445 21167 10461
rect 21339 10495 21539 10542
rect 21339 10461 21355 10495
rect 21523 10461 21539 10495
rect 21339 10445 21539 10461
rect 21711 10495 21911 10542
rect 21711 10461 21727 10495
rect 21895 10461 21911 10495
rect 21711 10445 21911 10461
rect 22083 10495 22283 10542
rect 22083 10461 22099 10495
rect 22267 10461 22283 10495
rect 22083 10445 22283 10461
rect 22455 10495 22655 10542
rect 22455 10461 22471 10495
rect 22639 10461 22655 10495
rect 22455 10445 22655 10461
rect 22827 10495 23027 10542
rect 22827 10461 22843 10495
rect 23011 10461 23027 10495
rect 22827 10445 23027 10461
rect 23199 10495 23399 10542
rect 23199 10461 23215 10495
rect 23383 10461 23399 10495
rect 23199 10445 23399 10461
rect 23571 10495 23771 10542
rect 23571 10461 23587 10495
rect 23755 10461 23771 10495
rect 23571 10445 23771 10461
rect 23943 10495 24143 10542
rect 23943 10461 23959 10495
rect 24127 10461 24143 10495
rect 23943 10445 24143 10461
rect 24315 10495 24515 10542
rect 24315 10461 24331 10495
rect 24499 10461 24515 10495
rect 24315 10445 24515 10461
rect 24687 10495 24887 10542
rect 24687 10461 24703 10495
rect 24871 10461 24887 10495
rect 24687 10445 24887 10461
rect 25059 10495 25259 10542
rect 25059 10461 25075 10495
rect 25243 10461 25259 10495
rect 25059 10445 25259 10461
rect 25431 10495 25631 10542
rect 25431 10461 25447 10495
rect 25615 10461 25631 10495
rect 25431 10445 25631 10461
rect 25803 10495 26003 10542
rect 25803 10461 25819 10495
rect 25987 10461 26003 10495
rect 25803 10445 26003 10461
rect 26175 10495 26375 10542
rect 26175 10461 26191 10495
rect 26359 10461 26375 10495
rect 26175 10445 26375 10461
rect 26547 10495 26747 10542
rect 26547 10461 26563 10495
rect 26731 10461 26747 10495
rect 26547 10445 26747 10461
rect 26919 10495 27119 10542
rect 26919 10461 26935 10495
rect 27103 10461 27119 10495
rect 26919 10445 27119 10461
rect 27291 10495 27491 10542
rect 27291 10461 27307 10495
rect 27475 10461 27491 10495
rect 27291 10445 27491 10461
rect 27663 10495 27863 10542
rect 27663 10461 27679 10495
rect 27847 10461 27863 10495
rect 27663 10445 27863 10461
rect 28035 10495 28235 10542
rect 28035 10461 28051 10495
rect 28219 10461 28235 10495
rect 28035 10445 28235 10461
rect 28407 10495 28607 10542
rect 28407 10461 28423 10495
rect 28591 10461 28607 10495
rect 28407 10445 28607 10461
rect 28779 10495 28979 10542
rect 28779 10461 28795 10495
rect 28963 10461 28979 10495
rect 28779 10445 28979 10461
rect 29151 10495 29351 10542
rect 29151 10461 29167 10495
rect 29335 10461 29351 10495
rect 29151 10445 29351 10461
rect 29523 10495 29723 10542
rect 29523 10461 29539 10495
rect 29707 10461 29723 10495
rect 29523 10445 29723 10461
rect 29895 10495 30095 10542
rect 29895 10461 29911 10495
rect 30079 10461 30095 10495
rect 29895 10445 30095 10461
rect 30267 10495 30467 10542
rect 30267 10461 30283 10495
rect 30451 10461 30467 10495
rect 30267 10445 30467 10461
rect 18735 10387 18935 10403
rect 18735 10353 18751 10387
rect 18919 10353 18935 10387
rect 18735 10306 18935 10353
rect 19107 10387 19307 10403
rect 19107 10353 19123 10387
rect 19291 10353 19307 10387
rect 19107 10306 19307 10353
rect 19479 10387 19679 10403
rect 19479 10353 19495 10387
rect 19663 10353 19679 10387
rect 19479 10306 19679 10353
rect 19851 10387 20051 10403
rect 19851 10353 19867 10387
rect 20035 10353 20051 10387
rect 19851 10306 20051 10353
rect 20223 10387 20423 10403
rect 20223 10353 20239 10387
rect 20407 10353 20423 10387
rect 20223 10306 20423 10353
rect 20595 10387 20795 10403
rect 20595 10353 20611 10387
rect 20779 10353 20795 10387
rect 20595 10306 20795 10353
rect 20967 10387 21167 10403
rect 20967 10353 20983 10387
rect 21151 10353 21167 10387
rect 20967 10306 21167 10353
rect 21339 10387 21539 10403
rect 21339 10353 21355 10387
rect 21523 10353 21539 10387
rect 21339 10306 21539 10353
rect 21711 10387 21911 10403
rect 21711 10353 21727 10387
rect 21895 10353 21911 10387
rect 21711 10306 21911 10353
rect 22083 10387 22283 10403
rect 22083 10353 22099 10387
rect 22267 10353 22283 10387
rect 22083 10306 22283 10353
rect 22455 10387 22655 10403
rect 22455 10353 22471 10387
rect 22639 10353 22655 10387
rect 22455 10306 22655 10353
rect 22827 10387 23027 10403
rect 22827 10353 22843 10387
rect 23011 10353 23027 10387
rect 22827 10306 23027 10353
rect 23199 10387 23399 10403
rect 23199 10353 23215 10387
rect 23383 10353 23399 10387
rect 23199 10306 23399 10353
rect 23571 10387 23771 10403
rect 23571 10353 23587 10387
rect 23755 10353 23771 10387
rect 23571 10306 23771 10353
rect 23943 10387 24143 10403
rect 23943 10353 23959 10387
rect 24127 10353 24143 10387
rect 23943 10306 24143 10353
rect 24315 10387 24515 10403
rect 24315 10353 24331 10387
rect 24499 10353 24515 10387
rect 24315 10306 24515 10353
rect 24687 10387 24887 10403
rect 24687 10353 24703 10387
rect 24871 10353 24887 10387
rect 24687 10306 24887 10353
rect 25059 10387 25259 10403
rect 25059 10353 25075 10387
rect 25243 10353 25259 10387
rect 25059 10306 25259 10353
rect 25431 10387 25631 10403
rect 25431 10353 25447 10387
rect 25615 10353 25631 10387
rect 25431 10306 25631 10353
rect 25803 10387 26003 10403
rect 25803 10353 25819 10387
rect 25987 10353 26003 10387
rect 25803 10306 26003 10353
rect 26175 10387 26375 10403
rect 26175 10353 26191 10387
rect 26359 10353 26375 10387
rect 26175 10306 26375 10353
rect 26547 10387 26747 10403
rect 26547 10353 26563 10387
rect 26731 10353 26747 10387
rect 26547 10306 26747 10353
rect 26919 10387 27119 10403
rect 26919 10353 26935 10387
rect 27103 10353 27119 10387
rect 26919 10306 27119 10353
rect 27291 10387 27491 10403
rect 27291 10353 27307 10387
rect 27475 10353 27491 10387
rect 27291 10306 27491 10353
rect 27663 10387 27863 10403
rect 27663 10353 27679 10387
rect 27847 10353 27863 10387
rect 27663 10306 27863 10353
rect 28035 10387 28235 10403
rect 28035 10353 28051 10387
rect 28219 10353 28235 10387
rect 28035 10306 28235 10353
rect 28407 10387 28607 10403
rect 28407 10353 28423 10387
rect 28591 10353 28607 10387
rect 28407 10306 28607 10353
rect 28779 10387 28979 10403
rect 28779 10353 28795 10387
rect 28963 10353 28979 10387
rect 28779 10306 28979 10353
rect 29151 10387 29351 10403
rect 29151 10353 29167 10387
rect 29335 10353 29351 10387
rect 29151 10306 29351 10353
rect 29523 10387 29723 10403
rect 29523 10353 29539 10387
rect 29707 10353 29723 10387
rect 29523 10306 29723 10353
rect 29895 10387 30095 10403
rect 29895 10353 29911 10387
rect 30079 10353 30095 10387
rect 29895 10306 30095 10353
rect 30267 10387 30467 10403
rect 30267 10353 30283 10387
rect 30451 10353 30467 10387
rect 30267 10306 30467 10353
rect 18735 9859 18935 9906
rect 18735 9825 18751 9859
rect 18919 9825 18935 9859
rect 18735 9809 18935 9825
rect 19107 9859 19307 9906
rect 19107 9825 19123 9859
rect 19291 9825 19307 9859
rect 19107 9809 19307 9825
rect 19479 9859 19679 9906
rect 19479 9825 19495 9859
rect 19663 9825 19679 9859
rect 19479 9809 19679 9825
rect 19851 9859 20051 9906
rect 19851 9825 19867 9859
rect 20035 9825 20051 9859
rect 19851 9809 20051 9825
rect 20223 9859 20423 9906
rect 20223 9825 20239 9859
rect 20407 9825 20423 9859
rect 20223 9809 20423 9825
rect 20595 9859 20795 9906
rect 20595 9825 20611 9859
rect 20779 9825 20795 9859
rect 20595 9809 20795 9825
rect 20967 9859 21167 9906
rect 20967 9825 20983 9859
rect 21151 9825 21167 9859
rect 20967 9809 21167 9825
rect 21339 9859 21539 9906
rect 21339 9825 21355 9859
rect 21523 9825 21539 9859
rect 21339 9809 21539 9825
rect 21711 9859 21911 9906
rect 21711 9825 21727 9859
rect 21895 9825 21911 9859
rect 21711 9809 21911 9825
rect 22083 9859 22283 9906
rect 22083 9825 22099 9859
rect 22267 9825 22283 9859
rect 22083 9809 22283 9825
rect 22455 9859 22655 9906
rect 22455 9825 22471 9859
rect 22639 9825 22655 9859
rect 22455 9809 22655 9825
rect 22827 9859 23027 9906
rect 22827 9825 22843 9859
rect 23011 9825 23027 9859
rect 22827 9809 23027 9825
rect 23199 9859 23399 9906
rect 23199 9825 23215 9859
rect 23383 9825 23399 9859
rect 23199 9809 23399 9825
rect 23571 9859 23771 9906
rect 23571 9825 23587 9859
rect 23755 9825 23771 9859
rect 23571 9809 23771 9825
rect 23943 9859 24143 9906
rect 23943 9825 23959 9859
rect 24127 9825 24143 9859
rect 23943 9809 24143 9825
rect 24315 9859 24515 9906
rect 24315 9825 24331 9859
rect 24499 9825 24515 9859
rect 24315 9809 24515 9825
rect 24687 9859 24887 9906
rect 24687 9825 24703 9859
rect 24871 9825 24887 9859
rect 24687 9809 24887 9825
rect 25059 9859 25259 9906
rect 25059 9825 25075 9859
rect 25243 9825 25259 9859
rect 25059 9809 25259 9825
rect 25431 9859 25631 9906
rect 25431 9825 25447 9859
rect 25615 9825 25631 9859
rect 25431 9809 25631 9825
rect 25803 9859 26003 9906
rect 25803 9825 25819 9859
rect 25987 9825 26003 9859
rect 25803 9809 26003 9825
rect 26175 9859 26375 9906
rect 26175 9825 26191 9859
rect 26359 9825 26375 9859
rect 26175 9809 26375 9825
rect 26547 9859 26747 9906
rect 26547 9825 26563 9859
rect 26731 9825 26747 9859
rect 26547 9809 26747 9825
rect 26919 9859 27119 9906
rect 26919 9825 26935 9859
rect 27103 9825 27119 9859
rect 26919 9809 27119 9825
rect 27291 9859 27491 9906
rect 27291 9825 27307 9859
rect 27475 9825 27491 9859
rect 27291 9809 27491 9825
rect 27663 9859 27863 9906
rect 27663 9825 27679 9859
rect 27847 9825 27863 9859
rect 27663 9809 27863 9825
rect 28035 9859 28235 9906
rect 28035 9825 28051 9859
rect 28219 9825 28235 9859
rect 28035 9809 28235 9825
rect 28407 9859 28607 9906
rect 28407 9825 28423 9859
rect 28591 9825 28607 9859
rect 28407 9809 28607 9825
rect 28779 9859 28979 9906
rect 28779 9825 28795 9859
rect 28963 9825 28979 9859
rect 28779 9809 28979 9825
rect 29151 9859 29351 9906
rect 29151 9825 29167 9859
rect 29335 9825 29351 9859
rect 29151 9809 29351 9825
rect 29523 9859 29723 9906
rect 29523 9825 29539 9859
rect 29707 9825 29723 9859
rect 29523 9809 29723 9825
rect 29895 9859 30095 9906
rect 29895 9825 29911 9859
rect 30079 9825 30095 9859
rect 29895 9809 30095 9825
rect 30267 9859 30467 9906
rect 30267 9825 30283 9859
rect 30451 9825 30467 9859
rect 30267 9809 30467 9825
rect 20223 9271 20423 9287
rect 20223 9237 20239 9271
rect 20407 9237 20423 9271
rect 20223 9190 20423 9237
rect 20595 9271 20795 9287
rect 20595 9237 20611 9271
rect 20779 9237 20795 9271
rect 20595 9190 20795 9237
rect 20967 9271 21167 9287
rect 20967 9237 20983 9271
rect 21151 9237 21167 9271
rect 20967 9190 21167 9237
rect 21339 9271 21539 9287
rect 21339 9237 21355 9271
rect 21523 9237 21539 9271
rect 21339 9190 21539 9237
rect 21711 9271 21911 9287
rect 21711 9237 21727 9271
rect 21895 9237 21911 9271
rect 21711 9190 21911 9237
rect 22083 9271 22283 9287
rect 22083 9237 22099 9271
rect 22267 9237 22283 9271
rect 22083 9190 22283 9237
rect 22455 9271 22655 9287
rect 22455 9237 22471 9271
rect 22639 9237 22655 9271
rect 22455 9190 22655 9237
rect 22827 9271 23027 9287
rect 22827 9237 22843 9271
rect 23011 9237 23027 9271
rect 22827 9190 23027 9237
rect 20223 8343 20423 8390
rect 20223 8309 20239 8343
rect 20407 8309 20423 8343
rect 20223 8293 20423 8309
rect 20595 8343 20795 8390
rect 20595 8309 20611 8343
rect 20779 8309 20795 8343
rect 20595 8293 20795 8309
rect 20967 8343 21167 8390
rect 20967 8309 20983 8343
rect 21151 8309 21167 8343
rect 20967 8293 21167 8309
rect 21339 8343 21539 8390
rect 21339 8309 21355 8343
rect 21523 8309 21539 8343
rect 21339 8293 21539 8309
rect 21711 8343 21911 8390
rect 21711 8309 21727 8343
rect 21895 8309 21911 8343
rect 21711 8293 21911 8309
rect 22083 8343 22283 8390
rect 22083 8309 22099 8343
rect 22267 8309 22283 8343
rect 22083 8293 22283 8309
rect 22455 8343 22655 8390
rect 22455 8309 22471 8343
rect 22639 8309 22655 8343
rect 22455 8293 22655 8309
rect 22827 8343 23027 8390
rect 22827 8309 22843 8343
rect 23011 8309 23027 8343
rect 22827 8293 23027 8309
rect 20223 8235 20423 8251
rect 20223 8201 20239 8235
rect 20407 8201 20423 8235
rect 20223 8154 20423 8201
rect 20595 8235 20795 8251
rect 20595 8201 20611 8235
rect 20779 8201 20795 8235
rect 20595 8154 20795 8201
rect 20967 8235 21167 8251
rect 20967 8201 20983 8235
rect 21151 8201 21167 8235
rect 20967 8154 21167 8201
rect 21339 8235 21539 8251
rect 21339 8201 21355 8235
rect 21523 8201 21539 8235
rect 21339 8154 21539 8201
rect 21711 8235 21911 8251
rect 21711 8201 21727 8235
rect 21895 8201 21911 8235
rect 21711 8154 21911 8201
rect 22083 8235 22283 8251
rect 22083 8201 22099 8235
rect 22267 8201 22283 8235
rect 22083 8154 22283 8201
rect 22455 8235 22655 8251
rect 22455 8201 22471 8235
rect 22639 8201 22655 8235
rect 22455 8154 22655 8201
rect 22827 8235 23027 8251
rect 22827 8201 22843 8235
rect 23011 8201 23027 8235
rect 22827 8154 23027 8201
rect 20223 7307 20423 7354
rect 20223 7273 20239 7307
rect 20407 7273 20423 7307
rect 20223 7257 20423 7273
rect 20595 7307 20795 7354
rect 20595 7273 20611 7307
rect 20779 7273 20795 7307
rect 20595 7257 20795 7273
rect 20967 7307 21167 7354
rect 20967 7273 20983 7307
rect 21151 7273 21167 7307
rect 20967 7257 21167 7273
rect 21339 7307 21539 7354
rect 21339 7273 21355 7307
rect 21523 7273 21539 7307
rect 21339 7257 21539 7273
rect 21711 7307 21911 7354
rect 21711 7273 21727 7307
rect 21895 7273 21911 7307
rect 21711 7257 21911 7273
rect 22083 7307 22283 7354
rect 22083 7273 22099 7307
rect 22267 7273 22283 7307
rect 22083 7257 22283 7273
rect 22455 7307 22655 7354
rect 22455 7273 22471 7307
rect 22639 7273 22655 7307
rect 22455 7257 22655 7273
rect 22827 7307 23027 7354
rect 22827 7273 22843 7307
rect 23011 7273 23027 7307
rect 22827 7257 23027 7273
rect 20223 7199 20423 7215
rect 20223 7165 20239 7199
rect 20407 7165 20423 7199
rect 20223 7118 20423 7165
rect 20595 7199 20795 7215
rect 20595 7165 20611 7199
rect 20779 7165 20795 7199
rect 20595 7118 20795 7165
rect 20967 7199 21167 7215
rect 20967 7165 20983 7199
rect 21151 7165 21167 7199
rect 20967 7118 21167 7165
rect 21339 7199 21539 7215
rect 21339 7165 21355 7199
rect 21523 7165 21539 7199
rect 21339 7118 21539 7165
rect 21711 7199 21911 7215
rect 21711 7165 21727 7199
rect 21895 7165 21911 7199
rect 21711 7118 21911 7165
rect 22083 7199 22283 7215
rect 22083 7165 22099 7199
rect 22267 7165 22283 7199
rect 22083 7118 22283 7165
rect 22455 7199 22655 7215
rect 22455 7165 22471 7199
rect 22639 7165 22655 7199
rect 22455 7118 22655 7165
rect 22827 7199 23027 7215
rect 22827 7165 22843 7199
rect 23011 7165 23027 7199
rect 22827 7118 23027 7165
rect 20223 6271 20423 6318
rect 20223 6237 20239 6271
rect 20407 6237 20423 6271
rect 20223 6221 20423 6237
rect 20595 6271 20795 6318
rect 20595 6237 20611 6271
rect 20779 6237 20795 6271
rect 20595 6221 20795 6237
rect 20967 6271 21167 6318
rect 20967 6237 20983 6271
rect 21151 6237 21167 6271
rect 20967 6221 21167 6237
rect 21339 6271 21539 6318
rect 21339 6237 21355 6271
rect 21523 6237 21539 6271
rect 21339 6221 21539 6237
rect 21711 6271 21911 6318
rect 21711 6237 21727 6271
rect 21895 6237 21911 6271
rect 21711 6221 21911 6237
rect 22083 6271 22283 6318
rect 22083 6237 22099 6271
rect 22267 6237 22283 6271
rect 22083 6221 22283 6237
rect 22455 6271 22655 6318
rect 22455 6237 22471 6271
rect 22639 6237 22655 6271
rect 22455 6221 22655 6237
rect 22827 6271 23027 6318
rect 22827 6237 22843 6271
rect 23011 6237 23027 6271
rect 22827 6221 23027 6237
rect 20223 6163 20423 6179
rect 20223 6129 20239 6163
rect 20407 6129 20423 6163
rect 20223 6082 20423 6129
rect 20595 6163 20795 6179
rect 20595 6129 20611 6163
rect 20779 6129 20795 6163
rect 20595 6082 20795 6129
rect 20967 6163 21167 6179
rect 20967 6129 20983 6163
rect 21151 6129 21167 6163
rect 20967 6082 21167 6129
rect 21339 6163 21539 6179
rect 21339 6129 21355 6163
rect 21523 6129 21539 6163
rect 21339 6082 21539 6129
rect 21711 6163 21911 6179
rect 21711 6129 21727 6163
rect 21895 6129 21911 6163
rect 21711 6082 21911 6129
rect 22083 6163 22283 6179
rect 22083 6129 22099 6163
rect 22267 6129 22283 6163
rect 22083 6082 22283 6129
rect 22455 6163 22655 6179
rect 22455 6129 22471 6163
rect 22639 6129 22655 6163
rect 22455 6082 22655 6129
rect 22827 6163 23027 6179
rect 22827 6129 22843 6163
rect 23011 6129 23027 6163
rect 22827 6082 23027 6129
rect 20223 5235 20423 5282
rect 20223 5201 20239 5235
rect 20407 5201 20423 5235
rect 20223 5185 20423 5201
rect 20595 5235 20795 5282
rect 20595 5201 20611 5235
rect 20779 5201 20795 5235
rect 20595 5185 20795 5201
rect 20967 5235 21167 5282
rect 20967 5201 20983 5235
rect 21151 5201 21167 5235
rect 20967 5185 21167 5201
rect 21339 5235 21539 5282
rect 21339 5201 21355 5235
rect 21523 5201 21539 5235
rect 21339 5185 21539 5201
rect 21711 5235 21911 5282
rect 21711 5201 21727 5235
rect 21895 5201 21911 5235
rect 21711 5185 21911 5201
rect 22083 5235 22283 5282
rect 22083 5201 22099 5235
rect 22267 5201 22283 5235
rect 22083 5185 22283 5201
rect 22455 5235 22655 5282
rect 22455 5201 22471 5235
rect 22639 5201 22655 5235
rect 22455 5185 22655 5201
rect 22827 5235 23027 5282
rect 22827 5201 22843 5235
rect 23011 5201 23027 5235
rect 22827 5185 23027 5201
rect 20223 4577 20423 4593
rect 20223 4543 20239 4577
rect 20407 4543 20423 4577
rect 20223 4505 20423 4543
rect 20595 4577 20795 4593
rect 20595 4543 20611 4577
rect 20779 4543 20795 4577
rect 20595 4505 20795 4543
rect 20967 4577 21167 4593
rect 20967 4543 20983 4577
rect 21151 4543 21167 4577
rect 20967 4505 21167 4543
rect 21339 4577 21539 4593
rect 21339 4543 21355 4577
rect 21523 4543 21539 4577
rect 21339 4505 21539 4543
rect 21711 4577 21911 4593
rect 21711 4543 21727 4577
rect 21895 4543 21911 4577
rect 21711 4505 21911 4543
rect 22083 4577 22283 4593
rect 22083 4543 22099 4577
rect 22267 4543 22283 4577
rect 22083 4505 22283 4543
rect 22455 4577 22655 4593
rect 22455 4543 22471 4577
rect 22639 4543 22655 4577
rect 22455 4505 22655 4543
rect 22827 4577 23027 4593
rect 22827 4543 22843 4577
rect 23011 4543 23027 4577
rect 22827 4505 23027 4543
rect 23199 4577 23399 4593
rect 23199 4543 23215 4577
rect 23383 4543 23399 4577
rect 23199 4505 23399 4543
rect 23571 4577 23771 4593
rect 23571 4543 23587 4577
rect 23755 4543 23771 4577
rect 23571 4505 23771 4543
rect 23943 4577 24143 4593
rect 23943 4543 23959 4577
rect 24127 4543 24143 4577
rect 23943 4505 24143 4543
rect 24315 4577 24515 4593
rect 24315 4543 24331 4577
rect 24499 4543 24515 4577
rect 24315 4505 24515 4543
rect 24687 4577 24887 4593
rect 24687 4543 24703 4577
rect 24871 4543 24887 4577
rect 24687 4505 24887 4543
rect 25059 4577 25259 4593
rect 25059 4543 25075 4577
rect 25243 4543 25259 4577
rect 25059 4505 25259 4543
rect 25431 4577 25631 4593
rect 25431 4543 25447 4577
rect 25615 4543 25631 4577
rect 25431 4505 25631 4543
rect 25803 4577 26003 4593
rect 25803 4543 25819 4577
rect 25987 4543 26003 4577
rect 25803 4505 26003 4543
rect 26175 4577 26375 4593
rect 26175 4543 26191 4577
rect 26359 4543 26375 4577
rect 26175 4505 26375 4543
rect 26547 4577 26747 4593
rect 26547 4543 26563 4577
rect 26731 4543 26747 4577
rect 26547 4505 26747 4543
rect 26919 4577 27119 4593
rect 26919 4543 26935 4577
rect 27103 4543 27119 4577
rect 26919 4505 27119 4543
rect 27291 4577 27491 4593
rect 27291 4543 27307 4577
rect 27475 4543 27491 4577
rect 27291 4505 27491 4543
rect 27663 4577 27863 4593
rect 27663 4543 27679 4577
rect 27847 4543 27863 4577
rect 27663 4505 27863 4543
rect 28035 4577 28235 4593
rect 28035 4543 28051 4577
rect 28219 4543 28235 4577
rect 28035 4505 28235 4543
rect 28407 4577 28607 4593
rect 28407 4543 28423 4577
rect 28591 4543 28607 4577
rect 28407 4505 28607 4543
rect 28779 4577 28979 4593
rect 28779 4543 28795 4577
rect 28963 4543 28979 4577
rect 28779 4505 28979 4543
rect 20223 4267 20423 4305
rect 20223 4233 20239 4267
rect 20407 4233 20423 4267
rect 20223 4217 20423 4233
rect 20595 4267 20795 4305
rect 20595 4233 20611 4267
rect 20779 4233 20795 4267
rect 20595 4217 20795 4233
rect 20967 4267 21167 4305
rect 20967 4233 20983 4267
rect 21151 4233 21167 4267
rect 20967 4217 21167 4233
rect 21339 4267 21539 4305
rect 21339 4233 21355 4267
rect 21523 4233 21539 4267
rect 21339 4217 21539 4233
rect 21711 4267 21911 4305
rect 21711 4233 21727 4267
rect 21895 4233 21911 4267
rect 21711 4217 21911 4233
rect 22083 4267 22283 4305
rect 22083 4233 22099 4267
rect 22267 4233 22283 4267
rect 22083 4217 22283 4233
rect 22455 4267 22655 4305
rect 22455 4233 22471 4267
rect 22639 4233 22655 4267
rect 22455 4217 22655 4233
rect 22827 4267 23027 4305
rect 22827 4233 22843 4267
rect 23011 4233 23027 4267
rect 22827 4217 23027 4233
rect 23199 4267 23399 4305
rect 23199 4233 23215 4267
rect 23383 4233 23399 4267
rect 23199 4217 23399 4233
rect 23571 4267 23771 4305
rect 23571 4233 23587 4267
rect 23755 4233 23771 4267
rect 23571 4217 23771 4233
rect 23943 4267 24143 4305
rect 23943 4233 23959 4267
rect 24127 4233 24143 4267
rect 23943 4217 24143 4233
rect 24315 4267 24515 4305
rect 24315 4233 24331 4267
rect 24499 4233 24515 4267
rect 24315 4217 24515 4233
rect 24687 4267 24887 4305
rect 24687 4233 24703 4267
rect 24871 4233 24887 4267
rect 24687 4217 24887 4233
rect 25059 4267 25259 4305
rect 25059 4233 25075 4267
rect 25243 4233 25259 4267
rect 25059 4217 25259 4233
rect 25431 4267 25631 4305
rect 25431 4233 25447 4267
rect 25615 4233 25631 4267
rect 25431 4217 25631 4233
rect 25803 4267 26003 4305
rect 25803 4233 25819 4267
rect 25987 4233 26003 4267
rect 25803 4217 26003 4233
rect 26175 4267 26375 4305
rect 26175 4233 26191 4267
rect 26359 4233 26375 4267
rect 26175 4217 26375 4233
rect 26547 4267 26747 4305
rect 26547 4233 26563 4267
rect 26731 4233 26747 4267
rect 26547 4217 26747 4233
rect 26919 4267 27119 4305
rect 26919 4233 26935 4267
rect 27103 4233 27119 4267
rect 26919 4217 27119 4233
rect 27291 4267 27491 4305
rect 27291 4233 27307 4267
rect 27475 4233 27491 4267
rect 27291 4217 27491 4233
rect 27663 4267 27863 4305
rect 27663 4233 27679 4267
rect 27847 4233 27863 4267
rect 27663 4217 27863 4233
rect 28035 4267 28235 4305
rect 28035 4233 28051 4267
rect 28219 4233 28235 4267
rect 28035 4217 28235 4233
rect 28407 4267 28607 4305
rect 28407 4233 28423 4267
rect 28591 4233 28607 4267
rect 28407 4217 28607 4233
rect 28779 4267 28979 4305
rect 28779 4233 28795 4267
rect 28963 4233 28979 4267
rect 28779 4217 28979 4233
rect 20223 4159 20423 4175
rect 20223 4125 20239 4159
rect 20407 4125 20423 4159
rect 20223 4087 20423 4125
rect 20595 4159 20795 4175
rect 20595 4125 20611 4159
rect 20779 4125 20795 4159
rect 20595 4087 20795 4125
rect 20967 4159 21167 4175
rect 20967 4125 20983 4159
rect 21151 4125 21167 4159
rect 20967 4087 21167 4125
rect 21339 4159 21539 4175
rect 21339 4125 21355 4159
rect 21523 4125 21539 4159
rect 21339 4087 21539 4125
rect 21711 4159 21911 4175
rect 21711 4125 21727 4159
rect 21895 4125 21911 4159
rect 21711 4087 21911 4125
rect 22083 4159 22283 4175
rect 22083 4125 22099 4159
rect 22267 4125 22283 4159
rect 22083 4087 22283 4125
rect 22455 4159 22655 4175
rect 22455 4125 22471 4159
rect 22639 4125 22655 4159
rect 22455 4087 22655 4125
rect 22827 4159 23027 4175
rect 22827 4125 22843 4159
rect 23011 4125 23027 4159
rect 22827 4087 23027 4125
rect 23199 4159 23399 4175
rect 23199 4125 23215 4159
rect 23383 4125 23399 4159
rect 23199 4087 23399 4125
rect 23571 4159 23771 4175
rect 23571 4125 23587 4159
rect 23755 4125 23771 4159
rect 23571 4087 23771 4125
rect 23943 4159 24143 4175
rect 23943 4125 23959 4159
rect 24127 4125 24143 4159
rect 23943 4087 24143 4125
rect 24315 4159 24515 4175
rect 24315 4125 24331 4159
rect 24499 4125 24515 4159
rect 24315 4087 24515 4125
rect 24687 4159 24887 4175
rect 24687 4125 24703 4159
rect 24871 4125 24887 4159
rect 24687 4087 24887 4125
rect 25059 4159 25259 4175
rect 25059 4125 25075 4159
rect 25243 4125 25259 4159
rect 25059 4087 25259 4125
rect 25431 4159 25631 4175
rect 25431 4125 25447 4159
rect 25615 4125 25631 4159
rect 25431 4087 25631 4125
rect 25803 4159 26003 4175
rect 25803 4125 25819 4159
rect 25987 4125 26003 4159
rect 25803 4087 26003 4125
rect 26175 4159 26375 4175
rect 26175 4125 26191 4159
rect 26359 4125 26375 4159
rect 26175 4087 26375 4125
rect 26547 4159 26747 4175
rect 26547 4125 26563 4159
rect 26731 4125 26747 4159
rect 26547 4087 26747 4125
rect 26919 4159 27119 4175
rect 26919 4125 26935 4159
rect 27103 4125 27119 4159
rect 26919 4087 27119 4125
rect 27291 4159 27491 4175
rect 27291 4125 27307 4159
rect 27475 4125 27491 4159
rect 27291 4087 27491 4125
rect 27663 4159 27863 4175
rect 27663 4125 27679 4159
rect 27847 4125 27863 4159
rect 27663 4087 27863 4125
rect 28035 4159 28235 4175
rect 28035 4125 28051 4159
rect 28219 4125 28235 4159
rect 28035 4087 28235 4125
rect 28407 4159 28607 4175
rect 28407 4125 28423 4159
rect 28591 4125 28607 4159
rect 28407 4087 28607 4125
rect 28779 4159 28979 4175
rect 28779 4125 28795 4159
rect 28963 4125 28979 4159
rect 28779 4087 28979 4125
rect 20223 3849 20423 3887
rect 20223 3815 20239 3849
rect 20407 3815 20423 3849
rect 20223 3799 20423 3815
rect 20595 3849 20795 3887
rect 20595 3815 20611 3849
rect 20779 3815 20795 3849
rect 20595 3799 20795 3815
rect 20967 3849 21167 3887
rect 20967 3815 20983 3849
rect 21151 3815 21167 3849
rect 20967 3799 21167 3815
rect 21339 3849 21539 3887
rect 21339 3815 21355 3849
rect 21523 3815 21539 3849
rect 21339 3799 21539 3815
rect 21711 3849 21911 3887
rect 21711 3815 21727 3849
rect 21895 3815 21911 3849
rect 21711 3799 21911 3815
rect 22083 3849 22283 3887
rect 22083 3815 22099 3849
rect 22267 3815 22283 3849
rect 22083 3799 22283 3815
rect 22455 3849 22655 3887
rect 22455 3815 22471 3849
rect 22639 3815 22655 3849
rect 22455 3799 22655 3815
rect 22827 3849 23027 3887
rect 22827 3815 22843 3849
rect 23011 3815 23027 3849
rect 22827 3799 23027 3815
rect 23199 3849 23399 3887
rect 23199 3815 23215 3849
rect 23383 3815 23399 3849
rect 23199 3799 23399 3815
rect 23571 3849 23771 3887
rect 23571 3815 23587 3849
rect 23755 3815 23771 3849
rect 23571 3799 23771 3815
rect 23943 3849 24143 3887
rect 23943 3815 23959 3849
rect 24127 3815 24143 3849
rect 23943 3799 24143 3815
rect 24315 3849 24515 3887
rect 24315 3815 24331 3849
rect 24499 3815 24515 3849
rect 24315 3799 24515 3815
rect 24687 3849 24887 3887
rect 24687 3815 24703 3849
rect 24871 3815 24887 3849
rect 24687 3799 24887 3815
rect 25059 3849 25259 3887
rect 25059 3815 25075 3849
rect 25243 3815 25259 3849
rect 25059 3799 25259 3815
rect 25431 3849 25631 3887
rect 25431 3815 25447 3849
rect 25615 3815 25631 3849
rect 25431 3799 25631 3815
rect 25803 3849 26003 3887
rect 25803 3815 25819 3849
rect 25987 3815 26003 3849
rect 25803 3799 26003 3815
rect 26175 3849 26375 3887
rect 26175 3815 26191 3849
rect 26359 3815 26375 3849
rect 26175 3799 26375 3815
rect 26547 3849 26747 3887
rect 26547 3815 26563 3849
rect 26731 3815 26747 3849
rect 26547 3799 26747 3815
rect 26919 3849 27119 3887
rect 26919 3815 26935 3849
rect 27103 3815 27119 3849
rect 26919 3799 27119 3815
rect 27291 3849 27491 3887
rect 27291 3815 27307 3849
rect 27475 3815 27491 3849
rect 27291 3799 27491 3815
rect 27663 3849 27863 3887
rect 27663 3815 27679 3849
rect 27847 3815 27863 3849
rect 27663 3799 27863 3815
rect 28035 3849 28235 3887
rect 28035 3815 28051 3849
rect 28219 3815 28235 3849
rect 28035 3799 28235 3815
rect 28407 3849 28607 3887
rect 28407 3815 28423 3849
rect 28591 3815 28607 3849
rect 28407 3799 28607 3815
rect 28779 3849 28979 3887
rect 28779 3815 28795 3849
rect 28963 3815 28979 3849
rect 28779 3799 28979 3815
rect 20223 3741 20423 3757
rect 20223 3707 20239 3741
rect 20407 3707 20423 3741
rect 20223 3669 20423 3707
rect 20595 3741 20795 3757
rect 20595 3707 20611 3741
rect 20779 3707 20795 3741
rect 20595 3669 20795 3707
rect 20967 3741 21167 3757
rect 20967 3707 20983 3741
rect 21151 3707 21167 3741
rect 20967 3669 21167 3707
rect 21339 3741 21539 3757
rect 21339 3707 21355 3741
rect 21523 3707 21539 3741
rect 21339 3669 21539 3707
rect 21711 3741 21911 3757
rect 21711 3707 21727 3741
rect 21895 3707 21911 3741
rect 21711 3669 21911 3707
rect 22083 3741 22283 3757
rect 22083 3707 22099 3741
rect 22267 3707 22283 3741
rect 22083 3669 22283 3707
rect 22455 3741 22655 3757
rect 22455 3707 22471 3741
rect 22639 3707 22655 3741
rect 22455 3669 22655 3707
rect 22827 3741 23027 3757
rect 22827 3707 22843 3741
rect 23011 3707 23027 3741
rect 22827 3669 23027 3707
rect 23199 3741 23399 3757
rect 23199 3707 23215 3741
rect 23383 3707 23399 3741
rect 23199 3669 23399 3707
rect 23571 3741 23771 3757
rect 23571 3707 23587 3741
rect 23755 3707 23771 3741
rect 23571 3669 23771 3707
rect 23943 3741 24143 3757
rect 23943 3707 23959 3741
rect 24127 3707 24143 3741
rect 23943 3669 24143 3707
rect 24315 3741 24515 3757
rect 24315 3707 24331 3741
rect 24499 3707 24515 3741
rect 24315 3669 24515 3707
rect 24687 3741 24887 3757
rect 24687 3707 24703 3741
rect 24871 3707 24887 3741
rect 24687 3669 24887 3707
rect 25059 3741 25259 3757
rect 25059 3707 25075 3741
rect 25243 3707 25259 3741
rect 25059 3669 25259 3707
rect 25431 3741 25631 3757
rect 25431 3707 25447 3741
rect 25615 3707 25631 3741
rect 25431 3669 25631 3707
rect 25803 3741 26003 3757
rect 25803 3707 25819 3741
rect 25987 3707 26003 3741
rect 25803 3669 26003 3707
rect 26175 3741 26375 3757
rect 26175 3707 26191 3741
rect 26359 3707 26375 3741
rect 26175 3669 26375 3707
rect 26547 3741 26747 3757
rect 26547 3707 26563 3741
rect 26731 3707 26747 3741
rect 26547 3669 26747 3707
rect 26919 3741 27119 3757
rect 26919 3707 26935 3741
rect 27103 3707 27119 3741
rect 26919 3669 27119 3707
rect 27291 3741 27491 3757
rect 27291 3707 27307 3741
rect 27475 3707 27491 3741
rect 27291 3669 27491 3707
rect 27663 3741 27863 3757
rect 27663 3707 27679 3741
rect 27847 3707 27863 3741
rect 27663 3669 27863 3707
rect 28035 3741 28235 3757
rect 28035 3707 28051 3741
rect 28219 3707 28235 3741
rect 28035 3669 28235 3707
rect 28407 3741 28607 3757
rect 28407 3707 28423 3741
rect 28591 3707 28607 3741
rect 28407 3669 28607 3707
rect 28779 3741 28979 3757
rect 28779 3707 28795 3741
rect 28963 3707 28979 3741
rect 28779 3669 28979 3707
rect 20223 3431 20423 3469
rect 20223 3397 20239 3431
rect 20407 3397 20423 3431
rect 20223 3381 20423 3397
rect 20595 3431 20795 3469
rect 20595 3397 20611 3431
rect 20779 3397 20795 3431
rect 20595 3381 20795 3397
rect 20967 3431 21167 3469
rect 20967 3397 20983 3431
rect 21151 3397 21167 3431
rect 20967 3381 21167 3397
rect 21339 3431 21539 3469
rect 21339 3397 21355 3431
rect 21523 3397 21539 3431
rect 21339 3381 21539 3397
rect 21711 3431 21911 3469
rect 21711 3397 21727 3431
rect 21895 3397 21911 3431
rect 21711 3381 21911 3397
rect 22083 3431 22283 3469
rect 22083 3397 22099 3431
rect 22267 3397 22283 3431
rect 22083 3381 22283 3397
rect 22455 3431 22655 3469
rect 22455 3397 22471 3431
rect 22639 3397 22655 3431
rect 22455 3381 22655 3397
rect 22827 3431 23027 3469
rect 22827 3397 22843 3431
rect 23011 3397 23027 3431
rect 22827 3381 23027 3397
rect 23199 3431 23399 3469
rect 23199 3397 23215 3431
rect 23383 3397 23399 3431
rect 23199 3381 23399 3397
rect 23571 3431 23771 3469
rect 23571 3397 23587 3431
rect 23755 3397 23771 3431
rect 23571 3381 23771 3397
rect 23943 3431 24143 3469
rect 23943 3397 23959 3431
rect 24127 3397 24143 3431
rect 23943 3381 24143 3397
rect 24315 3431 24515 3469
rect 24315 3397 24331 3431
rect 24499 3397 24515 3431
rect 24315 3381 24515 3397
rect 24687 3431 24887 3469
rect 24687 3397 24703 3431
rect 24871 3397 24887 3431
rect 24687 3381 24887 3397
rect 25059 3431 25259 3469
rect 25059 3397 25075 3431
rect 25243 3397 25259 3431
rect 25059 3381 25259 3397
rect 25431 3431 25631 3469
rect 25431 3397 25447 3431
rect 25615 3397 25631 3431
rect 25431 3381 25631 3397
rect 25803 3431 26003 3469
rect 25803 3397 25819 3431
rect 25987 3397 26003 3431
rect 25803 3381 26003 3397
rect 26175 3431 26375 3469
rect 26175 3397 26191 3431
rect 26359 3397 26375 3431
rect 26175 3381 26375 3397
rect 26547 3431 26747 3469
rect 26547 3397 26563 3431
rect 26731 3397 26747 3431
rect 26547 3381 26747 3397
rect 26919 3431 27119 3469
rect 26919 3397 26935 3431
rect 27103 3397 27119 3431
rect 26919 3381 27119 3397
rect 27291 3431 27491 3469
rect 27291 3397 27307 3431
rect 27475 3397 27491 3431
rect 27291 3381 27491 3397
rect 27663 3431 27863 3469
rect 27663 3397 27679 3431
rect 27847 3397 27863 3431
rect 27663 3381 27863 3397
rect 28035 3431 28235 3469
rect 28035 3397 28051 3431
rect 28219 3397 28235 3431
rect 28035 3381 28235 3397
rect 28407 3431 28607 3469
rect 28407 3397 28423 3431
rect 28591 3397 28607 3431
rect 28407 3381 28607 3397
rect 28779 3431 28979 3469
rect 28779 3397 28795 3431
rect 28963 3397 28979 3431
rect 28779 3381 28979 3397
rect 20223 3323 20423 3339
rect 20223 3289 20239 3323
rect 20407 3289 20423 3323
rect 20223 3251 20423 3289
rect 20595 3323 20795 3339
rect 20595 3289 20611 3323
rect 20779 3289 20795 3323
rect 20595 3251 20795 3289
rect 20967 3323 21167 3339
rect 20967 3289 20983 3323
rect 21151 3289 21167 3323
rect 20967 3251 21167 3289
rect 21339 3323 21539 3339
rect 21339 3289 21355 3323
rect 21523 3289 21539 3323
rect 21339 3251 21539 3289
rect 21711 3323 21911 3339
rect 21711 3289 21727 3323
rect 21895 3289 21911 3323
rect 21711 3251 21911 3289
rect 22083 3323 22283 3339
rect 22083 3289 22099 3323
rect 22267 3289 22283 3323
rect 22083 3251 22283 3289
rect 22455 3323 22655 3339
rect 22455 3289 22471 3323
rect 22639 3289 22655 3323
rect 22455 3251 22655 3289
rect 22827 3323 23027 3339
rect 22827 3289 22843 3323
rect 23011 3289 23027 3323
rect 22827 3251 23027 3289
rect 23199 3323 23399 3339
rect 23199 3289 23215 3323
rect 23383 3289 23399 3323
rect 23199 3251 23399 3289
rect 23571 3323 23771 3339
rect 23571 3289 23587 3323
rect 23755 3289 23771 3323
rect 23571 3251 23771 3289
rect 23943 3323 24143 3339
rect 23943 3289 23959 3323
rect 24127 3289 24143 3323
rect 23943 3251 24143 3289
rect 24315 3323 24515 3339
rect 24315 3289 24331 3323
rect 24499 3289 24515 3323
rect 24315 3251 24515 3289
rect 24687 3323 24887 3339
rect 24687 3289 24703 3323
rect 24871 3289 24887 3323
rect 24687 3251 24887 3289
rect 25059 3323 25259 3339
rect 25059 3289 25075 3323
rect 25243 3289 25259 3323
rect 25059 3251 25259 3289
rect 25431 3323 25631 3339
rect 25431 3289 25447 3323
rect 25615 3289 25631 3323
rect 25431 3251 25631 3289
rect 25803 3323 26003 3339
rect 25803 3289 25819 3323
rect 25987 3289 26003 3323
rect 25803 3251 26003 3289
rect 26175 3323 26375 3339
rect 26175 3289 26191 3323
rect 26359 3289 26375 3323
rect 26175 3251 26375 3289
rect 26547 3323 26747 3339
rect 26547 3289 26563 3323
rect 26731 3289 26747 3323
rect 26547 3251 26747 3289
rect 26919 3323 27119 3339
rect 26919 3289 26935 3323
rect 27103 3289 27119 3323
rect 26919 3251 27119 3289
rect 27291 3323 27491 3339
rect 27291 3289 27307 3323
rect 27475 3289 27491 3323
rect 27291 3251 27491 3289
rect 27663 3323 27863 3339
rect 27663 3289 27679 3323
rect 27847 3289 27863 3323
rect 27663 3251 27863 3289
rect 28035 3323 28235 3339
rect 28035 3289 28051 3323
rect 28219 3289 28235 3323
rect 28035 3251 28235 3289
rect 28407 3323 28607 3339
rect 28407 3289 28423 3323
rect 28591 3289 28607 3323
rect 28407 3251 28607 3289
rect 28779 3323 28979 3339
rect 28779 3289 28795 3323
rect 28963 3289 28979 3323
rect 28779 3251 28979 3289
rect 20223 3013 20423 3051
rect 20223 2979 20239 3013
rect 20407 2979 20423 3013
rect 20223 2963 20423 2979
rect 20595 3013 20795 3051
rect 20595 2979 20611 3013
rect 20779 2979 20795 3013
rect 20595 2963 20795 2979
rect 20967 3013 21167 3051
rect 20967 2979 20983 3013
rect 21151 2979 21167 3013
rect 20967 2963 21167 2979
rect 21339 3013 21539 3051
rect 21339 2979 21355 3013
rect 21523 2979 21539 3013
rect 21339 2963 21539 2979
rect 21711 3013 21911 3051
rect 21711 2979 21727 3013
rect 21895 2979 21911 3013
rect 21711 2963 21911 2979
rect 22083 3013 22283 3051
rect 22083 2979 22099 3013
rect 22267 2979 22283 3013
rect 22083 2963 22283 2979
rect 22455 3013 22655 3051
rect 22455 2979 22471 3013
rect 22639 2979 22655 3013
rect 22455 2963 22655 2979
rect 22827 3013 23027 3051
rect 22827 2979 22843 3013
rect 23011 2979 23027 3013
rect 22827 2963 23027 2979
rect 23199 3013 23399 3051
rect 23199 2979 23215 3013
rect 23383 2979 23399 3013
rect 23199 2963 23399 2979
rect 23571 3013 23771 3051
rect 23571 2979 23587 3013
rect 23755 2979 23771 3013
rect 23571 2963 23771 2979
rect 23943 3013 24143 3051
rect 23943 2979 23959 3013
rect 24127 2979 24143 3013
rect 23943 2963 24143 2979
rect 24315 3013 24515 3051
rect 24315 2979 24331 3013
rect 24499 2979 24515 3013
rect 24315 2963 24515 2979
rect 24687 3013 24887 3051
rect 24687 2979 24703 3013
rect 24871 2979 24887 3013
rect 24687 2963 24887 2979
rect 25059 3013 25259 3051
rect 25059 2979 25075 3013
rect 25243 2979 25259 3013
rect 25059 2963 25259 2979
rect 25431 3013 25631 3051
rect 25431 2979 25447 3013
rect 25615 2979 25631 3013
rect 25431 2963 25631 2979
rect 25803 3013 26003 3051
rect 25803 2979 25819 3013
rect 25987 2979 26003 3013
rect 25803 2963 26003 2979
rect 26175 3013 26375 3051
rect 26175 2979 26191 3013
rect 26359 2979 26375 3013
rect 26175 2963 26375 2979
rect 26547 3013 26747 3051
rect 26547 2979 26563 3013
rect 26731 2979 26747 3013
rect 26547 2963 26747 2979
rect 26919 3013 27119 3051
rect 26919 2979 26935 3013
rect 27103 2979 27119 3013
rect 26919 2963 27119 2979
rect 27291 3013 27491 3051
rect 27291 2979 27307 3013
rect 27475 2979 27491 3013
rect 27291 2963 27491 2979
rect 27663 3013 27863 3051
rect 27663 2979 27679 3013
rect 27847 2979 27863 3013
rect 27663 2963 27863 2979
rect 28035 3013 28235 3051
rect 28035 2979 28051 3013
rect 28219 2979 28235 3013
rect 28035 2963 28235 2979
rect 28407 3013 28607 3051
rect 28407 2979 28423 3013
rect 28591 2979 28607 3013
rect 28407 2963 28607 2979
rect 28779 3013 28979 3051
rect 28779 2979 28795 3013
rect 28963 2979 28979 3013
rect 28779 2963 28979 2979
<< polycont >>
rect 18751 11625 18919 11659
rect 19123 11625 19291 11659
rect 19495 11625 19663 11659
rect 19867 11625 20035 11659
rect 20239 11625 20407 11659
rect 20611 11625 20779 11659
rect 20983 11625 21151 11659
rect 21355 11625 21523 11659
rect 21727 11625 21895 11659
rect 22099 11625 22267 11659
rect 22471 11625 22639 11659
rect 22843 11625 23011 11659
rect 23215 11625 23383 11659
rect 23587 11625 23755 11659
rect 23959 11625 24127 11659
rect 24331 11625 24499 11659
rect 24703 11625 24871 11659
rect 25075 11625 25243 11659
rect 25447 11625 25615 11659
rect 25819 11625 25987 11659
rect 26191 11625 26359 11659
rect 26563 11625 26731 11659
rect 26935 11625 27103 11659
rect 27307 11625 27475 11659
rect 27679 11625 27847 11659
rect 28051 11625 28219 11659
rect 28423 11625 28591 11659
rect 28795 11625 28963 11659
rect 29167 11625 29335 11659
rect 29539 11625 29707 11659
rect 29911 11625 30079 11659
rect 30283 11625 30451 11659
rect 18751 11097 18919 11131
rect 19123 11097 19291 11131
rect 19495 11097 19663 11131
rect 19867 11097 20035 11131
rect 20239 11097 20407 11131
rect 20611 11097 20779 11131
rect 20983 11097 21151 11131
rect 21355 11097 21523 11131
rect 21727 11097 21895 11131
rect 22099 11097 22267 11131
rect 22471 11097 22639 11131
rect 22843 11097 23011 11131
rect 23215 11097 23383 11131
rect 23587 11097 23755 11131
rect 23959 11097 24127 11131
rect 24331 11097 24499 11131
rect 24703 11097 24871 11131
rect 25075 11097 25243 11131
rect 25447 11097 25615 11131
rect 25819 11097 25987 11131
rect 26191 11097 26359 11131
rect 26563 11097 26731 11131
rect 26935 11097 27103 11131
rect 27307 11097 27475 11131
rect 27679 11097 27847 11131
rect 28051 11097 28219 11131
rect 28423 11097 28591 11131
rect 28795 11097 28963 11131
rect 29167 11097 29335 11131
rect 29539 11097 29707 11131
rect 29911 11097 30079 11131
rect 30283 11097 30451 11131
rect 18751 10989 18919 11023
rect 19123 10989 19291 11023
rect 19495 10989 19663 11023
rect 19867 10989 20035 11023
rect 20239 10989 20407 11023
rect 20611 10989 20779 11023
rect 20983 10989 21151 11023
rect 21355 10989 21523 11023
rect 21727 10989 21895 11023
rect 22099 10989 22267 11023
rect 22471 10989 22639 11023
rect 22843 10989 23011 11023
rect 23215 10989 23383 11023
rect 23587 10989 23755 11023
rect 23959 10989 24127 11023
rect 24331 10989 24499 11023
rect 24703 10989 24871 11023
rect 25075 10989 25243 11023
rect 25447 10989 25615 11023
rect 25819 10989 25987 11023
rect 26191 10989 26359 11023
rect 26563 10989 26731 11023
rect 26935 10989 27103 11023
rect 27307 10989 27475 11023
rect 27679 10989 27847 11023
rect 28051 10989 28219 11023
rect 28423 10989 28591 11023
rect 28795 10989 28963 11023
rect 29167 10989 29335 11023
rect 29539 10989 29707 11023
rect 29911 10989 30079 11023
rect 30283 10989 30451 11023
rect 18751 10461 18919 10495
rect 19123 10461 19291 10495
rect 19495 10461 19663 10495
rect 19867 10461 20035 10495
rect 20239 10461 20407 10495
rect 20611 10461 20779 10495
rect 20983 10461 21151 10495
rect 21355 10461 21523 10495
rect 21727 10461 21895 10495
rect 22099 10461 22267 10495
rect 22471 10461 22639 10495
rect 22843 10461 23011 10495
rect 23215 10461 23383 10495
rect 23587 10461 23755 10495
rect 23959 10461 24127 10495
rect 24331 10461 24499 10495
rect 24703 10461 24871 10495
rect 25075 10461 25243 10495
rect 25447 10461 25615 10495
rect 25819 10461 25987 10495
rect 26191 10461 26359 10495
rect 26563 10461 26731 10495
rect 26935 10461 27103 10495
rect 27307 10461 27475 10495
rect 27679 10461 27847 10495
rect 28051 10461 28219 10495
rect 28423 10461 28591 10495
rect 28795 10461 28963 10495
rect 29167 10461 29335 10495
rect 29539 10461 29707 10495
rect 29911 10461 30079 10495
rect 30283 10461 30451 10495
rect 18751 10353 18919 10387
rect 19123 10353 19291 10387
rect 19495 10353 19663 10387
rect 19867 10353 20035 10387
rect 20239 10353 20407 10387
rect 20611 10353 20779 10387
rect 20983 10353 21151 10387
rect 21355 10353 21523 10387
rect 21727 10353 21895 10387
rect 22099 10353 22267 10387
rect 22471 10353 22639 10387
rect 22843 10353 23011 10387
rect 23215 10353 23383 10387
rect 23587 10353 23755 10387
rect 23959 10353 24127 10387
rect 24331 10353 24499 10387
rect 24703 10353 24871 10387
rect 25075 10353 25243 10387
rect 25447 10353 25615 10387
rect 25819 10353 25987 10387
rect 26191 10353 26359 10387
rect 26563 10353 26731 10387
rect 26935 10353 27103 10387
rect 27307 10353 27475 10387
rect 27679 10353 27847 10387
rect 28051 10353 28219 10387
rect 28423 10353 28591 10387
rect 28795 10353 28963 10387
rect 29167 10353 29335 10387
rect 29539 10353 29707 10387
rect 29911 10353 30079 10387
rect 30283 10353 30451 10387
rect 18751 9825 18919 9859
rect 19123 9825 19291 9859
rect 19495 9825 19663 9859
rect 19867 9825 20035 9859
rect 20239 9825 20407 9859
rect 20611 9825 20779 9859
rect 20983 9825 21151 9859
rect 21355 9825 21523 9859
rect 21727 9825 21895 9859
rect 22099 9825 22267 9859
rect 22471 9825 22639 9859
rect 22843 9825 23011 9859
rect 23215 9825 23383 9859
rect 23587 9825 23755 9859
rect 23959 9825 24127 9859
rect 24331 9825 24499 9859
rect 24703 9825 24871 9859
rect 25075 9825 25243 9859
rect 25447 9825 25615 9859
rect 25819 9825 25987 9859
rect 26191 9825 26359 9859
rect 26563 9825 26731 9859
rect 26935 9825 27103 9859
rect 27307 9825 27475 9859
rect 27679 9825 27847 9859
rect 28051 9825 28219 9859
rect 28423 9825 28591 9859
rect 28795 9825 28963 9859
rect 29167 9825 29335 9859
rect 29539 9825 29707 9859
rect 29911 9825 30079 9859
rect 30283 9825 30451 9859
rect 20239 9237 20407 9271
rect 20611 9237 20779 9271
rect 20983 9237 21151 9271
rect 21355 9237 21523 9271
rect 21727 9237 21895 9271
rect 22099 9237 22267 9271
rect 22471 9237 22639 9271
rect 22843 9237 23011 9271
rect 20239 8309 20407 8343
rect 20611 8309 20779 8343
rect 20983 8309 21151 8343
rect 21355 8309 21523 8343
rect 21727 8309 21895 8343
rect 22099 8309 22267 8343
rect 22471 8309 22639 8343
rect 22843 8309 23011 8343
rect 20239 8201 20407 8235
rect 20611 8201 20779 8235
rect 20983 8201 21151 8235
rect 21355 8201 21523 8235
rect 21727 8201 21895 8235
rect 22099 8201 22267 8235
rect 22471 8201 22639 8235
rect 22843 8201 23011 8235
rect 20239 7273 20407 7307
rect 20611 7273 20779 7307
rect 20983 7273 21151 7307
rect 21355 7273 21523 7307
rect 21727 7273 21895 7307
rect 22099 7273 22267 7307
rect 22471 7273 22639 7307
rect 22843 7273 23011 7307
rect 20239 7165 20407 7199
rect 20611 7165 20779 7199
rect 20983 7165 21151 7199
rect 21355 7165 21523 7199
rect 21727 7165 21895 7199
rect 22099 7165 22267 7199
rect 22471 7165 22639 7199
rect 22843 7165 23011 7199
rect 20239 6237 20407 6271
rect 20611 6237 20779 6271
rect 20983 6237 21151 6271
rect 21355 6237 21523 6271
rect 21727 6237 21895 6271
rect 22099 6237 22267 6271
rect 22471 6237 22639 6271
rect 22843 6237 23011 6271
rect 20239 6129 20407 6163
rect 20611 6129 20779 6163
rect 20983 6129 21151 6163
rect 21355 6129 21523 6163
rect 21727 6129 21895 6163
rect 22099 6129 22267 6163
rect 22471 6129 22639 6163
rect 22843 6129 23011 6163
rect 20239 5201 20407 5235
rect 20611 5201 20779 5235
rect 20983 5201 21151 5235
rect 21355 5201 21523 5235
rect 21727 5201 21895 5235
rect 22099 5201 22267 5235
rect 22471 5201 22639 5235
rect 22843 5201 23011 5235
rect 20239 4543 20407 4577
rect 20611 4543 20779 4577
rect 20983 4543 21151 4577
rect 21355 4543 21523 4577
rect 21727 4543 21895 4577
rect 22099 4543 22267 4577
rect 22471 4543 22639 4577
rect 22843 4543 23011 4577
rect 23215 4543 23383 4577
rect 23587 4543 23755 4577
rect 23959 4543 24127 4577
rect 24331 4543 24499 4577
rect 24703 4543 24871 4577
rect 25075 4543 25243 4577
rect 25447 4543 25615 4577
rect 25819 4543 25987 4577
rect 26191 4543 26359 4577
rect 26563 4543 26731 4577
rect 26935 4543 27103 4577
rect 27307 4543 27475 4577
rect 27679 4543 27847 4577
rect 28051 4543 28219 4577
rect 28423 4543 28591 4577
rect 28795 4543 28963 4577
rect 20239 4233 20407 4267
rect 20611 4233 20779 4267
rect 20983 4233 21151 4267
rect 21355 4233 21523 4267
rect 21727 4233 21895 4267
rect 22099 4233 22267 4267
rect 22471 4233 22639 4267
rect 22843 4233 23011 4267
rect 23215 4233 23383 4267
rect 23587 4233 23755 4267
rect 23959 4233 24127 4267
rect 24331 4233 24499 4267
rect 24703 4233 24871 4267
rect 25075 4233 25243 4267
rect 25447 4233 25615 4267
rect 25819 4233 25987 4267
rect 26191 4233 26359 4267
rect 26563 4233 26731 4267
rect 26935 4233 27103 4267
rect 27307 4233 27475 4267
rect 27679 4233 27847 4267
rect 28051 4233 28219 4267
rect 28423 4233 28591 4267
rect 28795 4233 28963 4267
rect 20239 4125 20407 4159
rect 20611 4125 20779 4159
rect 20983 4125 21151 4159
rect 21355 4125 21523 4159
rect 21727 4125 21895 4159
rect 22099 4125 22267 4159
rect 22471 4125 22639 4159
rect 22843 4125 23011 4159
rect 23215 4125 23383 4159
rect 23587 4125 23755 4159
rect 23959 4125 24127 4159
rect 24331 4125 24499 4159
rect 24703 4125 24871 4159
rect 25075 4125 25243 4159
rect 25447 4125 25615 4159
rect 25819 4125 25987 4159
rect 26191 4125 26359 4159
rect 26563 4125 26731 4159
rect 26935 4125 27103 4159
rect 27307 4125 27475 4159
rect 27679 4125 27847 4159
rect 28051 4125 28219 4159
rect 28423 4125 28591 4159
rect 28795 4125 28963 4159
rect 20239 3815 20407 3849
rect 20611 3815 20779 3849
rect 20983 3815 21151 3849
rect 21355 3815 21523 3849
rect 21727 3815 21895 3849
rect 22099 3815 22267 3849
rect 22471 3815 22639 3849
rect 22843 3815 23011 3849
rect 23215 3815 23383 3849
rect 23587 3815 23755 3849
rect 23959 3815 24127 3849
rect 24331 3815 24499 3849
rect 24703 3815 24871 3849
rect 25075 3815 25243 3849
rect 25447 3815 25615 3849
rect 25819 3815 25987 3849
rect 26191 3815 26359 3849
rect 26563 3815 26731 3849
rect 26935 3815 27103 3849
rect 27307 3815 27475 3849
rect 27679 3815 27847 3849
rect 28051 3815 28219 3849
rect 28423 3815 28591 3849
rect 28795 3815 28963 3849
rect 20239 3707 20407 3741
rect 20611 3707 20779 3741
rect 20983 3707 21151 3741
rect 21355 3707 21523 3741
rect 21727 3707 21895 3741
rect 22099 3707 22267 3741
rect 22471 3707 22639 3741
rect 22843 3707 23011 3741
rect 23215 3707 23383 3741
rect 23587 3707 23755 3741
rect 23959 3707 24127 3741
rect 24331 3707 24499 3741
rect 24703 3707 24871 3741
rect 25075 3707 25243 3741
rect 25447 3707 25615 3741
rect 25819 3707 25987 3741
rect 26191 3707 26359 3741
rect 26563 3707 26731 3741
rect 26935 3707 27103 3741
rect 27307 3707 27475 3741
rect 27679 3707 27847 3741
rect 28051 3707 28219 3741
rect 28423 3707 28591 3741
rect 28795 3707 28963 3741
rect 20239 3397 20407 3431
rect 20611 3397 20779 3431
rect 20983 3397 21151 3431
rect 21355 3397 21523 3431
rect 21727 3397 21895 3431
rect 22099 3397 22267 3431
rect 22471 3397 22639 3431
rect 22843 3397 23011 3431
rect 23215 3397 23383 3431
rect 23587 3397 23755 3431
rect 23959 3397 24127 3431
rect 24331 3397 24499 3431
rect 24703 3397 24871 3431
rect 25075 3397 25243 3431
rect 25447 3397 25615 3431
rect 25819 3397 25987 3431
rect 26191 3397 26359 3431
rect 26563 3397 26731 3431
rect 26935 3397 27103 3431
rect 27307 3397 27475 3431
rect 27679 3397 27847 3431
rect 28051 3397 28219 3431
rect 28423 3397 28591 3431
rect 28795 3397 28963 3431
rect 20239 3289 20407 3323
rect 20611 3289 20779 3323
rect 20983 3289 21151 3323
rect 21355 3289 21523 3323
rect 21727 3289 21895 3323
rect 22099 3289 22267 3323
rect 22471 3289 22639 3323
rect 22843 3289 23011 3323
rect 23215 3289 23383 3323
rect 23587 3289 23755 3323
rect 23959 3289 24127 3323
rect 24331 3289 24499 3323
rect 24703 3289 24871 3323
rect 25075 3289 25243 3323
rect 25447 3289 25615 3323
rect 25819 3289 25987 3323
rect 26191 3289 26359 3323
rect 26563 3289 26731 3323
rect 26935 3289 27103 3323
rect 27307 3289 27475 3323
rect 27679 3289 27847 3323
rect 28051 3289 28219 3323
rect 28423 3289 28591 3323
rect 28795 3289 28963 3323
rect 20239 2979 20407 3013
rect 20611 2979 20779 3013
rect 20983 2979 21151 3013
rect 21355 2979 21523 3013
rect 21727 2979 21895 3013
rect 22099 2979 22267 3013
rect 22471 2979 22639 3013
rect 22843 2979 23011 3013
rect 23215 2979 23383 3013
rect 23587 2979 23755 3013
rect 23959 2979 24127 3013
rect 24331 2979 24499 3013
rect 24703 2979 24871 3013
rect 25075 2979 25243 3013
rect 25447 2979 25615 3013
rect 25819 2979 25987 3013
rect 26191 2979 26359 3013
rect 26563 2979 26731 3013
rect 26935 2979 27103 3013
rect 27307 2979 27475 3013
rect 27679 2979 27847 3013
rect 28051 2979 28219 3013
rect 28423 2979 28591 3013
rect 28795 2979 28963 3013
<< xpolycontact >>
rect 23819 6897 23889 7329
rect 23819 5905 23889 6337
<< xpolyres >>
rect 23819 6337 23889 6897
<< locali >>
rect 18575 11727 18671 11761
rect 30534 11727 30627 11761
rect 18575 11665 18609 11727
rect 30593 11665 30627 11727
rect 18735 11625 18751 11659
rect 18919 11625 18935 11659
rect 19107 11625 19123 11659
rect 19291 11625 19307 11659
rect 19479 11625 19495 11659
rect 19663 11625 19679 11659
rect 19851 11625 19867 11659
rect 20035 11625 20051 11659
rect 20223 11625 20239 11659
rect 20407 11625 20423 11659
rect 20595 11625 20611 11659
rect 20779 11625 20795 11659
rect 20967 11625 20983 11659
rect 21151 11625 21167 11659
rect 21339 11625 21355 11659
rect 21523 11625 21539 11659
rect 21711 11625 21727 11659
rect 21895 11625 21911 11659
rect 22083 11625 22099 11659
rect 22267 11625 22283 11659
rect 22455 11625 22471 11659
rect 22639 11625 22655 11659
rect 22827 11625 22843 11659
rect 23011 11625 23027 11659
rect 23199 11625 23215 11659
rect 23383 11625 23399 11659
rect 23571 11625 23587 11659
rect 23755 11625 23771 11659
rect 23943 11625 23959 11659
rect 24127 11625 24143 11659
rect 24315 11625 24331 11659
rect 24499 11625 24515 11659
rect 24687 11625 24703 11659
rect 24871 11625 24887 11659
rect 25059 11625 25075 11659
rect 25243 11625 25259 11659
rect 25431 11625 25447 11659
rect 25615 11625 25631 11659
rect 25803 11625 25819 11659
rect 25987 11625 26003 11659
rect 26175 11625 26191 11659
rect 26359 11625 26375 11659
rect 26547 11625 26563 11659
rect 26731 11625 26747 11659
rect 26919 11625 26935 11659
rect 27103 11625 27119 11659
rect 27291 11625 27307 11659
rect 27475 11625 27491 11659
rect 27663 11625 27679 11659
rect 27847 11625 27863 11659
rect 28035 11625 28051 11659
rect 28219 11625 28235 11659
rect 28407 11625 28423 11659
rect 28591 11625 28607 11659
rect 28779 11625 28795 11659
rect 28963 11625 28979 11659
rect 29151 11625 29167 11659
rect 29335 11625 29351 11659
rect 29523 11625 29539 11659
rect 29707 11625 29723 11659
rect 29895 11625 29911 11659
rect 30079 11625 30095 11659
rect 30267 11625 30283 11659
rect 30451 11625 30467 11659
rect 18689 11566 18723 11582
rect 18689 11174 18723 11190
rect 18947 11566 18981 11582
rect 18947 11174 18981 11190
rect 19061 11566 19095 11582
rect 19061 11174 19095 11190
rect 19319 11566 19353 11582
rect 19319 11174 19353 11190
rect 19433 11566 19467 11582
rect 19433 11174 19467 11190
rect 19691 11566 19725 11582
rect 19691 11174 19725 11190
rect 19805 11566 19839 11582
rect 19805 11174 19839 11190
rect 20063 11566 20097 11582
rect 20063 11174 20097 11190
rect 20177 11566 20211 11582
rect 20177 11174 20211 11190
rect 20435 11566 20469 11582
rect 20435 11174 20469 11190
rect 20549 11566 20583 11582
rect 20549 11174 20583 11190
rect 20807 11566 20841 11582
rect 20807 11174 20841 11190
rect 20921 11566 20955 11582
rect 20921 11174 20955 11190
rect 21179 11566 21213 11582
rect 21179 11174 21213 11190
rect 21293 11566 21327 11582
rect 21293 11174 21327 11190
rect 21551 11566 21585 11582
rect 21551 11174 21585 11190
rect 21665 11566 21699 11582
rect 21665 11174 21699 11190
rect 21923 11566 21957 11582
rect 21923 11174 21957 11190
rect 22037 11566 22071 11582
rect 22037 11174 22071 11190
rect 22295 11566 22329 11582
rect 22295 11174 22329 11190
rect 22409 11566 22443 11582
rect 22409 11174 22443 11190
rect 22667 11566 22701 11582
rect 22667 11174 22701 11190
rect 22781 11566 22815 11582
rect 22781 11174 22815 11190
rect 23039 11566 23073 11582
rect 23039 11174 23073 11190
rect 23153 11566 23187 11582
rect 23153 11174 23187 11190
rect 23411 11566 23445 11582
rect 23411 11174 23445 11190
rect 23525 11566 23559 11582
rect 23525 11174 23559 11190
rect 23783 11566 23817 11582
rect 23783 11174 23817 11190
rect 23897 11566 23931 11582
rect 23897 11174 23931 11190
rect 24155 11566 24189 11582
rect 24155 11174 24189 11190
rect 24269 11566 24303 11582
rect 24269 11174 24303 11190
rect 24527 11566 24561 11582
rect 24527 11174 24561 11190
rect 24641 11566 24675 11582
rect 24641 11174 24675 11190
rect 24899 11566 24933 11582
rect 24899 11174 24933 11190
rect 25013 11566 25047 11582
rect 25013 11174 25047 11190
rect 25271 11566 25305 11582
rect 25271 11174 25305 11190
rect 25385 11566 25419 11582
rect 25385 11174 25419 11190
rect 25643 11566 25677 11582
rect 25643 11174 25677 11190
rect 25757 11566 25791 11582
rect 25757 11174 25791 11190
rect 26015 11566 26049 11582
rect 26015 11174 26049 11190
rect 26129 11566 26163 11582
rect 26129 11174 26163 11190
rect 26387 11566 26421 11582
rect 26387 11174 26421 11190
rect 26501 11566 26535 11582
rect 26501 11174 26535 11190
rect 26759 11566 26793 11582
rect 26759 11174 26793 11190
rect 26873 11566 26907 11582
rect 26873 11174 26907 11190
rect 27131 11566 27165 11582
rect 27131 11174 27165 11190
rect 27245 11566 27279 11582
rect 27245 11174 27279 11190
rect 27503 11566 27537 11582
rect 27503 11174 27537 11190
rect 27617 11566 27651 11582
rect 27617 11174 27651 11190
rect 27875 11566 27909 11582
rect 27875 11174 27909 11190
rect 27989 11566 28023 11582
rect 27989 11174 28023 11190
rect 28247 11566 28281 11582
rect 28247 11174 28281 11190
rect 28361 11566 28395 11582
rect 28361 11174 28395 11190
rect 28619 11566 28653 11582
rect 28619 11174 28653 11190
rect 28733 11566 28767 11582
rect 28733 11174 28767 11190
rect 28991 11566 29025 11582
rect 28991 11174 29025 11190
rect 29105 11566 29139 11582
rect 29105 11174 29139 11190
rect 29363 11566 29397 11582
rect 29363 11174 29397 11190
rect 29477 11566 29511 11582
rect 29477 11174 29511 11190
rect 29735 11566 29769 11582
rect 29735 11174 29769 11190
rect 29849 11566 29883 11582
rect 29849 11174 29883 11190
rect 30107 11566 30141 11582
rect 30107 11174 30141 11190
rect 30221 11566 30255 11582
rect 30221 11174 30255 11190
rect 30479 11566 30513 11582
rect 30479 11174 30513 11190
rect 18735 11097 18751 11131
rect 18919 11097 18935 11131
rect 19107 11097 19123 11131
rect 19291 11097 19307 11131
rect 19479 11097 19495 11131
rect 19663 11097 19679 11131
rect 19851 11097 19867 11131
rect 20035 11097 20051 11131
rect 20223 11097 20239 11131
rect 20407 11097 20423 11131
rect 20595 11097 20611 11131
rect 20779 11097 20795 11131
rect 20967 11097 20983 11131
rect 21151 11097 21167 11131
rect 21339 11097 21355 11131
rect 21523 11097 21539 11131
rect 21711 11097 21727 11131
rect 21895 11097 21911 11131
rect 22083 11097 22099 11131
rect 22267 11097 22283 11131
rect 22455 11097 22471 11131
rect 22639 11097 22655 11131
rect 22827 11097 22843 11131
rect 23011 11097 23027 11131
rect 23199 11097 23215 11131
rect 23383 11097 23399 11131
rect 23571 11097 23587 11131
rect 23755 11097 23771 11131
rect 23943 11097 23959 11131
rect 24127 11097 24143 11131
rect 24315 11097 24331 11131
rect 24499 11097 24515 11131
rect 24687 11097 24703 11131
rect 24871 11097 24887 11131
rect 25059 11097 25075 11131
rect 25243 11097 25259 11131
rect 25431 11097 25447 11131
rect 25615 11097 25631 11131
rect 25803 11097 25819 11131
rect 25987 11097 26003 11131
rect 26175 11097 26191 11131
rect 26359 11097 26375 11131
rect 26547 11097 26563 11131
rect 26731 11097 26747 11131
rect 26919 11097 26935 11131
rect 27103 11097 27119 11131
rect 27291 11097 27307 11131
rect 27475 11097 27491 11131
rect 27663 11097 27679 11131
rect 27847 11097 27863 11131
rect 28035 11097 28051 11131
rect 28219 11097 28235 11131
rect 28407 11097 28423 11131
rect 28591 11097 28607 11131
rect 28779 11097 28795 11131
rect 28963 11097 28979 11131
rect 29151 11097 29167 11131
rect 29335 11097 29351 11131
rect 29523 11097 29539 11131
rect 29707 11097 29723 11131
rect 29895 11097 29911 11131
rect 30079 11097 30095 11131
rect 30267 11097 30283 11131
rect 30451 11097 30467 11131
rect 18735 10989 18751 11023
rect 18919 10989 18935 11023
rect 19107 10989 19123 11023
rect 19291 10989 19307 11023
rect 19479 10989 19495 11023
rect 19663 10989 19679 11023
rect 19851 10989 19867 11023
rect 20035 10989 20051 11023
rect 20223 10989 20239 11023
rect 20407 10989 20423 11023
rect 20595 10989 20611 11023
rect 20779 10989 20795 11023
rect 20967 10989 20983 11023
rect 21151 10989 21167 11023
rect 21339 10989 21355 11023
rect 21523 10989 21539 11023
rect 21711 10989 21727 11023
rect 21895 10989 21911 11023
rect 22083 10989 22099 11023
rect 22267 10989 22283 11023
rect 22455 10989 22471 11023
rect 22639 10989 22655 11023
rect 22827 10989 22843 11023
rect 23011 10989 23027 11023
rect 23199 10989 23215 11023
rect 23383 10989 23399 11023
rect 23571 10989 23587 11023
rect 23755 10989 23771 11023
rect 23943 10989 23959 11023
rect 24127 10989 24143 11023
rect 24315 10989 24331 11023
rect 24499 10989 24515 11023
rect 24687 10989 24703 11023
rect 24871 10989 24887 11023
rect 25059 10989 25075 11023
rect 25243 10989 25259 11023
rect 25431 10989 25447 11023
rect 25615 10989 25631 11023
rect 25803 10989 25819 11023
rect 25987 10989 26003 11023
rect 26175 10989 26191 11023
rect 26359 10989 26375 11023
rect 26547 10989 26563 11023
rect 26731 10989 26747 11023
rect 26919 10989 26935 11023
rect 27103 10989 27119 11023
rect 27291 10989 27307 11023
rect 27475 10989 27491 11023
rect 27663 10989 27679 11023
rect 27847 10989 27863 11023
rect 28035 10989 28051 11023
rect 28219 10989 28235 11023
rect 28407 10989 28423 11023
rect 28591 10989 28607 11023
rect 28779 10989 28795 11023
rect 28963 10989 28979 11023
rect 29151 10989 29167 11023
rect 29335 10989 29351 11023
rect 29523 10989 29539 11023
rect 29707 10989 29723 11023
rect 29895 10989 29911 11023
rect 30079 10989 30095 11023
rect 30267 10989 30283 11023
rect 30451 10989 30467 11023
rect 18689 10930 18723 10946
rect 18689 10538 18723 10554
rect 18947 10930 18981 10946
rect 18947 10538 18981 10554
rect 19061 10930 19095 10946
rect 19061 10538 19095 10554
rect 19319 10930 19353 10946
rect 19319 10538 19353 10554
rect 19433 10930 19467 10946
rect 19433 10538 19467 10554
rect 19691 10930 19725 10946
rect 19691 10538 19725 10554
rect 19805 10930 19839 10946
rect 19805 10538 19839 10554
rect 20063 10930 20097 10946
rect 20063 10538 20097 10554
rect 20177 10930 20211 10946
rect 20177 10538 20211 10554
rect 20435 10930 20469 10946
rect 20435 10538 20469 10554
rect 20549 10930 20583 10946
rect 20549 10538 20583 10554
rect 20807 10930 20841 10946
rect 20807 10538 20841 10554
rect 20921 10930 20955 10946
rect 20921 10538 20955 10554
rect 21179 10930 21213 10946
rect 21179 10538 21213 10554
rect 21293 10930 21327 10946
rect 21293 10538 21327 10554
rect 21551 10930 21585 10946
rect 21551 10538 21585 10554
rect 21665 10930 21699 10946
rect 21665 10538 21699 10554
rect 21923 10930 21957 10946
rect 21923 10538 21957 10554
rect 22037 10930 22071 10946
rect 22037 10538 22071 10554
rect 22295 10930 22329 10946
rect 22295 10538 22329 10554
rect 22409 10930 22443 10946
rect 22409 10538 22443 10554
rect 22667 10930 22701 10946
rect 22667 10538 22701 10554
rect 22781 10930 22815 10946
rect 22781 10538 22815 10554
rect 23039 10930 23073 10946
rect 23039 10538 23073 10554
rect 23153 10930 23187 10946
rect 23153 10538 23187 10554
rect 23411 10930 23445 10946
rect 23411 10538 23445 10554
rect 23525 10930 23559 10946
rect 23525 10538 23559 10554
rect 23783 10930 23817 10946
rect 23783 10538 23817 10554
rect 23897 10930 23931 10946
rect 23897 10538 23931 10554
rect 24155 10930 24189 10946
rect 24155 10538 24189 10554
rect 24269 10930 24303 10946
rect 24269 10538 24303 10554
rect 24527 10930 24561 10946
rect 24527 10538 24561 10554
rect 24641 10930 24675 10946
rect 24641 10538 24675 10554
rect 24899 10930 24933 10946
rect 24899 10538 24933 10554
rect 25013 10930 25047 10946
rect 25013 10538 25047 10554
rect 25271 10930 25305 10946
rect 25271 10538 25305 10554
rect 25385 10930 25419 10946
rect 25385 10538 25419 10554
rect 25643 10930 25677 10946
rect 25643 10538 25677 10554
rect 25757 10930 25791 10946
rect 25757 10538 25791 10554
rect 26015 10930 26049 10946
rect 26015 10538 26049 10554
rect 26129 10930 26163 10946
rect 26129 10538 26163 10554
rect 26387 10930 26421 10946
rect 26387 10538 26421 10554
rect 26501 10930 26535 10946
rect 26501 10538 26535 10554
rect 26759 10930 26793 10946
rect 26759 10538 26793 10554
rect 26873 10930 26907 10946
rect 26873 10538 26907 10554
rect 27131 10930 27165 10946
rect 27131 10538 27165 10554
rect 27245 10930 27279 10946
rect 27245 10538 27279 10554
rect 27503 10930 27537 10946
rect 27503 10538 27537 10554
rect 27617 10930 27651 10946
rect 27617 10538 27651 10554
rect 27875 10930 27909 10946
rect 27875 10538 27909 10554
rect 27989 10930 28023 10946
rect 27989 10538 28023 10554
rect 28247 10930 28281 10946
rect 28247 10538 28281 10554
rect 28361 10930 28395 10946
rect 28361 10538 28395 10554
rect 28619 10930 28653 10946
rect 28619 10538 28653 10554
rect 28733 10930 28767 10946
rect 28733 10538 28767 10554
rect 28991 10930 29025 10946
rect 28991 10538 29025 10554
rect 29105 10930 29139 10946
rect 29105 10538 29139 10554
rect 29363 10930 29397 10946
rect 29363 10538 29397 10554
rect 29477 10930 29511 10946
rect 29477 10538 29511 10554
rect 29735 10930 29769 10946
rect 29735 10538 29769 10554
rect 29849 10930 29883 10946
rect 29849 10538 29883 10554
rect 30107 10930 30141 10946
rect 30107 10538 30141 10554
rect 30221 10930 30255 10946
rect 30221 10538 30255 10554
rect 30479 10930 30513 10946
rect 30479 10538 30513 10554
rect 18735 10461 18751 10495
rect 18919 10461 18935 10495
rect 19107 10461 19123 10495
rect 19291 10461 19307 10495
rect 19479 10461 19495 10495
rect 19663 10461 19679 10495
rect 19851 10461 19867 10495
rect 20035 10461 20051 10495
rect 20223 10461 20239 10495
rect 20407 10461 20423 10495
rect 20595 10461 20611 10495
rect 20779 10461 20795 10495
rect 20967 10461 20983 10495
rect 21151 10461 21167 10495
rect 21339 10461 21355 10495
rect 21523 10461 21539 10495
rect 21711 10461 21727 10495
rect 21895 10461 21911 10495
rect 22083 10461 22099 10495
rect 22267 10461 22283 10495
rect 22455 10461 22471 10495
rect 22639 10461 22655 10495
rect 22827 10461 22843 10495
rect 23011 10461 23027 10495
rect 23199 10461 23215 10495
rect 23383 10461 23399 10495
rect 23571 10461 23587 10495
rect 23755 10461 23771 10495
rect 23943 10461 23959 10495
rect 24127 10461 24143 10495
rect 24315 10461 24331 10495
rect 24499 10461 24515 10495
rect 24687 10461 24703 10495
rect 24871 10461 24887 10495
rect 25059 10461 25075 10495
rect 25243 10461 25259 10495
rect 25431 10461 25447 10495
rect 25615 10461 25631 10495
rect 25803 10461 25819 10495
rect 25987 10461 26003 10495
rect 26175 10461 26191 10495
rect 26359 10461 26375 10495
rect 26547 10461 26563 10495
rect 26731 10461 26747 10495
rect 26919 10461 26935 10495
rect 27103 10461 27119 10495
rect 27291 10461 27307 10495
rect 27475 10461 27491 10495
rect 27663 10461 27679 10495
rect 27847 10461 27863 10495
rect 28035 10461 28051 10495
rect 28219 10461 28235 10495
rect 28407 10461 28423 10495
rect 28591 10461 28607 10495
rect 28779 10461 28795 10495
rect 28963 10461 28979 10495
rect 29151 10461 29167 10495
rect 29335 10461 29351 10495
rect 29523 10461 29539 10495
rect 29707 10461 29723 10495
rect 29895 10461 29911 10495
rect 30079 10461 30095 10495
rect 30267 10461 30283 10495
rect 30451 10461 30467 10495
rect 18735 10353 18751 10387
rect 18919 10353 18935 10387
rect 19107 10353 19123 10387
rect 19291 10353 19307 10387
rect 19479 10353 19495 10387
rect 19663 10353 19679 10387
rect 19851 10353 19867 10387
rect 20035 10353 20051 10387
rect 20223 10353 20239 10387
rect 20407 10353 20423 10387
rect 20595 10353 20611 10387
rect 20779 10353 20795 10387
rect 20967 10353 20983 10387
rect 21151 10353 21167 10387
rect 21339 10353 21355 10387
rect 21523 10353 21539 10387
rect 21711 10353 21727 10387
rect 21895 10353 21911 10387
rect 22083 10353 22099 10387
rect 22267 10353 22283 10387
rect 22455 10353 22471 10387
rect 22639 10353 22655 10387
rect 22827 10353 22843 10387
rect 23011 10353 23027 10387
rect 23199 10353 23215 10387
rect 23383 10353 23399 10387
rect 23571 10353 23587 10387
rect 23755 10353 23771 10387
rect 23943 10353 23959 10387
rect 24127 10353 24143 10387
rect 24315 10353 24331 10387
rect 24499 10353 24515 10387
rect 24687 10353 24703 10387
rect 24871 10353 24887 10387
rect 25059 10353 25075 10387
rect 25243 10353 25259 10387
rect 25431 10353 25447 10387
rect 25615 10353 25631 10387
rect 25803 10353 25819 10387
rect 25987 10353 26003 10387
rect 26175 10353 26191 10387
rect 26359 10353 26375 10387
rect 26547 10353 26563 10387
rect 26731 10353 26747 10387
rect 26919 10353 26935 10387
rect 27103 10353 27119 10387
rect 27291 10353 27307 10387
rect 27475 10353 27491 10387
rect 27663 10353 27679 10387
rect 27847 10353 27863 10387
rect 28035 10353 28051 10387
rect 28219 10353 28235 10387
rect 28407 10353 28423 10387
rect 28591 10353 28607 10387
rect 28779 10353 28795 10387
rect 28963 10353 28979 10387
rect 29151 10353 29167 10387
rect 29335 10353 29351 10387
rect 29523 10353 29539 10387
rect 29707 10353 29723 10387
rect 29895 10353 29911 10387
rect 30079 10353 30095 10387
rect 30267 10353 30283 10387
rect 30451 10353 30467 10387
rect 18689 10294 18723 10310
rect 18689 9902 18723 9918
rect 18947 10294 18981 10310
rect 18947 9902 18981 9918
rect 19061 10294 19095 10310
rect 19061 9902 19095 9918
rect 19319 10294 19353 10310
rect 19319 9902 19353 9918
rect 19433 10294 19467 10310
rect 19433 9902 19467 9918
rect 19691 10294 19725 10310
rect 19691 9902 19725 9918
rect 19805 10294 19839 10310
rect 19805 9902 19839 9918
rect 20063 10294 20097 10310
rect 20063 9902 20097 9918
rect 20177 10294 20211 10310
rect 20177 9902 20211 9918
rect 20435 10294 20469 10310
rect 20435 9902 20469 9918
rect 20549 10294 20583 10310
rect 20549 9902 20583 9918
rect 20807 10294 20841 10310
rect 20807 9902 20841 9918
rect 20921 10294 20955 10310
rect 20921 9902 20955 9918
rect 21179 10294 21213 10310
rect 21179 9902 21213 9918
rect 21293 10294 21327 10310
rect 21293 9902 21327 9918
rect 21551 10294 21585 10310
rect 21551 9902 21585 9918
rect 21665 10294 21699 10310
rect 21665 9902 21699 9918
rect 21923 10294 21957 10310
rect 21923 9902 21957 9918
rect 22037 10294 22071 10310
rect 22037 9902 22071 9918
rect 22295 10294 22329 10310
rect 22295 9902 22329 9918
rect 22409 10294 22443 10310
rect 22409 9902 22443 9918
rect 22667 10294 22701 10310
rect 22667 9902 22701 9918
rect 22781 10294 22815 10310
rect 22781 9902 22815 9918
rect 23039 10294 23073 10310
rect 23039 9902 23073 9918
rect 23153 10294 23187 10310
rect 23153 9902 23187 9918
rect 23411 10294 23445 10310
rect 23411 9902 23445 9918
rect 23525 10294 23559 10310
rect 23525 9902 23559 9918
rect 23783 10294 23817 10310
rect 23783 9902 23817 9918
rect 23897 10294 23931 10310
rect 23897 9902 23931 9918
rect 24155 10294 24189 10310
rect 24155 9902 24189 9918
rect 24269 10294 24303 10310
rect 24269 9902 24303 9918
rect 24527 10294 24561 10310
rect 24527 9902 24561 9918
rect 24641 10294 24675 10310
rect 24641 9902 24675 9918
rect 24899 10294 24933 10310
rect 24899 9902 24933 9918
rect 25013 10294 25047 10310
rect 25013 9902 25047 9918
rect 25271 10294 25305 10310
rect 25271 9902 25305 9918
rect 25385 10294 25419 10310
rect 25385 9902 25419 9918
rect 25643 10294 25677 10310
rect 25643 9902 25677 9918
rect 25757 10294 25791 10310
rect 25757 9902 25791 9918
rect 26015 10294 26049 10310
rect 26015 9902 26049 9918
rect 26129 10294 26163 10310
rect 26129 9902 26163 9918
rect 26387 10294 26421 10310
rect 26387 9902 26421 9918
rect 26501 10294 26535 10310
rect 26501 9902 26535 9918
rect 26759 10294 26793 10310
rect 26759 9902 26793 9918
rect 26873 10294 26907 10310
rect 26873 9902 26907 9918
rect 27131 10294 27165 10310
rect 27131 9902 27165 9918
rect 27245 10294 27279 10310
rect 27245 9902 27279 9918
rect 27503 10294 27537 10310
rect 27503 9902 27537 9918
rect 27617 10294 27651 10310
rect 27617 9902 27651 9918
rect 27875 10294 27909 10310
rect 27875 9902 27909 9918
rect 27989 10294 28023 10310
rect 27989 9902 28023 9918
rect 28247 10294 28281 10310
rect 28247 9902 28281 9918
rect 28361 10294 28395 10310
rect 28361 9902 28395 9918
rect 28619 10294 28653 10310
rect 28619 9902 28653 9918
rect 28733 10294 28767 10310
rect 28733 9902 28767 9918
rect 28991 10294 29025 10310
rect 28991 9902 29025 9918
rect 29105 10294 29139 10310
rect 29105 9902 29139 9918
rect 29363 10294 29397 10310
rect 29363 9902 29397 9918
rect 29477 10294 29511 10310
rect 29477 9902 29511 9918
rect 29735 10294 29769 10310
rect 29735 9902 29769 9918
rect 29849 10294 29883 10310
rect 29849 9902 29883 9918
rect 30107 10294 30141 10310
rect 30107 9902 30141 9918
rect 30221 10294 30255 10310
rect 30221 9902 30255 9918
rect 30479 10294 30513 10310
rect 30479 9902 30513 9918
rect 18735 9825 18751 9859
rect 18919 9825 18935 9859
rect 19107 9825 19123 9859
rect 19291 9825 19307 9859
rect 19479 9825 19495 9859
rect 19663 9825 19679 9859
rect 19851 9825 19867 9859
rect 20035 9825 20051 9859
rect 20223 9825 20239 9859
rect 20407 9825 20423 9859
rect 20595 9825 20611 9859
rect 20779 9825 20795 9859
rect 20967 9825 20983 9859
rect 21151 9825 21167 9859
rect 21339 9825 21355 9859
rect 21523 9825 21539 9859
rect 21711 9825 21727 9859
rect 21895 9825 21911 9859
rect 22083 9825 22099 9859
rect 22267 9825 22283 9859
rect 22455 9825 22471 9859
rect 22639 9825 22655 9859
rect 22827 9825 22843 9859
rect 23011 9825 23027 9859
rect 23199 9825 23215 9859
rect 23383 9825 23399 9859
rect 23571 9825 23587 9859
rect 23755 9825 23771 9859
rect 23943 9825 23959 9859
rect 24127 9825 24143 9859
rect 24315 9825 24331 9859
rect 24499 9825 24515 9859
rect 24687 9825 24703 9859
rect 24871 9825 24887 9859
rect 25059 9825 25075 9859
rect 25243 9825 25259 9859
rect 25431 9825 25447 9859
rect 25615 9825 25631 9859
rect 25803 9825 25819 9859
rect 25987 9825 26003 9859
rect 26175 9825 26191 9859
rect 26359 9825 26375 9859
rect 26547 9825 26563 9859
rect 26731 9825 26747 9859
rect 26919 9825 26935 9859
rect 27103 9825 27119 9859
rect 27291 9825 27307 9859
rect 27475 9825 27491 9859
rect 27663 9825 27679 9859
rect 27847 9825 27863 9859
rect 28035 9825 28051 9859
rect 28219 9825 28235 9859
rect 28407 9825 28423 9859
rect 28591 9825 28607 9859
rect 28779 9825 28795 9859
rect 28963 9825 28979 9859
rect 29151 9825 29167 9859
rect 29335 9825 29351 9859
rect 29523 9825 29539 9859
rect 29707 9825 29723 9859
rect 29895 9825 29911 9859
rect 30079 9825 30095 9859
rect 30267 9825 30283 9859
rect 30451 9825 30467 9859
rect 18575 9757 18609 9819
rect 30593 9757 30627 9819
rect 18575 9723 18671 9757
rect 30531 9723 30627 9757
rect 20063 9339 20148 9373
rect 23091 9339 23187 9373
rect 20063 9277 20097 9339
rect 23153 9277 23187 9339
rect 20223 9237 20239 9271
rect 20407 9237 20423 9271
rect 20595 9237 20611 9271
rect 20779 9237 20795 9271
rect 20967 9237 20983 9271
rect 21151 9237 21167 9271
rect 21339 9237 21355 9271
rect 21523 9237 21539 9271
rect 21711 9237 21727 9271
rect 21895 9237 21911 9271
rect 22083 9237 22099 9271
rect 22267 9237 22283 9271
rect 22455 9237 22471 9271
rect 22639 9237 22655 9271
rect 22827 9237 22843 9271
rect 23011 9237 23027 9271
rect 20177 9178 20211 9194
rect 20177 8386 20211 8402
rect 20435 9178 20469 9194
rect 20435 8386 20469 8402
rect 20549 9178 20583 9194
rect 20549 8386 20583 8402
rect 20807 9178 20841 9194
rect 20807 8386 20841 8402
rect 20921 9178 20955 9194
rect 20921 8386 20955 8402
rect 21179 9178 21213 9194
rect 21179 8386 21213 8402
rect 21293 9178 21327 9194
rect 21293 8386 21327 8402
rect 21551 9178 21585 9194
rect 21551 8386 21585 8402
rect 21665 9178 21699 9194
rect 21665 8386 21699 8402
rect 21923 9178 21957 9194
rect 21923 8386 21957 8402
rect 22037 9178 22071 9194
rect 22037 8386 22071 8402
rect 22295 9178 22329 9194
rect 22295 8386 22329 8402
rect 22409 9178 22443 9194
rect 22409 8386 22443 8402
rect 22667 9178 22701 9194
rect 22667 8386 22701 8402
rect 22781 9178 22815 9194
rect 22781 8386 22815 8402
rect 23039 9178 23073 9194
rect 23039 8386 23073 8402
rect 20223 8309 20239 8343
rect 20407 8309 20423 8343
rect 20595 8309 20611 8343
rect 20779 8309 20795 8343
rect 20967 8309 20983 8343
rect 21151 8309 21167 8343
rect 21339 8309 21355 8343
rect 21523 8309 21539 8343
rect 21711 8309 21727 8343
rect 21895 8309 21911 8343
rect 22083 8309 22099 8343
rect 22267 8309 22283 8343
rect 22455 8309 22471 8343
rect 22639 8309 22655 8343
rect 22827 8309 22843 8343
rect 23011 8309 23027 8343
rect 20223 8201 20239 8235
rect 20407 8201 20423 8235
rect 20595 8201 20611 8235
rect 20779 8201 20795 8235
rect 20967 8201 20983 8235
rect 21151 8201 21167 8235
rect 21339 8201 21355 8235
rect 21523 8201 21539 8235
rect 21711 8201 21727 8235
rect 21895 8201 21911 8235
rect 22083 8201 22099 8235
rect 22267 8201 22283 8235
rect 22455 8201 22471 8235
rect 22639 8201 22655 8235
rect 22827 8201 22843 8235
rect 23011 8201 23027 8235
rect 20177 8142 20211 8158
rect 20177 7350 20211 7366
rect 20435 8142 20469 8158
rect 20435 7350 20469 7366
rect 20549 8142 20583 8158
rect 20549 7350 20583 7366
rect 20807 8142 20841 8158
rect 20807 7350 20841 7366
rect 20921 8142 20955 8158
rect 20921 7350 20955 7366
rect 21179 8142 21213 8158
rect 21179 7350 21213 7366
rect 21293 8142 21327 8158
rect 21293 7350 21327 7366
rect 21551 8142 21585 8158
rect 21551 7350 21585 7366
rect 21665 8142 21699 8158
rect 21665 7350 21699 7366
rect 21923 8142 21957 8158
rect 21923 7350 21957 7366
rect 22037 8142 22071 8158
rect 22037 7350 22071 7366
rect 22295 8142 22329 8158
rect 22295 7350 22329 7366
rect 22409 8142 22443 8158
rect 22409 7350 22443 7366
rect 22667 8142 22701 8158
rect 22667 7350 22701 7366
rect 22781 8142 22815 8158
rect 22781 7350 22815 7366
rect 23039 8142 23073 8158
rect 23039 7350 23073 7366
rect 20223 7273 20239 7307
rect 20407 7273 20423 7307
rect 20595 7273 20611 7307
rect 20779 7273 20795 7307
rect 20967 7273 20983 7307
rect 21151 7273 21167 7307
rect 21339 7273 21355 7307
rect 21523 7273 21539 7307
rect 21711 7273 21727 7307
rect 21895 7273 21911 7307
rect 22083 7273 22099 7307
rect 22267 7273 22283 7307
rect 22455 7273 22471 7307
rect 22639 7273 22655 7307
rect 22827 7273 22843 7307
rect 23011 7273 23027 7307
rect 20223 7165 20239 7199
rect 20407 7165 20423 7199
rect 20595 7165 20611 7199
rect 20779 7165 20795 7199
rect 20967 7165 20983 7199
rect 21151 7165 21167 7199
rect 21339 7165 21355 7199
rect 21523 7165 21539 7199
rect 21711 7165 21727 7199
rect 21895 7165 21911 7199
rect 22083 7165 22099 7199
rect 22267 7165 22283 7199
rect 22455 7165 22471 7199
rect 22639 7165 22655 7199
rect 22827 7165 22843 7199
rect 23011 7165 23027 7199
rect 20177 7106 20211 7122
rect 20177 6314 20211 6330
rect 20435 7106 20469 7122
rect 20435 6314 20469 6330
rect 20549 7106 20583 7122
rect 20549 6314 20583 6330
rect 20807 7106 20841 7122
rect 20807 6314 20841 6330
rect 20921 7106 20955 7122
rect 20921 6314 20955 6330
rect 21179 7106 21213 7122
rect 21179 6314 21213 6330
rect 21293 7106 21327 7122
rect 21293 6314 21327 6330
rect 21551 7106 21585 7122
rect 21551 6314 21585 6330
rect 21665 7106 21699 7122
rect 21665 6314 21699 6330
rect 21923 7106 21957 7122
rect 21923 6314 21957 6330
rect 22037 7106 22071 7122
rect 22037 6314 22071 6330
rect 22295 7106 22329 7122
rect 22295 6314 22329 6330
rect 22409 7106 22443 7122
rect 22409 6314 22443 6330
rect 22667 7106 22701 7122
rect 22667 6314 22701 6330
rect 22781 7106 22815 7122
rect 22781 6314 22815 6330
rect 23039 7106 23073 7122
rect 23039 6314 23073 6330
rect 20223 6237 20239 6271
rect 20407 6237 20423 6271
rect 20595 6237 20611 6271
rect 20779 6237 20795 6271
rect 20967 6237 20983 6271
rect 21151 6237 21167 6271
rect 21339 6237 21355 6271
rect 21523 6237 21539 6271
rect 21711 6237 21727 6271
rect 21895 6237 21911 6271
rect 22083 6237 22099 6271
rect 22267 6237 22283 6271
rect 22455 6237 22471 6271
rect 22639 6237 22655 6271
rect 22827 6237 22843 6271
rect 23011 6237 23027 6271
rect 20223 6129 20239 6163
rect 20407 6129 20423 6163
rect 20595 6129 20611 6163
rect 20779 6129 20795 6163
rect 20967 6129 20983 6163
rect 21151 6129 21167 6163
rect 21339 6129 21355 6163
rect 21523 6129 21539 6163
rect 21711 6129 21727 6163
rect 21895 6129 21911 6163
rect 22083 6129 22099 6163
rect 22267 6129 22283 6163
rect 22455 6129 22471 6163
rect 22639 6129 22655 6163
rect 22827 6129 22843 6163
rect 23011 6129 23027 6163
rect 20177 6070 20211 6086
rect 20177 5278 20211 5294
rect 20435 6070 20469 6086
rect 20435 5278 20469 5294
rect 20549 6070 20583 6086
rect 20549 5278 20583 5294
rect 20807 6070 20841 6086
rect 20807 5278 20841 5294
rect 20921 6070 20955 6086
rect 20921 5278 20955 5294
rect 21179 6070 21213 6086
rect 21179 5278 21213 5294
rect 21293 6070 21327 6086
rect 21293 5278 21327 5294
rect 21551 6070 21585 6086
rect 21551 5278 21585 5294
rect 21665 6070 21699 6086
rect 21665 5278 21699 5294
rect 21923 6070 21957 6086
rect 21923 5278 21957 5294
rect 22037 6070 22071 6086
rect 22037 5278 22071 5294
rect 22295 6070 22329 6086
rect 22295 5278 22329 5294
rect 22409 6070 22443 6086
rect 22409 5278 22443 5294
rect 22667 6070 22701 6086
rect 22667 5278 22701 5294
rect 22781 6070 22815 6086
rect 22781 5278 22815 5294
rect 23039 6070 23073 6086
rect 23039 5278 23073 5294
rect 20223 5201 20239 5235
rect 20407 5201 20423 5235
rect 20595 5201 20611 5235
rect 20779 5201 20795 5235
rect 20967 5201 20983 5235
rect 21151 5201 21167 5235
rect 21339 5201 21355 5235
rect 21523 5201 21539 5235
rect 21711 5201 21727 5235
rect 21895 5201 21911 5235
rect 22083 5201 22099 5235
rect 22267 5201 22283 5235
rect 22455 5201 22471 5235
rect 22639 5201 22655 5235
rect 22827 5201 22843 5235
rect 23011 5201 23027 5235
rect 20063 5133 20097 5195
rect 23689 7425 23785 7459
rect 23923 7425 24019 7459
rect 23689 7363 23723 7425
rect 23985 7363 24019 7425
rect 23689 5809 23723 5871
rect 23985 5809 24019 5871
rect 23689 5775 23785 5809
rect 23923 5775 24019 5809
rect 23153 5133 23187 5195
rect 20063 5099 20159 5133
rect 23091 5099 23187 5133
rect 20063 4645 20159 4679
rect 29043 4645 29139 4679
rect 20063 4583 20097 4645
rect 29105 4583 29139 4645
rect 20223 4543 20239 4577
rect 20407 4543 20423 4577
rect 20595 4543 20611 4577
rect 20779 4543 20795 4577
rect 20967 4543 20983 4577
rect 21151 4543 21167 4577
rect 21339 4543 21355 4577
rect 21523 4543 21539 4577
rect 21711 4543 21727 4577
rect 21895 4543 21911 4577
rect 22083 4543 22099 4577
rect 22267 4543 22283 4577
rect 22455 4543 22471 4577
rect 22639 4543 22655 4577
rect 22827 4543 22843 4577
rect 23011 4543 23027 4577
rect 23199 4543 23215 4577
rect 23383 4543 23399 4577
rect 23571 4543 23587 4577
rect 23755 4543 23771 4577
rect 23943 4543 23959 4577
rect 24127 4543 24143 4577
rect 24315 4543 24331 4577
rect 24499 4543 24515 4577
rect 24687 4543 24703 4577
rect 24871 4543 24887 4577
rect 25059 4543 25075 4577
rect 25243 4543 25259 4577
rect 25431 4543 25447 4577
rect 25615 4543 25631 4577
rect 25803 4543 25819 4577
rect 25987 4543 26003 4577
rect 26175 4543 26191 4577
rect 26359 4543 26375 4577
rect 26547 4543 26563 4577
rect 26731 4543 26747 4577
rect 26919 4543 26935 4577
rect 27103 4543 27119 4577
rect 27291 4543 27307 4577
rect 27475 4543 27491 4577
rect 27663 4543 27679 4577
rect 27847 4543 27863 4577
rect 28035 4543 28051 4577
rect 28219 4543 28235 4577
rect 28407 4543 28423 4577
rect 28591 4543 28607 4577
rect 28779 4543 28795 4577
rect 28963 4543 28979 4577
rect 20177 4493 20211 4509
rect 20177 4301 20211 4317
rect 20435 4493 20469 4509
rect 20435 4301 20469 4317
rect 20549 4493 20583 4509
rect 20549 4301 20583 4317
rect 20807 4493 20841 4509
rect 20807 4301 20841 4317
rect 20921 4493 20955 4509
rect 20921 4301 20955 4317
rect 21179 4493 21213 4509
rect 21179 4301 21213 4317
rect 21293 4493 21327 4509
rect 21293 4301 21327 4317
rect 21551 4493 21585 4509
rect 21551 4301 21585 4317
rect 21665 4493 21699 4509
rect 21665 4301 21699 4317
rect 21923 4493 21957 4509
rect 21923 4301 21957 4317
rect 22037 4493 22071 4509
rect 22037 4301 22071 4317
rect 22295 4493 22329 4509
rect 22295 4301 22329 4317
rect 22409 4493 22443 4509
rect 22409 4301 22443 4317
rect 22667 4493 22701 4509
rect 22667 4301 22701 4317
rect 22781 4493 22815 4509
rect 22781 4301 22815 4317
rect 23039 4493 23073 4509
rect 23039 4301 23073 4317
rect 23153 4493 23187 4509
rect 23153 4301 23187 4317
rect 23411 4493 23445 4509
rect 23411 4301 23445 4317
rect 23525 4493 23559 4509
rect 23525 4301 23559 4317
rect 23783 4493 23817 4509
rect 23783 4301 23817 4317
rect 23897 4493 23931 4509
rect 23897 4301 23931 4317
rect 24155 4493 24189 4509
rect 24155 4301 24189 4317
rect 24269 4493 24303 4509
rect 24269 4301 24303 4317
rect 24527 4493 24561 4509
rect 24527 4301 24561 4317
rect 24641 4493 24675 4509
rect 24641 4301 24675 4317
rect 24899 4493 24933 4509
rect 24899 4301 24933 4317
rect 25013 4493 25047 4509
rect 25013 4301 25047 4317
rect 25271 4493 25305 4509
rect 25271 4301 25305 4317
rect 25385 4493 25419 4509
rect 25385 4301 25419 4317
rect 25643 4493 25677 4509
rect 25643 4301 25677 4317
rect 25757 4493 25791 4509
rect 25757 4301 25791 4317
rect 26015 4493 26049 4509
rect 26015 4301 26049 4317
rect 26129 4493 26163 4509
rect 26129 4301 26163 4317
rect 26387 4493 26421 4509
rect 26387 4301 26421 4317
rect 26501 4493 26535 4509
rect 26501 4301 26535 4317
rect 26759 4493 26793 4509
rect 26759 4301 26793 4317
rect 26873 4493 26907 4509
rect 26873 4301 26907 4317
rect 27131 4493 27165 4509
rect 27131 4301 27165 4317
rect 27245 4493 27279 4509
rect 27245 4301 27279 4317
rect 27503 4493 27537 4509
rect 27503 4301 27537 4317
rect 27617 4493 27651 4509
rect 27617 4301 27651 4317
rect 27875 4493 27909 4509
rect 27875 4301 27909 4317
rect 27989 4493 28023 4509
rect 27989 4301 28023 4317
rect 28247 4493 28281 4509
rect 28247 4301 28281 4317
rect 28361 4493 28395 4509
rect 28361 4301 28395 4317
rect 28619 4493 28653 4509
rect 28619 4301 28653 4317
rect 28733 4493 28767 4509
rect 28733 4301 28767 4317
rect 28991 4493 29025 4509
rect 28991 4301 29025 4317
rect 20223 4233 20239 4267
rect 20407 4233 20423 4267
rect 20595 4233 20611 4267
rect 20779 4233 20795 4267
rect 20967 4233 20983 4267
rect 21151 4233 21167 4267
rect 21339 4233 21355 4267
rect 21523 4233 21539 4267
rect 21711 4233 21727 4267
rect 21895 4233 21911 4267
rect 22083 4233 22099 4267
rect 22267 4233 22283 4267
rect 22455 4233 22471 4267
rect 22639 4233 22655 4267
rect 22827 4233 22843 4267
rect 23011 4233 23027 4267
rect 23199 4233 23215 4267
rect 23383 4233 23399 4267
rect 23571 4233 23587 4267
rect 23755 4233 23771 4267
rect 23943 4233 23959 4267
rect 24127 4233 24143 4267
rect 24315 4233 24331 4267
rect 24499 4233 24515 4267
rect 24687 4233 24703 4267
rect 24871 4233 24887 4267
rect 25059 4233 25075 4267
rect 25243 4233 25259 4267
rect 25431 4233 25447 4267
rect 25615 4233 25631 4267
rect 25803 4233 25819 4267
rect 25987 4233 26003 4267
rect 26175 4233 26191 4267
rect 26359 4233 26375 4267
rect 26547 4233 26563 4267
rect 26731 4233 26747 4267
rect 26919 4233 26935 4267
rect 27103 4233 27119 4267
rect 27291 4233 27307 4267
rect 27475 4233 27491 4267
rect 27663 4233 27679 4267
rect 27847 4233 27863 4267
rect 28035 4233 28051 4267
rect 28219 4233 28235 4267
rect 28407 4233 28423 4267
rect 28591 4233 28607 4267
rect 28779 4233 28795 4267
rect 28963 4233 28979 4267
rect 20223 4125 20239 4159
rect 20407 4125 20423 4159
rect 20595 4125 20611 4159
rect 20779 4125 20795 4159
rect 20967 4125 20983 4159
rect 21151 4125 21167 4159
rect 21339 4125 21355 4159
rect 21523 4125 21539 4159
rect 21711 4125 21727 4159
rect 21895 4125 21911 4159
rect 22083 4125 22099 4159
rect 22267 4125 22283 4159
rect 22455 4125 22471 4159
rect 22639 4125 22655 4159
rect 22827 4125 22843 4159
rect 23011 4125 23027 4159
rect 23199 4125 23215 4159
rect 23383 4125 23399 4159
rect 23571 4125 23587 4159
rect 23755 4125 23771 4159
rect 23943 4125 23959 4159
rect 24127 4125 24143 4159
rect 24315 4125 24331 4159
rect 24499 4125 24515 4159
rect 24687 4125 24703 4159
rect 24871 4125 24887 4159
rect 25059 4125 25075 4159
rect 25243 4125 25259 4159
rect 25431 4125 25447 4159
rect 25615 4125 25631 4159
rect 25803 4125 25819 4159
rect 25987 4125 26003 4159
rect 26175 4125 26191 4159
rect 26359 4125 26375 4159
rect 26547 4125 26563 4159
rect 26731 4125 26747 4159
rect 26919 4125 26935 4159
rect 27103 4125 27119 4159
rect 27291 4125 27307 4159
rect 27475 4125 27491 4159
rect 27663 4125 27679 4159
rect 27847 4125 27863 4159
rect 28035 4125 28051 4159
rect 28219 4125 28235 4159
rect 28407 4125 28423 4159
rect 28591 4125 28607 4159
rect 28779 4125 28795 4159
rect 28963 4125 28979 4159
rect 20177 4075 20211 4091
rect 20177 3883 20211 3899
rect 20435 4075 20469 4091
rect 20435 3883 20469 3899
rect 20549 4075 20583 4091
rect 20549 3883 20583 3899
rect 20807 4075 20841 4091
rect 20807 3883 20841 3899
rect 20921 4075 20955 4091
rect 20921 3883 20955 3899
rect 21179 4075 21213 4091
rect 21179 3883 21213 3899
rect 21293 4075 21327 4091
rect 21293 3883 21327 3899
rect 21551 4075 21585 4091
rect 21551 3883 21585 3899
rect 21665 4075 21699 4091
rect 21665 3883 21699 3899
rect 21923 4075 21957 4091
rect 21923 3883 21957 3899
rect 22037 4075 22071 4091
rect 22037 3883 22071 3899
rect 22295 4075 22329 4091
rect 22295 3883 22329 3899
rect 22409 4075 22443 4091
rect 22409 3883 22443 3899
rect 22667 4075 22701 4091
rect 22667 3883 22701 3899
rect 22781 4075 22815 4091
rect 22781 3883 22815 3899
rect 23039 4075 23073 4091
rect 23039 3883 23073 3899
rect 23153 4075 23187 4091
rect 23153 3883 23187 3899
rect 23411 4075 23445 4091
rect 23411 3883 23445 3899
rect 23525 4075 23559 4091
rect 23525 3883 23559 3899
rect 23783 4075 23817 4091
rect 23783 3883 23817 3899
rect 23897 4075 23931 4091
rect 23897 3883 23931 3899
rect 24155 4075 24189 4091
rect 24155 3883 24189 3899
rect 24269 4075 24303 4091
rect 24269 3883 24303 3899
rect 24527 4075 24561 4091
rect 24527 3883 24561 3899
rect 24641 4075 24675 4091
rect 24641 3883 24675 3899
rect 24899 4075 24933 4091
rect 24899 3883 24933 3899
rect 25013 4075 25047 4091
rect 25013 3883 25047 3899
rect 25271 4075 25305 4091
rect 25271 3883 25305 3899
rect 25385 4075 25419 4091
rect 25385 3883 25419 3899
rect 25643 4075 25677 4091
rect 25643 3883 25677 3899
rect 25757 4075 25791 4091
rect 25757 3883 25791 3899
rect 26015 4075 26049 4091
rect 26015 3883 26049 3899
rect 26129 4075 26163 4091
rect 26129 3883 26163 3899
rect 26387 4075 26421 4091
rect 26387 3883 26421 3899
rect 26501 4075 26535 4091
rect 26501 3883 26535 3899
rect 26759 4075 26793 4091
rect 26759 3883 26793 3899
rect 26873 4075 26907 4091
rect 26873 3883 26907 3899
rect 27131 4075 27165 4091
rect 27131 3883 27165 3899
rect 27245 4075 27279 4091
rect 27245 3883 27279 3899
rect 27503 4075 27537 4091
rect 27503 3883 27537 3899
rect 27617 4075 27651 4091
rect 27617 3883 27651 3899
rect 27875 4075 27909 4091
rect 27875 3883 27909 3899
rect 27989 4075 28023 4091
rect 27989 3883 28023 3899
rect 28247 4075 28281 4091
rect 28247 3883 28281 3899
rect 28361 4075 28395 4091
rect 28361 3883 28395 3899
rect 28619 4075 28653 4091
rect 28619 3883 28653 3899
rect 28733 4075 28767 4091
rect 28733 3883 28767 3899
rect 28991 4075 29025 4091
rect 28991 3883 29025 3899
rect 20223 3815 20239 3849
rect 20407 3815 20423 3849
rect 20595 3815 20611 3849
rect 20779 3815 20795 3849
rect 20967 3815 20983 3849
rect 21151 3815 21167 3849
rect 21339 3815 21355 3849
rect 21523 3815 21539 3849
rect 21711 3815 21727 3849
rect 21895 3815 21911 3849
rect 22083 3815 22099 3849
rect 22267 3815 22283 3849
rect 22455 3815 22471 3849
rect 22639 3815 22655 3849
rect 22827 3815 22843 3849
rect 23011 3815 23027 3849
rect 23199 3815 23215 3849
rect 23383 3815 23399 3849
rect 23571 3815 23587 3849
rect 23755 3815 23771 3849
rect 23943 3815 23959 3849
rect 24127 3815 24143 3849
rect 24315 3815 24331 3849
rect 24499 3815 24515 3849
rect 24687 3815 24703 3849
rect 24871 3815 24887 3849
rect 25059 3815 25075 3849
rect 25243 3815 25259 3849
rect 25431 3815 25447 3849
rect 25615 3815 25631 3849
rect 25803 3815 25819 3849
rect 25987 3815 26003 3849
rect 26175 3815 26191 3849
rect 26359 3815 26375 3849
rect 26547 3815 26563 3849
rect 26731 3815 26747 3849
rect 26919 3815 26935 3849
rect 27103 3815 27119 3849
rect 27291 3815 27307 3849
rect 27475 3815 27491 3849
rect 27663 3815 27679 3849
rect 27847 3815 27863 3849
rect 28035 3815 28051 3849
rect 28219 3815 28235 3849
rect 28407 3815 28423 3849
rect 28591 3815 28607 3849
rect 28779 3815 28795 3849
rect 28963 3815 28979 3849
rect 20223 3707 20239 3741
rect 20407 3707 20423 3741
rect 20595 3707 20611 3741
rect 20779 3707 20795 3741
rect 20967 3707 20983 3741
rect 21151 3707 21167 3741
rect 21339 3707 21355 3741
rect 21523 3707 21539 3741
rect 21711 3707 21727 3741
rect 21895 3707 21911 3741
rect 22083 3707 22099 3741
rect 22267 3707 22283 3741
rect 22455 3707 22471 3741
rect 22639 3707 22655 3741
rect 22827 3707 22843 3741
rect 23011 3707 23027 3741
rect 23199 3707 23215 3741
rect 23383 3707 23399 3741
rect 23571 3707 23587 3741
rect 23755 3707 23771 3741
rect 23943 3707 23959 3741
rect 24127 3707 24143 3741
rect 24315 3707 24331 3741
rect 24499 3707 24515 3741
rect 24687 3707 24703 3741
rect 24871 3707 24887 3741
rect 25059 3707 25075 3741
rect 25243 3707 25259 3741
rect 25431 3707 25447 3741
rect 25615 3707 25631 3741
rect 25803 3707 25819 3741
rect 25987 3707 26003 3741
rect 26175 3707 26191 3741
rect 26359 3707 26375 3741
rect 26547 3707 26563 3741
rect 26731 3707 26747 3741
rect 26919 3707 26935 3741
rect 27103 3707 27119 3741
rect 27291 3707 27307 3741
rect 27475 3707 27491 3741
rect 27663 3707 27679 3741
rect 27847 3707 27863 3741
rect 28035 3707 28051 3741
rect 28219 3707 28235 3741
rect 28407 3707 28423 3741
rect 28591 3707 28607 3741
rect 28779 3707 28795 3741
rect 28963 3707 28979 3741
rect 20177 3657 20211 3673
rect 20177 3465 20211 3481
rect 20435 3657 20469 3673
rect 20435 3465 20469 3481
rect 20549 3657 20583 3673
rect 20549 3465 20583 3481
rect 20807 3657 20841 3673
rect 20807 3465 20841 3481
rect 20921 3657 20955 3673
rect 20921 3465 20955 3481
rect 21179 3657 21213 3673
rect 21179 3465 21213 3481
rect 21293 3657 21327 3673
rect 21293 3465 21327 3481
rect 21551 3657 21585 3673
rect 21551 3465 21585 3481
rect 21665 3657 21699 3673
rect 21665 3465 21699 3481
rect 21923 3657 21957 3673
rect 21923 3465 21957 3481
rect 22037 3657 22071 3673
rect 22037 3465 22071 3481
rect 22295 3657 22329 3673
rect 22295 3465 22329 3481
rect 22409 3657 22443 3673
rect 22409 3465 22443 3481
rect 22667 3657 22701 3673
rect 22667 3465 22701 3481
rect 22781 3657 22815 3673
rect 22781 3465 22815 3481
rect 23039 3657 23073 3673
rect 23039 3465 23073 3481
rect 23153 3657 23187 3673
rect 23153 3465 23187 3481
rect 23411 3657 23445 3673
rect 23411 3465 23445 3481
rect 23525 3657 23559 3673
rect 23525 3465 23559 3481
rect 23783 3657 23817 3673
rect 23783 3465 23817 3481
rect 23897 3657 23931 3673
rect 23897 3465 23931 3481
rect 24155 3657 24189 3673
rect 24155 3465 24189 3481
rect 24269 3657 24303 3673
rect 24269 3465 24303 3481
rect 24527 3657 24561 3673
rect 24527 3465 24561 3481
rect 24641 3657 24675 3673
rect 24641 3465 24675 3481
rect 24899 3657 24933 3673
rect 24899 3465 24933 3481
rect 25013 3657 25047 3673
rect 25013 3465 25047 3481
rect 25271 3657 25305 3673
rect 25271 3465 25305 3481
rect 25385 3657 25419 3673
rect 25385 3465 25419 3481
rect 25643 3657 25677 3673
rect 25643 3465 25677 3481
rect 25757 3657 25791 3673
rect 25757 3465 25791 3481
rect 26015 3657 26049 3673
rect 26015 3465 26049 3481
rect 26129 3657 26163 3673
rect 26129 3465 26163 3481
rect 26387 3657 26421 3673
rect 26387 3465 26421 3481
rect 26501 3657 26535 3673
rect 26501 3465 26535 3481
rect 26759 3657 26793 3673
rect 26759 3465 26793 3481
rect 26873 3657 26907 3673
rect 26873 3465 26907 3481
rect 27131 3657 27165 3673
rect 27131 3465 27165 3481
rect 27245 3657 27279 3673
rect 27245 3465 27279 3481
rect 27503 3657 27537 3673
rect 27503 3465 27537 3481
rect 27617 3657 27651 3673
rect 27617 3465 27651 3481
rect 27875 3657 27909 3673
rect 27875 3465 27909 3481
rect 27989 3657 28023 3673
rect 27989 3465 28023 3481
rect 28247 3657 28281 3673
rect 28247 3465 28281 3481
rect 28361 3657 28395 3673
rect 28361 3465 28395 3481
rect 28619 3657 28653 3673
rect 28619 3465 28653 3481
rect 28733 3657 28767 3673
rect 28733 3465 28767 3481
rect 28991 3657 29025 3673
rect 28991 3465 29025 3481
rect 20223 3397 20239 3431
rect 20407 3397 20423 3431
rect 20595 3397 20611 3431
rect 20779 3397 20795 3431
rect 20967 3397 20983 3431
rect 21151 3397 21167 3431
rect 21339 3397 21355 3431
rect 21523 3397 21539 3431
rect 21711 3397 21727 3431
rect 21895 3397 21911 3431
rect 22083 3397 22099 3431
rect 22267 3397 22283 3431
rect 22455 3397 22471 3431
rect 22639 3397 22655 3431
rect 22827 3397 22843 3431
rect 23011 3397 23027 3431
rect 23199 3397 23215 3431
rect 23383 3397 23399 3431
rect 23571 3397 23587 3431
rect 23755 3397 23771 3431
rect 23943 3397 23959 3431
rect 24127 3397 24143 3431
rect 24315 3397 24331 3431
rect 24499 3397 24515 3431
rect 24687 3397 24703 3431
rect 24871 3397 24887 3431
rect 25059 3397 25075 3431
rect 25243 3397 25259 3431
rect 25431 3397 25447 3431
rect 25615 3397 25631 3431
rect 25803 3397 25819 3431
rect 25987 3397 26003 3431
rect 26175 3397 26191 3431
rect 26359 3397 26375 3431
rect 26547 3397 26563 3431
rect 26731 3397 26747 3431
rect 26919 3397 26935 3431
rect 27103 3397 27119 3431
rect 27291 3397 27307 3431
rect 27475 3397 27491 3431
rect 27663 3397 27679 3431
rect 27847 3397 27863 3431
rect 28035 3397 28051 3431
rect 28219 3397 28235 3431
rect 28407 3397 28423 3431
rect 28591 3397 28607 3431
rect 28779 3397 28795 3431
rect 28963 3397 28979 3431
rect 20223 3289 20239 3323
rect 20407 3289 20423 3323
rect 20595 3289 20611 3323
rect 20779 3289 20795 3323
rect 20967 3289 20983 3323
rect 21151 3289 21167 3323
rect 21339 3289 21355 3323
rect 21523 3289 21539 3323
rect 21711 3289 21727 3323
rect 21895 3289 21911 3323
rect 22083 3289 22099 3323
rect 22267 3289 22283 3323
rect 22455 3289 22471 3323
rect 22639 3289 22655 3323
rect 22827 3289 22843 3323
rect 23011 3289 23027 3323
rect 23199 3289 23215 3323
rect 23383 3289 23399 3323
rect 23571 3289 23587 3323
rect 23755 3289 23771 3323
rect 23943 3289 23959 3323
rect 24127 3289 24143 3323
rect 24315 3289 24331 3323
rect 24499 3289 24515 3323
rect 24687 3289 24703 3323
rect 24871 3289 24887 3323
rect 25059 3289 25075 3323
rect 25243 3289 25259 3323
rect 25431 3289 25447 3323
rect 25615 3289 25631 3323
rect 25803 3289 25819 3323
rect 25987 3289 26003 3323
rect 26175 3289 26191 3323
rect 26359 3289 26375 3323
rect 26547 3289 26563 3323
rect 26731 3289 26747 3323
rect 26919 3289 26935 3323
rect 27103 3289 27119 3323
rect 27291 3289 27307 3323
rect 27475 3289 27491 3323
rect 27663 3289 27679 3323
rect 27847 3289 27863 3323
rect 28035 3289 28051 3323
rect 28219 3289 28235 3323
rect 28407 3289 28423 3323
rect 28591 3289 28607 3323
rect 28779 3289 28795 3323
rect 28963 3289 28979 3323
rect 20177 3239 20211 3255
rect 20177 3047 20211 3063
rect 20435 3239 20469 3255
rect 20435 3047 20469 3063
rect 20549 3239 20583 3255
rect 20549 3047 20583 3063
rect 20807 3239 20841 3255
rect 20807 3047 20841 3063
rect 20921 3239 20955 3255
rect 20921 3047 20955 3063
rect 21179 3239 21213 3255
rect 21179 3047 21213 3063
rect 21293 3239 21327 3255
rect 21293 3047 21327 3063
rect 21551 3239 21585 3255
rect 21551 3047 21585 3063
rect 21665 3239 21699 3255
rect 21665 3047 21699 3063
rect 21923 3239 21957 3255
rect 21923 3047 21957 3063
rect 22037 3239 22071 3255
rect 22037 3047 22071 3063
rect 22295 3239 22329 3255
rect 22295 3047 22329 3063
rect 22409 3239 22443 3255
rect 22409 3047 22443 3063
rect 22667 3239 22701 3255
rect 22667 3047 22701 3063
rect 22781 3239 22815 3255
rect 22781 3047 22815 3063
rect 23039 3239 23073 3255
rect 23039 3047 23073 3063
rect 23153 3239 23187 3255
rect 23153 3047 23187 3063
rect 23411 3239 23445 3255
rect 23411 3047 23445 3063
rect 23525 3239 23559 3255
rect 23525 3047 23559 3063
rect 23783 3239 23817 3255
rect 23783 3047 23817 3063
rect 23897 3239 23931 3255
rect 23897 3047 23931 3063
rect 24155 3239 24189 3255
rect 24155 3047 24189 3063
rect 24269 3239 24303 3255
rect 24269 3047 24303 3063
rect 24527 3239 24561 3255
rect 24527 3047 24561 3063
rect 24641 3239 24675 3255
rect 24641 3047 24675 3063
rect 24899 3239 24933 3255
rect 24899 3047 24933 3063
rect 25013 3239 25047 3255
rect 25013 3047 25047 3063
rect 25271 3239 25305 3255
rect 25271 3047 25305 3063
rect 25385 3239 25419 3255
rect 25385 3047 25419 3063
rect 25643 3239 25677 3255
rect 25643 3047 25677 3063
rect 25757 3239 25791 3255
rect 25757 3047 25791 3063
rect 26015 3239 26049 3255
rect 26015 3047 26049 3063
rect 26129 3239 26163 3255
rect 26129 3047 26163 3063
rect 26387 3239 26421 3255
rect 26387 3047 26421 3063
rect 26501 3239 26535 3255
rect 26501 3047 26535 3063
rect 26759 3239 26793 3255
rect 26759 3047 26793 3063
rect 26873 3239 26907 3255
rect 26873 3047 26907 3063
rect 27131 3239 27165 3255
rect 27131 3047 27165 3063
rect 27245 3239 27279 3255
rect 27245 3047 27279 3063
rect 27503 3239 27537 3255
rect 27503 3047 27537 3063
rect 27617 3239 27651 3255
rect 27617 3047 27651 3063
rect 27875 3239 27909 3255
rect 27875 3047 27909 3063
rect 27989 3239 28023 3255
rect 27989 3047 28023 3063
rect 28247 3239 28281 3255
rect 28247 3047 28281 3063
rect 28361 3239 28395 3255
rect 28361 3047 28395 3063
rect 28619 3239 28653 3255
rect 28619 3047 28653 3063
rect 28733 3239 28767 3255
rect 28733 3047 28767 3063
rect 28991 3239 29025 3255
rect 28991 3047 29025 3063
rect 20223 2979 20239 3013
rect 20407 2979 20423 3013
rect 20595 2979 20611 3013
rect 20779 2979 20795 3013
rect 20967 2979 20983 3013
rect 21151 2979 21167 3013
rect 21339 2979 21355 3013
rect 21523 2979 21539 3013
rect 21711 2979 21727 3013
rect 21895 2979 21911 3013
rect 22083 2979 22099 3013
rect 22267 2979 22283 3013
rect 22455 2979 22471 3013
rect 22639 2979 22655 3013
rect 22827 2979 22843 3013
rect 23011 2979 23027 3013
rect 23199 2979 23215 3013
rect 23383 2979 23399 3013
rect 23571 2979 23587 3013
rect 23755 2979 23771 3013
rect 23943 2979 23959 3013
rect 24127 2979 24143 3013
rect 24315 2979 24331 3013
rect 24499 2979 24515 3013
rect 24687 2979 24703 3013
rect 24871 2979 24887 3013
rect 25059 2979 25075 3013
rect 25243 2979 25259 3013
rect 25431 2979 25447 3013
rect 25615 2979 25631 3013
rect 25803 2979 25819 3013
rect 25987 2979 26003 3013
rect 26175 2979 26191 3013
rect 26359 2979 26375 3013
rect 26547 2979 26563 3013
rect 26731 2979 26747 3013
rect 26919 2979 26935 3013
rect 27103 2979 27119 3013
rect 27291 2979 27307 3013
rect 27475 2979 27491 3013
rect 27663 2979 27679 3013
rect 27847 2979 27863 3013
rect 28035 2979 28051 3013
rect 28219 2979 28235 3013
rect 28407 2979 28423 3013
rect 28591 2979 28607 3013
rect 28779 2979 28795 3013
rect 28963 2979 28979 3013
rect 20063 2911 20097 2973
rect 29105 2911 29139 2973
rect 20063 2877 20159 2911
rect 29043 2877 29139 2911
<< viali >>
rect 18986 11761 19056 11778
rect 19730 11761 19800 11778
rect 20474 11761 20544 11778
rect 21218 11761 21288 11778
rect 21962 11761 22032 11778
rect 22706 11761 22776 11778
rect 23450 11761 23520 11778
rect 24194 11761 24264 11778
rect 24566 11761 24636 11778
rect 25310 11761 25380 11778
rect 26054 11761 26124 11778
rect 26798 11761 26868 11778
rect 27542 11761 27612 11778
rect 28286 11761 28356 11778
rect 29030 11761 29100 11778
rect 29774 11761 29844 11778
rect 30464 11761 30534 11778
rect 18986 11727 19056 11761
rect 19730 11727 19800 11761
rect 20474 11727 20544 11761
rect 21218 11727 21288 11761
rect 21962 11727 22032 11761
rect 22706 11727 22776 11761
rect 23450 11727 23520 11761
rect 24194 11727 24264 11761
rect 24566 11727 24636 11761
rect 25310 11727 25380 11761
rect 26054 11727 26124 11761
rect 26798 11727 26868 11761
rect 27542 11727 27612 11761
rect 28286 11727 28356 11761
rect 29030 11727 29100 11761
rect 29774 11727 29844 11761
rect 30464 11727 30531 11761
rect 30531 11727 30534 11761
rect 18986 11708 19056 11727
rect 19730 11708 19800 11727
rect 20474 11708 20544 11727
rect 21218 11708 21288 11727
rect 21962 11708 22032 11727
rect 22706 11708 22776 11727
rect 23450 11708 23520 11727
rect 24194 11708 24264 11727
rect 24566 11708 24636 11727
rect 25310 11708 25380 11727
rect 26054 11708 26124 11727
rect 26798 11708 26868 11727
rect 27542 11708 27612 11727
rect 28286 11708 28356 11727
rect 29030 11708 29100 11727
rect 29774 11708 29844 11727
rect 30464 11708 30534 11727
rect 18751 11625 18919 11659
rect 19123 11625 19291 11659
rect 19495 11625 19663 11659
rect 19867 11625 20035 11659
rect 20239 11625 20407 11659
rect 20611 11625 20779 11659
rect 20983 11625 21151 11659
rect 21355 11625 21523 11659
rect 21727 11625 21895 11659
rect 22099 11625 22267 11659
rect 22471 11625 22639 11659
rect 22843 11625 23011 11659
rect 23215 11625 23383 11659
rect 23587 11625 23755 11659
rect 23959 11625 24127 11659
rect 24331 11625 24499 11659
rect 24703 11625 24871 11659
rect 25075 11625 25243 11659
rect 25447 11625 25615 11659
rect 25819 11625 25987 11659
rect 26191 11625 26359 11659
rect 26563 11625 26731 11659
rect 26935 11625 27103 11659
rect 27307 11625 27475 11659
rect 27679 11625 27847 11659
rect 28051 11625 28219 11659
rect 28423 11625 28591 11659
rect 28795 11625 28963 11659
rect 29167 11625 29335 11659
rect 29539 11625 29707 11659
rect 29911 11625 30079 11659
rect 30283 11625 30451 11659
rect 18689 11190 18723 11566
rect 18947 11190 18981 11566
rect 19061 11190 19095 11566
rect 19319 11190 19353 11566
rect 19433 11190 19467 11566
rect 19691 11190 19725 11566
rect 19805 11190 19839 11566
rect 20063 11190 20097 11566
rect 20177 11190 20211 11566
rect 20435 11190 20469 11566
rect 20549 11190 20583 11566
rect 20807 11190 20841 11566
rect 20921 11190 20955 11566
rect 21179 11190 21213 11566
rect 21293 11190 21327 11566
rect 21551 11190 21585 11566
rect 21665 11190 21699 11566
rect 21923 11190 21957 11566
rect 22037 11190 22071 11566
rect 22295 11190 22329 11566
rect 22409 11190 22443 11566
rect 22667 11190 22701 11566
rect 22781 11190 22815 11566
rect 23039 11190 23073 11566
rect 23153 11190 23187 11566
rect 23411 11190 23445 11566
rect 23525 11190 23559 11566
rect 23783 11190 23817 11566
rect 23897 11190 23931 11566
rect 24155 11190 24189 11566
rect 24269 11190 24303 11566
rect 24527 11190 24561 11566
rect 24641 11190 24675 11566
rect 24899 11190 24933 11566
rect 25013 11190 25047 11566
rect 25271 11190 25305 11566
rect 25385 11190 25419 11566
rect 25643 11190 25677 11566
rect 25757 11190 25791 11566
rect 26015 11190 26049 11566
rect 26129 11190 26163 11566
rect 26387 11190 26421 11566
rect 26501 11190 26535 11566
rect 26759 11190 26793 11566
rect 26873 11190 26907 11566
rect 27131 11190 27165 11566
rect 27245 11190 27279 11566
rect 27503 11190 27537 11566
rect 27617 11190 27651 11566
rect 27875 11190 27909 11566
rect 27989 11190 28023 11566
rect 28247 11190 28281 11566
rect 28361 11190 28395 11566
rect 28619 11190 28653 11566
rect 28733 11190 28767 11566
rect 28991 11190 29025 11566
rect 29105 11190 29139 11566
rect 29363 11190 29397 11566
rect 29477 11190 29511 11566
rect 29735 11190 29769 11566
rect 29849 11190 29883 11566
rect 30107 11190 30141 11566
rect 30221 11190 30255 11566
rect 30479 11190 30513 11566
rect 18751 11097 18919 11131
rect 19123 11097 19291 11131
rect 19495 11097 19663 11131
rect 19867 11097 20035 11131
rect 20239 11097 20407 11131
rect 20611 11097 20779 11131
rect 20983 11097 21151 11131
rect 21355 11097 21523 11131
rect 21727 11097 21895 11131
rect 22099 11097 22267 11131
rect 22471 11097 22639 11131
rect 22843 11097 23011 11131
rect 23215 11097 23383 11131
rect 23587 11097 23755 11131
rect 23959 11097 24127 11131
rect 24331 11097 24499 11131
rect 24703 11097 24871 11131
rect 25075 11097 25243 11131
rect 25447 11097 25615 11131
rect 25819 11097 25987 11131
rect 26191 11097 26359 11131
rect 26563 11097 26731 11131
rect 26935 11097 27103 11131
rect 27307 11097 27475 11131
rect 27679 11097 27847 11131
rect 28051 11097 28219 11131
rect 28423 11097 28591 11131
rect 28795 11097 28963 11131
rect 29167 11097 29335 11131
rect 29539 11097 29707 11131
rect 29911 11097 30079 11131
rect 30283 11097 30451 11131
rect 18751 10989 18919 11023
rect 19123 10989 19291 11023
rect 19495 10989 19663 11023
rect 19867 10989 20035 11023
rect 20239 10989 20407 11023
rect 20611 10989 20779 11023
rect 20983 10989 21151 11023
rect 21355 10989 21523 11023
rect 21727 10989 21895 11023
rect 22099 10989 22267 11023
rect 22471 10989 22639 11023
rect 22843 10989 23011 11023
rect 23215 10989 23383 11023
rect 23587 10989 23755 11023
rect 23959 10989 24127 11023
rect 24331 10989 24499 11023
rect 24703 10989 24871 11023
rect 25075 10989 25243 11023
rect 25447 10989 25615 11023
rect 25819 10989 25987 11023
rect 26191 10989 26359 11023
rect 26563 10989 26731 11023
rect 26935 10989 27103 11023
rect 27307 10989 27475 11023
rect 27679 10989 27847 11023
rect 28051 10989 28219 11023
rect 28423 10989 28591 11023
rect 28795 10989 28963 11023
rect 29167 10989 29335 11023
rect 29539 10989 29707 11023
rect 29911 10989 30079 11023
rect 30283 10989 30451 11023
rect 18689 10554 18723 10930
rect 18947 10554 18981 10930
rect 19061 10554 19095 10930
rect 19319 10554 19353 10930
rect 19433 10554 19467 10930
rect 19691 10554 19725 10930
rect 19805 10554 19839 10930
rect 20063 10554 20097 10930
rect 20177 10554 20211 10930
rect 20435 10554 20469 10930
rect 20549 10554 20583 10930
rect 20807 10554 20841 10930
rect 20921 10554 20955 10930
rect 21179 10554 21213 10930
rect 21293 10554 21327 10930
rect 21551 10554 21585 10930
rect 21665 10554 21699 10930
rect 21923 10554 21957 10930
rect 22037 10554 22071 10930
rect 22295 10554 22329 10930
rect 22409 10554 22443 10930
rect 22667 10554 22701 10930
rect 22781 10554 22815 10930
rect 23039 10554 23073 10930
rect 23153 10554 23187 10930
rect 23411 10554 23445 10930
rect 23525 10554 23559 10930
rect 23783 10554 23817 10930
rect 23897 10554 23931 10930
rect 24155 10554 24189 10930
rect 24269 10554 24303 10930
rect 24527 10554 24561 10930
rect 24641 10554 24675 10930
rect 24899 10554 24933 10930
rect 25013 10554 25047 10930
rect 25271 10554 25305 10930
rect 25385 10554 25419 10930
rect 25643 10554 25677 10930
rect 25757 10554 25791 10930
rect 26015 10554 26049 10930
rect 26129 10554 26163 10930
rect 26387 10554 26421 10930
rect 26501 10554 26535 10930
rect 26759 10554 26793 10930
rect 26873 10554 26907 10930
rect 27131 10554 27165 10930
rect 27245 10554 27279 10930
rect 27503 10554 27537 10930
rect 27617 10554 27651 10930
rect 27875 10554 27909 10930
rect 27989 10554 28023 10930
rect 28247 10554 28281 10930
rect 28361 10554 28395 10930
rect 28619 10554 28653 10930
rect 28733 10554 28767 10930
rect 28991 10554 29025 10930
rect 29105 10554 29139 10930
rect 29363 10554 29397 10930
rect 29477 10554 29511 10930
rect 29735 10554 29769 10930
rect 29849 10554 29883 10930
rect 30107 10554 30141 10930
rect 30221 10554 30255 10930
rect 30479 10554 30513 10930
rect 18751 10461 18919 10495
rect 19123 10461 19291 10495
rect 19495 10461 19663 10495
rect 19867 10461 20035 10495
rect 20239 10461 20407 10495
rect 20611 10461 20779 10495
rect 20983 10461 21151 10495
rect 21355 10461 21523 10495
rect 21727 10461 21895 10495
rect 22099 10461 22267 10495
rect 22471 10461 22639 10495
rect 22843 10461 23011 10495
rect 23215 10461 23383 10495
rect 23587 10461 23755 10495
rect 23959 10461 24127 10495
rect 24331 10461 24499 10495
rect 24703 10461 24871 10495
rect 25075 10461 25243 10495
rect 25447 10461 25615 10495
rect 25819 10461 25987 10495
rect 26191 10461 26359 10495
rect 26563 10461 26731 10495
rect 26935 10461 27103 10495
rect 27307 10461 27475 10495
rect 27679 10461 27847 10495
rect 28051 10461 28219 10495
rect 28423 10461 28591 10495
rect 28795 10461 28963 10495
rect 29167 10461 29335 10495
rect 29539 10461 29707 10495
rect 29911 10461 30079 10495
rect 30283 10461 30451 10495
rect 18751 10353 18919 10387
rect 19123 10353 19291 10387
rect 19495 10353 19663 10387
rect 19867 10353 20035 10387
rect 20239 10353 20407 10387
rect 20611 10353 20779 10387
rect 20983 10353 21151 10387
rect 21355 10353 21523 10387
rect 21727 10353 21895 10387
rect 22099 10353 22267 10387
rect 22471 10353 22639 10387
rect 22843 10353 23011 10387
rect 23215 10353 23383 10387
rect 23587 10353 23755 10387
rect 23959 10353 24127 10387
rect 24331 10353 24499 10387
rect 24703 10353 24871 10387
rect 25075 10353 25243 10387
rect 25447 10353 25615 10387
rect 25819 10353 25987 10387
rect 26191 10353 26359 10387
rect 26563 10353 26731 10387
rect 26935 10353 27103 10387
rect 27307 10353 27475 10387
rect 27679 10353 27847 10387
rect 28051 10353 28219 10387
rect 28423 10353 28591 10387
rect 28795 10353 28963 10387
rect 29167 10353 29335 10387
rect 29539 10353 29707 10387
rect 29911 10353 30079 10387
rect 30283 10353 30451 10387
rect 18689 9918 18723 10294
rect 18947 9918 18981 10294
rect 19061 9918 19095 10294
rect 19319 9918 19353 10294
rect 19433 9918 19467 10294
rect 19691 9918 19725 10294
rect 19805 9918 19839 10294
rect 20063 9918 20097 10294
rect 20177 9918 20211 10294
rect 20435 9918 20469 10294
rect 20549 9918 20583 10294
rect 20807 9918 20841 10294
rect 20921 9918 20955 10294
rect 21179 9918 21213 10294
rect 21293 9918 21327 10294
rect 21551 9918 21585 10294
rect 21665 9918 21699 10294
rect 21923 9918 21957 10294
rect 22037 9918 22071 10294
rect 22295 9918 22329 10294
rect 22409 9918 22443 10294
rect 22667 9918 22701 10294
rect 22781 9918 22815 10294
rect 23039 9918 23073 10294
rect 23153 9918 23187 10294
rect 23411 9918 23445 10294
rect 23525 9918 23559 10294
rect 23783 9918 23817 10294
rect 23897 9918 23931 10294
rect 24155 9918 24189 10294
rect 24269 9918 24303 10294
rect 24527 9918 24561 10294
rect 24641 9918 24675 10294
rect 24899 9918 24933 10294
rect 25013 9918 25047 10294
rect 25271 9918 25305 10294
rect 25385 9918 25419 10294
rect 25643 9918 25677 10294
rect 25757 9918 25791 10294
rect 26015 9918 26049 10294
rect 26129 9918 26163 10294
rect 26387 9918 26421 10294
rect 26501 9918 26535 10294
rect 26759 9918 26793 10294
rect 26873 9918 26907 10294
rect 27131 9918 27165 10294
rect 27245 9918 27279 10294
rect 27503 9918 27537 10294
rect 27617 9918 27651 10294
rect 27875 9918 27909 10294
rect 27989 9918 28023 10294
rect 28247 9918 28281 10294
rect 28361 9918 28395 10294
rect 28619 9918 28653 10294
rect 28733 9918 28767 10294
rect 28991 9918 29025 10294
rect 29105 9918 29139 10294
rect 29363 9918 29397 10294
rect 29477 9918 29511 10294
rect 29735 9918 29769 10294
rect 29849 9918 29883 10294
rect 30107 9918 30141 10294
rect 30221 9918 30255 10294
rect 30479 9918 30513 10294
rect 18751 9825 18919 9859
rect 19123 9825 19291 9859
rect 19495 9825 19663 9859
rect 19867 9825 20035 9859
rect 20239 9825 20407 9859
rect 20611 9825 20779 9859
rect 20983 9825 21151 9859
rect 21355 9825 21523 9859
rect 21727 9825 21895 9859
rect 22099 9825 22267 9859
rect 22471 9825 22639 9859
rect 22843 9825 23011 9859
rect 23215 9825 23383 9859
rect 23587 9825 23755 9859
rect 23959 9825 24127 9859
rect 24331 9825 24499 9859
rect 24703 9825 24871 9859
rect 25075 9825 25243 9859
rect 25447 9825 25615 9859
rect 25819 9825 25987 9859
rect 26191 9825 26359 9859
rect 26563 9825 26731 9859
rect 26935 9825 27103 9859
rect 27307 9825 27475 9859
rect 27679 9825 27847 9859
rect 28051 9825 28219 9859
rect 28423 9825 28591 9859
rect 28795 9825 28963 9859
rect 29167 9825 29335 9859
rect 29539 9825 29707 9859
rect 29911 9825 30079 9859
rect 30283 9825 30451 9859
rect 20148 9373 20218 9390
rect 20520 9373 20590 9390
rect 20892 9373 20962 9390
rect 21264 9373 21334 9390
rect 21636 9373 21706 9390
rect 22008 9373 22078 9390
rect 22380 9373 22450 9390
rect 22752 9373 22822 9390
rect 23014 9373 23084 9390
rect 20148 9339 20159 9373
rect 20159 9339 20218 9373
rect 20520 9339 20590 9373
rect 20892 9339 20962 9373
rect 21264 9339 21334 9373
rect 21636 9339 21706 9373
rect 22008 9339 22078 9373
rect 22380 9339 22450 9373
rect 22752 9339 22822 9373
rect 23014 9339 23084 9373
rect 20148 9320 20218 9339
rect 20520 9320 20590 9339
rect 20892 9320 20962 9339
rect 21264 9320 21334 9339
rect 21636 9320 21706 9339
rect 22008 9320 22078 9339
rect 22380 9320 22450 9339
rect 22752 9320 22822 9339
rect 23014 9320 23084 9339
rect 20239 9237 20407 9271
rect 20611 9237 20779 9271
rect 20983 9237 21151 9271
rect 21355 9237 21523 9271
rect 21727 9237 21895 9271
rect 22099 9237 22267 9271
rect 22471 9237 22639 9271
rect 22843 9237 23011 9271
rect 20177 8402 20211 9178
rect 20435 8402 20469 9178
rect 20549 8402 20583 9178
rect 20807 8402 20841 9178
rect 20921 8402 20955 9178
rect 21179 8402 21213 9178
rect 21293 8402 21327 9178
rect 21551 8402 21585 9178
rect 21665 8402 21699 9178
rect 21923 8402 21957 9178
rect 22037 8402 22071 9178
rect 22295 8402 22329 9178
rect 22409 8402 22443 9178
rect 22667 8402 22701 9178
rect 22781 8402 22815 9178
rect 23039 8402 23073 9178
rect 20239 8309 20407 8343
rect 20611 8309 20779 8343
rect 20983 8309 21151 8343
rect 21355 8309 21523 8343
rect 21727 8309 21895 8343
rect 22099 8309 22267 8343
rect 22471 8309 22639 8343
rect 22843 8309 23011 8343
rect 20239 8201 20407 8235
rect 20611 8201 20779 8235
rect 20983 8201 21151 8235
rect 21355 8201 21523 8235
rect 21727 8201 21895 8235
rect 22099 8201 22267 8235
rect 22471 8201 22639 8235
rect 22843 8201 23011 8235
rect 20177 7366 20211 8142
rect 20435 7366 20469 8142
rect 20549 7366 20583 8142
rect 20807 7366 20841 8142
rect 20921 7366 20955 8142
rect 21179 7366 21213 8142
rect 21293 7366 21327 8142
rect 21551 7366 21585 8142
rect 21665 7366 21699 8142
rect 21923 7366 21957 8142
rect 22037 7366 22071 8142
rect 22295 7366 22329 8142
rect 22409 7366 22443 8142
rect 22667 7366 22701 8142
rect 22781 7366 22815 8142
rect 23039 7366 23073 8142
rect 20239 7273 20407 7307
rect 20611 7273 20779 7307
rect 20983 7273 21151 7307
rect 21355 7273 21523 7307
rect 21727 7273 21895 7307
rect 22099 7273 22267 7307
rect 22471 7273 22639 7307
rect 22843 7273 23011 7307
rect 20239 7165 20407 7199
rect 20611 7165 20779 7199
rect 20983 7165 21151 7199
rect 21355 7165 21523 7199
rect 21727 7165 21895 7199
rect 22099 7165 22267 7199
rect 22471 7165 22639 7199
rect 22843 7165 23011 7199
rect 20177 6330 20211 7106
rect 20435 6330 20469 7106
rect 20549 6330 20583 7106
rect 20807 6330 20841 7106
rect 20921 6330 20955 7106
rect 21179 6330 21213 7106
rect 21293 6330 21327 7106
rect 21551 6330 21585 7106
rect 21665 6330 21699 7106
rect 21923 6330 21957 7106
rect 22037 6330 22071 7106
rect 22295 6330 22329 7106
rect 22409 6330 22443 7106
rect 22667 6330 22701 7106
rect 22781 6330 22815 7106
rect 23039 6330 23073 7106
rect 20239 6237 20407 6271
rect 20611 6237 20779 6271
rect 20983 6237 21151 6271
rect 21355 6237 21523 6271
rect 21727 6237 21895 6271
rect 22099 6237 22267 6271
rect 22471 6237 22639 6271
rect 22843 6237 23011 6271
rect 20239 6129 20407 6163
rect 20611 6129 20779 6163
rect 20983 6129 21151 6163
rect 21355 6129 21523 6163
rect 21727 6129 21895 6163
rect 22099 6129 22267 6163
rect 22471 6129 22639 6163
rect 22843 6129 23011 6163
rect 20177 5294 20211 6070
rect 20435 5294 20469 6070
rect 20549 5294 20583 6070
rect 20807 5294 20841 6070
rect 20921 5294 20955 6070
rect 21179 5294 21213 6070
rect 21293 5294 21327 6070
rect 21551 5294 21585 6070
rect 21665 5294 21699 6070
rect 21923 5294 21957 6070
rect 22037 5294 22071 6070
rect 22295 5294 22329 6070
rect 22409 5294 22443 6070
rect 22667 5294 22701 6070
rect 22781 5294 22815 6070
rect 23039 5294 23073 6070
rect 20239 5201 20407 5235
rect 20611 5201 20779 5235
rect 20983 5201 21151 5235
rect 21355 5201 21523 5235
rect 21727 5201 21895 5235
rect 22099 5201 22267 5235
rect 22471 5201 22639 5235
rect 22843 5201 23011 5235
rect 23835 6914 23873 7311
rect 23970 6756 23985 6816
rect 23985 6756 24019 6816
rect 24019 6756 24034 6816
rect 23970 6356 23985 6416
rect 23985 6356 24019 6416
rect 24019 6356 24034 6416
rect 23835 5923 23873 6320
rect 23970 5956 23985 6016
rect 23985 5956 24019 6016
rect 24019 5956 24034 6016
rect 20239 4543 20407 4577
rect 20611 4543 20779 4577
rect 20983 4543 21151 4577
rect 21355 4543 21523 4577
rect 21727 4543 21895 4577
rect 22099 4543 22267 4577
rect 22471 4543 22639 4577
rect 22843 4543 23011 4577
rect 23215 4543 23383 4577
rect 23587 4543 23755 4577
rect 23959 4543 24127 4577
rect 24331 4543 24499 4577
rect 24703 4543 24871 4577
rect 25075 4543 25243 4577
rect 25447 4543 25615 4577
rect 25819 4543 25987 4577
rect 26191 4543 26359 4577
rect 26563 4543 26731 4577
rect 26935 4543 27103 4577
rect 27307 4543 27475 4577
rect 27679 4543 27847 4577
rect 28051 4543 28219 4577
rect 28423 4543 28591 4577
rect 28795 4543 28963 4577
rect 20177 4317 20211 4493
rect 20435 4317 20469 4493
rect 20549 4317 20583 4493
rect 20807 4317 20841 4493
rect 20921 4317 20955 4493
rect 21179 4317 21213 4493
rect 21293 4317 21327 4493
rect 21551 4317 21585 4493
rect 21665 4317 21699 4493
rect 21923 4317 21957 4493
rect 22037 4317 22071 4493
rect 22295 4317 22329 4493
rect 22409 4317 22443 4493
rect 22667 4317 22701 4493
rect 22781 4317 22815 4493
rect 23039 4317 23073 4493
rect 23153 4317 23187 4493
rect 23411 4317 23445 4493
rect 23525 4317 23559 4493
rect 23783 4317 23817 4493
rect 23897 4317 23931 4493
rect 24155 4317 24189 4493
rect 24269 4317 24303 4493
rect 24527 4317 24561 4493
rect 24641 4317 24675 4493
rect 24899 4317 24933 4493
rect 25013 4317 25047 4493
rect 25271 4317 25305 4493
rect 25385 4317 25419 4493
rect 25643 4317 25677 4493
rect 25757 4317 25791 4493
rect 26015 4317 26049 4493
rect 26129 4317 26163 4493
rect 26387 4317 26421 4493
rect 26501 4317 26535 4493
rect 26759 4317 26793 4493
rect 26873 4317 26907 4493
rect 27131 4317 27165 4493
rect 27245 4317 27279 4493
rect 27503 4317 27537 4493
rect 27617 4317 27651 4493
rect 27875 4317 27909 4493
rect 27989 4317 28023 4493
rect 28247 4317 28281 4493
rect 28361 4317 28395 4493
rect 28619 4317 28653 4493
rect 28733 4317 28767 4493
rect 28991 4317 29025 4493
rect 20239 4233 20407 4267
rect 20611 4233 20779 4267
rect 20983 4233 21151 4267
rect 21355 4233 21523 4267
rect 21727 4233 21895 4267
rect 22099 4233 22267 4267
rect 22471 4233 22639 4267
rect 22843 4233 23011 4267
rect 23215 4233 23383 4267
rect 23587 4233 23755 4267
rect 23959 4233 24127 4267
rect 24331 4233 24499 4267
rect 24703 4233 24871 4267
rect 25075 4233 25243 4267
rect 25447 4233 25615 4267
rect 25819 4233 25987 4267
rect 26191 4233 26359 4267
rect 26563 4233 26731 4267
rect 26935 4233 27103 4267
rect 27307 4233 27475 4267
rect 27679 4233 27847 4267
rect 28051 4233 28219 4267
rect 28423 4233 28591 4267
rect 28795 4233 28963 4267
rect 20239 4125 20407 4159
rect 20611 4125 20779 4159
rect 20983 4125 21151 4159
rect 21355 4125 21523 4159
rect 21727 4125 21895 4159
rect 22099 4125 22267 4159
rect 22471 4125 22639 4159
rect 22843 4125 23011 4159
rect 23215 4125 23383 4159
rect 23587 4125 23755 4159
rect 23959 4125 24127 4159
rect 24331 4125 24499 4159
rect 24703 4125 24871 4159
rect 25075 4125 25243 4159
rect 25447 4125 25615 4159
rect 25819 4125 25987 4159
rect 26191 4125 26359 4159
rect 26563 4125 26731 4159
rect 26935 4125 27103 4159
rect 27307 4125 27475 4159
rect 27679 4125 27847 4159
rect 28051 4125 28219 4159
rect 28423 4125 28591 4159
rect 28795 4125 28963 4159
rect 20177 3899 20211 4075
rect 20435 3899 20469 4075
rect 20549 3899 20583 4075
rect 20807 3899 20841 4075
rect 20921 3899 20955 4075
rect 21179 3899 21213 4075
rect 21293 3899 21327 4075
rect 21551 3899 21585 4075
rect 21665 3899 21699 4075
rect 21923 3899 21957 4075
rect 22037 3899 22071 4075
rect 22295 3899 22329 4075
rect 22409 3899 22443 4075
rect 22667 3899 22701 4075
rect 22781 3899 22815 4075
rect 23039 3899 23073 4075
rect 23153 3899 23187 4075
rect 23411 3899 23445 4075
rect 23525 3899 23559 4075
rect 23783 3899 23817 4075
rect 23897 3899 23931 4075
rect 24155 3899 24189 4075
rect 24269 3899 24303 4075
rect 24527 3899 24561 4075
rect 24641 3899 24675 4075
rect 24899 3899 24933 4075
rect 25013 3899 25047 4075
rect 25271 3899 25305 4075
rect 25385 3899 25419 4075
rect 25643 3899 25677 4075
rect 25757 3899 25791 4075
rect 26015 3899 26049 4075
rect 26129 3899 26163 4075
rect 26387 3899 26421 4075
rect 26501 3899 26535 4075
rect 26759 3899 26793 4075
rect 26873 3899 26907 4075
rect 27131 3899 27165 4075
rect 27245 3899 27279 4075
rect 27503 3899 27537 4075
rect 27617 3899 27651 4075
rect 27875 3899 27909 4075
rect 27989 3899 28023 4075
rect 28247 3899 28281 4075
rect 28361 3899 28395 4075
rect 28619 3899 28653 4075
rect 28733 3899 28767 4075
rect 28991 3899 29025 4075
rect 20239 3815 20407 3849
rect 20611 3815 20779 3849
rect 20983 3815 21151 3849
rect 21355 3815 21523 3849
rect 21727 3815 21895 3849
rect 22099 3815 22267 3849
rect 22471 3815 22639 3849
rect 22843 3815 23011 3849
rect 23215 3815 23383 3849
rect 23587 3815 23755 3849
rect 23959 3815 24127 3849
rect 24331 3815 24499 3849
rect 24703 3815 24871 3849
rect 25075 3815 25243 3849
rect 25447 3815 25615 3849
rect 25819 3815 25987 3849
rect 26191 3815 26359 3849
rect 26563 3815 26731 3849
rect 26935 3815 27103 3849
rect 27307 3815 27475 3849
rect 27679 3815 27847 3849
rect 28051 3815 28219 3849
rect 28423 3815 28591 3849
rect 28795 3815 28963 3849
rect 20239 3707 20407 3741
rect 20611 3707 20779 3741
rect 20983 3707 21151 3741
rect 21355 3707 21523 3741
rect 21727 3707 21895 3741
rect 22099 3707 22267 3741
rect 22471 3707 22639 3741
rect 22843 3707 23011 3741
rect 23215 3707 23383 3741
rect 23587 3707 23755 3741
rect 23959 3707 24127 3741
rect 24331 3707 24499 3741
rect 24703 3707 24871 3741
rect 25075 3707 25243 3741
rect 25447 3707 25615 3741
rect 25819 3707 25987 3741
rect 26191 3707 26359 3741
rect 26563 3707 26731 3741
rect 26935 3707 27103 3741
rect 27307 3707 27475 3741
rect 27679 3707 27847 3741
rect 28051 3707 28219 3741
rect 28423 3707 28591 3741
rect 28795 3707 28963 3741
rect 20177 3481 20211 3657
rect 20435 3481 20469 3657
rect 20549 3481 20583 3657
rect 20807 3481 20841 3657
rect 20921 3481 20955 3657
rect 21179 3481 21213 3657
rect 21293 3481 21327 3657
rect 21551 3481 21585 3657
rect 21665 3481 21699 3657
rect 21923 3481 21957 3657
rect 22037 3481 22071 3657
rect 22295 3481 22329 3657
rect 22409 3481 22443 3657
rect 22667 3481 22701 3657
rect 22781 3481 22815 3657
rect 23039 3481 23073 3657
rect 23153 3481 23187 3657
rect 23411 3481 23445 3657
rect 23525 3481 23559 3657
rect 23783 3481 23817 3657
rect 23897 3481 23931 3657
rect 24155 3481 24189 3657
rect 24269 3481 24303 3657
rect 24527 3481 24561 3657
rect 24641 3481 24675 3657
rect 24899 3481 24933 3657
rect 25013 3481 25047 3657
rect 25271 3481 25305 3657
rect 25385 3481 25419 3657
rect 25643 3481 25677 3657
rect 25757 3481 25791 3657
rect 26015 3481 26049 3657
rect 26129 3481 26163 3657
rect 26387 3481 26421 3657
rect 26501 3481 26535 3657
rect 26759 3481 26793 3657
rect 26873 3481 26907 3657
rect 27131 3481 27165 3657
rect 27245 3481 27279 3657
rect 27503 3481 27537 3657
rect 27617 3481 27651 3657
rect 27875 3481 27909 3657
rect 27989 3481 28023 3657
rect 28247 3481 28281 3657
rect 28361 3481 28395 3657
rect 28619 3481 28653 3657
rect 28733 3481 28767 3657
rect 28991 3481 29025 3657
rect 20239 3397 20407 3431
rect 20611 3397 20779 3431
rect 20983 3397 21151 3431
rect 21355 3397 21523 3431
rect 21727 3397 21895 3431
rect 22099 3397 22267 3431
rect 22471 3397 22639 3431
rect 22843 3397 23011 3431
rect 23215 3397 23383 3431
rect 23587 3397 23755 3431
rect 23959 3397 24127 3431
rect 24331 3397 24499 3431
rect 24703 3397 24871 3431
rect 25075 3397 25243 3431
rect 25447 3397 25615 3431
rect 25819 3397 25987 3431
rect 26191 3397 26359 3431
rect 26563 3397 26731 3431
rect 26935 3397 27103 3431
rect 27307 3397 27475 3431
rect 27679 3397 27847 3431
rect 28051 3397 28219 3431
rect 28423 3397 28591 3431
rect 28795 3397 28963 3431
rect 20239 3289 20407 3323
rect 20611 3289 20779 3323
rect 20983 3289 21151 3323
rect 21355 3289 21523 3323
rect 21727 3289 21895 3323
rect 22099 3289 22267 3323
rect 22471 3289 22639 3323
rect 22843 3289 23011 3323
rect 23215 3289 23383 3323
rect 23587 3289 23755 3323
rect 23959 3289 24127 3323
rect 24331 3289 24499 3323
rect 24703 3289 24871 3323
rect 25075 3289 25243 3323
rect 25447 3289 25615 3323
rect 25819 3289 25987 3323
rect 26191 3289 26359 3323
rect 26563 3289 26731 3323
rect 26935 3289 27103 3323
rect 27307 3289 27475 3323
rect 27679 3289 27847 3323
rect 28051 3289 28219 3323
rect 28423 3289 28591 3323
rect 28795 3289 28963 3323
rect 20177 3063 20211 3239
rect 20435 3063 20469 3239
rect 20549 3063 20583 3239
rect 20807 3063 20841 3239
rect 20921 3063 20955 3239
rect 21179 3063 21213 3239
rect 21293 3063 21327 3239
rect 21551 3063 21585 3239
rect 21665 3063 21699 3239
rect 21923 3063 21957 3239
rect 22037 3063 22071 3239
rect 22295 3063 22329 3239
rect 22409 3063 22443 3239
rect 22667 3063 22701 3239
rect 22781 3063 22815 3239
rect 23039 3063 23073 3239
rect 23153 3063 23187 3239
rect 23411 3063 23445 3239
rect 23525 3063 23559 3239
rect 23783 3063 23817 3239
rect 23897 3063 23931 3239
rect 24155 3063 24189 3239
rect 24269 3063 24303 3239
rect 24527 3063 24561 3239
rect 24641 3063 24675 3239
rect 24899 3063 24933 3239
rect 25013 3063 25047 3239
rect 25271 3063 25305 3239
rect 25385 3063 25419 3239
rect 25643 3063 25677 3239
rect 25757 3063 25791 3239
rect 26015 3063 26049 3239
rect 26129 3063 26163 3239
rect 26387 3063 26421 3239
rect 26501 3063 26535 3239
rect 26759 3063 26793 3239
rect 26873 3063 26907 3239
rect 27131 3063 27165 3239
rect 27245 3063 27279 3239
rect 27503 3063 27537 3239
rect 27617 3063 27651 3239
rect 27875 3063 27909 3239
rect 27989 3063 28023 3239
rect 28247 3063 28281 3239
rect 28361 3063 28395 3239
rect 28619 3063 28653 3239
rect 28733 3063 28767 3239
rect 28991 3063 29025 3239
rect 20239 2979 20407 3013
rect 20611 2979 20779 3013
rect 20983 2979 21151 3013
rect 21355 2979 21523 3013
rect 21727 2979 21895 3013
rect 22099 2979 22267 3013
rect 22471 2979 22639 3013
rect 22843 2979 23011 3013
rect 23215 2979 23383 3013
rect 23587 2979 23755 3013
rect 23959 2979 24127 3013
rect 24331 2979 24499 3013
rect 24703 2979 24871 3013
rect 25075 2979 25243 3013
rect 25447 2979 25615 3013
rect 25819 2979 25987 3013
rect 26191 2979 26359 3013
rect 26563 2979 26731 3013
rect 26935 2979 27103 3013
rect 27307 2979 27475 3013
rect 27679 2979 27847 3013
rect 28051 2979 28219 3013
rect 28423 2979 28591 3013
rect 28795 2979 28963 3013
rect 20178 2911 20248 2922
rect 20846 2911 20916 2930
rect 21590 2911 21660 2930
rect 22334 2911 22404 2930
rect 23078 2911 23148 2930
rect 23822 2911 23892 2930
rect 24566 2911 24636 2930
rect 25310 2911 25380 2930
rect 26054 2911 26124 2930
rect 26798 2911 26868 2930
rect 27542 2911 27612 2930
rect 28286 2911 28356 2930
rect 28948 2911 29018 2926
rect 20178 2877 20248 2911
rect 20846 2877 20916 2911
rect 21590 2877 21660 2911
rect 22334 2877 22404 2911
rect 23078 2877 23148 2911
rect 23822 2877 23892 2911
rect 24566 2877 24636 2911
rect 25310 2877 25380 2911
rect 26054 2877 26124 2911
rect 26798 2877 26868 2911
rect 27542 2877 27612 2911
rect 28286 2877 28356 2911
rect 28948 2877 29018 2911
rect 20178 2852 20248 2877
rect 20846 2860 20916 2877
rect 21590 2860 21660 2877
rect 22334 2860 22404 2877
rect 23078 2860 23148 2877
rect 23822 2860 23892 2877
rect 24566 2860 24636 2877
rect 25310 2860 25380 2877
rect 26054 2860 26124 2877
rect 26798 2860 26868 2877
rect 27542 2860 27612 2877
rect 28286 2860 28356 2877
rect 28948 2856 29018 2877
<< metal1 >>
rect 18910 11860 18920 12060
rect 19120 11860 19130 12060
rect 19654 11860 19664 12060
rect 19864 11860 19874 12060
rect 20398 11860 20408 12060
rect 20608 11860 20618 12060
rect 21142 11860 21152 12060
rect 21352 11860 21362 12060
rect 21886 11860 21896 12060
rect 22096 11860 22106 12060
rect 22630 11860 22640 12060
rect 22840 11860 22850 12060
rect 23374 11860 23384 12060
rect 23584 11860 23594 12060
rect 24118 11860 24128 12060
rect 24328 11860 24338 12060
rect 24490 11860 24500 12060
rect 24700 11860 24710 12060
rect 25234 11860 25244 12060
rect 25444 11860 25454 12060
rect 25978 11860 25988 12060
rect 26188 11860 26198 12060
rect 26722 11860 26732 12060
rect 26932 11860 26942 12060
rect 27466 11860 27476 12060
rect 27676 11860 27686 12060
rect 28210 11860 28220 12060
rect 28420 11860 28430 12060
rect 28954 11860 28964 12060
rect 29164 11860 29174 12060
rect 29698 11860 29708 12060
rect 29908 11860 29918 12060
rect 30442 11860 30452 12060
rect 30652 11860 30662 12060
rect 18992 11784 19050 11860
rect 19736 11784 19794 11860
rect 20480 11784 20538 11860
rect 21224 11784 21282 11860
rect 21968 11784 22026 11860
rect 22712 11784 22770 11860
rect 23456 11784 23514 11860
rect 24180 11850 24258 11860
rect 24200 11784 24258 11850
rect 24610 11784 24662 11860
rect 25316 11784 25374 11860
rect 26060 11784 26118 11860
rect 26804 11784 26862 11860
rect 27548 11784 27606 11860
rect 28292 11784 28350 11860
rect 29036 11784 29094 11860
rect 29780 11784 29838 11860
rect 30506 11844 30582 11860
rect 30506 11784 30564 11844
rect 18974 11778 19068 11784
rect 18974 11708 18986 11778
rect 19056 11708 19068 11778
rect 18974 11702 19068 11708
rect 19718 11778 19812 11784
rect 19718 11708 19730 11778
rect 19800 11708 19812 11778
rect 19718 11702 19812 11708
rect 20462 11778 20556 11784
rect 20462 11708 20474 11778
rect 20544 11708 20556 11778
rect 20462 11702 20556 11708
rect 21206 11778 21300 11784
rect 21206 11708 21218 11778
rect 21288 11708 21300 11778
rect 21206 11702 21300 11708
rect 21950 11778 22044 11784
rect 21950 11708 21962 11778
rect 22032 11708 22044 11778
rect 21950 11702 22044 11708
rect 22694 11778 22788 11784
rect 22694 11708 22706 11778
rect 22776 11708 22788 11778
rect 22694 11702 22788 11708
rect 23438 11778 23532 11784
rect 23438 11708 23450 11778
rect 23520 11708 23532 11778
rect 23438 11702 23532 11708
rect 24182 11778 24276 11784
rect 24182 11708 24194 11778
rect 24264 11708 24276 11778
rect 24182 11702 24276 11708
rect 24554 11778 24662 11784
rect 24554 11708 24566 11778
rect 24636 11708 24662 11778
rect 24554 11702 24662 11708
rect 25298 11778 25392 11784
rect 25298 11708 25310 11778
rect 25380 11708 25392 11778
rect 25298 11702 25392 11708
rect 26042 11778 26136 11784
rect 26042 11708 26054 11778
rect 26124 11708 26136 11778
rect 26042 11702 26136 11708
rect 26786 11778 26880 11784
rect 26786 11708 26798 11778
rect 26868 11708 26880 11778
rect 26786 11702 26880 11708
rect 27530 11778 27624 11784
rect 27530 11708 27542 11778
rect 27612 11708 27624 11778
rect 27530 11702 27624 11708
rect 28274 11778 28368 11784
rect 28274 11708 28286 11778
rect 28356 11708 28368 11778
rect 28274 11702 28368 11708
rect 29018 11778 29112 11784
rect 29018 11708 29030 11778
rect 29100 11708 29112 11778
rect 29018 11702 29112 11708
rect 29762 11778 29856 11784
rect 29762 11708 29774 11778
rect 29844 11708 29856 11778
rect 29762 11702 29856 11708
rect 30452 11778 30564 11784
rect 30452 11708 30464 11778
rect 30534 11708 30564 11778
rect 30452 11702 30564 11708
rect 18682 11612 18750 11672
rect 18920 11665 18930 11672
rect 18920 11619 18931 11665
rect 18920 11612 18930 11619
rect 18682 11566 18730 11612
rect 18992 11578 19050 11702
rect 19112 11665 19122 11672
rect 19111 11619 19122 11665
rect 19292 11665 19302 11672
rect 19484 11665 19494 11672
rect 19112 11612 19122 11619
rect 19292 11619 19303 11665
rect 19483 11619 19494 11665
rect 19664 11665 19674 11672
rect 19292 11612 19302 11619
rect 19484 11612 19494 11619
rect 19664 11619 19675 11665
rect 19664 11612 19674 11619
rect 19736 11578 19794 11702
rect 19856 11665 19866 11672
rect 19855 11619 19866 11665
rect 19856 11612 19866 11619
rect 20036 11612 20238 11672
rect 20408 11665 20418 11672
rect 20408 11619 20419 11665
rect 20408 11612 20418 11619
rect 20108 11578 20166 11612
rect 20480 11578 20538 11702
rect 20600 11665 20610 11672
rect 20599 11619 20610 11665
rect 20780 11665 20790 11672
rect 20972 11665 20982 11672
rect 20600 11612 20610 11619
rect 20780 11619 20791 11665
rect 20971 11619 20982 11665
rect 21152 11665 21162 11672
rect 20780 11612 20790 11619
rect 20972 11612 20982 11619
rect 21152 11619 21163 11665
rect 21152 11612 21162 11619
rect 21224 11578 21282 11702
rect 21344 11665 21354 11672
rect 21343 11619 21354 11665
rect 21344 11612 21354 11619
rect 21524 11612 21726 11672
rect 21896 11665 21906 11672
rect 21896 11619 21907 11665
rect 21896 11612 21906 11619
rect 21596 11578 21654 11612
rect 21968 11578 22026 11702
rect 22088 11665 22098 11672
rect 22087 11619 22098 11665
rect 22268 11665 22278 11672
rect 22460 11665 22470 11672
rect 22088 11612 22098 11619
rect 22268 11619 22279 11665
rect 22459 11619 22470 11665
rect 22640 11665 22650 11672
rect 22268 11612 22278 11619
rect 22460 11612 22470 11619
rect 22640 11619 22651 11665
rect 22640 11612 22650 11619
rect 22712 11578 22770 11702
rect 22832 11665 22842 11672
rect 22831 11619 22842 11665
rect 22832 11612 22842 11619
rect 23012 11612 23214 11672
rect 23384 11665 23394 11672
rect 23384 11619 23395 11665
rect 23384 11612 23394 11619
rect 23084 11578 23142 11612
rect 23456 11578 23514 11702
rect 23576 11665 23586 11672
rect 23575 11619 23586 11665
rect 23756 11665 23766 11672
rect 23948 11665 23958 11672
rect 23576 11612 23586 11619
rect 23756 11619 23767 11665
rect 23947 11619 23958 11665
rect 24128 11665 24138 11672
rect 23756 11612 23766 11619
rect 23948 11612 23958 11619
rect 24128 11619 24139 11665
rect 24128 11612 24138 11619
rect 24200 11578 24258 11702
rect 24320 11665 24330 11672
rect 24319 11619 24330 11665
rect 24320 11612 24330 11619
rect 24500 11612 24572 11672
rect 18682 11190 18689 11566
rect 18723 11190 18730 11566
rect 18682 11138 18730 11190
rect 18941 11566 19101 11578
rect 18941 11190 18947 11566
rect 18981 11190 19061 11566
rect 19095 11190 19101 11566
rect 18941 11178 19101 11190
rect 19313 11566 19473 11578
rect 19313 11190 19319 11566
rect 19353 11190 19433 11566
rect 19467 11190 19473 11566
rect 19313 11178 19473 11190
rect 19685 11566 19845 11578
rect 19685 11190 19691 11566
rect 19725 11190 19805 11566
rect 19839 11190 19845 11566
rect 19685 11178 19845 11190
rect 20057 11566 20217 11578
rect 20057 11190 20063 11566
rect 20097 11190 20177 11566
rect 20211 11190 20217 11566
rect 20057 11178 20217 11190
rect 20429 11566 20589 11578
rect 20429 11190 20435 11566
rect 20469 11190 20549 11566
rect 20583 11190 20589 11566
rect 20429 11178 20589 11190
rect 20801 11566 20961 11578
rect 20801 11190 20807 11566
rect 20841 11190 20921 11566
rect 20955 11190 20961 11566
rect 20801 11178 20961 11190
rect 21173 11566 21333 11578
rect 21173 11190 21179 11566
rect 21213 11190 21293 11566
rect 21327 11190 21333 11566
rect 21173 11178 21333 11190
rect 21545 11566 21705 11578
rect 21545 11190 21551 11566
rect 21585 11190 21665 11566
rect 21699 11190 21705 11566
rect 21545 11178 21705 11190
rect 21917 11566 22077 11578
rect 21917 11190 21923 11566
rect 21957 11190 22037 11566
rect 22071 11190 22077 11566
rect 21917 11178 22077 11190
rect 22289 11566 22449 11578
rect 22289 11190 22295 11566
rect 22329 11190 22409 11566
rect 22443 11190 22449 11566
rect 22289 11178 22449 11190
rect 22661 11566 22821 11578
rect 22661 11190 22667 11566
rect 22701 11190 22781 11566
rect 22815 11190 22821 11566
rect 22661 11178 22821 11190
rect 23033 11566 23193 11578
rect 23033 11190 23039 11566
rect 23073 11190 23153 11566
rect 23187 11190 23193 11566
rect 23033 11178 23193 11190
rect 23405 11566 23565 11578
rect 23405 11190 23411 11566
rect 23445 11190 23525 11566
rect 23559 11190 23565 11566
rect 23405 11178 23565 11190
rect 23777 11566 23937 11578
rect 23777 11190 23783 11566
rect 23817 11190 23897 11566
rect 23931 11190 23937 11566
rect 23777 11178 23937 11190
rect 24149 11566 24309 11578
rect 24149 11190 24155 11566
rect 24189 11190 24269 11566
rect 24303 11190 24309 11566
rect 24149 11178 24309 11190
rect 24520 11566 24572 11612
rect 24520 11190 24527 11566
rect 24561 11190 24572 11566
rect 18682 11137 18770 11138
rect 18682 11132 18931 11137
rect 18682 10988 18750 11132
rect 18920 11091 18931 11132
rect 18920 11029 18930 11091
rect 18920 10988 18931 11029
rect 18682 10983 18931 10988
rect 18682 10982 18768 10983
rect 18682 10930 18730 10982
rect 18986 10942 19056 11178
rect 19111 11132 19303 11137
rect 19111 11091 19122 11132
rect 19112 11029 19122 11091
rect 19111 10988 19122 11029
rect 19292 11091 19303 11132
rect 19292 11029 19302 11091
rect 19292 10988 19303 11029
rect 19111 10983 19303 10988
rect 19358 10942 19428 11178
rect 19483 11132 19675 11137
rect 19483 11091 19494 11132
rect 19484 11029 19494 11091
rect 19483 10988 19494 11029
rect 19664 11091 19675 11132
rect 19664 11029 19674 11091
rect 19664 10988 19675 11029
rect 19483 10983 19675 10988
rect 19730 10942 19800 11178
rect 19855 11136 20047 11137
rect 20102 11136 20172 11178
rect 20227 11136 20419 11137
rect 19855 11132 20419 11136
rect 19855 11091 19866 11132
rect 19856 11029 19866 11091
rect 19855 10988 19866 11029
rect 20036 10988 20238 11132
rect 20408 11091 20419 11132
rect 20408 11029 20418 11091
rect 20408 10988 20419 11029
rect 19855 10984 20419 10988
rect 19855 10983 20047 10984
rect 20102 10942 20172 10984
rect 20227 10983 20419 10984
rect 20474 10942 20544 11178
rect 20599 11132 20791 11137
rect 20599 11091 20610 11132
rect 20600 11029 20610 11091
rect 20599 10988 20610 11029
rect 20780 11091 20791 11132
rect 20780 11029 20790 11091
rect 20780 10988 20791 11029
rect 20599 10983 20791 10988
rect 20846 10942 20916 11178
rect 20971 11132 21163 11137
rect 20971 11091 20982 11132
rect 20972 11029 20982 11091
rect 20971 10988 20982 11029
rect 21152 11091 21163 11132
rect 21152 11029 21162 11091
rect 21152 10988 21163 11029
rect 20971 10983 21163 10988
rect 21218 10942 21288 11178
rect 21590 11138 21660 11178
rect 21398 11137 21816 11138
rect 21343 11132 21907 11137
rect 21343 11091 21354 11132
rect 21344 11029 21354 11091
rect 21343 10988 21354 11029
rect 21524 10988 21726 11132
rect 21896 11091 21907 11132
rect 21896 11029 21906 11091
rect 21896 10988 21907 11029
rect 21343 10983 21907 10988
rect 21398 10982 21816 10983
rect 21590 10942 21660 10982
rect 21962 10942 22032 11178
rect 22087 11132 22279 11137
rect 22087 11091 22098 11132
rect 22088 11029 22098 11091
rect 22087 10988 22098 11029
rect 22268 11091 22279 11132
rect 22268 11029 22278 11091
rect 22268 10988 22279 11029
rect 22087 10983 22279 10988
rect 22334 10942 22404 11178
rect 22459 11132 22651 11137
rect 22459 11091 22470 11132
rect 22460 11029 22470 11091
rect 22459 10988 22470 11029
rect 22640 11091 22651 11132
rect 22640 11029 22650 11091
rect 22640 10988 22651 11029
rect 22459 10983 22651 10988
rect 22706 10942 22776 11178
rect 23078 11138 23148 11178
rect 22926 11137 23302 11138
rect 22831 11132 23395 11137
rect 22831 11091 22842 11132
rect 22832 11029 22842 11091
rect 22831 10988 22842 11029
rect 23012 10988 23214 11132
rect 23384 11091 23395 11132
rect 23384 11029 23394 11091
rect 23384 10988 23395 11029
rect 22831 10983 23395 10988
rect 22926 10982 23302 10983
rect 23078 10942 23148 10982
rect 23450 10942 23520 11178
rect 23575 11132 23767 11137
rect 23575 11091 23586 11132
rect 23576 11029 23586 11091
rect 23575 10988 23586 11029
rect 23756 11091 23767 11132
rect 23756 11029 23766 11091
rect 23756 10988 23767 11029
rect 23575 10983 23767 10988
rect 23822 10942 23892 11178
rect 23947 11132 24139 11137
rect 23947 11091 23958 11132
rect 23948 11029 23958 11091
rect 23947 10988 23958 11029
rect 24128 11091 24139 11132
rect 24128 11029 24138 11091
rect 24128 10988 24139 11029
rect 23947 10983 24139 10988
rect 24194 10942 24264 11178
rect 24520 11138 24572 11190
rect 24414 11137 24572 11138
rect 24319 11132 24572 11137
rect 24319 11091 24330 11132
rect 24320 11029 24330 11091
rect 24319 10988 24330 11029
rect 24500 10988 24572 11132
rect 24319 10983 24572 10988
rect 24414 10982 24572 10983
rect 18682 10554 18689 10930
rect 18723 10554 18730 10930
rect 18682 10502 18730 10554
rect 18941 10930 19101 10942
rect 18941 10554 18947 10930
rect 18981 10554 19061 10930
rect 19095 10554 19101 10930
rect 18941 10542 19101 10554
rect 19313 10930 19473 10942
rect 19313 10554 19319 10930
rect 19353 10554 19433 10930
rect 19467 10554 19473 10930
rect 19313 10542 19473 10554
rect 19685 10930 19845 10942
rect 19685 10554 19691 10930
rect 19725 10554 19805 10930
rect 19839 10554 19845 10930
rect 19685 10542 19845 10554
rect 20057 10930 20217 10942
rect 20057 10554 20063 10930
rect 20097 10554 20177 10930
rect 20211 10554 20217 10930
rect 20057 10542 20217 10554
rect 20429 10930 20589 10942
rect 20429 10554 20435 10930
rect 20469 10554 20549 10930
rect 20583 10554 20589 10930
rect 20429 10542 20589 10554
rect 20801 10930 20961 10942
rect 20801 10554 20807 10930
rect 20841 10554 20921 10930
rect 20955 10554 20961 10930
rect 20801 10542 20961 10554
rect 21173 10930 21333 10942
rect 21173 10554 21179 10930
rect 21213 10554 21293 10930
rect 21327 10554 21333 10930
rect 21173 10542 21333 10554
rect 21545 10930 21705 10942
rect 21545 10554 21551 10930
rect 21585 10554 21665 10930
rect 21699 10554 21705 10930
rect 21545 10542 21705 10554
rect 21917 10930 22077 10942
rect 21917 10554 21923 10930
rect 21957 10554 22037 10930
rect 22071 10554 22077 10930
rect 21917 10542 22077 10554
rect 22289 10930 22449 10942
rect 22289 10554 22295 10930
rect 22329 10554 22409 10930
rect 22443 10554 22449 10930
rect 22289 10542 22449 10554
rect 22661 10930 22821 10942
rect 22661 10554 22667 10930
rect 22701 10554 22781 10930
rect 22815 10554 22821 10930
rect 22661 10542 22821 10554
rect 23033 10930 23193 10942
rect 23033 10554 23039 10930
rect 23073 10554 23153 10930
rect 23187 10554 23193 10930
rect 23033 10542 23193 10554
rect 23405 10930 23565 10942
rect 23405 10554 23411 10930
rect 23445 10554 23525 10930
rect 23559 10554 23565 10930
rect 23405 10542 23565 10554
rect 23777 10930 23937 10942
rect 23777 10554 23783 10930
rect 23817 10554 23897 10930
rect 23931 10554 23937 10930
rect 23777 10542 23937 10554
rect 24149 10930 24309 10942
rect 24149 10554 24155 10930
rect 24189 10554 24269 10930
rect 24303 10554 24309 10930
rect 24149 10542 24309 10554
rect 24520 10930 24572 10982
rect 24520 10554 24527 10930
rect 24561 10554 24572 10930
rect 18682 10501 18772 10502
rect 18682 10496 18931 10501
rect 18682 10352 18750 10496
rect 18920 10455 18931 10496
rect 18920 10393 18930 10455
rect 18920 10352 18931 10393
rect 18682 10347 18931 10352
rect 18682 10342 18772 10347
rect 18682 10294 18730 10342
rect 18986 10306 19056 10542
rect 19111 10496 19303 10501
rect 19111 10455 19122 10496
rect 19112 10393 19122 10455
rect 19111 10352 19122 10393
rect 19292 10455 19303 10496
rect 19292 10393 19302 10455
rect 19292 10352 19303 10393
rect 19111 10347 19303 10352
rect 19358 10306 19428 10542
rect 19483 10496 19675 10501
rect 19483 10455 19494 10496
rect 19484 10393 19494 10455
rect 19483 10352 19494 10393
rect 19664 10455 19675 10496
rect 19664 10393 19674 10455
rect 19664 10352 19675 10393
rect 19483 10347 19675 10352
rect 19730 10306 19800 10542
rect 19855 10498 20047 10501
rect 20102 10498 20172 10542
rect 20227 10498 20419 10501
rect 19855 10496 20419 10498
rect 19855 10455 19866 10496
rect 19856 10393 19866 10455
rect 19855 10352 19866 10393
rect 20036 10352 20238 10496
rect 20408 10455 20419 10496
rect 20408 10393 20418 10455
rect 20408 10352 20419 10393
rect 19855 10347 20419 10352
rect 19896 10346 20372 10347
rect 20102 10306 20172 10346
rect 20474 10306 20544 10542
rect 20599 10496 20791 10501
rect 20599 10455 20610 10496
rect 20600 10393 20610 10455
rect 20599 10352 20610 10393
rect 20780 10455 20791 10496
rect 20780 10393 20790 10455
rect 20780 10352 20791 10393
rect 20599 10347 20791 10352
rect 20846 10306 20916 10542
rect 20971 10496 21163 10501
rect 20971 10455 20982 10496
rect 20972 10393 20982 10455
rect 20971 10352 20982 10393
rect 21152 10455 21163 10496
rect 21152 10393 21162 10455
rect 21152 10352 21163 10393
rect 20971 10347 21163 10352
rect 21218 10306 21288 10542
rect 21590 10502 21660 10542
rect 21418 10501 21836 10502
rect 21343 10496 21907 10501
rect 21343 10455 21354 10496
rect 21344 10393 21354 10455
rect 21343 10352 21354 10393
rect 21524 10352 21726 10496
rect 21896 10455 21907 10496
rect 21896 10393 21906 10455
rect 21896 10352 21907 10393
rect 21343 10347 21907 10352
rect 21418 10346 21836 10347
rect 21590 10306 21660 10346
rect 21962 10306 22032 10542
rect 22087 10496 22279 10501
rect 22087 10455 22098 10496
rect 22088 10393 22098 10455
rect 22087 10352 22098 10393
rect 22268 10455 22279 10496
rect 22268 10393 22278 10455
rect 22268 10352 22279 10393
rect 22087 10347 22279 10352
rect 22334 10306 22404 10542
rect 22459 10496 22651 10501
rect 22459 10455 22470 10496
rect 22460 10393 22470 10455
rect 22459 10352 22470 10393
rect 22640 10455 22651 10496
rect 22640 10393 22650 10455
rect 22640 10352 22651 10393
rect 22459 10347 22651 10352
rect 22706 10306 22776 10542
rect 23078 10502 23148 10542
rect 22914 10501 23290 10502
rect 22831 10496 23395 10501
rect 22831 10455 22842 10496
rect 22832 10393 22842 10455
rect 22831 10352 22842 10393
rect 23012 10352 23214 10496
rect 23384 10455 23395 10496
rect 23384 10393 23394 10455
rect 23384 10352 23395 10393
rect 22831 10347 23395 10352
rect 22914 10346 23290 10347
rect 23078 10306 23148 10346
rect 23450 10306 23520 10542
rect 23575 10496 23767 10501
rect 23575 10455 23586 10496
rect 23576 10393 23586 10455
rect 23575 10352 23586 10393
rect 23756 10455 23767 10496
rect 23756 10393 23766 10455
rect 23756 10352 23767 10393
rect 23575 10347 23767 10352
rect 23822 10306 23892 10542
rect 23947 10496 24139 10501
rect 23947 10455 23958 10496
rect 23948 10393 23958 10455
rect 23947 10352 23958 10393
rect 24128 10455 24139 10496
rect 24128 10393 24138 10455
rect 24128 10352 24139 10393
rect 23947 10347 24139 10352
rect 24194 10306 24264 10542
rect 24520 10502 24572 10554
rect 24430 10501 24572 10502
rect 24319 10496 24572 10501
rect 24319 10455 24330 10496
rect 24320 10393 24330 10455
rect 24319 10352 24330 10393
rect 24500 10352 24572 10496
rect 24319 10347 24572 10352
rect 24430 10346 24572 10347
rect 18682 9918 18689 10294
rect 18723 9918 18730 10294
rect 18682 9872 18730 9918
rect 18941 10294 19101 10306
rect 18941 9918 18947 10294
rect 18981 9918 19061 10294
rect 19095 9918 19101 10294
rect 18941 9906 19101 9918
rect 19313 10294 19473 10306
rect 19313 9918 19319 10294
rect 19353 9918 19433 10294
rect 19467 9918 19473 10294
rect 19313 9906 19473 9918
rect 19685 10294 19845 10306
rect 19685 9918 19691 10294
rect 19725 9918 19805 10294
rect 19839 9918 19845 10294
rect 19685 9906 19845 9918
rect 20057 10294 20217 10306
rect 20057 9918 20063 10294
rect 20097 9918 20177 10294
rect 20211 9918 20217 10294
rect 20057 9906 20217 9918
rect 20429 10294 20589 10306
rect 20429 9918 20435 10294
rect 20469 9918 20549 10294
rect 20583 9918 20589 10294
rect 20429 9906 20589 9918
rect 20801 10294 20961 10306
rect 20801 9918 20807 10294
rect 20841 9918 20921 10294
rect 20955 9918 20961 10294
rect 20801 9906 20961 9918
rect 21173 10294 21333 10306
rect 21173 9918 21179 10294
rect 21213 9918 21293 10294
rect 21327 9918 21333 10294
rect 21173 9906 21333 9918
rect 21545 10294 21705 10306
rect 21545 9918 21551 10294
rect 21585 9918 21665 10294
rect 21699 9918 21705 10294
rect 21545 9906 21705 9918
rect 21917 10294 22077 10306
rect 21917 9918 21923 10294
rect 21957 9918 22037 10294
rect 22071 9918 22077 10294
rect 21917 9906 22077 9918
rect 22289 10294 22449 10306
rect 22289 9918 22295 10294
rect 22329 9918 22409 10294
rect 22443 9918 22449 10294
rect 22289 9906 22449 9918
rect 22661 10294 22821 10306
rect 22661 9918 22667 10294
rect 22701 9918 22781 10294
rect 22815 9918 22821 10294
rect 22661 9906 22821 9918
rect 23033 10294 23193 10306
rect 23033 9918 23039 10294
rect 23073 9918 23153 10294
rect 23187 9918 23193 10294
rect 23033 9906 23193 9918
rect 23405 10294 23565 10306
rect 23405 9918 23411 10294
rect 23445 9918 23525 10294
rect 23559 9918 23565 10294
rect 23405 9906 23565 9918
rect 23777 10294 23937 10306
rect 23777 9918 23783 10294
rect 23817 9918 23897 10294
rect 23931 9918 23937 10294
rect 23777 9906 23937 9918
rect 24149 10294 24309 10306
rect 24149 9918 24155 10294
rect 24189 9918 24269 10294
rect 24303 9918 24309 10294
rect 24149 9906 24309 9918
rect 24520 10294 24572 10346
rect 24520 9918 24527 10294
rect 24561 9918 24572 10294
rect 18682 9812 18750 9872
rect 18920 9865 18930 9872
rect 19112 9865 19122 9872
rect 18920 9819 18931 9865
rect 19111 9819 19122 9865
rect 19292 9865 19302 9872
rect 18920 9812 18930 9819
rect 19112 9812 19122 9819
rect 19292 9819 19303 9865
rect 19292 9812 19302 9819
rect 19364 9564 19422 9906
rect 20108 9872 20166 9906
rect 19484 9865 19494 9872
rect 19483 9819 19494 9865
rect 19664 9865 19674 9872
rect 19856 9865 19866 9872
rect 19484 9812 19494 9819
rect 19664 9819 19675 9865
rect 19855 9819 19866 9865
rect 19664 9812 19674 9819
rect 19856 9812 19866 9819
rect 20036 9812 20238 9872
rect 20408 9865 20418 9872
rect 20600 9865 20610 9872
rect 20408 9819 20419 9865
rect 20599 9819 20610 9865
rect 20780 9865 20790 9872
rect 20408 9812 20418 9819
rect 20600 9812 20610 9819
rect 20780 9819 20791 9865
rect 20780 9812 20790 9819
rect 19982 9810 20312 9812
rect 20852 9564 20910 9906
rect 21596 9872 21654 9906
rect 20972 9865 20982 9872
rect 20971 9819 20982 9865
rect 21152 9865 21162 9872
rect 21344 9865 21354 9872
rect 20972 9812 20982 9819
rect 21152 9819 21163 9865
rect 21343 9819 21354 9865
rect 21152 9812 21162 9819
rect 21344 9812 21354 9819
rect 21524 9812 21726 9872
rect 21896 9865 21906 9872
rect 22088 9865 22098 9872
rect 21896 9819 21907 9865
rect 22087 9819 22098 9865
rect 22268 9865 22278 9872
rect 21896 9812 21906 9819
rect 22088 9812 22098 9819
rect 22268 9819 22279 9865
rect 22268 9812 22278 9819
rect 22340 9564 22398 9906
rect 23084 9872 23142 9906
rect 22460 9865 22470 9872
rect 22459 9819 22470 9865
rect 22640 9865 22650 9872
rect 22832 9865 22842 9872
rect 22460 9812 22470 9819
rect 22640 9819 22651 9865
rect 22831 9819 22842 9865
rect 22640 9812 22650 9819
rect 22832 9812 22842 9819
rect 23012 9812 23214 9872
rect 23384 9865 23394 9872
rect 23576 9865 23586 9872
rect 23384 9819 23395 9865
rect 23575 9819 23586 9865
rect 23756 9865 23766 9872
rect 23384 9812 23394 9819
rect 23576 9812 23586 9819
rect 23756 9819 23767 9865
rect 23756 9812 23766 9819
rect 23828 9564 23886 9906
rect 24520 9872 24572 9918
rect 24610 11578 24662 11702
rect 24696 11612 24702 11672
rect 24872 11665 24882 11672
rect 25064 11665 25074 11672
rect 24872 11619 24883 11665
rect 25063 11619 25074 11665
rect 25244 11665 25254 11672
rect 24872 11612 24882 11619
rect 25064 11612 25074 11619
rect 25244 11619 25255 11665
rect 25244 11612 25254 11619
rect 25316 11578 25374 11702
rect 25436 11665 25446 11672
rect 25435 11619 25446 11665
rect 25616 11665 25626 11672
rect 25808 11665 25818 11672
rect 25436 11612 25446 11619
rect 25616 11619 25627 11665
rect 25807 11619 25818 11665
rect 25988 11665 25998 11672
rect 25616 11612 25626 11619
rect 25808 11612 25818 11619
rect 25988 11619 25999 11665
rect 25988 11612 25998 11619
rect 26060 11578 26118 11702
rect 26180 11665 26190 11672
rect 26179 11619 26190 11665
rect 26360 11665 26370 11672
rect 26552 11665 26562 11672
rect 26180 11612 26190 11619
rect 26360 11619 26371 11665
rect 26551 11619 26562 11665
rect 26732 11665 26742 11672
rect 26360 11612 26370 11619
rect 26552 11612 26562 11619
rect 26732 11619 26743 11665
rect 26732 11612 26742 11619
rect 26804 11578 26862 11702
rect 26924 11665 26934 11672
rect 26923 11619 26934 11665
rect 27104 11665 27114 11672
rect 27296 11665 27306 11672
rect 26924 11612 26934 11619
rect 27104 11619 27115 11665
rect 27295 11619 27306 11665
rect 27476 11665 27486 11672
rect 27104 11612 27114 11619
rect 27296 11612 27306 11619
rect 27476 11619 27487 11665
rect 27476 11612 27486 11619
rect 27548 11578 27606 11702
rect 27668 11665 27678 11672
rect 27667 11619 27678 11665
rect 27848 11665 27858 11672
rect 28040 11665 28050 11672
rect 27668 11612 27678 11619
rect 27848 11619 27859 11665
rect 28039 11619 28050 11665
rect 28220 11665 28230 11672
rect 27848 11612 27858 11619
rect 28040 11612 28050 11619
rect 28220 11619 28231 11665
rect 28220 11612 28230 11619
rect 28292 11578 28350 11702
rect 28412 11665 28422 11672
rect 28411 11619 28422 11665
rect 28592 11665 28602 11672
rect 28784 11665 28794 11672
rect 28412 11612 28422 11619
rect 28592 11619 28603 11665
rect 28783 11619 28794 11665
rect 28964 11665 28974 11672
rect 28592 11612 28602 11619
rect 28784 11612 28794 11619
rect 28964 11619 28975 11665
rect 28964 11612 28974 11619
rect 29036 11578 29094 11702
rect 29156 11665 29166 11672
rect 29155 11619 29166 11665
rect 29336 11665 29346 11672
rect 29528 11665 29538 11672
rect 29156 11612 29166 11619
rect 29336 11619 29347 11665
rect 29527 11619 29538 11665
rect 29708 11665 29718 11672
rect 29336 11612 29346 11619
rect 29528 11612 29538 11619
rect 29708 11619 29719 11665
rect 29708 11612 29718 11619
rect 29780 11578 29838 11702
rect 29900 11665 29910 11672
rect 29899 11619 29910 11665
rect 30080 11665 30090 11672
rect 30272 11665 30282 11672
rect 29900 11612 29910 11619
rect 30080 11619 30091 11665
rect 30271 11619 30282 11665
rect 30452 11665 30462 11672
rect 30080 11612 30090 11619
rect 30272 11612 30282 11619
rect 30452 11619 30463 11665
rect 30452 11612 30462 11619
rect 30506 11578 30564 11702
rect 24610 11566 24681 11578
rect 24610 11190 24641 11566
rect 24675 11190 24681 11566
rect 24610 11178 24681 11190
rect 24893 11566 25053 11578
rect 24893 11190 24899 11566
rect 24933 11190 25013 11566
rect 25047 11190 25053 11566
rect 24893 11178 25053 11190
rect 25265 11566 25425 11578
rect 25265 11190 25271 11566
rect 25305 11190 25385 11566
rect 25419 11190 25425 11566
rect 25265 11178 25425 11190
rect 25637 11566 25797 11578
rect 25637 11190 25643 11566
rect 25677 11190 25757 11566
rect 25791 11190 25797 11566
rect 25637 11178 25797 11190
rect 26009 11566 26169 11578
rect 26009 11190 26015 11566
rect 26049 11190 26129 11566
rect 26163 11190 26169 11566
rect 26009 11178 26169 11190
rect 26381 11566 26541 11578
rect 26381 11190 26387 11566
rect 26421 11190 26501 11566
rect 26535 11190 26541 11566
rect 26381 11178 26541 11190
rect 26753 11566 26913 11578
rect 26753 11190 26759 11566
rect 26793 11190 26873 11566
rect 26907 11190 26913 11566
rect 26753 11178 26913 11190
rect 27125 11566 27285 11578
rect 27125 11190 27131 11566
rect 27165 11190 27245 11566
rect 27279 11190 27285 11566
rect 27125 11178 27285 11190
rect 27497 11566 27657 11578
rect 27497 11190 27503 11566
rect 27537 11190 27617 11566
rect 27651 11190 27657 11566
rect 27497 11178 27657 11190
rect 27869 11566 28029 11578
rect 27869 11190 27875 11566
rect 27909 11190 27989 11566
rect 28023 11190 28029 11566
rect 27869 11178 28029 11190
rect 28241 11566 28401 11578
rect 28241 11190 28247 11566
rect 28281 11190 28361 11566
rect 28395 11190 28401 11566
rect 28241 11178 28401 11190
rect 28613 11566 28773 11578
rect 28613 11190 28619 11566
rect 28653 11190 28733 11566
rect 28767 11190 28773 11566
rect 28613 11178 28773 11190
rect 28985 11566 29145 11578
rect 28985 11190 28991 11566
rect 29025 11190 29105 11566
rect 29139 11190 29145 11566
rect 28985 11178 29145 11190
rect 29357 11566 29517 11578
rect 29357 11190 29363 11566
rect 29397 11190 29477 11566
rect 29511 11190 29517 11566
rect 29357 11178 29517 11190
rect 29729 11566 29889 11578
rect 29729 11190 29735 11566
rect 29769 11190 29849 11566
rect 29883 11190 29889 11566
rect 29729 11178 29889 11190
rect 30101 11566 30261 11578
rect 30101 11190 30107 11566
rect 30141 11190 30221 11566
rect 30255 11190 30261 11566
rect 30101 11178 30261 11190
rect 30473 11566 30564 11578
rect 30473 11190 30479 11566
rect 30513 11190 30564 11566
rect 30473 11178 30564 11190
rect 24610 10942 24662 11178
rect 24690 11137 24816 11138
rect 24690 11132 24883 11137
rect 24690 10988 24702 11132
rect 24872 11091 24883 11132
rect 24872 11029 24882 11091
rect 24872 10988 24883 11029
rect 24690 10983 24883 10988
rect 24690 10982 24816 10983
rect 24938 10942 25008 11178
rect 25063 11132 25255 11137
rect 25063 11091 25074 11132
rect 25064 11029 25074 11091
rect 25063 10988 25074 11029
rect 25244 11091 25255 11132
rect 25244 11029 25254 11091
rect 25244 10988 25255 11029
rect 25063 10983 25255 10988
rect 25310 10942 25380 11178
rect 25435 11132 25627 11137
rect 25435 11091 25446 11132
rect 25436 11029 25446 11091
rect 25435 10988 25446 11029
rect 25616 11091 25627 11132
rect 25616 11029 25626 11091
rect 25616 10988 25627 11029
rect 25435 10983 25627 10988
rect 25682 10942 25752 11178
rect 25807 11132 25999 11137
rect 25807 11091 25818 11132
rect 25808 11029 25818 11091
rect 25807 10988 25818 11029
rect 25988 11091 25999 11132
rect 25988 11029 25998 11091
rect 25988 10988 25999 11029
rect 25807 10983 25999 10988
rect 26054 10942 26124 11178
rect 26179 11132 26371 11137
rect 26179 11091 26190 11132
rect 26180 11029 26190 11091
rect 26179 10988 26190 11029
rect 26360 11091 26371 11132
rect 26360 11029 26370 11091
rect 26360 10988 26371 11029
rect 26179 10983 26371 10988
rect 26426 10942 26496 11178
rect 26551 11132 26743 11137
rect 26551 11091 26562 11132
rect 26552 11029 26562 11091
rect 26551 10988 26562 11029
rect 26732 11091 26743 11132
rect 26732 11029 26742 11091
rect 26732 10988 26743 11029
rect 26551 10983 26743 10988
rect 26798 10942 26868 11178
rect 26923 11132 27115 11137
rect 26923 11091 26934 11132
rect 26924 11029 26934 11091
rect 26923 10988 26934 11029
rect 27104 11091 27115 11132
rect 27104 11029 27114 11091
rect 27104 10988 27115 11029
rect 26923 10983 27115 10988
rect 27170 10942 27240 11178
rect 27295 11132 27487 11137
rect 27295 11091 27306 11132
rect 27296 11029 27306 11091
rect 27295 10988 27306 11029
rect 27476 11091 27487 11132
rect 27476 11029 27486 11091
rect 27476 10988 27487 11029
rect 27295 10983 27487 10988
rect 27542 10942 27612 11178
rect 27667 11132 27859 11137
rect 27667 11091 27678 11132
rect 27668 11029 27678 11091
rect 27667 10988 27678 11029
rect 27848 11091 27859 11132
rect 27848 11029 27858 11091
rect 27848 10988 27859 11029
rect 27667 10983 27859 10988
rect 27914 10942 27984 11178
rect 28039 11132 28231 11137
rect 28039 11091 28050 11132
rect 28040 11029 28050 11091
rect 28039 10988 28050 11029
rect 28220 11091 28231 11132
rect 28220 11029 28230 11091
rect 28220 10988 28231 11029
rect 28039 10983 28231 10988
rect 28286 10942 28356 11178
rect 28411 11132 28603 11137
rect 28411 11091 28422 11132
rect 28412 11029 28422 11091
rect 28411 10988 28422 11029
rect 28592 11091 28603 11132
rect 28592 11029 28602 11091
rect 28592 10988 28603 11029
rect 28411 10983 28603 10988
rect 28658 10942 28728 11178
rect 28783 11132 28975 11137
rect 28783 11091 28794 11132
rect 28784 11029 28794 11091
rect 28783 10988 28794 11029
rect 28964 11091 28975 11132
rect 28964 11029 28974 11091
rect 28964 10988 28975 11029
rect 28783 10983 28975 10988
rect 29030 10942 29100 11178
rect 29155 11132 29347 11137
rect 29155 11091 29166 11132
rect 29156 11029 29166 11091
rect 29155 10988 29166 11029
rect 29336 11091 29347 11132
rect 29336 11029 29346 11091
rect 29336 10988 29347 11029
rect 29155 10983 29347 10988
rect 29402 10942 29472 11178
rect 29527 11132 29719 11137
rect 29527 11091 29538 11132
rect 29528 11029 29538 11091
rect 29527 10988 29538 11029
rect 29708 11091 29719 11132
rect 29708 11029 29718 11091
rect 29708 10988 29719 11029
rect 29527 10983 29719 10988
rect 29774 10942 29844 11178
rect 29899 11132 30091 11137
rect 29899 11091 29910 11132
rect 29900 11029 29910 11091
rect 29899 10988 29910 11029
rect 30080 11091 30091 11132
rect 30080 11029 30090 11091
rect 30080 10988 30091 11029
rect 29899 10983 30091 10988
rect 30146 10942 30216 11178
rect 30271 11132 30463 11137
rect 30271 11091 30282 11132
rect 30272 11029 30282 11091
rect 30271 10988 30282 11029
rect 30452 11091 30463 11132
rect 30452 11029 30462 11091
rect 30452 10988 30463 11029
rect 30271 10983 30463 10988
rect 30506 10942 30564 11178
rect 24610 10930 24681 10942
rect 24610 10554 24641 10930
rect 24675 10554 24681 10930
rect 24610 10542 24681 10554
rect 24893 10930 25053 10942
rect 24893 10554 24899 10930
rect 24933 10554 25013 10930
rect 25047 10554 25053 10930
rect 24893 10542 25053 10554
rect 25265 10930 25425 10942
rect 25265 10554 25271 10930
rect 25305 10554 25385 10930
rect 25419 10554 25425 10930
rect 25265 10542 25425 10554
rect 25637 10930 25797 10942
rect 25637 10554 25643 10930
rect 25677 10554 25757 10930
rect 25791 10554 25797 10930
rect 25637 10542 25797 10554
rect 26009 10930 26169 10942
rect 26009 10554 26015 10930
rect 26049 10554 26129 10930
rect 26163 10554 26169 10930
rect 26009 10542 26169 10554
rect 26381 10930 26541 10942
rect 26381 10554 26387 10930
rect 26421 10554 26501 10930
rect 26535 10554 26541 10930
rect 26381 10542 26541 10554
rect 26753 10930 26913 10942
rect 26753 10554 26759 10930
rect 26793 10554 26873 10930
rect 26907 10554 26913 10930
rect 26753 10542 26913 10554
rect 27125 10930 27285 10942
rect 27125 10554 27131 10930
rect 27165 10554 27245 10930
rect 27279 10554 27285 10930
rect 27125 10542 27285 10554
rect 27497 10930 27657 10942
rect 27497 10554 27503 10930
rect 27537 10554 27617 10930
rect 27651 10554 27657 10930
rect 27497 10542 27657 10554
rect 27869 10930 28029 10942
rect 27869 10554 27875 10930
rect 27909 10554 27989 10930
rect 28023 10554 28029 10930
rect 27869 10542 28029 10554
rect 28241 10930 28401 10942
rect 28241 10554 28247 10930
rect 28281 10554 28361 10930
rect 28395 10554 28401 10930
rect 28241 10542 28401 10554
rect 28613 10930 28773 10942
rect 28613 10554 28619 10930
rect 28653 10554 28733 10930
rect 28767 10554 28773 10930
rect 28613 10542 28773 10554
rect 28985 10930 29145 10942
rect 28985 10554 28991 10930
rect 29025 10554 29105 10930
rect 29139 10554 29145 10930
rect 28985 10542 29145 10554
rect 29357 10930 29517 10942
rect 29357 10554 29363 10930
rect 29397 10554 29477 10930
rect 29511 10554 29517 10930
rect 29357 10542 29517 10554
rect 29729 10930 29889 10942
rect 29729 10554 29735 10930
rect 29769 10554 29849 10930
rect 29883 10554 29889 10930
rect 29729 10542 29889 10554
rect 30101 10930 30261 10942
rect 30101 10554 30107 10930
rect 30141 10554 30221 10930
rect 30255 10554 30261 10930
rect 30101 10542 30261 10554
rect 30473 10930 30564 10942
rect 30473 10554 30479 10930
rect 30513 10554 30564 10930
rect 30473 10542 30564 10554
rect 24610 10306 24662 10542
rect 24690 10501 24832 10502
rect 24690 10496 24883 10501
rect 24690 10352 24702 10496
rect 24872 10455 24883 10496
rect 24872 10393 24882 10455
rect 24872 10352 24883 10393
rect 24690 10347 24883 10352
rect 24690 10346 24832 10347
rect 24938 10306 25008 10542
rect 25063 10496 25255 10501
rect 25063 10455 25074 10496
rect 25064 10393 25074 10455
rect 25063 10352 25074 10393
rect 25244 10455 25255 10496
rect 25244 10393 25254 10455
rect 25244 10352 25255 10393
rect 25063 10347 25255 10352
rect 25310 10306 25380 10542
rect 25435 10496 25627 10501
rect 25435 10455 25446 10496
rect 25436 10393 25446 10455
rect 25435 10352 25446 10393
rect 25616 10455 25627 10496
rect 25616 10393 25626 10455
rect 25616 10352 25627 10393
rect 25435 10347 25627 10352
rect 25682 10306 25752 10542
rect 25807 10496 25999 10501
rect 25807 10455 25818 10496
rect 25808 10393 25818 10455
rect 25807 10352 25818 10393
rect 25988 10455 25999 10496
rect 25988 10393 25998 10455
rect 25988 10352 25999 10393
rect 25807 10347 25999 10352
rect 26054 10306 26124 10542
rect 26179 10496 26371 10501
rect 26179 10455 26190 10496
rect 26180 10393 26190 10455
rect 26179 10352 26190 10393
rect 26360 10455 26371 10496
rect 26360 10393 26370 10455
rect 26360 10352 26371 10393
rect 26179 10347 26371 10352
rect 26426 10306 26496 10542
rect 26551 10496 26743 10501
rect 26551 10455 26562 10496
rect 26552 10393 26562 10455
rect 26551 10352 26562 10393
rect 26732 10455 26743 10496
rect 26732 10393 26742 10455
rect 26732 10352 26743 10393
rect 26551 10347 26743 10352
rect 26798 10306 26868 10542
rect 26923 10496 27115 10501
rect 26923 10455 26934 10496
rect 26924 10393 26934 10455
rect 26923 10352 26934 10393
rect 27104 10455 27115 10496
rect 27104 10393 27114 10455
rect 27104 10352 27115 10393
rect 26923 10347 27115 10352
rect 27170 10306 27240 10542
rect 27295 10496 27487 10501
rect 27295 10455 27306 10496
rect 27296 10393 27306 10455
rect 27295 10352 27306 10393
rect 27476 10455 27487 10496
rect 27476 10393 27486 10455
rect 27476 10352 27487 10393
rect 27295 10347 27487 10352
rect 27542 10306 27612 10542
rect 27667 10496 27859 10501
rect 27667 10455 27678 10496
rect 27668 10393 27678 10455
rect 27667 10352 27678 10393
rect 27848 10455 27859 10496
rect 27848 10393 27858 10455
rect 27848 10352 27859 10393
rect 27667 10347 27859 10352
rect 27914 10306 27984 10542
rect 28039 10496 28231 10501
rect 28039 10455 28050 10496
rect 28040 10393 28050 10455
rect 28039 10352 28050 10393
rect 28220 10455 28231 10496
rect 28220 10393 28230 10455
rect 28220 10352 28231 10393
rect 28039 10347 28231 10352
rect 28286 10306 28356 10542
rect 28411 10496 28603 10501
rect 28411 10455 28422 10496
rect 28412 10393 28422 10455
rect 28411 10352 28422 10393
rect 28592 10455 28603 10496
rect 28592 10393 28602 10455
rect 28592 10352 28603 10393
rect 28411 10347 28603 10352
rect 28658 10306 28728 10542
rect 28783 10496 28975 10501
rect 28783 10455 28794 10496
rect 28784 10393 28794 10455
rect 28783 10352 28794 10393
rect 28964 10455 28975 10496
rect 28964 10393 28974 10455
rect 28964 10352 28975 10393
rect 28783 10347 28975 10352
rect 29030 10306 29100 10542
rect 29155 10496 29347 10501
rect 29155 10455 29166 10496
rect 29156 10393 29166 10455
rect 29155 10352 29166 10393
rect 29336 10455 29347 10496
rect 29336 10393 29346 10455
rect 29336 10352 29347 10393
rect 29155 10347 29347 10352
rect 29402 10306 29472 10542
rect 29527 10496 29719 10501
rect 29527 10455 29538 10496
rect 29528 10393 29538 10455
rect 29527 10352 29538 10393
rect 29708 10455 29719 10496
rect 29708 10393 29718 10455
rect 29708 10352 29719 10393
rect 29527 10347 29719 10352
rect 29774 10306 29844 10542
rect 29899 10496 30091 10501
rect 29899 10455 29910 10496
rect 29900 10393 29910 10455
rect 29899 10352 29910 10393
rect 30080 10455 30091 10496
rect 30080 10393 30090 10455
rect 30080 10352 30091 10393
rect 29899 10347 30091 10352
rect 30146 10306 30216 10542
rect 30271 10496 30463 10501
rect 30271 10455 30282 10496
rect 30272 10393 30282 10455
rect 30271 10352 30282 10393
rect 30452 10455 30463 10496
rect 30452 10393 30462 10455
rect 30452 10352 30463 10393
rect 30271 10347 30463 10352
rect 30506 10306 30564 10542
rect 24610 10294 24681 10306
rect 24610 9918 24641 10294
rect 24675 9918 24681 10294
rect 24610 9906 24681 9918
rect 24893 10294 25053 10306
rect 24893 9918 24899 10294
rect 24933 9918 25013 10294
rect 25047 9918 25053 10294
rect 24893 9906 25053 9918
rect 25265 10294 25425 10306
rect 25265 9918 25271 10294
rect 25305 9918 25385 10294
rect 25419 9918 25425 10294
rect 25265 9906 25425 9918
rect 25637 10294 25797 10306
rect 25637 9918 25643 10294
rect 25677 9918 25757 10294
rect 25791 9918 25797 10294
rect 25637 9906 25797 9918
rect 26009 10294 26169 10306
rect 26009 9918 26015 10294
rect 26049 9918 26129 10294
rect 26163 9918 26169 10294
rect 26009 9906 26169 9918
rect 26381 10294 26541 10306
rect 26381 9918 26387 10294
rect 26421 9918 26501 10294
rect 26535 9918 26541 10294
rect 26381 9906 26541 9918
rect 26753 10294 26913 10306
rect 26753 9918 26759 10294
rect 26793 9918 26873 10294
rect 26907 9918 26913 10294
rect 26753 9906 26913 9918
rect 27125 10294 27285 10306
rect 27125 9918 27131 10294
rect 27165 9918 27245 10294
rect 27279 9918 27285 10294
rect 27125 9906 27285 9918
rect 27497 10294 27657 10306
rect 27497 9918 27503 10294
rect 27537 9918 27617 10294
rect 27651 9918 27657 10294
rect 27497 9906 27657 9918
rect 27869 10294 28029 10306
rect 27869 9918 27875 10294
rect 27909 9918 27989 10294
rect 28023 9918 28029 10294
rect 27869 9906 28029 9918
rect 28241 10294 28401 10306
rect 28241 9918 28247 10294
rect 28281 9918 28361 10294
rect 28395 9918 28401 10294
rect 28241 9906 28401 9918
rect 28613 10294 28773 10306
rect 28613 9918 28619 10294
rect 28653 9918 28733 10294
rect 28767 9918 28773 10294
rect 28613 9906 28773 9918
rect 28985 10294 29145 10306
rect 28985 9918 28991 10294
rect 29025 9918 29105 10294
rect 29139 9918 29145 10294
rect 28985 9906 29145 9918
rect 29357 10294 29517 10306
rect 29357 9918 29363 10294
rect 29397 9918 29477 10294
rect 29511 9918 29517 10294
rect 29357 9906 29517 9918
rect 29729 10294 29889 10306
rect 29729 9918 29735 10294
rect 29769 9918 29849 10294
rect 29883 9918 29889 10294
rect 29729 9906 29889 9918
rect 30101 10294 30261 10306
rect 30101 9918 30107 10294
rect 30141 9918 30221 10294
rect 30255 9918 30261 10294
rect 30101 9906 30261 9918
rect 30473 10294 30564 10306
rect 30473 9918 30479 10294
rect 30513 9918 30564 10294
rect 30473 9906 30564 9918
rect 23948 9865 23958 9872
rect 23947 9819 23958 9865
rect 24128 9865 24138 9872
rect 24320 9865 24330 9872
rect 23948 9812 23958 9819
rect 24128 9819 24139 9865
rect 24319 9819 24330 9865
rect 24128 9812 24138 9819
rect 24320 9812 24330 9819
rect 24500 9812 24572 9872
rect 24688 9812 24702 9872
rect 24872 9865 24882 9872
rect 24872 9819 24883 9865
rect 24872 9812 24882 9819
rect 19364 9500 23886 9564
rect 24938 9504 25008 9906
rect 25064 9865 25074 9872
rect 25063 9819 25074 9865
rect 25244 9865 25254 9872
rect 25436 9865 25446 9872
rect 25064 9812 25074 9819
rect 25244 9819 25255 9865
rect 25435 9819 25446 9865
rect 25616 9865 25626 9872
rect 25244 9812 25254 9819
rect 25436 9812 25446 9819
rect 25616 9819 25627 9865
rect 25616 9812 25626 9819
rect 25682 9504 25752 9906
rect 25808 9865 25818 9872
rect 25807 9819 25818 9865
rect 25988 9865 25998 9872
rect 26180 9865 26190 9872
rect 25808 9812 25818 9819
rect 25988 9819 25999 9865
rect 26179 9819 26190 9865
rect 26360 9865 26370 9872
rect 25988 9812 25998 9819
rect 26180 9812 26190 9819
rect 26360 9819 26371 9865
rect 26360 9812 26370 9819
rect 26426 9504 26496 9906
rect 26552 9865 26562 9872
rect 26551 9819 26562 9865
rect 26732 9865 26742 9872
rect 26924 9865 26934 9872
rect 26552 9812 26562 9819
rect 26732 9819 26743 9865
rect 26923 9819 26934 9865
rect 27104 9865 27114 9872
rect 26732 9812 26742 9819
rect 26924 9812 26934 9819
rect 27104 9819 27115 9865
rect 27104 9812 27114 9819
rect 27170 9504 27240 9906
rect 27296 9865 27306 9872
rect 27295 9819 27306 9865
rect 27476 9865 27486 9872
rect 27668 9865 27678 9872
rect 27296 9812 27306 9819
rect 27476 9819 27487 9865
rect 27667 9819 27678 9865
rect 27848 9865 27858 9872
rect 27476 9812 27486 9819
rect 27668 9812 27678 9819
rect 27848 9819 27859 9865
rect 27848 9812 27858 9819
rect 27914 9504 27984 9906
rect 28040 9865 28050 9872
rect 28039 9819 28050 9865
rect 28220 9865 28230 9872
rect 28412 9865 28422 9872
rect 28040 9812 28050 9819
rect 28220 9819 28231 9865
rect 28411 9819 28422 9865
rect 28592 9865 28602 9872
rect 28220 9812 28230 9819
rect 28412 9812 28422 9819
rect 28592 9819 28603 9865
rect 28592 9812 28602 9819
rect 28658 9504 28728 9906
rect 28784 9865 28794 9872
rect 28783 9819 28794 9865
rect 28964 9865 28974 9872
rect 29156 9865 29166 9872
rect 28784 9812 28794 9819
rect 28964 9819 28975 9865
rect 29155 9819 29166 9865
rect 29336 9865 29346 9872
rect 28964 9812 28974 9819
rect 29156 9812 29166 9819
rect 29336 9819 29347 9865
rect 29336 9812 29346 9819
rect 29402 9504 29472 9906
rect 29528 9865 29538 9872
rect 29527 9819 29538 9865
rect 29708 9865 29718 9872
rect 29900 9865 29910 9872
rect 29528 9812 29538 9819
rect 29708 9819 29719 9865
rect 29899 9819 29910 9865
rect 30080 9865 30090 9872
rect 29708 9812 29718 9819
rect 29900 9812 29910 9819
rect 30080 9819 30091 9865
rect 30080 9812 30090 9819
rect 30146 9504 30216 9906
rect 30272 9865 30282 9872
rect 30271 9819 30282 9865
rect 30452 9865 30462 9872
rect 30272 9812 30282 9819
rect 30452 9819 30463 9865
rect 30452 9812 30462 9819
rect 20124 9396 20178 9500
rect 20520 9396 20590 9500
rect 20852 9396 20910 9500
rect 21264 9396 21334 9500
rect 21596 9396 21654 9500
rect 22008 9396 22078 9500
rect 22340 9396 22398 9500
rect 22752 9396 22822 9500
rect 23072 9396 23126 9500
rect 20124 9390 20230 9396
rect 20124 9320 20148 9390
rect 20218 9320 20230 9390
rect 20124 9314 20230 9320
rect 20508 9390 20602 9396
rect 20508 9320 20520 9390
rect 20590 9320 20602 9390
rect 20508 9314 20602 9320
rect 20852 9390 20974 9396
rect 20852 9320 20892 9390
rect 20962 9320 20974 9390
rect 20852 9314 20974 9320
rect 21252 9390 21346 9396
rect 21252 9320 21264 9390
rect 21334 9320 21346 9390
rect 21252 9314 21346 9320
rect 21596 9390 21718 9396
rect 21596 9320 21636 9390
rect 21706 9320 21718 9390
rect 21596 9314 21718 9320
rect 21996 9390 22090 9396
rect 21996 9320 22008 9390
rect 22078 9320 22090 9390
rect 21996 9314 22090 9320
rect 22340 9390 22462 9396
rect 22340 9320 22380 9390
rect 22450 9320 22462 9390
rect 22340 9314 22462 9320
rect 22740 9390 22834 9396
rect 22740 9320 22752 9390
rect 22822 9320 22834 9390
rect 22740 9314 22834 9320
rect 23002 9390 23126 9396
rect 23002 9320 23014 9390
rect 23084 9320 23126 9390
rect 23002 9314 23126 9320
rect 20124 9190 20178 9314
rect 20228 9277 20238 9286
rect 20227 9231 20238 9277
rect 20408 9277 20418 9286
rect 20600 9277 20610 9286
rect 20228 9222 20238 9231
rect 20408 9231 20419 9277
rect 20599 9231 20610 9277
rect 20780 9277 20790 9286
rect 20408 9222 20418 9231
rect 20600 9222 20610 9231
rect 20780 9231 20791 9277
rect 20780 9222 20790 9231
rect 20852 9190 20910 9314
rect 20972 9277 20982 9286
rect 20971 9231 20982 9277
rect 21152 9277 21162 9286
rect 21344 9277 21354 9286
rect 20972 9222 20982 9231
rect 21152 9231 21163 9277
rect 21343 9231 21354 9277
rect 21524 9277 21534 9286
rect 21152 9222 21162 9231
rect 21344 9222 21354 9231
rect 21524 9231 21535 9277
rect 21524 9222 21534 9231
rect 21596 9190 21654 9314
rect 21716 9277 21726 9286
rect 21715 9231 21726 9277
rect 21896 9277 21906 9286
rect 22088 9277 22098 9286
rect 21716 9222 21726 9231
rect 21896 9231 21907 9277
rect 22087 9231 22098 9277
rect 22268 9277 22278 9286
rect 21896 9222 21906 9231
rect 22088 9222 22098 9231
rect 22268 9231 22279 9277
rect 22268 9222 22278 9231
rect 22340 9190 22398 9314
rect 22460 9277 22470 9286
rect 22459 9231 22470 9277
rect 22640 9277 22650 9286
rect 22832 9277 22842 9286
rect 22460 9222 22470 9231
rect 22640 9231 22651 9277
rect 22831 9231 22842 9277
rect 23012 9277 23022 9286
rect 22640 9222 22650 9231
rect 22832 9222 22842 9231
rect 23012 9231 23023 9277
rect 23012 9222 23022 9231
rect 23072 9190 23126 9314
rect 24824 9232 24834 9504
rect 25116 9232 25126 9504
rect 25568 9232 25578 9504
rect 25860 9232 25870 9504
rect 26312 9232 26322 9504
rect 26604 9232 26614 9504
rect 27056 9232 27066 9504
rect 27348 9232 27358 9504
rect 27800 9232 27810 9504
rect 28092 9232 28102 9504
rect 28544 9232 28554 9504
rect 28836 9232 28846 9504
rect 29288 9232 29298 9504
rect 29580 9232 29590 9504
rect 30032 9232 30042 9504
rect 30324 9232 30334 9504
rect 20124 9178 20217 9190
rect 20124 8402 20177 9178
rect 20211 8402 20217 9178
rect 20124 8390 20217 8402
rect 20429 9178 20589 9190
rect 20429 8402 20435 9178
rect 20469 8402 20549 9178
rect 20583 8402 20589 9178
rect 20429 8390 20589 8402
rect 20801 9178 20961 9190
rect 20801 8402 20807 9178
rect 20841 8402 20921 9178
rect 20955 8402 20961 9178
rect 20801 8390 20961 8402
rect 21173 9178 21333 9190
rect 21173 8402 21179 9178
rect 21213 8402 21293 9178
rect 21327 8402 21333 9178
rect 21173 8390 21333 8402
rect 21545 9178 21705 9190
rect 21545 8402 21551 9178
rect 21585 8402 21665 9178
rect 21699 8402 21705 9178
rect 21545 8390 21705 8402
rect 21917 9178 22077 9190
rect 21917 8402 21923 9178
rect 21957 8402 22037 9178
rect 22071 8402 22077 9178
rect 21917 8390 22077 8402
rect 22289 9178 22449 9190
rect 22289 8402 22295 9178
rect 22329 8402 22409 9178
rect 22443 8402 22449 9178
rect 22289 8390 22449 8402
rect 22661 9178 22821 9190
rect 22661 8402 22667 9178
rect 22701 8402 22781 9178
rect 22815 8402 22821 9178
rect 22661 8390 22821 8402
rect 23033 9178 23126 9190
rect 23033 8402 23039 9178
rect 23073 8402 23126 9178
rect 23033 8390 23126 8402
rect 20124 8154 20172 8390
rect 20227 8344 20419 8349
rect 20227 8303 20238 8344
rect 20228 8241 20238 8303
rect 20227 8200 20238 8241
rect 20408 8303 20419 8344
rect 20408 8241 20418 8303
rect 20408 8200 20419 8241
rect 20227 8195 20419 8200
rect 20474 8154 20544 8390
rect 20599 8344 20791 8349
rect 20599 8303 20610 8344
rect 20600 8241 20610 8303
rect 20599 8200 20610 8241
rect 20780 8303 20791 8344
rect 20780 8241 20790 8303
rect 20780 8200 20791 8241
rect 20599 8195 20791 8200
rect 20846 8154 20916 8390
rect 20971 8344 21163 8349
rect 20971 8303 20982 8344
rect 20972 8241 20982 8303
rect 20971 8200 20982 8241
rect 21152 8303 21163 8344
rect 21152 8241 21162 8303
rect 21152 8200 21163 8241
rect 20971 8195 21163 8200
rect 21218 8154 21288 8390
rect 21343 8344 21535 8349
rect 21343 8303 21354 8344
rect 21344 8241 21354 8303
rect 21343 8200 21354 8241
rect 21524 8303 21535 8344
rect 21524 8241 21534 8303
rect 21524 8200 21535 8241
rect 21343 8195 21535 8200
rect 21590 8154 21660 8390
rect 21715 8344 21907 8349
rect 21715 8303 21726 8344
rect 21716 8241 21726 8303
rect 21715 8200 21726 8241
rect 21896 8303 21907 8344
rect 21896 8241 21906 8303
rect 21896 8200 21907 8241
rect 21715 8195 21907 8200
rect 21962 8154 22032 8390
rect 22087 8344 22279 8349
rect 22087 8303 22098 8344
rect 22088 8241 22098 8303
rect 22087 8200 22098 8241
rect 22268 8303 22279 8344
rect 22268 8241 22278 8303
rect 22268 8200 22279 8241
rect 22087 8195 22279 8200
rect 22334 8154 22404 8390
rect 22459 8344 22651 8349
rect 22459 8303 22470 8344
rect 22460 8241 22470 8303
rect 22459 8200 22470 8241
rect 22640 8303 22651 8344
rect 22640 8241 22650 8303
rect 22640 8200 22651 8241
rect 22459 8195 22651 8200
rect 22706 8154 22776 8390
rect 22831 8344 23023 8349
rect 22831 8303 22842 8344
rect 22832 8241 22842 8303
rect 22831 8200 22842 8241
rect 23012 8303 23023 8344
rect 23012 8241 23022 8303
rect 23012 8200 23023 8241
rect 22831 8195 23023 8200
rect 23072 8154 23126 8390
rect 20124 8142 20217 8154
rect 20124 7366 20177 8142
rect 20211 7366 20217 8142
rect 20124 7354 20217 7366
rect 20429 8142 20589 8154
rect 20429 7366 20435 8142
rect 20469 7366 20549 8142
rect 20583 7366 20589 8142
rect 20429 7354 20589 7366
rect 20801 8142 20961 8154
rect 20801 7366 20807 8142
rect 20841 7366 20921 8142
rect 20955 7366 20961 8142
rect 20801 7354 20961 7366
rect 21173 8142 21333 8154
rect 21173 7366 21179 8142
rect 21213 7366 21293 8142
rect 21327 7366 21333 8142
rect 21173 7354 21333 7366
rect 21545 8142 21705 8154
rect 21545 7366 21551 8142
rect 21585 7366 21665 8142
rect 21699 7366 21705 8142
rect 21545 7354 21705 7366
rect 21917 8142 22077 8154
rect 21917 7366 21923 8142
rect 21957 7366 22037 8142
rect 22071 7366 22077 8142
rect 21917 7354 22077 7366
rect 22289 8142 22449 8154
rect 22289 7366 22295 8142
rect 22329 7366 22409 8142
rect 22443 7366 22449 8142
rect 22289 7354 22449 7366
rect 22661 8142 22821 8154
rect 22661 7366 22667 8142
rect 22701 7366 22781 8142
rect 22815 7366 22821 8142
rect 22661 7354 22821 7366
rect 23033 8142 23126 8154
rect 23033 7366 23039 8142
rect 23073 7366 23126 8142
rect 23706 7516 23716 7788
rect 23998 7516 24008 7788
rect 23033 7354 23126 7366
rect 20124 7118 20172 7354
rect 20227 7308 20419 7313
rect 20227 7267 20238 7308
rect 20228 7205 20238 7267
rect 20227 7164 20238 7205
rect 20408 7267 20419 7308
rect 20408 7205 20418 7267
rect 20408 7164 20419 7205
rect 20227 7159 20419 7164
rect 20474 7118 20544 7354
rect 20599 7308 20791 7313
rect 20599 7267 20610 7308
rect 20600 7205 20610 7267
rect 20599 7164 20610 7205
rect 20780 7267 20791 7308
rect 20780 7205 20790 7267
rect 20780 7164 20791 7205
rect 20599 7159 20791 7164
rect 20846 7118 20916 7354
rect 20971 7308 21163 7313
rect 20971 7267 20982 7308
rect 20972 7205 20982 7267
rect 20971 7164 20982 7205
rect 21152 7267 21163 7308
rect 21152 7205 21162 7267
rect 21152 7164 21163 7205
rect 20971 7159 21163 7164
rect 21218 7118 21288 7354
rect 21343 7308 21535 7313
rect 21343 7267 21354 7308
rect 21344 7205 21354 7267
rect 21343 7164 21354 7205
rect 21524 7267 21535 7308
rect 21524 7205 21534 7267
rect 21524 7164 21535 7205
rect 21343 7159 21535 7164
rect 21590 7118 21660 7354
rect 21715 7308 21907 7313
rect 21715 7267 21726 7308
rect 21716 7205 21726 7267
rect 21715 7164 21726 7205
rect 21896 7267 21907 7308
rect 21896 7205 21906 7267
rect 21896 7164 21907 7205
rect 21715 7159 21907 7164
rect 21962 7118 22032 7354
rect 22087 7308 22279 7313
rect 22087 7267 22098 7308
rect 22088 7205 22098 7267
rect 22087 7164 22098 7205
rect 22268 7267 22279 7308
rect 22268 7205 22278 7267
rect 22268 7164 22279 7205
rect 22087 7159 22279 7164
rect 22334 7118 22404 7354
rect 22459 7308 22651 7313
rect 22459 7267 22470 7308
rect 22460 7205 22470 7267
rect 22459 7164 22470 7205
rect 22640 7267 22651 7308
rect 22640 7205 22650 7267
rect 22640 7164 22651 7205
rect 22459 7159 22651 7164
rect 22706 7118 22776 7354
rect 22831 7308 23023 7313
rect 22831 7267 22842 7308
rect 22832 7205 22842 7267
rect 22831 7164 22842 7205
rect 23012 7267 23023 7308
rect 23012 7205 23022 7267
rect 23012 7164 23023 7205
rect 22831 7159 23023 7164
rect 23072 7118 23126 7354
rect 20124 7106 20217 7118
rect 20124 6330 20177 7106
rect 20211 6330 20217 7106
rect 20124 6318 20217 6330
rect 20429 7106 20589 7118
rect 20429 6330 20435 7106
rect 20469 6330 20549 7106
rect 20583 6330 20589 7106
rect 20429 6318 20589 6330
rect 20801 7106 20961 7118
rect 20801 6330 20807 7106
rect 20841 6330 20921 7106
rect 20955 6330 20961 7106
rect 20801 6318 20961 6330
rect 21173 7106 21333 7118
rect 21173 6330 21179 7106
rect 21213 6330 21293 7106
rect 21327 6330 21333 7106
rect 21173 6318 21333 6330
rect 21545 7106 21705 7118
rect 21545 6330 21551 7106
rect 21585 6330 21665 7106
rect 21699 6330 21705 7106
rect 21545 6318 21705 6330
rect 21917 7106 22077 7118
rect 21917 6330 21923 7106
rect 21957 6330 22037 7106
rect 22071 6330 22077 7106
rect 21917 6318 22077 6330
rect 22289 7106 22449 7118
rect 22289 6330 22295 7106
rect 22329 6330 22409 7106
rect 22443 6330 22449 7106
rect 22289 6318 22449 6330
rect 22661 7106 22821 7118
rect 22661 6330 22667 7106
rect 22701 6330 22781 7106
rect 22815 6330 22821 7106
rect 22661 6318 22821 6330
rect 23033 7106 23126 7118
rect 23033 6330 23039 7106
rect 23073 6330 23126 7106
rect 23818 7311 23890 7516
rect 23818 6914 23835 7311
rect 23873 6914 23890 7311
rect 23818 6896 23890 6914
rect 24122 6822 24132 6886
rect 23958 6816 24132 6822
rect 23958 6756 23970 6816
rect 24034 6756 24132 6816
rect 23958 6750 24132 6756
rect 24122 6688 24132 6750
rect 24330 6688 24340 6886
rect 24122 6422 24132 6486
rect 23958 6416 24132 6422
rect 23958 6356 23970 6416
rect 24034 6356 24132 6416
rect 23958 6350 24132 6356
rect 23033 6318 23126 6330
rect 20124 6082 20172 6318
rect 20227 6272 20419 6277
rect 20227 6231 20238 6272
rect 20228 6169 20238 6231
rect 20227 6128 20238 6169
rect 20408 6231 20419 6272
rect 20408 6169 20418 6231
rect 20408 6128 20419 6169
rect 20227 6123 20419 6128
rect 20474 6082 20544 6318
rect 20599 6272 20791 6277
rect 20599 6231 20610 6272
rect 20600 6169 20610 6231
rect 20599 6128 20610 6169
rect 20780 6231 20791 6272
rect 20780 6169 20790 6231
rect 20780 6128 20791 6169
rect 20599 6123 20791 6128
rect 20846 6082 20916 6318
rect 20971 6272 21163 6277
rect 20971 6231 20982 6272
rect 20972 6169 20982 6231
rect 20971 6128 20982 6169
rect 21152 6231 21163 6272
rect 21152 6169 21162 6231
rect 21152 6128 21163 6169
rect 20971 6123 21163 6128
rect 21218 6082 21288 6318
rect 21343 6272 21535 6277
rect 21343 6231 21354 6272
rect 21344 6169 21354 6231
rect 21343 6128 21354 6169
rect 21524 6231 21535 6272
rect 21524 6169 21534 6231
rect 21524 6128 21535 6169
rect 21343 6123 21535 6128
rect 21590 6082 21660 6318
rect 21715 6272 21907 6277
rect 21715 6231 21726 6272
rect 21716 6169 21726 6231
rect 21715 6128 21726 6169
rect 21896 6231 21907 6272
rect 21896 6169 21906 6231
rect 21896 6128 21907 6169
rect 21715 6123 21907 6128
rect 21962 6082 22032 6318
rect 22087 6272 22279 6277
rect 22087 6231 22098 6272
rect 22088 6169 22098 6231
rect 22087 6128 22098 6169
rect 22268 6231 22279 6272
rect 22268 6169 22278 6231
rect 22268 6128 22279 6169
rect 22087 6123 22279 6128
rect 22334 6082 22404 6318
rect 22459 6272 22651 6277
rect 22459 6231 22470 6272
rect 22460 6169 22470 6231
rect 22459 6128 22470 6169
rect 22640 6231 22651 6272
rect 22640 6169 22650 6231
rect 22640 6128 22651 6169
rect 22459 6123 22651 6128
rect 22706 6082 22776 6318
rect 22831 6272 23023 6277
rect 22831 6231 22842 6272
rect 22832 6169 22842 6231
rect 22831 6128 22842 6169
rect 23012 6231 23023 6272
rect 23012 6169 23022 6231
rect 23012 6128 23023 6169
rect 22831 6123 23023 6128
rect 23072 6082 23126 6318
rect 20124 6070 20217 6082
rect 20124 5294 20177 6070
rect 20211 5294 20217 6070
rect 20124 5282 20217 5294
rect 20429 6070 20589 6082
rect 20429 5294 20435 6070
rect 20469 5294 20549 6070
rect 20583 5294 20589 6070
rect 20429 5282 20589 5294
rect 20801 6070 20961 6082
rect 20801 5294 20807 6070
rect 20841 5294 20921 6070
rect 20955 5294 20961 6070
rect 20801 5282 20961 5294
rect 21173 6070 21333 6082
rect 21173 5294 21179 6070
rect 21213 5294 21293 6070
rect 21327 5294 21333 6070
rect 21173 5282 21333 5294
rect 21545 6070 21705 6082
rect 21545 5294 21551 6070
rect 21585 5294 21665 6070
rect 21699 5294 21705 6070
rect 21545 5282 21705 5294
rect 21917 6070 22077 6082
rect 21917 5294 21923 6070
rect 21957 5294 22037 6070
rect 22071 5294 22077 6070
rect 21917 5282 22077 5294
rect 22289 6070 22449 6082
rect 22289 5294 22295 6070
rect 22329 5294 22409 6070
rect 22443 5294 22449 6070
rect 22289 5282 22449 5294
rect 22661 6070 22821 6082
rect 22661 5294 22667 6070
rect 22701 5294 22781 6070
rect 22815 5294 22821 6070
rect 22661 5282 22821 5294
rect 23033 6070 23126 6082
rect 23033 5294 23039 6070
rect 23073 5294 23126 6070
rect 23818 6320 23890 6336
rect 23818 5923 23835 6320
rect 23873 5923 23890 6320
rect 24122 6288 24132 6350
rect 24330 6288 24340 6486
rect 24122 6022 24132 6086
rect 23958 6016 24132 6022
rect 23958 5956 23970 6016
rect 24034 5956 24132 6016
rect 23958 5950 24132 5956
rect 23033 5282 23126 5294
rect 20228 5241 20238 5246
rect 20227 5195 20238 5241
rect 20408 5241 20418 5246
rect 20228 5192 20238 5195
rect 20408 5195 20419 5241
rect 20408 5192 20418 5195
rect 20474 4598 20544 5282
rect 20600 5241 20610 5246
rect 20599 5195 20610 5241
rect 20780 5241 20790 5246
rect 20972 5241 20982 5246
rect 20600 5192 20610 5195
rect 20780 5195 20791 5241
rect 20971 5195 20982 5241
rect 21152 5241 21162 5246
rect 20780 5192 20790 5195
rect 20972 5192 20982 5195
rect 21152 5195 21163 5241
rect 21152 5192 21162 5195
rect 21218 4906 21288 5282
rect 21344 5241 21354 5246
rect 21343 5195 21354 5241
rect 21524 5241 21534 5246
rect 21716 5241 21726 5246
rect 21344 5192 21354 5195
rect 21524 5195 21535 5241
rect 21715 5195 21726 5241
rect 21896 5241 21906 5246
rect 21524 5192 21534 5195
rect 21716 5192 21726 5195
rect 21896 5195 21907 5241
rect 21896 5192 21906 5195
rect 21962 4906 22032 5282
rect 22088 5241 22098 5246
rect 22087 5195 22098 5241
rect 22268 5241 22278 5246
rect 22460 5241 22470 5246
rect 22088 5192 22098 5195
rect 22268 5195 22279 5241
rect 22459 5195 22470 5241
rect 22640 5241 22650 5246
rect 22268 5192 22278 5195
rect 22460 5192 22470 5195
rect 22640 5195 22651 5241
rect 22640 5192 22650 5195
rect 21208 4726 21218 4906
rect 22032 4726 22042 4906
rect 20226 4588 20792 4598
rect 20226 4542 20238 4588
rect 20227 4537 20238 4542
rect 20228 4532 20238 4537
rect 20408 4542 20610 4588
rect 20408 4537 20419 4542
rect 20408 4532 20418 4537
rect 20122 4505 20196 4506
rect 20474 4505 20544 4542
rect 20599 4537 20610 4542
rect 20600 4532 20610 4537
rect 20780 4542 20792 4588
rect 20972 4583 20982 4588
rect 20780 4537 20791 4542
rect 20971 4537 20982 4583
rect 21152 4583 21162 4588
rect 20780 4532 20790 4537
rect 20972 4532 20982 4537
rect 21152 4537 21163 4583
rect 21152 4532 21162 4537
rect 20846 4505 20916 4506
rect 21218 4505 21288 4726
rect 21344 4583 21354 4588
rect 21343 4537 21354 4583
rect 21524 4583 21534 4588
rect 21716 4583 21726 4588
rect 21344 4532 21354 4537
rect 21524 4537 21535 4583
rect 21715 4537 21726 4583
rect 21896 4583 21906 4588
rect 21524 4532 21534 4537
rect 21716 4532 21726 4537
rect 21896 4537 21907 4583
rect 21896 4532 21906 4537
rect 21590 4505 21660 4506
rect 21962 4505 22032 4726
rect 22706 4598 22776 5282
rect 22832 5241 22842 5246
rect 22831 5195 22842 5241
rect 23012 5241 23022 5246
rect 22832 5192 22842 5195
rect 23012 5195 23023 5241
rect 23012 5192 23022 5195
rect 23334 5050 23344 5322
rect 23626 5050 23636 5322
rect 22458 4588 23024 4598
rect 22088 4583 22098 4588
rect 22087 4537 22098 4583
rect 22268 4583 22278 4588
rect 22088 4532 22098 4537
rect 22268 4537 22279 4583
rect 22458 4542 22470 4588
rect 22459 4537 22470 4542
rect 22268 4532 22278 4537
rect 22460 4532 22470 4537
rect 22640 4542 22842 4588
rect 22640 4537 22651 4542
rect 22640 4532 22650 4537
rect 22334 4505 22404 4506
rect 22706 4505 22776 4542
rect 22831 4537 22842 4542
rect 22832 4532 22842 4537
rect 23012 4542 23024 4588
rect 23204 4583 23214 4588
rect 23012 4537 23023 4542
rect 23203 4537 23214 4583
rect 23384 4583 23394 4588
rect 23012 4532 23022 4537
rect 23204 4532 23214 4537
rect 23384 4537 23395 4583
rect 23384 4532 23394 4537
rect 23078 4505 23148 4506
rect 23450 4505 23520 5050
rect 23818 4976 23890 5923
rect 24122 5888 24132 5950
rect 24330 5888 24340 6086
rect 24078 5050 24088 5322
rect 24370 5050 24380 5322
rect 24822 5050 24832 5322
rect 25114 5050 25124 5322
rect 25566 5050 25576 5322
rect 25858 5050 25868 5322
rect 26310 5050 26320 5322
rect 26602 5050 26612 5322
rect 27054 5050 27064 5322
rect 27346 5050 27356 5322
rect 27798 5050 27808 5322
rect 28090 5050 28100 5322
rect 28542 5050 28552 5322
rect 28834 5050 28844 5322
rect 23714 4726 23724 4976
rect 23974 4726 23984 4976
rect 23576 4583 23586 4588
rect 23575 4537 23586 4583
rect 23756 4583 23766 4588
rect 23948 4583 23958 4588
rect 23576 4532 23586 4537
rect 23756 4537 23767 4583
rect 23947 4537 23958 4583
rect 24128 4583 24138 4588
rect 23756 4532 23766 4537
rect 23948 4532 23958 4537
rect 24128 4537 24139 4583
rect 24128 4532 24138 4537
rect 23822 4505 23892 4506
rect 24194 4505 24264 5050
rect 24320 4583 24330 4588
rect 24319 4537 24330 4583
rect 24500 4583 24510 4588
rect 24692 4583 24702 4588
rect 24320 4532 24330 4537
rect 24500 4537 24511 4583
rect 24691 4537 24702 4583
rect 24872 4583 24882 4588
rect 24500 4532 24510 4537
rect 24692 4532 24702 4537
rect 24872 4537 24883 4583
rect 24872 4532 24882 4537
rect 24566 4505 24636 4506
rect 24938 4505 25008 5050
rect 25064 4583 25074 4588
rect 25063 4537 25074 4583
rect 25244 4583 25254 4588
rect 25436 4583 25446 4588
rect 25064 4532 25074 4537
rect 25244 4537 25255 4583
rect 25435 4537 25446 4583
rect 25616 4583 25626 4588
rect 25244 4532 25254 4537
rect 25436 4532 25446 4537
rect 25616 4537 25627 4583
rect 25616 4532 25626 4537
rect 25310 4505 25380 4506
rect 25682 4505 25752 5050
rect 25808 4583 25818 4588
rect 25807 4537 25818 4583
rect 25988 4583 25998 4588
rect 26180 4583 26190 4588
rect 25808 4532 25818 4537
rect 25988 4537 25999 4583
rect 26179 4537 26190 4583
rect 26360 4583 26370 4588
rect 25988 4532 25998 4537
rect 26180 4532 26190 4537
rect 26360 4537 26371 4583
rect 26360 4532 26370 4537
rect 26054 4505 26124 4506
rect 26426 4505 26496 5050
rect 26552 4583 26562 4588
rect 26551 4537 26562 4583
rect 26732 4583 26742 4588
rect 26924 4583 26934 4588
rect 26552 4532 26562 4537
rect 26732 4537 26743 4583
rect 26923 4537 26934 4583
rect 27104 4583 27114 4588
rect 26732 4532 26742 4537
rect 26924 4532 26934 4537
rect 27104 4537 27115 4583
rect 27104 4532 27114 4537
rect 26798 4505 26868 4506
rect 27170 4505 27240 5050
rect 27296 4583 27306 4588
rect 27295 4537 27306 4583
rect 27476 4583 27486 4588
rect 27668 4583 27678 4588
rect 27296 4532 27306 4537
rect 27476 4537 27487 4583
rect 27667 4537 27678 4583
rect 27848 4583 27858 4588
rect 27476 4532 27486 4537
rect 27668 4532 27678 4537
rect 27848 4537 27859 4583
rect 27848 4532 27858 4537
rect 27542 4505 27612 4506
rect 27914 4505 27984 5050
rect 28040 4583 28050 4588
rect 28039 4537 28050 4583
rect 28220 4583 28230 4588
rect 28412 4583 28422 4588
rect 28040 4532 28050 4537
rect 28220 4537 28231 4583
rect 28411 4537 28422 4583
rect 28592 4583 28602 4588
rect 28220 4532 28230 4537
rect 28412 4532 28422 4537
rect 28592 4537 28603 4583
rect 28592 4532 28602 4537
rect 28286 4505 28356 4506
rect 28658 4505 28728 5050
rect 28784 4583 28794 4588
rect 28783 4537 28794 4583
rect 28964 4583 28974 4588
rect 28784 4532 28794 4537
rect 28964 4537 28975 4583
rect 28964 4532 28974 4537
rect 29006 4505 29080 4518
rect 20122 4493 20217 4505
rect 20122 4317 20177 4493
rect 20211 4317 20217 4493
rect 20122 4305 20217 4317
rect 20429 4493 20589 4505
rect 20429 4317 20435 4493
rect 20469 4317 20549 4493
rect 20583 4317 20589 4493
rect 20429 4305 20589 4317
rect 20801 4493 20961 4505
rect 20801 4317 20807 4493
rect 20841 4317 20921 4493
rect 20955 4317 20961 4493
rect 20801 4305 20961 4317
rect 21173 4493 21333 4505
rect 21173 4317 21179 4493
rect 21213 4317 21293 4493
rect 21327 4317 21333 4493
rect 21173 4305 21333 4317
rect 21545 4493 21705 4505
rect 21545 4317 21551 4493
rect 21585 4317 21665 4493
rect 21699 4317 21705 4493
rect 21545 4305 21705 4317
rect 21917 4493 22077 4505
rect 21917 4317 21923 4493
rect 21957 4317 22037 4493
rect 22071 4317 22077 4493
rect 21917 4305 22077 4317
rect 22289 4493 22449 4505
rect 22289 4317 22295 4493
rect 22329 4317 22409 4493
rect 22443 4317 22449 4493
rect 22289 4305 22449 4317
rect 22661 4493 22821 4505
rect 22661 4317 22667 4493
rect 22701 4317 22781 4493
rect 22815 4317 22821 4493
rect 22661 4305 22821 4317
rect 23033 4493 23193 4505
rect 23033 4317 23039 4493
rect 23073 4317 23153 4493
rect 23187 4317 23193 4493
rect 23033 4305 23193 4317
rect 23405 4493 23565 4505
rect 23405 4317 23411 4493
rect 23445 4317 23525 4493
rect 23559 4317 23565 4493
rect 23405 4305 23565 4317
rect 23777 4493 23937 4505
rect 23777 4317 23783 4493
rect 23817 4317 23897 4493
rect 23931 4317 23937 4493
rect 23777 4305 23937 4317
rect 24149 4493 24309 4505
rect 24149 4317 24155 4493
rect 24189 4317 24269 4493
rect 24303 4317 24309 4493
rect 24149 4305 24309 4317
rect 24521 4493 24681 4505
rect 24521 4317 24527 4493
rect 24561 4317 24641 4493
rect 24675 4317 24681 4493
rect 24521 4305 24681 4317
rect 24893 4493 25053 4505
rect 24893 4317 24899 4493
rect 24933 4317 25013 4493
rect 25047 4317 25053 4493
rect 24893 4305 25053 4317
rect 25265 4493 25425 4505
rect 25265 4317 25271 4493
rect 25305 4317 25385 4493
rect 25419 4317 25425 4493
rect 25265 4305 25425 4317
rect 25637 4493 25797 4505
rect 25637 4317 25643 4493
rect 25677 4317 25757 4493
rect 25791 4317 25797 4493
rect 25637 4305 25797 4317
rect 26009 4493 26169 4505
rect 26009 4317 26015 4493
rect 26049 4317 26129 4493
rect 26163 4317 26169 4493
rect 26009 4305 26169 4317
rect 26381 4493 26541 4505
rect 26381 4317 26387 4493
rect 26421 4317 26501 4493
rect 26535 4317 26541 4493
rect 26381 4305 26541 4317
rect 26753 4493 26913 4505
rect 26753 4317 26759 4493
rect 26793 4317 26873 4493
rect 26907 4317 26913 4493
rect 26753 4305 26913 4317
rect 27125 4493 27285 4505
rect 27125 4317 27131 4493
rect 27165 4317 27245 4493
rect 27279 4317 27285 4493
rect 27125 4305 27285 4317
rect 27497 4493 27657 4505
rect 27497 4317 27503 4493
rect 27537 4317 27617 4493
rect 27651 4317 27657 4493
rect 27497 4305 27657 4317
rect 27869 4493 28029 4505
rect 27869 4317 27875 4493
rect 27909 4317 27989 4493
rect 28023 4317 28029 4493
rect 27869 4305 28029 4317
rect 28241 4493 28401 4505
rect 28241 4317 28247 4493
rect 28281 4317 28361 4493
rect 28395 4317 28401 4493
rect 28241 4305 28401 4317
rect 28613 4493 28773 4505
rect 28613 4317 28619 4493
rect 28653 4317 28733 4493
rect 28767 4317 28773 4493
rect 28613 4305 28773 4317
rect 28985 4493 29080 4505
rect 28985 4317 28991 4493
rect 29025 4317 29080 4493
rect 28985 4305 29080 4317
rect 20122 4087 20196 4305
rect 20474 4274 20544 4305
rect 20226 4268 20792 4274
rect 20226 4124 20238 4268
rect 20408 4124 20610 4268
rect 20780 4124 20792 4268
rect 20226 4118 20792 4124
rect 20474 4087 20544 4118
rect 20846 4087 20916 4305
rect 20971 4268 21163 4273
rect 20971 4227 20982 4268
rect 20972 4165 20982 4227
rect 20971 4124 20982 4165
rect 21152 4227 21163 4268
rect 21152 4165 21162 4227
rect 21152 4124 21163 4165
rect 20971 4119 21163 4124
rect 21218 4087 21288 4305
rect 21343 4268 21535 4273
rect 21343 4227 21354 4268
rect 21344 4165 21354 4227
rect 21343 4124 21354 4165
rect 21524 4227 21535 4268
rect 21524 4165 21534 4227
rect 21524 4124 21535 4165
rect 21343 4119 21535 4124
rect 21590 4087 21660 4305
rect 21715 4268 21907 4273
rect 21715 4227 21726 4268
rect 21716 4165 21726 4227
rect 21715 4124 21726 4165
rect 21896 4227 21907 4268
rect 21896 4165 21906 4227
rect 21896 4124 21907 4165
rect 21715 4119 21907 4124
rect 21962 4087 22032 4305
rect 22087 4268 22279 4273
rect 22087 4227 22098 4268
rect 22088 4165 22098 4227
rect 22087 4124 22098 4165
rect 22268 4227 22279 4268
rect 22268 4165 22278 4227
rect 22268 4124 22279 4165
rect 22087 4119 22279 4124
rect 22334 4087 22404 4305
rect 22706 4274 22776 4305
rect 22458 4268 23024 4274
rect 22458 4124 22470 4268
rect 22640 4124 22842 4268
rect 23012 4124 23024 4268
rect 22458 4118 23024 4124
rect 22706 4087 22776 4118
rect 23078 4087 23148 4305
rect 23203 4268 23395 4273
rect 23203 4227 23214 4268
rect 23204 4165 23214 4227
rect 23203 4124 23214 4165
rect 23384 4227 23395 4268
rect 23384 4165 23394 4227
rect 23384 4124 23395 4165
rect 23203 4119 23395 4124
rect 23450 4087 23520 4305
rect 23575 4268 23767 4273
rect 23575 4227 23586 4268
rect 23576 4165 23586 4227
rect 23575 4124 23586 4165
rect 23756 4227 23767 4268
rect 23756 4165 23766 4227
rect 23756 4124 23767 4165
rect 23575 4119 23767 4124
rect 23822 4087 23892 4305
rect 23947 4268 24139 4273
rect 23947 4227 23958 4268
rect 23948 4165 23958 4227
rect 23947 4124 23958 4165
rect 24128 4227 24139 4268
rect 24128 4165 24138 4227
rect 24128 4124 24139 4165
rect 23947 4119 24139 4124
rect 24194 4087 24264 4305
rect 24319 4268 24511 4273
rect 24319 4227 24330 4268
rect 24320 4165 24330 4227
rect 24319 4124 24330 4165
rect 24500 4227 24511 4268
rect 24500 4165 24510 4227
rect 24500 4124 24511 4165
rect 24319 4119 24511 4124
rect 24566 4087 24636 4305
rect 24691 4268 24883 4273
rect 24691 4227 24702 4268
rect 24692 4165 24702 4227
rect 24691 4124 24702 4165
rect 24872 4227 24883 4268
rect 24872 4165 24882 4227
rect 24872 4124 24883 4165
rect 24691 4119 24883 4124
rect 24938 4087 25008 4305
rect 25063 4268 25255 4273
rect 25063 4227 25074 4268
rect 25064 4165 25074 4227
rect 25063 4124 25074 4165
rect 25244 4227 25255 4268
rect 25244 4165 25254 4227
rect 25244 4124 25255 4165
rect 25063 4119 25255 4124
rect 25310 4087 25380 4305
rect 25435 4268 25627 4273
rect 25435 4227 25446 4268
rect 25436 4165 25446 4227
rect 25435 4124 25446 4165
rect 25616 4227 25627 4268
rect 25616 4165 25626 4227
rect 25616 4124 25627 4165
rect 25435 4119 25627 4124
rect 25682 4087 25752 4305
rect 25807 4268 25999 4273
rect 25807 4227 25818 4268
rect 25808 4165 25818 4227
rect 25807 4124 25818 4165
rect 25988 4227 25999 4268
rect 25988 4165 25998 4227
rect 25988 4124 25999 4165
rect 25807 4119 25999 4124
rect 26054 4087 26124 4305
rect 26179 4268 26371 4273
rect 26179 4227 26190 4268
rect 26180 4165 26190 4227
rect 26179 4124 26190 4165
rect 26360 4227 26371 4268
rect 26360 4165 26370 4227
rect 26360 4124 26371 4165
rect 26179 4119 26371 4124
rect 26426 4087 26496 4305
rect 26551 4268 26743 4273
rect 26551 4227 26562 4268
rect 26552 4165 26562 4227
rect 26551 4124 26562 4165
rect 26732 4227 26743 4268
rect 26732 4165 26742 4227
rect 26732 4124 26743 4165
rect 26551 4119 26743 4124
rect 26798 4087 26868 4305
rect 26923 4268 27115 4273
rect 26923 4227 26934 4268
rect 26924 4165 26934 4227
rect 26923 4124 26934 4165
rect 27104 4227 27115 4268
rect 27104 4165 27114 4227
rect 27104 4124 27115 4165
rect 26923 4119 27115 4124
rect 27170 4087 27240 4305
rect 27295 4268 27487 4273
rect 27295 4227 27306 4268
rect 27296 4165 27306 4227
rect 27295 4124 27306 4165
rect 27476 4227 27487 4268
rect 27476 4165 27486 4227
rect 27476 4124 27487 4165
rect 27295 4119 27487 4124
rect 27542 4087 27612 4305
rect 27667 4268 27859 4273
rect 27667 4227 27678 4268
rect 27668 4165 27678 4227
rect 27667 4124 27678 4165
rect 27848 4227 27859 4268
rect 27848 4165 27858 4227
rect 27848 4124 27859 4165
rect 27667 4119 27859 4124
rect 27914 4087 27984 4305
rect 28039 4268 28231 4273
rect 28039 4227 28050 4268
rect 28040 4165 28050 4227
rect 28039 4124 28050 4165
rect 28220 4227 28231 4268
rect 28220 4165 28230 4227
rect 28220 4124 28231 4165
rect 28039 4119 28231 4124
rect 28286 4087 28356 4305
rect 28411 4268 28603 4273
rect 28411 4227 28422 4268
rect 28412 4165 28422 4227
rect 28411 4124 28422 4165
rect 28592 4227 28603 4268
rect 28592 4165 28602 4227
rect 28592 4124 28603 4165
rect 28411 4119 28603 4124
rect 28658 4087 28728 4305
rect 28783 4268 28975 4273
rect 28783 4227 28794 4268
rect 28784 4165 28794 4227
rect 28783 4124 28794 4165
rect 28964 4227 28975 4268
rect 28964 4165 28974 4227
rect 28964 4124 28975 4165
rect 28783 4119 28975 4124
rect 29006 4087 29080 4305
rect 20122 4075 20217 4087
rect 20122 3899 20177 4075
rect 20211 3899 20217 4075
rect 20122 3887 20217 3899
rect 20429 4075 20589 4087
rect 20429 3899 20435 4075
rect 20469 3899 20549 4075
rect 20583 3899 20589 4075
rect 20429 3887 20589 3899
rect 20801 4075 20961 4087
rect 20801 3899 20807 4075
rect 20841 3899 20921 4075
rect 20955 3899 20961 4075
rect 20801 3887 20961 3899
rect 21173 4075 21333 4087
rect 21173 3899 21179 4075
rect 21213 3899 21293 4075
rect 21327 3899 21333 4075
rect 21173 3887 21333 3899
rect 21545 4075 21705 4087
rect 21545 3899 21551 4075
rect 21585 3899 21665 4075
rect 21699 3899 21705 4075
rect 21545 3887 21705 3899
rect 21917 4075 22077 4087
rect 21917 3899 21923 4075
rect 21957 3899 22037 4075
rect 22071 3899 22077 4075
rect 21917 3887 22077 3899
rect 22289 4075 22449 4087
rect 22289 3899 22295 4075
rect 22329 3899 22409 4075
rect 22443 3899 22449 4075
rect 22289 3887 22449 3899
rect 22661 4075 22821 4087
rect 22661 3899 22667 4075
rect 22701 3899 22781 4075
rect 22815 3899 22821 4075
rect 22661 3887 22821 3899
rect 23033 4075 23193 4087
rect 23033 3899 23039 4075
rect 23073 3899 23153 4075
rect 23187 3899 23193 4075
rect 23033 3887 23193 3899
rect 23405 4075 23565 4087
rect 23405 3899 23411 4075
rect 23445 3899 23525 4075
rect 23559 3899 23565 4075
rect 23405 3887 23565 3899
rect 23777 4075 23937 4087
rect 23777 3899 23783 4075
rect 23817 3899 23897 4075
rect 23931 3899 23937 4075
rect 23777 3887 23937 3899
rect 24149 4075 24309 4087
rect 24149 3899 24155 4075
rect 24189 3899 24269 4075
rect 24303 3899 24309 4075
rect 24149 3887 24309 3899
rect 24521 4075 24681 4087
rect 24521 3899 24527 4075
rect 24561 3899 24641 4075
rect 24675 3899 24681 4075
rect 24521 3887 24681 3899
rect 24893 4075 25053 4087
rect 24893 3899 24899 4075
rect 24933 3899 25013 4075
rect 25047 3899 25053 4075
rect 24893 3887 25053 3899
rect 25265 4075 25425 4087
rect 25265 3899 25271 4075
rect 25305 3899 25385 4075
rect 25419 3899 25425 4075
rect 25265 3887 25425 3899
rect 25637 4075 25797 4087
rect 25637 3899 25643 4075
rect 25677 3899 25757 4075
rect 25791 3899 25797 4075
rect 25637 3887 25797 3899
rect 26009 4075 26169 4087
rect 26009 3899 26015 4075
rect 26049 3899 26129 4075
rect 26163 3899 26169 4075
rect 26009 3887 26169 3899
rect 26381 4075 26541 4087
rect 26381 3899 26387 4075
rect 26421 3899 26501 4075
rect 26535 3899 26541 4075
rect 26381 3887 26541 3899
rect 26753 4075 26913 4087
rect 26753 3899 26759 4075
rect 26793 3899 26873 4075
rect 26907 3899 26913 4075
rect 26753 3887 26913 3899
rect 27125 4075 27285 4087
rect 27125 3899 27131 4075
rect 27165 3899 27245 4075
rect 27279 3899 27285 4075
rect 27125 3887 27285 3899
rect 27497 4075 27657 4087
rect 27497 3899 27503 4075
rect 27537 3899 27617 4075
rect 27651 3899 27657 4075
rect 27497 3887 27657 3899
rect 27869 4075 28029 4087
rect 27869 3899 27875 4075
rect 27909 3899 27989 4075
rect 28023 3899 28029 4075
rect 27869 3887 28029 3899
rect 28241 4075 28401 4087
rect 28241 3899 28247 4075
rect 28281 3899 28361 4075
rect 28395 3899 28401 4075
rect 28241 3887 28401 3899
rect 28613 4075 28773 4087
rect 28613 3899 28619 4075
rect 28653 3899 28733 4075
rect 28767 3899 28773 4075
rect 28613 3887 28773 3899
rect 28985 4075 29080 4087
rect 28985 3899 28991 4075
rect 29025 3899 29080 4075
rect 28985 3887 29080 3899
rect 20122 3669 20196 3887
rect 20474 3856 20544 3887
rect 20226 3850 20792 3856
rect 20226 3706 20238 3850
rect 20408 3706 20610 3850
rect 20780 3706 20792 3850
rect 20226 3700 20792 3706
rect 20474 3669 20544 3700
rect 20846 3669 20916 3887
rect 20971 3850 21163 3855
rect 20971 3809 20982 3850
rect 20972 3747 20982 3809
rect 20971 3706 20982 3747
rect 21152 3809 21163 3850
rect 21152 3747 21162 3809
rect 21152 3706 21163 3747
rect 20971 3701 21163 3706
rect 21218 3669 21288 3887
rect 21343 3850 21535 3855
rect 21343 3809 21354 3850
rect 21344 3747 21354 3809
rect 21343 3706 21354 3747
rect 21524 3809 21535 3850
rect 21524 3747 21534 3809
rect 21524 3706 21535 3747
rect 21343 3701 21535 3706
rect 21590 3669 21660 3887
rect 21715 3850 21907 3855
rect 21715 3809 21726 3850
rect 21716 3747 21726 3809
rect 21715 3706 21726 3747
rect 21896 3809 21907 3850
rect 21896 3747 21906 3809
rect 21896 3706 21907 3747
rect 21715 3701 21907 3706
rect 21962 3669 22032 3887
rect 22087 3850 22279 3855
rect 22087 3809 22098 3850
rect 22088 3747 22098 3809
rect 22087 3706 22098 3747
rect 22268 3809 22279 3850
rect 22268 3747 22278 3809
rect 22268 3706 22279 3747
rect 22087 3701 22279 3706
rect 22334 3669 22404 3887
rect 22706 3856 22776 3887
rect 22458 3850 23024 3856
rect 22458 3706 22470 3850
rect 22640 3706 22842 3850
rect 23012 3706 23024 3850
rect 22458 3700 23024 3706
rect 22706 3669 22776 3700
rect 23078 3669 23148 3887
rect 23203 3850 23395 3855
rect 23203 3809 23214 3850
rect 23204 3747 23214 3809
rect 23203 3706 23214 3747
rect 23384 3809 23395 3850
rect 23384 3747 23394 3809
rect 23384 3706 23395 3747
rect 23203 3701 23395 3706
rect 23450 3669 23520 3887
rect 23575 3850 23767 3855
rect 23575 3809 23586 3850
rect 23576 3747 23586 3809
rect 23575 3706 23586 3747
rect 23756 3809 23767 3850
rect 23756 3747 23766 3809
rect 23756 3706 23767 3747
rect 23575 3701 23767 3706
rect 23822 3669 23892 3887
rect 23947 3850 24139 3855
rect 23947 3809 23958 3850
rect 23948 3747 23958 3809
rect 23947 3706 23958 3747
rect 24128 3809 24139 3850
rect 24128 3747 24138 3809
rect 24128 3706 24139 3747
rect 23947 3701 24139 3706
rect 24194 3669 24264 3887
rect 24319 3850 24511 3855
rect 24319 3809 24330 3850
rect 24320 3747 24330 3809
rect 24319 3706 24330 3747
rect 24500 3809 24511 3850
rect 24500 3747 24510 3809
rect 24500 3706 24511 3747
rect 24319 3701 24511 3706
rect 24566 3669 24636 3887
rect 24691 3850 24883 3855
rect 24691 3809 24702 3850
rect 24692 3747 24702 3809
rect 24691 3706 24702 3747
rect 24872 3809 24883 3850
rect 24872 3747 24882 3809
rect 24872 3706 24883 3747
rect 24691 3701 24883 3706
rect 24938 3669 25008 3887
rect 25063 3850 25255 3855
rect 25063 3809 25074 3850
rect 25064 3747 25074 3809
rect 25063 3706 25074 3747
rect 25244 3809 25255 3850
rect 25244 3747 25254 3809
rect 25244 3706 25255 3747
rect 25063 3701 25255 3706
rect 25310 3669 25380 3887
rect 25435 3850 25627 3855
rect 25435 3809 25446 3850
rect 25436 3747 25446 3809
rect 25435 3706 25446 3747
rect 25616 3809 25627 3850
rect 25616 3747 25626 3809
rect 25616 3706 25627 3747
rect 25435 3701 25627 3706
rect 25682 3669 25752 3887
rect 25807 3850 25999 3855
rect 25807 3809 25818 3850
rect 25808 3747 25818 3809
rect 25807 3706 25818 3747
rect 25988 3809 25999 3850
rect 25988 3747 25998 3809
rect 25988 3706 25999 3747
rect 25807 3701 25999 3706
rect 26054 3669 26124 3887
rect 26179 3850 26371 3855
rect 26179 3809 26190 3850
rect 26180 3747 26190 3809
rect 26179 3706 26190 3747
rect 26360 3809 26371 3850
rect 26360 3747 26370 3809
rect 26360 3706 26371 3747
rect 26179 3701 26371 3706
rect 26426 3669 26496 3887
rect 26551 3850 26743 3855
rect 26551 3809 26562 3850
rect 26552 3747 26562 3809
rect 26551 3706 26562 3747
rect 26732 3809 26743 3850
rect 26732 3747 26742 3809
rect 26732 3706 26743 3747
rect 26551 3701 26743 3706
rect 26798 3669 26868 3887
rect 26923 3850 27115 3855
rect 26923 3809 26934 3850
rect 26924 3747 26934 3809
rect 26923 3706 26934 3747
rect 27104 3809 27115 3850
rect 27104 3747 27114 3809
rect 27104 3706 27115 3747
rect 26923 3701 27115 3706
rect 27170 3669 27240 3887
rect 27295 3850 27487 3855
rect 27295 3809 27306 3850
rect 27296 3747 27306 3809
rect 27295 3706 27306 3747
rect 27476 3809 27487 3850
rect 27476 3747 27486 3809
rect 27476 3706 27487 3747
rect 27295 3701 27487 3706
rect 27542 3669 27612 3887
rect 27667 3850 27859 3855
rect 27667 3809 27678 3850
rect 27668 3747 27678 3809
rect 27667 3706 27678 3747
rect 27848 3809 27859 3850
rect 27848 3747 27858 3809
rect 27848 3706 27859 3747
rect 27667 3701 27859 3706
rect 27914 3669 27984 3887
rect 28039 3850 28231 3855
rect 28039 3809 28050 3850
rect 28040 3747 28050 3809
rect 28039 3706 28050 3747
rect 28220 3809 28231 3850
rect 28220 3747 28230 3809
rect 28220 3706 28231 3747
rect 28039 3701 28231 3706
rect 28286 3669 28356 3887
rect 28411 3850 28603 3855
rect 28411 3809 28422 3850
rect 28412 3747 28422 3809
rect 28411 3706 28422 3747
rect 28592 3809 28603 3850
rect 28592 3747 28602 3809
rect 28592 3706 28603 3747
rect 28411 3701 28603 3706
rect 28658 3669 28728 3887
rect 28783 3850 28975 3855
rect 28783 3809 28794 3850
rect 28784 3747 28794 3809
rect 28783 3706 28794 3747
rect 28964 3809 28975 3850
rect 28964 3747 28974 3809
rect 28964 3706 28975 3747
rect 28783 3701 28975 3706
rect 29006 3669 29080 3887
rect 20122 3657 20217 3669
rect 20122 3481 20177 3657
rect 20211 3481 20217 3657
rect 20122 3469 20217 3481
rect 20429 3657 20589 3669
rect 20429 3481 20435 3657
rect 20469 3481 20549 3657
rect 20583 3481 20589 3657
rect 20429 3469 20589 3481
rect 20801 3657 20961 3669
rect 20801 3481 20807 3657
rect 20841 3481 20921 3657
rect 20955 3481 20961 3657
rect 20801 3469 20961 3481
rect 21173 3657 21333 3669
rect 21173 3481 21179 3657
rect 21213 3481 21293 3657
rect 21327 3481 21333 3657
rect 21173 3469 21333 3481
rect 21545 3657 21705 3669
rect 21545 3481 21551 3657
rect 21585 3481 21665 3657
rect 21699 3481 21705 3657
rect 21545 3469 21705 3481
rect 21917 3657 22077 3669
rect 21917 3481 21923 3657
rect 21957 3481 22037 3657
rect 22071 3481 22077 3657
rect 21917 3469 22077 3481
rect 22289 3657 22449 3669
rect 22289 3481 22295 3657
rect 22329 3481 22409 3657
rect 22443 3481 22449 3657
rect 22289 3469 22449 3481
rect 22661 3657 22821 3669
rect 22661 3481 22667 3657
rect 22701 3481 22781 3657
rect 22815 3481 22821 3657
rect 22661 3469 22821 3481
rect 23033 3657 23193 3669
rect 23033 3481 23039 3657
rect 23073 3481 23153 3657
rect 23187 3481 23193 3657
rect 23033 3469 23193 3481
rect 23405 3657 23565 3669
rect 23405 3481 23411 3657
rect 23445 3481 23525 3657
rect 23559 3481 23565 3657
rect 23405 3469 23565 3481
rect 23777 3657 23937 3669
rect 23777 3481 23783 3657
rect 23817 3481 23897 3657
rect 23931 3481 23937 3657
rect 23777 3469 23937 3481
rect 24149 3657 24309 3669
rect 24149 3481 24155 3657
rect 24189 3481 24269 3657
rect 24303 3481 24309 3657
rect 24149 3469 24309 3481
rect 24521 3657 24681 3669
rect 24521 3481 24527 3657
rect 24561 3481 24641 3657
rect 24675 3481 24681 3657
rect 24521 3469 24681 3481
rect 24893 3657 25053 3669
rect 24893 3481 24899 3657
rect 24933 3481 25013 3657
rect 25047 3481 25053 3657
rect 24893 3469 25053 3481
rect 25265 3657 25425 3669
rect 25265 3481 25271 3657
rect 25305 3481 25385 3657
rect 25419 3481 25425 3657
rect 25265 3469 25425 3481
rect 25637 3657 25797 3669
rect 25637 3481 25643 3657
rect 25677 3481 25757 3657
rect 25791 3481 25797 3657
rect 25637 3469 25797 3481
rect 26009 3657 26169 3669
rect 26009 3481 26015 3657
rect 26049 3481 26129 3657
rect 26163 3481 26169 3657
rect 26009 3469 26169 3481
rect 26381 3657 26541 3669
rect 26381 3481 26387 3657
rect 26421 3481 26501 3657
rect 26535 3481 26541 3657
rect 26381 3469 26541 3481
rect 26753 3657 26913 3669
rect 26753 3481 26759 3657
rect 26793 3481 26873 3657
rect 26907 3481 26913 3657
rect 26753 3469 26913 3481
rect 27125 3657 27285 3669
rect 27125 3481 27131 3657
rect 27165 3481 27245 3657
rect 27279 3481 27285 3657
rect 27125 3469 27285 3481
rect 27497 3657 27657 3669
rect 27497 3481 27503 3657
rect 27537 3481 27617 3657
rect 27651 3481 27657 3657
rect 27497 3469 27657 3481
rect 27869 3657 28029 3669
rect 27869 3481 27875 3657
rect 27909 3481 27989 3657
rect 28023 3481 28029 3657
rect 27869 3469 28029 3481
rect 28241 3657 28401 3669
rect 28241 3481 28247 3657
rect 28281 3481 28361 3657
rect 28395 3481 28401 3657
rect 28241 3469 28401 3481
rect 28613 3657 28773 3669
rect 28613 3481 28619 3657
rect 28653 3481 28733 3657
rect 28767 3481 28773 3657
rect 28613 3469 28773 3481
rect 28985 3657 29080 3669
rect 28985 3481 28991 3657
rect 29025 3481 29080 3657
rect 28985 3469 29080 3481
rect 20122 3251 20196 3469
rect 20474 3438 20544 3469
rect 20226 3432 20792 3438
rect 20226 3288 20238 3432
rect 20408 3288 20610 3432
rect 20780 3288 20792 3432
rect 20226 3282 20792 3288
rect 20474 3251 20544 3282
rect 20846 3251 20916 3469
rect 20971 3432 21163 3437
rect 20971 3391 20982 3432
rect 20972 3329 20982 3391
rect 20971 3288 20982 3329
rect 21152 3391 21163 3432
rect 21152 3329 21162 3391
rect 21152 3288 21163 3329
rect 20971 3283 21163 3288
rect 21218 3251 21288 3469
rect 21343 3432 21535 3437
rect 21343 3391 21354 3432
rect 21344 3329 21354 3391
rect 21343 3288 21354 3329
rect 21524 3391 21535 3432
rect 21524 3329 21534 3391
rect 21524 3288 21535 3329
rect 21343 3283 21535 3288
rect 21590 3251 21660 3469
rect 21715 3432 21907 3437
rect 21715 3391 21726 3432
rect 21716 3329 21726 3391
rect 21715 3288 21726 3329
rect 21896 3391 21907 3432
rect 21896 3329 21906 3391
rect 21896 3288 21907 3329
rect 21715 3283 21907 3288
rect 21962 3251 22032 3469
rect 22087 3432 22279 3437
rect 22087 3391 22098 3432
rect 22088 3329 22098 3391
rect 22087 3288 22098 3329
rect 22268 3391 22279 3432
rect 22268 3329 22278 3391
rect 22268 3288 22279 3329
rect 22087 3283 22279 3288
rect 22334 3251 22404 3469
rect 22706 3438 22776 3469
rect 22458 3432 23024 3438
rect 22458 3288 22470 3432
rect 22640 3288 22842 3432
rect 23012 3288 23024 3432
rect 22458 3282 23024 3288
rect 22706 3251 22776 3282
rect 23078 3251 23148 3469
rect 23203 3432 23395 3437
rect 23203 3391 23214 3432
rect 23204 3329 23214 3391
rect 23203 3288 23214 3329
rect 23384 3391 23395 3432
rect 23384 3329 23394 3391
rect 23384 3288 23395 3329
rect 23203 3283 23395 3288
rect 23450 3251 23520 3469
rect 23575 3432 23767 3437
rect 23575 3391 23586 3432
rect 23576 3329 23586 3391
rect 23575 3288 23586 3329
rect 23756 3391 23767 3432
rect 23756 3329 23766 3391
rect 23756 3288 23767 3329
rect 23575 3283 23767 3288
rect 23822 3251 23892 3469
rect 23947 3432 24139 3437
rect 23947 3391 23958 3432
rect 23948 3329 23958 3391
rect 23947 3288 23958 3329
rect 24128 3391 24139 3432
rect 24128 3329 24138 3391
rect 24128 3288 24139 3329
rect 23947 3283 24139 3288
rect 24194 3251 24264 3469
rect 24319 3432 24511 3437
rect 24319 3391 24330 3432
rect 24320 3329 24330 3391
rect 24319 3288 24330 3329
rect 24500 3391 24511 3432
rect 24500 3329 24510 3391
rect 24500 3288 24511 3329
rect 24319 3283 24511 3288
rect 24566 3251 24636 3469
rect 24691 3432 24883 3437
rect 24691 3391 24702 3432
rect 24692 3329 24702 3391
rect 24691 3288 24702 3329
rect 24872 3391 24883 3432
rect 24872 3329 24882 3391
rect 24872 3288 24883 3329
rect 24691 3283 24883 3288
rect 24938 3251 25008 3469
rect 25063 3432 25255 3437
rect 25063 3391 25074 3432
rect 25064 3329 25074 3391
rect 25063 3288 25074 3329
rect 25244 3391 25255 3432
rect 25244 3329 25254 3391
rect 25244 3288 25255 3329
rect 25063 3283 25255 3288
rect 25310 3251 25380 3469
rect 25435 3432 25627 3437
rect 25435 3391 25446 3432
rect 25436 3329 25446 3391
rect 25435 3288 25446 3329
rect 25616 3391 25627 3432
rect 25616 3329 25626 3391
rect 25616 3288 25627 3329
rect 25435 3283 25627 3288
rect 25682 3251 25752 3469
rect 25807 3432 25999 3437
rect 25807 3391 25818 3432
rect 25808 3329 25818 3391
rect 25807 3288 25818 3329
rect 25988 3391 25999 3432
rect 25988 3329 25998 3391
rect 25988 3288 25999 3329
rect 25807 3283 25999 3288
rect 26054 3251 26124 3469
rect 26179 3432 26371 3437
rect 26179 3391 26190 3432
rect 26180 3329 26190 3391
rect 26179 3288 26190 3329
rect 26360 3391 26371 3432
rect 26360 3329 26370 3391
rect 26360 3288 26371 3329
rect 26179 3283 26371 3288
rect 26426 3251 26496 3469
rect 26551 3432 26743 3437
rect 26551 3391 26562 3432
rect 26552 3329 26562 3391
rect 26551 3288 26562 3329
rect 26732 3391 26743 3432
rect 26732 3329 26742 3391
rect 26732 3288 26743 3329
rect 26551 3283 26743 3288
rect 26798 3251 26868 3469
rect 26923 3432 27115 3437
rect 26923 3391 26934 3432
rect 26924 3329 26934 3391
rect 26923 3288 26934 3329
rect 27104 3391 27115 3432
rect 27104 3329 27114 3391
rect 27104 3288 27115 3329
rect 26923 3283 27115 3288
rect 27170 3251 27240 3469
rect 27295 3432 27487 3437
rect 27295 3391 27306 3432
rect 27296 3329 27306 3391
rect 27295 3288 27306 3329
rect 27476 3391 27487 3432
rect 27476 3329 27486 3391
rect 27476 3288 27487 3329
rect 27295 3283 27487 3288
rect 27542 3251 27612 3469
rect 27667 3432 27859 3437
rect 27667 3391 27678 3432
rect 27668 3329 27678 3391
rect 27667 3288 27678 3329
rect 27848 3391 27859 3432
rect 27848 3329 27858 3391
rect 27848 3288 27859 3329
rect 27667 3283 27859 3288
rect 27914 3251 27984 3469
rect 28039 3432 28231 3437
rect 28039 3391 28050 3432
rect 28040 3329 28050 3391
rect 28039 3288 28050 3329
rect 28220 3391 28231 3432
rect 28220 3329 28230 3391
rect 28220 3288 28231 3329
rect 28039 3283 28231 3288
rect 28286 3251 28356 3469
rect 28411 3432 28603 3437
rect 28411 3391 28422 3432
rect 28412 3329 28422 3391
rect 28411 3288 28422 3329
rect 28592 3391 28603 3432
rect 28592 3329 28602 3391
rect 28592 3288 28603 3329
rect 28411 3283 28603 3288
rect 28658 3251 28728 3469
rect 28783 3432 28975 3437
rect 28783 3391 28794 3432
rect 28784 3329 28794 3391
rect 28783 3288 28794 3329
rect 28964 3391 28975 3432
rect 28964 3329 28974 3391
rect 28964 3288 28975 3329
rect 28783 3283 28975 3288
rect 29006 3251 29080 3469
rect 20122 3239 20217 3251
rect 20122 3063 20177 3239
rect 20211 3063 20217 3239
rect 20122 3051 20217 3063
rect 20429 3239 20589 3251
rect 20429 3063 20435 3239
rect 20469 3063 20549 3239
rect 20583 3063 20589 3239
rect 20429 3051 20589 3063
rect 20801 3239 20961 3251
rect 20801 3063 20807 3239
rect 20841 3063 20921 3239
rect 20955 3063 20961 3239
rect 20801 3051 20961 3063
rect 21173 3239 21333 3251
rect 21173 3063 21179 3239
rect 21213 3063 21293 3239
rect 21327 3063 21333 3239
rect 21173 3051 21333 3063
rect 21545 3239 21705 3251
rect 21545 3063 21551 3239
rect 21585 3063 21665 3239
rect 21699 3063 21705 3239
rect 21545 3051 21705 3063
rect 21917 3239 22077 3251
rect 21917 3063 21923 3239
rect 21957 3063 22037 3239
rect 22071 3063 22077 3239
rect 21917 3051 22077 3063
rect 22289 3239 22449 3251
rect 22289 3063 22295 3239
rect 22329 3063 22409 3239
rect 22443 3063 22449 3239
rect 22289 3051 22449 3063
rect 22661 3239 22821 3251
rect 22661 3063 22667 3239
rect 22701 3063 22781 3239
rect 22815 3063 22821 3239
rect 22661 3051 22821 3063
rect 23033 3239 23193 3251
rect 23033 3063 23039 3239
rect 23073 3063 23153 3239
rect 23187 3063 23193 3239
rect 23033 3051 23193 3063
rect 23405 3239 23565 3251
rect 23405 3063 23411 3239
rect 23445 3063 23525 3239
rect 23559 3063 23565 3239
rect 23405 3051 23565 3063
rect 23777 3239 23937 3251
rect 23777 3063 23783 3239
rect 23817 3063 23897 3239
rect 23931 3063 23937 3239
rect 23777 3051 23937 3063
rect 24149 3239 24309 3251
rect 24149 3063 24155 3239
rect 24189 3063 24269 3239
rect 24303 3063 24309 3239
rect 24149 3051 24309 3063
rect 24521 3239 24681 3251
rect 24521 3063 24527 3239
rect 24561 3063 24641 3239
rect 24675 3063 24681 3239
rect 24521 3051 24681 3063
rect 24893 3239 25053 3251
rect 24893 3063 24899 3239
rect 24933 3063 25013 3239
rect 25047 3063 25053 3239
rect 24893 3051 25053 3063
rect 25265 3239 25425 3251
rect 25265 3063 25271 3239
rect 25305 3063 25385 3239
rect 25419 3063 25425 3239
rect 25265 3051 25425 3063
rect 25637 3239 25797 3251
rect 25637 3063 25643 3239
rect 25677 3063 25757 3239
rect 25791 3063 25797 3239
rect 25637 3051 25797 3063
rect 26009 3239 26169 3251
rect 26009 3063 26015 3239
rect 26049 3063 26129 3239
rect 26163 3063 26169 3239
rect 26009 3051 26169 3063
rect 26381 3239 26541 3251
rect 26381 3063 26387 3239
rect 26421 3063 26501 3239
rect 26535 3063 26541 3239
rect 26381 3051 26541 3063
rect 26753 3239 26913 3251
rect 26753 3063 26759 3239
rect 26793 3063 26873 3239
rect 26907 3063 26913 3239
rect 26753 3051 26913 3063
rect 27125 3239 27285 3251
rect 27125 3063 27131 3239
rect 27165 3063 27245 3239
rect 27279 3063 27285 3239
rect 27125 3051 27285 3063
rect 27497 3239 27657 3251
rect 27497 3063 27503 3239
rect 27537 3063 27617 3239
rect 27651 3063 27657 3239
rect 27497 3051 27657 3063
rect 27869 3239 28029 3251
rect 27869 3063 27875 3239
rect 27909 3063 27989 3239
rect 28023 3063 28029 3239
rect 27869 3051 28029 3063
rect 28241 3239 28401 3251
rect 28241 3063 28247 3239
rect 28281 3063 28361 3239
rect 28395 3063 28401 3239
rect 28241 3051 28401 3063
rect 28613 3239 28773 3251
rect 28613 3063 28619 3239
rect 28653 3063 28733 3239
rect 28767 3063 28773 3239
rect 28613 3051 28773 3063
rect 28985 3239 29080 3251
rect 28985 3063 28991 3239
rect 29025 3063 29080 3239
rect 28985 3051 29080 3063
rect 20122 2928 20196 3051
rect 20228 3019 20238 3024
rect 20227 3014 20238 3019
rect 20226 2968 20238 3014
rect 20408 3019 20418 3024
rect 20408 3014 20419 3019
rect 20474 3014 20544 3051
rect 20846 3050 20916 3051
rect 21218 3050 21288 3051
rect 21590 3050 21660 3051
rect 21962 3050 22032 3051
rect 22334 3050 22404 3051
rect 20600 3019 20610 3024
rect 20599 3014 20610 3019
rect 20408 2968 20610 3014
rect 20780 3019 20790 3024
rect 20780 3014 20791 3019
rect 20780 2968 20792 3014
rect 20226 2956 20792 2968
rect 20852 2936 20910 3050
rect 20972 3019 20982 3024
rect 20971 2973 20982 3019
rect 21152 3019 21162 3024
rect 21344 3019 21354 3024
rect 20972 2968 20982 2973
rect 21152 2973 21163 3019
rect 21343 2973 21354 3019
rect 21524 3019 21534 3024
rect 21152 2968 21162 2973
rect 21344 2968 21354 2973
rect 21524 2973 21535 3019
rect 21524 2968 21534 2973
rect 21596 2936 21654 3050
rect 21716 3019 21726 3024
rect 21715 2973 21726 3019
rect 21896 3019 21906 3024
rect 22088 3019 22098 3024
rect 21716 2968 21726 2973
rect 21896 2973 21907 3019
rect 22087 2973 22098 3019
rect 22268 3019 22278 3024
rect 21896 2968 21906 2973
rect 22088 2968 22098 2973
rect 22268 2973 22279 3019
rect 22268 2968 22278 2973
rect 22340 2936 22398 3050
rect 22460 3019 22470 3024
rect 22459 3014 22470 3019
rect 22458 2968 22470 3014
rect 22640 3019 22650 3024
rect 22640 3014 22651 3019
rect 22706 3014 22776 3051
rect 23078 3050 23148 3051
rect 23450 3050 23520 3051
rect 23822 3050 23892 3051
rect 24194 3050 24264 3051
rect 24566 3050 24636 3051
rect 24938 3050 25008 3051
rect 25310 3050 25380 3051
rect 25682 3050 25752 3051
rect 26054 3050 26124 3051
rect 26426 3050 26496 3051
rect 26798 3050 26868 3051
rect 27170 3050 27240 3051
rect 27542 3050 27612 3051
rect 27914 3050 27984 3051
rect 28286 3050 28356 3051
rect 28658 3050 28728 3051
rect 22832 3019 22842 3024
rect 22831 3014 22842 3019
rect 22640 2968 22842 3014
rect 23012 3019 23022 3024
rect 23012 3014 23023 3019
rect 23012 2968 23024 3014
rect 22458 2956 23024 2968
rect 23084 2936 23142 3050
rect 23204 3019 23214 3024
rect 23203 2973 23214 3019
rect 23384 3019 23394 3024
rect 23576 3019 23586 3024
rect 23204 2968 23214 2973
rect 23384 2973 23395 3019
rect 23575 2973 23586 3019
rect 23756 3019 23766 3024
rect 23384 2968 23394 2973
rect 23576 2968 23586 2973
rect 23756 2973 23767 3019
rect 23756 2968 23766 2973
rect 23828 2936 23886 3050
rect 23948 3019 23958 3024
rect 23947 2973 23958 3019
rect 24128 3019 24138 3024
rect 24320 3019 24330 3024
rect 23948 2968 23958 2973
rect 24128 2973 24139 3019
rect 24319 2973 24330 3019
rect 24500 3019 24510 3024
rect 24128 2968 24138 2973
rect 24320 2968 24330 2973
rect 24500 2973 24511 3019
rect 24500 2968 24510 2973
rect 24572 2936 24630 3050
rect 24692 3019 24702 3024
rect 24691 2973 24702 3019
rect 24872 3019 24882 3024
rect 25064 3019 25074 3024
rect 24692 2968 24702 2973
rect 24872 2973 24883 3019
rect 25063 2973 25074 3019
rect 25244 3019 25254 3024
rect 24872 2968 24882 2973
rect 25064 2968 25074 2973
rect 25244 2973 25255 3019
rect 25244 2968 25254 2973
rect 25316 2936 25374 3050
rect 25436 3019 25446 3024
rect 25435 2973 25446 3019
rect 25616 3019 25626 3024
rect 25808 3019 25818 3024
rect 25436 2968 25446 2973
rect 25616 2973 25627 3019
rect 25807 2973 25818 3019
rect 25988 3019 25998 3024
rect 25616 2968 25626 2973
rect 25808 2968 25818 2973
rect 25988 2973 25999 3019
rect 25988 2968 25998 2973
rect 26060 2936 26118 3050
rect 26180 3019 26190 3024
rect 26179 2973 26190 3019
rect 26360 3019 26370 3024
rect 26552 3019 26562 3024
rect 26180 2968 26190 2973
rect 26360 2973 26371 3019
rect 26551 2973 26562 3019
rect 26732 3019 26742 3024
rect 26360 2968 26370 2973
rect 26552 2968 26562 2973
rect 26732 2973 26743 3019
rect 26732 2968 26742 2973
rect 26804 2936 26862 3050
rect 26924 3019 26934 3024
rect 26923 2973 26934 3019
rect 27104 3019 27114 3024
rect 27296 3019 27306 3024
rect 26924 2968 26934 2973
rect 27104 2973 27115 3019
rect 27295 2973 27306 3019
rect 27476 3019 27486 3024
rect 27104 2968 27114 2973
rect 27296 2968 27306 2973
rect 27476 2973 27487 3019
rect 27476 2968 27486 2973
rect 27548 2936 27606 3050
rect 27668 3019 27678 3024
rect 27667 2973 27678 3019
rect 27848 3019 27858 3024
rect 28040 3019 28050 3024
rect 27668 2968 27678 2973
rect 27848 2973 27859 3019
rect 28039 2973 28050 3019
rect 28220 3019 28230 3024
rect 27848 2968 27858 2973
rect 28040 2968 28050 2973
rect 28220 2973 28231 3019
rect 28220 2968 28230 2973
rect 28292 2936 28350 3050
rect 28412 3019 28422 3024
rect 28411 2973 28422 3019
rect 28592 3019 28602 3024
rect 28784 3019 28794 3024
rect 28412 2968 28422 2973
rect 28592 2973 28603 3019
rect 28783 2973 28794 3019
rect 28964 3019 28974 3024
rect 28592 2968 28602 2973
rect 28784 2968 28794 2973
rect 28964 2973 28975 3019
rect 28964 2968 28974 2973
rect 20834 2930 20928 2936
rect 20122 2922 20260 2928
rect 20122 2852 20178 2922
rect 20248 2852 20260 2922
rect 20834 2860 20846 2930
rect 20916 2860 20928 2930
rect 20834 2854 20928 2860
rect 21578 2930 21672 2936
rect 21578 2860 21590 2930
rect 21660 2860 21672 2930
rect 21578 2854 21672 2860
rect 22322 2930 22416 2936
rect 22322 2860 22334 2930
rect 22404 2860 22416 2930
rect 22322 2854 22416 2860
rect 23066 2930 23160 2936
rect 23066 2860 23078 2930
rect 23148 2860 23160 2930
rect 23066 2854 23160 2860
rect 23810 2930 23904 2936
rect 23810 2860 23822 2930
rect 23892 2860 23904 2930
rect 23810 2854 23904 2860
rect 24554 2930 24648 2936
rect 24554 2860 24566 2930
rect 24636 2860 24648 2930
rect 24554 2854 24648 2860
rect 25298 2930 25392 2936
rect 25298 2860 25310 2930
rect 25380 2860 25392 2930
rect 25298 2854 25392 2860
rect 26042 2930 26136 2936
rect 26042 2860 26054 2930
rect 26124 2860 26136 2930
rect 26042 2854 26136 2860
rect 26786 2930 26880 2936
rect 26786 2860 26798 2930
rect 26868 2860 26880 2930
rect 26786 2854 26880 2860
rect 27530 2930 27624 2936
rect 27530 2860 27542 2930
rect 27612 2860 27624 2930
rect 27530 2854 27624 2860
rect 28274 2930 28368 2936
rect 29006 2932 29080 3051
rect 28274 2860 28286 2930
rect 28356 2860 28368 2930
rect 28274 2854 28368 2860
rect 28936 2926 29080 2932
rect 28936 2856 28948 2926
rect 29018 2856 29080 2926
rect 20122 2846 20260 2852
rect 20122 2814 20196 2846
rect 20852 2814 20910 2854
rect 21596 2814 21654 2854
rect 22340 2814 22398 2854
rect 23084 2814 23142 2854
rect 23828 2814 23886 2854
rect 24572 2814 24630 2854
rect 25316 2814 25374 2854
rect 26060 2814 26118 2854
rect 26804 2814 26862 2854
rect 27548 2814 27606 2854
rect 28292 2814 28350 2854
rect 28936 2850 29080 2856
rect 29006 2826 29080 2850
rect 29006 2814 29094 2826
rect 20048 2614 20058 2814
rect 20258 2614 20268 2814
rect 20772 2614 20782 2814
rect 20982 2614 20992 2814
rect 21516 2614 21526 2814
rect 21726 2614 21736 2814
rect 22260 2614 22270 2814
rect 22470 2614 22480 2814
rect 23004 2614 23014 2814
rect 23214 2614 23224 2814
rect 23748 2614 23758 2814
rect 23958 2614 23968 2814
rect 24492 2614 24502 2814
rect 24702 2614 24712 2814
rect 25236 2614 25246 2814
rect 25446 2614 25456 2814
rect 25980 2614 25990 2814
rect 26190 2614 26200 2814
rect 26724 2614 26734 2814
rect 26934 2614 26944 2814
rect 27468 2614 27478 2814
rect 27678 2614 27688 2814
rect 28212 2614 28222 2814
rect 28422 2614 28432 2814
rect 28956 2614 28966 2814
rect 29166 2614 29176 2814
<< via1 >>
rect 18920 11860 19120 12060
rect 19664 11860 19864 12060
rect 20408 11860 20608 12060
rect 21152 11860 21352 12060
rect 21896 11860 22096 12060
rect 22640 11860 22840 12060
rect 23384 11860 23584 12060
rect 24128 11860 24328 12060
rect 24500 11860 24700 12060
rect 25244 11860 25444 12060
rect 25988 11860 26188 12060
rect 26732 11860 26932 12060
rect 27476 11860 27676 12060
rect 28220 11860 28420 12060
rect 28964 11860 29164 12060
rect 29708 11860 29908 12060
rect 30452 11860 30652 12060
rect 18750 11659 18920 11672
rect 18750 11625 18751 11659
rect 18751 11625 18919 11659
rect 18919 11625 18920 11659
rect 18750 11612 18920 11625
rect 19122 11659 19292 11672
rect 19122 11625 19123 11659
rect 19123 11625 19291 11659
rect 19291 11625 19292 11659
rect 19122 11612 19292 11625
rect 19494 11659 19664 11672
rect 19494 11625 19495 11659
rect 19495 11625 19663 11659
rect 19663 11625 19664 11659
rect 19494 11612 19664 11625
rect 19866 11659 20036 11672
rect 19866 11625 19867 11659
rect 19867 11625 20035 11659
rect 20035 11625 20036 11659
rect 19866 11612 20036 11625
rect 20238 11659 20408 11672
rect 20238 11625 20239 11659
rect 20239 11625 20407 11659
rect 20407 11625 20408 11659
rect 20238 11612 20408 11625
rect 20610 11659 20780 11672
rect 20610 11625 20611 11659
rect 20611 11625 20779 11659
rect 20779 11625 20780 11659
rect 20610 11612 20780 11625
rect 20982 11659 21152 11672
rect 20982 11625 20983 11659
rect 20983 11625 21151 11659
rect 21151 11625 21152 11659
rect 20982 11612 21152 11625
rect 21354 11659 21524 11672
rect 21354 11625 21355 11659
rect 21355 11625 21523 11659
rect 21523 11625 21524 11659
rect 21354 11612 21524 11625
rect 21726 11659 21896 11672
rect 21726 11625 21727 11659
rect 21727 11625 21895 11659
rect 21895 11625 21896 11659
rect 21726 11612 21896 11625
rect 22098 11659 22268 11672
rect 22098 11625 22099 11659
rect 22099 11625 22267 11659
rect 22267 11625 22268 11659
rect 22098 11612 22268 11625
rect 22470 11659 22640 11672
rect 22470 11625 22471 11659
rect 22471 11625 22639 11659
rect 22639 11625 22640 11659
rect 22470 11612 22640 11625
rect 22842 11659 23012 11672
rect 22842 11625 22843 11659
rect 22843 11625 23011 11659
rect 23011 11625 23012 11659
rect 22842 11612 23012 11625
rect 23214 11659 23384 11672
rect 23214 11625 23215 11659
rect 23215 11625 23383 11659
rect 23383 11625 23384 11659
rect 23214 11612 23384 11625
rect 23586 11659 23756 11672
rect 23586 11625 23587 11659
rect 23587 11625 23755 11659
rect 23755 11625 23756 11659
rect 23586 11612 23756 11625
rect 23958 11659 24128 11672
rect 23958 11625 23959 11659
rect 23959 11625 24127 11659
rect 24127 11625 24128 11659
rect 23958 11612 24128 11625
rect 24330 11659 24500 11672
rect 24330 11625 24331 11659
rect 24331 11625 24499 11659
rect 24499 11625 24500 11659
rect 24330 11612 24500 11625
rect 18750 11131 18920 11132
rect 18750 11097 18751 11131
rect 18751 11097 18919 11131
rect 18919 11097 18920 11131
rect 18750 11023 18920 11097
rect 18750 10989 18751 11023
rect 18751 10989 18919 11023
rect 18919 10989 18920 11023
rect 18750 10988 18920 10989
rect 19122 11131 19292 11132
rect 19122 11097 19123 11131
rect 19123 11097 19291 11131
rect 19291 11097 19292 11131
rect 19122 11023 19292 11097
rect 19122 10989 19123 11023
rect 19123 10989 19291 11023
rect 19291 10989 19292 11023
rect 19122 10988 19292 10989
rect 19494 11131 19664 11132
rect 19494 11097 19495 11131
rect 19495 11097 19663 11131
rect 19663 11097 19664 11131
rect 19494 11023 19664 11097
rect 19494 10989 19495 11023
rect 19495 10989 19663 11023
rect 19663 10989 19664 11023
rect 19494 10988 19664 10989
rect 19866 11131 20036 11132
rect 19866 11097 19867 11131
rect 19867 11097 20035 11131
rect 20035 11097 20036 11131
rect 19866 11023 20036 11097
rect 19866 10989 19867 11023
rect 19867 10989 20035 11023
rect 20035 10989 20036 11023
rect 19866 10988 20036 10989
rect 20238 11131 20408 11132
rect 20238 11097 20239 11131
rect 20239 11097 20407 11131
rect 20407 11097 20408 11131
rect 20238 11023 20408 11097
rect 20238 10989 20239 11023
rect 20239 10989 20407 11023
rect 20407 10989 20408 11023
rect 20238 10988 20408 10989
rect 20610 11131 20780 11132
rect 20610 11097 20611 11131
rect 20611 11097 20779 11131
rect 20779 11097 20780 11131
rect 20610 11023 20780 11097
rect 20610 10989 20611 11023
rect 20611 10989 20779 11023
rect 20779 10989 20780 11023
rect 20610 10988 20780 10989
rect 20982 11131 21152 11132
rect 20982 11097 20983 11131
rect 20983 11097 21151 11131
rect 21151 11097 21152 11131
rect 20982 11023 21152 11097
rect 20982 10989 20983 11023
rect 20983 10989 21151 11023
rect 21151 10989 21152 11023
rect 20982 10988 21152 10989
rect 21354 11131 21524 11132
rect 21354 11097 21355 11131
rect 21355 11097 21523 11131
rect 21523 11097 21524 11131
rect 21354 11023 21524 11097
rect 21354 10989 21355 11023
rect 21355 10989 21523 11023
rect 21523 10989 21524 11023
rect 21354 10988 21524 10989
rect 21726 11131 21896 11132
rect 21726 11097 21727 11131
rect 21727 11097 21895 11131
rect 21895 11097 21896 11131
rect 21726 11023 21896 11097
rect 21726 10989 21727 11023
rect 21727 10989 21895 11023
rect 21895 10989 21896 11023
rect 21726 10988 21896 10989
rect 22098 11131 22268 11132
rect 22098 11097 22099 11131
rect 22099 11097 22267 11131
rect 22267 11097 22268 11131
rect 22098 11023 22268 11097
rect 22098 10989 22099 11023
rect 22099 10989 22267 11023
rect 22267 10989 22268 11023
rect 22098 10988 22268 10989
rect 22470 11131 22640 11132
rect 22470 11097 22471 11131
rect 22471 11097 22639 11131
rect 22639 11097 22640 11131
rect 22470 11023 22640 11097
rect 22470 10989 22471 11023
rect 22471 10989 22639 11023
rect 22639 10989 22640 11023
rect 22470 10988 22640 10989
rect 22842 11131 23012 11132
rect 22842 11097 22843 11131
rect 22843 11097 23011 11131
rect 23011 11097 23012 11131
rect 22842 11023 23012 11097
rect 22842 10989 22843 11023
rect 22843 10989 23011 11023
rect 23011 10989 23012 11023
rect 22842 10988 23012 10989
rect 23214 11131 23384 11132
rect 23214 11097 23215 11131
rect 23215 11097 23383 11131
rect 23383 11097 23384 11131
rect 23214 11023 23384 11097
rect 23214 10989 23215 11023
rect 23215 10989 23383 11023
rect 23383 10989 23384 11023
rect 23214 10988 23384 10989
rect 23586 11131 23756 11132
rect 23586 11097 23587 11131
rect 23587 11097 23755 11131
rect 23755 11097 23756 11131
rect 23586 11023 23756 11097
rect 23586 10989 23587 11023
rect 23587 10989 23755 11023
rect 23755 10989 23756 11023
rect 23586 10988 23756 10989
rect 23958 11131 24128 11132
rect 23958 11097 23959 11131
rect 23959 11097 24127 11131
rect 24127 11097 24128 11131
rect 23958 11023 24128 11097
rect 23958 10989 23959 11023
rect 23959 10989 24127 11023
rect 24127 10989 24128 11023
rect 23958 10988 24128 10989
rect 24330 11131 24500 11132
rect 24330 11097 24331 11131
rect 24331 11097 24499 11131
rect 24499 11097 24500 11131
rect 24330 11023 24500 11097
rect 24330 10989 24331 11023
rect 24331 10989 24499 11023
rect 24499 10989 24500 11023
rect 24330 10988 24500 10989
rect 18750 10495 18920 10496
rect 18750 10461 18751 10495
rect 18751 10461 18919 10495
rect 18919 10461 18920 10495
rect 18750 10387 18920 10461
rect 18750 10353 18751 10387
rect 18751 10353 18919 10387
rect 18919 10353 18920 10387
rect 18750 10352 18920 10353
rect 19122 10495 19292 10496
rect 19122 10461 19123 10495
rect 19123 10461 19291 10495
rect 19291 10461 19292 10495
rect 19122 10387 19292 10461
rect 19122 10353 19123 10387
rect 19123 10353 19291 10387
rect 19291 10353 19292 10387
rect 19122 10352 19292 10353
rect 19494 10495 19664 10496
rect 19494 10461 19495 10495
rect 19495 10461 19663 10495
rect 19663 10461 19664 10495
rect 19494 10387 19664 10461
rect 19494 10353 19495 10387
rect 19495 10353 19663 10387
rect 19663 10353 19664 10387
rect 19494 10352 19664 10353
rect 19866 10495 20036 10496
rect 19866 10461 19867 10495
rect 19867 10461 20035 10495
rect 20035 10461 20036 10495
rect 19866 10387 20036 10461
rect 19866 10353 19867 10387
rect 19867 10353 20035 10387
rect 20035 10353 20036 10387
rect 19866 10352 20036 10353
rect 20238 10495 20408 10496
rect 20238 10461 20239 10495
rect 20239 10461 20407 10495
rect 20407 10461 20408 10495
rect 20238 10387 20408 10461
rect 20238 10353 20239 10387
rect 20239 10353 20407 10387
rect 20407 10353 20408 10387
rect 20238 10352 20408 10353
rect 20610 10495 20780 10496
rect 20610 10461 20611 10495
rect 20611 10461 20779 10495
rect 20779 10461 20780 10495
rect 20610 10387 20780 10461
rect 20610 10353 20611 10387
rect 20611 10353 20779 10387
rect 20779 10353 20780 10387
rect 20610 10352 20780 10353
rect 20982 10495 21152 10496
rect 20982 10461 20983 10495
rect 20983 10461 21151 10495
rect 21151 10461 21152 10495
rect 20982 10387 21152 10461
rect 20982 10353 20983 10387
rect 20983 10353 21151 10387
rect 21151 10353 21152 10387
rect 20982 10352 21152 10353
rect 21354 10495 21524 10496
rect 21354 10461 21355 10495
rect 21355 10461 21523 10495
rect 21523 10461 21524 10495
rect 21354 10387 21524 10461
rect 21354 10353 21355 10387
rect 21355 10353 21523 10387
rect 21523 10353 21524 10387
rect 21354 10352 21524 10353
rect 21726 10495 21896 10496
rect 21726 10461 21727 10495
rect 21727 10461 21895 10495
rect 21895 10461 21896 10495
rect 21726 10387 21896 10461
rect 21726 10353 21727 10387
rect 21727 10353 21895 10387
rect 21895 10353 21896 10387
rect 21726 10352 21896 10353
rect 22098 10495 22268 10496
rect 22098 10461 22099 10495
rect 22099 10461 22267 10495
rect 22267 10461 22268 10495
rect 22098 10387 22268 10461
rect 22098 10353 22099 10387
rect 22099 10353 22267 10387
rect 22267 10353 22268 10387
rect 22098 10352 22268 10353
rect 22470 10495 22640 10496
rect 22470 10461 22471 10495
rect 22471 10461 22639 10495
rect 22639 10461 22640 10495
rect 22470 10387 22640 10461
rect 22470 10353 22471 10387
rect 22471 10353 22639 10387
rect 22639 10353 22640 10387
rect 22470 10352 22640 10353
rect 22842 10495 23012 10496
rect 22842 10461 22843 10495
rect 22843 10461 23011 10495
rect 23011 10461 23012 10495
rect 22842 10387 23012 10461
rect 22842 10353 22843 10387
rect 22843 10353 23011 10387
rect 23011 10353 23012 10387
rect 22842 10352 23012 10353
rect 23214 10495 23384 10496
rect 23214 10461 23215 10495
rect 23215 10461 23383 10495
rect 23383 10461 23384 10495
rect 23214 10387 23384 10461
rect 23214 10353 23215 10387
rect 23215 10353 23383 10387
rect 23383 10353 23384 10387
rect 23214 10352 23384 10353
rect 23586 10495 23756 10496
rect 23586 10461 23587 10495
rect 23587 10461 23755 10495
rect 23755 10461 23756 10495
rect 23586 10387 23756 10461
rect 23586 10353 23587 10387
rect 23587 10353 23755 10387
rect 23755 10353 23756 10387
rect 23586 10352 23756 10353
rect 23958 10495 24128 10496
rect 23958 10461 23959 10495
rect 23959 10461 24127 10495
rect 24127 10461 24128 10495
rect 23958 10387 24128 10461
rect 23958 10353 23959 10387
rect 23959 10353 24127 10387
rect 24127 10353 24128 10387
rect 23958 10352 24128 10353
rect 24330 10495 24500 10496
rect 24330 10461 24331 10495
rect 24331 10461 24499 10495
rect 24499 10461 24500 10495
rect 24330 10387 24500 10461
rect 24330 10353 24331 10387
rect 24331 10353 24499 10387
rect 24499 10353 24500 10387
rect 24330 10352 24500 10353
rect 18750 9859 18920 9872
rect 18750 9825 18751 9859
rect 18751 9825 18919 9859
rect 18919 9825 18920 9859
rect 18750 9812 18920 9825
rect 19122 9859 19292 9872
rect 19122 9825 19123 9859
rect 19123 9825 19291 9859
rect 19291 9825 19292 9859
rect 19122 9812 19292 9825
rect 19494 9859 19664 9872
rect 19494 9825 19495 9859
rect 19495 9825 19663 9859
rect 19663 9825 19664 9859
rect 19494 9812 19664 9825
rect 19866 9859 20036 9872
rect 19866 9825 19867 9859
rect 19867 9825 20035 9859
rect 20035 9825 20036 9859
rect 19866 9812 20036 9825
rect 20238 9859 20408 9872
rect 20238 9825 20239 9859
rect 20239 9825 20407 9859
rect 20407 9825 20408 9859
rect 20238 9812 20408 9825
rect 20610 9859 20780 9872
rect 20610 9825 20611 9859
rect 20611 9825 20779 9859
rect 20779 9825 20780 9859
rect 20610 9812 20780 9825
rect 20982 9859 21152 9872
rect 20982 9825 20983 9859
rect 20983 9825 21151 9859
rect 21151 9825 21152 9859
rect 20982 9812 21152 9825
rect 21354 9859 21524 9872
rect 21354 9825 21355 9859
rect 21355 9825 21523 9859
rect 21523 9825 21524 9859
rect 21354 9812 21524 9825
rect 21726 9859 21896 9872
rect 21726 9825 21727 9859
rect 21727 9825 21895 9859
rect 21895 9825 21896 9859
rect 21726 9812 21896 9825
rect 22098 9859 22268 9872
rect 22098 9825 22099 9859
rect 22099 9825 22267 9859
rect 22267 9825 22268 9859
rect 22098 9812 22268 9825
rect 22470 9859 22640 9872
rect 22470 9825 22471 9859
rect 22471 9825 22639 9859
rect 22639 9825 22640 9859
rect 22470 9812 22640 9825
rect 22842 9859 23012 9872
rect 22842 9825 22843 9859
rect 22843 9825 23011 9859
rect 23011 9825 23012 9859
rect 22842 9812 23012 9825
rect 23214 9859 23384 9872
rect 23214 9825 23215 9859
rect 23215 9825 23383 9859
rect 23383 9825 23384 9859
rect 23214 9812 23384 9825
rect 23586 9859 23756 9872
rect 23586 9825 23587 9859
rect 23587 9825 23755 9859
rect 23755 9825 23756 9859
rect 23586 9812 23756 9825
rect 24702 11659 24872 11672
rect 24702 11625 24703 11659
rect 24703 11625 24871 11659
rect 24871 11625 24872 11659
rect 24702 11612 24872 11625
rect 25074 11659 25244 11672
rect 25074 11625 25075 11659
rect 25075 11625 25243 11659
rect 25243 11625 25244 11659
rect 25074 11612 25244 11625
rect 25446 11659 25616 11672
rect 25446 11625 25447 11659
rect 25447 11625 25615 11659
rect 25615 11625 25616 11659
rect 25446 11612 25616 11625
rect 25818 11659 25988 11672
rect 25818 11625 25819 11659
rect 25819 11625 25987 11659
rect 25987 11625 25988 11659
rect 25818 11612 25988 11625
rect 26190 11659 26360 11672
rect 26190 11625 26191 11659
rect 26191 11625 26359 11659
rect 26359 11625 26360 11659
rect 26190 11612 26360 11625
rect 26562 11659 26732 11672
rect 26562 11625 26563 11659
rect 26563 11625 26731 11659
rect 26731 11625 26732 11659
rect 26562 11612 26732 11625
rect 26934 11659 27104 11672
rect 26934 11625 26935 11659
rect 26935 11625 27103 11659
rect 27103 11625 27104 11659
rect 26934 11612 27104 11625
rect 27306 11659 27476 11672
rect 27306 11625 27307 11659
rect 27307 11625 27475 11659
rect 27475 11625 27476 11659
rect 27306 11612 27476 11625
rect 27678 11659 27848 11672
rect 27678 11625 27679 11659
rect 27679 11625 27847 11659
rect 27847 11625 27848 11659
rect 27678 11612 27848 11625
rect 28050 11659 28220 11672
rect 28050 11625 28051 11659
rect 28051 11625 28219 11659
rect 28219 11625 28220 11659
rect 28050 11612 28220 11625
rect 28422 11659 28592 11672
rect 28422 11625 28423 11659
rect 28423 11625 28591 11659
rect 28591 11625 28592 11659
rect 28422 11612 28592 11625
rect 28794 11659 28964 11672
rect 28794 11625 28795 11659
rect 28795 11625 28963 11659
rect 28963 11625 28964 11659
rect 28794 11612 28964 11625
rect 29166 11659 29336 11672
rect 29166 11625 29167 11659
rect 29167 11625 29335 11659
rect 29335 11625 29336 11659
rect 29166 11612 29336 11625
rect 29538 11659 29708 11672
rect 29538 11625 29539 11659
rect 29539 11625 29707 11659
rect 29707 11625 29708 11659
rect 29538 11612 29708 11625
rect 29910 11659 30080 11672
rect 29910 11625 29911 11659
rect 29911 11625 30079 11659
rect 30079 11625 30080 11659
rect 29910 11612 30080 11625
rect 30282 11659 30452 11672
rect 30282 11625 30283 11659
rect 30283 11625 30451 11659
rect 30451 11625 30452 11659
rect 30282 11612 30452 11625
rect 24702 11131 24872 11132
rect 24702 11097 24703 11131
rect 24703 11097 24871 11131
rect 24871 11097 24872 11131
rect 24702 11023 24872 11097
rect 24702 10989 24703 11023
rect 24703 10989 24871 11023
rect 24871 10989 24872 11023
rect 24702 10988 24872 10989
rect 25074 11131 25244 11132
rect 25074 11097 25075 11131
rect 25075 11097 25243 11131
rect 25243 11097 25244 11131
rect 25074 11023 25244 11097
rect 25074 10989 25075 11023
rect 25075 10989 25243 11023
rect 25243 10989 25244 11023
rect 25074 10988 25244 10989
rect 25446 11131 25616 11132
rect 25446 11097 25447 11131
rect 25447 11097 25615 11131
rect 25615 11097 25616 11131
rect 25446 11023 25616 11097
rect 25446 10989 25447 11023
rect 25447 10989 25615 11023
rect 25615 10989 25616 11023
rect 25446 10988 25616 10989
rect 25818 11131 25988 11132
rect 25818 11097 25819 11131
rect 25819 11097 25987 11131
rect 25987 11097 25988 11131
rect 25818 11023 25988 11097
rect 25818 10989 25819 11023
rect 25819 10989 25987 11023
rect 25987 10989 25988 11023
rect 25818 10988 25988 10989
rect 26190 11131 26360 11132
rect 26190 11097 26191 11131
rect 26191 11097 26359 11131
rect 26359 11097 26360 11131
rect 26190 11023 26360 11097
rect 26190 10989 26191 11023
rect 26191 10989 26359 11023
rect 26359 10989 26360 11023
rect 26190 10988 26360 10989
rect 26562 11131 26732 11132
rect 26562 11097 26563 11131
rect 26563 11097 26731 11131
rect 26731 11097 26732 11131
rect 26562 11023 26732 11097
rect 26562 10989 26563 11023
rect 26563 10989 26731 11023
rect 26731 10989 26732 11023
rect 26562 10988 26732 10989
rect 26934 11131 27104 11132
rect 26934 11097 26935 11131
rect 26935 11097 27103 11131
rect 27103 11097 27104 11131
rect 26934 11023 27104 11097
rect 26934 10989 26935 11023
rect 26935 10989 27103 11023
rect 27103 10989 27104 11023
rect 26934 10988 27104 10989
rect 27306 11131 27476 11132
rect 27306 11097 27307 11131
rect 27307 11097 27475 11131
rect 27475 11097 27476 11131
rect 27306 11023 27476 11097
rect 27306 10989 27307 11023
rect 27307 10989 27475 11023
rect 27475 10989 27476 11023
rect 27306 10988 27476 10989
rect 27678 11131 27848 11132
rect 27678 11097 27679 11131
rect 27679 11097 27847 11131
rect 27847 11097 27848 11131
rect 27678 11023 27848 11097
rect 27678 10989 27679 11023
rect 27679 10989 27847 11023
rect 27847 10989 27848 11023
rect 27678 10988 27848 10989
rect 28050 11131 28220 11132
rect 28050 11097 28051 11131
rect 28051 11097 28219 11131
rect 28219 11097 28220 11131
rect 28050 11023 28220 11097
rect 28050 10989 28051 11023
rect 28051 10989 28219 11023
rect 28219 10989 28220 11023
rect 28050 10988 28220 10989
rect 28422 11131 28592 11132
rect 28422 11097 28423 11131
rect 28423 11097 28591 11131
rect 28591 11097 28592 11131
rect 28422 11023 28592 11097
rect 28422 10989 28423 11023
rect 28423 10989 28591 11023
rect 28591 10989 28592 11023
rect 28422 10988 28592 10989
rect 28794 11131 28964 11132
rect 28794 11097 28795 11131
rect 28795 11097 28963 11131
rect 28963 11097 28964 11131
rect 28794 11023 28964 11097
rect 28794 10989 28795 11023
rect 28795 10989 28963 11023
rect 28963 10989 28964 11023
rect 28794 10988 28964 10989
rect 29166 11131 29336 11132
rect 29166 11097 29167 11131
rect 29167 11097 29335 11131
rect 29335 11097 29336 11131
rect 29166 11023 29336 11097
rect 29166 10989 29167 11023
rect 29167 10989 29335 11023
rect 29335 10989 29336 11023
rect 29166 10988 29336 10989
rect 29538 11131 29708 11132
rect 29538 11097 29539 11131
rect 29539 11097 29707 11131
rect 29707 11097 29708 11131
rect 29538 11023 29708 11097
rect 29538 10989 29539 11023
rect 29539 10989 29707 11023
rect 29707 10989 29708 11023
rect 29538 10988 29708 10989
rect 29910 11131 30080 11132
rect 29910 11097 29911 11131
rect 29911 11097 30079 11131
rect 30079 11097 30080 11131
rect 29910 11023 30080 11097
rect 29910 10989 29911 11023
rect 29911 10989 30079 11023
rect 30079 10989 30080 11023
rect 29910 10988 30080 10989
rect 30282 11131 30452 11132
rect 30282 11097 30283 11131
rect 30283 11097 30451 11131
rect 30451 11097 30452 11131
rect 30282 11023 30452 11097
rect 30282 10989 30283 11023
rect 30283 10989 30451 11023
rect 30451 10989 30452 11023
rect 30282 10988 30452 10989
rect 24702 10495 24872 10496
rect 24702 10461 24703 10495
rect 24703 10461 24871 10495
rect 24871 10461 24872 10495
rect 24702 10387 24872 10461
rect 24702 10353 24703 10387
rect 24703 10353 24871 10387
rect 24871 10353 24872 10387
rect 24702 10352 24872 10353
rect 25074 10495 25244 10496
rect 25074 10461 25075 10495
rect 25075 10461 25243 10495
rect 25243 10461 25244 10495
rect 25074 10387 25244 10461
rect 25074 10353 25075 10387
rect 25075 10353 25243 10387
rect 25243 10353 25244 10387
rect 25074 10352 25244 10353
rect 25446 10495 25616 10496
rect 25446 10461 25447 10495
rect 25447 10461 25615 10495
rect 25615 10461 25616 10495
rect 25446 10387 25616 10461
rect 25446 10353 25447 10387
rect 25447 10353 25615 10387
rect 25615 10353 25616 10387
rect 25446 10352 25616 10353
rect 25818 10495 25988 10496
rect 25818 10461 25819 10495
rect 25819 10461 25987 10495
rect 25987 10461 25988 10495
rect 25818 10387 25988 10461
rect 25818 10353 25819 10387
rect 25819 10353 25987 10387
rect 25987 10353 25988 10387
rect 25818 10352 25988 10353
rect 26190 10495 26360 10496
rect 26190 10461 26191 10495
rect 26191 10461 26359 10495
rect 26359 10461 26360 10495
rect 26190 10387 26360 10461
rect 26190 10353 26191 10387
rect 26191 10353 26359 10387
rect 26359 10353 26360 10387
rect 26190 10352 26360 10353
rect 26562 10495 26732 10496
rect 26562 10461 26563 10495
rect 26563 10461 26731 10495
rect 26731 10461 26732 10495
rect 26562 10387 26732 10461
rect 26562 10353 26563 10387
rect 26563 10353 26731 10387
rect 26731 10353 26732 10387
rect 26562 10352 26732 10353
rect 26934 10495 27104 10496
rect 26934 10461 26935 10495
rect 26935 10461 27103 10495
rect 27103 10461 27104 10495
rect 26934 10387 27104 10461
rect 26934 10353 26935 10387
rect 26935 10353 27103 10387
rect 27103 10353 27104 10387
rect 26934 10352 27104 10353
rect 27306 10495 27476 10496
rect 27306 10461 27307 10495
rect 27307 10461 27475 10495
rect 27475 10461 27476 10495
rect 27306 10387 27476 10461
rect 27306 10353 27307 10387
rect 27307 10353 27475 10387
rect 27475 10353 27476 10387
rect 27306 10352 27476 10353
rect 27678 10495 27848 10496
rect 27678 10461 27679 10495
rect 27679 10461 27847 10495
rect 27847 10461 27848 10495
rect 27678 10387 27848 10461
rect 27678 10353 27679 10387
rect 27679 10353 27847 10387
rect 27847 10353 27848 10387
rect 27678 10352 27848 10353
rect 28050 10495 28220 10496
rect 28050 10461 28051 10495
rect 28051 10461 28219 10495
rect 28219 10461 28220 10495
rect 28050 10387 28220 10461
rect 28050 10353 28051 10387
rect 28051 10353 28219 10387
rect 28219 10353 28220 10387
rect 28050 10352 28220 10353
rect 28422 10495 28592 10496
rect 28422 10461 28423 10495
rect 28423 10461 28591 10495
rect 28591 10461 28592 10495
rect 28422 10387 28592 10461
rect 28422 10353 28423 10387
rect 28423 10353 28591 10387
rect 28591 10353 28592 10387
rect 28422 10352 28592 10353
rect 28794 10495 28964 10496
rect 28794 10461 28795 10495
rect 28795 10461 28963 10495
rect 28963 10461 28964 10495
rect 28794 10387 28964 10461
rect 28794 10353 28795 10387
rect 28795 10353 28963 10387
rect 28963 10353 28964 10387
rect 28794 10352 28964 10353
rect 29166 10495 29336 10496
rect 29166 10461 29167 10495
rect 29167 10461 29335 10495
rect 29335 10461 29336 10495
rect 29166 10387 29336 10461
rect 29166 10353 29167 10387
rect 29167 10353 29335 10387
rect 29335 10353 29336 10387
rect 29166 10352 29336 10353
rect 29538 10495 29708 10496
rect 29538 10461 29539 10495
rect 29539 10461 29707 10495
rect 29707 10461 29708 10495
rect 29538 10387 29708 10461
rect 29538 10353 29539 10387
rect 29539 10353 29707 10387
rect 29707 10353 29708 10387
rect 29538 10352 29708 10353
rect 29910 10495 30080 10496
rect 29910 10461 29911 10495
rect 29911 10461 30079 10495
rect 30079 10461 30080 10495
rect 29910 10387 30080 10461
rect 29910 10353 29911 10387
rect 29911 10353 30079 10387
rect 30079 10353 30080 10387
rect 29910 10352 30080 10353
rect 30282 10495 30452 10496
rect 30282 10461 30283 10495
rect 30283 10461 30451 10495
rect 30451 10461 30452 10495
rect 30282 10387 30452 10461
rect 30282 10353 30283 10387
rect 30283 10353 30451 10387
rect 30451 10353 30452 10387
rect 30282 10352 30452 10353
rect 23958 9859 24128 9872
rect 23958 9825 23959 9859
rect 23959 9825 24127 9859
rect 24127 9825 24128 9859
rect 23958 9812 24128 9825
rect 24330 9859 24500 9872
rect 24330 9825 24331 9859
rect 24331 9825 24499 9859
rect 24499 9825 24500 9859
rect 24330 9812 24500 9825
rect 24702 9859 24872 9872
rect 24702 9825 24703 9859
rect 24703 9825 24871 9859
rect 24871 9825 24872 9859
rect 24702 9812 24872 9825
rect 25074 9859 25244 9872
rect 25074 9825 25075 9859
rect 25075 9825 25243 9859
rect 25243 9825 25244 9859
rect 25074 9812 25244 9825
rect 25446 9859 25616 9872
rect 25446 9825 25447 9859
rect 25447 9825 25615 9859
rect 25615 9825 25616 9859
rect 25446 9812 25616 9825
rect 25818 9859 25988 9872
rect 25818 9825 25819 9859
rect 25819 9825 25987 9859
rect 25987 9825 25988 9859
rect 25818 9812 25988 9825
rect 26190 9859 26360 9872
rect 26190 9825 26191 9859
rect 26191 9825 26359 9859
rect 26359 9825 26360 9859
rect 26190 9812 26360 9825
rect 26562 9859 26732 9872
rect 26562 9825 26563 9859
rect 26563 9825 26731 9859
rect 26731 9825 26732 9859
rect 26562 9812 26732 9825
rect 26934 9859 27104 9872
rect 26934 9825 26935 9859
rect 26935 9825 27103 9859
rect 27103 9825 27104 9859
rect 26934 9812 27104 9825
rect 27306 9859 27476 9872
rect 27306 9825 27307 9859
rect 27307 9825 27475 9859
rect 27475 9825 27476 9859
rect 27306 9812 27476 9825
rect 27678 9859 27848 9872
rect 27678 9825 27679 9859
rect 27679 9825 27847 9859
rect 27847 9825 27848 9859
rect 27678 9812 27848 9825
rect 28050 9859 28220 9872
rect 28050 9825 28051 9859
rect 28051 9825 28219 9859
rect 28219 9825 28220 9859
rect 28050 9812 28220 9825
rect 28422 9859 28592 9872
rect 28422 9825 28423 9859
rect 28423 9825 28591 9859
rect 28591 9825 28592 9859
rect 28422 9812 28592 9825
rect 28794 9859 28964 9872
rect 28794 9825 28795 9859
rect 28795 9825 28963 9859
rect 28963 9825 28964 9859
rect 28794 9812 28964 9825
rect 29166 9859 29336 9872
rect 29166 9825 29167 9859
rect 29167 9825 29335 9859
rect 29335 9825 29336 9859
rect 29166 9812 29336 9825
rect 29538 9859 29708 9872
rect 29538 9825 29539 9859
rect 29539 9825 29707 9859
rect 29707 9825 29708 9859
rect 29538 9812 29708 9825
rect 29910 9859 30080 9872
rect 29910 9825 29911 9859
rect 29911 9825 30079 9859
rect 30079 9825 30080 9859
rect 29910 9812 30080 9825
rect 30282 9859 30452 9872
rect 30282 9825 30283 9859
rect 30283 9825 30451 9859
rect 30451 9825 30452 9859
rect 30282 9812 30452 9825
rect 20238 9271 20408 9286
rect 20238 9237 20239 9271
rect 20239 9237 20407 9271
rect 20407 9237 20408 9271
rect 20238 9222 20408 9237
rect 20610 9271 20780 9286
rect 20610 9237 20611 9271
rect 20611 9237 20779 9271
rect 20779 9237 20780 9271
rect 20610 9222 20780 9237
rect 20982 9271 21152 9286
rect 20982 9237 20983 9271
rect 20983 9237 21151 9271
rect 21151 9237 21152 9271
rect 20982 9222 21152 9237
rect 21354 9271 21524 9286
rect 21354 9237 21355 9271
rect 21355 9237 21523 9271
rect 21523 9237 21524 9271
rect 21354 9222 21524 9237
rect 21726 9271 21896 9286
rect 21726 9237 21727 9271
rect 21727 9237 21895 9271
rect 21895 9237 21896 9271
rect 21726 9222 21896 9237
rect 22098 9271 22268 9286
rect 22098 9237 22099 9271
rect 22099 9237 22267 9271
rect 22267 9237 22268 9271
rect 22098 9222 22268 9237
rect 22470 9271 22640 9286
rect 22470 9237 22471 9271
rect 22471 9237 22639 9271
rect 22639 9237 22640 9271
rect 22470 9222 22640 9237
rect 22842 9271 23012 9286
rect 22842 9237 22843 9271
rect 22843 9237 23011 9271
rect 23011 9237 23012 9271
rect 22842 9222 23012 9237
rect 24834 9232 25116 9504
rect 25578 9232 25860 9504
rect 26322 9232 26604 9504
rect 27066 9232 27348 9504
rect 27810 9232 28092 9504
rect 28554 9232 28836 9504
rect 29298 9232 29580 9504
rect 30042 9232 30324 9504
rect 20238 8343 20408 8344
rect 20238 8309 20239 8343
rect 20239 8309 20407 8343
rect 20407 8309 20408 8343
rect 20238 8235 20408 8309
rect 20238 8201 20239 8235
rect 20239 8201 20407 8235
rect 20407 8201 20408 8235
rect 20238 8200 20408 8201
rect 20610 8343 20780 8344
rect 20610 8309 20611 8343
rect 20611 8309 20779 8343
rect 20779 8309 20780 8343
rect 20610 8235 20780 8309
rect 20610 8201 20611 8235
rect 20611 8201 20779 8235
rect 20779 8201 20780 8235
rect 20610 8200 20780 8201
rect 20982 8343 21152 8344
rect 20982 8309 20983 8343
rect 20983 8309 21151 8343
rect 21151 8309 21152 8343
rect 20982 8235 21152 8309
rect 20982 8201 20983 8235
rect 20983 8201 21151 8235
rect 21151 8201 21152 8235
rect 20982 8200 21152 8201
rect 21354 8343 21524 8344
rect 21354 8309 21355 8343
rect 21355 8309 21523 8343
rect 21523 8309 21524 8343
rect 21354 8235 21524 8309
rect 21354 8201 21355 8235
rect 21355 8201 21523 8235
rect 21523 8201 21524 8235
rect 21354 8200 21524 8201
rect 21726 8343 21896 8344
rect 21726 8309 21727 8343
rect 21727 8309 21895 8343
rect 21895 8309 21896 8343
rect 21726 8235 21896 8309
rect 21726 8201 21727 8235
rect 21727 8201 21895 8235
rect 21895 8201 21896 8235
rect 21726 8200 21896 8201
rect 22098 8343 22268 8344
rect 22098 8309 22099 8343
rect 22099 8309 22267 8343
rect 22267 8309 22268 8343
rect 22098 8235 22268 8309
rect 22098 8201 22099 8235
rect 22099 8201 22267 8235
rect 22267 8201 22268 8235
rect 22098 8200 22268 8201
rect 22470 8343 22640 8344
rect 22470 8309 22471 8343
rect 22471 8309 22639 8343
rect 22639 8309 22640 8343
rect 22470 8235 22640 8309
rect 22470 8201 22471 8235
rect 22471 8201 22639 8235
rect 22639 8201 22640 8235
rect 22470 8200 22640 8201
rect 22842 8343 23012 8344
rect 22842 8309 22843 8343
rect 22843 8309 23011 8343
rect 23011 8309 23012 8343
rect 22842 8235 23012 8309
rect 22842 8201 22843 8235
rect 22843 8201 23011 8235
rect 23011 8201 23012 8235
rect 22842 8200 23012 8201
rect 23716 7516 23998 7788
rect 20238 7307 20408 7308
rect 20238 7273 20239 7307
rect 20239 7273 20407 7307
rect 20407 7273 20408 7307
rect 20238 7199 20408 7273
rect 20238 7165 20239 7199
rect 20239 7165 20407 7199
rect 20407 7165 20408 7199
rect 20238 7164 20408 7165
rect 20610 7307 20780 7308
rect 20610 7273 20611 7307
rect 20611 7273 20779 7307
rect 20779 7273 20780 7307
rect 20610 7199 20780 7273
rect 20610 7165 20611 7199
rect 20611 7165 20779 7199
rect 20779 7165 20780 7199
rect 20610 7164 20780 7165
rect 20982 7307 21152 7308
rect 20982 7273 20983 7307
rect 20983 7273 21151 7307
rect 21151 7273 21152 7307
rect 20982 7199 21152 7273
rect 20982 7165 20983 7199
rect 20983 7165 21151 7199
rect 21151 7165 21152 7199
rect 20982 7164 21152 7165
rect 21354 7307 21524 7308
rect 21354 7273 21355 7307
rect 21355 7273 21523 7307
rect 21523 7273 21524 7307
rect 21354 7199 21524 7273
rect 21354 7165 21355 7199
rect 21355 7165 21523 7199
rect 21523 7165 21524 7199
rect 21354 7164 21524 7165
rect 21726 7307 21896 7308
rect 21726 7273 21727 7307
rect 21727 7273 21895 7307
rect 21895 7273 21896 7307
rect 21726 7199 21896 7273
rect 21726 7165 21727 7199
rect 21727 7165 21895 7199
rect 21895 7165 21896 7199
rect 21726 7164 21896 7165
rect 22098 7307 22268 7308
rect 22098 7273 22099 7307
rect 22099 7273 22267 7307
rect 22267 7273 22268 7307
rect 22098 7199 22268 7273
rect 22098 7165 22099 7199
rect 22099 7165 22267 7199
rect 22267 7165 22268 7199
rect 22098 7164 22268 7165
rect 22470 7307 22640 7308
rect 22470 7273 22471 7307
rect 22471 7273 22639 7307
rect 22639 7273 22640 7307
rect 22470 7199 22640 7273
rect 22470 7165 22471 7199
rect 22471 7165 22639 7199
rect 22639 7165 22640 7199
rect 22470 7164 22640 7165
rect 22842 7307 23012 7308
rect 22842 7273 22843 7307
rect 22843 7273 23011 7307
rect 23011 7273 23012 7307
rect 22842 7199 23012 7273
rect 22842 7165 22843 7199
rect 22843 7165 23011 7199
rect 23011 7165 23012 7199
rect 22842 7164 23012 7165
rect 24132 6688 24330 6886
rect 20238 6271 20408 6272
rect 20238 6237 20239 6271
rect 20239 6237 20407 6271
rect 20407 6237 20408 6271
rect 20238 6163 20408 6237
rect 20238 6129 20239 6163
rect 20239 6129 20407 6163
rect 20407 6129 20408 6163
rect 20238 6128 20408 6129
rect 20610 6271 20780 6272
rect 20610 6237 20611 6271
rect 20611 6237 20779 6271
rect 20779 6237 20780 6271
rect 20610 6163 20780 6237
rect 20610 6129 20611 6163
rect 20611 6129 20779 6163
rect 20779 6129 20780 6163
rect 20610 6128 20780 6129
rect 20982 6271 21152 6272
rect 20982 6237 20983 6271
rect 20983 6237 21151 6271
rect 21151 6237 21152 6271
rect 20982 6163 21152 6237
rect 20982 6129 20983 6163
rect 20983 6129 21151 6163
rect 21151 6129 21152 6163
rect 20982 6128 21152 6129
rect 21354 6271 21524 6272
rect 21354 6237 21355 6271
rect 21355 6237 21523 6271
rect 21523 6237 21524 6271
rect 21354 6163 21524 6237
rect 21354 6129 21355 6163
rect 21355 6129 21523 6163
rect 21523 6129 21524 6163
rect 21354 6128 21524 6129
rect 21726 6271 21896 6272
rect 21726 6237 21727 6271
rect 21727 6237 21895 6271
rect 21895 6237 21896 6271
rect 21726 6163 21896 6237
rect 21726 6129 21727 6163
rect 21727 6129 21895 6163
rect 21895 6129 21896 6163
rect 21726 6128 21896 6129
rect 22098 6271 22268 6272
rect 22098 6237 22099 6271
rect 22099 6237 22267 6271
rect 22267 6237 22268 6271
rect 22098 6163 22268 6237
rect 22098 6129 22099 6163
rect 22099 6129 22267 6163
rect 22267 6129 22268 6163
rect 22098 6128 22268 6129
rect 22470 6271 22640 6272
rect 22470 6237 22471 6271
rect 22471 6237 22639 6271
rect 22639 6237 22640 6271
rect 22470 6163 22640 6237
rect 22470 6129 22471 6163
rect 22471 6129 22639 6163
rect 22639 6129 22640 6163
rect 22470 6128 22640 6129
rect 22842 6271 23012 6272
rect 22842 6237 22843 6271
rect 22843 6237 23011 6271
rect 23011 6237 23012 6271
rect 22842 6163 23012 6237
rect 22842 6129 22843 6163
rect 22843 6129 23011 6163
rect 23011 6129 23012 6163
rect 22842 6128 23012 6129
rect 24132 6288 24330 6486
rect 20238 5235 20408 5246
rect 20238 5201 20239 5235
rect 20239 5201 20407 5235
rect 20407 5201 20408 5235
rect 20238 5192 20408 5201
rect 20610 5235 20780 5246
rect 20610 5201 20611 5235
rect 20611 5201 20779 5235
rect 20779 5201 20780 5235
rect 20610 5192 20780 5201
rect 20982 5235 21152 5246
rect 20982 5201 20983 5235
rect 20983 5201 21151 5235
rect 21151 5201 21152 5235
rect 20982 5192 21152 5201
rect 21354 5235 21524 5246
rect 21354 5201 21355 5235
rect 21355 5201 21523 5235
rect 21523 5201 21524 5235
rect 21354 5192 21524 5201
rect 21726 5235 21896 5246
rect 21726 5201 21727 5235
rect 21727 5201 21895 5235
rect 21895 5201 21896 5235
rect 21726 5192 21896 5201
rect 22098 5235 22268 5246
rect 22098 5201 22099 5235
rect 22099 5201 22267 5235
rect 22267 5201 22268 5235
rect 22098 5192 22268 5201
rect 22470 5235 22640 5246
rect 22470 5201 22471 5235
rect 22471 5201 22639 5235
rect 22639 5201 22640 5235
rect 22470 5192 22640 5201
rect 21218 4726 22032 4906
rect 20238 4577 20408 4588
rect 20238 4543 20239 4577
rect 20239 4543 20407 4577
rect 20407 4543 20408 4577
rect 20238 4532 20408 4543
rect 20610 4577 20780 4588
rect 20610 4543 20611 4577
rect 20611 4543 20779 4577
rect 20779 4543 20780 4577
rect 20610 4532 20780 4543
rect 20982 4577 21152 4588
rect 20982 4543 20983 4577
rect 20983 4543 21151 4577
rect 21151 4543 21152 4577
rect 20982 4532 21152 4543
rect 21354 4577 21524 4588
rect 21354 4543 21355 4577
rect 21355 4543 21523 4577
rect 21523 4543 21524 4577
rect 21354 4532 21524 4543
rect 21726 4577 21896 4588
rect 21726 4543 21727 4577
rect 21727 4543 21895 4577
rect 21895 4543 21896 4577
rect 21726 4532 21896 4543
rect 22842 5235 23012 5246
rect 22842 5201 22843 5235
rect 22843 5201 23011 5235
rect 23011 5201 23012 5235
rect 22842 5192 23012 5201
rect 23344 5050 23626 5322
rect 22098 4577 22268 4588
rect 22098 4543 22099 4577
rect 22099 4543 22267 4577
rect 22267 4543 22268 4577
rect 22098 4532 22268 4543
rect 22470 4577 22640 4588
rect 22470 4543 22471 4577
rect 22471 4543 22639 4577
rect 22639 4543 22640 4577
rect 22470 4532 22640 4543
rect 22842 4577 23012 4588
rect 22842 4543 22843 4577
rect 22843 4543 23011 4577
rect 23011 4543 23012 4577
rect 22842 4532 23012 4543
rect 23214 4577 23384 4588
rect 23214 4543 23215 4577
rect 23215 4543 23383 4577
rect 23383 4543 23384 4577
rect 23214 4532 23384 4543
rect 24132 5888 24330 6086
rect 24088 5050 24370 5322
rect 24832 5050 25114 5322
rect 25576 5050 25858 5322
rect 26320 5050 26602 5322
rect 27064 5050 27346 5322
rect 27808 5050 28090 5322
rect 28552 5050 28834 5322
rect 23724 4726 23974 4976
rect 23586 4577 23756 4588
rect 23586 4543 23587 4577
rect 23587 4543 23755 4577
rect 23755 4543 23756 4577
rect 23586 4532 23756 4543
rect 23958 4577 24128 4588
rect 23958 4543 23959 4577
rect 23959 4543 24127 4577
rect 24127 4543 24128 4577
rect 23958 4532 24128 4543
rect 24330 4577 24500 4588
rect 24330 4543 24331 4577
rect 24331 4543 24499 4577
rect 24499 4543 24500 4577
rect 24330 4532 24500 4543
rect 24702 4577 24872 4588
rect 24702 4543 24703 4577
rect 24703 4543 24871 4577
rect 24871 4543 24872 4577
rect 24702 4532 24872 4543
rect 25074 4577 25244 4588
rect 25074 4543 25075 4577
rect 25075 4543 25243 4577
rect 25243 4543 25244 4577
rect 25074 4532 25244 4543
rect 25446 4577 25616 4588
rect 25446 4543 25447 4577
rect 25447 4543 25615 4577
rect 25615 4543 25616 4577
rect 25446 4532 25616 4543
rect 25818 4577 25988 4588
rect 25818 4543 25819 4577
rect 25819 4543 25987 4577
rect 25987 4543 25988 4577
rect 25818 4532 25988 4543
rect 26190 4577 26360 4588
rect 26190 4543 26191 4577
rect 26191 4543 26359 4577
rect 26359 4543 26360 4577
rect 26190 4532 26360 4543
rect 26562 4577 26732 4588
rect 26562 4543 26563 4577
rect 26563 4543 26731 4577
rect 26731 4543 26732 4577
rect 26562 4532 26732 4543
rect 26934 4577 27104 4588
rect 26934 4543 26935 4577
rect 26935 4543 27103 4577
rect 27103 4543 27104 4577
rect 26934 4532 27104 4543
rect 27306 4577 27476 4588
rect 27306 4543 27307 4577
rect 27307 4543 27475 4577
rect 27475 4543 27476 4577
rect 27306 4532 27476 4543
rect 27678 4577 27848 4588
rect 27678 4543 27679 4577
rect 27679 4543 27847 4577
rect 27847 4543 27848 4577
rect 27678 4532 27848 4543
rect 28050 4577 28220 4588
rect 28050 4543 28051 4577
rect 28051 4543 28219 4577
rect 28219 4543 28220 4577
rect 28050 4532 28220 4543
rect 28422 4577 28592 4588
rect 28422 4543 28423 4577
rect 28423 4543 28591 4577
rect 28591 4543 28592 4577
rect 28422 4532 28592 4543
rect 28794 4577 28964 4588
rect 28794 4543 28795 4577
rect 28795 4543 28963 4577
rect 28963 4543 28964 4577
rect 28794 4532 28964 4543
rect 20238 4267 20408 4268
rect 20238 4233 20239 4267
rect 20239 4233 20407 4267
rect 20407 4233 20408 4267
rect 20238 4159 20408 4233
rect 20238 4125 20239 4159
rect 20239 4125 20407 4159
rect 20407 4125 20408 4159
rect 20238 4124 20408 4125
rect 20610 4267 20780 4268
rect 20610 4233 20611 4267
rect 20611 4233 20779 4267
rect 20779 4233 20780 4267
rect 20610 4159 20780 4233
rect 20610 4125 20611 4159
rect 20611 4125 20779 4159
rect 20779 4125 20780 4159
rect 20610 4124 20780 4125
rect 20982 4267 21152 4268
rect 20982 4233 20983 4267
rect 20983 4233 21151 4267
rect 21151 4233 21152 4267
rect 20982 4159 21152 4233
rect 20982 4125 20983 4159
rect 20983 4125 21151 4159
rect 21151 4125 21152 4159
rect 20982 4124 21152 4125
rect 21354 4267 21524 4268
rect 21354 4233 21355 4267
rect 21355 4233 21523 4267
rect 21523 4233 21524 4267
rect 21354 4159 21524 4233
rect 21354 4125 21355 4159
rect 21355 4125 21523 4159
rect 21523 4125 21524 4159
rect 21354 4124 21524 4125
rect 21726 4267 21896 4268
rect 21726 4233 21727 4267
rect 21727 4233 21895 4267
rect 21895 4233 21896 4267
rect 21726 4159 21896 4233
rect 21726 4125 21727 4159
rect 21727 4125 21895 4159
rect 21895 4125 21896 4159
rect 21726 4124 21896 4125
rect 22098 4267 22268 4268
rect 22098 4233 22099 4267
rect 22099 4233 22267 4267
rect 22267 4233 22268 4267
rect 22098 4159 22268 4233
rect 22098 4125 22099 4159
rect 22099 4125 22267 4159
rect 22267 4125 22268 4159
rect 22098 4124 22268 4125
rect 22470 4267 22640 4268
rect 22470 4233 22471 4267
rect 22471 4233 22639 4267
rect 22639 4233 22640 4267
rect 22470 4159 22640 4233
rect 22470 4125 22471 4159
rect 22471 4125 22639 4159
rect 22639 4125 22640 4159
rect 22470 4124 22640 4125
rect 22842 4267 23012 4268
rect 22842 4233 22843 4267
rect 22843 4233 23011 4267
rect 23011 4233 23012 4267
rect 22842 4159 23012 4233
rect 22842 4125 22843 4159
rect 22843 4125 23011 4159
rect 23011 4125 23012 4159
rect 22842 4124 23012 4125
rect 23214 4267 23384 4268
rect 23214 4233 23215 4267
rect 23215 4233 23383 4267
rect 23383 4233 23384 4267
rect 23214 4159 23384 4233
rect 23214 4125 23215 4159
rect 23215 4125 23383 4159
rect 23383 4125 23384 4159
rect 23214 4124 23384 4125
rect 23586 4267 23756 4268
rect 23586 4233 23587 4267
rect 23587 4233 23755 4267
rect 23755 4233 23756 4267
rect 23586 4159 23756 4233
rect 23586 4125 23587 4159
rect 23587 4125 23755 4159
rect 23755 4125 23756 4159
rect 23586 4124 23756 4125
rect 23958 4267 24128 4268
rect 23958 4233 23959 4267
rect 23959 4233 24127 4267
rect 24127 4233 24128 4267
rect 23958 4159 24128 4233
rect 23958 4125 23959 4159
rect 23959 4125 24127 4159
rect 24127 4125 24128 4159
rect 23958 4124 24128 4125
rect 24330 4267 24500 4268
rect 24330 4233 24331 4267
rect 24331 4233 24499 4267
rect 24499 4233 24500 4267
rect 24330 4159 24500 4233
rect 24330 4125 24331 4159
rect 24331 4125 24499 4159
rect 24499 4125 24500 4159
rect 24330 4124 24500 4125
rect 24702 4267 24872 4268
rect 24702 4233 24703 4267
rect 24703 4233 24871 4267
rect 24871 4233 24872 4267
rect 24702 4159 24872 4233
rect 24702 4125 24703 4159
rect 24703 4125 24871 4159
rect 24871 4125 24872 4159
rect 24702 4124 24872 4125
rect 25074 4267 25244 4268
rect 25074 4233 25075 4267
rect 25075 4233 25243 4267
rect 25243 4233 25244 4267
rect 25074 4159 25244 4233
rect 25074 4125 25075 4159
rect 25075 4125 25243 4159
rect 25243 4125 25244 4159
rect 25074 4124 25244 4125
rect 25446 4267 25616 4268
rect 25446 4233 25447 4267
rect 25447 4233 25615 4267
rect 25615 4233 25616 4267
rect 25446 4159 25616 4233
rect 25446 4125 25447 4159
rect 25447 4125 25615 4159
rect 25615 4125 25616 4159
rect 25446 4124 25616 4125
rect 25818 4267 25988 4268
rect 25818 4233 25819 4267
rect 25819 4233 25987 4267
rect 25987 4233 25988 4267
rect 25818 4159 25988 4233
rect 25818 4125 25819 4159
rect 25819 4125 25987 4159
rect 25987 4125 25988 4159
rect 25818 4124 25988 4125
rect 26190 4267 26360 4268
rect 26190 4233 26191 4267
rect 26191 4233 26359 4267
rect 26359 4233 26360 4267
rect 26190 4159 26360 4233
rect 26190 4125 26191 4159
rect 26191 4125 26359 4159
rect 26359 4125 26360 4159
rect 26190 4124 26360 4125
rect 26562 4267 26732 4268
rect 26562 4233 26563 4267
rect 26563 4233 26731 4267
rect 26731 4233 26732 4267
rect 26562 4159 26732 4233
rect 26562 4125 26563 4159
rect 26563 4125 26731 4159
rect 26731 4125 26732 4159
rect 26562 4124 26732 4125
rect 26934 4267 27104 4268
rect 26934 4233 26935 4267
rect 26935 4233 27103 4267
rect 27103 4233 27104 4267
rect 26934 4159 27104 4233
rect 26934 4125 26935 4159
rect 26935 4125 27103 4159
rect 27103 4125 27104 4159
rect 26934 4124 27104 4125
rect 27306 4267 27476 4268
rect 27306 4233 27307 4267
rect 27307 4233 27475 4267
rect 27475 4233 27476 4267
rect 27306 4159 27476 4233
rect 27306 4125 27307 4159
rect 27307 4125 27475 4159
rect 27475 4125 27476 4159
rect 27306 4124 27476 4125
rect 27678 4267 27848 4268
rect 27678 4233 27679 4267
rect 27679 4233 27847 4267
rect 27847 4233 27848 4267
rect 27678 4159 27848 4233
rect 27678 4125 27679 4159
rect 27679 4125 27847 4159
rect 27847 4125 27848 4159
rect 27678 4124 27848 4125
rect 28050 4267 28220 4268
rect 28050 4233 28051 4267
rect 28051 4233 28219 4267
rect 28219 4233 28220 4267
rect 28050 4159 28220 4233
rect 28050 4125 28051 4159
rect 28051 4125 28219 4159
rect 28219 4125 28220 4159
rect 28050 4124 28220 4125
rect 28422 4267 28592 4268
rect 28422 4233 28423 4267
rect 28423 4233 28591 4267
rect 28591 4233 28592 4267
rect 28422 4159 28592 4233
rect 28422 4125 28423 4159
rect 28423 4125 28591 4159
rect 28591 4125 28592 4159
rect 28422 4124 28592 4125
rect 28794 4267 28964 4268
rect 28794 4233 28795 4267
rect 28795 4233 28963 4267
rect 28963 4233 28964 4267
rect 28794 4159 28964 4233
rect 28794 4125 28795 4159
rect 28795 4125 28963 4159
rect 28963 4125 28964 4159
rect 28794 4124 28964 4125
rect 20238 3849 20408 3850
rect 20238 3815 20239 3849
rect 20239 3815 20407 3849
rect 20407 3815 20408 3849
rect 20238 3741 20408 3815
rect 20238 3707 20239 3741
rect 20239 3707 20407 3741
rect 20407 3707 20408 3741
rect 20238 3706 20408 3707
rect 20610 3849 20780 3850
rect 20610 3815 20611 3849
rect 20611 3815 20779 3849
rect 20779 3815 20780 3849
rect 20610 3741 20780 3815
rect 20610 3707 20611 3741
rect 20611 3707 20779 3741
rect 20779 3707 20780 3741
rect 20610 3706 20780 3707
rect 20982 3849 21152 3850
rect 20982 3815 20983 3849
rect 20983 3815 21151 3849
rect 21151 3815 21152 3849
rect 20982 3741 21152 3815
rect 20982 3707 20983 3741
rect 20983 3707 21151 3741
rect 21151 3707 21152 3741
rect 20982 3706 21152 3707
rect 21354 3849 21524 3850
rect 21354 3815 21355 3849
rect 21355 3815 21523 3849
rect 21523 3815 21524 3849
rect 21354 3741 21524 3815
rect 21354 3707 21355 3741
rect 21355 3707 21523 3741
rect 21523 3707 21524 3741
rect 21354 3706 21524 3707
rect 21726 3849 21896 3850
rect 21726 3815 21727 3849
rect 21727 3815 21895 3849
rect 21895 3815 21896 3849
rect 21726 3741 21896 3815
rect 21726 3707 21727 3741
rect 21727 3707 21895 3741
rect 21895 3707 21896 3741
rect 21726 3706 21896 3707
rect 22098 3849 22268 3850
rect 22098 3815 22099 3849
rect 22099 3815 22267 3849
rect 22267 3815 22268 3849
rect 22098 3741 22268 3815
rect 22098 3707 22099 3741
rect 22099 3707 22267 3741
rect 22267 3707 22268 3741
rect 22098 3706 22268 3707
rect 22470 3849 22640 3850
rect 22470 3815 22471 3849
rect 22471 3815 22639 3849
rect 22639 3815 22640 3849
rect 22470 3741 22640 3815
rect 22470 3707 22471 3741
rect 22471 3707 22639 3741
rect 22639 3707 22640 3741
rect 22470 3706 22640 3707
rect 22842 3849 23012 3850
rect 22842 3815 22843 3849
rect 22843 3815 23011 3849
rect 23011 3815 23012 3849
rect 22842 3741 23012 3815
rect 22842 3707 22843 3741
rect 22843 3707 23011 3741
rect 23011 3707 23012 3741
rect 22842 3706 23012 3707
rect 23214 3849 23384 3850
rect 23214 3815 23215 3849
rect 23215 3815 23383 3849
rect 23383 3815 23384 3849
rect 23214 3741 23384 3815
rect 23214 3707 23215 3741
rect 23215 3707 23383 3741
rect 23383 3707 23384 3741
rect 23214 3706 23384 3707
rect 23586 3849 23756 3850
rect 23586 3815 23587 3849
rect 23587 3815 23755 3849
rect 23755 3815 23756 3849
rect 23586 3741 23756 3815
rect 23586 3707 23587 3741
rect 23587 3707 23755 3741
rect 23755 3707 23756 3741
rect 23586 3706 23756 3707
rect 23958 3849 24128 3850
rect 23958 3815 23959 3849
rect 23959 3815 24127 3849
rect 24127 3815 24128 3849
rect 23958 3741 24128 3815
rect 23958 3707 23959 3741
rect 23959 3707 24127 3741
rect 24127 3707 24128 3741
rect 23958 3706 24128 3707
rect 24330 3849 24500 3850
rect 24330 3815 24331 3849
rect 24331 3815 24499 3849
rect 24499 3815 24500 3849
rect 24330 3741 24500 3815
rect 24330 3707 24331 3741
rect 24331 3707 24499 3741
rect 24499 3707 24500 3741
rect 24330 3706 24500 3707
rect 24702 3849 24872 3850
rect 24702 3815 24703 3849
rect 24703 3815 24871 3849
rect 24871 3815 24872 3849
rect 24702 3741 24872 3815
rect 24702 3707 24703 3741
rect 24703 3707 24871 3741
rect 24871 3707 24872 3741
rect 24702 3706 24872 3707
rect 25074 3849 25244 3850
rect 25074 3815 25075 3849
rect 25075 3815 25243 3849
rect 25243 3815 25244 3849
rect 25074 3741 25244 3815
rect 25074 3707 25075 3741
rect 25075 3707 25243 3741
rect 25243 3707 25244 3741
rect 25074 3706 25244 3707
rect 25446 3849 25616 3850
rect 25446 3815 25447 3849
rect 25447 3815 25615 3849
rect 25615 3815 25616 3849
rect 25446 3741 25616 3815
rect 25446 3707 25447 3741
rect 25447 3707 25615 3741
rect 25615 3707 25616 3741
rect 25446 3706 25616 3707
rect 25818 3849 25988 3850
rect 25818 3815 25819 3849
rect 25819 3815 25987 3849
rect 25987 3815 25988 3849
rect 25818 3741 25988 3815
rect 25818 3707 25819 3741
rect 25819 3707 25987 3741
rect 25987 3707 25988 3741
rect 25818 3706 25988 3707
rect 26190 3849 26360 3850
rect 26190 3815 26191 3849
rect 26191 3815 26359 3849
rect 26359 3815 26360 3849
rect 26190 3741 26360 3815
rect 26190 3707 26191 3741
rect 26191 3707 26359 3741
rect 26359 3707 26360 3741
rect 26190 3706 26360 3707
rect 26562 3849 26732 3850
rect 26562 3815 26563 3849
rect 26563 3815 26731 3849
rect 26731 3815 26732 3849
rect 26562 3741 26732 3815
rect 26562 3707 26563 3741
rect 26563 3707 26731 3741
rect 26731 3707 26732 3741
rect 26562 3706 26732 3707
rect 26934 3849 27104 3850
rect 26934 3815 26935 3849
rect 26935 3815 27103 3849
rect 27103 3815 27104 3849
rect 26934 3741 27104 3815
rect 26934 3707 26935 3741
rect 26935 3707 27103 3741
rect 27103 3707 27104 3741
rect 26934 3706 27104 3707
rect 27306 3849 27476 3850
rect 27306 3815 27307 3849
rect 27307 3815 27475 3849
rect 27475 3815 27476 3849
rect 27306 3741 27476 3815
rect 27306 3707 27307 3741
rect 27307 3707 27475 3741
rect 27475 3707 27476 3741
rect 27306 3706 27476 3707
rect 27678 3849 27848 3850
rect 27678 3815 27679 3849
rect 27679 3815 27847 3849
rect 27847 3815 27848 3849
rect 27678 3741 27848 3815
rect 27678 3707 27679 3741
rect 27679 3707 27847 3741
rect 27847 3707 27848 3741
rect 27678 3706 27848 3707
rect 28050 3849 28220 3850
rect 28050 3815 28051 3849
rect 28051 3815 28219 3849
rect 28219 3815 28220 3849
rect 28050 3741 28220 3815
rect 28050 3707 28051 3741
rect 28051 3707 28219 3741
rect 28219 3707 28220 3741
rect 28050 3706 28220 3707
rect 28422 3849 28592 3850
rect 28422 3815 28423 3849
rect 28423 3815 28591 3849
rect 28591 3815 28592 3849
rect 28422 3741 28592 3815
rect 28422 3707 28423 3741
rect 28423 3707 28591 3741
rect 28591 3707 28592 3741
rect 28422 3706 28592 3707
rect 28794 3849 28964 3850
rect 28794 3815 28795 3849
rect 28795 3815 28963 3849
rect 28963 3815 28964 3849
rect 28794 3741 28964 3815
rect 28794 3707 28795 3741
rect 28795 3707 28963 3741
rect 28963 3707 28964 3741
rect 28794 3706 28964 3707
rect 20238 3431 20408 3432
rect 20238 3397 20239 3431
rect 20239 3397 20407 3431
rect 20407 3397 20408 3431
rect 20238 3323 20408 3397
rect 20238 3289 20239 3323
rect 20239 3289 20407 3323
rect 20407 3289 20408 3323
rect 20238 3288 20408 3289
rect 20610 3431 20780 3432
rect 20610 3397 20611 3431
rect 20611 3397 20779 3431
rect 20779 3397 20780 3431
rect 20610 3323 20780 3397
rect 20610 3289 20611 3323
rect 20611 3289 20779 3323
rect 20779 3289 20780 3323
rect 20610 3288 20780 3289
rect 20982 3431 21152 3432
rect 20982 3397 20983 3431
rect 20983 3397 21151 3431
rect 21151 3397 21152 3431
rect 20982 3323 21152 3397
rect 20982 3289 20983 3323
rect 20983 3289 21151 3323
rect 21151 3289 21152 3323
rect 20982 3288 21152 3289
rect 21354 3431 21524 3432
rect 21354 3397 21355 3431
rect 21355 3397 21523 3431
rect 21523 3397 21524 3431
rect 21354 3323 21524 3397
rect 21354 3289 21355 3323
rect 21355 3289 21523 3323
rect 21523 3289 21524 3323
rect 21354 3288 21524 3289
rect 21726 3431 21896 3432
rect 21726 3397 21727 3431
rect 21727 3397 21895 3431
rect 21895 3397 21896 3431
rect 21726 3323 21896 3397
rect 21726 3289 21727 3323
rect 21727 3289 21895 3323
rect 21895 3289 21896 3323
rect 21726 3288 21896 3289
rect 22098 3431 22268 3432
rect 22098 3397 22099 3431
rect 22099 3397 22267 3431
rect 22267 3397 22268 3431
rect 22098 3323 22268 3397
rect 22098 3289 22099 3323
rect 22099 3289 22267 3323
rect 22267 3289 22268 3323
rect 22098 3288 22268 3289
rect 22470 3431 22640 3432
rect 22470 3397 22471 3431
rect 22471 3397 22639 3431
rect 22639 3397 22640 3431
rect 22470 3323 22640 3397
rect 22470 3289 22471 3323
rect 22471 3289 22639 3323
rect 22639 3289 22640 3323
rect 22470 3288 22640 3289
rect 22842 3431 23012 3432
rect 22842 3397 22843 3431
rect 22843 3397 23011 3431
rect 23011 3397 23012 3431
rect 22842 3323 23012 3397
rect 22842 3289 22843 3323
rect 22843 3289 23011 3323
rect 23011 3289 23012 3323
rect 22842 3288 23012 3289
rect 23214 3431 23384 3432
rect 23214 3397 23215 3431
rect 23215 3397 23383 3431
rect 23383 3397 23384 3431
rect 23214 3323 23384 3397
rect 23214 3289 23215 3323
rect 23215 3289 23383 3323
rect 23383 3289 23384 3323
rect 23214 3288 23384 3289
rect 23586 3431 23756 3432
rect 23586 3397 23587 3431
rect 23587 3397 23755 3431
rect 23755 3397 23756 3431
rect 23586 3323 23756 3397
rect 23586 3289 23587 3323
rect 23587 3289 23755 3323
rect 23755 3289 23756 3323
rect 23586 3288 23756 3289
rect 23958 3431 24128 3432
rect 23958 3397 23959 3431
rect 23959 3397 24127 3431
rect 24127 3397 24128 3431
rect 23958 3323 24128 3397
rect 23958 3289 23959 3323
rect 23959 3289 24127 3323
rect 24127 3289 24128 3323
rect 23958 3288 24128 3289
rect 24330 3431 24500 3432
rect 24330 3397 24331 3431
rect 24331 3397 24499 3431
rect 24499 3397 24500 3431
rect 24330 3323 24500 3397
rect 24330 3289 24331 3323
rect 24331 3289 24499 3323
rect 24499 3289 24500 3323
rect 24330 3288 24500 3289
rect 24702 3431 24872 3432
rect 24702 3397 24703 3431
rect 24703 3397 24871 3431
rect 24871 3397 24872 3431
rect 24702 3323 24872 3397
rect 24702 3289 24703 3323
rect 24703 3289 24871 3323
rect 24871 3289 24872 3323
rect 24702 3288 24872 3289
rect 25074 3431 25244 3432
rect 25074 3397 25075 3431
rect 25075 3397 25243 3431
rect 25243 3397 25244 3431
rect 25074 3323 25244 3397
rect 25074 3289 25075 3323
rect 25075 3289 25243 3323
rect 25243 3289 25244 3323
rect 25074 3288 25244 3289
rect 25446 3431 25616 3432
rect 25446 3397 25447 3431
rect 25447 3397 25615 3431
rect 25615 3397 25616 3431
rect 25446 3323 25616 3397
rect 25446 3289 25447 3323
rect 25447 3289 25615 3323
rect 25615 3289 25616 3323
rect 25446 3288 25616 3289
rect 25818 3431 25988 3432
rect 25818 3397 25819 3431
rect 25819 3397 25987 3431
rect 25987 3397 25988 3431
rect 25818 3323 25988 3397
rect 25818 3289 25819 3323
rect 25819 3289 25987 3323
rect 25987 3289 25988 3323
rect 25818 3288 25988 3289
rect 26190 3431 26360 3432
rect 26190 3397 26191 3431
rect 26191 3397 26359 3431
rect 26359 3397 26360 3431
rect 26190 3323 26360 3397
rect 26190 3289 26191 3323
rect 26191 3289 26359 3323
rect 26359 3289 26360 3323
rect 26190 3288 26360 3289
rect 26562 3431 26732 3432
rect 26562 3397 26563 3431
rect 26563 3397 26731 3431
rect 26731 3397 26732 3431
rect 26562 3323 26732 3397
rect 26562 3289 26563 3323
rect 26563 3289 26731 3323
rect 26731 3289 26732 3323
rect 26562 3288 26732 3289
rect 26934 3431 27104 3432
rect 26934 3397 26935 3431
rect 26935 3397 27103 3431
rect 27103 3397 27104 3431
rect 26934 3323 27104 3397
rect 26934 3289 26935 3323
rect 26935 3289 27103 3323
rect 27103 3289 27104 3323
rect 26934 3288 27104 3289
rect 27306 3431 27476 3432
rect 27306 3397 27307 3431
rect 27307 3397 27475 3431
rect 27475 3397 27476 3431
rect 27306 3323 27476 3397
rect 27306 3289 27307 3323
rect 27307 3289 27475 3323
rect 27475 3289 27476 3323
rect 27306 3288 27476 3289
rect 27678 3431 27848 3432
rect 27678 3397 27679 3431
rect 27679 3397 27847 3431
rect 27847 3397 27848 3431
rect 27678 3323 27848 3397
rect 27678 3289 27679 3323
rect 27679 3289 27847 3323
rect 27847 3289 27848 3323
rect 27678 3288 27848 3289
rect 28050 3431 28220 3432
rect 28050 3397 28051 3431
rect 28051 3397 28219 3431
rect 28219 3397 28220 3431
rect 28050 3323 28220 3397
rect 28050 3289 28051 3323
rect 28051 3289 28219 3323
rect 28219 3289 28220 3323
rect 28050 3288 28220 3289
rect 28422 3431 28592 3432
rect 28422 3397 28423 3431
rect 28423 3397 28591 3431
rect 28591 3397 28592 3431
rect 28422 3323 28592 3397
rect 28422 3289 28423 3323
rect 28423 3289 28591 3323
rect 28591 3289 28592 3323
rect 28422 3288 28592 3289
rect 28794 3431 28964 3432
rect 28794 3397 28795 3431
rect 28795 3397 28963 3431
rect 28963 3397 28964 3431
rect 28794 3323 28964 3397
rect 28794 3289 28795 3323
rect 28795 3289 28963 3323
rect 28963 3289 28964 3323
rect 28794 3288 28964 3289
rect 20238 3013 20408 3024
rect 20238 2979 20239 3013
rect 20239 2979 20407 3013
rect 20407 2979 20408 3013
rect 20238 2968 20408 2979
rect 20610 3013 20780 3024
rect 20610 2979 20611 3013
rect 20611 2979 20779 3013
rect 20779 2979 20780 3013
rect 20610 2968 20780 2979
rect 20982 3013 21152 3024
rect 20982 2979 20983 3013
rect 20983 2979 21151 3013
rect 21151 2979 21152 3013
rect 20982 2968 21152 2979
rect 21354 3013 21524 3024
rect 21354 2979 21355 3013
rect 21355 2979 21523 3013
rect 21523 2979 21524 3013
rect 21354 2968 21524 2979
rect 21726 3013 21896 3024
rect 21726 2979 21727 3013
rect 21727 2979 21895 3013
rect 21895 2979 21896 3013
rect 21726 2968 21896 2979
rect 22098 3013 22268 3024
rect 22098 2979 22099 3013
rect 22099 2979 22267 3013
rect 22267 2979 22268 3013
rect 22098 2968 22268 2979
rect 22470 3013 22640 3024
rect 22470 2979 22471 3013
rect 22471 2979 22639 3013
rect 22639 2979 22640 3013
rect 22470 2968 22640 2979
rect 22842 3013 23012 3024
rect 22842 2979 22843 3013
rect 22843 2979 23011 3013
rect 23011 2979 23012 3013
rect 22842 2968 23012 2979
rect 23214 3013 23384 3024
rect 23214 2979 23215 3013
rect 23215 2979 23383 3013
rect 23383 2979 23384 3013
rect 23214 2968 23384 2979
rect 23586 3013 23756 3024
rect 23586 2979 23587 3013
rect 23587 2979 23755 3013
rect 23755 2979 23756 3013
rect 23586 2968 23756 2979
rect 23958 3013 24128 3024
rect 23958 2979 23959 3013
rect 23959 2979 24127 3013
rect 24127 2979 24128 3013
rect 23958 2968 24128 2979
rect 24330 3013 24500 3024
rect 24330 2979 24331 3013
rect 24331 2979 24499 3013
rect 24499 2979 24500 3013
rect 24330 2968 24500 2979
rect 24702 3013 24872 3024
rect 24702 2979 24703 3013
rect 24703 2979 24871 3013
rect 24871 2979 24872 3013
rect 24702 2968 24872 2979
rect 25074 3013 25244 3024
rect 25074 2979 25075 3013
rect 25075 2979 25243 3013
rect 25243 2979 25244 3013
rect 25074 2968 25244 2979
rect 25446 3013 25616 3024
rect 25446 2979 25447 3013
rect 25447 2979 25615 3013
rect 25615 2979 25616 3013
rect 25446 2968 25616 2979
rect 25818 3013 25988 3024
rect 25818 2979 25819 3013
rect 25819 2979 25987 3013
rect 25987 2979 25988 3013
rect 25818 2968 25988 2979
rect 26190 3013 26360 3024
rect 26190 2979 26191 3013
rect 26191 2979 26359 3013
rect 26359 2979 26360 3013
rect 26190 2968 26360 2979
rect 26562 3013 26732 3024
rect 26562 2979 26563 3013
rect 26563 2979 26731 3013
rect 26731 2979 26732 3013
rect 26562 2968 26732 2979
rect 26934 3013 27104 3024
rect 26934 2979 26935 3013
rect 26935 2979 27103 3013
rect 27103 2979 27104 3013
rect 26934 2968 27104 2979
rect 27306 3013 27476 3024
rect 27306 2979 27307 3013
rect 27307 2979 27475 3013
rect 27475 2979 27476 3013
rect 27306 2968 27476 2979
rect 27678 3013 27848 3024
rect 27678 2979 27679 3013
rect 27679 2979 27847 3013
rect 27847 2979 27848 3013
rect 27678 2968 27848 2979
rect 28050 3013 28220 3024
rect 28050 2979 28051 3013
rect 28051 2979 28219 3013
rect 28219 2979 28220 3013
rect 28050 2968 28220 2979
rect 28422 3013 28592 3024
rect 28422 2979 28423 3013
rect 28423 2979 28591 3013
rect 28591 2979 28592 3013
rect 28422 2968 28592 2979
rect 28794 3013 28964 3024
rect 28794 2979 28795 3013
rect 28795 2979 28963 3013
rect 28963 2979 28964 3013
rect 28794 2968 28964 2979
rect 20058 2614 20258 2814
rect 20782 2614 20982 2814
rect 21526 2614 21726 2814
rect 22270 2614 22470 2814
rect 23014 2614 23214 2814
rect 23758 2614 23958 2814
rect 24502 2614 24702 2814
rect 25246 2614 25446 2814
rect 25990 2614 26190 2814
rect 26734 2614 26934 2814
rect 27478 2614 27678 2814
rect 28222 2614 28422 2814
rect 28966 2614 29166 2814
<< metal2 >>
rect 18920 12060 19120 12070
rect 18920 11850 19120 11860
rect 19664 12060 19864 12070
rect 19664 11850 19864 11860
rect 20408 12060 20608 12070
rect 20408 11850 20608 11860
rect 21152 12060 21352 12070
rect 21152 11850 21352 11860
rect 21896 12060 22096 12070
rect 21896 11850 22096 11860
rect 22640 12060 22840 12070
rect 22640 11850 22840 11860
rect 23384 12060 23584 12070
rect 23384 11850 23584 11860
rect 24128 12060 24328 12070
rect 24128 11850 24328 11860
rect 24500 12060 24700 12070
rect 24500 11850 24700 11860
rect 25244 12060 25444 12070
rect 25244 11850 25444 11860
rect 25988 12060 26188 12070
rect 25988 11850 26188 11860
rect 26732 12060 26932 12070
rect 26732 11850 26932 11860
rect 27476 12060 27676 12070
rect 27476 11850 27676 11860
rect 28220 12060 28420 12070
rect 28220 11850 28420 11860
rect 28964 12060 29164 12070
rect 28964 11850 29164 11860
rect 29708 12060 29908 12070
rect 29708 11850 29908 11860
rect 30452 12060 30652 12070
rect 30452 11850 30652 11860
rect 18750 11672 30462 11682
rect 18920 11612 19122 11672
rect 19292 11612 19494 11672
rect 19664 11612 19866 11672
rect 20036 11612 20238 11672
rect 20408 11612 20610 11672
rect 20780 11612 20982 11672
rect 21152 11612 21354 11672
rect 21524 11612 21726 11672
rect 21896 11612 22098 11672
rect 22268 11612 22470 11672
rect 22640 11612 22842 11672
rect 23012 11612 23214 11672
rect 23384 11612 23586 11672
rect 23756 11612 23958 11672
rect 24128 11612 24330 11672
rect 24500 11612 24702 11672
rect 24872 11612 25074 11672
rect 25244 11612 25446 11672
rect 25616 11612 25818 11672
rect 25988 11612 26190 11672
rect 26360 11612 26562 11672
rect 26732 11612 26934 11672
rect 27104 11612 27306 11672
rect 27476 11612 27678 11672
rect 27848 11612 28050 11672
rect 28220 11612 28422 11672
rect 28592 11612 28794 11672
rect 28964 11612 29166 11672
rect 29336 11612 29538 11672
rect 29708 11612 29910 11672
rect 30080 11612 30282 11672
rect 30452 11612 30462 11672
rect 18750 11602 30462 11612
rect 18750 11132 30452 11142
rect 18920 10988 19122 11132
rect 19292 10988 19494 11132
rect 19664 10988 19866 11132
rect 20036 10988 20238 11132
rect 20408 10988 20610 11132
rect 20780 10988 20982 11132
rect 21152 10988 21354 11132
rect 21524 10988 21726 11132
rect 21896 10988 22098 11132
rect 22268 10988 22470 11132
rect 22640 10988 22842 11132
rect 23012 10988 23214 11132
rect 23384 10988 23586 11132
rect 23756 10988 23958 11132
rect 24128 10988 24330 11132
rect 24500 10988 24702 11132
rect 24872 10988 25074 11132
rect 25244 10988 25446 11132
rect 25616 10988 25818 11132
rect 25988 10988 26190 11132
rect 26360 10988 26562 11132
rect 26732 10988 26934 11132
rect 27104 10988 27306 11132
rect 27476 10988 27678 11132
rect 27848 10988 28050 11132
rect 28220 10988 28422 11132
rect 28592 10988 28794 11132
rect 28964 10988 29166 11132
rect 29336 10988 29538 11132
rect 29708 10988 29910 11132
rect 30080 10988 30282 11132
rect 18750 10978 30452 10988
rect 18750 10496 30452 10506
rect 18920 10352 19122 10496
rect 19292 10352 19494 10496
rect 19664 10352 19866 10496
rect 20036 10352 20238 10496
rect 20408 10352 20610 10496
rect 20780 10352 20982 10496
rect 21152 10352 21354 10496
rect 21524 10352 21726 10496
rect 21896 10352 22098 10496
rect 22268 10352 22470 10496
rect 22640 10352 22842 10496
rect 23012 10352 23214 10496
rect 23384 10352 23586 10496
rect 23756 10352 23958 10496
rect 24128 10352 24330 10496
rect 24500 10352 24702 10496
rect 24872 10352 25074 10496
rect 25244 10352 25446 10496
rect 25616 10352 25818 10496
rect 25988 10352 26190 10496
rect 26360 10352 26562 10496
rect 26732 10352 26934 10496
rect 27104 10352 27306 10496
rect 27476 10352 27678 10496
rect 27848 10352 28050 10496
rect 28220 10352 28422 10496
rect 28592 10352 28794 10496
rect 28964 10352 29166 10496
rect 29336 10352 29538 10496
rect 29708 10352 29910 10496
rect 30080 10352 30282 10496
rect 18750 10342 30452 10352
rect 18750 9872 30452 9882
rect 18920 9812 19122 9872
rect 19292 9812 19494 9872
rect 19664 9812 19866 9872
rect 20036 9812 20238 9872
rect 20408 9812 20610 9872
rect 20780 9812 20982 9872
rect 21152 9812 21354 9872
rect 21524 9812 21726 9872
rect 21896 9812 22098 9872
rect 22268 9812 22470 9872
rect 22640 9812 22842 9872
rect 23012 9812 23214 9872
rect 23384 9812 23586 9872
rect 23756 9812 23958 9872
rect 24128 9812 24330 9872
rect 24500 9812 24702 9872
rect 24872 9812 25074 9872
rect 25244 9812 25446 9872
rect 25616 9812 25818 9872
rect 25988 9812 26190 9872
rect 26360 9812 26562 9872
rect 26732 9812 26934 9872
rect 27104 9812 27306 9872
rect 27476 9812 27678 9872
rect 27848 9812 28050 9872
rect 28220 9812 28422 9872
rect 28592 9812 28794 9872
rect 28964 9812 29166 9872
rect 29336 9812 29538 9872
rect 29708 9812 29910 9872
rect 30080 9812 30282 9872
rect 18750 9802 30452 9812
rect 24834 9504 30324 9514
rect 19758 9386 22826 9484
rect 20424 9296 20594 9386
rect 22656 9296 22826 9386
rect 20238 9286 20780 9296
rect 20408 9222 20610 9286
rect 20238 9212 20780 9222
rect 20982 9286 22268 9296
rect 21152 9222 21354 9286
rect 21524 9222 21726 9286
rect 21896 9222 22098 9286
rect 20982 9212 22268 9222
rect 22470 9286 23012 9296
rect 22640 9222 22842 9286
rect 25116 9232 25578 9504
rect 25860 9232 26322 9504
rect 26604 9232 27066 9504
rect 27348 9232 27810 9504
rect 28092 9232 28554 9504
rect 28836 9232 29298 9504
rect 29580 9232 30042 9504
rect 24834 9222 30324 9232
rect 22470 9212 23012 9222
rect 20482 8354 20536 9212
rect 21226 8354 21280 9212
rect 21970 8354 22024 9212
rect 22714 8354 22768 9212
rect 20238 8344 20780 8354
rect 20408 8200 20610 8344
rect 20238 8190 20780 8200
rect 20982 8344 22268 8354
rect 21152 8200 21354 8344
rect 21524 8200 21726 8344
rect 21896 8200 22098 8344
rect 20982 8190 22268 8200
rect 22470 8344 23012 8354
rect 22640 8200 22842 8344
rect 22470 8190 23012 8200
rect 20482 7318 20536 8190
rect 21226 7318 21280 8190
rect 21970 7318 22024 8190
rect 22714 7318 22768 8190
rect 23716 7788 23998 7798
rect 23716 7506 23998 7516
rect 20238 7308 20780 7318
rect 20408 7164 20610 7308
rect 20238 7154 20780 7164
rect 20982 7308 22268 7318
rect 21152 7164 21354 7308
rect 21524 7164 21726 7308
rect 21896 7164 22098 7308
rect 20982 7154 22268 7164
rect 22470 7308 23012 7318
rect 22640 7164 22842 7308
rect 22470 7154 23012 7164
rect 20482 6282 20536 7154
rect 21226 6282 21280 7154
rect 21970 6282 22024 7154
rect 22714 6282 22768 7154
rect 24132 6886 24330 6896
rect 24132 6678 24330 6688
rect 24132 6486 24330 6496
rect 20238 6272 20780 6282
rect 20408 6128 20610 6272
rect 20238 6118 20780 6128
rect 20982 6272 22268 6282
rect 21152 6128 21354 6272
rect 21524 6128 21726 6272
rect 21896 6128 22098 6272
rect 20982 6118 22268 6128
rect 22470 6272 23012 6282
rect 24132 6278 24330 6288
rect 22640 6128 22842 6272
rect 22470 6118 23012 6128
rect 20482 5256 20536 6118
rect 21226 5256 21280 6118
rect 21970 5256 22024 6118
rect 22714 5256 22768 6118
rect 24132 6086 24330 6096
rect 24132 5878 24330 5888
rect 23344 5322 28844 5332
rect 20238 5246 20780 5256
rect 20408 5192 20610 5246
rect 20238 5182 20780 5192
rect 20982 5246 22268 5256
rect 21152 5192 21354 5246
rect 21524 5192 21726 5246
rect 21896 5192 22098 5246
rect 20982 5182 22268 5192
rect 22470 5246 23012 5256
rect 22640 5192 22842 5246
rect 22470 5182 23012 5192
rect 21168 5082 21338 5182
rect 21912 5082 22082 5182
rect 19758 4984 22082 5082
rect 23626 5158 24088 5322
rect 23344 5040 23626 5050
rect 24370 5158 24832 5322
rect 24088 5040 24370 5050
rect 25114 5158 25576 5322
rect 24832 5040 25114 5050
rect 25858 5158 26320 5322
rect 25576 5040 25858 5050
rect 26602 5158 27064 5322
rect 26320 5040 26602 5050
rect 27346 5158 27808 5322
rect 27064 5040 27346 5050
rect 28090 5158 28552 5322
rect 27808 5040 28090 5050
rect 28834 5158 28844 5322
rect 28552 5040 28834 5050
rect 23724 4976 23974 4986
rect 21218 4906 23724 4916
rect 22032 4772 23724 4906
rect 22032 4726 23198 4772
rect 21218 4716 23198 4726
rect 23724 4716 23974 4726
rect 23072 4598 23198 4716
rect 20238 4588 23024 4598
rect 20408 4532 20610 4588
rect 20780 4532 20982 4588
rect 21152 4532 21354 4588
rect 21524 4532 21726 4588
rect 21896 4532 22098 4588
rect 22268 4532 22470 4588
rect 22640 4532 22842 4588
rect 23012 4532 23024 4588
rect 20238 4522 23024 4532
rect 23072 4588 28964 4598
rect 23072 4532 23214 4588
rect 23384 4532 23586 4588
rect 23756 4532 23958 4588
rect 24128 4532 24330 4588
rect 24500 4532 24702 4588
rect 24872 4532 25074 4588
rect 25244 4532 25446 4588
rect 25616 4532 25818 4588
rect 25988 4532 26190 4588
rect 26360 4532 26562 4588
rect 26732 4532 26934 4588
rect 27104 4532 27306 4588
rect 27476 4532 27678 4588
rect 27848 4532 28050 4588
rect 28220 4532 28422 4588
rect 28592 4532 28794 4588
rect 23072 4522 28964 4532
rect 23072 4278 23198 4522
rect 20238 4268 23024 4278
rect 20408 4124 20610 4268
rect 20780 4124 20982 4268
rect 21152 4124 21354 4268
rect 21524 4124 21726 4268
rect 21896 4124 22098 4268
rect 22268 4124 22470 4268
rect 22640 4124 22842 4268
rect 23012 4124 23024 4268
rect 20238 4114 23024 4124
rect 23072 4268 28964 4278
rect 23072 4124 23214 4268
rect 23384 4124 23586 4268
rect 23756 4124 23958 4268
rect 24128 4124 24330 4268
rect 24500 4124 24702 4268
rect 24872 4124 25074 4268
rect 25244 4124 25446 4268
rect 25616 4124 25818 4268
rect 25988 4124 26190 4268
rect 26360 4124 26562 4268
rect 26732 4124 26934 4268
rect 27104 4124 27306 4268
rect 27476 4124 27678 4268
rect 27848 4124 28050 4268
rect 28220 4124 28422 4268
rect 28592 4124 28794 4268
rect 23072 4114 28964 4124
rect 23072 3860 23198 4114
rect 20238 3850 23024 3860
rect 20408 3706 20610 3850
rect 20780 3706 20982 3850
rect 21152 3706 21354 3850
rect 21524 3706 21726 3850
rect 21896 3706 22098 3850
rect 22268 3706 22470 3850
rect 22640 3706 22842 3850
rect 23012 3706 23024 3850
rect 20238 3696 23024 3706
rect 23072 3850 28964 3860
rect 23072 3706 23214 3850
rect 23384 3706 23586 3850
rect 23756 3706 23958 3850
rect 24128 3706 24330 3850
rect 24500 3706 24702 3850
rect 24872 3706 25074 3850
rect 25244 3706 25446 3850
rect 25616 3706 25818 3850
rect 25988 3706 26190 3850
rect 26360 3706 26562 3850
rect 26732 3706 26934 3850
rect 27104 3706 27306 3850
rect 27476 3706 27678 3850
rect 27848 3706 28050 3850
rect 28220 3706 28422 3850
rect 28592 3706 28794 3850
rect 23072 3696 28964 3706
rect 23072 3442 23198 3696
rect 20238 3432 23024 3442
rect 20408 3288 20610 3432
rect 20780 3288 20982 3432
rect 21152 3288 21354 3432
rect 21524 3288 21726 3432
rect 21896 3288 22098 3432
rect 22268 3288 22470 3432
rect 22640 3288 22842 3432
rect 23012 3288 23024 3432
rect 20238 3278 23024 3288
rect 23072 3432 28964 3442
rect 23072 3288 23214 3432
rect 23384 3288 23586 3432
rect 23756 3288 23958 3432
rect 24128 3288 24330 3432
rect 24500 3288 24702 3432
rect 24872 3288 25074 3432
rect 25244 3288 25446 3432
rect 25616 3288 25818 3432
rect 25988 3288 26190 3432
rect 26360 3288 26562 3432
rect 26732 3288 26934 3432
rect 27104 3288 27306 3432
rect 27476 3288 27678 3432
rect 27848 3288 28050 3432
rect 28220 3288 28422 3432
rect 28592 3288 28794 3432
rect 23072 3278 28964 3288
rect 23072 3034 23198 3278
rect 20238 3024 23024 3034
rect 20408 2968 20610 3024
rect 20780 2968 20982 3024
rect 21152 2968 21354 3024
rect 21524 2968 21726 3024
rect 21896 2968 22098 3024
rect 22268 2968 22470 3024
rect 22640 2968 22842 3024
rect 23012 2968 23024 3024
rect 20238 2958 23024 2968
rect 23072 3024 28964 3034
rect 23072 2968 23214 3024
rect 23384 2968 23586 3024
rect 23756 2968 23958 3024
rect 24128 2968 24330 3024
rect 24500 2968 24702 3024
rect 24872 2968 25074 3024
rect 25244 2968 25446 3024
rect 25616 2968 25818 3024
rect 25988 2968 26190 3024
rect 26360 2968 26562 3024
rect 26732 2968 26934 3024
rect 27104 2968 27306 3024
rect 27476 2968 27678 3024
rect 27848 2968 28050 3024
rect 28220 2968 28422 3024
rect 28592 2968 28794 3024
rect 23072 2958 28964 2968
rect 20058 2814 20258 2824
rect 20058 2604 20258 2614
rect 20782 2814 20982 2824
rect 20782 2604 20982 2614
rect 21526 2814 21726 2824
rect 21526 2604 21726 2614
rect 22270 2814 22470 2824
rect 22270 2604 22470 2614
rect 23014 2814 23214 2824
rect 23014 2604 23214 2614
rect 23758 2814 23958 2824
rect 23758 2604 23958 2614
rect 24502 2814 24702 2824
rect 24502 2604 24702 2614
rect 25246 2814 25446 2824
rect 25246 2604 25446 2614
rect 25990 2814 26190 2824
rect 25990 2604 26190 2614
rect 26734 2814 26934 2824
rect 26734 2604 26934 2614
rect 27478 2814 27678 2824
rect 27478 2604 27678 2614
rect 28222 2814 28422 2824
rect 28222 2604 28422 2614
rect 28966 2814 29166 2824
rect 28966 2604 29166 2614
<< via2 >>
rect 18920 11860 19120 12060
rect 19664 11860 19864 12060
rect 20408 11860 20608 12060
rect 21152 11860 21352 12060
rect 21896 11860 22096 12060
rect 22640 11860 22840 12060
rect 23384 11860 23584 12060
rect 24128 11860 24328 12060
rect 24500 11860 24700 12060
rect 25244 11860 25444 12060
rect 25988 11860 26188 12060
rect 26732 11860 26932 12060
rect 27476 11860 27676 12060
rect 28220 11860 28420 12060
rect 28964 11860 29164 12060
rect 29708 11860 29908 12060
rect 30452 11860 30652 12060
rect 26322 9232 26604 9504
rect 27066 9232 27348 9504
rect 27810 9232 28092 9504
rect 28554 9232 28836 9504
rect 23716 7516 23998 7788
rect 24132 6688 24330 6886
rect 24132 6288 24330 6486
rect 24132 5888 24330 6086
rect 26320 5050 26602 5322
rect 27064 5050 27346 5322
rect 27808 5050 28090 5322
rect 28552 5050 28834 5322
rect 20058 2614 20258 2814
rect 20782 2614 20982 2814
rect 21526 2614 21726 2814
rect 22270 2614 22470 2814
rect 23014 2614 23214 2814
rect 23758 2614 23958 2814
rect 24502 2614 24702 2814
rect 25246 2614 25446 2814
rect 25990 2614 26190 2814
rect 26734 2614 26934 2814
rect 27478 2614 27678 2814
rect 28222 2614 28422 2814
rect 28966 2614 29166 2814
<< metal3 >>
rect 18910 12060 19130 12065
rect 18910 11860 18920 12060
rect 19120 11860 19130 12060
rect 18910 11855 19130 11860
rect 19654 12060 19874 12065
rect 19654 11860 19664 12060
rect 19864 11860 19874 12060
rect 19654 11855 19874 11860
rect 20398 12060 20618 12065
rect 20398 11860 20408 12060
rect 20608 11860 20618 12060
rect 20398 11855 20618 11860
rect 21142 12060 21362 12065
rect 21142 11860 21152 12060
rect 21352 11860 21362 12060
rect 21142 11855 21362 11860
rect 21886 12060 22106 12065
rect 21886 11860 21896 12060
rect 22096 11860 22106 12060
rect 21886 11855 22106 11860
rect 22630 12060 22850 12065
rect 22630 11860 22640 12060
rect 22840 11860 22850 12060
rect 22630 11855 22850 11860
rect 23374 12060 23594 12065
rect 23374 11860 23384 12060
rect 23584 11860 23594 12060
rect 23374 11855 23594 11860
rect 24118 12060 24338 12065
rect 24118 11860 24128 12060
rect 24328 11860 24338 12060
rect 24118 11855 24338 11860
rect 24490 12060 24710 12065
rect 24490 11860 24500 12060
rect 24700 11860 24710 12060
rect 24490 11855 24710 11860
rect 25234 12060 25454 12065
rect 25234 11860 25244 12060
rect 25444 11860 25454 12060
rect 25234 11855 25454 11860
rect 25978 12060 26198 12065
rect 25978 11860 25988 12060
rect 26188 11860 26198 12060
rect 25978 11855 26198 11860
rect 26722 12060 26942 12065
rect 26722 11860 26732 12060
rect 26932 11860 26942 12060
rect 26722 11855 26942 11860
rect 27466 12060 27686 12065
rect 27466 11860 27476 12060
rect 27676 11860 27686 12060
rect 27466 11855 27686 11860
rect 28210 12060 28430 12065
rect 28210 11860 28220 12060
rect 28420 11860 28430 12060
rect 28210 11855 28430 11860
rect 28954 12060 29174 12065
rect 28954 11860 28964 12060
rect 29164 11860 29174 12060
rect 28954 11855 29174 11860
rect 29698 12060 29918 12065
rect 29698 11860 29708 12060
rect 29908 11860 29918 12060
rect 29698 11855 29918 11860
rect 30442 12060 30662 12065
rect 30442 11860 30452 12060
rect 30652 11860 30662 12060
rect 30442 11855 30662 11860
rect 26312 9504 26614 9509
rect 26312 9232 26322 9504
rect 26604 9232 26614 9504
rect 26312 9026 26614 9232
rect 27056 9504 27358 9509
rect 27056 9232 27066 9504
rect 27348 9232 27358 9504
rect 27056 9026 27358 9232
rect 27800 9504 28102 9509
rect 27800 9232 27810 9504
rect 28092 9232 28102 9504
rect 27800 9026 28102 9232
rect 28544 9504 28846 9509
rect 28544 9232 28554 9504
rect 28836 9232 28846 9504
rect 28544 9026 28846 9232
rect 30712 9026 33688 9538
rect 23706 7788 24008 7793
rect 23706 7516 23716 7788
rect 23998 7516 24008 7788
rect 23706 7511 24008 7516
rect 24482 7050 33688 9026
rect 24122 6886 24340 6891
rect 24122 6688 24132 6886
rect 24330 6688 24340 6886
rect 24122 6683 24340 6688
rect 24482 6564 34162 7050
rect 24122 6486 24340 6491
rect 24122 6288 24132 6486
rect 24330 6288 24340 6486
rect 24122 6283 24340 6288
rect 24122 6086 24340 6091
rect 24122 5888 24132 6086
rect 24330 5888 24340 6086
rect 24482 6026 33688 6564
rect 24122 5883 24340 5888
rect 26310 5322 26612 6026
rect 26310 5050 26320 5322
rect 26602 5050 26612 5322
rect 26310 5045 26612 5050
rect 27054 5322 27356 6026
rect 27054 5050 27064 5322
rect 27346 5050 27356 5322
rect 27054 5045 27356 5050
rect 27798 5322 28100 6026
rect 27798 5050 27808 5322
rect 28090 5050 28100 5322
rect 27798 5045 28100 5050
rect 28542 5322 28844 6026
rect 28542 5050 28552 5322
rect 28834 5050 28844 5322
rect 28542 5045 28844 5050
rect 30712 3338 33688 6026
rect 20048 2814 20268 2819
rect 20048 2614 20058 2814
rect 20258 2614 20268 2814
rect 20048 2609 20268 2614
rect 20772 2814 20992 2819
rect 20772 2614 20782 2814
rect 20982 2614 20992 2814
rect 20772 2609 20992 2614
rect 21516 2814 21736 2819
rect 21516 2614 21526 2814
rect 21726 2614 21736 2814
rect 21516 2609 21736 2614
rect 22260 2814 22480 2819
rect 22260 2614 22270 2814
rect 22470 2614 22480 2814
rect 22260 2609 22480 2614
rect 23004 2814 23224 2819
rect 23004 2614 23014 2814
rect 23214 2614 23224 2814
rect 23004 2609 23224 2614
rect 23748 2814 23968 2819
rect 23748 2614 23758 2814
rect 23958 2614 23968 2814
rect 23748 2609 23968 2614
rect 24492 2814 24712 2819
rect 24492 2614 24502 2814
rect 24702 2614 24712 2814
rect 24492 2609 24712 2614
rect 25236 2814 25456 2819
rect 25236 2614 25246 2814
rect 25446 2614 25456 2814
rect 25236 2609 25456 2614
rect 25980 2814 26200 2819
rect 25980 2614 25990 2814
rect 26190 2614 26200 2814
rect 25980 2609 26200 2614
rect 26724 2814 26944 2819
rect 26724 2614 26734 2814
rect 26934 2614 26944 2814
rect 26724 2609 26944 2614
rect 27468 2814 27688 2819
rect 27468 2614 27478 2814
rect 27678 2614 27688 2814
rect 27468 2609 27688 2614
rect 28212 2814 28432 2819
rect 28212 2614 28222 2814
rect 28422 2614 28432 2814
rect 28212 2609 28432 2614
rect 28956 2814 29176 2819
rect 28956 2614 28966 2814
rect 29166 2614 29176 2814
rect 28956 2609 29176 2614
<< via3 >>
rect 18920 11860 19120 12060
rect 19664 11860 19864 12060
rect 20408 11860 20608 12060
rect 21152 11860 21352 12060
rect 21896 11860 22096 12060
rect 22640 11860 22840 12060
rect 23384 11860 23584 12060
rect 24128 11860 24328 12060
rect 24500 11860 24700 12060
rect 25244 11860 25444 12060
rect 25988 11860 26188 12060
rect 26732 11860 26932 12060
rect 27476 11860 27676 12060
rect 28220 11860 28420 12060
rect 28964 11860 29164 12060
rect 29708 11860 29908 12060
rect 30452 11860 30652 12060
rect 23716 7516 23998 7788
rect 24132 6688 24330 6886
rect 24132 6288 24330 6486
rect 24132 5888 24330 6086
rect 20058 2614 20258 2814
rect 20782 2614 20982 2814
rect 21526 2614 21726 2814
rect 22270 2614 22470 2814
rect 23014 2614 23214 2814
rect 23758 2614 23958 2814
rect 24502 2614 24702 2814
rect 25246 2614 25446 2814
rect 25990 2614 26190 2814
rect 26734 2614 26934 2814
rect 27478 2614 27678 2814
rect 28222 2614 28422 2814
rect 28966 2614 29166 2814
<< mimcap >>
rect 30812 9398 33612 9438
rect 24582 8886 30582 8926
rect 24582 6166 24622 8886
rect 30542 6166 30582 8886
rect 24582 6126 30582 6166
rect 30812 3478 30852 9398
rect 33572 3478 33612 9398
rect 30812 3438 33612 3478
<< mimcapcontact >>
rect 24622 6166 30542 8886
rect 30852 3478 33572 9398
<< metal4 >>
rect 18314 12060 30838 12838
rect 18314 11860 18920 12060
rect 19120 11860 19664 12060
rect 19864 11860 20408 12060
rect 20608 11860 21152 12060
rect 21352 11860 21896 12060
rect 22096 11860 22640 12060
rect 22840 11860 23384 12060
rect 23584 11860 24128 12060
rect 24328 11860 24500 12060
rect 24700 11860 25244 12060
rect 25444 11860 25988 12060
rect 26188 11860 26732 12060
rect 26932 11860 27476 12060
rect 27676 11860 28220 12060
rect 28420 11860 28964 12060
rect 29164 11860 29708 12060
rect 29908 11860 30452 12060
rect 30652 11860 30838 12060
rect 18314 11834 30838 11860
rect 30851 9398 33573 9399
rect 30851 8888 30852 9398
rect 30496 8887 30852 8888
rect 24621 8886 30852 8887
rect 23715 7788 23999 7789
rect 23715 7516 23716 7788
rect 23998 7760 23999 7788
rect 24621 7760 24622 8886
rect 23998 7542 24622 7760
rect 23998 7516 23999 7542
rect 23715 7515 23999 7516
rect 24104 6886 24364 6914
rect 24104 6688 24132 6886
rect 24330 6688 24364 6886
rect 24104 6486 24364 6688
rect 24104 6288 24132 6486
rect 24330 6288 24364 6486
rect 24104 6086 24364 6288
rect 24621 6166 24622 7542
rect 30542 6166 30852 8886
rect 24621 6165 30852 6166
rect 30496 6164 30852 6165
rect 24104 5888 24132 6086
rect 24330 5888 24364 6086
rect 24104 2838 24364 5888
rect 30851 3478 30852 6164
rect 33572 3478 33573 9398
rect 30851 3477 33573 3478
rect 18314 2814 30838 2838
rect 18314 2614 20058 2814
rect 20258 2614 20782 2814
rect 20982 2614 21526 2814
rect 21726 2614 22270 2814
rect 22470 2614 23014 2814
rect 23214 2614 23758 2814
rect 23958 2614 24502 2814
rect 24702 2614 25246 2814
rect 25446 2614 25990 2814
rect 26190 2614 26734 2814
rect 26934 2614 27478 2814
rect 27678 2614 28222 2814
rect 28422 2614 28966 2814
rect 29166 2614 30838 2814
rect 18314 1834 30838 2614
<< labels >>
flabel metal4 19510 12512 19510 12512 0 FreeSans 8000 0 0 0 vdd
port 0 nsew
flabel metal4 19076 1998 19076 1998 0 FreeSans 8000 0 0 0 vss
port 4 nsew
flabel metal2 19788 9416 19788 9416 0 FreeSans 8000 0 0 0 vn
port 2 nsew
flabel metal2 19824 5016 19824 5016 0 FreeSans 8000 0 0 0 vp
port 1 nsew
flabel metal1 18700 10416 18700 10416 0 FreeSans 8000 0 0 0 vbias
port 3 nsew
flabel metal3 33908 6768 33908 6768 0 FreeSans 8000 0 0 0 vout
port 5 nsew
<< end >>
